module tt_um_Coline3003_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire clknet_0_clk;
 wire \top1.FSM1.SL ;
 wire \top1.FSM1.counter_register[0] ;
 wire \top1.FSM1.counter_register[1] ;
 wire \top1.FSM1.counter_register[2] ;
 wire \top1.FSM1.counter_register[3] ;
 wire \top1.FSM1.ovf ;
 wire \top1.FSM1.state_next[0] ;
 wire \top1.FSM1.state_next[1] ;
 wire \top1.FSM1.state_next[2] ;
 wire \top1.FSM1.state_next[3] ;
 wire \top1.FSM1.state_next[4] ;
 wire \top1.FSM1.state_reg[0] ;
 wire \top1.FSM1.state_reg[1] ;
 wire \top1.FSM1.state_reg[2] ;
 wire \top1.FSM1.state_reg[3] ;
 wire \top1.FSM1.state_reg[4] ;
 wire \top1.PISO_register1.register[0] ;
 wire \top1.PISO_register1.register[10] ;
 wire \top1.PISO_register1.register[1] ;
 wire \top1.PISO_register1.register[2] ;
 wire \top1.PISO_register1.register[3] ;
 wire \top1.PISO_register1.register[4] ;
 wire \top1.PISO_register1.register[5] ;
 wire \top1.PISO_register1.register[6] ;
 wire \top1.PISO_register1.register[7] ;
 wire \top1.PISO_register1.register[8] ;
 wire \top1.PISO_register1.register[9] ;
 wire \top1.PISO_register1.serial_out ;
 wire \top1.a0_out ;
 wire \top1.a1_out ;
 wire \top1.a2_out ;
 wire \top1.a3_out ;
 wire \top1.ch10c.data[0] ;
 wire \top1.ch10c.data[10] ;
 wire \top1.ch10c.data[11] ;
 wire \top1.ch10c.data[1] ;
 wire \top1.ch10c.data[2] ;
 wire \top1.ch10c.data[3] ;
 wire \top1.ch10c.data[4] ;
 wire \top1.ch10c.data[5] ;
 wire \top1.ch10c.data[6] ;
 wire \top1.ch10c.data[7] ;
 wire \top1.ch10c.data[8] ;
 wire \top1.ch10c.data[9] ;
 wire \top1.ch10c.ovf ;
 wire \top1.ch11c.data[0] ;
 wire \top1.ch11c.data[10] ;
 wire \top1.ch11c.data[11] ;
 wire \top1.ch11c.data[1] ;
 wire \top1.ch11c.data[2] ;
 wire \top1.ch11c.data[3] ;
 wire \top1.ch11c.data[4] ;
 wire \top1.ch11c.data[5] ;
 wire \top1.ch11c.data[6] ;
 wire \top1.ch11c.data[7] ;
 wire \top1.ch11c.data[8] ;
 wire \top1.ch11c.data[9] ;
 wire \top1.ch11c.ovf ;
 wire \top1.ch12c.data[0] ;
 wire \top1.ch12c.data[10] ;
 wire \top1.ch12c.data[11] ;
 wire \top1.ch12c.data[1] ;
 wire \top1.ch12c.data[2] ;
 wire \top1.ch12c.data[3] ;
 wire \top1.ch12c.data[4] ;
 wire \top1.ch12c.data[5] ;
 wire \top1.ch12c.data[6] ;
 wire \top1.ch12c.data[7] ;
 wire \top1.ch12c.data[8] ;
 wire \top1.ch12c.data[9] ;
 wire \top1.ch12c.ovf ;
 wire \top1.ch13c.data[0] ;
 wire \top1.ch13c.data[10] ;
 wire \top1.ch13c.data[11] ;
 wire \top1.ch13c.data[1] ;
 wire \top1.ch13c.data[2] ;
 wire \top1.ch13c.data[3] ;
 wire \top1.ch13c.data[4] ;
 wire \top1.ch13c.data[5] ;
 wire \top1.ch13c.data[6] ;
 wire \top1.ch13c.data[7] ;
 wire \top1.ch13c.data[8] ;
 wire \top1.ch13c.data[9] ;
 wire \top1.ch13c.ovf ;
 wire \top1.ch14c.data[0] ;
 wire \top1.ch14c.data[10] ;
 wire \top1.ch14c.data[11] ;
 wire \top1.ch14c.data[1] ;
 wire \top1.ch14c.data[2] ;
 wire \top1.ch14c.data[3] ;
 wire \top1.ch14c.data[4] ;
 wire \top1.ch14c.data[5] ;
 wire \top1.ch14c.data[6] ;
 wire \top1.ch14c.data[7] ;
 wire \top1.ch14c.data[8] ;
 wire \top1.ch14c.data[9] ;
 wire \top1.ch14c.ovf ;
 wire \top1.ch15c.data[0] ;
 wire \top1.ch15c.data[10] ;
 wire \top1.ch15c.data[11] ;
 wire \top1.ch15c.data[1] ;
 wire \top1.ch15c.data[2] ;
 wire \top1.ch15c.data[3] ;
 wire \top1.ch15c.data[4] ;
 wire \top1.ch15c.data[5] ;
 wire \top1.ch15c.data[6] ;
 wire \top1.ch15c.data[7] ;
 wire \top1.ch15c.data[8] ;
 wire \top1.ch15c.data[9] ;
 wire \top1.ch15c.ovf ;
 wire \top1.ch1c.data[0] ;
 wire \top1.ch1c.data[10] ;
 wire \top1.ch1c.data[11] ;
 wire \top1.ch1c.data[1] ;
 wire \top1.ch1c.data[2] ;
 wire \top1.ch1c.data[3] ;
 wire \top1.ch1c.data[4] ;
 wire \top1.ch1c.data[5] ;
 wire \top1.ch1c.data[6] ;
 wire \top1.ch1c.data[7] ;
 wire \top1.ch1c.data[8] ;
 wire \top1.ch1c.data[9] ;
 wire \top1.ch1c.ovf ;
 wire \top1.ch2c.data[0] ;
 wire \top1.ch2c.data[10] ;
 wire \top1.ch2c.data[11] ;
 wire \top1.ch2c.data[1] ;
 wire \top1.ch2c.data[2] ;
 wire \top1.ch2c.data[3] ;
 wire \top1.ch2c.data[4] ;
 wire \top1.ch2c.data[5] ;
 wire \top1.ch2c.data[6] ;
 wire \top1.ch2c.data[7] ;
 wire \top1.ch2c.data[8] ;
 wire \top1.ch2c.data[9] ;
 wire \top1.ch2c.ovf ;
 wire \top1.ch3c.data[0] ;
 wire \top1.ch3c.data[10] ;
 wire \top1.ch3c.data[11] ;
 wire \top1.ch3c.data[1] ;
 wire \top1.ch3c.data[2] ;
 wire \top1.ch3c.data[3] ;
 wire \top1.ch3c.data[4] ;
 wire \top1.ch3c.data[5] ;
 wire \top1.ch3c.data[6] ;
 wire \top1.ch3c.data[7] ;
 wire \top1.ch3c.data[8] ;
 wire \top1.ch3c.data[9] ;
 wire \top1.ch3c.ovf ;
 wire \top1.ch4c.data[0] ;
 wire \top1.ch4c.data[10] ;
 wire \top1.ch4c.data[11] ;
 wire \top1.ch4c.data[1] ;
 wire \top1.ch4c.data[2] ;
 wire \top1.ch4c.data[3] ;
 wire \top1.ch4c.data[4] ;
 wire \top1.ch4c.data[5] ;
 wire \top1.ch4c.data[6] ;
 wire \top1.ch4c.data[7] ;
 wire \top1.ch4c.data[8] ;
 wire \top1.ch4c.data[9] ;
 wire \top1.ch4c.ovf ;
 wire \top1.ch5c.data[0] ;
 wire \top1.ch5c.data[10] ;
 wire \top1.ch5c.data[11] ;
 wire \top1.ch5c.data[1] ;
 wire \top1.ch5c.data[2] ;
 wire \top1.ch5c.data[3] ;
 wire \top1.ch5c.data[4] ;
 wire \top1.ch5c.data[5] ;
 wire \top1.ch5c.data[6] ;
 wire \top1.ch5c.data[7] ;
 wire \top1.ch5c.data[8] ;
 wire \top1.ch5c.data[9] ;
 wire \top1.ch5c.ovf ;
 wire \top1.ch6c.data[0] ;
 wire \top1.ch6c.data[10] ;
 wire \top1.ch6c.data[11] ;
 wire \top1.ch6c.data[1] ;
 wire \top1.ch6c.data[2] ;
 wire \top1.ch6c.data[3] ;
 wire \top1.ch6c.data[4] ;
 wire \top1.ch6c.data[5] ;
 wire \top1.ch6c.data[6] ;
 wire \top1.ch6c.data[7] ;
 wire \top1.ch6c.data[8] ;
 wire \top1.ch6c.data[9] ;
 wire \top1.ch6c.ovf ;
 wire \top1.ch7c.data[0] ;
 wire \top1.ch7c.data[10] ;
 wire \top1.ch7c.data[11] ;
 wire \top1.ch7c.data[1] ;
 wire \top1.ch7c.data[2] ;
 wire \top1.ch7c.data[3] ;
 wire \top1.ch7c.data[4] ;
 wire \top1.ch7c.data[5] ;
 wire \top1.ch7c.data[6] ;
 wire \top1.ch7c.data[7] ;
 wire \top1.ch7c.data[8] ;
 wire \top1.ch7c.data[9] ;
 wire \top1.ch7c.ovf ;
 wire \top1.ch8c.data[0] ;
 wire \top1.ch8c.data[10] ;
 wire \top1.ch8c.data[11] ;
 wire \top1.ch8c.data[1] ;
 wire \top1.ch8c.data[2] ;
 wire \top1.ch8c.data[3] ;
 wire \top1.ch8c.data[4] ;
 wire \top1.ch8c.data[5] ;
 wire \top1.ch8c.data[6] ;
 wire \top1.ch8c.data[7] ;
 wire \top1.ch8c.data[8] ;
 wire \top1.ch8c.data[9] ;
 wire \top1.ch8c.ovf ;
 wire \top1.ch9c.data[0] ;
 wire \top1.ch9c.data[10] ;
 wire \top1.ch9c.data[11] ;
 wire \top1.ch9c.data[1] ;
 wire \top1.ch9c.data[2] ;
 wire \top1.ch9c.data[3] ;
 wire \top1.ch9c.data[4] ;
 wire \top1.ch9c.data[5] ;
 wire \top1.ch9c.data[6] ;
 wire \top1.ch9c.data[7] ;
 wire \top1.ch9c.data[8] ;
 wire \top1.ch9c.data[9] ;
 wire \top1.ch9c.ovf ;
 wire \top1.data[0][0] ;
 wire \top1.data[0][10] ;
 wire \top1.data[0][11] ;
 wire \top1.data[0][1] ;
 wire \top1.data[0][2] ;
 wire \top1.data[0][3] ;
 wire \top1.data[0][4] ;
 wire \top1.data[0][5] ;
 wire \top1.data[0][6] ;
 wire \top1.data[0][7] ;
 wire \top1.data[0][8] ;
 wire \top1.data[0][9] ;
 wire \top1.ovf_RTC ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net1;
 wire net2;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;

 sg13g2_inv_1 _1247_ (.Y(_0807_),
    .A(\top1.ch9c.data[7] ));
 sg13g2_inv_1 _1248_ (.Y(_0808_),
    .A(\top1.ch9c.data[2] ));
 sg13g2_inv_1 _1249_ (.Y(_0809_),
    .A(\top1.ch15c.data[7] ));
 sg13g2_inv_1 _1250_ (.Y(_0810_),
    .A(\top1.ch15c.data[2] ));
 sg13g2_inv_1 _1251_ (.Y(_0811_),
    .A(\top1.ch1c.data[7] ));
 sg13g2_inv_1 _1252_ (.Y(_0812_),
    .A(\top1.ch1c.data[2] ));
 sg13g2_inv_1 _1253_ (.Y(_0813_),
    .A(\top1.ch2c.data[7] ));
 sg13g2_inv_1 _1254_ (.Y(_0814_),
    .A(\top1.ch2c.data[2] ));
 sg13g2_inv_1 _1255_ (.Y(_0815_),
    .A(\top1.ch3c.data[7] ));
 sg13g2_inv_1 _1256_ (.Y(_0816_),
    .A(\top1.ch3c.data[2] ));
 sg13g2_inv_1 _1257_ (.Y(_0817_),
    .A(\top1.ch4c.data[3] ));
 sg13g2_inv_1 _1258_ (.Y(_0818_),
    .A(\top1.ch5c.data[7] ));
 sg13g2_inv_1 _1259_ (.Y(_0819_),
    .A(\top1.ch5c.data[2] ));
 sg13g2_inv_1 _1260_ (.Y(_0820_),
    .A(\top1.ch6c.data[6] ));
 sg13g2_inv_1 _1261_ (.Y(_0821_),
    .A(\top1.ch6c.data[2] ));
 sg13g2_inv_1 _1262_ (.Y(_0822_),
    .A(\top1.ch7c.data[6] ));
 sg13g2_inv_1 _1263_ (.Y(_0823_),
    .A(\top1.ch7c.data[2] ));
 sg13g2_inv_1 _1264_ (.Y(_0824_),
    .A(\top1.ch8c.data[7] ));
 sg13g2_inv_1 _1265_ (.Y(_0825_),
    .A(\top1.ch8c.data[2] ));
 sg13g2_inv_1 _1266_ (.Y(_0826_),
    .A(\top1.ch10c.data[7] ));
 sg13g2_inv_1 _1267_ (.Y(_0827_),
    .A(\top1.ch10c.data[2] ));
 sg13g2_inv_1 _1268_ (.Y(_0828_),
    .A(\top1.ch11c.data[7] ));
 sg13g2_inv_1 _1269_ (.Y(_0829_),
    .A(\top1.ch11c.data[2] ));
 sg13g2_inv_1 _1270_ (.Y(_0830_),
    .A(\top1.ch12c.data[7] ));
 sg13g2_inv_1 _1271_ (.Y(_0831_),
    .A(\top1.ch12c.data[2] ));
 sg13g2_inv_1 _1272_ (.Y(_0832_),
    .A(\top1.ch13c.data[7] ));
 sg13g2_inv_1 _1273_ (.Y(_0833_),
    .A(\top1.ch13c.data[2] ));
 sg13g2_inv_1 _1274_ (.Y(_0834_),
    .A(\top1.ch14c.data[7] ));
 sg13g2_inv_1 _1275_ (.Y(_0835_),
    .A(\top1.ch14c.data[2] ));
 sg13g2_inv_1 _1276_ (.Y(_0836_),
    .A(net607));
 sg13g2_inv_1 _1277_ (.Y(_0837_),
    .A(\top1.FSM1.state_reg[4] ));
 sg13g2_inv_1 _1278_ (.Y(_0838_),
    .A(net600));
 sg13g2_inv_1 _1279_ (.Y(_0011_),
    .A(\top1.data[0][0] ));
 sg13g2_inv_1 _1280_ (.Y(_0839_),
    .A(\top1.data[0][11] ));
 sg13g2_inv_1 _1281_ (.Y(_0840_),
    .A(net43));
 sg13g2_nand4_1 _1282_ (.B(\top1.ch1c.data[2] ),
    .C(\top1.ch1c.data[1] ),
    .A(\top1.ch1c.data[3] ),
    .Y(_0841_),
    .D(\top1.ch1c.data[0] ));
 sg13g2_and2_1 _1283_ (.A(\top1.ch1c.data[10] ),
    .B(\top1.ch1c.data[9] ),
    .X(_0842_));
 sg13g2_nand2_1 _1284_ (.Y(_0843_),
    .A(\top1.ch1c.data[10] ),
    .B(\top1.ch1c.data[9] ));
 sg13g2_nand4_1 _1285_ (.B(\top1.ch1c.data[6] ),
    .C(\top1.ch1c.data[5] ),
    .A(\top1.ch1c.data[7] ),
    .Y(_0844_),
    .D(\top1.ch1c.data[4] ));
 sg13g2_nand2_1 _1286_ (.Y(_0845_),
    .A(\top1.ch1c.data[11] ),
    .B(\top1.ch1c.data[8] ));
 sg13g2_nor4_1 _1287_ (.A(_0841_),
    .B(_0843_),
    .C(_0844_),
    .D(_0845_),
    .Y(_0846_));
 sg13g2_or2_1 _1288_ (.X(_0435_),
    .B(_0846_),
    .A(\top1.ch1c.ovf ));
 sg13g2_nand4_1 _1289_ (.B(\top1.ch2c.data[2] ),
    .C(\top1.ch2c.data[1] ),
    .A(\top1.ch2c.data[3] ),
    .Y(_0847_),
    .D(\top1.ch2c.data[0] ));
 sg13g2_and2_1 _1290_ (.A(\top1.ch2c.data[10] ),
    .B(\top1.ch2c.data[9] ),
    .X(_0848_));
 sg13g2_nand2_1 _1291_ (.Y(_0849_),
    .A(\top1.ch2c.data[10] ),
    .B(\top1.ch2c.data[9] ));
 sg13g2_nand4_1 _1292_ (.B(\top1.ch2c.data[6] ),
    .C(\top1.ch2c.data[5] ),
    .A(\top1.ch2c.data[7] ),
    .Y(_0850_),
    .D(\top1.ch2c.data[4] ));
 sg13g2_nand2_1 _1293_ (.Y(_0851_),
    .A(\top1.ch2c.data[11] ),
    .B(\top1.ch2c.data[8] ));
 sg13g2_nor4_1 _1294_ (.A(_0847_),
    .B(_0849_),
    .C(_0850_),
    .D(_0851_),
    .Y(_0852_));
 sg13g2_or2_1 _1295_ (.X(_0434_),
    .B(_0852_),
    .A(\top1.ch2c.ovf ));
 sg13g2_nand4_1 _1296_ (.B(\top1.ch3c.data[2] ),
    .C(\top1.ch3c.data[1] ),
    .A(\top1.ch3c.data[3] ),
    .Y(_0853_),
    .D(\top1.ch3c.data[0] ));
 sg13g2_and2_1 _1297_ (.A(\top1.ch3c.data[10] ),
    .B(\top1.ch3c.data[9] ),
    .X(_0854_));
 sg13g2_nand2_1 _1298_ (.Y(_0855_),
    .A(\top1.ch3c.data[10] ),
    .B(\top1.ch3c.data[9] ));
 sg13g2_nand4_1 _1299_ (.B(\top1.ch3c.data[6] ),
    .C(\top1.ch3c.data[5] ),
    .A(\top1.ch3c.data[7] ),
    .Y(_0856_),
    .D(\top1.ch3c.data[4] ));
 sg13g2_nand2_1 _1300_ (.Y(_0857_),
    .A(\top1.ch3c.data[11] ),
    .B(\top1.ch3c.data[8] ));
 sg13g2_nor4_1 _1301_ (.A(_0853_),
    .B(_0855_),
    .C(_0856_),
    .D(_0857_),
    .Y(_0858_));
 sg13g2_or2_1 _1302_ (.X(_0433_),
    .B(_0858_),
    .A(\top1.ch3c.ovf ));
 sg13g2_nand4_1 _1303_ (.B(\top1.ch4c.data[2] ),
    .C(\top1.ch4c.data[1] ),
    .A(\top1.ch4c.data[3] ),
    .Y(_0859_),
    .D(\top1.ch4c.data[0] ));
 sg13g2_nand2_1 _1304_ (.Y(_0860_),
    .A(\top1.ch4c.data[11] ),
    .B(\top1.ch4c.data[8] ));
 sg13g2_nand4_1 _1305_ (.B(\top1.ch4c.data[6] ),
    .C(\top1.ch4c.data[5] ),
    .A(\top1.ch4c.data[7] ),
    .Y(_0861_),
    .D(\top1.ch4c.data[4] ));
 sg13g2_nand2_1 _1306_ (.Y(_0862_),
    .A(\top1.ch4c.data[10] ),
    .B(\top1.ch4c.data[9] ));
 sg13g2_nor4_1 _1307_ (.A(_0859_),
    .B(_0860_),
    .C(_0861_),
    .D(_0862_),
    .Y(_0863_));
 sg13g2_or2_1 _1308_ (.X(_0432_),
    .B(_0863_),
    .A(\top1.ch4c.ovf ));
 sg13g2_nand4_1 _1309_ (.B(\top1.ch5c.data[2] ),
    .C(\top1.ch5c.data[1] ),
    .A(\top1.ch5c.data[3] ),
    .Y(_0864_),
    .D(\top1.ch5c.data[0] ));
 sg13g2_nand2_1 _1310_ (.Y(_0865_),
    .A(\top1.ch5c.data[11] ),
    .B(\top1.ch5c.data[8] ));
 sg13g2_nand4_1 _1311_ (.B(\top1.ch5c.data[6] ),
    .C(\top1.ch5c.data[5] ),
    .A(\top1.ch5c.data[7] ),
    .Y(_0866_),
    .D(\top1.ch5c.data[4] ));
 sg13g2_and2_1 _1312_ (.A(\top1.ch5c.data[10] ),
    .B(\top1.ch5c.data[9] ),
    .X(_0867_));
 sg13g2_nand2_1 _1313_ (.Y(_0868_),
    .A(\top1.ch5c.data[10] ),
    .B(\top1.ch5c.data[9] ));
 sg13g2_nor4_2 _1314_ (.A(_0864_),
    .B(_0865_),
    .C(_0866_),
    .Y(_0869_),
    .D(_0868_));
 sg13g2_or2_1 _1315_ (.X(_0431_),
    .B(_0869_),
    .A(\top1.ch5c.ovf ));
 sg13g2_nand4_1 _1316_ (.B(\top1.ch6c.data[2] ),
    .C(\top1.ch6c.data[1] ),
    .A(\top1.ch6c.data[3] ),
    .Y(_0870_),
    .D(\top1.ch6c.data[0] ));
 sg13g2_nand2_1 _1317_ (.Y(_0871_),
    .A(\top1.ch6c.data[10] ),
    .B(\top1.ch6c.data[9] ));
 sg13g2_nand4_1 _1318_ (.B(\top1.ch6c.data[6] ),
    .C(\top1.ch6c.data[5] ),
    .A(\top1.ch6c.data[7] ),
    .Y(_0872_),
    .D(\top1.ch6c.data[4] ));
 sg13g2_nand2_1 _1319_ (.Y(_0873_),
    .A(\top1.ch6c.data[11] ),
    .B(\top1.ch6c.data[8] ));
 sg13g2_nor4_1 _1320_ (.A(_0870_),
    .B(_0871_),
    .C(_0872_),
    .D(_0873_),
    .Y(_0874_));
 sg13g2_or2_1 _1321_ (.X(_0430_),
    .B(_0874_),
    .A(\top1.ch6c.ovf ));
 sg13g2_nand4_1 _1322_ (.B(\top1.ch7c.data[2] ),
    .C(\top1.ch7c.data[1] ),
    .A(\top1.ch7c.data[3] ),
    .Y(_0875_),
    .D(\top1.ch7c.data[0] ));
 sg13g2_nand2_1 _1323_ (.Y(_0876_),
    .A(\top1.ch7c.data[10] ),
    .B(\top1.ch7c.data[9] ));
 sg13g2_nand4_1 _1324_ (.B(\top1.ch7c.data[6] ),
    .C(\top1.ch7c.data[5] ),
    .A(\top1.ch7c.data[7] ),
    .Y(_0877_),
    .D(\top1.ch7c.data[4] ));
 sg13g2_nand2_1 _1325_ (.Y(_0878_),
    .A(\top1.ch7c.data[11] ),
    .B(\top1.ch7c.data[8] ));
 sg13g2_nor4_1 _1326_ (.A(_0875_),
    .B(_0876_),
    .C(_0877_),
    .D(_0878_),
    .Y(_0879_));
 sg13g2_or2_1 _1327_ (.X(_0429_),
    .B(_0879_),
    .A(\top1.ch7c.ovf ));
 sg13g2_nand2_1 _1328_ (.Y(_0880_),
    .A(\top1.ch8c.data[9] ),
    .B(\top1.ch8c.data[8] ));
 sg13g2_nand4_1 _1329_ (.B(\top1.ch8c.data[4] ),
    .C(\top1.ch8c.data[1] ),
    .A(\top1.ch8c.data[5] ),
    .Y(_0881_),
    .D(\top1.ch8c.data[0] ));
 sg13g2_nand4_1 _1330_ (.B(\top1.ch8c.data[6] ),
    .C(\top1.ch8c.data[3] ),
    .A(\top1.ch8c.data[7] ),
    .Y(_0882_),
    .D(\top1.ch8c.data[2] ));
 sg13g2_nor3_1 _1331_ (.A(_0880_),
    .B(_0881_),
    .C(_0882_),
    .Y(_0883_));
 sg13g2_nand4_1 _1332_ (.B(\top1.ch8c.data[2] ),
    .C(\top1.ch8c.data[1] ),
    .A(\top1.ch8c.data[3] ),
    .Y(_0884_),
    .D(\top1.ch8c.data[0] ));
 sg13g2_nand4_1 _1333_ (.B(\top1.ch8c.data[6] ),
    .C(\top1.ch8c.data[5] ),
    .A(\top1.ch8c.data[7] ),
    .Y(_0885_),
    .D(\top1.ch8c.data[4] ));
 sg13g2_nand3_1 _1334_ (.B(\top1.ch8c.data[10] ),
    .C(_0883_),
    .A(\top1.ch8c.data[11] ),
    .Y(_0886_));
 sg13g2_nand2b_1 _1335_ (.Y(_0428_),
    .B(_0886_),
    .A_N(\top1.ch8c.ovf ));
 sg13g2_nand4_1 _1336_ (.B(\top1.ch9c.data[2] ),
    .C(\top1.ch9c.data[1] ),
    .A(\top1.ch9c.data[3] ),
    .Y(_0887_),
    .D(\top1.ch9c.data[0] ));
 sg13g2_and2_1 _1337_ (.A(\top1.ch9c.data[10] ),
    .B(\top1.ch9c.data[9] ),
    .X(_0888_));
 sg13g2_nand2_1 _1338_ (.Y(_0889_),
    .A(\top1.ch9c.data[10] ),
    .B(\top1.ch9c.data[9] ));
 sg13g2_nand4_1 _1339_ (.B(\top1.ch9c.data[6] ),
    .C(\top1.ch9c.data[5] ),
    .A(\top1.ch9c.data[7] ),
    .Y(_0890_),
    .D(\top1.ch9c.data[4] ));
 sg13g2_nand2_1 _1340_ (.Y(_0891_),
    .A(\top1.ch9c.data[11] ),
    .B(\top1.ch9c.data[8] ));
 sg13g2_nor4_1 _1341_ (.A(_0887_),
    .B(_0889_),
    .C(_0890_),
    .D(_0891_),
    .Y(_0892_));
 sg13g2_or2_1 _1342_ (.X(_0427_),
    .B(_0892_),
    .A(\top1.ch9c.ovf ));
 sg13g2_nand4_1 _1343_ (.B(\top1.ch10c.data[2] ),
    .C(\top1.ch10c.data[1] ),
    .A(\top1.ch10c.data[3] ),
    .Y(_0893_),
    .D(\top1.ch10c.data[0] ));
 sg13g2_nand2_1 _1344_ (.Y(_0894_),
    .A(\top1.ch10c.data[11] ),
    .B(\top1.ch10c.data[8] ));
 sg13g2_nand4_1 _1345_ (.B(\top1.ch10c.data[6] ),
    .C(\top1.ch10c.data[5] ),
    .A(\top1.ch10c.data[7] ),
    .Y(_0895_),
    .D(\top1.ch10c.data[4] ));
 sg13g2_and2_1 _1346_ (.A(\top1.ch10c.data[10] ),
    .B(\top1.ch10c.data[9] ),
    .X(_0896_));
 sg13g2_nand2_1 _1347_ (.Y(_0897_),
    .A(\top1.ch10c.data[10] ),
    .B(\top1.ch10c.data[9] ));
 sg13g2_nor4_1 _1348_ (.A(_0893_),
    .B(_0894_),
    .C(_0895_),
    .D(_0897_),
    .Y(_0898_));
 sg13g2_or2_1 _1349_ (.X(_0426_),
    .B(_0898_),
    .A(\top1.ch10c.ovf ));
 sg13g2_nand4_1 _1350_ (.B(\top1.ch11c.data[2] ),
    .C(\top1.ch11c.data[1] ),
    .A(\top1.ch11c.data[3] ),
    .Y(_0899_),
    .D(\top1.ch11c.data[0] ));
 sg13g2_nand2_1 _1351_ (.Y(_0900_),
    .A(\top1.ch11c.data[11] ),
    .B(\top1.ch11c.data[8] ));
 sg13g2_nand4_1 _1352_ (.B(\top1.ch11c.data[6] ),
    .C(\top1.ch11c.data[5] ),
    .A(\top1.ch11c.data[7] ),
    .Y(_0901_),
    .D(\top1.ch11c.data[4] ));
 sg13g2_and2_1 _1353_ (.A(\top1.ch11c.data[10] ),
    .B(\top1.ch11c.data[9] ),
    .X(_0902_));
 sg13g2_nand2_1 _1354_ (.Y(_0903_),
    .A(\top1.ch11c.data[10] ),
    .B(\top1.ch11c.data[9] ));
 sg13g2_nor4_2 _1355_ (.A(_0899_),
    .B(_0900_),
    .C(_0901_),
    .Y(_0904_),
    .D(_0903_));
 sg13g2_or2_1 _1356_ (.X(_0425_),
    .B(_0904_),
    .A(\top1.ch11c.ovf ));
 sg13g2_nand4_1 _1357_ (.B(\top1.ch12c.data[2] ),
    .C(\top1.ch12c.data[1] ),
    .A(\top1.ch12c.data[3] ),
    .Y(_0905_),
    .D(\top1.ch12c.data[0] ));
 sg13g2_and2_1 _1358_ (.A(\top1.ch12c.data[10] ),
    .B(\top1.ch12c.data[9] ),
    .X(_0906_));
 sg13g2_nand2_1 _1359_ (.Y(_0907_),
    .A(\top1.ch12c.data[10] ),
    .B(\top1.ch12c.data[9] ));
 sg13g2_nand4_1 _1360_ (.B(\top1.ch12c.data[6] ),
    .C(\top1.ch12c.data[5] ),
    .A(\top1.ch12c.data[7] ),
    .Y(_0908_),
    .D(\top1.ch12c.data[4] ));
 sg13g2_nand2_1 _1361_ (.Y(_0909_),
    .A(\top1.ch12c.data[11] ),
    .B(\top1.ch12c.data[8] ));
 sg13g2_nor4_1 _1362_ (.A(_0905_),
    .B(_0907_),
    .C(_0908_),
    .D(_0909_),
    .Y(_0910_));
 sg13g2_or2_1 _1363_ (.X(_0424_),
    .B(_0910_),
    .A(\top1.ch12c.ovf ));
 sg13g2_nand4_1 _1364_ (.B(\top1.ch13c.data[2] ),
    .C(\top1.ch13c.data[1] ),
    .A(\top1.ch13c.data[3] ),
    .Y(_0911_),
    .D(\top1.ch13c.data[0] ));
 sg13g2_and2_1 _1365_ (.A(\top1.ch13c.data[10] ),
    .B(\top1.ch13c.data[9] ),
    .X(_0912_));
 sg13g2_nand2_1 _1366_ (.Y(_0913_),
    .A(\top1.ch13c.data[10] ),
    .B(\top1.ch13c.data[9] ));
 sg13g2_nand4_1 _1367_ (.B(\top1.ch13c.data[6] ),
    .C(\top1.ch13c.data[5] ),
    .A(\top1.ch13c.data[7] ),
    .Y(_0914_),
    .D(\top1.ch13c.data[4] ));
 sg13g2_nand2_1 _1368_ (.Y(_0915_),
    .A(\top1.ch13c.data[11] ),
    .B(\top1.ch13c.data[8] ));
 sg13g2_nor4_1 _1369_ (.A(_0911_),
    .B(_0913_),
    .C(_0914_),
    .D(_0915_),
    .Y(_0916_));
 sg13g2_or2_1 _1370_ (.X(_0423_),
    .B(_0916_),
    .A(\top1.ch13c.ovf ));
 sg13g2_nand4_1 _1371_ (.B(\top1.ch14c.data[2] ),
    .C(\top1.ch14c.data[1] ),
    .A(\top1.ch14c.data[3] ),
    .Y(_0917_),
    .D(\top1.ch14c.data[0] ));
 sg13g2_and2_1 _1372_ (.A(\top1.ch14c.data[10] ),
    .B(\top1.ch14c.data[9] ),
    .X(_0918_));
 sg13g2_nand2_1 _1373_ (.Y(_0919_),
    .A(\top1.ch14c.data[10] ),
    .B(\top1.ch14c.data[9] ));
 sg13g2_nand4_1 _1374_ (.B(\top1.ch14c.data[6] ),
    .C(\top1.ch14c.data[5] ),
    .A(\top1.ch14c.data[7] ),
    .Y(_0920_),
    .D(\top1.ch14c.data[4] ));
 sg13g2_nand2_1 _1375_ (.Y(_0921_),
    .A(\top1.ch14c.data[11] ),
    .B(\top1.ch14c.data[8] ));
 sg13g2_nor4_1 _1376_ (.A(_0917_),
    .B(_0919_),
    .C(_0920_),
    .D(_0921_),
    .Y(_0922_));
 sg13g2_or2_1 _1377_ (.X(_0422_),
    .B(_0922_),
    .A(\top1.ch14c.ovf ));
 sg13g2_nand4_1 _1378_ (.B(\top1.ch15c.data[2] ),
    .C(\top1.ch15c.data[1] ),
    .A(\top1.ch15c.data[3] ),
    .Y(_0923_),
    .D(\top1.ch15c.data[0] ));
 sg13g2_and2_1 _1379_ (.A(\top1.ch15c.data[10] ),
    .B(\top1.ch15c.data[9] ),
    .X(_0924_));
 sg13g2_nand2_1 _1380_ (.Y(_0925_),
    .A(\top1.ch15c.data[10] ),
    .B(\top1.ch15c.data[9] ));
 sg13g2_nand4_1 _1381_ (.B(\top1.ch15c.data[6] ),
    .C(\top1.ch15c.data[5] ),
    .A(\top1.ch15c.data[7] ),
    .Y(_0926_),
    .D(\top1.ch15c.data[4] ));
 sg13g2_nand2_1 _1382_ (.Y(_0927_),
    .A(\top1.ch15c.data[11] ),
    .B(\top1.ch15c.data[8] ));
 sg13g2_nor4_1 _1383_ (.A(_0923_),
    .B(_0925_),
    .C(_0926_),
    .D(_0927_),
    .Y(_0928_));
 sg13g2_or2_1 _1384_ (.X(_0421_),
    .B(_0928_),
    .A(\top1.ch15c.ovf ));
 sg13g2_nor4_1 _1385_ (.A(\top1.ch5c.ovf ),
    .B(\top1.ch6c.ovf ),
    .C(\top1.ch7c.ovf ),
    .D(\top1.ch8c.ovf ),
    .Y(_0929_));
 sg13g2_nor4_2 _1386_ (.A(\top1.ch1c.ovf ),
    .B(\top1.ch2c.ovf ),
    .C(\top1.ch3c.ovf ),
    .Y(_0930_),
    .D(\top1.ch4c.ovf ));
 sg13g2_nor4_1 _1387_ (.A(\top1.ch9c.ovf ),
    .B(\top1.ch10c.ovf ),
    .C(\top1.ch11c.ovf ),
    .D(\top1.ch12c.ovf ),
    .Y(_0931_));
 sg13g2_nor4_2 _1388_ (.A(\top1.ch13c.ovf ),
    .B(\top1.ch14c.ovf ),
    .C(\top1.ch15c.ovf ),
    .Y(_0932_),
    .D(\top1.ovf_RTC ));
 sg13g2_and4_1 _1389_ (.A(_0929_),
    .B(_0930_),
    .C(_0931_),
    .D(_0932_),
    .X(_0933_));
 sg13g2_inv_1 _1390_ (.Y(\top1.FSM1.ovf ),
    .A(net594));
 sg13g2_nor2_2 _1391_ (.A(_0887_),
    .B(net537),
    .Y(_0934_));
 sg13g2_nor3_2 _1392_ (.A(_0887_),
    .B(_0890_),
    .C(net537),
    .Y(_0935_));
 sg13g2_and2_1 _1393_ (.A(\top1.ch9c.data[8] ),
    .B(_0935_),
    .X(_0936_));
 sg13g2_nand2_1 _1394_ (.Y(_0937_),
    .A(_0888_),
    .B(_0936_));
 sg13g2_nand3_1 _1395_ (.B(\top1.ch9c.data[0] ),
    .C(net598),
    .A(\top1.ch9c.data[1] ),
    .Y(_0938_));
 sg13g2_nor2_1 _1396_ (.A(_0808_),
    .B(_0938_),
    .Y(_0939_));
 sg13g2_nand4_1 _1397_ (.B(\top1.ch9c.data[4] ),
    .C(\top1.ch9c.data[3] ),
    .A(\top1.ch9c.data[5] ),
    .Y(_0940_),
    .D(_0939_));
 sg13g2_xnor2_1 _1398_ (.Y(_0416_),
    .A(\top1.ch9c.data[11] ),
    .B(_0937_));
 sg13g2_a21oi_1 _1399_ (.A1(\top1.ch9c.data[9] ),
    .A2(_0936_),
    .Y(_0941_),
    .B1(\top1.ch9c.data[10] ));
 sg13g2_a21oi_1 _1400_ (.A1(_0888_),
    .A2(_0936_),
    .Y(_0415_),
    .B1(_0941_));
 sg13g2_xor2_1 _1401_ (.B(_0936_),
    .A(\top1.ch9c.data[9] ),
    .X(_0414_));
 sg13g2_xor2_1 _1402_ (.B(_0935_),
    .A(\top1.ch9c.data[8] ),
    .X(_0413_));
 sg13g2_nand2_1 _1403_ (.Y(_0942_),
    .A(\top1.ch9c.data[4] ),
    .B(_0934_));
 sg13g2_nand4_1 _1404_ (.B(\top1.ch9c.data[5] ),
    .C(\top1.ch9c.data[4] ),
    .A(\top1.ch9c.data[6] ),
    .Y(_0943_),
    .D(_0934_));
 sg13g2_a21oi_1 _1405_ (.A1(_0807_),
    .A2(_0943_),
    .Y(_0412_),
    .B1(_0935_));
 sg13g2_xnor2_1 _1406_ (.Y(_0411_),
    .A(\top1.ch9c.data[6] ),
    .B(_0940_));
 sg13g2_xnor2_1 _1407_ (.Y(_0410_),
    .A(\top1.ch9c.data[5] ),
    .B(_0942_));
 sg13g2_xor2_1 _1408_ (.B(_0934_),
    .A(\top1.ch9c.data[4] ),
    .X(_0409_));
 sg13g2_xor2_1 _1409_ (.B(_0939_),
    .A(\top1.ch9c.data[3] ),
    .X(_0408_));
 sg13g2_xnor2_1 _1410_ (.Y(_0407_),
    .A(\top1.ch9c.data[2] ),
    .B(_0938_));
 sg13g2_a21o_1 _1411_ (.A2(net598),
    .A1(\top1.ch9c.data[0] ),
    .B1(\top1.ch9c.data[1] ),
    .X(_0944_));
 sg13g2_and2_1 _1412_ (.A(_0938_),
    .B(_0944_),
    .X(_0406_));
 sg13g2_mux2_1 _1413_ (.A0(_0018_),
    .A1(\top1.ch9c.data[0] ),
    .S(net537),
    .X(_0405_));
 sg13g2_nor2_1 _1414_ (.A(_0923_),
    .B(net540),
    .Y(_0945_));
 sg13g2_nor3_2 _1415_ (.A(_0923_),
    .B(_0926_),
    .C(net540),
    .Y(_0946_));
 sg13g2_and2_1 _1416_ (.A(\top1.ch15c.data[8] ),
    .B(_0946_),
    .X(_0947_));
 sg13g2_nand2_1 _1417_ (.Y(_0948_),
    .A(_0924_),
    .B(_0947_));
 sg13g2_nand3_1 _1418_ (.B(\top1.ch15c.data[0] ),
    .C(net596),
    .A(\top1.ch15c.data[1] ),
    .Y(_0949_));
 sg13g2_nor2_1 _1419_ (.A(_0810_),
    .B(_0949_),
    .Y(_0950_));
 sg13g2_nand4_1 _1420_ (.B(\top1.ch15c.data[4] ),
    .C(\top1.ch15c.data[3] ),
    .A(\top1.ch15c.data[5] ),
    .Y(_0951_),
    .D(_0950_));
 sg13g2_xnor2_1 _1421_ (.Y(_0398_),
    .A(\top1.ch15c.data[11] ),
    .B(_0948_));
 sg13g2_a21oi_1 _1422_ (.A1(\top1.ch15c.data[9] ),
    .A2(_0947_),
    .Y(_0952_),
    .B1(\top1.ch15c.data[10] ));
 sg13g2_a21oi_1 _1423_ (.A1(_0924_),
    .A2(_0947_),
    .Y(_0397_),
    .B1(_0952_));
 sg13g2_xor2_1 _1424_ (.B(_0947_),
    .A(\top1.ch15c.data[9] ),
    .X(_0396_));
 sg13g2_xor2_1 _1425_ (.B(_0946_),
    .A(\top1.ch15c.data[8] ),
    .X(_0395_));
 sg13g2_nand2_1 _1426_ (.Y(_0953_),
    .A(\top1.ch15c.data[4] ),
    .B(_0945_));
 sg13g2_nand4_1 _1427_ (.B(\top1.ch15c.data[5] ),
    .C(\top1.ch15c.data[4] ),
    .A(\top1.ch15c.data[6] ),
    .Y(_0954_),
    .D(_0945_));
 sg13g2_a21oi_1 _1428_ (.A1(_0809_),
    .A2(_0954_),
    .Y(_0394_),
    .B1(_0946_));
 sg13g2_xnor2_1 _1429_ (.Y(_0393_),
    .A(\top1.ch15c.data[6] ),
    .B(_0951_));
 sg13g2_xnor2_1 _1430_ (.Y(_0392_),
    .A(\top1.ch15c.data[5] ),
    .B(_0953_));
 sg13g2_xor2_1 _1431_ (.B(_0945_),
    .A(\top1.ch15c.data[4] ),
    .X(_0391_));
 sg13g2_xor2_1 _1432_ (.B(_0950_),
    .A(\top1.ch15c.data[3] ),
    .X(_0390_));
 sg13g2_xnor2_1 _1433_ (.Y(_0389_),
    .A(\top1.ch15c.data[2] ),
    .B(_0949_));
 sg13g2_a21o_1 _1434_ (.A2(net596),
    .A1(\top1.ch15c.data[0] ),
    .B1(\top1.ch15c.data[1] ),
    .X(_0955_));
 sg13g2_and2_1 _1435_ (.A(_0949_),
    .B(_0955_),
    .X(_0388_));
 sg13g2_mux2_1 _1436_ (.A0(_0019_),
    .A1(\top1.ch15c.data[0] ),
    .S(net535),
    .X(_0387_));
 sg13g2_nor2_1 _1437_ (.A(_0841_),
    .B(net539),
    .Y(_0956_));
 sg13g2_nor3_2 _1438_ (.A(_0841_),
    .B(_0844_),
    .C(net539),
    .Y(_0957_));
 sg13g2_and2_1 _1439_ (.A(\top1.ch1c.data[8] ),
    .B(_0957_),
    .X(_0958_));
 sg13g2_nand2_1 _1440_ (.Y(_0959_),
    .A(_0842_),
    .B(_0958_));
 sg13g2_nand3_1 _1441_ (.B(\top1.ch1c.data[0] ),
    .C(net597),
    .A(\top1.ch1c.data[1] ),
    .Y(_0960_));
 sg13g2_nor2_1 _1442_ (.A(_0812_),
    .B(_0960_),
    .Y(_0961_));
 sg13g2_nand4_1 _1443_ (.B(\top1.ch1c.data[4] ),
    .C(\top1.ch1c.data[3] ),
    .A(\top1.ch1c.data[5] ),
    .Y(_0962_),
    .D(_0961_));
 sg13g2_xnor2_1 _1444_ (.Y(_0386_),
    .A(\top1.ch1c.data[11] ),
    .B(_0959_));
 sg13g2_a21oi_1 _1445_ (.A1(\top1.ch1c.data[9] ),
    .A2(_0958_),
    .Y(_0963_),
    .B1(\top1.ch1c.data[10] ));
 sg13g2_a21oi_1 _1446_ (.A1(_0842_),
    .A2(_0958_),
    .Y(_0385_),
    .B1(_0963_));
 sg13g2_xor2_1 _1447_ (.B(_0958_),
    .A(\top1.ch1c.data[9] ),
    .X(_0384_));
 sg13g2_xor2_1 _1448_ (.B(_0957_),
    .A(\top1.ch1c.data[8] ),
    .X(_0383_));
 sg13g2_nand2_1 _1449_ (.Y(_0964_),
    .A(\top1.ch1c.data[4] ),
    .B(_0956_));
 sg13g2_nand4_1 _1450_ (.B(\top1.ch1c.data[5] ),
    .C(\top1.ch1c.data[4] ),
    .A(\top1.ch1c.data[6] ),
    .Y(_0965_),
    .D(_0956_));
 sg13g2_a21oi_1 _1451_ (.A1(_0811_),
    .A2(_0965_),
    .Y(_0382_),
    .B1(_0957_));
 sg13g2_xnor2_1 _1452_ (.Y(_0381_),
    .A(\top1.ch1c.data[6] ),
    .B(_0962_));
 sg13g2_xnor2_1 _1453_ (.Y(_0380_),
    .A(\top1.ch1c.data[5] ),
    .B(_0964_));
 sg13g2_xor2_1 _1454_ (.B(_0956_),
    .A(\top1.ch1c.data[4] ),
    .X(_0379_));
 sg13g2_xor2_1 _1455_ (.B(_0961_),
    .A(\top1.ch1c.data[3] ),
    .X(_0378_));
 sg13g2_xnor2_1 _1456_ (.Y(_0377_),
    .A(\top1.ch1c.data[2] ),
    .B(_0960_));
 sg13g2_a21o_1 _1457_ (.A2(net597),
    .A1(\top1.ch1c.data[0] ),
    .B1(\top1.ch1c.data[1] ),
    .X(_0966_));
 sg13g2_and2_1 _1458_ (.A(_0960_),
    .B(_0966_),
    .X(_0376_));
 sg13g2_mux2_1 _1459_ (.A0(_0020_),
    .A1(\top1.ch1c.data[0] ),
    .S(net539),
    .X(_0375_));
 sg13g2_nor2_1 _1460_ (.A(_0847_),
    .B(net539),
    .Y(_0967_));
 sg13g2_nor3_2 _1461_ (.A(_0847_),
    .B(_0850_),
    .C(net539),
    .Y(_0968_));
 sg13g2_and2_1 _1462_ (.A(\top1.ch2c.data[8] ),
    .B(_0968_),
    .X(_0969_));
 sg13g2_nand2_1 _1463_ (.Y(_0970_),
    .A(_0848_),
    .B(_0969_));
 sg13g2_nand3_1 _1464_ (.B(\top1.ch2c.data[0] ),
    .C(net599),
    .A(\top1.ch2c.data[1] ),
    .Y(_0971_));
 sg13g2_nor2_1 _1465_ (.A(_0814_),
    .B(_0971_),
    .Y(_0972_));
 sg13g2_nand4_1 _1466_ (.B(\top1.ch2c.data[4] ),
    .C(\top1.ch2c.data[3] ),
    .A(\top1.ch2c.data[5] ),
    .Y(_0973_),
    .D(_0972_));
 sg13g2_xnor2_1 _1467_ (.Y(_0374_),
    .A(\top1.ch2c.data[11] ),
    .B(_0970_));
 sg13g2_a21oi_1 _1468_ (.A1(\top1.ch2c.data[9] ),
    .A2(_0969_),
    .Y(_0974_),
    .B1(\top1.ch2c.data[10] ));
 sg13g2_a21oi_1 _1469_ (.A1(_0848_),
    .A2(_0969_),
    .Y(_0373_),
    .B1(_0974_));
 sg13g2_xor2_1 _1470_ (.B(_0969_),
    .A(\top1.ch2c.data[9] ),
    .X(_0372_));
 sg13g2_xor2_1 _1471_ (.B(_0968_),
    .A(\top1.ch2c.data[8] ),
    .X(_0371_));
 sg13g2_nand2_1 _1472_ (.Y(_0975_),
    .A(\top1.ch2c.data[4] ),
    .B(_0967_));
 sg13g2_nand4_1 _1473_ (.B(\top1.ch2c.data[5] ),
    .C(\top1.ch2c.data[4] ),
    .A(\top1.ch2c.data[6] ),
    .Y(_0976_),
    .D(_0967_));
 sg13g2_a21oi_1 _1474_ (.A1(_0813_),
    .A2(_0976_),
    .Y(_0370_),
    .B1(_0968_));
 sg13g2_xnor2_1 _1475_ (.Y(_0369_),
    .A(\top1.ch2c.data[6] ),
    .B(_0973_));
 sg13g2_xnor2_1 _1476_ (.Y(_0368_),
    .A(\top1.ch2c.data[5] ),
    .B(_0975_));
 sg13g2_xor2_1 _1477_ (.B(_0967_),
    .A(\top1.ch2c.data[4] ),
    .X(_0367_));
 sg13g2_xor2_1 _1478_ (.B(_0972_),
    .A(\top1.ch2c.data[3] ),
    .X(_0366_));
 sg13g2_xnor2_1 _1479_ (.Y(_0365_),
    .A(\top1.ch2c.data[2] ),
    .B(_0971_));
 sg13g2_a21o_1 _1480_ (.A2(net597),
    .A1(\top1.ch2c.data[0] ),
    .B1(\top1.ch2c.data[1] ),
    .X(_0977_));
 sg13g2_and2_1 _1481_ (.A(_0971_),
    .B(_0977_),
    .X(_0364_));
 sg13g2_mux2_1 _1482_ (.A0(_0021_),
    .A1(\top1.ch2c.data[0] ),
    .S(net539),
    .X(_0363_));
 sg13g2_nor2_1 _1483_ (.A(_0853_),
    .B(net541),
    .Y(_0978_));
 sg13g2_nor3_2 _1484_ (.A(_0853_),
    .B(_0856_),
    .C(net541),
    .Y(_0979_));
 sg13g2_and2_1 _1485_ (.A(\top1.ch3c.data[8] ),
    .B(_0979_),
    .X(_0980_));
 sg13g2_nand2_1 _1486_ (.Y(_0981_),
    .A(_0854_),
    .B(_0980_));
 sg13g2_nand3_1 _1487_ (.B(\top1.ch3c.data[0] ),
    .C(net597),
    .A(\top1.ch3c.data[1] ),
    .Y(_0982_));
 sg13g2_nor2_1 _1488_ (.A(_0816_),
    .B(_0982_),
    .Y(_0983_));
 sg13g2_nand4_1 _1489_ (.B(\top1.ch3c.data[4] ),
    .C(\top1.ch3c.data[3] ),
    .A(\top1.ch3c.data[5] ),
    .Y(_0984_),
    .D(_0983_));
 sg13g2_xnor2_1 _1490_ (.Y(_0362_),
    .A(\top1.ch3c.data[11] ),
    .B(_0981_));
 sg13g2_a21oi_1 _1491_ (.A1(\top1.ch3c.data[9] ),
    .A2(_0980_),
    .Y(_0985_),
    .B1(\top1.ch3c.data[10] ));
 sg13g2_a21oi_1 _1492_ (.A1(_0854_),
    .A2(_0980_),
    .Y(_0361_),
    .B1(_0985_));
 sg13g2_xor2_1 _1493_ (.B(_0980_),
    .A(\top1.ch3c.data[9] ),
    .X(_0360_));
 sg13g2_xor2_1 _1494_ (.B(_0979_),
    .A(\top1.ch3c.data[8] ),
    .X(_0359_));
 sg13g2_nand2_1 _1495_ (.Y(_0986_),
    .A(\top1.ch3c.data[4] ),
    .B(_0978_));
 sg13g2_nand4_1 _1496_ (.B(\top1.ch3c.data[5] ),
    .C(\top1.ch3c.data[4] ),
    .A(\top1.ch3c.data[6] ),
    .Y(_0987_),
    .D(_0978_));
 sg13g2_a21oi_1 _1497_ (.A1(_0815_),
    .A2(_0987_),
    .Y(_0358_),
    .B1(_0979_));
 sg13g2_xnor2_1 _1498_ (.Y(_0357_),
    .A(\top1.ch3c.data[6] ),
    .B(_0984_));
 sg13g2_xnor2_1 _1499_ (.Y(_0356_),
    .A(\top1.ch3c.data[5] ),
    .B(_0986_));
 sg13g2_xor2_1 _1500_ (.B(_0978_),
    .A(\top1.ch3c.data[4] ),
    .X(_0355_));
 sg13g2_xor2_1 _1501_ (.B(_0983_),
    .A(\top1.ch3c.data[3] ),
    .X(_0354_));
 sg13g2_xnor2_1 _1502_ (.Y(_0353_),
    .A(\top1.ch3c.data[2] ),
    .B(_0982_));
 sg13g2_a21o_1 _1503_ (.A2(net597),
    .A1(\top1.ch3c.data[0] ),
    .B1(\top1.ch3c.data[1] ),
    .X(_0988_));
 sg13g2_and2_1 _1504_ (.A(_0982_),
    .B(_0988_),
    .X(_0352_));
 sg13g2_mux2_1 _1505_ (.A0(_0022_),
    .A1(\top1.ch3c.data[0] ),
    .S(net539),
    .X(_0351_));
 sg13g2_nor2_1 _1506_ (.A(_0859_),
    .B(net540),
    .Y(_0989_));
 sg13g2_nor3_2 _1507_ (.A(_0859_),
    .B(_0861_),
    .C(net540),
    .Y(_0990_));
 sg13g2_nand4_1 _1508_ (.B(\top1.ch4c.data[9] ),
    .C(\top1.ch4c.data[8] ),
    .A(\top1.ch4c.data[10] ),
    .Y(_0991_),
    .D(_0990_));
 sg13g2_nand3_1 _1509_ (.B(\top1.ch4c.data[0] ),
    .C(net594),
    .A(\top1.ch4c.data[1] ),
    .Y(_0992_));
 sg13g2_nand4_1 _1510_ (.B(\top1.ch4c.data[1] ),
    .C(\top1.ch4c.data[0] ),
    .A(\top1.ch4c.data[2] ),
    .Y(_0993_),
    .D(net594));
 sg13g2_nor2_1 _1511_ (.A(_0817_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_and4_1 _1512_ (.A(\top1.ch4c.data[6] ),
    .B(\top1.ch4c.data[5] ),
    .C(\top1.ch4c.data[4] ),
    .D(_0994_),
    .X(_0995_));
 sg13g2_nand4_1 _1513_ (.B(\top1.ch4c.data[8] ),
    .C(\top1.ch4c.data[7] ),
    .A(\top1.ch4c.data[9] ),
    .Y(_0996_),
    .D(_0995_));
 sg13g2_xnor2_1 _1514_ (.Y(_0350_),
    .A(\top1.ch4c.data[11] ),
    .B(_0991_));
 sg13g2_xnor2_1 _1515_ (.Y(_0349_),
    .A(\top1.ch4c.data[10] ),
    .B(_0996_));
 sg13g2_a21o_1 _1516_ (.A2(_0990_),
    .A1(\top1.ch4c.data[8] ),
    .B1(\top1.ch4c.data[9] ),
    .X(_0997_));
 sg13g2_and2_1 _1517_ (.A(_0996_),
    .B(_0997_),
    .X(_0348_));
 sg13g2_xor2_1 _1518_ (.B(_0990_),
    .A(\top1.ch4c.data[8] ),
    .X(_0347_));
 sg13g2_and2_1 _1519_ (.A(\top1.ch4c.data[4] ),
    .B(_0989_),
    .X(_0998_));
 sg13g2_xor2_1 _1520_ (.B(_0995_),
    .A(\top1.ch4c.data[7] ),
    .X(_0346_));
 sg13g2_a21oi_1 _1521_ (.A1(\top1.ch4c.data[5] ),
    .A2(_0998_),
    .Y(_0999_),
    .B1(\top1.ch4c.data[6] ));
 sg13g2_nor2_1 _1522_ (.A(_0995_),
    .B(_0999_),
    .Y(_0345_));
 sg13g2_xor2_1 _1523_ (.B(_0998_),
    .A(\top1.ch4c.data[5] ),
    .X(_0344_));
 sg13g2_xor2_1 _1524_ (.B(_0989_),
    .A(\top1.ch4c.data[4] ),
    .X(_0343_));
 sg13g2_xnor2_1 _1525_ (.Y(_0342_),
    .A(\top1.ch4c.data[3] ),
    .B(_0993_));
 sg13g2_xnor2_1 _1526_ (.Y(_0341_),
    .A(\top1.ch4c.data[2] ),
    .B(_0992_));
 sg13g2_a21o_1 _1527_ (.A2(net594),
    .A1(\top1.ch4c.data[0] ),
    .B1(\top1.ch4c.data[1] ),
    .X(_1000_));
 sg13g2_and2_1 _1528_ (.A(_0992_),
    .B(_1000_),
    .X(_0340_));
 sg13g2_mux2_1 _1529_ (.A0(_0023_),
    .A1(\top1.ch4c.data[0] ),
    .S(net538),
    .X(_0339_));
 sg13g2_nor2_2 _1530_ (.A(_0864_),
    .B(net538),
    .Y(_1001_));
 sg13g2_nor3_2 _1531_ (.A(_0864_),
    .B(_0866_),
    .C(net538),
    .Y(_1002_));
 sg13g2_and2_1 _1532_ (.A(\top1.ch5c.data[8] ),
    .B(_1002_),
    .X(_1003_));
 sg13g2_nand2_1 _1533_ (.Y(_1004_),
    .A(_0867_),
    .B(_1003_));
 sg13g2_nand3_1 _1534_ (.B(\top1.ch5c.data[0] ),
    .C(net597),
    .A(\top1.ch5c.data[1] ),
    .Y(_1005_));
 sg13g2_nor2_1 _1535_ (.A(_0819_),
    .B(_1005_),
    .Y(_1006_));
 sg13g2_nand4_1 _1536_ (.B(\top1.ch5c.data[4] ),
    .C(\top1.ch5c.data[3] ),
    .A(\top1.ch5c.data[5] ),
    .Y(_1007_),
    .D(_1006_));
 sg13g2_xnor2_1 _1537_ (.Y(_0338_),
    .A(\top1.ch5c.data[11] ),
    .B(_1004_));
 sg13g2_a21oi_1 _1538_ (.A1(\top1.ch5c.data[9] ),
    .A2(_1003_),
    .Y(_1008_),
    .B1(\top1.ch5c.data[10] ));
 sg13g2_a21oi_1 _1539_ (.A1(_0867_),
    .A2(_1003_),
    .Y(_0337_),
    .B1(_1008_));
 sg13g2_xor2_1 _1540_ (.B(_1003_),
    .A(\top1.ch5c.data[9] ),
    .X(_0336_));
 sg13g2_xor2_1 _1541_ (.B(_1002_),
    .A(\top1.ch5c.data[8] ),
    .X(_0335_));
 sg13g2_nand2_1 _1542_ (.Y(_1009_),
    .A(\top1.ch5c.data[4] ),
    .B(_1001_));
 sg13g2_nand4_1 _1543_ (.B(\top1.ch5c.data[5] ),
    .C(\top1.ch5c.data[4] ),
    .A(\top1.ch5c.data[6] ),
    .Y(_1010_),
    .D(_1001_));
 sg13g2_a21oi_1 _1544_ (.A1(_0818_),
    .A2(_1010_),
    .Y(_0334_),
    .B1(_1002_));
 sg13g2_xnor2_1 _1545_ (.Y(_0333_),
    .A(\top1.ch5c.data[6] ),
    .B(_1007_));
 sg13g2_xnor2_1 _1546_ (.Y(_0332_),
    .A(\top1.ch5c.data[5] ),
    .B(_1009_));
 sg13g2_xor2_1 _1547_ (.B(_1001_),
    .A(\top1.ch5c.data[4] ),
    .X(_0331_));
 sg13g2_xor2_1 _1548_ (.B(_1006_),
    .A(\top1.ch5c.data[3] ),
    .X(_0330_));
 sg13g2_xnor2_1 _1549_ (.Y(_0329_),
    .A(\top1.ch5c.data[2] ),
    .B(_1005_));
 sg13g2_a21o_1 _1550_ (.A2(net597),
    .A1(\top1.ch5c.data[0] ),
    .B1(\top1.ch5c.data[1] ),
    .X(_1011_));
 sg13g2_and2_1 _1551_ (.A(_1005_),
    .B(_1011_),
    .X(_0328_));
 sg13g2_mux2_1 _1552_ (.A0(_0024_),
    .A1(\top1.ch5c.data[0] ),
    .S(net536),
    .X(_0327_));
 sg13g2_nor2_1 _1553_ (.A(_0870_),
    .B(net536),
    .Y(_1012_));
 sg13g2_nor3_1 _1554_ (.A(_0870_),
    .B(_0872_),
    .C(net536),
    .Y(_1013_));
 sg13g2_and2_1 _1555_ (.A(\top1.ch6c.data[8] ),
    .B(_1013_),
    .X(_1014_));
 sg13g2_nand2b_1 _1556_ (.Y(_1015_),
    .B(_1014_),
    .A_N(_0871_));
 sg13g2_nand3_1 _1557_ (.B(\top1.ch6c.data[0] ),
    .C(net598),
    .A(\top1.ch6c.data[1] ),
    .Y(_1016_));
 sg13g2_nor2_1 _1558_ (.A(_0821_),
    .B(_1016_),
    .Y(_1017_));
 sg13g2_nand4_1 _1559_ (.B(\top1.ch6c.data[4] ),
    .C(\top1.ch6c.data[3] ),
    .A(\top1.ch6c.data[5] ),
    .Y(_1018_),
    .D(_1017_));
 sg13g2_nor2_1 _1560_ (.A(_0820_),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_xnor2_1 _1561_ (.Y(_0326_),
    .A(\top1.ch6c.data[11] ),
    .B(_1015_));
 sg13g2_a21o_1 _1562_ (.A2(_1014_),
    .A1(\top1.ch6c.data[9] ),
    .B1(\top1.ch6c.data[10] ),
    .X(_1020_));
 sg13g2_and2_1 _1563_ (.A(_1015_),
    .B(_1020_),
    .X(_0325_));
 sg13g2_xor2_1 _1564_ (.B(_1014_),
    .A(\top1.ch6c.data[9] ),
    .X(_0324_));
 sg13g2_xor2_1 _1565_ (.B(_1013_),
    .A(\top1.ch6c.data[8] ),
    .X(_0323_));
 sg13g2_nand2_1 _1566_ (.Y(_1021_),
    .A(\top1.ch6c.data[4] ),
    .B(_1012_));
 sg13g2_xor2_1 _1567_ (.B(_1019_),
    .A(\top1.ch6c.data[7] ),
    .X(_0322_));
 sg13g2_xnor2_1 _1568_ (.Y(_0321_),
    .A(\top1.ch6c.data[6] ),
    .B(_1018_));
 sg13g2_xnor2_1 _1569_ (.Y(_0320_),
    .A(\top1.ch6c.data[5] ),
    .B(_1021_));
 sg13g2_xor2_1 _1570_ (.B(_1012_),
    .A(\top1.ch6c.data[4] ),
    .X(_0319_));
 sg13g2_xor2_1 _1571_ (.B(_1017_),
    .A(\top1.ch6c.data[3] ),
    .X(_0318_));
 sg13g2_xnor2_1 _1572_ (.Y(_0317_),
    .A(\top1.ch6c.data[2] ),
    .B(_1016_));
 sg13g2_a21o_1 _1573_ (.A2(net598),
    .A1(\top1.ch6c.data[0] ),
    .B1(\top1.ch6c.data[1] ),
    .X(_0436_));
 sg13g2_and2_1 _1574_ (.A(_1016_),
    .B(_0436_),
    .X(_0316_));
 sg13g2_mux2_1 _1575_ (.A0(_0025_),
    .A1(\top1.ch6c.data[0] ),
    .S(net537),
    .X(_0315_));
 sg13g2_nor2_1 _1576_ (.A(_0875_),
    .B(net537),
    .Y(_0437_));
 sg13g2_nor3_1 _1577_ (.A(_0875_),
    .B(_0877_),
    .C(net537),
    .Y(_0438_));
 sg13g2_and2_1 _1578_ (.A(\top1.ch7c.data[8] ),
    .B(_0438_),
    .X(_0439_));
 sg13g2_nand2b_1 _1579_ (.Y(_0440_),
    .B(_0439_),
    .A_N(_0876_));
 sg13g2_nand3_1 _1580_ (.B(\top1.ch7c.data[0] ),
    .C(net598),
    .A(\top1.ch7c.data[1] ),
    .Y(_0441_));
 sg13g2_nor2_1 _1581_ (.A(_0823_),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_nand4_1 _1582_ (.B(\top1.ch7c.data[4] ),
    .C(\top1.ch7c.data[3] ),
    .A(\top1.ch7c.data[5] ),
    .Y(_0443_),
    .D(_0442_));
 sg13g2_nor2_1 _1583_ (.A(_0822_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_xnor2_1 _1584_ (.Y(_0314_),
    .A(\top1.ch7c.data[11] ),
    .B(_0440_));
 sg13g2_a21o_1 _1585_ (.A2(_0439_),
    .A1(\top1.ch7c.data[9] ),
    .B1(\top1.ch7c.data[10] ),
    .X(_0445_));
 sg13g2_and2_1 _1586_ (.A(_0440_),
    .B(_0445_),
    .X(_0313_));
 sg13g2_xor2_1 _1587_ (.B(_0439_),
    .A(\top1.ch7c.data[9] ),
    .X(_0312_));
 sg13g2_xor2_1 _1588_ (.B(_0438_),
    .A(\top1.ch7c.data[8] ),
    .X(_0311_));
 sg13g2_nand2_1 _1589_ (.Y(_0446_),
    .A(\top1.ch7c.data[4] ),
    .B(_0437_));
 sg13g2_xor2_1 _1590_ (.B(_0444_),
    .A(\top1.ch7c.data[7] ),
    .X(_0310_));
 sg13g2_xnor2_1 _1591_ (.Y(_0309_),
    .A(\top1.ch7c.data[6] ),
    .B(_0443_));
 sg13g2_xnor2_1 _1592_ (.Y(_0308_),
    .A(\top1.ch7c.data[5] ),
    .B(_0446_));
 sg13g2_xor2_1 _1593_ (.B(_0437_),
    .A(\top1.ch7c.data[4] ),
    .X(_0307_));
 sg13g2_xor2_1 _1594_ (.B(_0442_),
    .A(\top1.ch7c.data[3] ),
    .X(_0306_));
 sg13g2_xnor2_1 _1595_ (.Y(_0305_),
    .A(\top1.ch7c.data[2] ),
    .B(_0441_));
 sg13g2_a21o_1 _1596_ (.A2(net598),
    .A1(\top1.ch7c.data[0] ),
    .B1(\top1.ch7c.data[1] ),
    .X(_0447_));
 sg13g2_and2_1 _1597_ (.A(_0441_),
    .B(_0447_),
    .X(_0304_));
 sg13g2_mux2_1 _1598_ (.A0(_0026_),
    .A1(\top1.ch7c.data[0] ),
    .S(net537),
    .X(_0303_));
 sg13g2_nor2_2 _1599_ (.A(_0884_),
    .B(net535),
    .Y(_0448_));
 sg13g2_nor3_2 _1600_ (.A(_0884_),
    .B(_0885_),
    .C(net535),
    .Y(_0449_));
 sg13g2_and2_1 _1601_ (.A(\top1.ch8c.data[8] ),
    .B(_0449_),
    .X(_0450_));
 sg13g2_nand3_1 _1602_ (.B(\top1.ch8c.data[9] ),
    .C(_0450_),
    .A(\top1.ch8c.data[10] ),
    .Y(_0451_));
 sg13g2_nand3_1 _1603_ (.B(\top1.ch8c.data[0] ),
    .C(net595),
    .A(\top1.ch8c.data[1] ),
    .Y(_0452_));
 sg13g2_nor2_1 _1604_ (.A(_0825_),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_nand4_1 _1605_ (.B(\top1.ch8c.data[4] ),
    .C(\top1.ch8c.data[3] ),
    .A(\top1.ch8c.data[5] ),
    .Y(_0454_),
    .D(_0453_));
 sg13g2_xnor2_1 _1606_ (.Y(_0302_),
    .A(\top1.ch8c.data[11] ),
    .B(_0451_));
 sg13g2_a21o_1 _1607_ (.A2(net595),
    .A1(_0883_),
    .B1(\top1.ch8c.data[10] ),
    .X(_0455_));
 sg13g2_and2_1 _1608_ (.A(_0451_),
    .B(_0455_),
    .X(_0301_));
 sg13g2_xor2_1 _1609_ (.B(_0450_),
    .A(\top1.ch8c.data[9] ),
    .X(_0300_));
 sg13g2_xor2_1 _1610_ (.B(_0449_),
    .A(\top1.ch8c.data[8] ),
    .X(_0299_));
 sg13g2_nand2_1 _1611_ (.Y(_0456_),
    .A(\top1.ch8c.data[4] ),
    .B(_0448_));
 sg13g2_nand4_1 _1612_ (.B(\top1.ch8c.data[5] ),
    .C(\top1.ch8c.data[4] ),
    .A(\top1.ch8c.data[6] ),
    .Y(_0457_),
    .D(_0448_));
 sg13g2_a21oi_1 _1613_ (.A1(_0824_),
    .A2(_0457_),
    .Y(_0298_),
    .B1(_0449_));
 sg13g2_xnor2_1 _1614_ (.Y(_0297_),
    .A(\top1.ch8c.data[6] ),
    .B(_0454_));
 sg13g2_xnor2_1 _1615_ (.Y(_0296_),
    .A(\top1.ch8c.data[5] ),
    .B(_0456_));
 sg13g2_xor2_1 _1616_ (.B(_0448_),
    .A(\top1.ch8c.data[4] ),
    .X(_0295_));
 sg13g2_xor2_1 _1617_ (.B(_0453_),
    .A(\top1.ch8c.data[3] ),
    .X(_0294_));
 sg13g2_xnor2_1 _1618_ (.Y(_0293_),
    .A(\top1.ch8c.data[2] ),
    .B(_0452_));
 sg13g2_a21o_1 _1619_ (.A2(net595),
    .A1(\top1.ch8c.data[0] ),
    .B1(\top1.ch8c.data[1] ),
    .X(_0458_));
 sg13g2_and2_1 _1620_ (.A(_0452_),
    .B(_0458_),
    .X(_0292_));
 sg13g2_mux2_1 _1621_ (.A0(_0027_),
    .A1(\top1.ch8c.data[0] ),
    .S(net535),
    .X(_0291_));
 sg13g2_nor2_1 _1622_ (.A(_0893_),
    .B(net536),
    .Y(_0459_));
 sg13g2_nor3_2 _1623_ (.A(_0893_),
    .B(_0895_),
    .C(net536),
    .Y(_0460_));
 sg13g2_and2_1 _1624_ (.A(\top1.ch10c.data[8] ),
    .B(_0460_),
    .X(_0461_));
 sg13g2_nand2_1 _1625_ (.Y(_0462_),
    .A(_0896_),
    .B(_0461_));
 sg13g2_nand3_1 _1626_ (.B(\top1.ch10c.data[0] ),
    .C(net595),
    .A(\top1.ch10c.data[1] ),
    .Y(_0463_));
 sg13g2_nor2_1 _1627_ (.A(_0827_),
    .B(_0463_),
    .Y(_0464_));
 sg13g2_nand4_1 _1628_ (.B(\top1.ch10c.data[4] ),
    .C(\top1.ch10c.data[3] ),
    .A(\top1.ch10c.data[5] ),
    .Y(_0465_),
    .D(_0464_));
 sg13g2_xnor2_1 _1629_ (.Y(_0289_),
    .A(\top1.ch10c.data[11] ),
    .B(_0462_));
 sg13g2_a21oi_1 _1630_ (.A1(\top1.ch10c.data[9] ),
    .A2(_0461_),
    .Y(_0466_),
    .B1(\top1.ch10c.data[10] ));
 sg13g2_a21oi_1 _1631_ (.A1(_0896_),
    .A2(_0461_),
    .Y(_0288_),
    .B1(_0466_));
 sg13g2_xor2_1 _1632_ (.B(_0461_),
    .A(\top1.ch10c.data[9] ),
    .X(_0287_));
 sg13g2_xor2_1 _1633_ (.B(_0460_),
    .A(\top1.ch10c.data[8] ),
    .X(_0286_));
 sg13g2_nand2_1 _1634_ (.Y(_0467_),
    .A(\top1.ch10c.data[4] ),
    .B(_0459_));
 sg13g2_nand4_1 _1635_ (.B(\top1.ch10c.data[5] ),
    .C(\top1.ch10c.data[4] ),
    .A(\top1.ch10c.data[6] ),
    .Y(_0468_),
    .D(_0459_));
 sg13g2_a21oi_1 _1636_ (.A1(_0826_),
    .A2(_0468_),
    .Y(_0285_),
    .B1(_0460_));
 sg13g2_xnor2_1 _1637_ (.Y(_0284_),
    .A(\top1.ch10c.data[6] ),
    .B(_0465_));
 sg13g2_xnor2_1 _1638_ (.Y(_0283_),
    .A(\top1.ch10c.data[5] ),
    .B(_0467_));
 sg13g2_xor2_1 _1639_ (.B(_0459_),
    .A(\top1.ch10c.data[4] ),
    .X(_0282_));
 sg13g2_xor2_1 _1640_ (.B(_0464_),
    .A(\top1.ch10c.data[3] ),
    .X(_0281_));
 sg13g2_xnor2_1 _1641_ (.Y(_0280_),
    .A(\top1.ch10c.data[2] ),
    .B(_0463_));
 sg13g2_a21o_1 _1642_ (.A2(net595),
    .A1(\top1.ch10c.data[0] ),
    .B1(\top1.ch10c.data[1] ),
    .X(_0469_));
 sg13g2_and2_1 _1643_ (.A(_0463_),
    .B(_0469_),
    .X(_0279_));
 sg13g2_mux2_1 _1644_ (.A0(_0028_),
    .A1(\top1.ch10c.data[0] ),
    .S(net538),
    .X(_0278_));
 sg13g2_nor2_1 _1645_ (.A(_0899_),
    .B(net536),
    .Y(_0470_));
 sg13g2_nor3_2 _1646_ (.A(_0899_),
    .B(_0901_),
    .C(net536),
    .Y(_0471_));
 sg13g2_and2_1 _1647_ (.A(\top1.ch11c.data[8] ),
    .B(_0471_),
    .X(_0472_));
 sg13g2_nand2_1 _1648_ (.Y(_0473_),
    .A(_0902_),
    .B(_0472_));
 sg13g2_nand3_1 _1649_ (.B(\top1.ch11c.data[0] ),
    .C(net598),
    .A(\top1.ch11c.data[1] ),
    .Y(_0474_));
 sg13g2_nor2_1 _1650_ (.A(_0829_),
    .B(_0474_),
    .Y(_0475_));
 sg13g2_nand4_1 _1651_ (.B(\top1.ch11c.data[4] ),
    .C(\top1.ch11c.data[3] ),
    .A(\top1.ch11c.data[5] ),
    .Y(_0476_),
    .D(_0475_));
 sg13g2_xnor2_1 _1652_ (.Y(_0277_),
    .A(\top1.ch11c.data[11] ),
    .B(_0473_));
 sg13g2_a21oi_1 _1653_ (.A1(\top1.ch11c.data[9] ),
    .A2(_0472_),
    .Y(_0477_),
    .B1(\top1.ch11c.data[10] ));
 sg13g2_a21oi_1 _1654_ (.A1(_0902_),
    .A2(_0472_),
    .Y(_0276_),
    .B1(_0477_));
 sg13g2_xor2_1 _1655_ (.B(_0472_),
    .A(\top1.ch11c.data[9] ),
    .X(_0275_));
 sg13g2_xor2_1 _1656_ (.B(_0471_),
    .A(\top1.ch11c.data[8] ),
    .X(_0274_));
 sg13g2_nand2_1 _1657_ (.Y(_0478_),
    .A(\top1.ch11c.data[4] ),
    .B(_0470_));
 sg13g2_nand4_1 _1658_ (.B(\top1.ch11c.data[5] ),
    .C(\top1.ch11c.data[4] ),
    .A(\top1.ch11c.data[6] ),
    .Y(_0479_),
    .D(_0470_));
 sg13g2_a21oi_1 _1659_ (.A1(_0828_),
    .A2(_0479_),
    .Y(_0273_),
    .B1(_0471_));
 sg13g2_xnor2_1 _1660_ (.Y(_0272_),
    .A(\top1.ch11c.data[6] ),
    .B(_0476_));
 sg13g2_xnor2_1 _1661_ (.Y(_0271_),
    .A(\top1.ch11c.data[5] ),
    .B(_0478_));
 sg13g2_xor2_1 _1662_ (.B(_0470_),
    .A(\top1.ch11c.data[4] ),
    .X(_0270_));
 sg13g2_xor2_1 _1663_ (.B(_0475_),
    .A(\top1.ch11c.data[3] ),
    .X(_0269_));
 sg13g2_xnor2_1 _1664_ (.Y(_0268_),
    .A(\top1.ch11c.data[2] ),
    .B(_0474_));
 sg13g2_a21o_1 _1665_ (.A2(net598),
    .A1(\top1.ch11c.data[0] ),
    .B1(\top1.ch11c.data[1] ),
    .X(_0480_));
 sg13g2_and2_1 _1666_ (.A(_0474_),
    .B(_0480_),
    .X(_0267_));
 sg13g2_mux2_1 _1667_ (.A0(_0029_),
    .A1(\top1.ch11c.data[0] ),
    .S(net536),
    .X(_0266_));
 sg13g2_nor2_1 _1668_ (.A(_0905_),
    .B(net538),
    .Y(_0481_));
 sg13g2_nor3_2 _1669_ (.A(_0905_),
    .B(_0908_),
    .C(net535),
    .Y(_0482_));
 sg13g2_and2_1 _1670_ (.A(\top1.ch12c.data[8] ),
    .B(_0482_),
    .X(_0483_));
 sg13g2_nand2_1 _1671_ (.Y(_0484_),
    .A(_0906_),
    .B(_0483_));
 sg13g2_nand3_1 _1672_ (.B(\top1.ch12c.data[0] ),
    .C(net594),
    .A(\top1.ch12c.data[1] ),
    .Y(_0485_));
 sg13g2_nor2_1 _1673_ (.A(_0831_),
    .B(_0485_),
    .Y(_0486_));
 sg13g2_nand4_1 _1674_ (.B(\top1.ch12c.data[4] ),
    .C(\top1.ch12c.data[3] ),
    .A(\top1.ch12c.data[5] ),
    .Y(_0487_),
    .D(_0486_));
 sg13g2_xnor2_1 _1675_ (.Y(_0265_),
    .A(\top1.ch12c.data[11] ),
    .B(_0484_));
 sg13g2_a21oi_1 _1676_ (.A1(\top1.ch12c.data[9] ),
    .A2(_0483_),
    .Y(_0488_),
    .B1(\top1.ch12c.data[10] ));
 sg13g2_a21oi_1 _1677_ (.A1(_0906_),
    .A2(_0483_),
    .Y(_0264_),
    .B1(_0488_));
 sg13g2_xor2_1 _1678_ (.B(_0483_),
    .A(\top1.ch12c.data[9] ),
    .X(_0263_));
 sg13g2_xor2_1 _1679_ (.B(_0482_),
    .A(\top1.ch12c.data[8] ),
    .X(_0262_));
 sg13g2_nand2_1 _1680_ (.Y(_0489_),
    .A(\top1.ch12c.data[4] ),
    .B(_0481_));
 sg13g2_nand4_1 _1681_ (.B(\top1.ch12c.data[5] ),
    .C(\top1.ch12c.data[4] ),
    .A(\top1.ch12c.data[6] ),
    .Y(_0490_),
    .D(_0481_));
 sg13g2_a21oi_1 _1682_ (.A1(_0830_),
    .A2(_0490_),
    .Y(_0261_),
    .B1(_0482_));
 sg13g2_xnor2_1 _1683_ (.Y(_0260_),
    .A(\top1.ch12c.data[6] ),
    .B(_0487_));
 sg13g2_xnor2_1 _1684_ (.Y(_0259_),
    .A(\top1.ch12c.data[5] ),
    .B(_0489_));
 sg13g2_xor2_1 _1685_ (.B(_0481_),
    .A(\top1.ch12c.data[4] ),
    .X(_0258_));
 sg13g2_xor2_1 _1686_ (.B(_0486_),
    .A(\top1.ch12c.data[3] ),
    .X(_0257_));
 sg13g2_xnor2_1 _1687_ (.Y(_0256_),
    .A(\top1.ch12c.data[2] ),
    .B(_0485_));
 sg13g2_a21o_1 _1688_ (.A2(net594),
    .A1(\top1.ch12c.data[0] ),
    .B1(\top1.ch12c.data[1] ),
    .X(_0491_));
 sg13g2_and2_1 _1689_ (.A(_0485_),
    .B(_0491_),
    .X(_0255_));
 sg13g2_mux2_1 _1690_ (.A0(_0030_),
    .A1(\top1.ch12c.data[0] ),
    .S(net535),
    .X(_0254_));
 sg13g2_nor2_2 _1691_ (.A(_0911_),
    .B(net540),
    .Y(_0492_));
 sg13g2_nor3_2 _1692_ (.A(_0911_),
    .B(_0914_),
    .C(net540),
    .Y(_0493_));
 sg13g2_and2_1 _1693_ (.A(\top1.ch13c.data[8] ),
    .B(_0493_),
    .X(_0494_));
 sg13g2_nand2_1 _1694_ (.Y(_0495_),
    .A(_0912_),
    .B(_0494_));
 sg13g2_nand3_1 _1695_ (.B(\top1.ch13c.data[0] ),
    .C(net596),
    .A(\top1.ch13c.data[1] ),
    .Y(_0496_));
 sg13g2_nor2_1 _1696_ (.A(_0833_),
    .B(_0496_),
    .Y(_0497_));
 sg13g2_nand4_1 _1697_ (.B(\top1.ch13c.data[4] ),
    .C(\top1.ch13c.data[3] ),
    .A(\top1.ch13c.data[5] ),
    .Y(_0498_),
    .D(_0497_));
 sg13g2_xnor2_1 _1698_ (.Y(_0253_),
    .A(\top1.ch13c.data[11] ),
    .B(_0495_));
 sg13g2_a21oi_1 _1699_ (.A1(\top1.ch13c.data[9] ),
    .A2(_0494_),
    .Y(_0499_),
    .B1(\top1.ch13c.data[10] ));
 sg13g2_a21oi_1 _1700_ (.A1(_0912_),
    .A2(_0494_),
    .Y(_0252_),
    .B1(_0499_));
 sg13g2_xor2_1 _1701_ (.B(_0494_),
    .A(\top1.ch13c.data[9] ),
    .X(_0251_));
 sg13g2_xor2_1 _1702_ (.B(_0493_),
    .A(\top1.ch13c.data[8] ),
    .X(_0250_));
 sg13g2_nand2_1 _1703_ (.Y(_0500_),
    .A(\top1.ch13c.data[4] ),
    .B(_0492_));
 sg13g2_nand4_1 _1704_ (.B(\top1.ch13c.data[5] ),
    .C(\top1.ch13c.data[4] ),
    .A(\top1.ch13c.data[6] ),
    .Y(_0501_),
    .D(_0492_));
 sg13g2_a21oi_1 _1705_ (.A1(_0832_),
    .A2(_0501_),
    .Y(_0249_),
    .B1(_0493_));
 sg13g2_xnor2_1 _1706_ (.Y(_0248_),
    .A(\top1.ch13c.data[6] ),
    .B(_0498_));
 sg13g2_xnor2_1 _1707_ (.Y(_0247_),
    .A(\top1.ch13c.data[5] ),
    .B(_0500_));
 sg13g2_xor2_1 _1708_ (.B(_0492_),
    .A(\top1.ch13c.data[4] ),
    .X(_0246_));
 sg13g2_xor2_1 _1709_ (.B(_0497_),
    .A(\top1.ch13c.data[3] ),
    .X(_0245_));
 sg13g2_xnor2_1 _1710_ (.Y(_0244_),
    .A(\top1.ch13c.data[2] ),
    .B(_0496_));
 sg13g2_a21o_1 _1711_ (.A2(net596),
    .A1(\top1.ch13c.data[0] ),
    .B1(\top1.ch13c.data[1] ),
    .X(_0502_));
 sg13g2_and2_1 _1712_ (.A(_0496_),
    .B(_0502_),
    .X(_0243_));
 sg13g2_mux2_1 _1713_ (.A0(_0031_),
    .A1(\top1.ch13c.data[0] ),
    .S(net540),
    .X(_0242_));
 sg13g2_nor2_1 _1714_ (.A(_0917_),
    .B(net535),
    .Y(_0503_));
 sg13g2_nor3_2 _1715_ (.A(_0917_),
    .B(_0920_),
    .C(net540),
    .Y(_0504_));
 sg13g2_and2_1 _1716_ (.A(\top1.ch14c.data[8] ),
    .B(_0504_),
    .X(_0505_));
 sg13g2_nand2_1 _1717_ (.Y(_0506_),
    .A(_0918_),
    .B(_0505_));
 sg13g2_nand3_1 _1718_ (.B(\top1.ch14c.data[0] ),
    .C(net594),
    .A(\top1.ch14c.data[1] ),
    .Y(_0507_));
 sg13g2_nor2_1 _1719_ (.A(_0835_),
    .B(_0507_),
    .Y(_0508_));
 sg13g2_nand4_1 _1720_ (.B(\top1.ch14c.data[4] ),
    .C(\top1.ch14c.data[3] ),
    .A(\top1.ch14c.data[5] ),
    .Y(_0509_),
    .D(_0508_));
 sg13g2_xnor2_1 _1721_ (.Y(_0241_),
    .A(\top1.ch14c.data[11] ),
    .B(_0506_));
 sg13g2_a21oi_1 _1722_ (.A1(\top1.ch14c.data[9] ),
    .A2(_0505_),
    .Y(_0510_),
    .B1(\top1.ch14c.data[10] ));
 sg13g2_a21oi_1 _1723_ (.A1(_0918_),
    .A2(_0505_),
    .Y(_0240_),
    .B1(_0510_));
 sg13g2_xor2_1 _1724_ (.B(_0505_),
    .A(\top1.ch14c.data[9] ),
    .X(_0239_));
 sg13g2_xor2_1 _1725_ (.B(_0504_),
    .A(\top1.ch14c.data[8] ),
    .X(_0238_));
 sg13g2_nand2_1 _1726_ (.Y(_0511_),
    .A(\top1.ch14c.data[4] ),
    .B(_0503_));
 sg13g2_nand4_1 _1727_ (.B(\top1.ch14c.data[5] ),
    .C(\top1.ch14c.data[4] ),
    .A(\top1.ch14c.data[6] ),
    .Y(_0512_),
    .D(_0503_));
 sg13g2_a21oi_1 _1728_ (.A1(_0834_),
    .A2(_0512_),
    .Y(_0237_),
    .B1(_0504_));
 sg13g2_xnor2_1 _1729_ (.Y(_0236_),
    .A(\top1.ch14c.data[6] ),
    .B(_0509_));
 sg13g2_xnor2_1 _1730_ (.Y(_0235_),
    .A(\top1.ch14c.data[5] ),
    .B(_0511_));
 sg13g2_xor2_1 _1731_ (.B(_0503_),
    .A(\top1.ch14c.data[4] ),
    .X(_0234_));
 sg13g2_xor2_1 _1732_ (.B(_0508_),
    .A(\top1.ch14c.data[3] ),
    .X(_0233_));
 sg13g2_xnor2_1 _1733_ (.Y(_0232_),
    .A(\top1.ch14c.data[2] ),
    .B(_0507_));
 sg13g2_a21o_1 _1734_ (.A2(net594),
    .A1(\top1.ch14c.data[0] ),
    .B1(\top1.ch14c.data[1] ),
    .X(_0513_));
 sg13g2_and2_1 _1735_ (.A(_0507_),
    .B(_0513_),
    .X(_0231_));
 sg13g2_mux2_1 _1736_ (.A0(_0032_),
    .A1(\top1.ch14c.data[0] ),
    .S(net535),
    .X(_0230_));
 sg13g2_and2_1 _1737_ (.A(\top1.data[0][1] ),
    .B(\top1.data[0][0] ),
    .X(_0514_));
 sg13g2_nand4_1 _1738_ (.B(\top1.data[0][4] ),
    .C(\top1.data[0][5] ),
    .A(\top1.data[0][3] ),
    .Y(_0515_),
    .D(_0514_));
 sg13g2_nor2_2 _1739_ (.A(\top1.data[0][2] ),
    .B(_0515_),
    .Y(_0516_));
 sg13g2_and3_1 _1740_ (.X(_0517_),
    .A(\top1.data[0][7] ),
    .B(\top1.data[0][6] ),
    .C(_0516_));
 sg13g2_and4_1 _1741_ (.A(\top1.data[0][9] ),
    .B(\top1.data[0][10] ),
    .C(\top1.data[0][11] ),
    .D(_0517_),
    .X(_0518_));
 sg13g2_nor2b_1 _1742_ (.A(\top1.data[0][8] ),
    .B_N(_0518_),
    .Y(_0519_));
 sg13g2_or2_1 _1743_ (.X(_0229_),
    .B(_0519_),
    .A(\top1.ovf_RTC ));
 sg13g2_nor2_1 _1744_ (.A(net607),
    .B(net604),
    .Y(_0520_));
 sg13g2_or2_1 _1745_ (.X(_0521_),
    .B(\top1.FSM1.state_reg[3] ),
    .A(net602));
 sg13g2_nor4_2 _1746_ (.A(net607),
    .B(net604),
    .C(net602),
    .Y(_0522_),
    .D(net601));
 sg13g2_or4_2 _1747_ (.A(net607),
    .B(net604),
    .C(net602),
    .D(net601),
    .X(_0523_));
 sg13g2_nand2_1 _1748_ (.Y(_0524_),
    .A(\top1.FSM1.state_reg[4] ),
    .B(_0523_));
 sg13g2_nand2_2 _1749_ (.Y(_0525_),
    .A(net602),
    .B(net601));
 sg13g2_and2_1 _1750_ (.A(net606),
    .B(net604),
    .X(_0526_));
 sg13g2_and4_1 _1751_ (.A(net606),
    .B(net604),
    .C(net602),
    .D(net601),
    .X(_0527_));
 sg13g2_nand4_1 _1752_ (.B(net604),
    .C(net602),
    .A(net607),
    .Y(_0528_),
    .D(net601));
 sg13g2_mux2_1 _1753_ (.A0(_0522_),
    .A1(_0527_),
    .S(_0837_),
    .X(_0529_));
 sg13g2_mux2_2 _1754_ (.A0(_0523_),
    .A1(_0528_),
    .S(_0837_),
    .X(_0530_));
 sg13g2_o21ai_1 _1755_ (.B1(net600),
    .Y(_0531_),
    .A1(net606),
    .A2(net604));
 sg13g2_nor2_1 _1756_ (.A(_0526_),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_nor3_1 _1757_ (.A(_0525_),
    .B(_0526_),
    .C(_0531_),
    .Y(_0533_));
 sg13g2_or3_1 _1758_ (.A(_0525_),
    .B(_0526_),
    .C(_0531_),
    .X(_0534_));
 sg13g2_nor2_1 _1759_ (.A(_0529_),
    .B(_0533_),
    .Y(_0535_));
 sg13g2_nand2_1 _1760_ (.Y(_0536_),
    .A(_0530_),
    .B(_0534_));
 sg13g2_and2_1 _1761_ (.A(net600),
    .B(_0520_),
    .X(_0537_));
 sg13g2_and3_1 _1762_ (.X(_0538_),
    .A(net603),
    .B(net600),
    .C(_0520_));
 sg13g2_nand3_1 _1763_ (.B(net600),
    .C(_0520_),
    .A(net602),
    .Y(_0539_));
 sg13g2_nor4_1 _1764_ (.A(net606),
    .B(net605),
    .C(_0838_),
    .D(_0525_),
    .Y(_0540_));
 sg13g2_nand2b_1 _1765_ (.Y(_0541_),
    .B(net601),
    .A_N(net603));
 sg13g2_nor2_1 _1766_ (.A(_0531_),
    .B(_0541_),
    .Y(_0542_));
 sg13g2_nand3_1 _1767_ (.B(net605),
    .C(net600),
    .A(net606),
    .Y(_0543_));
 sg13g2_nor2_1 _1768_ (.A(net603),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_o21ai_1 _1769_ (.B1(_0539_),
    .Y(_0545_),
    .A1(net602),
    .A2(_0531_));
 sg13g2_nor2_1 _1770_ (.A(net593),
    .B(_0542_),
    .Y(_0546_));
 sg13g2_or2_1 _1771_ (.X(_0547_),
    .B(_0542_),
    .A(net593));
 sg13g2_nand2_1 _1772_ (.Y(\top1.a3_out ),
    .A(_0535_),
    .B(_0546_));
 sg13g2_nand2b_2 _1773_ (.Y(_0548_),
    .B(net603),
    .A_N(net601));
 sg13g2_nor3_1 _1774_ (.A(_0526_),
    .B(_0531_),
    .C(_0548_),
    .Y(_0549_));
 sg13g2_or3_1 _1775_ (.A(_0526_),
    .B(_0531_),
    .C(_0548_),
    .X(_0550_));
 sg13g2_nor4_1 _1776_ (.A(net606),
    .B(net605),
    .C(_0838_),
    .D(_0541_),
    .Y(_0551_));
 sg13g2_nor2_1 _1777_ (.A(_0543_),
    .B(_0548_),
    .Y(_0552_));
 sg13g2_or3_1 _1778_ (.A(_0549_),
    .B(net590),
    .C(net588),
    .X(_0553_));
 sg13g2_or2_1 _1779_ (.X(\top1.a2_out ),
    .B(_0553_),
    .A(_0536_));
 sg13g2_nor4_2 _1780_ (.A(_0538_),
    .B(_0544_),
    .C(net590),
    .Y(_0554_),
    .D(net588));
 sg13g2_and2_1 _1781_ (.A(_0530_),
    .B(_0554_),
    .X(_0555_));
 sg13g2_inv_1 _1782_ (.Y(\top1.a1_out ),
    .A(_0555_));
 sg13g2_nand2b_1 _1783_ (.Y(_0556_),
    .B(net604),
    .A_N(net606));
 sg13g2_o21ai_1 _1784_ (.B1(_0837_),
    .Y(_0557_),
    .A1(_0525_),
    .A2(_0556_));
 sg13g2_nand3b_1 _1785_ (.B(net605),
    .C(net600),
    .Y(_0558_),
    .A_N(net606));
 sg13g2_nor2b_1 _1786_ (.A(_0558_),
    .B_N(_0525_),
    .Y(_0559_));
 sg13g2_nand2_1 _1787_ (.Y(_0560_),
    .A(_0521_),
    .B(_0537_));
 sg13g2_nand2_1 _1788_ (.Y(_0561_),
    .A(_0558_),
    .B(_0560_));
 sg13g2_a221oi_1 _1789_ (.B2(_0524_),
    .C1(_0559_),
    .B1(_0557_),
    .A1(_0521_),
    .Y(_0562_),
    .A2(_0537_));
 sg13g2_a21o_1 _1790_ (.A2(_0535_),
    .A1(_0838_),
    .B1(_0562_),
    .X(_0563_));
 sg13g2_inv_1 _1791_ (.Y(\top1.a0_out ),
    .A(net532));
 sg13g2_nor3_1 _1792_ (.A(_0536_),
    .B(_0547_),
    .C(_0553_),
    .Y(_0564_));
 sg13g2_or3_2 _1793_ (.A(_0536_),
    .B(_0545_),
    .C(_0553_),
    .X(_0565_));
 sg13g2_nor4_1 _1794_ (.A(\top1.FSM1.counter_register[1] ),
    .B(\top1.FSM1.counter_register[0] ),
    .C(\top1.FSM1.counter_register[3] ),
    .D(\top1.FSM1.counter_register[2] ),
    .Y(_0566_));
 sg13g2_nand2_1 _1795_ (.Y(_0567_),
    .A(_0565_),
    .B(_0566_));
 sg13g2_inv_1 _1796_ (.Y(\top1.FSM1.SL ),
    .A(net520));
 sg13g2_nand2_1 _1797_ (.Y(_0568_),
    .A(net34),
    .B(net520));
 sg13g2_nand3_1 _1798_ (.B(net532),
    .C(_0564_),
    .A(_0555_),
    .Y(_0569_));
 sg13g2_nor2_1 _1799_ (.A(_0530_),
    .B(_0562_),
    .Y(_0570_));
 sg13g2_nand2_1 _1800_ (.Y(_0571_),
    .A(\top1.ch15c.data[1] ),
    .B(net528));
 sg13g2_and2_1 _1801_ (.A(_0529_),
    .B(_0562_),
    .X(_0572_));
 sg13g2_and2_1 _1802_ (.A(_0533_),
    .B(_0562_),
    .X(_0573_));
 sg13g2_a22oi_1 _1803_ (.Y(_0574_),
    .B1(net524),
    .B2(\top1.ch12c.data[1] ),
    .A2(net526),
    .A1(\top1.ch14c.data[1] ));
 sg13g2_and3_1 _1804_ (.X(_0575_),
    .A(net516),
    .B(_0571_),
    .C(_0574_));
 sg13g2_and3_1 _1805_ (.X(_0576_),
    .A(_0553_),
    .B(_0555_),
    .C(net532));
 sg13g2_nand2_1 _1806_ (.Y(_0577_),
    .A(\top1.ch4c.data[1] ),
    .B(net513));
 sg13g2_and3_1 _1807_ (.X(_0578_),
    .A(_0547_),
    .B(_0555_),
    .C(net532));
 sg13g2_nand2_1 _1808_ (.Y(_0579_),
    .A(\top1.ch8c.data[1] ),
    .B(net511));
 sg13g2_nor2_1 _1809_ (.A(_0534_),
    .B(_0562_),
    .Y(_0580_));
 sg13g2_a21oi_2 _1810_ (.B1(_0546_),
    .Y(_0581_),
    .A2(_0554_),
    .A1(_0530_));
 sg13g2_and2_1 _1811_ (.A(net530),
    .B(net521),
    .X(_0582_));
 sg13g2_nor2_1 _1812_ (.A(_0541_),
    .B(_0558_),
    .Y(_0583_));
 sg13g2_and2_1 _1813_ (.A(\top1.ch9c.data[1] ),
    .B(net585),
    .X(_0584_));
 sg13g2_nor2_1 _1814_ (.A(_0548_),
    .B(_0558_),
    .Y(_0585_));
 sg13g2_nand2_1 _1815_ (.Y(_0586_),
    .A(\top1.ch11c.data[1] ),
    .B(net591));
 sg13g2_nor2_1 _1816_ (.A(_0521_),
    .B(_0558_),
    .Y(_0587_));
 sg13g2_nor2_1 _1817_ (.A(net601),
    .B(_0539_),
    .Y(_0588_));
 sg13g2_nor2_1 _1818_ (.A(_0521_),
    .B(_0543_),
    .Y(_0589_));
 sg13g2_a221oi_1 _1819_ (.B2(\top1.ch3c.data[1] ),
    .C1(_0584_),
    .B1(net533),
    .A1(\top1.ch7c.data[1] ),
    .Y(_0590_),
    .A2(net590));
 sg13g2_a22oi_1 _1820_ (.Y(_0591_),
    .B1(net581),
    .B2(\top1.ch1c.data[1] ),
    .A2(net583),
    .A1(\top1.ch5c.data[1] ));
 sg13g2_a22oi_1 _1821_ (.Y(_0592_),
    .B1(net579),
    .B2(\top1.ch2c.data[1] ),
    .A2(net587),
    .A1(\top1.ch6c.data[1] ));
 sg13g2_nand4_1 _1822_ (.B(_0590_),
    .C(_0591_),
    .A(_0586_),
    .Y(_0593_),
    .D(_0592_));
 sg13g2_a221oi_1 _1823_ (.B2(\top1.ch10c.data[1] ),
    .C1(_0593_),
    .B1(_0582_),
    .A1(\top1.ch13c.data[1] ),
    .Y(_0594_),
    .A2(net523));
 sg13g2_and4_2 _1824_ (.A(_0575_),
    .B(_0577_),
    .C(_0579_),
    .D(_0594_),
    .X(_0595_));
 sg13g2_o21ai_1 _1825_ (.B1(net509),
    .Y(_0596_),
    .A1(\top1.data[0][1] ),
    .A2(net517));
 sg13g2_o21ai_1 _1826_ (.B1(_0568_),
    .Y(_0000_),
    .A1(_0595_),
    .A2(_0596_));
 sg13g2_a22oi_1 _1827_ (.Y(_0597_),
    .B1(net522),
    .B2(\top1.ch13c.data[2] ),
    .A2(net526),
    .A1(\top1.ch14c.data[2] ));
 sg13g2_a22oi_1 _1828_ (.Y(_0598_),
    .B1(net524),
    .B2(\top1.ch12c.data[2] ),
    .A2(net528),
    .A1(\top1.ch15c.data[2] ));
 sg13g2_nand2_1 _1829_ (.Y(_0599_),
    .A(_0597_),
    .B(_0598_));
 sg13g2_and2_1 _1830_ (.A(\top1.ch4c.data[2] ),
    .B(net513),
    .X(_0600_));
 sg13g2_and2_1 _1831_ (.A(\top1.ch8c.data[2] ),
    .B(net511),
    .X(_0601_));
 sg13g2_nand3_1 _1832_ (.B(net530),
    .C(net521),
    .A(\top1.ch10c.data[2] ),
    .Y(_0602_));
 sg13g2_nand2_1 _1833_ (.Y(_0603_),
    .A(\top1.ch1c.data[2] ),
    .B(net581));
 sg13g2_nand2_1 _1834_ (.Y(_0604_),
    .A(\top1.ch11c.data[2] ),
    .B(net591));
 sg13g2_a22oi_1 _1835_ (.Y(_0605_),
    .B1(net584),
    .B2(\top1.ch9c.data[2] ),
    .A2(net590),
    .A1(\top1.ch7c.data[2] ));
 sg13g2_a22oi_1 _1836_ (.Y(_0606_),
    .B1(net582),
    .B2(\top1.ch5c.data[2] ),
    .A2(net586),
    .A1(\top1.ch6c.data[2] ));
 sg13g2_nand4_1 _1837_ (.B(_0604_),
    .C(_0605_),
    .A(_0603_),
    .Y(_0607_),
    .D(_0606_));
 sg13g2_a221oi_1 _1838_ (.B2(\top1.ch2c.data[2] ),
    .C1(_0607_),
    .B1(net578),
    .A1(\top1.ch3c.data[2] ),
    .Y(_0608_),
    .A2(net534));
 sg13g2_nand3_1 _1839_ (.B(_0602_),
    .C(_0608_),
    .A(net515),
    .Y(_0609_));
 sg13g2_nor4_2 _1840_ (.A(_0599_),
    .B(_0600_),
    .C(_0601_),
    .Y(_0610_),
    .D(_0609_));
 sg13g2_o21ai_1 _1841_ (.B1(net509),
    .Y(_0611_),
    .A1(\top1.data[0][2] ),
    .A2(net517));
 sg13g2_nand2_1 _1842_ (.Y(_0612_),
    .A(net36),
    .B(net519));
 sg13g2_o21ai_1 _1843_ (.B1(_0612_),
    .Y(_0001_),
    .A1(_0610_),
    .A2(_0611_));
 sg13g2_a22oi_1 _1844_ (.Y(_0613_),
    .B1(net522),
    .B2(\top1.ch13c.data[3] ),
    .A2(net526),
    .A1(\top1.ch14c.data[3] ));
 sg13g2_a22oi_1 _1845_ (.Y(_0614_),
    .B1(net524),
    .B2(\top1.ch12c.data[3] ),
    .A2(net528),
    .A1(\top1.ch15c.data[3] ));
 sg13g2_nand2_1 _1846_ (.Y(_0615_),
    .A(_0613_),
    .B(_0614_));
 sg13g2_and2_1 _1847_ (.A(\top1.ch8c.data[3] ),
    .B(net511),
    .X(_0616_));
 sg13g2_and2_1 _1848_ (.A(\top1.ch4c.data[3] ),
    .B(net513),
    .X(_0617_));
 sg13g2_nand3_1 _1849_ (.B(net530),
    .C(net521),
    .A(\top1.ch10c.data[3] ),
    .Y(_0618_));
 sg13g2_nand2_2 _1850_ (.Y(_0619_),
    .A(\top1.ch1c.data[3] ),
    .B(net580));
 sg13g2_nand2_1 _1851_ (.Y(_0620_),
    .A(\top1.ch11c.data[3] ),
    .B(net591));
 sg13g2_a22oi_1 _1852_ (.Y(_0621_),
    .B1(net584),
    .B2(\top1.ch9c.data[3] ),
    .A2(net589),
    .A1(\top1.ch7c.data[3] ));
 sg13g2_a22oi_1 _1853_ (.Y(_0622_),
    .B1(net582),
    .B2(\top1.ch5c.data[3] ),
    .A2(net586),
    .A1(\top1.ch6c.data[3] ));
 sg13g2_nand4_1 _1854_ (.B(_0620_),
    .C(_0621_),
    .A(_0619_),
    .Y(_0623_),
    .D(_0622_));
 sg13g2_a221oi_1 _1855_ (.B2(\top1.ch2c.data[3] ),
    .C1(_0623_),
    .B1(net578),
    .A1(\top1.ch3c.data[3] ),
    .Y(_0624_),
    .A2(net533));
 sg13g2_nand3_1 _1856_ (.B(_0618_),
    .C(_0624_),
    .A(net515),
    .Y(_0625_));
 sg13g2_nor4_2 _1857_ (.A(_0615_),
    .B(_0616_),
    .C(_0617_),
    .Y(_0626_),
    .D(_0625_));
 sg13g2_o21ai_1 _1858_ (.B1(net509),
    .Y(_0627_),
    .A1(\top1.data[0][3] ),
    .A2(net517));
 sg13g2_nand2_1 _1859_ (.Y(_0628_),
    .A(net31),
    .B(net519));
 sg13g2_o21ai_1 _1860_ (.B1(_0628_),
    .Y(_0002_),
    .A1(_0626_),
    .A2(_0627_));
 sg13g2_nand2_1 _1861_ (.Y(_0629_),
    .A(net39),
    .B(net519));
 sg13g2_a22oi_1 _1862_ (.Y(_0630_),
    .B1(net523),
    .B2(\top1.ch13c.data[4] ),
    .A2(net528),
    .A1(\top1.ch15c.data[4] ));
 sg13g2_a22oi_1 _1863_ (.Y(_0631_),
    .B1(net524),
    .B2(\top1.ch12c.data[4] ),
    .A2(net526),
    .A1(\top1.ch14c.data[4] ));
 sg13g2_nand2_1 _1864_ (.Y(_0632_),
    .A(_0630_),
    .B(_0631_));
 sg13g2_and2_1 _1865_ (.A(\top1.ch8c.data[4] ),
    .B(net511),
    .X(_0633_));
 sg13g2_and2_1 _1866_ (.A(\top1.ch4c.data[4] ),
    .B(net514),
    .X(_0634_));
 sg13g2_nand3_1 _1867_ (.B(net531),
    .C(_0581_),
    .A(\top1.ch10c.data[4] ),
    .Y(_0635_));
 sg13g2_nand2_1 _1868_ (.Y(_0636_),
    .A(\top1.ch11c.data[4] ),
    .B(net591));
 sg13g2_nand2_1 _1869_ (.Y(_0637_),
    .A(\top1.ch2c.data[4] ),
    .B(net579));
 sg13g2_a22oi_1 _1870_ (.Y(_0638_),
    .B1(net584),
    .B2(\top1.ch9c.data[4] ),
    .A2(net589),
    .A1(\top1.ch7c.data[4] ));
 sg13g2_a22oi_1 _1871_ (.Y(_0639_),
    .B1(net582),
    .B2(\top1.ch5c.data[4] ),
    .A2(net586),
    .A1(\top1.ch6c.data[4] ));
 sg13g2_nand4_1 _1872_ (.B(_0637_),
    .C(_0638_),
    .A(_0636_),
    .Y(_0640_),
    .D(_0639_));
 sg13g2_a221oi_1 _1873_ (.B2(\top1.ch3c.data[4] ),
    .C1(_0640_),
    .B1(net534),
    .A1(\top1.ch1c.data[4] ),
    .Y(_0641_),
    .A2(net581));
 sg13g2_nand3_1 _1874_ (.B(_0635_),
    .C(_0641_),
    .A(net516),
    .Y(_0642_));
 sg13g2_nor4_2 _1875_ (.A(_0632_),
    .B(_0633_),
    .C(_0634_),
    .Y(_0643_),
    .D(_0642_));
 sg13g2_o21ai_1 _1876_ (.B1(net509),
    .Y(_0644_),
    .A1(\top1.data[0][4] ),
    .A2(net517));
 sg13g2_o21ai_1 _1877_ (.B1(_0629_),
    .Y(_0003_),
    .A1(_0643_),
    .A2(_0644_));
 sg13g2_nand2_1 _1878_ (.Y(_0645_),
    .A(net32),
    .B(net519));
 sg13g2_a22oi_1 _1879_ (.Y(_0646_),
    .B1(net522),
    .B2(\top1.ch13c.data[5] ),
    .A2(net527),
    .A1(\top1.ch14c.data[5] ));
 sg13g2_a22oi_1 _1880_ (.Y(_0647_),
    .B1(net524),
    .B2(\top1.ch12c.data[5] ),
    .A2(net528),
    .A1(\top1.ch15c.data[5] ));
 sg13g2_nand2_1 _1881_ (.Y(_0648_),
    .A(_0646_),
    .B(_0647_));
 sg13g2_and2_1 _1882_ (.A(\top1.ch4c.data[5] ),
    .B(net513),
    .X(_0649_));
 sg13g2_and2_1 _1883_ (.A(\top1.ch8c.data[5] ),
    .B(net511),
    .X(_0650_));
 sg13g2_nand3_1 _1884_ (.B(net530),
    .C(net521),
    .A(\top1.ch10c.data[5] ),
    .Y(_0651_));
 sg13g2_nand2_2 _1885_ (.Y(_0652_),
    .A(\top1.ch1c.data[5] ),
    .B(net580));
 sg13g2_nand2_1 _1886_ (.Y(_0653_),
    .A(\top1.ch2c.data[5] ),
    .B(net578));
 sg13g2_a22oi_1 _1887_ (.Y(_0654_),
    .B1(net584),
    .B2(\top1.ch9c.data[5] ),
    .A2(net589),
    .A1(\top1.ch7c.data[5] ));
 sg13g2_a22oi_1 _1888_ (.Y(_0655_),
    .B1(net582),
    .B2(\top1.ch5c.data[5] ),
    .A2(net586),
    .A1(\top1.ch6c.data[5] ));
 sg13g2_nand4_1 _1889_ (.B(_0653_),
    .C(_0654_),
    .A(_0652_),
    .Y(_0656_),
    .D(_0655_));
 sg13g2_a221oi_1 _1890_ (.B2(\top1.ch3c.data[5] ),
    .C1(_0656_),
    .B1(net533),
    .A1(\top1.ch11c.data[5] ),
    .Y(_0657_),
    .A2(net592));
 sg13g2_nand3_1 _1891_ (.B(_0651_),
    .C(_0657_),
    .A(net515),
    .Y(_0658_));
 sg13g2_nor4_2 _1892_ (.A(_0648_),
    .B(_0649_),
    .C(_0650_),
    .Y(_0659_),
    .D(_0658_));
 sg13g2_o21ai_1 _1893_ (.B1(net509),
    .Y(_0660_),
    .A1(\top1.data[0][5] ),
    .A2(net517));
 sg13g2_o21ai_1 _1894_ (.B1(_0645_),
    .Y(_0004_),
    .A1(_0659_),
    .A2(_0660_));
 sg13g2_a22oi_1 _1895_ (.Y(_0661_),
    .B1(net522),
    .B2(\top1.ch13c.data[6] ),
    .A2(net529),
    .A1(\top1.ch15c.data[6] ));
 sg13g2_a22oi_1 _1896_ (.Y(_0662_),
    .B1(net524),
    .B2(\top1.ch12c.data[6] ),
    .A2(net526),
    .A1(\top1.ch14c.data[6] ));
 sg13g2_nand2_1 _1897_ (.Y(_0663_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_and2_1 _1898_ (.A(\top1.ch8c.data[6] ),
    .B(net511),
    .X(_0664_));
 sg13g2_and2_1 _1899_ (.A(\top1.ch4c.data[6] ),
    .B(net513),
    .X(_0665_));
 sg13g2_nand3_1 _1900_ (.B(net530),
    .C(net521),
    .A(\top1.ch10c.data[6] ),
    .Y(_0666_));
 sg13g2_nand2_2 _1901_ (.Y(_0667_),
    .A(\top1.ch1c.data[6] ),
    .B(net580));
 sg13g2_a22oi_1 _1902_ (.Y(_0668_),
    .B1(net533),
    .B2(\top1.ch3c.data[6] ),
    .A2(net591),
    .A1(\top1.ch11c.data[6] ));
 sg13g2_nand2_1 _1903_ (.Y(_0669_),
    .A(\top1.ch2c.data[6] ),
    .B(net578));
 sg13g2_a22oi_1 _1904_ (.Y(_0670_),
    .B1(net584),
    .B2(\top1.ch9c.data[6] ),
    .A2(net589),
    .A1(\top1.ch7c.data[6] ));
 sg13g2_a22oi_1 _1905_ (.Y(_0671_),
    .B1(net582),
    .B2(\top1.ch5c.data[6] ),
    .A2(net586),
    .A1(\top1.ch6c.data[6] ));
 sg13g2_and4_1 _1906_ (.A(_0667_),
    .B(_0669_),
    .C(_0670_),
    .D(_0671_),
    .X(_0672_));
 sg13g2_nand4_1 _1907_ (.B(_0666_),
    .C(_0668_),
    .A(net515),
    .Y(_0673_),
    .D(_0672_));
 sg13g2_nor4_2 _1908_ (.A(_0663_),
    .B(_0664_),
    .C(_0665_),
    .Y(_0674_),
    .D(_0673_));
 sg13g2_o21ai_1 _1909_ (.B1(net509),
    .Y(_0675_),
    .A1(\top1.data[0][6] ),
    .A2(net517));
 sg13g2_nand2_1 _1910_ (.Y(_0676_),
    .A(net37),
    .B(net519));
 sg13g2_o21ai_1 _1911_ (.B1(_0676_),
    .Y(_0005_),
    .A1(_0674_),
    .A2(_0675_));
 sg13g2_nand2_1 _1912_ (.Y(_0677_),
    .A(net30),
    .B(net519));
 sg13g2_a22oi_1 _1913_ (.Y(_0678_),
    .B1(net526),
    .B2(\top1.ch14c.data[7] ),
    .A2(net528),
    .A1(\top1.ch15c.data[7] ));
 sg13g2_a22oi_1 _1914_ (.Y(_0679_),
    .B1(net522),
    .B2(\top1.ch13c.data[7] ),
    .A2(net525),
    .A1(\top1.ch12c.data[7] ));
 sg13g2_nand2_1 _1915_ (.Y(_0680_),
    .A(_0678_),
    .B(_0679_));
 sg13g2_and2_1 _1916_ (.A(\top1.ch8c.data[7] ),
    .B(net512),
    .X(_0681_));
 sg13g2_and2_1 _1917_ (.A(\top1.ch4c.data[7] ),
    .B(net513),
    .X(_0682_));
 sg13g2_nand3_1 _1918_ (.B(net530),
    .C(net521),
    .A(\top1.ch10c.data[7] ),
    .Y(_0683_));
 sg13g2_nand2_2 _1919_ (.Y(_0684_),
    .A(\top1.ch1c.data[7] ),
    .B(net580));
 sg13g2_nand2_1 _1920_ (.Y(_0685_),
    .A(\top1.ch11c.data[7] ),
    .B(net591));
 sg13g2_a22oi_1 _1921_ (.Y(_0686_),
    .B1(net533),
    .B2(\top1.ch3c.data[7] ),
    .A2(net585),
    .A1(\top1.ch9c.data[7] ));
 sg13g2_a22oi_1 _1922_ (.Y(_0687_),
    .B1(net578),
    .B2(\top1.ch2c.data[7] ),
    .A2(net590),
    .A1(\top1.ch7c.data[7] ));
 sg13g2_a22oi_1 _1923_ (.Y(_0688_),
    .B1(net582),
    .B2(\top1.ch5c.data[7] ),
    .A2(net586),
    .A1(\top1.ch6c.data[7] ));
 sg13g2_and4_1 _1924_ (.A(_0684_),
    .B(_0685_),
    .C(_0687_),
    .D(_0688_),
    .X(_0689_));
 sg13g2_nand4_1 _1925_ (.B(_0683_),
    .C(_0686_),
    .A(net515),
    .Y(_0690_),
    .D(_0689_));
 sg13g2_nor4_2 _1926_ (.A(_0680_),
    .B(_0681_),
    .C(_0682_),
    .Y(_0691_),
    .D(_0690_));
 sg13g2_o21ai_1 _1927_ (.B1(net509),
    .Y(_0692_),
    .A1(\top1.data[0][7] ),
    .A2(net518));
 sg13g2_o21ai_1 _1928_ (.B1(_0677_),
    .Y(_0006_),
    .A1(_0691_),
    .A2(_0692_));
 sg13g2_nand2_1 _1929_ (.Y(_0693_),
    .A(net33),
    .B(net520));
 sg13g2_a22oi_1 _1930_ (.Y(_0694_),
    .B1(net522),
    .B2(\top1.ch13c.data[8] ),
    .A2(net527),
    .A1(\top1.ch14c.data[8] ));
 sg13g2_a22oi_1 _1931_ (.Y(_0695_),
    .B1(net524),
    .B2(\top1.ch12c.data[8] ),
    .A2(net529),
    .A1(\top1.ch15c.data[8] ));
 sg13g2_nand2_1 _1932_ (.Y(_0696_),
    .A(_0694_),
    .B(_0695_));
 sg13g2_and2_1 _1933_ (.A(\top1.ch4c.data[8] ),
    .B(net513),
    .X(_0697_));
 sg13g2_and2_1 _1934_ (.A(\top1.ch8c.data[8] ),
    .B(net512),
    .X(_0698_));
 sg13g2_nand3_1 _1935_ (.B(net531),
    .C(_0581_),
    .A(\top1.ch10c.data[8] ),
    .Y(_0699_));
 sg13g2_nand2_1 _1936_ (.Y(_0700_),
    .A(\top1.ch11c.data[8] ),
    .B(net592));
 sg13g2_nand2_1 _1937_ (.Y(_0701_),
    .A(\top1.ch2c.data[8] ),
    .B(net578));
 sg13g2_a22oi_1 _1938_ (.Y(_0702_),
    .B1(net584),
    .B2(\top1.ch9c.data[8] ),
    .A2(net589),
    .A1(\top1.ch7c.data[8] ));
 sg13g2_a22oi_1 _1939_ (.Y(_0703_),
    .B1(net582),
    .B2(\top1.ch5c.data[8] ),
    .A2(net586),
    .A1(\top1.ch6c.data[8] ));
 sg13g2_nand4_1 _1940_ (.B(_0701_),
    .C(_0702_),
    .A(_0700_),
    .Y(_0704_),
    .D(_0703_));
 sg13g2_a221oi_1 _1941_ (.B2(\top1.ch3c.data[8] ),
    .C1(_0704_),
    .B1(net534),
    .A1(\top1.ch1c.data[8] ),
    .Y(_0705_),
    .A2(net580));
 sg13g2_nand3_1 _1942_ (.B(_0699_),
    .C(_0705_),
    .A(net516),
    .Y(_0706_));
 sg13g2_nor4_2 _1943_ (.A(_0696_),
    .B(_0697_),
    .C(_0698_),
    .Y(_0707_),
    .D(_0706_));
 sg13g2_o21ai_1 _1944_ (.B1(net510),
    .Y(_0708_),
    .A1(\top1.data[0][8] ),
    .A2(net518));
 sg13g2_o21ai_1 _1945_ (.B1(_0693_),
    .Y(_0007_),
    .A1(_0707_),
    .A2(_0708_));
 sg13g2_a22oi_1 _1946_ (.Y(_0709_),
    .B1(net523),
    .B2(\top1.ch13c.data[9] ),
    .A2(net529),
    .A1(\top1.ch15c.data[9] ));
 sg13g2_a22oi_1 _1947_ (.Y(_0710_),
    .B1(net525),
    .B2(\top1.ch12c.data[9] ),
    .A2(net526),
    .A1(\top1.ch14c.data[9] ));
 sg13g2_nand2_1 _1948_ (.Y(_0711_),
    .A(_0709_),
    .B(_0710_));
 sg13g2_and2_1 _1949_ (.A(\top1.ch4c.data[9] ),
    .B(net514),
    .X(_0712_));
 sg13g2_and2_1 _1950_ (.A(\top1.ch8c.data[9] ),
    .B(net511),
    .X(_0713_));
 sg13g2_nand3_1 _1951_ (.B(net531),
    .C(_0581_),
    .A(\top1.ch10c.data[9] ),
    .Y(_0714_));
 sg13g2_nand2_1 _1952_ (.Y(_0715_),
    .A(\top1.ch9c.data[9] ),
    .B(net585));
 sg13g2_nand2_1 _1953_ (.Y(_0716_),
    .A(\top1.ch11c.data[9] ),
    .B(net591));
 sg13g2_a22oi_1 _1954_ (.Y(_0717_),
    .B1(net579),
    .B2(\top1.ch2c.data[9] ),
    .A2(net590),
    .A1(\top1.ch7c.data[9] ));
 sg13g2_a22oi_1 _1955_ (.Y(_0718_),
    .B1(net582),
    .B2(\top1.ch5c.data[9] ),
    .A2(net586),
    .A1(\top1.ch6c.data[9] ));
 sg13g2_nand3_1 _1956_ (.B(_0716_),
    .C(_0718_),
    .A(_0715_),
    .Y(_0719_));
 sg13g2_a221oi_1 _1957_ (.B2(\top1.ch3c.data[9] ),
    .C1(_0719_),
    .B1(net534),
    .A1(\top1.ch1c.data[9] ),
    .Y(_0720_),
    .A2(net580));
 sg13g2_nand4_1 _1958_ (.B(_0714_),
    .C(_0717_),
    .A(net516),
    .Y(_0721_),
    .D(_0720_));
 sg13g2_nor4_2 _1959_ (.A(_0711_),
    .B(_0712_),
    .C(_0713_),
    .Y(_0722_),
    .D(_0721_));
 sg13g2_o21ai_1 _1960_ (.B1(net510),
    .Y(_0723_),
    .A1(\top1.data[0][9] ),
    .A2(net518));
 sg13g2_nand2_1 _1961_ (.Y(_0724_),
    .A(net35),
    .B(net520));
 sg13g2_o21ai_1 _1962_ (.B1(_0724_),
    .Y(_0008_),
    .A1(_0722_),
    .A2(_0723_));
 sg13g2_nand2_1 _1963_ (.Y(_0725_),
    .A(net38),
    .B(net519));
 sg13g2_a22oi_1 _1964_ (.Y(_0726_),
    .B1(net523),
    .B2(\top1.ch13c.data[10] ),
    .A2(net527),
    .A1(\top1.ch14c.data[10] ));
 sg13g2_a22oi_1 _1965_ (.Y(_0727_),
    .B1(net525),
    .B2(\top1.ch12c.data[10] ),
    .A2(net529),
    .A1(\top1.ch15c.data[10] ));
 sg13g2_nand2_1 _1966_ (.Y(_0728_),
    .A(_0726_),
    .B(_0727_));
 sg13g2_and2_1 _1967_ (.A(\top1.ch4c.data[10] ),
    .B(net514),
    .X(_0729_));
 sg13g2_and2_1 _1968_ (.A(\top1.ch8c.data[10] ),
    .B(net512),
    .X(_0730_));
 sg13g2_nand3_1 _1969_ (.B(net530),
    .C(net521),
    .A(\top1.ch10c.data[10] ),
    .Y(_0731_));
 sg13g2_nand2_2 _1970_ (.Y(_0732_),
    .A(\top1.ch1c.data[10] ),
    .B(net580));
 sg13g2_nand2_1 _1971_ (.Y(_0733_),
    .A(\top1.ch2c.data[10] ),
    .B(net578));
 sg13g2_a22oi_1 _1972_ (.Y(_0734_),
    .B1(net584),
    .B2(\top1.ch9c.data[10] ),
    .A2(net589),
    .A1(\top1.ch7c.data[10] ));
 sg13g2_a22oi_1 _1973_ (.Y(_0735_),
    .B1(net583),
    .B2(\top1.ch5c.data[10] ),
    .A2(net587),
    .A1(\top1.ch6c.data[10] ));
 sg13g2_nand4_1 _1974_ (.B(_0733_),
    .C(_0734_),
    .A(_0732_),
    .Y(_0736_),
    .D(_0735_));
 sg13g2_a221oi_1 _1975_ (.B2(\top1.ch3c.data[10] ),
    .C1(_0736_),
    .B1(net533),
    .A1(\top1.ch11c.data[10] ),
    .Y(_0737_),
    .A2(net591));
 sg13g2_nand3_1 _1976_ (.B(_0731_),
    .C(_0737_),
    .A(net515),
    .Y(_0738_));
 sg13g2_nor4_2 _1977_ (.A(_0728_),
    .B(_0729_),
    .C(_0730_),
    .Y(_0739_),
    .D(_0738_));
 sg13g2_o21ai_1 _1978_ (.B1(net510),
    .Y(_0740_),
    .A1(\top1.data[0][10] ),
    .A2(net517));
 sg13g2_o21ai_1 _1979_ (.B1(_0725_),
    .Y(_0009_),
    .A1(_0739_),
    .A2(_0740_));
 sg13g2_a22oi_1 _1980_ (.Y(_0741_),
    .B1(net522),
    .B2(\top1.ch13c.data[0] ),
    .A2(net526),
    .A1(\top1.ch14c.data[0] ));
 sg13g2_a22oi_1 _1981_ (.Y(_0742_),
    .B1(net524),
    .B2(\top1.ch12c.data[0] ),
    .A2(net528),
    .A1(\top1.ch15c.data[0] ));
 sg13g2_nand2_1 _1982_ (.Y(_0743_),
    .A(_0741_),
    .B(_0742_));
 sg13g2_and2_1 _1983_ (.A(\top1.ch8c.data[0] ),
    .B(net511),
    .X(_0744_));
 sg13g2_and2_1 _1984_ (.A(\top1.ch4c.data[0] ),
    .B(net513),
    .X(_0745_));
 sg13g2_nand3_1 _1985_ (.B(net530),
    .C(net521),
    .A(\top1.ch10c.data[0] ),
    .Y(_0746_));
 sg13g2_nand2_2 _1986_ (.Y(_0747_),
    .A(\top1.ch1c.data[0] ),
    .B(net580));
 sg13g2_a22oi_1 _1987_ (.Y(_0748_),
    .B1(net533),
    .B2(\top1.ch3c.data[0] ),
    .A2(net592),
    .A1(\top1.ch11c.data[0] ));
 sg13g2_nand2_1 _1988_ (.Y(_0749_),
    .A(\top1.ch2c.data[0] ),
    .B(net578));
 sg13g2_a22oi_1 _1989_ (.Y(_0750_),
    .B1(net584),
    .B2(\top1.ch9c.data[0] ),
    .A2(net589),
    .A1(\top1.ch7c.data[0] ));
 sg13g2_a22oi_1 _1990_ (.Y(_0751_),
    .B1(net583),
    .B2(\top1.ch5c.data[0] ),
    .A2(net587),
    .A1(\top1.ch6c.data[0] ));
 sg13g2_and4_1 _1991_ (.A(_0747_),
    .B(_0749_),
    .C(_0750_),
    .D(_0751_),
    .X(_0752_));
 sg13g2_nand4_1 _1992_ (.B(_0746_),
    .C(_0748_),
    .A(net515),
    .Y(_0753_),
    .D(_0752_));
 sg13g2_nor4_2 _1993_ (.A(_0743_),
    .B(_0744_),
    .C(_0745_),
    .Y(_0754_),
    .D(_0753_));
 sg13g2_o21ai_1 _1994_ (.B1(net509),
    .Y(_0755_),
    .A1(\top1.data[0][0] ),
    .A2(net517));
 sg13g2_nand2_1 _1995_ (.Y(_0756_),
    .A(net40),
    .B(net519));
 sg13g2_o21ai_1 _1996_ (.B1(_0756_),
    .Y(_0010_),
    .A1(_0754_),
    .A2(_0755_));
 sg13g2_xor2_1 _1997_ (.B(\top1.data[0][0] ),
    .A(\top1.data[0][1] ),
    .X(_0012_));
 sg13g2_and2_1 _1998_ (.A(\top1.data[0][2] ),
    .B(_0514_),
    .X(_0757_));
 sg13g2_o21ai_1 _1999_ (.B1(_0515_),
    .Y(_0758_),
    .A1(\top1.data[0][2] ),
    .A2(_0514_));
 sg13g2_nor2_1 _2000_ (.A(_0757_),
    .B(_0758_),
    .Y(_0013_));
 sg13g2_a21oi_1 _2001_ (.A1(\top1.data[0][3] ),
    .A2(_0515_),
    .Y(_0759_),
    .B1(_0757_));
 sg13g2_a21oi_1 _2002_ (.A1(\top1.data[0][3] ),
    .A2(_0757_),
    .Y(_0014_),
    .B1(_0759_));
 sg13g2_nand3_1 _2003_ (.B(\top1.data[0][4] ),
    .C(_0757_),
    .A(\top1.data[0][3] ),
    .Y(_0760_));
 sg13g2_a21oi_1 _2004_ (.A1(\top1.data[0][3] ),
    .A2(_0757_),
    .Y(_0761_),
    .B1(\top1.data[0][4] ));
 sg13g2_nor2_1 _2005_ (.A(_0516_),
    .B(_0761_),
    .Y(_0762_));
 sg13g2_and2_1 _2006_ (.A(_0760_),
    .B(_0762_),
    .X(_0015_));
 sg13g2_nand2b_1 _2007_ (.Y(_0763_),
    .B(_0760_),
    .A_N(\top1.data[0][5] ));
 sg13g2_and2_1 _2008_ (.A(_0515_),
    .B(_0763_),
    .X(_0016_));
 sg13g2_a21oi_2 _2009_ (.B1(_0565_),
    .Y(_0764_),
    .A2(_0522_),
    .A1(net46));
 sg13g2_nand3_1 _2010_ (.B(net55),
    .C(net51),
    .A(net41),
    .Y(_0765_));
 sg13g2_nor2_2 _2011_ (.A(net49),
    .B(_0765_),
    .Y(_0766_));
 sg13g2_nor2_1 _2012_ (.A(net46),
    .B(_0523_),
    .Y(_0767_));
 sg13g2_o21ai_1 _2013_ (.B1(_0766_),
    .Y(_0768_),
    .A1(_0561_),
    .A2(_0767_));
 sg13g2_o21ai_1 _2014_ (.B1(net52),
    .Y(_0769_),
    .A1(\top1.FSM1.counter_register[2] ),
    .A2(_0765_));
 sg13g2_o21ai_1 _2015_ (.B1(_0769_),
    .Y(_0770_),
    .A1(net597),
    .A2(_0523_));
 sg13g2_nand2_1 _2016_ (.Y(_0771_),
    .A(net46),
    .B(_0770_));
 sg13g2_a21oi_1 _2017_ (.A1(_0768_),
    .A2(net47),
    .Y(\top1.FSM1.state_next[0] ),
    .B1(_0764_));
 sg13g2_nor2_1 _2018_ (.A(_0543_),
    .B(_0766_),
    .Y(_0772_));
 sg13g2_a21oi_1 _2019_ (.A1(_0532_),
    .A2(net53),
    .Y(_0773_),
    .B1(_0772_));
 sg13g2_nor2_1 _2020_ (.A(_0764_),
    .B(_0773_),
    .Y(\top1.FSM1.state_next[1] ));
 sg13g2_nor2_1 _2021_ (.A(_0532_),
    .B(_0772_),
    .Y(_0774_));
 sg13g2_nor2_1 _2022_ (.A(_0525_),
    .B(_0543_),
    .Y(_0775_));
 sg13g2_nor2_1 _2023_ (.A(_0525_),
    .B(_0774_),
    .Y(_0776_));
 sg13g2_mux2_1 _2024_ (.A0(net588),
    .A1(_0544_),
    .S(_0766_),
    .X(_0777_));
 sg13g2_nor3_1 _2025_ (.A(_0538_),
    .B(_0776_),
    .C(_0777_),
    .Y(_0778_));
 sg13g2_a21oi_1 _2026_ (.A1(_0550_),
    .A2(_0778_),
    .Y(\top1.FSM1.state_next[2] ),
    .B1(_0764_));
 sg13g2_and2_1 _2027_ (.A(net588),
    .B(_0766_),
    .X(_0779_));
 sg13g2_nor4_2 _2028_ (.A(_0547_),
    .B(net590),
    .C(_0776_),
    .Y(_0780_),
    .D(_0779_));
 sg13g2_nor2_1 _2029_ (.A(_0764_),
    .B(_0780_),
    .Y(\top1.FSM1.state_next[3] ));
 sg13g2_a21oi_1 _2030_ (.A1(_0766_),
    .A2(_0775_),
    .Y(_0781_),
    .B1(_0767_));
 sg13g2_nor2_1 _2031_ (.A(_0764_),
    .B(_0781_),
    .Y(\top1.FSM1.state_next[4] ));
 sg13g2_nor4_1 _2032_ (.A(_0836_),
    .B(net605),
    .C(net600),
    .D(_0521_),
    .Y(_0782_));
 sg13g2_nor2b_1 _2033_ (.A(net576),
    .B_N(net667),
    .Y(_0033_));
 sg13g2_nand2_1 _2034_ (.Y(_0783_),
    .A(\top1.ch5c.data[11] ),
    .B(net583));
 sg13g2_a22oi_1 _2035_ (.Y(_0784_),
    .B1(_0582_),
    .B2(\top1.ch10c.data[11] ),
    .A2(net588),
    .A1(\top1.ch6c.data[11] ));
 sg13g2_and2_1 _2036_ (.A(net515),
    .B(_0783_),
    .X(_0785_));
 sg13g2_a22oi_1 _2037_ (.Y(_0786_),
    .B1(net579),
    .B2(\top1.ch2c.data[11] ),
    .A2(net514),
    .A1(\top1.ch4c.data[11] ));
 sg13g2_a22oi_1 _2038_ (.Y(_0787_),
    .B1(net533),
    .B2(\top1.ch3c.data[11] ),
    .A2(_0573_),
    .A1(\top1.ch12c.data[11] ));
 sg13g2_and4_1 _2039_ (.A(_0784_),
    .B(_0785_),
    .C(_0786_),
    .D(_0787_),
    .X(_0788_));
 sg13g2_a22oi_1 _2040_ (.Y(_0789_),
    .B1(net585),
    .B2(\top1.ch9c.data[11] ),
    .A2(net527),
    .A1(\top1.ch14c.data[11] ));
 sg13g2_a22oi_1 _2041_ (.Y(_0790_),
    .B1(net581),
    .B2(\top1.ch1c.data[11] ),
    .A2(net593),
    .A1(\top1.ch11c.data[11] ));
 sg13g2_a22oi_1 _2042_ (.Y(_0791_),
    .B1(net512),
    .B2(\top1.ch8c.data[11] ),
    .A2(net589),
    .A1(\top1.ch7c.data[11] ));
 sg13g2_a22oi_1 _2043_ (.Y(_0792_),
    .B1(net522),
    .B2(\top1.ch13c.data[11] ),
    .A2(net528),
    .A1(\top1.ch15c.data[11] ));
 sg13g2_and4_1 _2044_ (.A(_0789_),
    .B(_0790_),
    .C(_0791_),
    .D(_0792_),
    .X(_0793_));
 sg13g2_o21ai_1 _2045_ (.B1(net510),
    .Y(_0794_),
    .A1(\top1.data[0][11] ),
    .A2(net518));
 sg13g2_a21oi_2 _2046_ (.B1(_0794_),
    .Y(_0290_),
    .A2(_0793_),
    .A1(_0788_));
 sg13g2_xor2_1 _2047_ (.B(_0516_),
    .A(\top1.data[0][6] ),
    .X(_0399_));
 sg13g2_a21oi_1 _2048_ (.A1(\top1.data[0][6] ),
    .A2(_0516_),
    .Y(_0795_),
    .B1(\top1.data[0][7] ));
 sg13g2_nor2_1 _2049_ (.A(_0517_),
    .B(_0795_),
    .Y(_0400_));
 sg13g2_nor2_1 _2050_ (.A(\top1.data[0][8] ),
    .B(_0517_),
    .Y(_0796_));
 sg13g2_and2_1 _2051_ (.A(\top1.data[0][8] ),
    .B(_0517_),
    .X(_0797_));
 sg13g2_nor3_1 _2052_ (.A(_0518_),
    .B(_0796_),
    .C(_0797_),
    .Y(_0401_));
 sg13g2_xnor2_1 _2053_ (.Y(_0798_),
    .A(\top1.data[0][9] ),
    .B(_0797_));
 sg13g2_nor2_1 _2054_ (.A(_0519_),
    .B(_0798_),
    .Y(_0402_));
 sg13g2_a21oi_1 _2055_ (.A1(\top1.data[0][9] ),
    .A2(_0797_),
    .Y(_0799_),
    .B1(\top1.data[0][10] ));
 sg13g2_nand3_1 _2056_ (.B(\top1.data[0][10] ),
    .C(_0797_),
    .A(\top1.data[0][9] ),
    .Y(_0800_));
 sg13g2_nand2b_1 _2057_ (.Y(_0801_),
    .B(_0800_),
    .A_N(_0799_));
 sg13g2_nor2_1 _2058_ (.A(_0519_),
    .B(_0801_),
    .Y(_0403_));
 sg13g2_a21oi_1 _2059_ (.A1(_0839_),
    .A2(_0800_),
    .Y(_0404_),
    .B1(_0518_));
 sg13g2_or2_1 _2060_ (.X(_0802_),
    .B(_0766_),
    .A(_0565_));
 sg13g2_xor2_1 _2061_ (.B(_0802_),
    .A(net45),
    .X(_0417_));
 sg13g2_and3_1 _2062_ (.X(_0803_),
    .A(net41),
    .B(net54),
    .C(_0802_));
 sg13g2_a21oi_1 _2063_ (.A1(\top1.FSM1.counter_register[0] ),
    .A2(_0565_),
    .Y(_0804_),
    .B1(net41));
 sg13g2_nor2_1 _2064_ (.A(_0803_),
    .B(net42),
    .Y(_0418_));
 sg13g2_a21oi_1 _2065_ (.A1(_0840_),
    .A2(_0803_),
    .Y(_0805_),
    .B1(net49));
 sg13g2_a21oi_1 _2066_ (.A1(net49),
    .A2(_0803_),
    .Y(_0419_),
    .B1(_0805_));
 sg13g2_a21oi_1 _2067_ (.A1(\top1.FSM1.counter_register[2] ),
    .A2(_0803_),
    .Y(_0806_),
    .B1(net43));
 sg13g2_a21oi_1 _2068_ (.A1(net43),
    .A2(_0803_),
    .Y(_0420_),
    .B1(_0806_));
 sg13g2_nor2b_1 _2069_ (.A(net545),
    .B_N(net643),
    .Y(_0034_));
 sg13g2_nor2b_1 _2070_ (.A(net545),
    .B_N(net643),
    .Y(_0035_));
 sg13g2_nor2b_1 _2071_ (.A(net545),
    .B_N(net643),
    .Y(_0036_));
 sg13g2_nor2b_1 _2072_ (.A(net545),
    .B_N(net643),
    .Y(_0037_));
 sg13g2_nor2b_1 _2073_ (.A(net546),
    .B_N(net644),
    .Y(_0038_));
 sg13g2_nor2b_1 _2074_ (.A(net561),
    .B_N(net659),
    .Y(_0039_));
 sg13g2_nor2b_1 _2075_ (.A(net545),
    .B_N(net643),
    .Y(_0040_));
 sg13g2_nor2b_1 _2076_ (.A(net561),
    .B_N(net659),
    .Y(_0041_));
 sg13g2_nor2b_1 _2077_ (.A(net563),
    .B_N(net661),
    .Y(_0042_));
 sg13g2_nor2b_1 _2078_ (.A(net563),
    .B_N(net661),
    .Y(_0043_));
 sg13g2_nor2b_1 _2079_ (.A(net561),
    .B_N(net659),
    .Y(_0044_));
 sg13g2_nor2b_1 _2080_ (.A(net563),
    .B_N(net661),
    .Y(_0045_));
 sg13g2_nor2b_1 _2081_ (.A(net562),
    .B_N(net660),
    .Y(_0046_));
 sg13g2_nor2b_1 _2082_ (.A(net562),
    .B_N(net660),
    .Y(_0047_));
 sg13g2_nor2b_1 _2083_ (.A(net561),
    .B_N(net659),
    .Y(_0048_));
 sg13g2_nor2b_1 _2084_ (.A(net562),
    .B_N(net660),
    .Y(_0049_));
 sg13g2_nor2b_1 _2085_ (.A(net566),
    .B_N(net664),
    .Y(_0050_));
 sg13g2_nor2b_1 _2086_ (.A(net566),
    .B_N(net664),
    .Y(_0051_));
 sg13g2_nor2b_1 _2087_ (.A(net566),
    .B_N(net664),
    .Y(_0052_));
 sg13g2_nor2b_1 _2088_ (.A(net567),
    .B_N(net666),
    .Y(_0053_));
 sg13g2_nor2b_1 _2089_ (.A(net566),
    .B_N(net664),
    .Y(_0054_));
 sg13g2_nor2b_1 _2090_ (.A(net567),
    .B_N(net665),
    .Y(_0055_));
 sg13g2_nor2b_1 _2091_ (.A(net567),
    .B_N(net665),
    .Y(_0056_));
 sg13g2_nor2b_1 _2092_ (.A(net567),
    .B_N(net665),
    .Y(_0057_));
 sg13g2_nor2b_1 _2093_ (.A(net544),
    .B_N(net642),
    .Y(_0058_));
 sg13g2_nor2b_1 _2094_ (.A(net544),
    .B_N(net642),
    .Y(_0059_));
 sg13g2_nor2b_1 _2095_ (.A(net544),
    .B_N(net642),
    .Y(_0060_));
 sg13g2_nor2b_1 _2096_ (.A(net544),
    .B_N(net642),
    .Y(_0061_));
 sg13g2_nor2b_1 _2097_ (.A(net549),
    .B_N(net647),
    .Y(_0062_));
 sg13g2_nor2b_1 _2098_ (.A(net549),
    .B_N(net647),
    .Y(_0063_));
 sg13g2_nor2b_1 _2099_ (.A(net546),
    .B_N(net642),
    .Y(_0064_));
 sg13g2_nor2b_1 _2100_ (.A(net544),
    .B_N(net644),
    .Y(_0065_));
 sg13g2_nor2b_1 _2101_ (.A(net544),
    .B_N(net642),
    .Y(_0066_));
 sg13g2_nor2b_1 _2102_ (.A(net544),
    .B_N(net642),
    .Y(_0067_));
 sg13g2_nor2b_1 _2103_ (.A(net544),
    .B_N(net642),
    .Y(_0068_));
 sg13g2_nor2b_1 _2104_ (.A(net547),
    .B_N(net645),
    .Y(_0069_));
 sg13g2_nor2b_1 _2105_ (.A(net557),
    .B_N(net655),
    .Y(_0070_));
 sg13g2_nor2b_1 _2106_ (.A(net557),
    .B_N(net655),
    .Y(_0071_));
 sg13g2_nor2b_1 _2107_ (.A(net556),
    .B_N(net654),
    .Y(_0072_));
 sg13g2_nor2b_1 _2108_ (.A(net557),
    .B_N(net655),
    .Y(_0073_));
 sg13g2_nor2b_1 _2109_ (.A(net557),
    .B_N(net655),
    .Y(_0074_));
 sg13g2_nor2b_1 _2110_ (.A(net556),
    .B_N(net654),
    .Y(_0075_));
 sg13g2_nor2b_1 _2111_ (.A(net556),
    .B_N(net654),
    .Y(_0076_));
 sg13g2_nor2b_1 _2112_ (.A(net568),
    .B_N(net668),
    .Y(_0077_));
 sg13g2_nor2b_1 _2113_ (.A(net568),
    .B_N(net668),
    .Y(_0078_));
 sg13g2_nor2b_1 _2114_ (.A(net568),
    .B_N(net668),
    .Y(_0079_));
 sg13g2_nor2b_1 _2115_ (.A(net568),
    .B_N(net668),
    .Y(_0080_));
 sg13g2_nor2b_1 _2116_ (.A(net568),
    .B_N(net668),
    .Y(_0081_));
 sg13g2_nor2b_1 _2117_ (.A(net547),
    .B_N(net645),
    .Y(_0082_));
 sg13g2_nor2b_1 _2118_ (.A(net547),
    .B_N(net645),
    .Y(_0083_));
 sg13g2_nor2b_1 _2119_ (.A(net547),
    .B_N(net645),
    .Y(_0084_));
 sg13g2_nor2b_1 _2120_ (.A(net547),
    .B_N(net645),
    .Y(_0085_));
 sg13g2_nor2b_1 _2121_ (.A(net547),
    .B_N(net645),
    .Y(_0086_));
 sg13g2_nor2b_1 _2122_ (.A(net547),
    .B_N(net645),
    .Y(_0087_));
 sg13g2_nor2b_1 _2123_ (.A(net568),
    .B_N(net668),
    .Y(_0088_));
 sg13g2_nor2b_1 _2124_ (.A(net568),
    .B_N(net668),
    .Y(_0089_));
 sg13g2_nor2b_1 _2125_ (.A(net557),
    .B_N(net655),
    .Y(_0090_));
 sg13g2_nor2b_1 _2126_ (.A(net556),
    .B_N(net654),
    .Y(_0091_));
 sg13g2_nor2b_1 _2127_ (.A(net556),
    .B_N(net654),
    .Y(_0092_));
 sg13g2_nor2b_1 _2128_ (.A(net556),
    .B_N(net654),
    .Y(_0093_));
 sg13g2_nor2b_1 _2129_ (.A(net542),
    .B_N(net640),
    .Y(_0094_));
 sg13g2_nor2b_1 _2130_ (.A(net542),
    .B_N(net640),
    .Y(_0095_));
 sg13g2_nor2b_1 _2131_ (.A(net542),
    .B_N(net640),
    .Y(_0096_));
 sg13g2_nor2b_1 _2132_ (.A(net542),
    .B_N(net640),
    .Y(_0097_));
 sg13g2_nor2b_1 _2133_ (.A(net542),
    .B_N(net640),
    .Y(_0098_));
 sg13g2_nor2b_1 _2134_ (.A(net542),
    .B_N(net640),
    .Y(_0099_));
 sg13g2_nor2b_1 _2135_ (.A(net543),
    .B_N(net641),
    .Y(_0100_));
 sg13g2_nor2b_1 _2136_ (.A(net543),
    .B_N(net641),
    .Y(_0101_));
 sg13g2_nor2b_1 _2137_ (.A(net543),
    .B_N(net641),
    .Y(_0102_));
 sg13g2_nor2b_1 _2138_ (.A(net542),
    .B_N(net640),
    .Y(_0103_));
 sg13g2_nor2b_1 _2139_ (.A(net542),
    .B_N(net640),
    .Y(_0104_));
 sg13g2_nor2b_1 _2140_ (.A(net555),
    .B_N(net653),
    .Y(_0105_));
 sg13g2_nor2b_1 _2141_ (.A(net553),
    .B_N(net651),
    .Y(_0106_));
 sg13g2_nor2b_1 _2142_ (.A(net553),
    .B_N(net651),
    .Y(_0107_));
 sg13g2_nor2b_1 _2143_ (.A(net553),
    .B_N(net651),
    .Y(_0108_));
 sg13g2_nor2b_1 _2144_ (.A(net553),
    .B_N(net651),
    .Y(_0109_));
 sg13g2_nor2b_1 _2145_ (.A(net553),
    .B_N(net651),
    .Y(_0110_));
 sg13g2_nor2b_1 _2146_ (.A(net553),
    .B_N(net651),
    .Y(_0111_));
 sg13g2_nor2b_1 _2147_ (.A(net553),
    .B_N(net651),
    .Y(_0112_));
 sg13g2_nor2b_1 _2148_ (.A(net553),
    .B_N(net651),
    .Y(_0113_));
 sg13g2_nor2b_1 _2149_ (.A(net552),
    .B_N(net650),
    .Y(_0114_));
 sg13g2_nor2b_1 _2150_ (.A(net552),
    .B_N(net650),
    .Y(_0115_));
 sg13g2_nor2b_1 _2151_ (.A(net552),
    .B_N(net650),
    .Y(_0116_));
 sg13g2_nor2b_1 _2152_ (.A(net552),
    .B_N(net650),
    .Y(_0117_));
 sg13g2_nor2b_1 _2153_ (.A(net554),
    .B_N(net652),
    .Y(_0118_));
 sg13g2_nor2b_1 _2154_ (.A(net554),
    .B_N(net652),
    .Y(_0119_));
 sg13g2_nor2b_1 _2155_ (.A(net554),
    .B_N(net652),
    .Y(_0120_));
 sg13g2_nor2b_1 _2156_ (.A(net558),
    .B_N(net656),
    .Y(_0121_));
 sg13g2_nor2b_1 _2157_ (.A(net554),
    .B_N(net652),
    .Y(_0122_));
 sg13g2_nor2b_1 _2158_ (.A(net554),
    .B_N(net652),
    .Y(_0123_));
 sg13g2_nor2b_1 _2159_ (.A(net558),
    .B_N(net656),
    .Y(_0124_));
 sg13g2_nor2b_1 _2160_ (.A(net558),
    .B_N(net656),
    .Y(_0125_));
 sg13g2_nor2b_1 _2161_ (.A(net558),
    .B_N(net656),
    .Y(_0126_));
 sg13g2_nor2b_1 _2162_ (.A(net559),
    .B_N(net657),
    .Y(_0127_));
 sg13g2_nor2b_1 _2163_ (.A(net559),
    .B_N(net657),
    .Y(_0128_));
 sg13g2_nor2b_1 _2164_ (.A(net558),
    .B_N(net656),
    .Y(_0129_));
 sg13g2_nor2b_1 _2165_ (.A(net570),
    .B_N(net670),
    .Y(_0130_));
 sg13g2_nor2b_1 _2166_ (.A(net570),
    .B_N(net670),
    .Y(_0131_));
 sg13g2_nor2b_1 _2167_ (.A(net570),
    .B_N(net670),
    .Y(_0132_));
 sg13g2_nor2b_1 _2168_ (.A(net559),
    .B_N(net657),
    .Y(_0133_));
 sg13g2_nor2b_1 _2169_ (.A(net559),
    .B_N(net657),
    .Y(_0134_));
 sg13g2_nor2b_1 _2170_ (.A(net559),
    .B_N(net657),
    .Y(_0135_));
 sg13g2_nor2b_1 _2171_ (.A(net559),
    .B_N(net657),
    .Y(_0136_));
 sg13g2_nor2b_1 _2172_ (.A(net558),
    .B_N(net657),
    .Y(_0137_));
 sg13g2_nor2b_1 _2173_ (.A(net559),
    .B_N(net656),
    .Y(_0138_));
 sg13g2_nor2b_1 _2174_ (.A(net570),
    .B_N(net670),
    .Y(_0139_));
 sg13g2_nor2b_1 _2175_ (.A(net570),
    .B_N(net670),
    .Y(_0140_));
 sg13g2_nor2b_1 _2176_ (.A(net570),
    .B_N(net670),
    .Y(_0141_));
 sg13g2_nor2b_1 _2177_ (.A(net548),
    .B_N(net646),
    .Y(_0142_));
 sg13g2_nor2b_1 _2178_ (.A(net548),
    .B_N(net646),
    .Y(_0143_));
 sg13g2_nor2b_1 _2179_ (.A(net548),
    .B_N(net646),
    .Y(_0144_));
 sg13g2_nor2b_1 _2180_ (.A(net548),
    .B_N(net646),
    .Y(_0145_));
 sg13g2_nor2b_1 _2181_ (.A(net563),
    .B_N(net661),
    .Y(_0146_));
 sg13g2_nor2b_1 _2182_ (.A(net563),
    .B_N(net661),
    .Y(_0147_));
 sg13g2_nor2b_1 _2183_ (.A(net563),
    .B_N(net661),
    .Y(_0148_));
 sg13g2_nor2b_1 _2184_ (.A(net563),
    .B_N(net661),
    .Y(_0149_));
 sg13g2_nor2b_1 _2185_ (.A(net564),
    .B_N(net662),
    .Y(_0150_));
 sg13g2_nor2b_1 _2186_ (.A(net564),
    .B_N(net662),
    .Y(_0151_));
 sg13g2_nor2b_1 _2187_ (.A(net563),
    .B_N(net661),
    .Y(_0152_));
 sg13g2_nor2b_1 _2188_ (.A(net564),
    .B_N(net662),
    .Y(_0153_));
 sg13g2_nor2b_1 _2189_ (.A(net571),
    .B_N(net671),
    .Y(_0154_));
 sg13g2_nor2b_1 _2190_ (.A(net568),
    .B_N(net668),
    .Y(_0155_));
 sg13g2_nor2b_1 _2191_ (.A(net569),
    .B_N(net669),
    .Y(_0156_));
 sg13g2_nor2b_1 _2192_ (.A(net569),
    .B_N(net669),
    .Y(_0157_));
 sg13g2_nor2b_1 _2193_ (.A(net574),
    .B_N(net676),
    .Y(_0158_));
 sg13g2_nor2b_1 _2194_ (.A(net574),
    .B_N(net676),
    .Y(_0159_));
 sg13g2_nor2b_1 _2195_ (.A(net575),
    .B_N(net673),
    .Y(_0160_));
 sg13g2_nor2b_1 _2196_ (.A(net575),
    .B_N(net672),
    .Y(_0161_));
 sg13g2_nor2b_1 _2197_ (.A(net575),
    .B_N(net673),
    .Y(_0162_));
 sg13g2_nor2b_1 _2198_ (.A(net575),
    .B_N(net677),
    .Y(_0163_));
 sg13g2_nor2b_1 _2199_ (.A(net575),
    .B_N(net673),
    .Y(_0164_));
 sg13g2_nor2b_1 _2200_ (.A(net575),
    .B_N(net672),
    .Y(_0165_));
 sg13g2_nor2b_1 _2201_ (.A(net569),
    .B_N(net669),
    .Y(_0166_));
 sg13g2_nor2b_1 _2202_ (.A(net571),
    .B_N(net671),
    .Y(_0167_));
 sg13g2_nor2b_1 _2203_ (.A(net569),
    .B_N(net669),
    .Y(_0168_));
 sg13g2_nor2b_1 _2204_ (.A(net569),
    .B_N(net669),
    .Y(_0169_));
 sg13g2_nor2b_1 _2205_ (.A(net570),
    .B_N(net670),
    .Y(_0170_));
 sg13g2_nor2b_1 _2206_ (.A(net571),
    .B_N(net671),
    .Y(_0171_));
 sg13g2_nor2b_1 _2207_ (.A(net569),
    .B_N(net669),
    .Y(_0172_));
 sg13g2_nor2b_1 _2208_ (.A(net569),
    .B_N(net669),
    .Y(_0173_));
 sg13g2_nor2b_1 _2209_ (.A(net574),
    .B_N(net676),
    .Y(_0174_));
 sg13g2_nor2b_1 _2210_ (.A(net574),
    .B_N(net676),
    .Y(_0175_));
 sg13g2_nor2b_1 _2211_ (.A(net574),
    .B_N(net676),
    .Y(_0176_));
 sg13g2_nor2b_1 _2212_ (.A(net569),
    .B_N(net669),
    .Y(_0177_));
 sg13g2_nor2b_1 _2213_ (.A(net572),
    .B_N(net674),
    .Y(_0178_));
 sg13g2_nor2b_1 _2214_ (.A(net572),
    .B_N(net674),
    .Y(_0179_));
 sg13g2_nor2b_1 _2215_ (.A(net572),
    .B_N(net674),
    .Y(_0180_));
 sg13g2_nor2b_1 _2216_ (.A(net572),
    .B_N(net674),
    .Y(_0181_));
 sg13g2_nor2b_1 _2217_ (.A(net572),
    .B_N(net674),
    .Y(_0182_));
 sg13g2_nor2b_1 _2218_ (.A(net572),
    .B_N(net674),
    .Y(_0183_));
 sg13g2_nor2b_1 _2219_ (.A(net572),
    .B_N(net674),
    .Y(_0184_));
 sg13g2_nor2b_1 _2220_ (.A(net572),
    .B_N(net675),
    .Y(_0185_));
 sg13g2_nor2b_1 _2221_ (.A(net573),
    .B_N(net674),
    .Y(_0186_));
 sg13g2_nor2b_1 _2222_ (.A(net573),
    .B_N(net675),
    .Y(_0187_));
 sg13g2_nor2b_1 _2223_ (.A(net573),
    .B_N(net675),
    .Y(_0188_));
 sg13g2_nor2b_1 _2224_ (.A(net573),
    .B_N(net675),
    .Y(_0189_));
 sg13g2_nor2b_1 _2225_ (.A(net545),
    .B_N(net643),
    .Y(_0190_));
 sg13g2_nor2b_1 _2226_ (.A(net545),
    .B_N(net643),
    .Y(_0191_));
 sg13g2_nor2b_1 _2227_ (.A(net545),
    .B_N(net643),
    .Y(_0192_));
 sg13g2_nor2b_1 _2228_ (.A(net561),
    .B_N(net659),
    .Y(_0193_));
 sg13g2_nor2b_1 _2229_ (.A(net562),
    .B_N(net660),
    .Y(_0194_));
 sg13g2_nor2b_1 _2230_ (.A(net561),
    .B_N(net659),
    .Y(_0195_));
 sg13g2_nor2b_1 _2231_ (.A(net561),
    .B_N(net659),
    .Y(_0196_));
 sg13g2_nor2b_1 _2232_ (.A(net562),
    .B_N(net660),
    .Y(_0197_));
 sg13g2_nor2b_1 _2233_ (.A(net562),
    .B_N(net660),
    .Y(_0198_));
 sg13g2_nor2b_1 _2234_ (.A(net566),
    .B_N(net664),
    .Y(_0199_));
 sg13g2_nor2b_1 _2235_ (.A(net566),
    .B_N(net664),
    .Y(_0200_));
 sg13g2_nor2b_1 _2236_ (.A(net566),
    .B_N(net664),
    .Y(_0201_));
 sg13g2_nor2b_1 _2237_ (.A(net550),
    .B_N(net648),
    .Y(_0202_));
 sg13g2_nor2b_1 _2238_ (.A(net550),
    .B_N(net648),
    .Y(_0203_));
 sg13g2_nor2b_1 _2239_ (.A(net551),
    .B_N(net649),
    .Y(_0204_));
 sg13g2_nor2b_1 _2240_ (.A(net551),
    .B_N(net649),
    .Y(_0205_));
 sg13g2_nor2b_1 _2241_ (.A(net551),
    .B_N(net649),
    .Y(_0206_));
 sg13g2_nor2b_1 _2242_ (.A(net551),
    .B_N(net649),
    .Y(_0207_));
 sg13g2_nor2b_1 _2243_ (.A(net550),
    .B_N(net648),
    .Y(_0208_));
 sg13g2_nor2b_1 _2244_ (.A(net550),
    .B_N(net648),
    .Y(_0209_));
 sg13g2_nor2b_1 _2245_ (.A(net550),
    .B_N(net648),
    .Y(_0210_));
 sg13g2_nor2b_1 _2246_ (.A(net550),
    .B_N(net648),
    .Y(_0211_));
 sg13g2_nor2b_1 _2247_ (.A(net550),
    .B_N(net648),
    .Y(_0212_));
 sg13g2_nor2b_1 _2248_ (.A(net550),
    .B_N(net648),
    .Y(_0213_));
 sg13g2_nor2b_1 _2249_ (.A(net561),
    .B_N(net659),
    .Y(_0214_));
 sg13g2_nor2b_1 _2250_ (.A(net564),
    .B_N(net662),
    .Y(_0215_));
 sg13g2_nor2b_1 _2251_ (.A(net566),
    .B_N(net664),
    .Y(_0216_));
 sg13g2_nor2b_1 _2252_ (.A(net547),
    .B_N(net645),
    .Y(_0217_));
 sg13g2_nor2b_1 _2253_ (.A(net556),
    .B_N(net654),
    .Y(_0218_));
 sg13g2_nor2b_1 _2254_ (.A(net556),
    .B_N(net654),
    .Y(_0219_));
 sg13g2_nor2b_1 _2255_ (.A(net552),
    .B_N(net650),
    .Y(_0220_));
 sg13g2_nor2b_1 _2256_ (.A(net552),
    .B_N(net650),
    .Y(_0221_));
 sg13g2_nor2b_1 _2257_ (.A(net554),
    .B_N(net652),
    .Y(_0222_));
 sg13g2_nor2b_1 _2258_ (.A(net558),
    .B_N(net656),
    .Y(_0223_));
 sg13g2_nor2b_1 _2259_ (.A(net558),
    .B_N(net656),
    .Y(_0224_));
 sg13g2_nor2b_2 _2260_ (.A(net575),
    .B_N(net672),
    .Y(_0225_));
 sg13g2_nor2b_1 _2261_ (.A(net573),
    .B_N(net675),
    .Y(_0226_));
 sg13g2_nor2b_1 _2262_ (.A(net573),
    .B_N(net675),
    .Y(_0227_));
 sg13g2_nor2b_1 _2263_ (.A(net573),
    .B_N(net675),
    .Y(_0228_));
 sg13g2_dfrbp_1 _2264_ (.CLK(net639),
    .RESET_B(_0033_),
    .D(_0229_),
    .Q_N(_1213_),
    .Q(\top1.ovf_RTC ));
 sg13g2_dfrbp_1 _2265_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net18),
    .D(_0000_),
    .Q_N(_1214_),
    .Q(\top1.PISO_register1.register[0] ));
 sg13g2_dfrbp_1 _2266_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net19),
    .D(_0001_),
    .Q_N(_1215_),
    .Q(\top1.PISO_register1.register[1] ));
 sg13g2_dfrbp_1 _2267_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net20),
    .D(_0002_),
    .Q_N(_1216_),
    .Q(\top1.PISO_register1.register[2] ));
 sg13g2_dfrbp_1 _2268_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net21),
    .D(_0003_),
    .Q_N(_1217_),
    .Q(\top1.PISO_register1.register[3] ));
 sg13g2_dfrbp_1 _2269_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net22),
    .D(_0004_),
    .Q_N(_1218_),
    .Q(\top1.PISO_register1.register[4] ));
 sg13g2_dfrbp_1 _2270_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net23),
    .D(_0005_),
    .Q_N(_1219_),
    .Q(\top1.PISO_register1.register[5] ));
 sg13g2_dfrbp_1 _2271_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net24),
    .D(_0006_),
    .Q_N(_1220_),
    .Q(\top1.PISO_register1.register[6] ));
 sg13g2_dfrbp_1 _2272_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net25),
    .D(_0007_),
    .Q_N(_1221_),
    .Q(\top1.PISO_register1.register[7] ));
 sg13g2_dfrbp_1 _2273_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net26),
    .D(_0008_),
    .Q_N(_1222_),
    .Q(\top1.PISO_register1.register[8] ));
 sg13g2_dfrbp_1 _2274_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net27),
    .D(_0009_),
    .Q_N(_1223_),
    .Q(\top1.PISO_register1.register[9] ));
 sg13g2_dfrbp_1 _2275_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net28),
    .D(_0010_),
    .Q_N(_1224_),
    .Q(\top1.PISO_register1.serial_out ));
 sg13g2_dfrbp_1 _2276_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net672),
    .D(net48),
    .Q_N(_1225_),
    .Q(\top1.FSM1.state_reg[0] ));
 sg13g2_dfrbp_1 _2277_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net673),
    .D(\top1.FSM1.state_next[1] ),
    .Q_N(_1226_),
    .Q(\top1.FSM1.state_reg[1] ));
 sg13g2_dfrbp_1 _2278_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net673),
    .D(\top1.FSM1.state_next[2] ),
    .Q_N(_1227_),
    .Q(\top1.FSM1.state_reg[2] ));
 sg13g2_dfrbp_1 _2279_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net673),
    .D(\top1.FSM1.state_next[3] ),
    .Q_N(_1228_),
    .Q(\top1.FSM1.state_reg[3] ));
 sg13g2_dfrbp_1 _2280_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net673),
    .D(\top1.FSM1.state_next[4] ),
    .Q_N(_0017_),
    .Q(\top1.FSM1.state_reg[4] ));
 sg13g2_dfrbp_1 _2281_ (.CLK(net610),
    .RESET_B(_0034_),
    .D(_0230_),
    .Q_N(_0032_),
    .Q(\top1.ch14c.data[0] ));
 sg13g2_dfrbp_1 _2282_ (.CLK(net610),
    .RESET_B(_0035_),
    .D(_0231_),
    .Q_N(_1212_),
    .Q(\top1.ch14c.data[1] ));
 sg13g2_dfrbp_1 _2283_ (.CLK(net610),
    .RESET_B(_0036_),
    .D(_0232_),
    .Q_N(_1211_),
    .Q(\top1.ch14c.data[2] ));
 sg13g2_dfrbp_1 _2284_ (.CLK(net610),
    .RESET_B(_0037_),
    .D(_0233_),
    .Q_N(_1210_),
    .Q(\top1.ch14c.data[3] ));
 sg13g2_dfrbp_1 _2285_ (.CLK(net610),
    .RESET_B(_0038_),
    .D(_0234_),
    .Q_N(_1209_),
    .Q(\top1.ch14c.data[4] ));
 sg13g2_dfrbp_1 _2286_ (.CLK(net611),
    .RESET_B(_0039_),
    .D(_0235_),
    .Q_N(_1208_),
    .Q(\top1.ch14c.data[5] ));
 sg13g2_dfrbp_1 _2287_ (.CLK(net610),
    .RESET_B(_0040_),
    .D(_0236_),
    .Q_N(_1207_),
    .Q(\top1.ch14c.data[6] ));
 sg13g2_dfrbp_1 _2288_ (.CLK(net611),
    .RESET_B(_0041_),
    .D(_0237_),
    .Q_N(_1206_),
    .Q(\top1.ch14c.data[7] ));
 sg13g2_dfrbp_1 _2289_ (.CLK(net611),
    .RESET_B(_0042_),
    .D(_0238_),
    .Q_N(_1205_),
    .Q(\top1.ch14c.data[8] ));
 sg13g2_dfrbp_1 _2290_ (.CLK(net610),
    .RESET_B(_0043_),
    .D(_0239_),
    .Q_N(_1204_),
    .Q(\top1.ch14c.data[9] ));
 sg13g2_dfrbp_1 _2291_ (.CLK(net610),
    .RESET_B(_0044_),
    .D(_0240_),
    .Q_N(_1203_),
    .Q(\top1.ch14c.data[10] ));
 sg13g2_dfrbp_1 _2292_ (.CLK(net611),
    .RESET_B(_0045_),
    .D(_0241_),
    .Q_N(_1202_),
    .Q(\top1.ch14c.data[11] ));
 sg13g2_dfrbp_1 _2293_ (.CLK(net612),
    .RESET_B(_0046_),
    .D(_0242_),
    .Q_N(_0031_),
    .Q(\top1.ch13c.data[0] ));
 sg13g2_dfrbp_1 _2294_ (.CLK(net612),
    .RESET_B(_0047_),
    .D(_0243_),
    .Q_N(_1201_),
    .Q(\top1.ch13c.data[1] ));
 sg13g2_dfrbp_1 _2295_ (.CLK(net612),
    .RESET_B(_0048_),
    .D(_0244_),
    .Q_N(_1200_),
    .Q(\top1.ch13c.data[2] ));
 sg13g2_dfrbp_1 _2296_ (.CLK(net612),
    .RESET_B(_0049_),
    .D(_0245_),
    .Q_N(_1199_),
    .Q(\top1.ch13c.data[3] ));
 sg13g2_dfrbp_1 _2297_ (.CLK(net613),
    .RESET_B(_0050_),
    .D(_0246_),
    .Q_N(_1198_),
    .Q(\top1.ch13c.data[4] ));
 sg13g2_dfrbp_1 _2298_ (.CLK(net613),
    .RESET_B(_0051_),
    .D(_0247_),
    .Q_N(_1197_),
    .Q(\top1.ch13c.data[5] ));
 sg13g2_dfrbp_1 _2299_ (.CLK(net612),
    .RESET_B(_0052_),
    .D(_0248_),
    .Q_N(_1196_),
    .Q(\top1.ch13c.data[6] ));
 sg13g2_dfrbp_1 _2300_ (.CLK(net612),
    .RESET_B(_0053_),
    .D(_0249_),
    .Q_N(_1195_),
    .Q(\top1.ch13c.data[7] ));
 sg13g2_dfrbp_1 _2301_ (.CLK(net613),
    .RESET_B(_0054_),
    .D(_0250_),
    .Q_N(_1194_),
    .Q(\top1.ch13c.data[8] ));
 sg13g2_dfrbp_1 _2302_ (.CLK(net613),
    .RESET_B(_0055_),
    .D(_0251_),
    .Q_N(_1193_),
    .Q(\top1.ch13c.data[9] ));
 sg13g2_dfrbp_1 _2303_ (.CLK(net612),
    .RESET_B(_0056_),
    .D(_0252_),
    .Q_N(_1192_),
    .Q(\top1.ch13c.data[10] ));
 sg13g2_dfrbp_1 _2304_ (.CLK(net613),
    .RESET_B(_0057_),
    .D(_0253_),
    .Q_N(_1191_),
    .Q(\top1.ch13c.data[11] ));
 sg13g2_dfrbp_1 _2305_ (.CLK(net614),
    .RESET_B(_0058_),
    .D(_0254_),
    .Q_N(_0030_),
    .Q(\top1.ch12c.data[0] ));
 sg13g2_dfrbp_1 _2306_ (.CLK(net614),
    .RESET_B(_0059_),
    .D(_0255_),
    .Q_N(_1190_),
    .Q(\top1.ch12c.data[1] ));
 sg13g2_dfrbp_1 _2307_ (.CLK(net614),
    .RESET_B(_0060_),
    .D(_0256_),
    .Q_N(_1189_),
    .Q(\top1.ch12c.data[2] ));
 sg13g2_dfrbp_1 _2308_ (.CLK(net614),
    .RESET_B(_0061_),
    .D(_0257_),
    .Q_N(_1188_),
    .Q(\top1.ch12c.data[3] ));
 sg13g2_dfrbp_1 _2309_ (.CLK(net615),
    .RESET_B(_0062_),
    .D(_0258_),
    .Q_N(_1187_),
    .Q(\top1.ch12c.data[4] ));
 sg13g2_dfrbp_1 _2310_ (.CLK(net614),
    .RESET_B(_0063_),
    .D(_0259_),
    .Q_N(_1186_),
    .Q(\top1.ch12c.data[5] ));
 sg13g2_dfrbp_1 _2311_ (.CLK(net614),
    .RESET_B(_0064_),
    .D(_0260_),
    .Q_N(_1185_),
    .Q(\top1.ch12c.data[6] ));
 sg13g2_dfrbp_1 _2312_ (.CLK(net614),
    .RESET_B(_0065_),
    .D(_0261_),
    .Q_N(_1184_),
    .Q(\top1.ch12c.data[7] ));
 sg13g2_dfrbp_1 _2313_ (.CLK(net614),
    .RESET_B(_0066_),
    .D(_0262_),
    .Q_N(_1183_),
    .Q(\top1.ch12c.data[8] ));
 sg13g2_dfrbp_1 _2314_ (.CLK(net615),
    .RESET_B(_0067_),
    .D(_0263_),
    .Q_N(_1182_),
    .Q(\top1.ch12c.data[9] ));
 sg13g2_dfrbp_1 _2315_ (.CLK(net615),
    .RESET_B(_0068_),
    .D(_0264_),
    .Q_N(_1181_),
    .Q(\top1.ch12c.data[10] ));
 sg13g2_dfrbp_1 _2316_ (.CLK(net615),
    .RESET_B(_0069_),
    .D(_0265_),
    .Q_N(_1180_),
    .Q(\top1.ch12c.data[11] ));
 sg13g2_dfrbp_1 _2317_ (.CLK(net616),
    .RESET_B(_0070_),
    .D(_0266_),
    .Q_N(_0029_),
    .Q(\top1.ch11c.data[0] ));
 sg13g2_dfrbp_1 _2318_ (.CLK(net616),
    .RESET_B(_0071_),
    .D(_0267_),
    .Q_N(_1179_),
    .Q(\top1.ch11c.data[1] ));
 sg13g2_dfrbp_1 _2319_ (.CLK(net616),
    .RESET_B(_0072_),
    .D(_0268_),
    .Q_N(_1178_),
    .Q(\top1.ch11c.data[2] ));
 sg13g2_dfrbp_1 _2320_ (.CLK(net616),
    .RESET_B(_0073_),
    .D(_0269_),
    .Q_N(_1177_),
    .Q(\top1.ch11c.data[3] ));
 sg13g2_dfrbp_1 _2321_ (.CLK(net616),
    .RESET_B(_0074_),
    .D(_0270_),
    .Q_N(_1176_),
    .Q(\top1.ch11c.data[4] ));
 sg13g2_dfrbp_1 _2322_ (.CLK(net617),
    .RESET_B(_0075_),
    .D(_0271_),
    .Q_N(_1175_),
    .Q(\top1.ch11c.data[5] ));
 sg13g2_dfrbp_1 _2323_ (.CLK(net617),
    .RESET_B(_0076_),
    .D(_0272_),
    .Q_N(_1174_),
    .Q(\top1.ch11c.data[6] ));
 sg13g2_dfrbp_1 _2324_ (.CLK(net617),
    .RESET_B(_0077_),
    .D(_0273_),
    .Q_N(_1173_),
    .Q(\top1.ch11c.data[7] ));
 sg13g2_dfrbp_1 _2325_ (.CLK(net617),
    .RESET_B(_0078_),
    .D(_0274_),
    .Q_N(_1172_),
    .Q(\top1.ch11c.data[8] ));
 sg13g2_dfrbp_1 _2326_ (.CLK(net616),
    .RESET_B(_0079_),
    .D(_0275_),
    .Q_N(_1171_),
    .Q(\top1.ch11c.data[9] ));
 sg13g2_dfrbp_1 _2327_ (.CLK(net616),
    .RESET_B(_0080_),
    .D(_0276_),
    .Q_N(_1170_),
    .Q(\top1.ch11c.data[10] ));
 sg13g2_dfrbp_1 _2328_ (.CLK(net617),
    .RESET_B(_0081_),
    .D(_0277_),
    .Q_N(_1169_),
    .Q(\top1.ch11c.data[11] ));
 sg13g2_dfrbp_1 _2329_ (.CLK(net618),
    .RESET_B(_0082_),
    .D(_0278_),
    .Q_N(_0028_),
    .Q(\top1.ch10c.data[0] ));
 sg13g2_dfrbp_1 _2330_ (.CLK(net618),
    .RESET_B(_0083_),
    .D(_0279_),
    .Q_N(_1168_),
    .Q(\top1.ch10c.data[1] ));
 sg13g2_dfrbp_1 _2331_ (.CLK(net618),
    .RESET_B(_0084_),
    .D(_0280_),
    .Q_N(_1167_),
    .Q(\top1.ch10c.data[2] ));
 sg13g2_dfrbp_1 _2332_ (.CLK(net619),
    .RESET_B(_0085_),
    .D(_0281_),
    .Q_N(_1166_),
    .Q(\top1.ch10c.data[3] ));
 sg13g2_dfrbp_1 _2333_ (.CLK(net619),
    .RESET_B(_0086_),
    .D(_0282_),
    .Q_N(_1165_),
    .Q(\top1.ch10c.data[4] ));
 sg13g2_dfrbp_1 _2334_ (.CLK(net618),
    .RESET_B(_0087_),
    .D(_0283_),
    .Q_N(_1164_),
    .Q(\top1.ch10c.data[5] ));
 sg13g2_dfrbp_1 _2335_ (.CLK(net619),
    .RESET_B(_0088_),
    .D(_0284_),
    .Q_N(_1163_),
    .Q(\top1.ch10c.data[6] ));
 sg13g2_dfrbp_1 _2336_ (.CLK(net619),
    .RESET_B(_0089_),
    .D(_0285_),
    .Q_N(_1162_),
    .Q(\top1.ch10c.data[7] ));
 sg13g2_dfrbp_1 _2337_ (.CLK(net619),
    .RESET_B(_0090_),
    .D(_0286_),
    .Q_N(_1161_),
    .Q(\top1.ch10c.data[8] ));
 sg13g2_dfrbp_1 _2338_ (.CLK(net618),
    .RESET_B(_0091_),
    .D(_0287_),
    .Q_N(_1160_),
    .Q(\top1.ch10c.data[9] ));
 sg13g2_dfrbp_1 _2339_ (.CLK(net618),
    .RESET_B(_0092_),
    .D(_0288_),
    .Q_N(_1159_),
    .Q(\top1.ch10c.data[10] ));
 sg13g2_dfrbp_1 _2340_ (.CLK(net618),
    .RESET_B(_0093_),
    .D(_0289_),
    .Q_N(_1158_),
    .Q(\top1.ch10c.data[11] ));
 sg13g2_dfrbp_1 _2341_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net29),
    .D(_0290_),
    .Q_N(_1157_),
    .Q(\top1.PISO_register1.register[10] ));
 sg13g2_dfrbp_1 _2342_ (.CLK(net622),
    .RESET_B(_0094_),
    .D(_0291_),
    .Q_N(_0027_),
    .Q(\top1.ch8c.data[0] ));
 sg13g2_dfrbp_1 _2343_ (.CLK(net622),
    .RESET_B(_0095_),
    .D(_0292_),
    .Q_N(_1156_),
    .Q(\top1.ch8c.data[1] ));
 sg13g2_dfrbp_1 _2344_ (.CLK(net622),
    .RESET_B(_0096_),
    .D(_0293_),
    .Q_N(_1155_),
    .Q(\top1.ch8c.data[2] ));
 sg13g2_dfrbp_1 _2345_ (.CLK(net622),
    .RESET_B(_0097_),
    .D(_0294_),
    .Q_N(_1154_),
    .Q(\top1.ch8c.data[3] ));
 sg13g2_dfrbp_1 _2346_ (.CLK(net622),
    .RESET_B(_0098_),
    .D(_0295_),
    .Q_N(_1153_),
    .Q(\top1.ch8c.data[4] ));
 sg13g2_dfrbp_1 _2347_ (.CLK(net622),
    .RESET_B(_0099_),
    .D(_0296_),
    .Q_N(_1152_),
    .Q(\top1.ch8c.data[5] ));
 sg13g2_dfrbp_1 _2348_ (.CLK(net622),
    .RESET_B(_0100_),
    .D(_0297_),
    .Q_N(_1151_),
    .Q(\top1.ch8c.data[6] ));
 sg13g2_dfrbp_1 _2349_ (.CLK(net623),
    .RESET_B(_0101_),
    .D(_0298_),
    .Q_N(_1150_),
    .Q(\top1.ch8c.data[7] ));
 sg13g2_dfrbp_1 _2350_ (.CLK(net622),
    .RESET_B(_0102_),
    .D(_0299_),
    .Q_N(_1149_),
    .Q(\top1.ch8c.data[8] ));
 sg13g2_dfrbp_1 _2351_ (.CLK(net623),
    .RESET_B(_0103_),
    .D(_0300_),
    .Q_N(_1148_),
    .Q(\top1.ch8c.data[9] ));
 sg13g2_dfrbp_1 _2352_ (.CLK(net623),
    .RESET_B(_0104_),
    .D(_0301_),
    .Q_N(_1147_),
    .Q(\top1.ch8c.data[10] ));
 sg13g2_dfrbp_1 _2353_ (.CLK(net623),
    .RESET_B(_0105_),
    .D(_0302_),
    .Q_N(_1146_),
    .Q(\top1.ch8c.data[11] ));
 sg13g2_dfrbp_1 _2354_ (.CLK(net624),
    .RESET_B(_0106_),
    .D(_0303_),
    .Q_N(_0026_),
    .Q(\top1.ch7c.data[0] ));
 sg13g2_dfrbp_1 _2355_ (.CLK(net624),
    .RESET_B(_0107_),
    .D(_0304_),
    .Q_N(_1145_),
    .Q(\top1.ch7c.data[1] ));
 sg13g2_dfrbp_1 _2356_ (.CLK(net624),
    .RESET_B(_0108_),
    .D(_0305_),
    .Q_N(_1144_),
    .Q(\top1.ch7c.data[2] ));
 sg13g2_dfrbp_1 _2357_ (.CLK(net624),
    .RESET_B(_0109_),
    .D(_0306_),
    .Q_N(_1143_),
    .Q(\top1.ch7c.data[3] ));
 sg13g2_dfrbp_1 _2358_ (.CLK(net624),
    .RESET_B(_0110_),
    .D(_0307_),
    .Q_N(_1142_),
    .Q(\top1.ch7c.data[4] ));
 sg13g2_dfrbp_1 _2359_ (.CLK(net624),
    .RESET_B(_0111_),
    .D(_0308_),
    .Q_N(_1141_),
    .Q(\top1.ch7c.data[5] ));
 sg13g2_dfrbp_1 _2360_ (.CLK(net624),
    .RESET_B(_0112_),
    .D(_0309_),
    .Q_N(_1140_),
    .Q(\top1.ch7c.data[6] ));
 sg13g2_dfrbp_1 _2361_ (.CLK(net624),
    .RESET_B(_0113_),
    .D(_0310_),
    .Q_N(_1139_),
    .Q(\top1.ch7c.data[7] ));
 sg13g2_dfrbp_1 _2362_ (.CLK(net625),
    .RESET_B(_0114_),
    .D(_0311_),
    .Q_N(_1138_),
    .Q(\top1.ch7c.data[8] ));
 sg13g2_dfrbp_1 _2363_ (.CLK(net625),
    .RESET_B(_0115_),
    .D(_0312_),
    .Q_N(_1137_),
    .Q(\top1.ch7c.data[9] ));
 sg13g2_dfrbp_1 _2364_ (.CLK(net625),
    .RESET_B(_0116_),
    .D(_0313_),
    .Q_N(_1136_),
    .Q(\top1.ch7c.data[10] ));
 sg13g2_dfrbp_1 _2365_ (.CLK(net625),
    .RESET_B(_0117_),
    .D(_0314_),
    .Q_N(_1135_),
    .Q(\top1.ch7c.data[11] ));
 sg13g2_dfrbp_1 _2366_ (.CLK(net626),
    .RESET_B(_0118_),
    .D(_0315_),
    .Q_N(_0025_),
    .Q(\top1.ch6c.data[0] ));
 sg13g2_dfrbp_1 _2367_ (.CLK(net626),
    .RESET_B(_0119_),
    .D(_0316_),
    .Q_N(_1134_),
    .Q(\top1.ch6c.data[1] ));
 sg13g2_dfrbp_1 _2368_ (.CLK(net626),
    .RESET_B(_0120_),
    .D(_0317_),
    .Q_N(_1133_),
    .Q(\top1.ch6c.data[2] ));
 sg13g2_dfrbp_1 _2369_ (.CLK(net626),
    .RESET_B(_0121_),
    .D(_0318_),
    .Q_N(_1132_),
    .Q(\top1.ch6c.data[3] ));
 sg13g2_dfrbp_1 _2370_ (.CLK(net626),
    .RESET_B(_0122_),
    .D(_0319_),
    .Q_N(_1131_),
    .Q(\top1.ch6c.data[4] ));
 sg13g2_dfrbp_1 _2371_ (.CLK(net626),
    .RESET_B(_0123_),
    .D(_0320_),
    .Q_N(_1130_),
    .Q(\top1.ch6c.data[5] ));
 sg13g2_dfrbp_1 _2372_ (.CLK(net626),
    .RESET_B(_0124_),
    .D(_0321_),
    .Q_N(_1129_),
    .Q(\top1.ch6c.data[6] ));
 sg13g2_dfrbp_1 _2373_ (.CLK(net627),
    .RESET_B(_0125_),
    .D(_0322_),
    .Q_N(_1128_),
    .Q(\top1.ch6c.data[7] ));
 sg13g2_dfrbp_1 _2374_ (.CLK(net627),
    .RESET_B(_0126_),
    .D(_0323_),
    .Q_N(_1127_),
    .Q(\top1.ch6c.data[8] ));
 sg13g2_dfrbp_1 _2375_ (.CLK(net627),
    .RESET_B(_0127_),
    .D(_0324_),
    .Q_N(_1126_),
    .Q(\top1.ch6c.data[9] ));
 sg13g2_dfrbp_1 _2376_ (.CLK(net627),
    .RESET_B(_0128_),
    .D(_0325_),
    .Q_N(_1125_),
    .Q(\top1.ch6c.data[10] ));
 sg13g2_dfrbp_1 _2377_ (.CLK(net627),
    .RESET_B(_0129_),
    .D(_0326_),
    .Q_N(_1124_),
    .Q(\top1.ch6c.data[11] ));
 sg13g2_dfrbp_1 _2378_ (.CLK(net629),
    .RESET_B(_0130_),
    .D(_0327_),
    .Q_N(_0024_),
    .Q(\top1.ch5c.data[0] ));
 sg13g2_dfrbp_1 _2379_ (.CLK(net629),
    .RESET_B(_0131_),
    .D(_0328_),
    .Q_N(_1123_),
    .Q(\top1.ch5c.data[1] ));
 sg13g2_dfrbp_1 _2380_ (.CLK(net628),
    .RESET_B(_0132_),
    .D(_0329_),
    .Q_N(_1122_),
    .Q(\top1.ch5c.data[2] ));
 sg13g2_dfrbp_1 _2381_ (.CLK(net628),
    .RESET_B(_0133_),
    .D(_0330_),
    .Q_N(_1121_),
    .Q(\top1.ch5c.data[3] ));
 sg13g2_dfrbp_1 _2382_ (.CLK(net628),
    .RESET_B(_0134_),
    .D(_0331_),
    .Q_N(_1120_),
    .Q(\top1.ch5c.data[4] ));
 sg13g2_dfrbp_1 _2383_ (.CLK(net628),
    .RESET_B(_0135_),
    .D(_0332_),
    .Q_N(_1119_),
    .Q(\top1.ch5c.data[5] ));
 sg13g2_dfrbp_1 _2384_ (.CLK(net628),
    .RESET_B(_0136_),
    .D(_0333_),
    .Q_N(_1118_),
    .Q(\top1.ch5c.data[6] ));
 sg13g2_dfrbp_1 _2385_ (.CLK(net628),
    .RESET_B(_0137_),
    .D(_0334_),
    .Q_N(_1117_),
    .Q(\top1.ch5c.data[7] ));
 sg13g2_dfrbp_1 _2386_ (.CLK(net629),
    .RESET_B(_0138_),
    .D(_0335_),
    .Q_N(_1116_),
    .Q(\top1.ch5c.data[8] ));
 sg13g2_dfrbp_1 _2387_ (.CLK(net629),
    .RESET_B(_0139_),
    .D(_0336_),
    .Q_N(_1115_),
    .Q(\top1.ch5c.data[9] ));
 sg13g2_dfrbp_1 _2388_ (.CLK(net629),
    .RESET_B(_0140_),
    .D(_0337_),
    .Q_N(_1114_),
    .Q(\top1.ch5c.data[10] ));
 sg13g2_dfrbp_1 _2389_ (.CLK(net628),
    .RESET_B(_0141_),
    .D(_0338_),
    .Q_N(_1113_),
    .Q(\top1.ch5c.data[11] ));
 sg13g2_dfrbp_1 _2390_ (.CLK(net630),
    .RESET_B(_0142_),
    .D(_0339_),
    .Q_N(_0023_),
    .Q(\top1.ch4c.data[0] ));
 sg13g2_dfrbp_1 _2391_ (.CLK(net630),
    .RESET_B(_0143_),
    .D(_0340_),
    .Q_N(_1112_),
    .Q(\top1.ch4c.data[1] ));
 sg13g2_dfrbp_1 _2392_ (.CLK(net630),
    .RESET_B(_0144_),
    .D(_0341_),
    .Q_N(_1111_),
    .Q(\top1.ch4c.data[2] ));
 sg13g2_dfrbp_1 _2393_ (.CLK(net630),
    .RESET_B(_0145_),
    .D(_0342_),
    .Q_N(_1110_),
    .Q(\top1.ch4c.data[3] ));
 sg13g2_dfrbp_1 _2394_ (.CLK(net631),
    .RESET_B(_0146_),
    .D(_0343_),
    .Q_N(_1109_),
    .Q(\top1.ch4c.data[4] ));
 sg13g2_dfrbp_1 _2395_ (.CLK(net631),
    .RESET_B(_0147_),
    .D(_0344_),
    .Q_N(_1108_),
    .Q(\top1.ch4c.data[5] ));
 sg13g2_dfrbp_1 _2396_ (.CLK(net631),
    .RESET_B(_0148_),
    .D(_0345_),
    .Q_N(_1107_),
    .Q(\top1.ch4c.data[6] ));
 sg13g2_dfrbp_1 _2397_ (.CLK(net630),
    .RESET_B(_0149_),
    .D(_0346_),
    .Q_N(_1106_),
    .Q(\top1.ch4c.data[7] ));
 sg13g2_dfrbp_1 _2398_ (.CLK(net630),
    .RESET_B(_0150_),
    .D(_0347_),
    .Q_N(_1105_),
    .Q(\top1.ch4c.data[8] ));
 sg13g2_dfrbp_1 _2399_ (.CLK(net630),
    .RESET_B(_0151_),
    .D(_0348_),
    .Q_N(_1104_),
    .Q(\top1.ch4c.data[9] ));
 sg13g2_dfrbp_1 _2400_ (.CLK(net630),
    .RESET_B(_0152_),
    .D(_0349_),
    .Q_N(_1103_),
    .Q(\top1.ch4c.data[10] ));
 sg13g2_dfrbp_1 _2401_ (.CLK(net631),
    .RESET_B(_0153_),
    .D(_0350_),
    .Q_N(_1102_),
    .Q(\top1.ch4c.data[11] ));
 sg13g2_dfrbp_1 _2402_ (.CLK(net632),
    .RESET_B(_0154_),
    .D(_0351_),
    .Q_N(_0022_),
    .Q(\top1.ch3c.data[0] ));
 sg13g2_dfrbp_1 _2403_ (.CLK(net632),
    .RESET_B(_0155_),
    .D(_0352_),
    .Q_N(_1101_),
    .Q(\top1.ch3c.data[1] ));
 sg13g2_dfrbp_1 _2404_ (.CLK(net632),
    .RESET_B(_0156_),
    .D(_0353_),
    .Q_N(_1100_),
    .Q(\top1.ch3c.data[2] ));
 sg13g2_dfrbp_1 _2405_ (.CLK(net632),
    .RESET_B(_0157_),
    .D(_0354_),
    .Q_N(_1099_),
    .Q(\top1.ch3c.data[3] ));
 sg13g2_dfrbp_1 _2406_ (.CLK(net632),
    .RESET_B(_0158_),
    .D(_0355_),
    .Q_N(_1098_),
    .Q(\top1.ch3c.data[4] ));
 sg13g2_dfrbp_1 _2407_ (.CLK(net633),
    .RESET_B(_0159_),
    .D(_0356_),
    .Q_N(_1097_),
    .Q(\top1.ch3c.data[5] ));
 sg13g2_dfrbp_1 _2408_ (.CLK(net632),
    .RESET_B(_0160_),
    .D(_0357_),
    .Q_N(_1096_),
    .Q(\top1.ch3c.data[6] ));
 sg13g2_dfrbp_1 _2409_ (.CLK(net633),
    .RESET_B(_0161_),
    .D(_0358_),
    .Q_N(_1095_),
    .Q(\top1.ch3c.data[7] ));
 sg13g2_dfrbp_1 _2410_ (.CLK(net633),
    .RESET_B(_0162_),
    .D(_0359_),
    .Q_N(_1094_),
    .Q(\top1.ch3c.data[8] ));
 sg13g2_dfrbp_1 _2411_ (.CLK(net633),
    .RESET_B(_0163_),
    .D(_0360_),
    .Q_N(_1093_),
    .Q(\top1.ch3c.data[9] ));
 sg13g2_dfrbp_1 _2412_ (.CLK(net633),
    .RESET_B(_0164_),
    .D(_0361_),
    .Q_N(_1092_),
    .Q(\top1.ch3c.data[10] ));
 sg13g2_dfrbp_1 _2413_ (.CLK(net632),
    .RESET_B(_0165_),
    .D(_0362_),
    .Q_N(_1091_),
    .Q(\top1.ch3c.data[11] ));
 sg13g2_dfrbp_1 _2414_ (.CLK(net634),
    .RESET_B(_0166_),
    .D(_0363_),
    .Q_N(_0021_),
    .Q(\top1.ch2c.data[0] ));
 sg13g2_dfrbp_1 _2415_ (.CLK(net634),
    .RESET_B(_0167_),
    .D(_0364_),
    .Q_N(_1090_),
    .Q(\top1.ch2c.data[1] ));
 sg13g2_dfrbp_1 _2416_ (.CLK(net634),
    .RESET_B(_0168_),
    .D(_0365_),
    .Q_N(_1089_),
    .Q(\top1.ch2c.data[2] ));
 sg13g2_dfrbp_1 _2417_ (.CLK(net635),
    .RESET_B(_0169_),
    .D(_0366_),
    .Q_N(_1088_),
    .Q(\top1.ch2c.data[3] ));
 sg13g2_dfrbp_1 _2418_ (.CLK(net634),
    .RESET_B(_0170_),
    .D(_0367_),
    .Q_N(_1087_),
    .Q(\top1.ch2c.data[4] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(net634),
    .RESET_B(_0171_),
    .D(_0368_),
    .Q_N(_1086_),
    .Q(\top1.ch2c.data[5] ));
 sg13g2_dfrbp_1 _2420_ (.CLK(net635),
    .RESET_B(_0172_),
    .D(_0369_),
    .Q_N(_1085_),
    .Q(\top1.ch2c.data[6] ));
 sg13g2_dfrbp_1 _2421_ (.CLK(net635),
    .RESET_B(_0173_),
    .D(_0370_),
    .Q_N(_1084_),
    .Q(\top1.ch2c.data[7] ));
 sg13g2_dfrbp_1 _2422_ (.CLK(net634),
    .RESET_B(_0174_),
    .D(_0371_),
    .Q_N(_1083_),
    .Q(\top1.ch2c.data[8] ));
 sg13g2_dfrbp_1 _2423_ (.CLK(net635),
    .RESET_B(_0175_),
    .D(_0372_),
    .Q_N(_1082_),
    .Q(\top1.ch2c.data[9] ));
 sg13g2_dfrbp_1 _2424_ (.CLK(net634),
    .RESET_B(_0176_),
    .D(_0373_),
    .Q_N(_1081_),
    .Q(\top1.ch2c.data[10] ));
 sg13g2_dfrbp_1 _2425_ (.CLK(net634),
    .RESET_B(_0177_),
    .D(_0374_),
    .Q_N(_1080_),
    .Q(\top1.ch2c.data[11] ));
 sg13g2_dfrbp_1 _2426_ (.CLK(net636),
    .RESET_B(_0178_),
    .D(_0375_),
    .Q_N(_0020_),
    .Q(\top1.ch1c.data[0] ));
 sg13g2_dfrbp_1 _2427_ (.CLK(net637),
    .RESET_B(_0179_),
    .D(_0376_),
    .Q_N(_1079_),
    .Q(\top1.ch1c.data[1] ));
 sg13g2_dfrbp_1 _2428_ (.CLK(net637),
    .RESET_B(_0180_),
    .D(_0377_),
    .Q_N(_1078_),
    .Q(\top1.ch1c.data[2] ));
 sg13g2_dfrbp_1 _2429_ (.CLK(net636),
    .RESET_B(_0181_),
    .D(_0378_),
    .Q_N(_1077_),
    .Q(\top1.ch1c.data[3] ));
 sg13g2_dfrbp_1 _2430_ (.CLK(net637),
    .RESET_B(_0182_),
    .D(_0379_),
    .Q_N(_1076_),
    .Q(\top1.ch1c.data[4] ));
 sg13g2_dfrbp_1 _2431_ (.CLK(net637),
    .RESET_B(_0183_),
    .D(_0380_),
    .Q_N(_1075_),
    .Q(\top1.ch1c.data[5] ));
 sg13g2_dfrbp_1 _2432_ (.CLK(net636),
    .RESET_B(_0184_),
    .D(_0381_),
    .Q_N(_1074_),
    .Q(\top1.ch1c.data[6] ));
 sg13g2_dfrbp_1 _2433_ (.CLK(net637),
    .RESET_B(_0185_),
    .D(_0382_),
    .Q_N(_1073_),
    .Q(\top1.ch1c.data[7] ));
 sg13g2_dfrbp_1 _2434_ (.CLK(net636),
    .RESET_B(_0186_),
    .D(_0383_),
    .Q_N(_1072_),
    .Q(\top1.ch1c.data[8] ));
 sg13g2_dfrbp_1 _2435_ (.CLK(net636),
    .RESET_B(_0187_),
    .D(_0384_),
    .Q_N(_1071_),
    .Q(\top1.ch1c.data[9] ));
 sg13g2_dfrbp_1 _2436_ (.CLK(net636),
    .RESET_B(_0188_),
    .D(_0385_),
    .Q_N(_1070_),
    .Q(\top1.ch1c.data[10] ));
 sg13g2_dfrbp_1 _2437_ (.CLK(net636),
    .RESET_B(_0189_),
    .D(_0386_),
    .Q_N(_1069_),
    .Q(\top1.ch1c.data[11] ));
 sg13g2_dfrbp_1 _2438_ (.CLK(net608),
    .RESET_B(_0190_),
    .D(_0387_),
    .Q_N(_0019_),
    .Q(\top1.ch15c.data[0] ));
 sg13g2_dfrbp_1 _2439_ (.CLK(net608),
    .RESET_B(_0191_),
    .D(_0388_),
    .Q_N(_1068_),
    .Q(\top1.ch15c.data[1] ));
 sg13g2_dfrbp_1 _2440_ (.CLK(net608),
    .RESET_B(_0192_),
    .D(_0389_),
    .Q_N(_1067_),
    .Q(\top1.ch15c.data[2] ));
 sg13g2_dfrbp_1 _2441_ (.CLK(net608),
    .RESET_B(_0193_),
    .D(_0390_),
    .Q_N(_1066_),
    .Q(\top1.ch15c.data[3] ));
 sg13g2_dfrbp_1 _2442_ (.CLK(net609),
    .RESET_B(_0194_),
    .D(_0391_),
    .Q_N(_1065_),
    .Q(\top1.ch15c.data[4] ));
 sg13g2_dfrbp_1 _2443_ (.CLK(net608),
    .RESET_B(_0195_),
    .D(_0392_),
    .Q_N(_1064_),
    .Q(\top1.ch15c.data[5] ));
 sg13g2_dfrbp_1 _2444_ (.CLK(net608),
    .RESET_B(_0196_),
    .D(_0393_),
    .Q_N(_1063_),
    .Q(\top1.ch15c.data[6] ));
 sg13g2_dfrbp_1 _2445_ (.CLK(net609),
    .RESET_B(_0197_),
    .D(_0394_),
    .Q_N(_1062_),
    .Q(\top1.ch15c.data[7] ));
 sg13g2_dfrbp_1 _2446_ (.CLK(net609),
    .RESET_B(_0198_),
    .D(_0395_),
    .Q_N(_1061_),
    .Q(\top1.ch15c.data[8] ));
 sg13g2_dfrbp_1 _2447_ (.CLK(net609),
    .RESET_B(_0199_),
    .D(_0396_),
    .Q_N(_1060_),
    .Q(\top1.ch15c.data[9] ));
 sg13g2_dfrbp_1 _2448_ (.CLK(net608),
    .RESET_B(_0200_),
    .D(_0397_),
    .Q_N(_1059_),
    .Q(\top1.ch15c.data[10] ));
 sg13g2_dfrbp_1 _2449_ (.CLK(net608),
    .RESET_B(_0201_),
    .D(_0398_),
    .Q_N(_1058_),
    .Q(\top1.ch15c.data[11] ));
 sg13g2_dfrbp_1 _2450_ (.CLK(net638),
    .RESET_B(net667),
    .D(_0399_),
    .Q_N(_1057_),
    .Q(\top1.data[0][6] ));
 sg13g2_dfrbp_1 _2451_ (.CLK(net638),
    .RESET_B(net667),
    .D(_0400_),
    .Q_N(_1056_),
    .Q(\top1.data[0][7] ));
 sg13g2_dfrbp_1 _2452_ (.CLK(net639),
    .RESET_B(net667),
    .D(_0401_),
    .Q_N(_1055_),
    .Q(\top1.data[0][8] ));
 sg13g2_dfrbp_1 _2453_ (.CLK(net639),
    .RESET_B(net667),
    .D(_0402_),
    .Q_N(_1054_),
    .Q(\top1.data[0][9] ));
 sg13g2_dfrbp_1 _2454_ (.CLK(net639),
    .RESET_B(net667),
    .D(_0403_),
    .Q_N(_1053_),
    .Q(\top1.data[0][10] ));
 sg13g2_dfrbp_1 _2455_ (.CLK(net639),
    .RESET_B(net667),
    .D(_0404_),
    .Q_N(_1052_),
    .Q(\top1.data[0][11] ));
 sg13g2_dfrbp_1 _2456_ (.CLK(net621),
    .RESET_B(_0202_),
    .D(_0405_),
    .Q_N(_0018_),
    .Q(\top1.ch9c.data[0] ));
 sg13g2_dfrbp_1 _2457_ (.CLK(net620),
    .RESET_B(_0203_),
    .D(_0406_),
    .Q_N(_1051_),
    .Q(\top1.ch9c.data[1] ));
 sg13g2_dfrbp_1 _2458_ (.CLK(net620),
    .RESET_B(_0204_),
    .D(_0407_),
    .Q_N(_1050_),
    .Q(\top1.ch9c.data[2] ));
 sg13g2_dfrbp_1 _2459_ (.CLK(net620),
    .RESET_B(_0205_),
    .D(_0408_),
    .Q_N(_1049_),
    .Q(\top1.ch9c.data[3] ));
 sg13g2_dfrbp_1 _2460_ (.CLK(net620),
    .RESET_B(_0206_),
    .D(_0409_),
    .Q_N(_1048_),
    .Q(\top1.ch9c.data[4] ));
 sg13g2_dfrbp_1 _2461_ (.CLK(net620),
    .RESET_B(_0207_),
    .D(_0410_),
    .Q_N(_1047_),
    .Q(\top1.ch9c.data[5] ));
 sg13g2_dfrbp_1 _2462_ (.CLK(net620),
    .RESET_B(_0208_),
    .D(_0411_),
    .Q_N(_1046_),
    .Q(\top1.ch9c.data[6] ));
 sg13g2_dfrbp_1 _2463_ (.CLK(net620),
    .RESET_B(_0209_),
    .D(_0412_),
    .Q_N(_1045_),
    .Q(\top1.ch9c.data[7] ));
 sg13g2_dfrbp_1 _2464_ (.CLK(net620),
    .RESET_B(_0210_),
    .D(_0413_),
    .Q_N(_1044_),
    .Q(\top1.ch9c.data[8] ));
 sg13g2_dfrbp_1 _2465_ (.CLK(net621),
    .RESET_B(_0211_),
    .D(_0414_),
    .Q_N(_1043_),
    .Q(\top1.ch9c.data[9] ));
 sg13g2_dfrbp_1 _2466_ (.CLK(net621),
    .RESET_B(_0212_),
    .D(_0415_),
    .Q_N(_1042_),
    .Q(\top1.ch9c.data[10] ));
 sg13g2_dfrbp_1 _2467_ (.CLK(net621),
    .RESET_B(_0213_),
    .D(_0416_),
    .Q_N(_1229_),
    .Q(\top1.ch9c.data[11] ));
 sg13g2_dfrbp_1 _2468_ (.CLK(net638),
    .RESET_B(net665),
    .D(_0011_),
    .Q_N(_1230_),
    .Q(\top1.data[0][0] ));
 sg13g2_dfrbp_1 _2469_ (.CLK(net638),
    .RESET_B(net665),
    .D(_0012_),
    .Q_N(_1231_),
    .Q(\top1.data[0][1] ));
 sg13g2_dfrbp_1 _2470_ (.CLK(net638),
    .RESET_B(net665),
    .D(_0013_),
    .Q_N(_1232_),
    .Q(\top1.data[0][2] ));
 sg13g2_dfrbp_1 _2471_ (.CLK(net638),
    .RESET_B(net666),
    .D(_0014_),
    .Q_N(_1233_),
    .Q(\top1.data[0][3] ));
 sg13g2_dfrbp_1 _2472_ (.CLK(net638),
    .RESET_B(net665),
    .D(_0015_),
    .Q_N(_1234_),
    .Q(\top1.data[0][4] ));
 sg13g2_dfrbp_1 _2473_ (.CLK(net638),
    .RESET_B(net665),
    .D(_0016_),
    .Q_N(_1041_),
    .Q(\top1.data[0][5] ));
 sg13g2_dfrbp_1 _2474_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net672),
    .D(_0417_),
    .Q_N(_1040_),
    .Q(\top1.FSM1.counter_register[0] ));
 sg13g2_dfrbp_1 _2475_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net672),
    .D(_0418_),
    .Q_N(_1039_),
    .Q(\top1.FSM1.counter_register[1] ));
 sg13g2_dfrbp_1 _2476_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net672),
    .D(net50),
    .Q_N(_1038_),
    .Q(\top1.FSM1.counter_register[2] ));
 sg13g2_dfrbp_1 _2477_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net672),
    .D(net44),
    .Q_N(_1037_),
    .Q(\top1.FSM1.counter_register[3] ));
 sg13g2_dfrbp_1 _2478_ (.CLK(net609),
    .RESET_B(_0214_),
    .D(_0421_),
    .Q_N(_1036_),
    .Q(\top1.ch15c.ovf ));
 sg13g2_dfrbp_1 _2479_ (.CLK(net611),
    .RESET_B(_0215_),
    .D(_0422_),
    .Q_N(_1035_),
    .Q(\top1.ch14c.ovf ));
 sg13g2_dfrbp_1 _2480_ (.CLK(net612),
    .RESET_B(_0216_),
    .D(_0423_),
    .Q_N(_1034_),
    .Q(\top1.ch13c.ovf ));
 sg13g2_dfrbp_1 _2481_ (.CLK(net615),
    .RESET_B(_0217_),
    .D(_0424_),
    .Q_N(_1033_),
    .Q(\top1.ch12c.ovf ));
 sg13g2_dfrbp_1 _2482_ (.CLK(net616),
    .RESET_B(_0218_),
    .D(_0425_),
    .Q_N(_1032_),
    .Q(\top1.ch11c.ovf ));
 sg13g2_dfrbp_1 _2483_ (.CLK(net618),
    .RESET_B(_0219_),
    .D(_0426_),
    .Q_N(_1031_),
    .Q(\top1.ch10c.ovf ));
 sg13g2_dfrbp_1 _2484_ (.CLK(net621),
    .RESET_B(_0220_),
    .D(_0427_),
    .Q_N(_1030_),
    .Q(\top1.ch9c.ovf ));
 sg13g2_dfrbp_1 _2485_ (.CLK(net623),
    .RESET_B(_0221_),
    .D(_0428_),
    .Q_N(_1029_),
    .Q(\top1.ch8c.ovf ));
 sg13g2_dfrbp_1 _2486_ (.CLK(net625),
    .RESET_B(_0222_),
    .D(_0429_),
    .Q_N(_1028_),
    .Q(\top1.ch7c.ovf ));
 sg13g2_dfrbp_1 _2487_ (.CLK(net626),
    .RESET_B(_0223_),
    .D(_0430_),
    .Q_N(_1027_),
    .Q(\top1.ch6c.ovf ));
 sg13g2_dfrbp_1 _2488_ (.CLK(net628),
    .RESET_B(_0224_),
    .D(_0431_),
    .Q_N(_1026_),
    .Q(\top1.ch5c.ovf ));
 sg13g2_dfrbp_1 _2489_ (.CLK(net1),
    .RESET_B(_0225_),
    .D(_0432_),
    .Q_N(_1025_),
    .Q(\top1.ch4c.ovf ));
 sg13g2_dfrbp_1 _2490_ (.CLK(net632),
    .RESET_B(_0226_),
    .D(_0433_),
    .Q_N(_1024_),
    .Q(\top1.ch3c.ovf ));
 sg13g2_dfrbp_1 _2491_ (.CLK(net635),
    .RESET_B(_0227_),
    .D(_0434_),
    .Q_N(_1023_),
    .Q(\top1.ch2c.ovf ));
 sg13g2_dfrbp_1 _2492_ (.CLK(net636),
    .RESET_B(_0228_),
    .D(_0435_),
    .Q_N(_1022_),
    .Q(\top1.ch1c.ovf ));
 sg13g2_tiehi _2266__19 (.L_HI(net19));
 sg13g2_tiehi _2267__20 (.L_HI(net20));
 sg13g2_tiehi _2268__21 (.L_HI(net21));
 sg13g2_tiehi _2269__22 (.L_HI(net22));
 sg13g2_tiehi _2270__23 (.L_HI(net23));
 sg13g2_tiehi _2271__24 (.L_HI(net24));
 sg13g2_tiehi _2272__25 (.L_HI(net25));
 sg13g2_tiehi _2273__26 (.L_HI(net26));
 sg13g2_tiehi _2274__27 (.L_HI(net27));
 sg13g2_tiehi _2275__28 (.L_HI(net28));
 sg13g2_tiehi _2341__29 (.L_HI(net29));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_Coline3003_top_3 (.L_LO(net3));
 sg13g2_tielo tt_um_Coline3003_top_4 (.L_LO(net4));
 sg13g2_tielo tt_um_Coline3003_top_5 (.L_LO(net5));
 sg13g2_tielo tt_um_Coline3003_top_6 (.L_LO(net6));
 sg13g2_tielo tt_um_Coline3003_top_7 (.L_LO(net7));
 sg13g2_tielo tt_um_Coline3003_top_8 (.L_LO(net8));
 sg13g2_tielo tt_um_Coline3003_top_9 (.L_LO(net9));
 sg13g2_tielo tt_um_Coline3003_top_10 (.L_LO(net10));
 sg13g2_tielo tt_um_Coline3003_top_11 (.L_LO(net11));
 sg13g2_tielo tt_um_Coline3003_top_12 (.L_LO(net12));
 sg13g2_tielo tt_um_Coline3003_top_13 (.L_LO(net13));
 sg13g2_tielo tt_um_Coline3003_top_14 (.L_LO(net14));
 sg13g2_tielo tt_um_Coline3003_top_15 (.L_LO(net15));
 sg13g2_tielo tt_um_Coline3003_top_16 (.L_LO(net16));
 sg13g2_tielo tt_um_Coline3003_top_17 (.L_LO(net17));
 sg13g2_tiehi _2265__18 (.L_HI(net18));
 sg13g2_buf_1 _2521_ (.A(\top1.PISO_register1.serial_out ),
    .X(uo_out[0]));
 sg13g2_buf_1 _2522_ (.A(net539),
    .X(uo_out[1]));
 sg13g2_buf_2 _2523_ (.A(\top1.ovf_RTC ),
    .X(uo_out[2]));
 sg13g2_buf_2 _2524_ (.A(\top1.a0_out ),
    .X(uo_out[3]));
 sg13g2_buf_2 _2525_ (.A(\top1.a1_out ),
    .X(uo_out[4]));
 sg13g2_buf_2 _2526_ (.A(\top1.a2_out ),
    .X(uo_out[5]));
 sg13g2_buf_2 _2527_ (.A(\top1.a3_out ),
    .X(uo_out[6]));
 sg13g2_buf_1 _2528_ (.A(\top1.FSM1.SL ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout509 (.A(\top1.FSM1.SL ),
    .X(net509));
 sg13g2_buf_1 fanout510 (.A(\top1.FSM1.SL ),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net512),
    .X(net511));
 sg13g2_buf_1 fanout512 (.A(_0578_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net514),
    .X(net513));
 sg13g2_buf_1 fanout514 (.A(_0576_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(net516),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_0569_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_0569_),
    .X(net517));
 sg13g2_buf_1 fanout518 (.A(_0569_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_0567_),
    .X(net519));
 sg13g2_buf_1 fanout520 (.A(_0567_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_0581_),
    .X(net521));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(net523));
 sg13g2_buf_2 fanout523 (.A(_0580_),
    .X(net523));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(net525));
 sg13g2_buf_2 fanout525 (.A(_0573_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(net527),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_0572_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_0570_),
    .X(net528));
 sg13g2_buf_1 fanout529 (.A(_0570_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(net531),
    .X(net530));
 sg13g2_buf_1 fanout531 (.A(net532),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_0563_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_0588_),
    .X(net534));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(net538));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net537));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(net538));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(net541));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(net541));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(net541));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(\top1.FSM1.ovf ));
 sg13g2_buf_2 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_1 fanout543 (.A(net549),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(net546),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net546),
    .X(net545));
 sg13g2_buf_1 fanout546 (.A(net549),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net549),
    .X(net547));
 sg13g2_buf_1 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(net577),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net552),
    .X(net550));
 sg13g2_buf_1 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(net555),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net555),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(net577),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net560),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(net560),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net560),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(net560),
    .X(net559));
 sg13g2_buf_1 fanout560 (.A(net577),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net565),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net565),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(net565),
    .X(net563));
 sg13g2_buf_1 fanout564 (.A(net565),
    .X(net564));
 sg13g2_buf_1 fanout565 (.A(net576),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(net576),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net571),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net576),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net575),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_0782_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_0589_),
    .X(net579));
 sg13g2_buf_4 fanout580 (.X(net580),
    .A(net581));
 sg13g2_buf_2 fanout581 (.A(_0587_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_0585_),
    .X(net583));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(net585));
 sg13g2_buf_2 fanout585 (.A(_0583_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_1 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_0552_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(_0551_));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_1 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_1 fanout593 (.A(_0540_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(net596),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(net596),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(net599),
    .X(net596));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(net599));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_0933_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_0017_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(\top1.FSM1.state_reg[3] ),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(\top1.FSM1.state_reg[2] ),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(\top1.FSM1.state_reg[2] ),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(\top1.FSM1.state_reg[1] ),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(\top1.FSM1.state_reg[0] ),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(\top1.FSM1.state_reg[0] ),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(uio_in[7]),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(uio_in[7]),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(uio_in[6]),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(uio_in[6]),
    .X(net611));
 sg13g2_buf_4 fanout612 (.X(net612),
    .A(uio_in[5]));
 sg13g2_buf_1 fanout613 (.A(uio_in[5]),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(uio_in[4]),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(uio_in[3]),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(uio_in[3]),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(uio_in[2]),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(uio_in[2]),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(uio_in[1]),
    .X(net620));
 sg13g2_buf_1 fanout621 (.A(uio_in[1]),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(uio_in[0]),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(ui_in[7]),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(ui_in[7]),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(ui_in[6]),
    .X(net626));
 sg13g2_buf_1 fanout627 (.A(ui_in[6]),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(ui_in[5]),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(ui_in[5]),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(net631),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(net1),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(ui_in[3]),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(ui_in[3]),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(ui_in[2]),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(ui_in[1]),
    .X(net636));
 sg13g2_buf_1 fanout637 (.A(ui_in[1]),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(ui_in[0]),
    .X(net638));
 sg13g2_buf_1 fanout639 (.A(ui_in[0]),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_1 fanout641 (.A(net647),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(net644),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_1 fanout644 (.A(net647),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(net647),
    .X(net645));
 sg13g2_buf_1 fanout646 (.A(net647),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(net678),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(net650),
    .X(net648));
 sg13g2_buf_1 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(net653),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(net653),
    .X(net651));
 sg13g2_buf_1 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(net678),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(net658),
    .X(net654));
 sg13g2_buf_1 fanout655 (.A(net658),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(net658),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_1 fanout658 (.A(net678),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(net663),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net663),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(net663),
    .X(net661));
 sg13g2_buf_1 fanout662 (.A(net663),
    .X(net662));
 sg13g2_buf_1 fanout663 (.A(net678),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net666),
    .X(net664));
 sg13g2_buf_4 fanout665 (.X(net665),
    .A(net666));
 sg13g2_buf_2 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(net678));
 sg13g2_buf_2 fanout668 (.A(net671),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_1 fanout671 (.A(net677),
    .X(net671));
 sg13g2_buf_4 fanout672 (.X(net672),
    .A(net673));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(net677));
 sg13g2_buf_2 fanout674 (.A(net675),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(net676),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_tielo tt_um_Coline3003_top_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\top1.PISO_register1.register[7] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold2 (.A(\top1.PISO_register1.register[3] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold3 (.A(\top1.PISO_register1.register[5] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold4 (.A(\top1.PISO_register1.register[8] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold5 (.A(\top1.PISO_register1.register[1] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold6 (.A(\top1.PISO_register1.register[9] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold7 (.A(\top1.PISO_register1.register[2] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold8 (.A(\top1.PISO_register1.register[6] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold9 (.A(\top1.PISO_register1.register[10] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold10 (.A(\top1.PISO_register1.register[4] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold11 (.A(\top1.PISO_register1.register[0] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold12 (.A(\top1.FSM1.counter_register[1] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0804_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold14 (.A(\top1.FSM1.counter_register[3] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0420_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold16 (.A(\top1.FSM1.counter_register[0] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0017_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0771_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold19 (.A(\top1.FSM1.state_next[0] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold20 (.A(\top1.FSM1.counter_register[2] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0419_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold22 (.A(\top1.FSM1.counter_register[3] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold23 (.A(\top1.FSM1.state_reg[0] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0769_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold25 (.A(\top1.FSM1.counter_register[0] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold26 (.A(\top1.FSM1.counter_register[0] ),
    .X(net55));
 sg13g2_antennanp ANTENNA_1 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_2 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_3 (.A(uio_in[4]));
 sg13g2_antennanp ANTENNA_4 (.A(uio_in[4]));
 sg13g2_antennanp ANTENNA_5 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_6 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_7 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_8 (.A(uio_in[0]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_4 FILLER_12_301 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_fill_1 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_4 FILLER_14_301 ();
 sg13g2_fill_2 FILLER_14_313 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_4 FILLER_15_273 ();
 sg13g2_fill_2 FILLER_15_277 ();
 sg13g2_fill_2 FILLER_15_305 ();
 sg13g2_fill_1 FILLER_15_307 ();
 sg13g2_decap_4 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_4 FILLER_16_266 ();
 sg13g2_fill_1 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_211 ();
 sg13g2_decap_8 FILLER_18_218 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_239 ();
 sg13g2_decap_8 FILLER_18_246 ();
 sg13g2_decap_8 FILLER_18_253 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_decap_4 FILLER_18_267 ();
 sg13g2_fill_1 FILLER_18_271 ();
 sg13g2_fill_1 FILLER_18_300 ();
 sg13g2_fill_2 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_fill_2 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_fill_2 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_198 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_decap_8 FILLER_19_236 ();
 sg13g2_decap_8 FILLER_19_243 ();
 sg13g2_decap_8 FILLER_19_250 ();
 sg13g2_decap_8 FILLER_19_257 ();
 sg13g2_decap_8 FILLER_19_264 ();
 sg13g2_decap_8 FILLER_19_271 ();
 sg13g2_decap_4 FILLER_19_282 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_decap_8 FILLER_19_293 ();
 sg13g2_decap_8 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_314 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_4 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_decap_8 FILLER_20_260 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_decap_4 FILLER_20_288 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_fill_2 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_259 ();
 sg13g2_decap_4 FILLER_21_317 ();
 sg13g2_fill_2 FILLER_21_321 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_fill_2 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_359 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_208 ();
 sg13g2_fill_1 FILLER_22_215 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_254 ();
 sg13g2_decap_4 FILLER_22_294 ();
 sg13g2_fill_2 FILLER_22_308 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_decap_4 FILLER_22_324 ();
 sg13g2_decap_8 FILLER_22_332 ();
 sg13g2_decap_8 FILLER_22_339 ();
 sg13g2_fill_2 FILLER_22_346 ();
 sg13g2_fill_1 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_fill_2 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_230 ();
 sg13g2_decap_8 FILLER_23_237 ();
 sg13g2_decap_8 FILLER_23_244 ();
 sg13g2_decap_8 FILLER_23_251 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_4 FILLER_23_291 ();
 sg13g2_decap_4 FILLER_23_304 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_decap_4 FILLER_23_320 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_4 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_171 ();
 sg13g2_decap_8 FILLER_24_178 ();
 sg13g2_decap_4 FILLER_24_185 ();
 sg13g2_fill_1 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_240 ();
 sg13g2_decap_8 FILLER_24_247 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_284 ();
 sg13g2_fill_1 FILLER_24_291 ();
 sg13g2_fill_2 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_306 ();
 sg13g2_fill_1 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_153 ();
 sg13g2_fill_2 FILLER_25_194 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_decap_8 FILLER_25_247 ();
 sg13g2_fill_2 FILLER_25_254 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_decap_4 FILLER_25_283 ();
 sg13g2_fill_1 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_fill_2 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_123 ();
 sg13g2_decap_4 FILLER_26_156 ();
 sg13g2_fill_2 FILLER_26_160 ();
 sg13g2_decap_4 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_decap_4 FILLER_26_218 ();
 sg13g2_fill_2 FILLER_26_227 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_decap_8 FILLER_26_253 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_fill_2 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_fill_1 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_192 ();
 sg13g2_decap_8 FILLER_27_199 ();
 sg13g2_decap_4 FILLER_27_206 ();
 sg13g2_fill_2 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_4 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_254 ();
 sg13g2_decap_8 FILLER_27_265 ();
 sg13g2_fill_2 FILLER_27_272 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_decap_4 FILLER_27_285 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_4 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_139 ();
 sg13g2_decap_8 FILLER_28_146 ();
 sg13g2_decap_8 FILLER_28_153 ();
 sg13g2_decap_8 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_fill_1 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_decap_4 FILLER_28_309 ();
 sg13g2_decap_4 FILLER_28_319 ();
 sg13g2_fill_2 FILLER_28_323 ();
 sg13g2_fill_2 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_338 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_4 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_142 ();
 sg13g2_decap_4 FILLER_29_149 ();
 sg13g2_fill_2 FILLER_29_153 ();
 sg13g2_fill_2 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_decap_4 FILLER_29_184 ();
 sg13g2_fill_1 FILLER_29_188 ();
 sg13g2_fill_2 FILLER_29_299 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_decap_4 FILLER_29_312 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_334 ();
 sg13g2_decap_4 FILLER_29_341 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_fill_2 FILLER_30_126 ();
 sg13g2_decap_4 FILLER_30_154 ();
 sg13g2_decap_4 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_188 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_245 ();
 sg13g2_fill_1 FILLER_30_251 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_4 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_decap_8 FILLER_31_190 ();
 sg13g2_decap_4 FILLER_31_201 ();
 sg13g2_fill_1 FILLER_31_205 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_4 FILLER_31_245 ();
 sg13g2_fill_2 FILLER_31_249 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_fill_2 FILLER_31_269 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_decap_8 FILLER_32_205 ();
 sg13g2_decap_8 FILLER_32_212 ();
 sg13g2_decap_8 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_226 ();
 sg13g2_fill_1 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_244 ();
 sg13g2_decap_8 FILLER_32_251 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_265 ();
 sg13g2_decap_4 FILLER_32_272 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_fill_2 FILLER_32_282 ();
 sg13g2_fill_1 FILLER_32_284 ();
 sg13g2_decap_4 FILLER_32_298 ();
 sg13g2_decap_4 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_356 ();
 sg13g2_fill_1 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_4 FILLER_33_126 ();
 sg13g2_fill_2 FILLER_33_130 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_decap_4 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_181 ();
 sg13g2_decap_4 FILLER_33_188 ();
 sg13g2_decap_8 FILLER_33_197 ();
 sg13g2_decap_8 FILLER_33_204 ();
 sg13g2_decap_8 FILLER_33_211 ();
 sg13g2_decap_4 FILLER_33_218 ();
 sg13g2_decap_8 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_257 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_268 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_decap_4 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_300 ();
 sg13g2_decap_8 FILLER_33_307 ();
 sg13g2_decap_8 FILLER_33_314 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_4 FILLER_33_343 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_153 ();
 sg13g2_decap_4 FILLER_34_160 ();
 sg13g2_fill_1 FILLER_34_168 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_fill_1 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_234 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_247 ();
 sg13g2_fill_1 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_254 ();
 sg13g2_decap_4 FILLER_34_282 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_decap_8 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_300 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_fill_1 FILLER_34_326 ();
 sg13g2_fill_2 FILLER_34_359 ();
 sg13g2_fill_2 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_fill_2 FILLER_35_120 ();
 sg13g2_decap_4 FILLER_35_132 ();
 sg13g2_fill_1 FILLER_35_136 ();
 sg13g2_decap_8 FILLER_35_142 ();
 sg13g2_fill_2 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_228 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_fill_2 FILLER_35_312 ();
 sg13g2_fill_1 FILLER_35_314 ();
 sg13g2_fill_2 FILLER_35_320 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_decap_4 FILLER_36_168 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_fill_2 FILLER_36_190 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_204 ();
 sg13g2_fill_1 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_249 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_4 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_4 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_102 ();
 sg13g2_fill_2 FILLER_37_150 ();
 sg13g2_decap_8 FILLER_37_157 ();
 sg13g2_decap_8 FILLER_37_164 ();
 sg13g2_decap_8 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_178 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_decap_8 FILLER_37_200 ();
 sg13g2_decap_8 FILLER_37_207 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_decap_4 FILLER_37_221 ();
 sg13g2_fill_1 FILLER_37_225 ();
 sg13g2_fill_2 FILLER_37_252 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_decap_4 FILLER_37_280 ();
 sg13g2_fill_1 FILLER_37_284 ();
 sg13g2_decap_4 FILLER_37_342 ();
 sg13g2_decap_8 FILLER_37_356 ();
 sg13g2_decap_8 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_370 ();
 sg13g2_fill_2 FILLER_37_382 ();
 sg13g2_fill_1 FILLER_37_384 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_fill_1 FILLER_38_112 ();
 sg13g2_fill_2 FILLER_38_118 ();
 sg13g2_fill_1 FILLER_38_120 ();
 sg13g2_fill_2 FILLER_38_131 ();
 sg13g2_fill_1 FILLER_38_138 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_150 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_4 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_4 FILLER_38_301 ();
 sg13g2_fill_2 FILLER_38_305 ();
 sg13g2_decap_4 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_fill_1 FILLER_38_345 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_2 FILLER_38_365 ();
 sg13g2_fill_1 FILLER_38_372 ();
 sg13g2_decap_4 FILLER_38_378 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_fill_1 FILLER_39_105 ();
 sg13g2_fill_2 FILLER_39_132 ();
 sg13g2_fill_2 FILLER_39_184 ();
 sg13g2_fill_1 FILLER_39_186 ();
 sg13g2_decap_4 FILLER_39_249 ();
 sg13g2_fill_2 FILLER_39_263 ();
 sg13g2_fill_1 FILLER_39_265 ();
 sg13g2_decap_8 FILLER_39_292 ();
 sg13g2_fill_1 FILLER_39_299 ();
 sg13g2_decap_4 FILLER_39_304 ();
 sg13g2_fill_2 FILLER_39_308 ();
 sg13g2_fill_1 FILLER_39_327 ();
 sg13g2_fill_1 FILLER_39_349 ();
 sg13g2_fill_1 FILLER_39_362 ();
 sg13g2_decap_8 FILLER_39_389 ();
 sg13g2_decap_8 FILLER_39_396 ();
 sg13g2_decap_4 FILLER_39_403 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_4 FILLER_40_91 ();
 sg13g2_fill_2 FILLER_40_95 ();
 sg13g2_fill_2 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_169 ();
 sg13g2_decap_4 FILLER_40_176 ();
 sg13g2_fill_2 FILLER_40_200 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_fill_2 FILLER_40_217 ();
 sg13g2_fill_1 FILLER_40_219 ();
 sg13g2_decap_4 FILLER_40_289 ();
 sg13g2_fill_2 FILLER_40_293 ();
 sg13g2_fill_2 FILLER_40_309 ();
 sg13g2_fill_2 FILLER_40_342 ();
 sg13g2_fill_1 FILLER_40_344 ();
 sg13g2_decap_4 FILLER_40_381 ();
 sg13g2_decap_8 FILLER_40_400 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_fill_1 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_132 ();
 sg13g2_decap_4 FILLER_41_139 ();
 sg13g2_decap_4 FILLER_41_149 ();
 sg13g2_fill_2 FILLER_41_159 ();
 sg13g2_decap_8 FILLER_41_165 ();
 sg13g2_decap_8 FILLER_41_172 ();
 sg13g2_fill_1 FILLER_41_179 ();
 sg13g2_decap_4 FILLER_41_185 ();
 sg13g2_decap_8 FILLER_41_194 ();
 sg13g2_fill_1 FILLER_41_201 ();
 sg13g2_decap_8 FILLER_41_208 ();
 sg13g2_decap_8 FILLER_41_215 ();
 sg13g2_decap_8 FILLER_41_222 ();
 sg13g2_decap_4 FILLER_41_256 ();
 sg13g2_decap_8 FILLER_41_278 ();
 sg13g2_fill_2 FILLER_41_285 ();
 sg13g2_decap_8 FILLER_41_297 ();
 sg13g2_decap_4 FILLER_41_304 ();
 sg13g2_fill_1 FILLER_41_308 ();
 sg13g2_fill_2 FILLER_41_320 ();
 sg13g2_fill_2 FILLER_41_332 ();
 sg13g2_decap_8 FILLER_41_339 ();
 sg13g2_fill_1 FILLER_41_346 ();
 sg13g2_decap_4 FILLER_41_357 ();
 sg13g2_fill_1 FILLER_41_361 ();
 sg13g2_fill_2 FILLER_41_372 ();
 sg13g2_fill_1 FILLER_41_374 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_fill_2 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_108 ();
 sg13g2_fill_1 FILLER_42_110 ();
 sg13g2_decap_8 FILLER_42_123 ();
 sg13g2_decap_8 FILLER_42_130 ();
 sg13g2_fill_2 FILLER_42_137 ();
 sg13g2_fill_2 FILLER_42_147 ();
 sg13g2_decap_4 FILLER_42_155 ();
 sg13g2_decap_4 FILLER_42_163 ();
 sg13g2_fill_2 FILLER_42_167 ();
 sg13g2_decap_4 FILLER_42_181 ();
 sg13g2_fill_1 FILLER_42_185 ();
 sg13g2_decap_8 FILLER_42_219 ();
 sg13g2_decap_8 FILLER_42_226 ();
 sg13g2_fill_1 FILLER_42_233 ();
 sg13g2_decap_4 FILLER_42_260 ();
 sg13g2_fill_1 FILLER_42_264 ();
 sg13g2_fill_2 FILLER_42_279 ();
 sg13g2_decap_4 FILLER_42_307 ();
 sg13g2_fill_1 FILLER_42_311 ();
 sg13g2_decap_4 FILLER_42_335 ();
 sg13g2_fill_1 FILLER_42_339 ();
 sg13g2_fill_1 FILLER_42_349 ();
 sg13g2_fill_2 FILLER_42_376 ();
 sg13g2_fill_1 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_fill_2 FILLER_43_110 ();
 sg13g2_decap_8 FILLER_43_118 ();
 sg13g2_decap_4 FILLER_43_125 ();
 sg13g2_fill_2 FILLER_43_129 ();
 sg13g2_fill_2 FILLER_43_161 ();
 sg13g2_fill_1 FILLER_43_163 ();
 sg13g2_decap_8 FILLER_43_233 ();
 sg13g2_decap_4 FILLER_43_240 ();
 sg13g2_fill_1 FILLER_43_252 ();
 sg13g2_decap_4 FILLER_43_275 ();
 sg13g2_fill_2 FILLER_43_279 ();
 sg13g2_fill_1 FILLER_43_315 ();
 sg13g2_fill_2 FILLER_43_342 ();
 sg13g2_fill_1 FILLER_43_344 ();
 sg13g2_fill_2 FILLER_43_376 ();
 sg13g2_fill_1 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_4 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_121 ();
 sg13g2_decap_8 FILLER_44_128 ();
 sg13g2_fill_2 FILLER_44_135 ();
 sg13g2_fill_1 FILLER_44_137 ();
 sg13g2_fill_2 FILLER_44_242 ();
 sg13g2_fill_2 FILLER_44_250 ();
 sg13g2_fill_1 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_285 ();
 sg13g2_fill_2 FILLER_44_292 ();
 sg13g2_fill_1 FILLER_44_294 ();
 sg13g2_fill_2 FILLER_44_303 ();
 sg13g2_decap_8 FILLER_44_339 ();
 sg13g2_decap_4 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_370 ();
 sg13g2_decap_4 FILLER_44_377 ();
 sg13g2_fill_2 FILLER_44_387 ();
 sg13g2_fill_1 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_400 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_132 ();
 sg13g2_fill_2 FILLER_45_139 ();
 sg13g2_fill_1 FILLER_45_141 ();
 sg13g2_fill_2 FILLER_45_148 ();
 sg13g2_fill_1 FILLER_45_155 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_fill_2 FILLER_45_203 ();
 sg13g2_fill_1 FILLER_45_205 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_decap_4 FILLER_45_306 ();
 sg13g2_decap_8 FILLER_45_316 ();
 sg13g2_decap_8 FILLER_45_323 ();
 sg13g2_decap_8 FILLER_45_330 ();
 sg13g2_decap_8 FILLER_45_337 ();
 sg13g2_decap_8 FILLER_45_344 ();
 sg13g2_decap_4 FILLER_45_351 ();
 sg13g2_fill_2 FILLER_45_355 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_4 FILLER_46_131 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_fill_2 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_fill_1 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_172 ();
 sg13g2_decap_8 FILLER_46_179 ();
 sg13g2_decap_8 FILLER_46_186 ();
 sg13g2_decap_8 FILLER_46_193 ();
 sg13g2_decap_8 FILLER_46_200 ();
 sg13g2_decap_8 FILLER_46_207 ();
 sg13g2_decap_8 FILLER_46_214 ();
 sg13g2_decap_8 FILLER_46_221 ();
 sg13g2_decap_4 FILLER_46_228 ();
 sg13g2_fill_2 FILLER_46_232 ();
 sg13g2_fill_2 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_261 ();
 sg13g2_decap_8 FILLER_46_268 ();
 sg13g2_fill_1 FILLER_46_275 ();
 sg13g2_decap_8 FILLER_46_286 ();
 sg13g2_decap_4 FILLER_46_293 ();
 sg13g2_fill_1 FILLER_46_297 ();
 sg13g2_fill_1 FILLER_46_313 ();
 sg13g2_decap_4 FILLER_46_328 ();
 sg13g2_fill_2 FILLER_46_332 ();
 sg13g2_decap_8 FILLER_46_342 ();
 sg13g2_decap_4 FILLER_46_349 ();
 sg13g2_fill_2 FILLER_46_353 ();
 sg13g2_decap_4 FILLER_46_367 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_98 ();
 sg13g2_fill_1 FILLER_47_100 ();
 sg13g2_fill_2 FILLER_47_120 ();
 sg13g2_fill_1 FILLER_47_122 ();
 sg13g2_decap_8 FILLER_47_149 ();
 sg13g2_decap_8 FILLER_47_160 ();
 sg13g2_decap_4 FILLER_47_182 ();
 sg13g2_fill_1 FILLER_47_186 ();
 sg13g2_decap_4 FILLER_47_213 ();
 sg13g2_fill_1 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_235 ();
 sg13g2_decap_8 FILLER_47_242 ();
 sg13g2_decap_8 FILLER_47_254 ();
 sg13g2_decap_4 FILLER_47_261 ();
 sg13g2_decap_8 FILLER_47_270 ();
 sg13g2_fill_2 FILLER_47_277 ();
 sg13g2_fill_1 FILLER_47_279 ();
 sg13g2_fill_1 FILLER_47_321 ();
 sg13g2_fill_1 FILLER_47_330 ();
 sg13g2_fill_2 FILLER_47_349 ();
 sg13g2_fill_1 FILLER_47_351 ();
 sg13g2_fill_2 FILLER_47_358 ();
 sg13g2_fill_2 FILLER_47_366 ();
 sg13g2_fill_1 FILLER_47_382 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_fill_2 FILLER_48_98 ();
 sg13g2_fill_2 FILLER_48_158 ();
 sg13g2_fill_1 FILLER_48_186 ();
 sg13g2_fill_2 FILLER_48_233 ();
 sg13g2_fill_2 FILLER_48_268 ();
 sg13g2_fill_1 FILLER_48_270 ();
 sg13g2_fill_2 FILLER_48_282 ();
 sg13g2_fill_1 FILLER_48_284 ();
 sg13g2_decap_8 FILLER_48_290 ();
 sg13g2_fill_1 FILLER_48_297 ();
 sg13g2_fill_1 FILLER_48_319 ();
 sg13g2_decap_4 FILLER_48_338 ();
 sg13g2_fill_1 FILLER_48_342 ();
 sg13g2_fill_1 FILLER_48_349 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_394 ();
 sg13g2_decap_8 FILLER_48_401 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_4 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_fill_1 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_118 ();
 sg13g2_fill_2 FILLER_49_162 ();
 sg13g2_fill_2 FILLER_49_196 ();
 sg13g2_fill_1 FILLER_49_211 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_fill_1 FILLER_49_230 ();
 sg13g2_fill_2 FILLER_49_248 ();
 sg13g2_fill_1 FILLER_49_250 ();
 sg13g2_fill_1 FILLER_49_266 ();
 sg13g2_decap_4 FILLER_49_285 ();
 sg13g2_decap_8 FILLER_49_303 ();
 sg13g2_fill_2 FILLER_49_310 ();
 sg13g2_fill_1 FILLER_49_331 ();
 sg13g2_fill_1 FILLER_49_336 ();
 sg13g2_fill_2 FILLER_49_343 ();
 sg13g2_fill_1 FILLER_49_345 ();
 sg13g2_fill_2 FILLER_49_379 ();
 sg13g2_decap_8 FILLER_49_386 ();
 sg13g2_decap_8 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_400 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_4 FILLER_50_91 ();
 sg13g2_fill_1 FILLER_50_95 ();
 sg13g2_fill_1 FILLER_50_104 ();
 sg13g2_decap_8 FILLER_50_117 ();
 sg13g2_decap_8 FILLER_50_124 ();
 sg13g2_fill_2 FILLER_50_131 ();
 sg13g2_fill_1 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_141 ();
 sg13g2_decap_8 FILLER_50_148 ();
 sg13g2_fill_2 FILLER_50_170 ();
 sg13g2_fill_2 FILLER_50_180 ();
 sg13g2_decap_8 FILLER_50_235 ();
 sg13g2_decap_8 FILLER_50_242 ();
 sg13g2_decap_4 FILLER_50_249 ();
 sg13g2_decap_8 FILLER_50_263 ();
 sg13g2_decap_4 FILLER_50_270 ();
 sg13g2_fill_2 FILLER_50_274 ();
 sg13g2_fill_2 FILLER_50_311 ();
 sg13g2_fill_1 FILLER_50_313 ();
 sg13g2_fill_2 FILLER_50_323 ();
 sg13g2_fill_1 FILLER_50_325 ();
 sg13g2_fill_2 FILLER_50_344 ();
 sg13g2_fill_1 FILLER_50_362 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_fill_2 FILLER_51_128 ();
 sg13g2_fill_1 FILLER_51_130 ();
 sg13g2_decap_8 FILLER_51_144 ();
 sg13g2_decap_4 FILLER_51_151 ();
 sg13g2_decap_4 FILLER_51_161 ();
 sg13g2_fill_2 FILLER_51_165 ();
 sg13g2_decap_8 FILLER_51_182 ();
 sg13g2_decap_8 FILLER_51_189 ();
 sg13g2_fill_1 FILLER_51_196 ();
 sg13g2_decap_8 FILLER_51_202 ();
 sg13g2_decap_8 FILLER_51_213 ();
 sg13g2_fill_2 FILLER_51_220 ();
 sg13g2_decap_8 FILLER_51_239 ();
 sg13g2_decap_4 FILLER_51_246 ();
 sg13g2_fill_1 FILLER_51_250 ();
 sg13g2_decap_8 FILLER_51_271 ();
 sg13g2_decap_4 FILLER_51_278 ();
 sg13g2_fill_2 FILLER_51_297 ();
 sg13g2_fill_2 FILLER_51_303 ();
 sg13g2_decap_8 FILLER_51_322 ();
 sg13g2_decap_4 FILLER_51_329 ();
 sg13g2_fill_2 FILLER_51_339 ();
 sg13g2_decap_4 FILLER_51_345 ();
 sg13g2_decap_8 FILLER_51_359 ();
 sg13g2_decap_4 FILLER_51_366 ();
 sg13g2_fill_2 FILLER_51_370 ();
 sg13g2_fill_2 FILLER_51_380 ();
 sg13g2_fill_1 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_4 FILLER_52_91 ();
 sg13g2_fill_1 FILLER_52_95 ();
 sg13g2_fill_2 FILLER_52_153 ();
 sg13g2_fill_1 FILLER_52_155 ();
 sg13g2_decap_8 FILLER_52_189 ();
 sg13g2_fill_1 FILLER_52_196 ();
 sg13g2_fill_1 FILLER_52_205 ();
 sg13g2_decap_8 FILLER_52_212 ();
 sg13g2_fill_2 FILLER_52_219 ();
 sg13g2_decap_4 FILLER_52_238 ();
 sg13g2_fill_2 FILLER_52_242 ();
 sg13g2_fill_1 FILLER_52_247 ();
 sg13g2_fill_1 FILLER_52_257 ();
 sg13g2_fill_2 FILLER_52_268 ();
 sg13g2_fill_1 FILLER_52_270 ();
 sg13g2_fill_2 FILLER_52_287 ();
 sg13g2_fill_1 FILLER_52_289 ();
 sg13g2_fill_2 FILLER_52_298 ();
 sg13g2_fill_1 FILLER_52_300 ();
 sg13g2_fill_1 FILLER_52_332 ();
 sg13g2_fill_1 FILLER_52_341 ();
 sg13g2_fill_2 FILLER_52_350 ();
 sg13g2_fill_2 FILLER_52_379 ();
 sg13g2_fill_1 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_400 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_fill_2 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_124 ();
 sg13g2_fill_1 FILLER_53_131 ();
 sg13g2_decap_4 FILLER_53_148 ();
 sg13g2_fill_1 FILLER_53_165 ();
 sg13g2_fill_2 FILLER_53_178 ();
 sg13g2_fill_2 FILLER_53_185 ();
 sg13g2_fill_2 FILLER_53_218 ();
 sg13g2_fill_1 FILLER_53_220 ();
 sg13g2_fill_2 FILLER_53_226 ();
 sg13g2_fill_1 FILLER_53_233 ();
 sg13g2_fill_2 FILLER_53_257 ();
 sg13g2_fill_2 FILLER_53_265 ();
 sg13g2_fill_1 FILLER_53_267 ();
 sg13g2_fill_2 FILLER_53_346 ();
 sg13g2_fill_1 FILLER_53_348 ();
 sg13g2_fill_2 FILLER_53_380 ();
 sg13g2_fill_1 FILLER_53_382 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_4 FILLER_54_98 ();
 sg13g2_fill_2 FILLER_54_102 ();
 sg13g2_fill_2 FILLER_54_130 ();
 sg13g2_fill_2 FILLER_54_163 ();
 sg13g2_fill_1 FILLER_54_165 ();
 sg13g2_fill_2 FILLER_54_200 ();
 sg13g2_fill_1 FILLER_54_202 ();
 sg13g2_decap_8 FILLER_54_211 ();
 sg13g2_fill_2 FILLER_54_218 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_fill_2 FILLER_54_243 ();
 sg13g2_decap_8 FILLER_54_253 ();
 sg13g2_fill_2 FILLER_54_260 ();
 sg13g2_fill_1 FILLER_54_262 ();
 sg13g2_decap_8 FILLER_54_274 ();
 sg13g2_decap_4 FILLER_54_281 ();
 sg13g2_fill_2 FILLER_54_296 ();
 sg13g2_decap_8 FILLER_54_321 ();
 sg13g2_decap_4 FILLER_54_328 ();
 sg13g2_fill_1 FILLER_54_332 ();
 sg13g2_fill_1 FILLER_54_385 ();
 sg13g2_decap_8 FILLER_54_401 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_4 FILLER_55_91 ();
 sg13g2_fill_1 FILLER_55_95 ();
 sg13g2_fill_1 FILLER_55_113 ();
 sg13g2_fill_2 FILLER_55_119 ();
 sg13g2_fill_2 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_221 ();
 sg13g2_decap_8 FILLER_55_228 ();
 sg13g2_decap_4 FILLER_55_235 ();
 sg13g2_fill_1 FILLER_55_239 ();
 sg13g2_fill_2 FILLER_55_248 ();
 sg13g2_fill_1 FILLER_55_250 ();
 sg13g2_decap_4 FILLER_55_264 ();
 sg13g2_fill_2 FILLER_55_268 ();
 sg13g2_decap_8 FILLER_55_275 ();
 sg13g2_decap_4 FILLER_55_282 ();
 sg13g2_decap_8 FILLER_55_291 ();
 sg13g2_fill_2 FILLER_55_304 ();
 sg13g2_fill_1 FILLER_55_306 ();
 sg13g2_decap_8 FILLER_55_311 ();
 sg13g2_decap_8 FILLER_55_318 ();
 sg13g2_decap_8 FILLER_55_325 ();
 sg13g2_fill_2 FILLER_55_332 ();
 sg13g2_fill_2 FILLER_55_339 ();
 sg13g2_fill_1 FILLER_55_341 ();
 sg13g2_decap_8 FILLER_55_347 ();
 sg13g2_fill_1 FILLER_55_354 ();
 sg13g2_decap_8 FILLER_55_359 ();
 sg13g2_fill_2 FILLER_55_366 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_4 FILLER_56_98 ();
 sg13g2_fill_1 FILLER_56_102 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_fill_1 FILLER_56_140 ();
 sg13g2_fill_2 FILLER_56_162 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_fill_1 FILLER_56_175 ();
 sg13g2_fill_2 FILLER_56_180 ();
 sg13g2_fill_1 FILLER_56_182 ();
 sg13g2_decap_8 FILLER_56_193 ();
 sg13g2_decap_8 FILLER_56_200 ();
 sg13g2_decap_8 FILLER_56_207 ();
 sg13g2_decap_8 FILLER_56_232 ();
 sg13g2_fill_1 FILLER_56_239 ();
 sg13g2_decap_8 FILLER_56_243 ();
 sg13g2_decap_4 FILLER_56_250 ();
 sg13g2_fill_1 FILLER_56_254 ();
 sg13g2_decap_4 FILLER_56_264 ();
 sg13g2_fill_1 FILLER_56_285 ();
 sg13g2_decap_8 FILLER_56_294 ();
 sg13g2_decap_4 FILLER_56_301 ();
 sg13g2_fill_1 FILLER_56_305 ();
 sg13g2_decap_4 FILLER_56_311 ();
 sg13g2_decap_8 FILLER_56_320 ();
 sg13g2_decap_8 FILLER_56_327 ();
 sg13g2_fill_2 FILLER_56_334 ();
 sg13g2_fill_1 FILLER_56_336 ();
 sg13g2_decap_4 FILLER_56_352 ();
 sg13g2_decap_8 FILLER_56_359 ();
 sg13g2_decap_8 FILLER_56_366 ();
 sg13g2_fill_2 FILLER_56_373 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_4 FILLER_57_105 ();
 sg13g2_fill_1 FILLER_57_109 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_fill_2 FILLER_57_140 ();
 sg13g2_fill_1 FILLER_57_142 ();
 sg13g2_decap_8 FILLER_57_148 ();
 sg13g2_decap_8 FILLER_57_155 ();
 sg13g2_fill_1 FILLER_57_162 ();
 sg13g2_fill_2 FILLER_57_169 ();
 sg13g2_fill_1 FILLER_57_171 ();
 sg13g2_decap_4 FILLER_57_181 ();
 sg13g2_decap_4 FILLER_57_199 ();
 sg13g2_fill_2 FILLER_57_208 ();
 sg13g2_fill_1 FILLER_57_210 ();
 sg13g2_fill_2 FILLER_57_246 ();
 sg13g2_fill_1 FILLER_57_248 ();
 sg13g2_fill_2 FILLER_57_260 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_fill_2 FILLER_57_281 ();
 sg13g2_fill_2 FILLER_57_297 ();
 sg13g2_fill_1 FILLER_57_299 ();
 sg13g2_fill_1 FILLER_57_310 ();
 sg13g2_decap_8 FILLER_57_370 ();
 sg13g2_decap_8 FILLER_57_377 ();
 sg13g2_fill_1 FILLER_57_384 ();
 sg13g2_fill_2 FILLER_57_389 ();
 sg13g2_decap_8 FILLER_57_401 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_4 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_135 ();
 sg13g2_decap_8 FILLER_58_142 ();
 sg13g2_decap_8 FILLER_58_149 ();
 sg13g2_decap_8 FILLER_58_160 ();
 sg13g2_fill_2 FILLER_58_167 ();
 sg13g2_fill_1 FILLER_58_169 ();
 sg13g2_decap_4 FILLER_58_240 ();
 sg13g2_fill_2 FILLER_58_249 ();
 sg13g2_fill_1 FILLER_58_251 ();
 sg13g2_fill_2 FILLER_58_299 ();
 sg13g2_fill_1 FILLER_58_301 ();
 sg13g2_fill_1 FILLER_58_337 ();
 sg13g2_decap_8 FILLER_58_380 ();
 sg13g2_decap_8 FILLER_58_387 ();
 sg13g2_decap_8 FILLER_58_394 ();
 sg13g2_decap_8 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_fill_1 FILLER_59_98 ();
 sg13g2_fill_1 FILLER_59_135 ();
 sg13g2_fill_2 FILLER_59_144 ();
 sg13g2_fill_2 FILLER_59_164 ();
 sg13g2_fill_1 FILLER_59_166 ();
 sg13g2_fill_2 FILLER_59_223 ();
 sg13g2_fill_1 FILLER_59_225 ();
 sg13g2_fill_2 FILLER_59_306 ();
 sg13g2_fill_1 FILLER_59_308 ();
 sg13g2_decap_4 FILLER_59_326 ();
 sg13g2_fill_2 FILLER_59_330 ();
 sg13g2_decap_4 FILLER_59_337 ();
 sg13g2_fill_2 FILLER_59_346 ();
 sg13g2_decap_4 FILLER_59_403 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_fill_1 FILLER_60_113 ();
 sg13g2_fill_2 FILLER_60_176 ();
 sg13g2_fill_1 FILLER_60_178 ();
 sg13g2_fill_1 FILLER_60_183 ();
 sg13g2_decap_4 FILLER_60_203 ();
 sg13g2_decap_8 FILLER_60_223 ();
 sg13g2_decap_8 FILLER_60_230 ();
 sg13g2_decap_8 FILLER_60_237 ();
 sg13g2_fill_2 FILLER_60_244 ();
 sg13g2_fill_1 FILLER_60_246 ();
 sg13g2_fill_2 FILLER_60_299 ();
 sg13g2_fill_1 FILLER_60_301 ();
 sg13g2_decap_8 FILLER_60_322 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_decap_8 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_343 ();
 sg13g2_decap_8 FILLER_60_350 ();
 sg13g2_fill_1 FILLER_60_357 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_fill_2 FILLER_61_91 ();
 sg13g2_fill_2 FILLER_61_134 ();
 sg13g2_fill_2 FILLER_61_141 ();
 sg13g2_decap_8 FILLER_61_174 ();
 sg13g2_decap_8 FILLER_61_181 ();
 sg13g2_decap_8 FILLER_61_188 ();
 sg13g2_decap_8 FILLER_61_195 ();
 sg13g2_decap_8 FILLER_61_202 ();
 sg13g2_decap_8 FILLER_61_209 ();
 sg13g2_decap_8 FILLER_61_216 ();
 sg13g2_decap_8 FILLER_61_223 ();
 sg13g2_decap_8 FILLER_61_230 ();
 sg13g2_fill_2 FILLER_61_237 ();
 sg13g2_decap_8 FILLER_61_243 ();
 sg13g2_decap_8 FILLER_61_250 ();
 sg13g2_fill_1 FILLER_61_284 ();
 sg13g2_fill_1 FILLER_61_290 ();
 sg13g2_decap_4 FILLER_61_295 ();
 sg13g2_fill_2 FILLER_61_299 ();
 sg13g2_decap_8 FILLER_61_327 ();
 sg13g2_decap_4 FILLER_61_334 ();
 sg13g2_decap_8 FILLER_61_348 ();
 sg13g2_decap_8 FILLER_61_355 ();
 sg13g2_decap_4 FILLER_61_362 ();
 sg13g2_fill_1 FILLER_61_374 ();
 sg13g2_fill_2 FILLER_61_387 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_4 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_136 ();
 sg13g2_fill_2 FILLER_62_143 ();
 sg13g2_fill_1 FILLER_62_145 ();
 sg13g2_fill_1 FILLER_62_152 ();
 sg13g2_fill_2 FILLER_62_179 ();
 sg13g2_fill_2 FILLER_62_194 ();
 sg13g2_fill_1 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_202 ();
 sg13g2_decap_8 FILLER_62_209 ();
 sg13g2_decap_4 FILLER_62_216 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_decap_4 FILLER_62_266 ();
 sg13g2_fill_2 FILLER_62_270 ();
 sg13g2_decap_4 FILLER_62_297 ();
 sg13g2_fill_2 FILLER_62_310 ();
 sg13g2_fill_1 FILLER_62_312 ();
 sg13g2_fill_2 FILLER_62_324 ();
 sg13g2_fill_1 FILLER_62_326 ();
 sg13g2_fill_2 FILLER_62_373 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_4 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_113 ();
 sg13g2_fill_1 FILLER_63_120 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_4 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_142 ();
 sg13g2_decap_4 FILLER_63_149 ();
 sg13g2_decap_8 FILLER_63_158 ();
 sg13g2_decap_8 FILLER_63_165 ();
 sg13g2_decap_8 FILLER_63_172 ();
 sg13g2_decap_8 FILLER_63_179 ();
 sg13g2_fill_2 FILLER_63_212 ();
 sg13g2_fill_1 FILLER_63_245 ();
 sg13g2_fill_1 FILLER_63_255 ();
 sg13g2_fill_2 FILLER_63_279 ();
 sg13g2_fill_1 FILLER_63_281 ();
 sg13g2_fill_2 FILLER_63_296 ();
 sg13g2_fill_1 FILLER_63_298 ();
 sg13g2_decap_4 FILLER_63_304 ();
 sg13g2_fill_1 FILLER_63_308 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_4 FILLER_64_126 ();
 sg13g2_fill_2 FILLER_64_130 ();
 sg13g2_fill_2 FILLER_64_168 ();
 sg13g2_fill_2 FILLER_64_178 ();
 sg13g2_fill_1 FILLER_64_180 ();
 sg13g2_fill_2 FILLER_64_217 ();
 sg13g2_fill_1 FILLER_64_219 ();
 sg13g2_fill_2 FILLER_64_269 ();
 sg13g2_fill_2 FILLER_64_291 ();
 sg13g2_fill_2 FILLER_64_297 ();
 sg13g2_fill_2 FILLER_64_304 ();
 sg13g2_fill_1 FILLER_64_306 ();
 sg13g2_decap_8 FILLER_64_315 ();
 sg13g2_fill_2 FILLER_64_322 ();
 sg13g2_fill_1 FILLER_64_324 ();
 sg13g2_fill_2 FILLER_64_372 ();
 sg13g2_fill_1 FILLER_64_374 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_fill_1 FILLER_65_119 ();
 sg13g2_fill_1 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_243 ();
 sg13g2_fill_1 FILLER_65_286 ();
 sg13g2_decap_8 FILLER_65_306 ();
 sg13g2_fill_1 FILLER_65_313 ();
 sg13g2_decap_8 FILLER_65_322 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_fill_2 FILLER_65_336 ();
 sg13g2_fill_1 FILLER_65_338 ();
 sg13g2_fill_2 FILLER_65_347 ();
 sg13g2_fill_1 FILLER_65_362 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_4 FILLER_65_378 ();
 sg13g2_fill_2 FILLER_65_382 ();
 sg13g2_decap_8 FILLER_65_394 ();
 sg13g2_decap_8 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_4 FILLER_66_126 ();
 sg13g2_decap_4 FILLER_66_169 ();
 sg13g2_fill_1 FILLER_66_173 ();
 sg13g2_decap_4 FILLER_66_179 ();
 sg13g2_fill_2 FILLER_66_198 ();
 sg13g2_fill_2 FILLER_66_216 ();
 sg13g2_fill_1 FILLER_66_218 ();
 sg13g2_fill_2 FILLER_66_256 ();
 sg13g2_fill_1 FILLER_66_288 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_decap_8 FILLER_66_327 ();
 sg13g2_decap_8 FILLER_66_334 ();
 sg13g2_fill_1 FILLER_66_382 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_4 FILLER_67_133 ();
 sg13g2_fill_1 FILLER_67_137 ();
 sg13g2_decap_8 FILLER_67_142 ();
 sg13g2_fill_2 FILLER_67_149 ();
 sg13g2_fill_1 FILLER_67_151 ();
 sg13g2_decap_8 FILLER_67_157 ();
 sg13g2_decap_8 FILLER_67_164 ();
 sg13g2_decap_4 FILLER_67_171 ();
 sg13g2_fill_2 FILLER_67_175 ();
 sg13g2_decap_4 FILLER_67_208 ();
 sg13g2_fill_2 FILLER_67_212 ();
 sg13g2_decap_4 FILLER_67_254 ();
 sg13g2_fill_2 FILLER_67_306 ();
 sg13g2_fill_1 FILLER_67_308 ();
 sg13g2_fill_2 FILLER_67_319 ();
 sg13g2_fill_1 FILLER_67_321 ();
 sg13g2_fill_2 FILLER_67_331 ();
 sg13g2_decap_8 FILLER_67_402 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_fill_1 FILLER_68_147 ();
 sg13g2_fill_2 FILLER_68_156 ();
 sg13g2_decap_8 FILLER_68_163 ();
 sg13g2_fill_1 FILLER_68_170 ();
 sg13g2_decap_8 FILLER_68_176 ();
 sg13g2_decap_4 FILLER_68_183 ();
 sg13g2_fill_1 FILLER_68_187 ();
 sg13g2_decap_8 FILLER_68_192 ();
 sg13g2_decap_8 FILLER_68_199 ();
 sg13g2_decap_8 FILLER_68_206 ();
 sg13g2_decap_8 FILLER_68_213 ();
 sg13g2_fill_1 FILLER_68_220 ();
 sg13g2_fill_2 FILLER_68_319 ();
 sg13g2_fill_2 FILLER_68_347 ();
 sg13g2_fill_1 FILLER_68_349 ();
 sg13g2_decap_8 FILLER_68_365 ();
 sg13g2_decap_4 FILLER_68_372 ();
 sg13g2_decap_8 FILLER_68_386 ();
 sg13g2_decap_8 FILLER_68_393 ();
 sg13g2_decap_8 FILLER_68_400 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_fill_2 FILLER_69_133 ();
 sg13g2_fill_1 FILLER_69_135 ();
 sg13g2_fill_1 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_203 ();
 sg13g2_fill_2 FILLER_69_210 ();
 sg13g2_decap_4 FILLER_69_217 ();
 sg13g2_decap_8 FILLER_69_226 ();
 sg13g2_fill_1 FILLER_69_233 ();
 sg13g2_decap_4 FILLER_69_250 ();
 sg13g2_fill_1 FILLER_69_254 ();
 sg13g2_fill_1 FILLER_69_292 ();
 sg13g2_decap_8 FILLER_69_298 ();
 sg13g2_decap_8 FILLER_69_320 ();
 sg13g2_decap_8 FILLER_69_327 ();
 sg13g2_fill_1 FILLER_69_334 ();
 sg13g2_fill_2 FILLER_69_340 ();
 sg13g2_fill_1 FILLER_69_342 ();
 sg13g2_decap_8 FILLER_69_354 ();
 sg13g2_decap_8 FILLER_69_361 ();
 sg13g2_decap_8 FILLER_69_368 ();
 sg13g2_decap_4 FILLER_69_380 ();
 sg13g2_decap_8 FILLER_69_388 ();
 sg13g2_decap_8 FILLER_69_395 ();
 sg13g2_decap_8 FILLER_69_402 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_4 FILLER_70_126 ();
 sg13g2_fill_2 FILLER_70_130 ();
 sg13g2_fill_1 FILLER_70_205 ();
 sg13g2_decap_4 FILLER_70_216 ();
 sg13g2_fill_1 FILLER_70_294 ();
 sg13g2_fill_2 FILLER_70_344 ();
 sg13g2_fill_1 FILLER_70_346 ();
 sg13g2_fill_1 FILLER_70_353 ();
 sg13g2_decap_8 FILLER_70_360 ();
 sg13g2_fill_1 FILLER_70_367 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_fill_2 FILLER_71_140 ();
 sg13g2_fill_1 FILLER_71_142 ();
 sg13g2_fill_2 FILLER_71_174 ();
 sg13g2_fill_1 FILLER_71_176 ();
 sg13g2_decap_4 FILLER_71_188 ();
 sg13g2_fill_1 FILLER_71_218 ();
 sg13g2_fill_1 FILLER_71_224 ();
 sg13g2_fill_1 FILLER_71_269 ();
 sg13g2_decap_4 FILLER_71_348 ();
 sg13g2_fill_1 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_fill_1 FILLER_72_147 ();
 sg13g2_fill_1 FILLER_72_157 ();
 sg13g2_decap_8 FILLER_72_163 ();
 sg13g2_decap_8 FILLER_72_170 ();
 sg13g2_decap_8 FILLER_72_177 ();
 sg13g2_fill_2 FILLER_72_184 ();
 sg13g2_fill_1 FILLER_72_186 ();
 sg13g2_fill_1 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_223 ();
 sg13g2_decap_8 FILLER_72_230 ();
 sg13g2_decap_8 FILLER_72_237 ();
 sg13g2_fill_1 FILLER_72_244 ();
 sg13g2_fill_1 FILLER_72_253 ();
 sg13g2_decap_4 FILLER_72_302 ();
 sg13g2_fill_2 FILLER_72_336 ();
 sg13g2_fill_1 FILLER_72_338 ();
 sg13g2_fill_1 FILLER_72_391 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_4 FILLER_73_168 ();
 sg13g2_fill_2 FILLER_73_172 ();
 sg13g2_decap_8 FILLER_73_188 ();
 sg13g2_fill_1 FILLER_73_195 ();
 sg13g2_fill_2 FILLER_73_216 ();
 sg13g2_fill_2 FILLER_73_230 ();
 sg13g2_fill_1 FILLER_73_271 ();
 sg13g2_decap_8 FILLER_73_300 ();
 sg13g2_decap_8 FILLER_73_307 ();
 sg13g2_decap_8 FILLER_73_314 ();
 sg13g2_decap_8 FILLER_73_321 ();
 sg13g2_decap_8 FILLER_73_328 ();
 sg13g2_fill_1 FILLER_73_335 ();
 sg13g2_fill_1 FILLER_73_342 ();
 sg13g2_decap_8 FILLER_73_360 ();
 sg13g2_decap_4 FILLER_73_367 ();
 sg13g2_fill_1 FILLER_73_371 ();
 sg13g2_decap_8 FILLER_73_382 ();
 sg13g2_fill_2 FILLER_73_389 ();
 sg13g2_decap_8 FILLER_73_396 ();
 sg13g2_decap_4 FILLER_73_403 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_4 FILLER_74_161 ();
 sg13g2_fill_1 FILLER_74_165 ();
 sg13g2_decap_8 FILLER_74_192 ();
 sg13g2_decap_8 FILLER_74_199 ();
 sg13g2_decap_4 FILLER_74_206 ();
 sg13g2_fill_1 FILLER_74_210 ();
 sg13g2_fill_1 FILLER_74_220 ();
 sg13g2_fill_2 FILLER_74_247 ();
 sg13g2_fill_1 FILLER_74_254 ();
 sg13g2_fill_1 FILLER_74_264 ();
 sg13g2_fill_2 FILLER_74_274 ();
 sg13g2_fill_1 FILLER_74_281 ();
 sg13g2_decap_4 FILLER_74_314 ();
 sg13g2_fill_2 FILLER_74_323 ();
 sg13g2_fill_1 FILLER_74_334 ();
 sg13g2_decap_4 FILLER_74_340 ();
 sg13g2_fill_1 FILLER_74_357 ();
 sg13g2_decap_4 FILLER_74_368 ();
 sg13g2_fill_2 FILLER_74_372 ();
 sg13g2_fill_1 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_fill_1 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_181 ();
 sg13g2_decap_4 FILLER_75_188 ();
 sg13g2_fill_1 FILLER_75_192 ();
 sg13g2_decap_8 FILLER_75_208 ();
 sg13g2_decap_4 FILLER_75_215 ();
 sg13g2_fill_1 FILLER_75_219 ();
 sg13g2_fill_2 FILLER_75_260 ();
 sg13g2_fill_2 FILLER_75_282 ();
 sg13g2_decap_8 FILLER_75_346 ();
 sg13g2_fill_2 FILLER_75_353 ();
 sg13g2_fill_1 FILLER_75_355 ();
 sg13g2_fill_1 FILLER_75_365 ();
 sg13g2_fill_1 FILLER_75_378 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_4 FILLER_76_168 ();
 sg13g2_fill_1 FILLER_76_172 ();
 sg13g2_fill_1 FILLER_76_215 ();
 sg13g2_fill_2 FILLER_76_248 ();
 sg13g2_fill_1 FILLER_76_250 ();
 sg13g2_fill_2 FILLER_76_297 ();
 sg13g2_fill_2 FILLER_76_327 ();
 sg13g2_fill_1 FILLER_76_329 ();
 sg13g2_fill_2 FILLER_76_356 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_4 FILLER_77_168 ();
 sg13g2_fill_2 FILLER_77_172 ();
 sg13g2_fill_1 FILLER_77_247 ();
 sg13g2_fill_2 FILLER_77_305 ();
 sg13g2_fill_2 FILLER_77_346 ();
 sg13g2_decap_4 FILLER_77_357 ();
 sg13g2_fill_1 FILLER_77_361 ();
 sg13g2_fill_1 FILLER_77_370 ();
 sg13g2_fill_1 FILLER_77_386 ();
 sg13g2_decap_8 FILLER_77_400 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_4 FILLER_78_175 ();
 sg13g2_fill_1 FILLER_78_179 ();
 sg13g2_fill_1 FILLER_78_184 ();
 sg13g2_fill_2 FILLER_78_221 ();
 sg13g2_fill_1 FILLER_78_324 ();
 sg13g2_fill_2 FILLER_78_367 ();
 sg13g2_fill_1 FILLER_78_374 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_fill_2 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_207 ();
 sg13g2_decap_4 FILLER_79_214 ();
 sg13g2_fill_2 FILLER_79_244 ();
 sg13g2_fill_1 FILLER_79_246 ();
 sg13g2_decap_8 FILLER_79_321 ();
 sg13g2_decap_4 FILLER_79_328 ();
 sg13g2_decap_4 FILLER_79_384 ();
 sg13g2_fill_2 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_8 FILLER_80_233 ();
 sg13g2_fill_2 FILLER_80_240 ();
 sg13g2_fill_1 FILLER_80_242 ();
 sg13g2_fill_2 FILLER_80_251 ();
 sg13g2_fill_1 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_307 ();
 sg13g2_decap_8 FILLER_80_314 ();
 sg13g2_decap_8 FILLER_80_321 ();
 sg13g2_decap_8 FILLER_80_328 ();
 sg13g2_decap_8 FILLER_80_350 ();
 sg13g2_decap_8 FILLER_80_357 ();
 sg13g2_decap_8 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_371 ();
 sg13g2_decap_4 FILLER_80_378 ();
 sg13g2_fill_1 FILLER_80_382 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
endmodule

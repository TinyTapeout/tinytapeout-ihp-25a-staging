module tt_um_tiny_shader_mole99 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire clk_regs;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire hsync;
 wire next_frame;
 wire next_vertical;
 wire rst_n_sync;
 wire spi_miso;
 wire \tiny_shader_top_inst.capture ;
 wire \tiny_shader_top_inst.counter_h[0] ;
 wire \tiny_shader_top_inst.counter_h[10] ;
 wire \tiny_shader_top_inst.counter_h[1] ;
 wire \tiny_shader_top_inst.counter_h[2] ;
 wire \tiny_shader_top_inst.counter_h[3] ;
 wire \tiny_shader_top_inst.counter_h[4] ;
 wire \tiny_shader_top_inst.counter_h[5] ;
 wire \tiny_shader_top_inst.counter_h[6] ;
 wire \tiny_shader_top_inst.counter_h[7] ;
 wire \tiny_shader_top_inst.counter_h[8] ;
 wire \tiny_shader_top_inst.counter_h[9] ;
 wire \tiny_shader_top_inst.counter_v[0] ;
 wire \tiny_shader_top_inst.counter_v[10] ;
 wire \tiny_shader_top_inst.counter_v[1] ;
 wire \tiny_shader_top_inst.counter_v[2] ;
 wire \tiny_shader_top_inst.counter_v[3] ;
 wire \tiny_shader_top_inst.counter_v[4] ;
 wire \tiny_shader_top_inst.counter_v[5] ;
 wire \tiny_shader_top_inst.counter_v[6] ;
 wire \tiny_shader_top_inst.counter_v[7] ;
 wire \tiny_shader_top_inst.counter_v[8] ;
 wire \tiny_shader_top_inst.counter_v[9] ;
 wire \tiny_shader_top_inst.cur_time[0] ;
 wire \tiny_shader_top_inst.cur_time[1] ;
 wire \tiny_shader_top_inst.cur_time[2] ;
 wire \tiny_shader_top_inst.cur_time[3] ;
 wire \tiny_shader_top_inst.cur_time[4] ;
 wire \tiny_shader_top_inst.cur_time[5] ;
 wire \tiny_shader_top_inst.cur_time[6] ;
 wire \tiny_shader_top_inst.cur_time[7] ;
 wire \tiny_shader_top_inst.cur_time[8] ;
 wire \tiny_shader_top_inst.hsync ;
 wire \tiny_shader_top_inst.instr[0] ;
 wire \tiny_shader_top_inst.instr[1] ;
 wire \tiny_shader_top_inst.instr[2] ;
 wire \tiny_shader_top_inst.instr[3] ;
 wire \tiny_shader_top_inst.instr[4] ;
 wire \tiny_shader_top_inst.instr[5] ;
 wire \tiny_shader_top_inst.instr[6] ;
 wire \tiny_shader_top_inst.instr[7] ;
 wire \tiny_shader_top_inst.memory_instr[0] ;
 wire \tiny_shader_top_inst.memory_instr[1] ;
 wire \tiny_shader_top_inst.memory_instr[2] ;
 wire \tiny_shader_top_inst.memory_instr[3] ;
 wire \tiny_shader_top_inst.memory_instr[4] ;
 wire \tiny_shader_top_inst.memory_instr[5] ;
 wire \tiny_shader_top_inst.memory_instr[6] ;
 wire \tiny_shader_top_inst.memory_instr[7] ;
 wire \tiny_shader_top_inst.memory_load ;
 wire \tiny_shader_top_inst.next_frame ;
 wire \tiny_shader_top_inst.next_vertical ;
 wire \tiny_shader_top_inst.rgb_o[0] ;
 wire \tiny_shader_top_inst.rgb_o[1] ;
 wire \tiny_shader_top_inst.rgb_o[2] ;
 wire \tiny_shader_top_inst.rgb_o[3] ;
 wire \tiny_shader_top_inst.rgb_o[4] ;
 wire \tiny_shader_top_inst.rgb_o[5] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[0][0] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[0][1] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[0][2] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[0][3] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[0][4] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[0][5] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[1][0] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[1][1] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[1][2] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[1][3] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[1][4] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[1][5] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[2][0] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[2][1] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[2][2] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[2][3] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[2][4] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[2][5] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[3][0] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[3][1] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[3][2] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[3][3] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[3][4] ;
 wire \tiny_shader_top_inst.shader_execute_inst.regs[3][5] ;
 wire \tiny_shader_top_inst.shader_execute_inst.skip ;
 wire \tiny_shader_top_inst.shader_execute_inst.user_i[0] ;
 wire \tiny_shader_top_inst.shader_execute_inst.user_i[1] ;
 wire \tiny_shader_top_inst.shader_execute_inst.user_i[2] ;
 wire \tiny_shader_top_inst.shader_execute_inst.user_i[3] ;
 wire \tiny_shader_top_inst.shader_execute_inst.user_i[4] ;
 wire \tiny_shader_top_inst.shader_execute_inst.user_i[5] ;
 wire \tiny_shader_top_inst.shader_execute_inst.x_pos_i[0] ;
 wire \tiny_shader_top_inst.shader_execute_inst.x_pos_i[1] ;
 wire \tiny_shader_top_inst.shader_execute_inst.x_pos_i[2] ;
 wire \tiny_shader_top_inst.shader_execute_inst.x_pos_i[3] ;
 wire \tiny_shader_top_inst.shader_execute_inst.x_pos_i[4] ;
 wire \tiny_shader_top_inst.shader_execute_inst.x_pos_i[5] ;
 wire \tiny_shader_top_inst.shader_execute_inst.y_pos_i[0] ;
 wire \tiny_shader_top_inst.shader_execute_inst.y_pos_i[1] ;
 wire \tiny_shader_top_inst.shader_execute_inst.y_pos_i[2] ;
 wire \tiny_shader_top_inst.shader_execute_inst.y_pos_i[3] ;
 wire \tiny_shader_top_inst.shader_execute_inst.y_pos_i[4] ;
 wire \tiny_shader_top_inst.shader_execute_inst.y_pos_i[5] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[1][0] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[1][1] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[1][2] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[1][3] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[1][4] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[1][5] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[1][6] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[1][7] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[2][0] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[2][1] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[2][2] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[2][3] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[2][4] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[2][5] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[2][6] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[2][7] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[3][0] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[3][1] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[3][2] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[3][3] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[3][4] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[3][5] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[3][6] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[3][7] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[4][0] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[4][1] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[4][2] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[4][3] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[4][4] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[4][5] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[4][6] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[4][7] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[5][0] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[5][1] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[5][2] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[5][3] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[5][4] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[5][5] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[5][6] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[5][7] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[6][0] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[6][1] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[6][2] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[6][3] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[6][4] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[6][5] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[6][6] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[6][7] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[7][0] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[7][1] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[7][2] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[7][3] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[7][4] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[7][5] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[7][6] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[7][7] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[8][0] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[8][1] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[8][2] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[8][3] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[8][4] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[8][5] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[8][6] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[8][7] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[9][0] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[9][1] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[9][2] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[9][3] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[9][4] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[9][5] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[9][6] ;
 wire \tiny_shader_top_inst.shader_memory_inst.memory[9][7] ;
 wire \tiny_shader_top_inst.spi_receiver_inst.mode_sync ;
 wire \tiny_shader_top_inst.spi_receiver_inst.spi_cnt[0] ;
 wire \tiny_shader_top_inst.spi_receiver_inst.spi_cnt[1] ;
 wire \tiny_shader_top_inst.spi_receiver_inst.spi_cnt[2] ;
 wire \tiny_shader_top_inst.spi_receiver_inst.spi_cs_sync ;
 wire \tiny_shader_top_inst.spi_receiver_inst.spi_mosi_sync ;
 wire \tiny_shader_top_inst.spi_receiver_inst.spi_sclk_delayed ;
 wire \tiny_shader_top_inst.spi_receiver_inst.spi_sclk_sync ;
 wire \tiny_shader_top_inst.spi_receiver_inst.synchronizer_mode.pipe[0] ;
 wire \tiny_shader_top_inst.spi_receiver_inst.synchronizer_spi_cs.pipe[0] ;
 wire \tiny_shader_top_inst.spi_receiver_inst.synchronizer_spi_mosi.pipe[0] ;
 wire \tiny_shader_top_inst.spi_receiver_inst.synchronizer_spi_sclk.pipe[0] ;
 wire \tiny_shader_top_inst.time_dir ;
 wire \tiny_shader_top_inst.timing_ver.sync ;
 wire \tiny_shader_top_inst.vsync_o ;
 wire \tiny_shader_top_inst.x_subpos[0] ;
 wire \tiny_shader_top_inst.x_subpos[1] ;
 wire \tiny_shader_top_inst.x_subpos[2] ;
 wire \tiny_shader_top_inst.x_subpos[3] ;
 wire \tiny_shader_top_inst.y_subpos[0] ;
 wire \tiny_shader_top_inst.y_subpos[1] ;
 wire \tiny_shader_top_inst.y_subpos[2] ;
 wire \tiny_shader_top_inst.y_subpos[3] ;
 wire net9;
 wire net10;
 wire net21;
 wire net11;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net12;
 wire net13;
 wire net14;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_3_0__leaf_clk_regs;
 wire clknet_3_1__leaf_clk_regs;
 wire clknet_3_2__leaf_clk_regs;
 wire clknet_3_3__leaf_clk_regs;
 wire clknet_3_4__leaf_clk_regs;
 wire clknet_3_5__leaf_clk_regs;
 wire clknet_3_6__leaf_clk_regs;
 wire clknet_3_7__leaf_clk_regs;
 wire delaynet_0_clk;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;

 sg13g2_inv_1 _1062_ (.Y(_0427_),
    .A(\tiny_shader_top_inst.spi_receiver_inst.spi_cnt[0] ));
 sg13g2_inv_1 _1063_ (.Y(_0428_),
    .A(net316));
 sg13g2_inv_1 _1064_ (.Y(_0429_),
    .A(net435));
 sg13g2_inv_1 _1065_ (.Y(_0430_),
    .A(\tiny_shader_top_inst.counter_h[10] ));
 sg13g2_inv_1 _1066_ (.Y(_0431_),
    .A(net318));
 sg13g2_inv_4 _1067_ (.A(net455),
    .Y(_0432_));
 sg13g2_inv_1 _1068_ (.Y(_0433_),
    .A(net451));
 sg13g2_inv_1 _1069_ (.Y(_0434_),
    .A(\tiny_shader_top_inst.counter_v[8] ));
 sg13g2_inv_1 _1070_ (.Y(_0435_),
    .A(\tiny_shader_top_inst.counter_v[7] ));
 sg13g2_inv_1 _1071_ (.Y(_0436_),
    .A(\tiny_shader_top_inst.counter_v[4] ));
 sg13g2_inv_1 _1072_ (.Y(_0437_),
    .A(net205));
 sg13g2_inv_2 _1073_ (.Y(_0438_),
    .A(\tiny_shader_top_inst.shader_execute_inst.regs[0][4] ));
 sg13g2_inv_1 _1074_ (.Y(_0439_),
    .A(_0017_));
 sg13g2_inv_1 _1075_ (.Y(_0440_),
    .A(net276));
 sg13g2_inv_1 _1076_ (.Y(_0441_),
    .A(net438));
 sg13g2_inv_1 _1077_ (.Y(_0442_),
    .A(\tiny_shader_top_inst.cur_time[8] ));
 sg13g2_inv_1 _1078_ (.Y(_0443_),
    .A(net284));
 sg13g2_inv_1 _1079_ (.Y(_0444_),
    .A(_0020_));
 sg13g2_inv_1 _1080_ (.Y(_0445_),
    .A(net302));
 sg13g2_inv_1 _1081_ (.Y(_0446_),
    .A(net298));
 sg13g2_inv_1 _1082_ (.Y(_0447_),
    .A(net462));
 sg13g2_inv_1 _1083_ (.Y(_0448_),
    .A(\tiny_shader_top_inst.shader_execute_inst.regs[0][5] ));
 sg13g2_inv_1 _1084_ (.Y(_0449_),
    .A(_0021_));
 sg13g2_inv_1 _1085_ (.Y(_0450_),
    .A(_0022_));
 sg13g2_inv_1 _1086_ (.Y(_0451_),
    .A(_0023_));
 sg13g2_inv_1 _1087_ (.Y(_0452_),
    .A(net458));
 sg13g2_inv_1 _1088_ (.Y(_0453_),
    .A(_0025_));
 sg13g2_inv_1 _1089_ (.Y(_0454_),
    .A(_0024_));
 sg13g2_inv_2 _1090_ (.Y(_0455_),
    .A(net457));
 sg13g2_inv_1 _1091_ (.Y(_0456_),
    .A(_0026_));
 sg13g2_inv_1 _1092_ (.Y(_0457_),
    .A(_0027_));
 sg13g2_inv_1 _1093_ (.Y(_0458_),
    .A(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[1] ));
 sg13g2_inv_1 _1094_ (.Y(_0459_),
    .A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[1] ));
 sg13g2_inv_1 _1095_ (.Y(_0460_),
    .A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[2] ));
 sg13g2_inv_1 _1096_ (.Y(_0461_),
    .A(net331));
 sg13g2_inv_1 _1097_ (.Y(_0462_),
    .A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[3] ));
 sg13g2_inv_1 _1098_ (.Y(_0463_),
    .A(net306));
 sg13g2_inv_1 _1099_ (.Y(_0464_),
    .A(net337));
 sg13g2_inv_1 _1100_ (.Y(_0465_),
    .A(net465));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_nor2b_1 _1102_ (.A(\tiny_shader_top_inst.counter_h[8] ),
    .B_N(_0013_),
    .Y(_0466_));
 sg13g2_nand2_1 _1103_ (.Y(_0467_),
    .A(net319),
    .B(net299));
 sg13g2_and2_1 _1104_ (.A(net264),
    .B(net130),
    .X(_0468_));
 sg13g2_nand2_1 _1105_ (.Y(_0469_),
    .A(\tiny_shader_top_inst.counter_h[2] ),
    .B(_0468_));
 sg13g2_nand4_1 _1106_ (.B(\tiny_shader_top_inst.counter_h[2] ),
    .C(\tiny_shader_top_inst.counter_h[1] ),
    .A(\tiny_shader_top_inst.counter_h[3] ),
    .Y(_0470_),
    .D(net130));
 sg13g2_nand3_1 _1107_ (.B(\tiny_shader_top_inst.counter_h[4] ),
    .C(\tiny_shader_top_inst.counter_h[5] ),
    .A(net316),
    .Y(_0471_));
 sg13g2_nor2_2 _1108_ (.A(_0470_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_inv_1 _1109_ (.Y(_0473_),
    .A(_0472_));
 sg13g2_o21ai_1 _1110_ (.B1(_0466_),
    .Y(_0474_),
    .A1(\tiny_shader_top_inst.counter_h[7] ),
    .A2(_0473_));
 sg13g2_nand3_1 _1111_ (.B(\tiny_shader_top_inst.counter_h[9] ),
    .C(_0474_),
    .A(_0430_),
    .Y(_0475_));
 sg13g2_inv_1 _1112_ (.Y(\tiny_shader_top_inst.next_vertical ),
    .A(net378));
 sg13g2_nand3_1 _1113_ (.B(net329),
    .C(_0472_),
    .A(net435),
    .Y(_0476_));
 sg13g2_nand4_1 _1114_ (.B(net332),
    .C(net329),
    .A(net435),
    .Y(_0477_),
    .D(_0472_));
 sg13g2_a21oi_1 _1115_ (.A1(net85),
    .A2(_0477_),
    .Y(_0081_),
    .B1(net376));
 sg13g2_nand2b_1 _1116_ (.Y(_0478_),
    .B(_0476_),
    .A_N(net332));
 sg13g2_a21oi_1 _1117_ (.A1(net333),
    .A2(_0478_),
    .Y(_0080_),
    .B1(net376));
 sg13g2_a21o_1 _1118_ (.A2(_0472_),
    .A1(net435),
    .B1(net329),
    .X(_0479_));
 sg13g2_a21oi_1 _1119_ (.A1(net330),
    .A2(_0479_),
    .Y(_0079_),
    .B1(net376));
 sg13g2_o21ai_1 _1120_ (.B1(_0428_),
    .Y(_0480_),
    .A1(_0467_),
    .A2(_0470_));
 sg13g2_a21oi_1 _1121_ (.A1(_0473_),
    .A2(net320),
    .Y(_0078_),
    .B1(net375));
 sg13g2_nor2_1 _1122_ (.A(net139),
    .B(_0470_),
    .Y(_0481_));
 sg13g2_xor2_1 _1123_ (.B(_0481_),
    .A(net299),
    .X(_0482_));
 sg13g2_nor2_1 _1124_ (.A(net375),
    .B(net300),
    .Y(_0077_));
 sg13g2_and3_1 _1125_ (.X(_0483_),
    .A(\tiny_shader_top_inst.counter_v[8] ),
    .B(\tiny_shader_top_inst.counter_v[7] ),
    .C(\tiny_shader_top_inst.counter_v[6] ));
 sg13g2_and2_1 _1126_ (.A(\tiny_shader_top_inst.counter_v[5] ),
    .B(_0483_),
    .X(_0484_));
 sg13g2_nor3_2 _1127_ (.A(\tiny_shader_top_inst.counter_v[9] ),
    .B(\tiny_shader_top_inst.counter_v[10] ),
    .C(_0484_),
    .Y(_0485_));
 sg13g2_nor2_1 _1128_ (.A(\tiny_shader_top_inst.counter_v[10] ),
    .B(_0485_),
    .Y(_0486_));
 sg13g2_and2_1 _1129_ (.A(\tiny_shader_top_inst.counter_v[1] ),
    .B(net119),
    .X(_0487_));
 sg13g2_nand3_1 _1130_ (.B(\tiny_shader_top_inst.counter_v[2] ),
    .C(_0487_),
    .A(\tiny_shader_top_inst.counter_v[3] ),
    .Y(_0488_));
 sg13g2_nor2_2 _1131_ (.A(_0436_),
    .B(_0488_),
    .Y(_0489_));
 sg13g2_nor3_1 _1132_ (.A(\tiny_shader_top_inst.counter_v[9] ),
    .B(\tiny_shader_top_inst.counter_v[5] ),
    .C(\tiny_shader_top_inst.counter_v[10] ),
    .Y(_0490_));
 sg13g2_nand3_1 _1133_ (.B(_0489_),
    .C(_0490_),
    .A(_0483_),
    .Y(_0491_));
 sg13g2_nor2b_1 _1134_ (.A(_0486_),
    .B_N(_0491_),
    .Y(_0492_));
 sg13g2_nand2b_2 _1135_ (.Y(_0493_),
    .B(net375),
    .A_N(_0492_));
 sg13g2_inv_4 _1136_ (.A(_0493_),
    .Y(\tiny_shader_top_inst.next_frame ));
 sg13g2_nand2_1 _1137_ (.Y(_0494_),
    .A(\tiny_shader_top_inst.x_subpos[0] ),
    .B(net205));
 sg13g2_nor3_2 _1138_ (.A(\tiny_shader_top_inst.x_subpos[1] ),
    .B(net262),
    .C(_0494_),
    .Y(_0000_));
 sg13g2_mux4_1 _1139_ (.S0(net3),
    .A0(\tiny_shader_top_inst.cur_time[0] ),
    .A1(\tiny_shader_top_inst.cur_time[7] ),
    .A2(_0485_),
    .A3(net438),
    .S1(net4),
    .X(uio_out[6]));
 sg13g2_a21oi_1 _1140_ (.A1(\tiny_shader_top_inst.counter_h[2] ),
    .A2(\tiny_shader_top_inst.counter_h[1] ),
    .Y(_0495_),
    .B1(\tiny_shader_top_inst.counter_h[3] ));
 sg13g2_nor2_1 _1141_ (.A(_0471_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_nand2_1 _1142_ (.Y(_0497_),
    .A(net435),
    .B(\tiny_shader_top_inst.counter_h[8] ));
 sg13g2_nor3_2 _1143_ (.A(_0471_),
    .B(_0495_),
    .C(_0497_),
    .Y(_0498_));
 sg13g2_nand2_1 _1144_ (.Y(_0499_),
    .A(\tiny_shader_top_inst.counter_h[9] ),
    .B(_0498_));
 sg13g2_nor2b_1 _1145_ (.A(_0013_),
    .B_N(\tiny_shader_top_inst.counter_h[8] ),
    .Y(_0500_));
 sg13g2_mux2_1 _1146_ (.A0(_0466_),
    .A1(_0500_),
    .S(_0496_),
    .X(_0501_));
 sg13g2_nor2_1 _1147_ (.A(\tiny_shader_top_inst.counter_h[9] ),
    .B(_0498_),
    .Y(_0502_));
 sg13g2_a21o_1 _1148_ (.A2(_0501_),
    .A1(_0499_),
    .B1(\tiny_shader_top_inst.counter_h[10] ),
    .X(_0503_));
 sg13g2_a21oi_1 _1149_ (.A1(\tiny_shader_top_inst.counter_h[9] ),
    .A2(_0498_),
    .Y(_0504_),
    .B1(_0430_));
 sg13g2_nor2b_1 _1150_ (.A(_0504_),
    .B_N(_0485_),
    .Y(_0505_));
 sg13g2_o21ai_1 _1151_ (.B1(_0505_),
    .Y(_0506_),
    .A1(_0502_),
    .A2(_0503_));
 sg13g2_mux4_1 _1152_ (.S0(net4),
    .A0(_0443_),
    .A1(_0506_),
    .A2(_0442_),
    .A3(_0441_),
    .S1(net3),
    .X(_0507_));
 sg13g2_inv_1 _1153_ (.Y(uio_out[7]),
    .A(_0507_));
 sg13g2_nor2_1 _1154_ (.A(net130),
    .B(net374),
    .Y(_0002_));
 sg13g2_nor2_1 _1155_ (.A(net264),
    .B(net130),
    .Y(_0508_));
 sg13g2_nor3_1 _1156_ (.A(_0468_),
    .B(net374),
    .C(_0508_),
    .Y(_0003_));
 sg13g2_xnor2_1 _1157_ (.Y(_0509_),
    .A(net303),
    .B(_0468_));
 sg13g2_nor2_1 _1158_ (.A(net374),
    .B(_0509_),
    .Y(_0004_));
 sg13g2_xnor2_1 _1159_ (.Y(_0510_),
    .A(net107),
    .B(_0469_));
 sg13g2_nor2_1 _1160_ (.A(net374),
    .B(net108),
    .Y(_0005_));
 sg13g2_and2_1 _1161_ (.A(net139),
    .B(_0470_),
    .X(_0511_));
 sg13g2_nor3_1 _1162_ (.A(net375),
    .B(_0481_),
    .C(net140),
    .Y(_0006_));
 sg13g2_xor2_1 _1163_ (.B(_0472_),
    .A(net269),
    .X(_0512_));
 sg13g2_nor2_1 _1164_ (.A(net376),
    .B(net270),
    .Y(_0007_));
 sg13g2_nand3_1 _1165_ (.B(\tiny_shader_top_inst.counter_v[10] ),
    .C(_0483_),
    .A(\tiny_shader_top_inst.counter_v[9] ),
    .Y(_0513_));
 sg13g2_or2_1 _1166_ (.X(_0514_),
    .B(net119),
    .A(\tiny_shader_top_inst.counter_v[1] ));
 sg13g2_nand4_1 _1167_ (.B(net258),
    .C(net287),
    .A(net334),
    .Y(_0515_),
    .D(_0514_));
 sg13g2_or4_1 _1168_ (.A(net326),
    .B(_0489_),
    .C(_0513_),
    .D(net335),
    .X(\tiny_shader_top_inst.timing_ver.sync ));
 sg13g2_nand3_1 _1169_ (.B(\tiny_shader_top_inst.counter_h[9] ),
    .C(\tiny_shader_top_inst.counter_h[8] ),
    .A(net85),
    .Y(_0516_));
 sg13g2_a21oi_1 _1170_ (.A1(_0428_),
    .A2(_0429_),
    .Y(_0517_),
    .B1(_0516_));
 sg13g2_a21oi_1 _1171_ (.A1(\tiny_shader_top_inst.counter_h[4] ),
    .A2(net299),
    .Y(_0518_),
    .B1(net435));
 sg13g2_o21ai_1 _1172_ (.B1(net435),
    .Y(_0519_),
    .A1(\tiny_shader_top_inst.counter_h[4] ),
    .A2(\tiny_shader_top_inst.counter_h[5] ));
 sg13g2_nor2b_1 _1173_ (.A(_0518_),
    .B_N(_0519_),
    .Y(_0520_));
 sg13g2_o21ai_1 _1174_ (.B1(_0517_),
    .Y(\tiny_shader_top_inst.hsync ),
    .A1(_0428_),
    .A2(_0520_));
 sg13g2_nand3b_1 _1175_ (.B(\tiny_shader_top_inst.spi_receiver_inst.spi_sclk_delayed ),
    .C(_0018_),
    .Y(_0521_),
    .A_N(\tiny_shader_top_inst.spi_receiver_inst.spi_sclk_sync ));
 sg13g2_nor2_1 _1176_ (.A(_0427_),
    .B(net431),
    .Y(_0522_));
 sg13g2_nand2_1 _1177_ (.Y(_0523_),
    .A(\tiny_shader_top_inst.spi_receiver_inst.spi_cnt[0] ),
    .B(net134));
 sg13g2_nor2_1 _1178_ (.A(net431),
    .B(_0523_),
    .Y(_0524_));
 sg13g2_nor4_1 _1179_ (.A(_0440_),
    .B(net47),
    .C(net431),
    .D(_0523_),
    .Y(_0001_));
 sg13g2_or2_2 _1180_ (.X(_0525_),
    .B(_0506_),
    .A(\tiny_shader_top_inst.shader_execute_inst.skip ));
 sg13g2_nor2_2 _1181_ (.A(net441),
    .B(net439),
    .Y(_0526_));
 sg13g2_or2_2 _1182_ (.X(_0527_),
    .B(\tiny_shader_top_inst.instr[7] ),
    .A(net440));
 sg13g2_nor3_2 _1183_ (.A(net448),
    .B(net446),
    .C(_0527_),
    .Y(_0528_));
 sg13g2_nor2_2 _1184_ (.A(net444),
    .B(net442),
    .Y(_0529_));
 sg13g2_or2_2 _1185_ (.X(_0530_),
    .B(net442),
    .A(net445));
 sg13g2_nor2b_1 _1186_ (.A(net448),
    .B_N(net446),
    .Y(_0531_));
 sg13g2_nand3_1 _1187_ (.B(_0529_),
    .C(_0531_),
    .A(_0526_),
    .Y(_0532_));
 sg13g2_nor4_2 _1188_ (.A(net448),
    .B(_0525_),
    .C(_0527_),
    .Y(_0533_),
    .D(_0530_));
 sg13g2_nand3_1 _1189_ (.B(net452),
    .C(_0444_),
    .A(net455),
    .Y(_0534_));
 sg13g2_nor2_2 _1190_ (.A(net454),
    .B(net451),
    .Y(_0535_));
 sg13g2_or2_1 _1191_ (.X(_0536_),
    .B(net451),
    .A(net454));
 sg13g2_a22oi_1 _1192_ (.Y(_0537_),
    .B1(\tiny_shader_top_inst.shader_execute_inst.regs[1][0] ),
    .B2(net432),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[2][0] ),
    .A1(_0432_));
 sg13g2_mux4_1 _1193_ (.S0(_0432_),
    .A0(_0444_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[2][0] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[1][0] ),
    .A3(net462),
    .S1(net432),
    .X(_0538_));
 sg13g2_nand3b_1 _1194_ (.B(net452),
    .C(net455),
    .Y(_0539_),
    .A_N(_0025_));
 sg13g2_nor2b_1 _1195_ (.A(net451),
    .B_N(net454),
    .Y(_0540_));
 sg13g2_nand3b_1 _1196_ (.B(\tiny_shader_top_inst.shader_execute_inst.regs[1][2] ),
    .C(net455),
    .Y(_0541_),
    .A_N(net452));
 sg13g2_nand2b_1 _1197_ (.Y(_0542_),
    .B(\tiny_shader_top_inst.shader_execute_inst.regs[2][2] ),
    .A_N(net455));
 sg13g2_nand4_1 _1198_ (.B(_0539_),
    .C(_0541_),
    .A(net428),
    .Y(_0543_),
    .D(_0542_));
 sg13g2_and2_1 _1199_ (.A(_0454_),
    .B(_0543_),
    .X(_0544_));
 sg13g2_mux4_1 _1200_ (.S0(_0432_),
    .A0(_0453_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[2][2] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[1][2] ),
    .A3(_0454_),
    .S1(net432),
    .X(_0545_));
 sg13g2_mux2_1 _1201_ (.A0(net393),
    .A1(_0545_),
    .S(_0532_),
    .X(_0546_));
 sg13g2_mux2_1 _1202_ (.A0(net175),
    .A1(_0546_),
    .S(_0533_),
    .X(_0082_));
 sg13g2_nand3_1 _1203_ (.B(net452),
    .C(\tiny_shader_top_inst.shader_execute_inst.regs[3][3] ),
    .A(net454),
    .Y(_0547_));
 sg13g2_o21ai_1 _1204_ (.B1(_0432_),
    .Y(_0548_),
    .A1(_0433_),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[2][3] ));
 sg13g2_nand2_1 _1205_ (.Y(_0549_),
    .A(net432),
    .B(\tiny_shader_top_inst.shader_execute_inst.regs[1][3] ));
 sg13g2_nand3_1 _1206_ (.B(_0548_),
    .C(_0549_),
    .A(_0547_),
    .Y(_0550_));
 sg13g2_mux4_1 _1207_ (.S0(_0432_),
    .A0(\tiny_shader_top_inst.shader_execute_inst.regs[3][3] ),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[2][3] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[1][3] ),
    .A3(_0456_),
    .S1(net432),
    .X(_0551_));
 sg13g2_nand3_1 _1208_ (.B(net452),
    .C(_0450_),
    .A(net455),
    .Y(_0552_));
 sg13g2_nor2b_1 _1209_ (.A(net454),
    .B_N(net451),
    .Y(_0553_));
 sg13g2_a22oi_1 _1210_ (.Y(_0554_),
    .B1(_0553_),
    .B2(\tiny_shader_top_inst.shader_execute_inst.regs[2][1] ),
    .A2(_0540_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[1][1] ));
 sg13g2_mux4_1 _1211_ (.S0(_0432_),
    .A0(_0450_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[2][1] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[1][1] ),
    .A3(net461),
    .S1(net432),
    .X(_0555_));
 sg13g2_mux2_1 _1212_ (.A0(net389),
    .A1(net390),
    .S(_0532_),
    .X(_0556_));
 sg13g2_mux2_1 _1213_ (.A0(net246),
    .A1(_0556_),
    .S(_0533_),
    .X(_0083_));
 sg13g2_nor2b_2 _1214_ (.A(net446),
    .B_N(net448),
    .Y(_0557_));
 sg13g2_nand2_1 _1215_ (.Y(_0558_),
    .A(_0526_),
    .B(_0557_));
 sg13g2_nand3_1 _1216_ (.B(_0529_),
    .C(_0557_),
    .A(_0526_),
    .Y(_0559_));
 sg13g2_nor4_2 _1217_ (.A(net447),
    .B(_0525_),
    .C(_0527_),
    .Y(_0560_),
    .D(_0530_));
 sg13g2_and3_1 _1218_ (.X(_0561_),
    .A(net454),
    .B(net451),
    .C(\tiny_shader_top_inst.shader_execute_inst.regs[3][4] ));
 sg13g2_nor2b_1 _1219_ (.A(net454),
    .B_N(\tiny_shader_top_inst.shader_execute_inst.regs[2][4] ),
    .Y(_0562_));
 sg13g2_nor2b_1 _1220_ (.A(net451),
    .B_N(\tiny_shader_top_inst.shader_execute_inst.regs[1][4] ),
    .Y(_0563_));
 sg13g2_nor4_2 _1221_ (.A(_0535_),
    .B(_0561_),
    .C(_0562_),
    .Y(_0564_),
    .D(_0563_));
 sg13g2_mux4_1 _1222_ (.S0(net453),
    .A0(_0439_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[2][4] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[1][4] ),
    .A3(\tiny_shader_top_inst.shader_execute_inst.regs[3][4] ),
    .S1(net456),
    .X(_0565_));
 sg13g2_mux2_1 _1223_ (.A0(net393),
    .A1(net387),
    .S(_0559_),
    .X(_0566_));
 sg13g2_mux2_1 _1224_ (.A0(net172),
    .A1(_0566_),
    .S(_0560_),
    .X(_0084_));
 sg13g2_nand3_1 _1225_ (.B(net451),
    .C(\tiny_shader_top_inst.shader_execute_inst.regs[3][5] ),
    .A(net454),
    .Y(_0567_));
 sg13g2_a22oi_1 _1226_ (.Y(_0568_),
    .B1(\tiny_shader_top_inst.shader_execute_inst.regs[1][5] ),
    .B2(net432),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[2][5] ),
    .A1(_0432_));
 sg13g2_nand2_1 _1227_ (.Y(_0569_),
    .A(_0567_),
    .B(_0568_));
 sg13g2_o21ai_1 _1228_ (.B1(_0457_),
    .Y(_0570_),
    .A1(_0535_),
    .A2(_0569_));
 sg13g2_mux4_1 _1229_ (.S0(_0432_),
    .A0(\tiny_shader_top_inst.shader_execute_inst.regs[3][5] ),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[2][5] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[1][5] ),
    .A3(_0457_),
    .S1(net432),
    .X(_0571_));
 sg13g2_mux2_1 _1230_ (.A0(net389),
    .A1(net386),
    .S(_0559_),
    .X(_0572_));
 sg13g2_mux2_1 _1231_ (.A0(net212),
    .A1(_0572_),
    .S(_0560_),
    .X(_0085_));
 sg13g2_or2_1 _1232_ (.X(_0573_),
    .B(_0506_),
    .A(_0431_));
 sg13g2_and2_2 _1233_ (.A(net440),
    .B(net439),
    .X(_0574_));
 sg13g2_nand2_1 _1234_ (.Y(_0575_),
    .A(net440),
    .B(net439));
 sg13g2_nand2_2 _1235_ (.Y(_0576_),
    .A(net444),
    .B(net442));
 sg13g2_nand2_1 _1236_ (.Y(_0577_),
    .A(net448),
    .B(net446));
 sg13g2_nor2_1 _1237_ (.A(_0527_),
    .B(_0577_),
    .Y(_0578_));
 sg13g2_nor3_1 _1238_ (.A(_0527_),
    .B(_0576_),
    .C(_0577_),
    .Y(_0579_));
 sg13g2_nor2b_1 _1239_ (.A(net442),
    .B_N(net444),
    .Y(_0580_));
 sg13g2_nand2b_2 _1240_ (.Y(_0581_),
    .B(net444),
    .A_N(net442));
 sg13g2_nand3b_1 _1241_ (.B(net445),
    .C(net443),
    .Y(_0582_),
    .A_N(net448));
 sg13g2_a21oi_1 _1242_ (.A1(_0526_),
    .A2(_0582_),
    .Y(_0583_),
    .B1(_0574_));
 sg13g2_and3_1 _1243_ (.X(_0584_),
    .A(net444),
    .B(_0526_),
    .C(_0557_));
 sg13g2_nor3_2 _1244_ (.A(_0527_),
    .B(_0577_),
    .C(_0581_),
    .Y(_0585_));
 sg13g2_and3_2 _1245_ (.X(_0586_),
    .A(_0526_),
    .B(_0531_),
    .C(_0580_));
 sg13g2_or4_1 _1246_ (.A(_0583_),
    .B(_0584_),
    .C(_0585_),
    .D(_0586_),
    .X(_0587_));
 sg13g2_a21o_1 _1247_ (.A2(_0580_),
    .A1(_0528_),
    .B1(_0587_),
    .X(_0588_));
 sg13g2_or2_2 _1248_ (.X(_0589_),
    .B(_0587_),
    .A(net385));
 sg13g2_inv_2 _1249_ (.Y(_0590_),
    .A(_0589_));
 sg13g2_nor2_2 _1250_ (.A(net385),
    .B(_0588_),
    .Y(_0591_));
 sg13g2_a22oi_1 _1251_ (.Y(_0592_),
    .B1(_0591_),
    .B2(_0575_),
    .A2(_0588_),
    .A1(net429));
 sg13g2_nand2b_1 _1252_ (.Y(_0593_),
    .B(_0592_),
    .A_N(_0573_));
 sg13g2_mux4_1 _1253_ (.S0(net446),
    .A0(\tiny_shader_top_inst.shader_execute_inst.regs[0][4] ),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[2][4] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[1][4] ),
    .A3(\tiny_shader_top_inst.shader_execute_inst.regs[3][4] ),
    .S1(net449),
    .X(_0594_));
 sg13g2_nand2_1 _1254_ (.Y(_0595_),
    .A(net387),
    .B(_0594_));
 sg13g2_xnor2_1 _1255_ (.Y(_0596_),
    .A(net387),
    .B(_0594_));
 sg13g2_mux4_1 _1256_ (.S0(net450),
    .A0(_0451_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[1][1] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[2][1] ),
    .A3(_0450_),
    .S1(net447),
    .X(_0597_));
 sg13g2_nand2_1 _1257_ (.Y(_0598_),
    .A(net388),
    .B(net384));
 sg13g2_mux4_1 _1258_ (.S0(net450),
    .A0(_0449_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[1][0] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[2][0] ),
    .A3(_0444_),
    .S1(net447),
    .X(_0599_));
 sg13g2_mux4_1 _1259_ (.S0(net450),
    .A0(_0021_),
    .A1(_0446_),
    .A2(_0445_),
    .A3(_0020_),
    .S1(net447),
    .X(_0600_));
 sg13g2_nand2_2 _1260_ (.Y(_0601_),
    .A(_0538_),
    .B(_0599_));
 sg13g2_nor2_1 _1261_ (.A(net388),
    .B(net384),
    .Y(_0602_));
 sg13g2_or2_1 _1262_ (.X(_0603_),
    .B(net384),
    .A(net388));
 sg13g2_and2_1 _1263_ (.A(_0598_),
    .B(_0603_),
    .X(_0604_));
 sg13g2_o21ai_1 _1264_ (.B1(_0598_),
    .Y(_0605_),
    .A1(_0601_),
    .A2(_0602_));
 sg13g2_mux4_1 _1265_ (.S0(net450),
    .A0(_0454_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[1][2] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[2][2] ),
    .A3(_0453_),
    .S1(net447),
    .X(_0606_));
 sg13g2_and2_1 _1266_ (.A(net392),
    .B(net381),
    .X(_0607_));
 sg13g2_xor2_1 _1267_ (.B(net381),
    .A(net392),
    .X(_0608_));
 sg13g2_mux4_1 _1268_ (.S0(net447),
    .A0(\tiny_shader_top_inst.shader_execute_inst.regs[0][3] ),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[2][3] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[1][3] ),
    .A3(\tiny_shader_top_inst.shader_execute_inst.regs[3][3] ),
    .S1(net449),
    .X(_0609_));
 sg13g2_and2_1 _1269_ (.A(net390),
    .B(net427),
    .X(_0610_));
 sg13g2_nor2_1 _1270_ (.A(net390),
    .B(net427),
    .Y(_0611_));
 sg13g2_or2_1 _1271_ (.X(_0612_),
    .B(net427),
    .A(net390));
 sg13g2_xor2_1 _1272_ (.B(net427),
    .A(net390),
    .X(_0613_));
 sg13g2_and2_1 _1273_ (.A(_0608_),
    .B(_0613_),
    .X(_0614_));
 sg13g2_a221oi_1 _1274_ (.B2(_0605_),
    .C1(_0610_),
    .B1(_0614_),
    .A1(_0607_),
    .Y(_0615_),
    .A2(_0612_));
 sg13g2_nand2b_2 _1275_ (.Y(_0616_),
    .B(net439),
    .A_N(net440));
 sg13g2_nor2_2 _1276_ (.A(_0581_),
    .B(_0616_),
    .Y(_0617_));
 sg13g2_or2_1 _1277_ (.X(_0618_),
    .B(_0616_),
    .A(_0581_));
 sg13g2_xor2_1 _1278_ (.B(_0615_),
    .A(_0596_),
    .X(_0619_));
 sg13g2_nor2_2 _1279_ (.A(_0530_),
    .B(_0616_),
    .Y(_0620_));
 sg13g2_nor2b_1 _1280_ (.A(net444),
    .B_N(net442),
    .Y(_0621_));
 sg13g2_nand2b_1 _1281_ (.Y(_0622_),
    .B(net442),
    .A_N(net444));
 sg13g2_nor2_2 _1282_ (.A(_0616_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_and2_1 _1283_ (.A(net382),
    .B(_0623_),
    .X(_0624_));
 sg13g2_nor2_2 _1284_ (.A(_0576_),
    .B(_0616_),
    .Y(_0625_));
 sg13g2_nand2b_2 _1285_ (.Y(_0626_),
    .B(_0625_),
    .A_N(net384));
 sg13g2_mux4_1 _1286_ (.S0(net449),
    .A0(\tiny_shader_top_inst.shader_execute_inst.regs[0][5] ),
    .A1(\tiny_shader_top_inst.shader_execute_inst.regs[1][5] ),
    .A2(\tiny_shader_top_inst.shader_execute_inst.regs[2][5] ),
    .A3(\tiny_shader_top_inst.shader_execute_inst.regs[3][5] ),
    .S1(net446),
    .X(_0627_));
 sg13g2_nor2_1 _1287_ (.A(_0594_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_a21oi_1 _1288_ (.A1(net387),
    .A2(net379),
    .Y(_0629_),
    .B1(_0599_));
 sg13g2_a21oi_1 _1289_ (.A1(net386),
    .A2(net379),
    .Y(_0630_),
    .B1(net383));
 sg13g2_or2_1 _1290_ (.X(_0631_),
    .B(_0630_),
    .A(_0629_));
 sg13g2_nor2_1 _1291_ (.A(_0626_),
    .B(_0631_),
    .Y(_0632_));
 sg13g2_nand2b_2 _1292_ (.Y(_0633_),
    .B(_0623_),
    .A_N(_0597_));
 sg13g2_a21oi_1 _1293_ (.A1(net390),
    .A2(net379),
    .Y(_0634_),
    .B1(net383));
 sg13g2_nor3_1 _1294_ (.A(_0629_),
    .B(_0633_),
    .C(_0634_),
    .Y(_0635_));
 sg13g2_nand2_2 _1295_ (.Y(_0636_),
    .A(net384),
    .B(_0623_));
 sg13g2_nand2_1 _1296_ (.Y(_0637_),
    .A(net388),
    .B(net379));
 sg13g2_nand2_1 _1297_ (.Y(_0638_),
    .A(net392),
    .B(net379));
 sg13g2_mux2_1 _1298_ (.A0(_0637_),
    .A1(_0638_),
    .S(net383),
    .X(_0639_));
 sg13g2_nor2_1 _1299_ (.A(_0636_),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_nor4_1 _1300_ (.A(_0624_),
    .B(_0632_),
    .C(_0635_),
    .D(_0640_),
    .Y(_0641_));
 sg13g2_nand3_1 _1301_ (.B(net383),
    .C(net379),
    .A(_0538_),
    .Y(_0642_));
 sg13g2_o21ai_1 _1302_ (.B1(net381),
    .Y(_0643_),
    .A1(_0633_),
    .A2(_0642_));
 sg13g2_inv_1 _1303_ (.Y(_0644_),
    .A(_0643_));
 sg13g2_nor3_1 _1304_ (.A(net427),
    .B(_0641_),
    .C(_0644_),
    .Y(_0645_));
 sg13g2_a221oi_1 _1305_ (.B2(_0594_),
    .C1(_0645_),
    .B1(_0620_),
    .A1(_0617_),
    .Y(_0646_),
    .A2(_0619_));
 sg13g2_nor2b_1 _1306_ (.A(net439),
    .B_N(net440),
    .Y(_0647_));
 sg13g2_nand2b_2 _1307_ (.Y(_0648_),
    .B(net440),
    .A_N(net439));
 sg13g2_nor2_2 _1308_ (.A(_0576_),
    .B(_0648_),
    .Y(_0649_));
 sg13g2_nor2b_1 _1309_ (.A(_0596_),
    .B_N(_0649_),
    .Y(_0650_));
 sg13g2_nor2_2 _1310_ (.A(_0558_),
    .B(_0576_),
    .Y(_0651_));
 sg13g2_nand2_2 _1311_ (.Y(_0652_),
    .A(_0621_),
    .B(_0647_));
 sg13g2_nand3_1 _1312_ (.B(_0557_),
    .C(_0580_),
    .A(_0526_),
    .Y(_0653_));
 sg13g2_nor2_1 _1313_ (.A(_0010_),
    .B(_0653_),
    .Y(_0654_));
 sg13g2_a221oi_1 _1314_ (.B2(\tiny_shader_top_inst.cur_time[7] ),
    .C1(_0654_),
    .B1(_0586_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.user_i[4] ),
    .Y(_0655_),
    .A2(_0585_));
 sg13g2_o21ai_1 _1315_ (.B1(_0655_),
    .Y(_0656_),
    .A1(_0594_),
    .A2(_0652_));
 sg13g2_nor4_2 _1316_ (.A(net448),
    .B(net446),
    .C(_0527_),
    .Y(_0657_),
    .D(_0576_));
 sg13g2_a22oi_1 _1317_ (.Y(_0658_),
    .B1(_0657_),
    .B2(net390),
    .A2(_0651_),
    .A1(_0571_));
 sg13g2_inv_1 _1318_ (.Y(_0659_),
    .A(_0658_));
 sg13g2_nor2_1 _1319_ (.A(_0530_),
    .B(_0648_),
    .Y(_0660_));
 sg13g2_nand2_2 _1320_ (.Y(_0661_),
    .A(_0529_),
    .B(_0647_));
 sg13g2_nor2_2 _1321_ (.A(_0581_),
    .B(_0648_),
    .Y(_0662_));
 sg13g2_o21ai_1 _1322_ (.B1(_0662_),
    .Y(_0663_),
    .A1(net387),
    .A2(_0594_));
 sg13g2_o21ai_1 _1323_ (.B1(_0663_),
    .Y(_0664_),
    .A1(_0595_),
    .A2(_0661_));
 sg13g2_nor4_2 _1324_ (.A(_0650_),
    .B(_0656_),
    .C(_0659_),
    .Y(_0665_),
    .D(_0664_));
 sg13g2_nor2_2 _1325_ (.A(net440),
    .B(_0589_),
    .Y(_0666_));
 sg13g2_or2_1 _1326_ (.X(_0667_),
    .B(_0589_),
    .A(net440));
 sg13g2_nand2_2 _1327_ (.Y(_0668_),
    .A(net462),
    .B(net459));
 sg13g2_inv_1 _1328_ (.Y(_0669_),
    .A(_0668_));
 sg13g2_nand2_1 _1329_ (.Y(_0670_),
    .A(_0452_),
    .B(_0455_));
 sg13g2_nand2_2 _1330_ (.Y(_0671_),
    .A(net458),
    .B(net457));
 sg13g2_nand2b_1 _1331_ (.Y(_0672_),
    .B(net458),
    .A_N(net459));
 sg13g2_nand2_1 _1332_ (.Y(_0673_),
    .A(_0671_),
    .B(_0672_));
 sg13g2_nor2b_2 _1333_ (.A(net458),
    .B_N(net457),
    .Y(_0674_));
 sg13g2_nor2_2 _1334_ (.A(net462),
    .B(net459),
    .Y(_0675_));
 sg13g2_nand2b_1 _1335_ (.Y(_0676_),
    .B(_0674_),
    .A_N(_0675_));
 sg13g2_o21ai_1 _1336_ (.B1(_0676_),
    .Y(_0677_),
    .A1(_0668_),
    .A2(_0670_));
 sg13g2_or3_1 _1337_ (.A(net466),
    .B(_0673_),
    .C(_0677_),
    .X(_0678_));
 sg13g2_and2_1 _1338_ (.A(net385),
    .B(_0678_),
    .X(_0679_));
 sg13g2_nand2_1 _1339_ (.Y(_0680_),
    .A(net459),
    .B(_0674_));
 sg13g2_nand3_1 _1340_ (.B(_0670_),
    .C(_0680_),
    .A(net466),
    .Y(_0681_));
 sg13g2_nor2_2 _1341_ (.A(_0452_),
    .B(net457),
    .Y(_0682_));
 sg13g2_nor2b_1 _1342_ (.A(_0671_),
    .B_N(_0675_),
    .Y(_0683_));
 sg13g2_a21oi_1 _1343_ (.A1(_0668_),
    .A2(_0682_),
    .Y(_0684_),
    .B1(_0683_));
 sg13g2_nand2b_1 _1344_ (.Y(_0685_),
    .B(_0684_),
    .A_N(_0681_));
 sg13g2_nor2_1 _1345_ (.A(net429),
    .B(_0685_),
    .Y(_0686_));
 sg13g2_a21oi_1 _1346_ (.A1(_0438_),
    .A2(net428),
    .Y(_0687_),
    .B1(_0686_));
 sg13g2_a22oi_1 _1347_ (.Y(_0688_),
    .B1(_0679_),
    .B2(_0687_),
    .A2(_0574_),
    .A1(net444));
 sg13g2_and3_1 _1348_ (.X(_0689_),
    .A(_0665_),
    .B(_0667_),
    .C(_0688_));
 sg13g2_a221oi_1 _1349_ (.B2(_0646_),
    .C1(_0593_),
    .B1(_0689_),
    .A1(_0463_),
    .Y(_0690_),
    .A2(_0666_));
 sg13g2_a21o_1 _1350_ (.A2(_0593_),
    .A1(net466),
    .B1(_0690_),
    .X(_0086_));
 sg13g2_nand2_1 _1351_ (.Y(_0691_),
    .A(net375),
    .B(_0492_));
 sg13g2_inv_1 _1352_ (.Y(_0692_),
    .A(net353));
 sg13g2_a22oi_1 _1353_ (.Y(_0693_),
    .B1(_0692_),
    .B2(net119),
    .A2(net378),
    .A1(_0042_));
 sg13g2_inv_1 _1354_ (.Y(_0087_),
    .A(net120));
 sg13g2_nand2_1 _1355_ (.Y(_0694_),
    .A(net117),
    .B(net377));
 sg13g2_nor2b_1 _1356_ (.A(_0487_),
    .B_N(_0514_),
    .Y(_0695_));
 sg13g2_o21ai_1 _1357_ (.B1(_0694_),
    .Y(_0088_),
    .A1(_0691_),
    .A2(_0695_));
 sg13g2_and3_1 _1358_ (.X(_0696_),
    .A(net287),
    .B(net375),
    .C(_0487_));
 sg13g2_a21oi_1 _1359_ (.A1(net375),
    .A2(_0487_),
    .Y(_0697_),
    .B1(net287));
 sg13g2_nor3_1 _1360_ (.A(\tiny_shader_top_inst.next_frame ),
    .B(_0696_),
    .C(net288),
    .Y(_0089_));
 sg13g2_o21ai_1 _1361_ (.B1(_0493_),
    .Y(_0698_),
    .A1(net258),
    .A2(_0696_));
 sg13g2_a21oi_1 _1362_ (.A1(net258),
    .A2(_0696_),
    .Y(_0090_),
    .B1(_0698_));
 sg13g2_nand2_1 _1363_ (.Y(_0699_),
    .A(net95),
    .B(net377));
 sg13g2_xnor2_1 _1364_ (.Y(_0700_),
    .A(\tiny_shader_top_inst.counter_v[4] ),
    .B(_0488_));
 sg13g2_o21ai_1 _1365_ (.B1(_0699_),
    .Y(_0091_),
    .A1(net353),
    .A2(_0700_));
 sg13g2_nand2_1 _1366_ (.Y(_0701_),
    .A(net326),
    .B(net377));
 sg13g2_xnor2_1 _1367_ (.Y(_0702_),
    .A(net326),
    .B(_0489_));
 sg13g2_o21ai_1 _1368_ (.B1(_0701_),
    .Y(_0092_),
    .A1(net353),
    .A2(_0702_));
 sg13g2_nand2_1 _1369_ (.Y(_0703_),
    .A(net121),
    .B(net377));
 sg13g2_nand3_1 _1370_ (.B(\tiny_shader_top_inst.counter_v[5] ),
    .C(_0489_),
    .A(\tiny_shader_top_inst.counter_v[6] ),
    .Y(_0704_));
 sg13g2_a21o_1 _1371_ (.A2(_0489_),
    .A1(\tiny_shader_top_inst.counter_v[5] ),
    .B1(\tiny_shader_top_inst.counter_v[6] ),
    .X(_0705_));
 sg13g2_and2_1 _1372_ (.A(_0704_),
    .B(_0705_),
    .X(_0706_));
 sg13g2_o21ai_1 _1373_ (.B1(_0703_),
    .Y(_0093_),
    .A1(net353),
    .A2(_0706_));
 sg13g2_nand2_1 _1374_ (.Y(_0707_),
    .A(net97),
    .B(net377));
 sg13g2_xnor2_1 _1375_ (.Y(_0708_),
    .A(\tiny_shader_top_inst.counter_v[7] ),
    .B(_0704_));
 sg13g2_o21ai_1 _1376_ (.B1(_0707_),
    .Y(_0094_),
    .A1(net353),
    .A2(_0708_));
 sg13g2_nand2_1 _1377_ (.Y(_0709_),
    .A(_0484_),
    .B(_0489_));
 sg13g2_o21ai_1 _1378_ (.B1(_0434_),
    .Y(_0710_),
    .A1(_0435_),
    .A2(_0704_));
 sg13g2_a21oi_1 _1379_ (.A1(_0709_),
    .A2(_0710_),
    .Y(_0711_),
    .B1(net353));
 sg13g2_a21o_1 _1380_ (.A2(net377),
    .A1(net145),
    .B1(_0711_),
    .X(_0095_));
 sg13g2_nand2_1 _1381_ (.Y(_0712_),
    .A(net113),
    .B(net377));
 sg13g2_nand3_1 _1382_ (.B(_0484_),
    .C(_0489_),
    .A(\tiny_shader_top_inst.counter_v[9] ),
    .Y(_0713_));
 sg13g2_xnor2_1 _1383_ (.Y(_0714_),
    .A(\tiny_shader_top_inst.counter_v[9] ),
    .B(_0709_));
 sg13g2_o21ai_1 _1384_ (.B1(_0712_),
    .Y(_0096_),
    .A1(net353),
    .A2(_0714_));
 sg13g2_nand2_1 _1385_ (.Y(_0715_),
    .A(net101),
    .B(net377));
 sg13g2_xnor2_1 _1386_ (.Y(_0716_),
    .A(\tiny_shader_top_inst.counter_v[10] ),
    .B(_0713_));
 sg13g2_o21ai_1 _1387_ (.B1(_0715_),
    .Y(_0097_),
    .A1(net353),
    .A2(_0716_));
 sg13g2_nor4_1 _1388_ (.A(\tiny_shader_top_inst.cur_time[1] ),
    .B(\tiny_shader_top_inst.cur_time[3] ),
    .C(\tiny_shader_top_inst.cur_time[4] ),
    .D(\tiny_shader_top_inst.cur_time[5] ),
    .Y(_0717_));
 sg13g2_nand3b_1 _1389_ (.B(_0717_),
    .C(\tiny_shader_top_inst.cur_time[0] ),
    .Y(_0718_),
    .A_N(\tiny_shader_top_inst.cur_time[7] ));
 sg13g2_nor4_1 _1390_ (.A(net331),
    .B(_0464_),
    .C(net250),
    .D(_0718_),
    .Y(_0719_));
 sg13g2_a21oi_1 _1391_ (.A1(\tiny_shader_top_inst.next_frame ),
    .A2(net338),
    .Y(_0098_),
    .B1(_0465_));
 sg13g2_o21ai_1 _1392_ (.B1(_0529_),
    .Y(_0720_),
    .A1(_0528_),
    .A2(_0578_));
 sg13g2_nor2_2 _1393_ (.A(_0525_),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_mux2_1 _1394_ (.A0(net216),
    .A1(net393),
    .S(_0721_),
    .X(_0099_));
 sg13g2_mux2_1 _1395_ (.A0(net232),
    .A1(net388),
    .S(_0721_),
    .X(_0100_));
 sg13g2_and2_1 _1396_ (.A(net241),
    .B(_0506_),
    .X(_0722_));
 sg13g2_nor2_1 _1397_ (.A(_0448_),
    .B(net386),
    .Y(_0723_));
 sg13g2_nand2b_1 _1398_ (.Y(_0724_),
    .B(\tiny_shader_top_inst.shader_execute_inst.regs[0][3] ),
    .A_N(net391));
 sg13g2_nand2_1 _1399_ (.Y(_0725_),
    .A(_0455_),
    .B(net391));
 sg13g2_a21oi_1 _1400_ (.A1(net428),
    .A2(_0543_),
    .Y(_0726_),
    .B1(_0454_));
 sg13g2_nor2_1 _1401_ (.A(_0544_),
    .B(_0726_),
    .Y(_0727_));
 sg13g2_o21ai_1 _1402_ (.B1(_0725_),
    .Y(_0728_),
    .A1(_0544_),
    .A2(_0726_));
 sg13g2_nor2_1 _1403_ (.A(_0023_),
    .B(net389),
    .Y(_0729_));
 sg13g2_or2_1 _1404_ (.X(_0730_),
    .B(net389),
    .A(_0023_));
 sg13g2_a22oi_1 _1405_ (.Y(_0731_),
    .B1(net389),
    .B2(_0023_),
    .A2(net393),
    .A1(_0447_));
 sg13g2_nor2_1 _1406_ (.A(_0729_),
    .B(_0731_),
    .Y(_0732_));
 sg13g2_nor2_1 _1407_ (.A(_0452_),
    .B(net392),
    .Y(_0733_));
 sg13g2_nor2_1 _1408_ (.A(_0438_),
    .B(net387),
    .Y(_0734_));
 sg13g2_a21oi_1 _1409_ (.A1(_0725_),
    .A2(_0733_),
    .Y(_0735_),
    .B1(_0734_));
 sg13g2_o21ai_1 _1410_ (.B1(_0735_),
    .Y(_0736_),
    .A1(_0728_),
    .A2(_0732_));
 sg13g2_o21ai_1 _1411_ (.B1(_0017_),
    .Y(_0737_),
    .A1(_0535_),
    .A2(_0564_));
 sg13g2_o21ai_1 _1412_ (.B1(_0737_),
    .Y(_0738_),
    .A1(_0017_),
    .A2(_0564_));
 sg13g2_nand4_1 _1413_ (.B(_0534_),
    .C(net428),
    .A(net462),
    .Y(_0739_),
    .D(_0537_));
 sg13g2_nand4_1 _1414_ (.B(_0731_),
    .C(_0738_),
    .A(_0730_),
    .Y(_0740_),
    .D(_0739_));
 sg13g2_o21ai_1 _1415_ (.B1(_0736_),
    .Y(_0741_),
    .A1(_0728_),
    .A2(_0740_));
 sg13g2_nor2_1 _1416_ (.A(_0734_),
    .B(_0738_),
    .Y(_0742_));
 sg13g2_a221oi_1 _1417_ (.B2(_0741_),
    .C1(_0742_),
    .B1(_0724_),
    .A1(_0448_),
    .Y(_0743_),
    .A2(net386));
 sg13g2_nand2_1 _1418_ (.Y(_0744_),
    .A(_0578_),
    .B(_0621_));
 sg13g2_or3_1 _1419_ (.A(_0723_),
    .B(_0743_),
    .C(_0744_),
    .X(_0745_));
 sg13g2_and2_1 _1420_ (.A(net447),
    .B(_0744_),
    .X(_0746_));
 sg13g2_o21ai_1 _1421_ (.B1(_0746_),
    .Y(_0747_),
    .A1(_0723_),
    .A2(_0743_));
 sg13g2_nand2_1 _1422_ (.Y(_0748_),
    .A(_0026_),
    .B(net391));
 sg13g2_o21ai_1 _1423_ (.B1(_0570_),
    .Y(_0749_),
    .A1(_0457_),
    .A2(net386));
 sg13g2_xnor2_1 _1424_ (.Y(_0750_),
    .A(_0021_),
    .B(net393));
 sg13g2_nor2b_1 _1425_ (.A(net461),
    .B_N(net389),
    .Y(_0751_));
 sg13g2_nand4_1 _1426_ (.B(net429),
    .C(_0552_),
    .A(net461),
    .Y(_0752_),
    .D(_0554_));
 sg13g2_o21ai_1 _1427_ (.B1(_0752_),
    .Y(_0753_),
    .A1(_0026_),
    .A2(_0550_));
 sg13g2_nor4_1 _1428_ (.A(_0727_),
    .B(_0750_),
    .C(_0751_),
    .D(_0753_),
    .Y(_0754_));
 sg13g2_nand4_1 _1429_ (.B(_0748_),
    .C(_0749_),
    .A(_0738_),
    .Y(_0755_),
    .D(_0754_));
 sg13g2_nand2b_1 _1430_ (.Y(_0756_),
    .B(_0755_),
    .A_N(_0528_));
 sg13g2_nand2b_1 _1431_ (.Y(_0757_),
    .B(_0558_),
    .A_N(_0755_));
 sg13g2_nand3_1 _1432_ (.B(_0756_),
    .C(_0757_),
    .A(_0621_),
    .Y(_0758_));
 sg13g2_nand3_1 _1433_ (.B(_0747_),
    .C(_0758_),
    .A(_0745_),
    .Y(_0759_));
 sg13g2_nor3_1 _1434_ (.A(_0527_),
    .B(_0573_),
    .C(_0622_),
    .Y(_0760_));
 sg13g2_a21o_1 _1435_ (.A2(_0760_),
    .A1(_0759_),
    .B1(_0722_),
    .X(_0101_));
 sg13g2_a21oi_1 _1436_ (.A1(\tiny_shader_top_inst.shader_execute_inst.regs[0][4] ),
    .A2(_0017_),
    .Y(_0761_),
    .B1(_0535_));
 sg13g2_a21oi_1 _1437_ (.A1(net385),
    .A2(_0761_),
    .Y(_0762_),
    .B1(_0593_));
 sg13g2_nor2_1 _1438_ (.A(net462),
    .B(net352),
    .Y(_0763_));
 sg13g2_o21ai_1 _1439_ (.B1(_0626_),
    .Y(_0764_),
    .A1(_0633_),
    .A2(_0642_));
 sg13g2_o21ai_1 _1440_ (.B1(_0642_),
    .Y(_0765_),
    .A1(net383),
    .A2(_0637_));
 sg13g2_nand2_2 _1441_ (.Y(_0766_),
    .A(net384),
    .B(_0625_));
 sg13g2_a21o_1 _1442_ (.A2(_0638_),
    .A1(net383),
    .B1(_0634_),
    .X(_0767_));
 sg13g2_and2_1 _1443_ (.A(net381),
    .B(_0625_),
    .X(_0768_));
 sg13g2_a21oi_1 _1444_ (.A1(_0764_),
    .A2(_0765_),
    .Y(_0769_),
    .B1(_0768_));
 sg13g2_o21ai_1 _1445_ (.B1(_0769_),
    .Y(_0770_),
    .A1(_0766_),
    .A2(_0767_));
 sg13g2_o21ai_1 _1446_ (.B1(net381),
    .Y(_0771_),
    .A1(_0626_),
    .A2(_0631_));
 sg13g2_nor2b_1 _1447_ (.A(_0609_),
    .B_N(_0771_),
    .Y(_0772_));
 sg13g2_nand2b_1 _1448_ (.Y(_0773_),
    .B(net383),
    .A_N(net393));
 sg13g2_o21ai_1 _1449_ (.B1(_0601_),
    .Y(_0774_),
    .A1(_0617_),
    .A2(_0649_));
 sg13g2_a21oi_1 _1450_ (.A1(_0599_),
    .A2(_0620_),
    .Y(_0775_),
    .B1(_0662_));
 sg13g2_o21ai_1 _1451_ (.B1(_0775_),
    .Y(_0776_),
    .A1(_0601_),
    .A2(_0661_));
 sg13g2_nand2b_1 _1452_ (.Y(_0777_),
    .B(_0774_),
    .A_N(_0776_));
 sg13g2_a22oi_1 _1453_ (.Y(_0778_),
    .B1(_0586_),
    .B2(\tiny_shader_top_inst.cur_time[3] ),
    .A2(_0585_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.user_i[0] ));
 sg13g2_o21ai_1 _1454_ (.B1(_0778_),
    .Y(_0779_),
    .A1(_0028_),
    .A2(_0653_));
 sg13g2_a21oi_1 _1455_ (.A1(net388),
    .A2(_0651_),
    .Y(_0780_),
    .B1(_0779_));
 sg13g2_o21ai_1 _1456_ (.B1(_0780_),
    .Y(_0781_),
    .A1(_0599_),
    .A2(_0652_));
 sg13g2_a221oi_1 _1457_ (.B2(_0777_),
    .C1(_0781_),
    .B1(_0773_),
    .A1(_0770_),
    .Y(_0782_),
    .A2(_0772_));
 sg13g2_a21oi_1 _1458_ (.A1(_0455_),
    .A2(_0675_),
    .Y(_0783_),
    .B1(_0438_));
 sg13g2_o21ai_1 _1459_ (.B1(_0438_),
    .Y(_0784_),
    .A1(_0447_),
    .A2(_0680_));
 sg13g2_nand2_1 _1460_ (.Y(_0785_),
    .A(net460),
    .B(net458));
 sg13g2_nor2_1 _1461_ (.A(_0455_),
    .B(_0785_),
    .Y(_0786_));
 sg13g2_a221oi_1 _1462_ (.B2(net462),
    .C1(_0784_),
    .B1(_0786_),
    .A1(_0668_),
    .Y(_0787_),
    .A2(_0682_));
 sg13g2_a21oi_1 _1463_ (.A1(_0676_),
    .A2(_0783_),
    .Y(_0788_),
    .B1(_0787_));
 sg13g2_nand3_1 _1464_ (.B(_0452_),
    .C(_0455_),
    .A(net459),
    .Y(_0789_));
 sg13g2_nor2_1 _1465_ (.A(net459),
    .B(_0671_),
    .Y(_0790_));
 sg13g2_o21ai_1 _1466_ (.B1(_0789_),
    .Y(_0791_),
    .A1(net460),
    .A2(_0671_));
 sg13g2_o21ai_1 _1467_ (.B1(net385),
    .Y(_0792_),
    .A1(_0788_),
    .A2(_0791_));
 sg13g2_or2_1 _1468_ (.X(_0793_),
    .B(_0792_),
    .A(net428));
 sg13g2_nand2_1 _1469_ (.Y(_0794_),
    .A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[0] ),
    .B(_0590_));
 sg13g2_a22oi_1 _1470_ (.Y(_0795_),
    .B1(_0666_),
    .B2(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[0] ),
    .A2(_0574_),
    .A1(net455));
 sg13g2_nand4_1 _1471_ (.B(_0782_),
    .C(_0793_),
    .A(net352),
    .Y(_0796_),
    .D(_0795_));
 sg13g2_nor2b_1 _1472_ (.A(_0763_),
    .B_N(_0796_),
    .Y(_0102_));
 sg13g2_nand2b_1 _1473_ (.Y(_0797_),
    .B(net461),
    .A_N(net352));
 sg13g2_a21oi_2 _1474_ (.B1(_0599_),
    .Y(_0798_),
    .A2(net380),
    .A1(net388));
 sg13g2_a21oi_1 _1475_ (.A1(net392),
    .A2(net379),
    .Y(_0799_),
    .B1(net383));
 sg13g2_nor3_1 _1476_ (.A(_0626_),
    .B(_0798_),
    .C(_0799_),
    .Y(_0800_));
 sg13g2_nand3_1 _1477_ (.B(_0599_),
    .C(net380),
    .A(net387),
    .Y(_0801_));
 sg13g2_a21oi_2 _1478_ (.B1(_0599_),
    .Y(_0802_),
    .A2(net379),
    .A1(net390));
 sg13g2_a21oi_1 _1479_ (.A1(net387),
    .A2(net380),
    .Y(_0803_),
    .B1(_0600_));
 sg13g2_nor3_1 _1480_ (.A(_0766_),
    .B(_0802_),
    .C(_0803_),
    .Y(_0804_));
 sg13g2_a21oi_1 _1481_ (.A1(net393),
    .A2(net380),
    .Y(_0805_),
    .B1(_0600_));
 sg13g2_nor3_1 _1482_ (.A(_0633_),
    .B(_0798_),
    .C(_0805_),
    .Y(_0806_));
 sg13g2_or3_1 _1483_ (.A(_0633_),
    .B(_0798_),
    .C(_0805_),
    .X(_0807_));
 sg13g2_nor4_1 _1484_ (.A(_0768_),
    .B(_0800_),
    .C(_0804_),
    .D(_0806_),
    .Y(_0808_));
 sg13g2_nand3_1 _1485_ (.B(_0600_),
    .C(net380),
    .A(net386),
    .Y(_0809_));
 sg13g2_o21ai_1 _1486_ (.B1(net381),
    .Y(_0810_),
    .A1(_0626_),
    .A2(_0809_));
 sg13g2_nand2b_1 _1487_ (.Y(_0811_),
    .B(_0810_),
    .A_N(net427));
 sg13g2_xnor2_1 _1488_ (.Y(_0812_),
    .A(_0601_),
    .B(_0604_));
 sg13g2_a22oi_1 _1489_ (.Y(_0813_),
    .B1(_0812_),
    .B2(_0617_),
    .A2(_0620_),
    .A1(net384));
 sg13g2_o21ai_1 _1490_ (.B1(_0813_),
    .Y(_0814_),
    .A1(_0808_),
    .A2(_0811_));
 sg13g2_and2_1 _1491_ (.A(_0604_),
    .B(_0649_),
    .X(_0815_));
 sg13g2_a22oi_1 _1492_ (.Y(_0816_),
    .B1(_0586_),
    .B2(\tiny_shader_top_inst.cur_time[4] ),
    .A2(_0585_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.user_i[1] ));
 sg13g2_o21ai_1 _1493_ (.B1(_0816_),
    .Y(_0817_),
    .A1(_0458_),
    .A2(_0653_));
 sg13g2_a21oi_1 _1494_ (.A1(net393),
    .A2(_0657_),
    .Y(_0818_),
    .B1(_0817_));
 sg13g2_o21ai_1 _1495_ (.B1(_0818_),
    .Y(_0819_),
    .A1(net384),
    .A2(_0652_));
 sg13g2_a22oi_1 _1496_ (.Y(_0820_),
    .B1(_0662_),
    .B2(_0603_),
    .A2(_0651_),
    .A1(net392));
 sg13g2_o21ai_1 _1497_ (.B1(_0820_),
    .Y(_0821_),
    .A1(_0598_),
    .A2(_0661_));
 sg13g2_nor3_2 _1498_ (.A(_0815_),
    .B(_0819_),
    .C(_0821_),
    .Y(_0822_));
 sg13g2_inv_1 _1499_ (.Y(_0823_),
    .A(_0822_));
 sg13g2_nor2_1 _1500_ (.A(net459),
    .B(net458),
    .Y(_0824_));
 sg13g2_xnor2_1 _1501_ (.Y(_0825_),
    .A(net459),
    .B(\tiny_shader_top_inst.shader_execute_inst.regs[0][2] ));
 sg13g2_a21oi_1 _1502_ (.A1(net466),
    .A2(_0825_),
    .Y(_0826_),
    .B1(net457));
 sg13g2_nor2_1 _1503_ (.A(net466),
    .B(_0455_),
    .Y(_0827_));
 sg13g2_o21ai_1 _1504_ (.B1(net457),
    .Y(_0828_),
    .A1(net466),
    .A2(_0785_));
 sg13g2_a22oi_1 _1505_ (.Y(_0829_),
    .B1(_0828_),
    .B2(net463),
    .A2(_0827_),
    .A1(_0824_));
 sg13g2_o21ai_1 _1506_ (.B1(_0829_),
    .Y(_0830_),
    .A1(net462),
    .A2(_0826_));
 sg13g2_nand2_1 _1507_ (.Y(_0831_),
    .A(net385),
    .B(_0830_));
 sg13g2_a21oi_1 _1508_ (.A1(net452),
    .A2(_0574_),
    .Y(_0832_),
    .B1(_0666_));
 sg13g2_o21ai_1 _1509_ (.B1(_0832_),
    .Y(_0833_),
    .A1(net428),
    .A2(_0831_));
 sg13g2_nor3_1 _1510_ (.A(_0814_),
    .B(_0823_),
    .C(_0833_),
    .Y(_0834_));
 sg13g2_o21ai_1 _1511_ (.B1(net352),
    .Y(_0835_),
    .A1(net314),
    .A2(_0667_));
 sg13g2_o21ai_1 _1512_ (.B1(_0797_),
    .Y(_0103_),
    .A1(_0834_),
    .A2(_0835_));
 sg13g2_nor2_1 _1513_ (.A(net458),
    .B(net352),
    .Y(_0836_));
 sg13g2_or2_1 _1514_ (.X(_0837_),
    .B(_0609_),
    .A(net381));
 sg13g2_nor2_1 _1515_ (.A(_0636_),
    .B(_0642_),
    .Y(_0838_));
 sg13g2_nor2_1 _1516_ (.A(_0633_),
    .B(_0639_),
    .Y(_0839_));
 sg13g2_nor2_1 _1517_ (.A(_0631_),
    .B(_0766_),
    .Y(_0840_));
 sg13g2_nor2_1 _1518_ (.A(_0626_),
    .B(_0767_),
    .Y(_0841_));
 sg13g2_nor4_1 _1519_ (.A(_0838_),
    .B(_0839_),
    .C(_0840_),
    .D(_0841_),
    .Y(_0842_));
 sg13g2_nor2_1 _1520_ (.A(_0837_),
    .B(_0842_),
    .Y(_0843_));
 sg13g2_nand2_1 _1521_ (.Y(_0844_),
    .A(_0607_),
    .B(_0660_));
 sg13g2_o21ai_1 _1522_ (.B1(_0662_),
    .Y(_0845_),
    .A1(net392),
    .A2(net382));
 sg13g2_nor2_1 _1523_ (.A(net382),
    .B(_0652_),
    .Y(_0846_));
 sg13g2_a221oi_1 _1524_ (.B2(net388),
    .C1(_0846_),
    .B1(_0657_),
    .A1(net391),
    .Y(_0847_),
    .A2(_0651_));
 sg13g2_a22oi_1 _1525_ (.Y(_0848_),
    .B1(_0586_),
    .B2(\tiny_shader_top_inst.cur_time[5] ),
    .A2(_0585_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.user_i[2] ));
 sg13g2_o21ai_1 _1526_ (.B1(_0848_),
    .Y(_0849_),
    .A1(_0008_),
    .A2(_0653_));
 sg13g2_a221oi_1 _1527_ (.B2(_0608_),
    .C1(_0849_),
    .B1(_0649_),
    .A1(net381),
    .Y(_0850_),
    .A2(_0620_));
 sg13g2_nand4_1 _1528_ (.B(_0845_),
    .C(_0847_),
    .A(_0844_),
    .Y(_0851_),
    .D(_0850_));
 sg13g2_o21ai_1 _1529_ (.B1(_0617_),
    .Y(_0852_),
    .A1(_0605_),
    .A2(_0608_));
 sg13g2_a21oi_1 _1530_ (.A1(_0605_),
    .A2(_0608_),
    .Y(_0853_),
    .B1(_0852_));
 sg13g2_nor3_1 _1531_ (.A(_0843_),
    .B(_0851_),
    .C(_0853_),
    .Y(_0854_));
 sg13g2_nand2_1 _1532_ (.Y(_0855_),
    .A(_0670_),
    .B(_0676_));
 sg13g2_o21ai_1 _1533_ (.B1(_0668_),
    .Y(_0856_),
    .A1(_0786_),
    .A2(_0855_));
 sg13g2_o21ai_1 _1534_ (.B1(net463),
    .Y(_0857_),
    .A1(_0682_),
    .A2(_0790_));
 sg13g2_nand3_1 _1535_ (.B(_0856_),
    .C(_0857_),
    .A(net466),
    .Y(_0858_));
 sg13g2_and2_1 _1536_ (.A(net457),
    .B(_0672_),
    .X(_0859_));
 sg13g2_nor3_1 _1537_ (.A(_0669_),
    .B(_0675_),
    .C(_0859_),
    .Y(_0860_));
 sg13g2_and2_1 _1538_ (.A(_0447_),
    .B(_0674_),
    .X(_0861_));
 sg13g2_or4_1 _1539_ (.A(net466),
    .B(_0786_),
    .C(_0860_),
    .D(_0861_),
    .X(_0862_));
 sg13g2_nand3_1 _1540_ (.B(_0858_),
    .C(_0862_),
    .A(net385),
    .Y(_0863_));
 sg13g2_or2_1 _1541_ (.X(_0864_),
    .B(_0863_),
    .A(net428));
 sg13g2_a22oi_1 _1542_ (.Y(_0865_),
    .B1(_0666_),
    .B2(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[2] ),
    .A2(_0574_),
    .A1(net450));
 sg13g2_nand4_1 _1543_ (.B(_0854_),
    .C(_0864_),
    .A(net352),
    .Y(_0866_),
    .D(_0865_));
 sg13g2_nor2b_1 _1544_ (.A(_0836_),
    .B_N(_0866_),
    .Y(_0104_));
 sg13g2_a21oi_1 _1545_ (.A1(_0605_),
    .A2(_0608_),
    .Y(_0867_),
    .B1(_0607_));
 sg13g2_xnor2_1 _1546_ (.Y(_0868_),
    .A(_0613_),
    .B(_0867_));
 sg13g2_nor2_1 _1547_ (.A(_0766_),
    .B(_0809_),
    .Y(_0869_));
 sg13g2_nor3_1 _1548_ (.A(_0626_),
    .B(_0802_),
    .C(_0803_),
    .Y(_0870_));
 sg13g2_nor3_1 _1549_ (.A(_0636_),
    .B(_0798_),
    .C(_0805_),
    .Y(_0871_));
 sg13g2_nor3_1 _1550_ (.A(_0633_),
    .B(_0799_),
    .C(_0802_),
    .Y(_0872_));
 sg13g2_nor4_1 _1551_ (.A(_0869_),
    .B(_0870_),
    .C(_0871_),
    .D(_0872_),
    .Y(_0873_));
 sg13g2_nor2_1 _1552_ (.A(_0837_),
    .B(_0873_),
    .Y(_0874_));
 sg13g2_a221oi_1 _1553_ (.B2(_0617_),
    .C1(_0874_),
    .B1(_0868_),
    .A1(net427),
    .Y(_0875_),
    .A2(_0620_));
 sg13g2_nor2b_1 _1554_ (.A(_0611_),
    .B_N(_0662_),
    .Y(_0876_));
 sg13g2_a221oi_1 _1555_ (.B2(_0610_),
    .C1(_0876_),
    .B1(_0660_),
    .A1(_0613_),
    .Y(_0877_),
    .A2(_0649_));
 sg13g2_o21ai_1 _1556_ (.B1(_0877_),
    .Y(_0878_),
    .A1(net427),
    .A2(_0652_));
 sg13g2_a22oi_1 _1557_ (.Y(_0879_),
    .B1(_0682_),
    .B2(_0669_),
    .A2(_0675_),
    .A1(_0674_));
 sg13g2_a221oi_1 _1558_ (.B2(net463),
    .C1(_0681_),
    .B1(_0790_),
    .A1(_0455_),
    .Y(_0880_),
    .A2(_0675_));
 sg13g2_nor2_1 _1559_ (.A(net463),
    .B(_0789_),
    .Y(_0881_));
 sg13g2_nor3_1 _1560_ (.A(_0673_),
    .B(_0784_),
    .C(_0881_),
    .Y(_0882_));
 sg13g2_o21ai_1 _1561_ (.B1(_0879_),
    .Y(_0883_),
    .A1(_0880_),
    .A2(_0882_));
 sg13g2_nand2_1 _1562_ (.Y(_0884_),
    .A(net385),
    .B(_0883_));
 sg13g2_nor2_1 _1563_ (.A(_0009_),
    .B(_0653_),
    .Y(_0885_));
 sg13g2_a221oi_1 _1564_ (.B2(net392),
    .C1(_0885_),
    .B1(_0657_),
    .A1(\tiny_shader_top_inst.cur_time[6] ),
    .Y(_0886_),
    .A2(_0586_));
 sg13g2_a22oi_1 _1565_ (.Y(_0887_),
    .B1(_0651_),
    .B2(_0565_),
    .A2(_0585_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.user_i[3] ));
 sg13g2_nand2_1 _1566_ (.Y(_0888_),
    .A(_0886_),
    .B(_0887_));
 sg13g2_nand2_1 _1567_ (.Y(_0889_),
    .A(net447),
    .B(_0574_));
 sg13g2_o21ai_1 _1568_ (.B1(_0889_),
    .Y(_0890_),
    .A1(net428),
    .A2(_0884_));
 sg13g2_nor4_1 _1569_ (.A(_0666_),
    .B(_0878_),
    .C(_0888_),
    .D(_0890_),
    .Y(_0891_));
 sg13g2_and2_1 _1570_ (.A(_0875_),
    .B(_0891_),
    .X(_0892_));
 sg13g2_o21ai_1 _1571_ (.B1(_0762_),
    .Y(_0893_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[3] ),
    .A2(_0667_));
 sg13g2_nand2b_1 _1572_ (.Y(_0894_),
    .B(net292),
    .A_N(_0762_));
 sg13g2_o21ai_1 _1573_ (.B1(_0894_),
    .Y(_0105_),
    .A1(_0892_),
    .A2(_0893_));
 sg13g2_xnor2_1 _1574_ (.Y(_0895_),
    .A(_0571_),
    .B(_0627_));
 sg13g2_o21ai_1 _1575_ (.B1(_0595_),
    .Y(_0896_),
    .A1(_0596_),
    .A2(_0615_));
 sg13g2_xor2_1 _1576_ (.B(_0896_),
    .A(_0895_),
    .X(_0897_));
 sg13g2_o21ai_1 _1577_ (.B1(_0633_),
    .Y(_0898_),
    .A1(_0626_),
    .A2(_0809_));
 sg13g2_nand2_1 _1578_ (.Y(_0899_),
    .A(_0801_),
    .B(_0809_));
 sg13g2_nand2_1 _1579_ (.Y(_0900_),
    .A(_0898_),
    .B(_0899_));
 sg13g2_nor3_1 _1580_ (.A(_0636_),
    .B(_0799_),
    .C(_0802_),
    .Y(_0901_));
 sg13g2_nor2_1 _1581_ (.A(_0624_),
    .B(_0901_),
    .Y(_0902_));
 sg13g2_a221oi_1 _1582_ (.B2(_0902_),
    .C1(_0609_),
    .B1(_0900_),
    .A1(net382),
    .Y(_0903_),
    .A2(_0807_));
 sg13g2_nor3_1 _1583_ (.A(_0576_),
    .B(_0648_),
    .C(_0895_),
    .Y(_0904_));
 sg13g2_nand2_1 _1584_ (.Y(_0905_),
    .A(\tiny_shader_top_inst.shader_execute_inst.user_i[5] ),
    .B(_0585_));
 sg13g2_o21ai_1 _1585_ (.B1(_0905_),
    .Y(_0906_),
    .A1(_0012_),
    .A2(_0653_));
 sg13g2_a22oi_1 _1586_ (.Y(_0907_),
    .B1(_0620_),
    .B2(_0627_),
    .A2(_0586_),
    .A1(_0464_));
 sg13g2_o21ai_1 _1587_ (.B1(_0907_),
    .Y(_0908_),
    .A1(_0627_),
    .A2(_0652_));
 sg13g2_nand2_1 _1588_ (.Y(_0909_),
    .A(_0565_),
    .B(_0657_));
 sg13g2_nand3_1 _1589_ (.B(_0627_),
    .C(_0660_),
    .A(net386),
    .Y(_0910_));
 sg13g2_o21ai_1 _1590_ (.B1(_0662_),
    .Y(_0911_),
    .A1(net386),
    .A2(_0627_));
 sg13g2_nor3_1 _1591_ (.A(_0904_),
    .B(_0906_),
    .C(_0908_),
    .Y(_0912_));
 sg13g2_nand4_1 _1592_ (.B(_0910_),
    .C(_0911_),
    .A(_0909_),
    .Y(_0913_),
    .D(_0912_));
 sg13g2_nand2_1 _1593_ (.Y(_0914_),
    .A(net442),
    .B(_0574_));
 sg13g2_o21ai_1 _1594_ (.B1(net457),
    .Y(_0915_),
    .A1(net460),
    .A2(net458));
 sg13g2_nand2_1 _1595_ (.Y(_0916_),
    .A(_0438_),
    .B(_0785_));
 sg13g2_a21oi_1 _1596_ (.A1(_0915_),
    .A2(_0916_),
    .Y(_0917_),
    .B1(_0827_));
 sg13g2_nand2b_1 _1597_ (.Y(_0918_),
    .B(_0579_),
    .A_N(_0917_));
 sg13g2_o21ai_1 _1598_ (.B1(_0914_),
    .Y(_0919_),
    .A1(net429),
    .A2(_0918_));
 sg13g2_nor4_1 _1599_ (.A(_0666_),
    .B(_0903_),
    .C(_0913_),
    .D(_0919_),
    .Y(_0920_));
 sg13g2_o21ai_1 _1600_ (.B1(_0920_),
    .Y(_0258_),
    .A1(_0618_),
    .A2(_0897_));
 sg13g2_o21ai_1 _1601_ (.B1(_0258_),
    .Y(_0259_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[5] ),
    .A2(_0667_));
 sg13g2_nor2_1 _1602_ (.A(net225),
    .B(net352),
    .Y(_0260_));
 sg13g2_a21oi_1 _1603_ (.A1(net352),
    .A2(_0259_),
    .Y(_0106_),
    .B1(_0260_));
 sg13g2_nor2_1 _1604_ (.A(_0573_),
    .B(_0591_),
    .Y(_0261_));
 sg13g2_nor3_2 _1605_ (.A(_0438_),
    .B(_0439_),
    .C(_0588_),
    .Y(_0262_));
 sg13g2_o21ai_1 _1606_ (.B1(_0261_),
    .Y(_0263_),
    .A1(_0540_),
    .A2(_0262_));
 sg13g2_nand3_1 _1607_ (.B(_0792_),
    .C(_0794_),
    .A(_0782_),
    .Y(_0264_));
 sg13g2_nor2_1 _1608_ (.A(_0263_),
    .B(_0264_),
    .Y(_0265_));
 sg13g2_a21oi_1 _1609_ (.A1(_0446_),
    .A2(_0263_),
    .Y(_0107_),
    .B1(_0265_));
 sg13g2_nand2_1 _1610_ (.Y(_0266_),
    .A(_0589_),
    .B(_0831_));
 sg13g2_nor2_1 _1611_ (.A(_0814_),
    .B(_0266_),
    .Y(_0267_));
 sg13g2_a22oi_1 _1612_ (.Y(_0268_),
    .B1(_0822_),
    .B2(_0267_),
    .A2(_0590_),
    .A1(_0459_));
 sg13g2_mux2_1 _1613_ (.A0(_0268_),
    .A1(net308),
    .S(_0263_),
    .X(_0108_));
 sg13g2_and2_1 _1614_ (.A(_0589_),
    .B(_0863_),
    .X(_0269_));
 sg13g2_a22oi_1 _1615_ (.Y(_0270_),
    .B1(_0854_),
    .B2(_0269_),
    .A2(_0590_),
    .A1(_0460_));
 sg13g2_mux2_1 _1616_ (.A0(_0270_),
    .A1(net310),
    .S(_0263_),
    .X(_0109_));
 sg13g2_nand2_1 _1617_ (.Y(_0271_),
    .A(_0589_),
    .B(_0884_));
 sg13g2_nor3_1 _1618_ (.A(_0878_),
    .B(_0888_),
    .C(_0271_),
    .Y(_0272_));
 sg13g2_a22oi_1 _1619_ (.Y(_0273_),
    .B1(_0875_),
    .B2(_0272_),
    .A2(_0590_),
    .A1(_0462_));
 sg13g2_mux2_1 _1620_ (.A0(_0273_),
    .A1(net312),
    .S(_0263_),
    .X(_0110_));
 sg13g2_a21oi_1 _1621_ (.A1(_0679_),
    .A2(_0685_),
    .Y(_0274_),
    .B1(_0590_));
 sg13g2_and2_1 _1622_ (.A(_0665_),
    .B(_0274_),
    .X(_0275_));
 sg13g2_a22oi_1 _1623_ (.Y(_0276_),
    .B1(_0646_),
    .B2(_0275_),
    .A2(_0590_),
    .A1(_0463_));
 sg13g2_mux2_1 _1624_ (.A0(_0276_),
    .A1(net311),
    .S(_0263_),
    .X(_0111_));
 sg13g2_nand2_1 _1625_ (.Y(_0277_),
    .A(_0589_),
    .B(_0918_));
 sg13g2_nor3_1 _1626_ (.A(_0903_),
    .B(_0913_),
    .C(_0277_),
    .Y(_0278_));
 sg13g2_o21ai_1 _1627_ (.B1(_0278_),
    .Y(_0279_),
    .A1(_0618_),
    .A2(_0897_));
 sg13g2_o21ai_1 _1628_ (.B1(_0279_),
    .Y(_0280_),
    .A1(net344),
    .A2(_0589_));
 sg13g2_nand2_1 _1629_ (.Y(_0281_),
    .A(net244),
    .B(_0263_));
 sg13g2_o21ai_1 _1630_ (.B1(_0281_),
    .Y(_0112_),
    .A1(_0263_),
    .A2(_0280_));
 sg13g2_o21ai_1 _1631_ (.B1(_0261_),
    .Y(_0282_),
    .A1(_0553_),
    .A2(_0262_));
 sg13g2_nor2_1 _1632_ (.A(_0264_),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_a21oi_1 _1633_ (.A1(_0445_),
    .A2(_0282_),
    .Y(_0113_),
    .B1(_0283_));
 sg13g2_mux2_1 _1634_ (.A0(_0268_),
    .A1(net301),
    .S(_0282_),
    .X(_0114_));
 sg13g2_mux2_1 _1635_ (.A0(_0270_),
    .A1(net305),
    .S(_0282_),
    .X(_0115_));
 sg13g2_mux2_1 _1636_ (.A0(_0273_),
    .A1(net313),
    .S(_0282_),
    .X(_0116_));
 sg13g2_mux2_1 _1637_ (.A0(_0276_),
    .A1(net315),
    .S(_0282_),
    .X(_0117_));
 sg13g2_nand2_1 _1638_ (.Y(_0284_),
    .A(net227),
    .B(_0282_));
 sg13g2_o21ai_1 _1639_ (.B1(_0284_),
    .Y(_0118_),
    .A1(_0280_),
    .A2(_0282_));
 sg13g2_nor4_2 _1640_ (.A(net274),
    .B(\tiny_shader_top_inst.x_subpos[1] ),
    .C(net262),
    .Y(_0285_),
    .D(net205));
 sg13g2_and3_1 _1641_ (.X(_0286_),
    .A(_0441_),
    .B(_0506_),
    .C(_0285_));
 sg13g2_mux2_1 _1642_ (.A0(net128),
    .A1(net159),
    .S(net372),
    .X(_0119_));
 sg13g2_mux2_1 _1643_ (.A0(net105),
    .A1(net208),
    .S(net366),
    .X(_0120_));
 sg13g2_mux2_1 _1644_ (.A0(net125),
    .A1(net127),
    .S(net358),
    .X(_0121_));
 sg13g2_mux2_1 _1645_ (.A0(net115),
    .A1(net161),
    .S(net365),
    .X(_0122_));
 sg13g2_mux2_1 _1646_ (.A0(net137),
    .A1(net197),
    .S(net360),
    .X(_0123_));
 sg13g2_mux2_1 _1647_ (.A0(net99),
    .A1(net149),
    .S(net369),
    .X(_0124_));
 sg13g2_nand2_1 _1648_ (.Y(_0287_),
    .A(_0050_),
    .B(net369));
 sg13g2_o21ai_1 _1649_ (.B1(_0287_),
    .Y(_0125_),
    .A1(net31),
    .A2(net370));
 sg13g2_mux2_1 _1650_ (.A0(net123),
    .A1(net150),
    .S(net360),
    .X(_0126_));
 sg13g2_a21oi_1 _1651_ (.A1(net456),
    .A2(net452),
    .Y(_0288_),
    .B1(_0262_));
 sg13g2_nor3_2 _1652_ (.A(_0525_),
    .B(_0591_),
    .C(_0288_),
    .Y(_0289_));
 sg13g2_mux2_1 _1653_ (.A0(net132),
    .A1(_0264_),
    .S(_0289_),
    .X(_0127_));
 sg13g2_mux2_1 _1654_ (.A0(net131),
    .A1(_0268_),
    .S(_0289_),
    .X(_0128_));
 sg13g2_mux2_1 _1655_ (.A0(net133),
    .A1(_0270_),
    .S(_0289_),
    .X(_0129_));
 sg13g2_mux2_1 _1656_ (.A0(net291),
    .A1(_0273_),
    .S(_0289_),
    .X(_0130_));
 sg13g2_mux2_1 _1657_ (.A0(net289),
    .A1(_0276_),
    .S(_0289_),
    .X(_0131_));
 sg13g2_nor2_1 _1658_ (.A(net268),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_a21oi_1 _1659_ (.A1(_0280_),
    .A2(_0289_),
    .Y(_0132_),
    .B1(_0290_));
 sg13g2_mux2_1 _1660_ (.A0(net61),
    .A1(net456),
    .S(net371),
    .X(_0133_));
 sg13g2_mux2_1 _1661_ (.A0(net220),
    .A1(net453),
    .S(net364),
    .X(_0134_));
 sg13g2_mux2_1 _1662_ (.A0(net49),
    .A1(net450),
    .S(net357),
    .X(_0135_));
 sg13g2_mux2_1 _1663_ (.A0(net157),
    .A1(net446),
    .S(net361),
    .X(_0136_));
 sg13g2_nand2_1 _1664_ (.Y(_0291_),
    .A(_0051_),
    .B(net362));
 sg13g2_o21ai_1 _1665_ (.B1(_0291_),
    .Y(_0137_),
    .A1(net43),
    .A2(net362));
 sg13g2_mux2_1 _1666_ (.A0(net170),
    .A1(net443),
    .S(net365),
    .X(_0138_));
 sg13g2_mux2_1 _1667_ (.A0(net179),
    .A1(net441),
    .S(net369),
    .X(_0139_));
 sg13g2_mux2_1 _1668_ (.A0(net173),
    .A1(net439),
    .S(net358),
    .X(_0140_));
 sg13g2_mux2_1 _1669_ (.A0(net159),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[7][0] ),
    .S(net372),
    .X(_0141_));
 sg13g2_mux2_1 _1670_ (.A0(\tiny_shader_top_inst.shader_memory_inst.memory[8][1] ),
    .A1(net183),
    .S(net364),
    .X(_0142_));
 sg13g2_mux2_1 _1671_ (.A0(net127),
    .A1(net166),
    .S(net357),
    .X(_0143_));
 sg13g2_mux2_1 _1672_ (.A0(net161),
    .A1(net196),
    .S(net365),
    .X(_0144_));
 sg13g2_mux2_1 _1673_ (.A0(net197),
    .A1(net167),
    .S(net361),
    .X(_0145_));
 sg13g2_mux2_1 _1674_ (.A0(net149),
    .A1(net153),
    .S(net366),
    .X(_0146_));
 sg13g2_nand2_1 _1675_ (.Y(_0292_),
    .A(_0052_),
    .B(net370));
 sg13g2_o21ai_1 _1676_ (.B1(_0292_),
    .Y(_0147_),
    .A1(net33),
    .A2(net370));
 sg13g2_mux2_1 _1677_ (.A0(net150),
    .A1(net181),
    .S(net360),
    .X(_0148_));
 sg13g2_mux2_1 _1678_ (.A0(net65),
    .A1(_0053_),
    .S(net372),
    .X(_0149_));
 sg13g2_mux2_1 _1679_ (.A0(net231),
    .A1(net220),
    .S(net364),
    .X(_0150_));
 sg13g2_nand2_1 _1680_ (.Y(_0293_),
    .A(_0054_),
    .B(net357));
 sg13g2_o21ai_1 _1681_ (.B1(_0293_),
    .Y(_0151_),
    .A1(net57),
    .A2(net357));
 sg13g2_mux2_1 _1682_ (.A0(net222),
    .A1(net157),
    .S(net361),
    .X(_0152_));
 sg13g2_nand2_1 _1683_ (.Y(_0294_),
    .A(_0055_),
    .B(net368));
 sg13g2_o21ai_1 _1684_ (.B1(_0294_),
    .Y(_0153_),
    .A1(net45),
    .A2(net368));
 sg13g2_mux2_1 _1685_ (.A0(net81),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[1][5] ),
    .S(net365),
    .X(_0154_));
 sg13g2_mux2_1 _1686_ (.A0(net71),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[1][6] ),
    .S(net369),
    .X(_0155_));
 sg13g2_mux2_1 _1687_ (.A0(net230),
    .A1(net173),
    .S(net358),
    .X(_0156_));
 sg13g2_mux2_1 _1688_ (.A0(net187),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[5][0] ),
    .S(net371),
    .X(_0157_));
 sg13g2_mux2_1 _1689_ (.A0(net199),
    .A1(net219),
    .S(net363),
    .X(_0158_));
 sg13g2_mux2_1 _1690_ (.A0(net176),
    .A1(net200),
    .S(net359),
    .X(_0159_));
 sg13g2_mux2_1 _1691_ (.A0(net147),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[5][3] ),
    .S(net363),
    .X(_0160_));
 sg13g2_mux2_1 _1692_ (.A0(net155),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[5][4] ),
    .S(net361),
    .X(_0161_));
 sg13g2_mux2_1 _1693_ (.A0(net168),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[5][5] ),
    .S(net366),
    .X(_0162_));
 sg13g2_mux2_1 _1694_ (.A0(net77),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[5][6] ),
    .S(net371),
    .X(_0163_));
 sg13g2_mux2_1 _1695_ (.A0(net194),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[5][7] ),
    .S(net359),
    .X(_0164_));
 sg13g2_mux2_1 _1696_ (.A0(net185),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[2][0] ),
    .S(net372),
    .X(_0165_));
 sg13g2_mux2_1 _1697_ (.A0(net63),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[2][1] ),
    .S(net364),
    .X(_0166_));
 sg13g2_mux2_1 _1698_ (.A0(net73),
    .A1(_0056_),
    .S(net357),
    .X(_0167_));
 sg13g2_mux2_1 _1699_ (.A0(net51),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[2][3] ),
    .S(net363),
    .X(_0168_));
 sg13g2_nand2_1 _1700_ (.Y(_0295_),
    .A(_0057_),
    .B(net361));
 sg13g2_o21ai_1 _1701_ (.B1(_0295_),
    .Y(_0169_),
    .A1(net39),
    .A2(net360));
 sg13g2_mux2_1 _1702_ (.A0(net55),
    .A1(_0058_),
    .S(net365),
    .X(_0170_));
 sg13g2_mux2_1 _1703_ (.A0(net67),
    .A1(_0059_),
    .S(net369),
    .X(_0171_));
 sg13g2_mux2_1 _1704_ (.A0(net151),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[2][7] ),
    .S(net358),
    .X(_0172_));
 sg13g2_mux2_1 _1705_ (.A0(net207),
    .A1(net185),
    .S(net371),
    .X(_0173_));
 sg13g2_mux2_1 _1706_ (.A0(net59),
    .A1(_0060_),
    .S(net364),
    .X(_0174_));
 sg13g2_mux2_1 _1707_ (.A0(net233),
    .A1(net240),
    .S(net357),
    .X(_0175_));
 sg13g2_nand2_1 _1708_ (.Y(_0296_),
    .A(_0061_),
    .B(net363));
 sg13g2_o21ai_1 _1709_ (.B1(_0296_),
    .Y(_0176_),
    .A1(net37),
    .A2(net363));
 sg13g2_nand2_1 _1710_ (.Y(_0297_),
    .A(_0062_),
    .B(net360));
 sg13g2_o21ai_1 _1711_ (.B1(_0297_),
    .Y(_0177_),
    .A1(net41),
    .A2(net360));
 sg13g2_mux2_1 _1712_ (.A0(net217),
    .A1(net237),
    .S(net366),
    .X(_0178_));
 sg13g2_mux2_1 _1713_ (.A0(\tiny_shader_top_inst.shader_memory_inst.memory[4][6] ),
    .A1(net223),
    .S(net369),
    .X(_0179_));
 sg13g2_mux2_1 _1714_ (.A0(net69),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[3][7] ),
    .S(net358),
    .X(_0180_));
 sg13g2_mux2_1 _1715_ (.A0(net198),
    .A1(net187),
    .S(net371),
    .X(_0181_));
 sg13g2_mux2_1 _1716_ (.A0(net183),
    .A1(net199),
    .S(net363),
    .X(_0182_));
 sg13g2_mux2_1 _1717_ (.A0(net166),
    .A1(net176),
    .S(net357),
    .X(_0183_));
 sg13g2_mux2_1 _1718_ (.A0(net196),
    .A1(net147),
    .S(net363),
    .X(_0184_));
 sg13g2_mux2_1 _1719_ (.A0(net167),
    .A1(net155),
    .S(net361),
    .X(_0185_));
 sg13g2_mux2_1 _1720_ (.A0(net153),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[6][5] ),
    .S(net366),
    .X(_0186_));
 sg13g2_nand2_1 _1721_ (.Y(_0298_),
    .A(_0063_),
    .B(net371));
 sg13g2_o21ai_1 _1722_ (.B1(_0298_),
    .Y(_0187_),
    .A1(net35),
    .A2(net369));
 sg13g2_mux2_1 _1723_ (.A0(net181),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[6][7] ),
    .S(net360),
    .X(_0188_));
 sg13g2_mux2_1 _1724_ (.A0(net189),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[4][0] ),
    .S(net371),
    .X(_0189_));
 sg13g2_mux2_1 _1725_ (.A0(\tiny_shader_top_inst.shader_memory_inst.memory[5][1] ),
    .A1(net177),
    .S(net364),
    .X(_0190_));
 sg13g2_mux2_1 _1726_ (.A0(net200),
    .A1(net233),
    .S(net357),
    .X(_0191_));
 sg13g2_mux2_1 _1727_ (.A0(net89),
    .A1(_0064_),
    .S(net363),
    .X(_0192_));
 sg13g2_mux2_1 _1728_ (.A0(net53),
    .A1(_0065_),
    .S(net360),
    .X(_0193_));
 sg13g2_mux2_1 _1729_ (.A0(\tiny_shader_top_inst.shader_memory_inst.memory[5][5] ),
    .A1(net217),
    .S(net366),
    .X(_0194_));
 sg13g2_mux2_1 _1730_ (.A0(net164),
    .A1(\tiny_shader_top_inst.shader_memory_inst.memory[4][6] ),
    .S(net371),
    .X(_0195_));
 sg13g2_mux2_1 _1731_ (.A0(net75),
    .A1(_0066_),
    .S(net358),
    .X(_0196_));
 sg13g2_nand2b_1 _1732_ (.Y(_0299_),
    .B(net438),
    .A_N(\tiny_shader_top_inst.memory_instr[0] ));
 sg13g2_o21ai_1 _1733_ (.B1(_0299_),
    .Y(_0300_),
    .A1(net456),
    .A2(net438));
 sg13g2_nand2_1 _1734_ (.Y(_0301_),
    .A(net128),
    .B(net372));
 sg13g2_o21ai_1 _1735_ (.B1(_0301_),
    .Y(_0197_),
    .A1(net372),
    .A2(_0300_));
 sg13g2_nand2b_1 _1736_ (.Y(_0302_),
    .B(net437),
    .A_N(\tiny_shader_top_inst.memory_instr[1] ));
 sg13g2_o21ai_1 _1737_ (.B1(_0302_),
    .Y(_0303_),
    .A1(net453),
    .A2(net437));
 sg13g2_nand2_1 _1738_ (.Y(_0304_),
    .A(net105),
    .B(net365));
 sg13g2_o21ai_1 _1739_ (.B1(_0304_),
    .Y(_0198_),
    .A1(net365),
    .A2(_0303_));
 sg13g2_nand2b_1 _1740_ (.Y(_0305_),
    .B(net436),
    .A_N(\tiny_shader_top_inst.memory_instr[2] ));
 sg13g2_o21ai_1 _1741_ (.B1(_0305_),
    .Y(_0306_),
    .A1(net448),
    .A2(net436));
 sg13g2_nand2_1 _1742_ (.Y(_0307_),
    .A(net125),
    .B(net358));
 sg13g2_o21ai_1 _1743_ (.B1(_0307_),
    .Y(_0199_),
    .A1(net358),
    .A2(_0306_));
 sg13g2_nand2b_1 _1744_ (.Y(_0308_),
    .B(net437),
    .A_N(\tiny_shader_top_inst.memory_instr[3] ));
 sg13g2_o21ai_1 _1745_ (.B1(_0308_),
    .Y(_0309_),
    .A1(\tiny_shader_top_inst.instr[3] ),
    .A2(net436));
 sg13g2_nand2_1 _1746_ (.Y(_0310_),
    .A(net115),
    .B(net365));
 sg13g2_o21ai_1 _1747_ (.B1(_0310_),
    .Y(_0200_),
    .A1(net362),
    .A2(_0309_));
 sg13g2_nand2b_1 _1748_ (.Y(_0311_),
    .B(net437),
    .A_N(\tiny_shader_top_inst.memory_instr[4] ));
 sg13g2_o21ai_1 _1749_ (.B1(_0311_),
    .Y(_0312_),
    .A1(net445),
    .A2(net436));
 sg13g2_nand2_1 _1750_ (.Y(_0313_),
    .A(net137),
    .B(net362));
 sg13g2_o21ai_1 _1751_ (.B1(_0313_),
    .Y(_0201_),
    .A1(net362),
    .A2(_0312_));
 sg13g2_nand2b_1 _1752_ (.Y(_0314_),
    .B(net436),
    .A_N(\tiny_shader_top_inst.memory_instr[5] ));
 sg13g2_o21ai_1 _1753_ (.B1(_0314_),
    .Y(_0315_),
    .A1(net443),
    .A2(net437));
 sg13g2_nand2_1 _1754_ (.Y(_0316_),
    .A(net99),
    .B(net369));
 sg13g2_o21ai_1 _1755_ (.B1(_0316_),
    .Y(_0202_),
    .A1(net370),
    .A2(_0315_));
 sg13g2_mux2_1 _1756_ (.A0(net441),
    .A1(\tiny_shader_top_inst.memory_instr[6] ),
    .S(net436),
    .X(_0317_));
 sg13g2_nand2_1 _1757_ (.Y(_0318_),
    .A(net109),
    .B(net370));
 sg13g2_o21ai_1 _1758_ (.B1(_0318_),
    .Y(_0203_),
    .A1(net370),
    .A2(_0317_));
 sg13g2_nand2b_1 _1759_ (.Y(_0319_),
    .B(net436),
    .A_N(\tiny_shader_top_inst.memory_instr[7] ));
 sg13g2_o21ai_1 _1760_ (.B1(_0319_),
    .Y(_0320_),
    .A1(net439),
    .A2(net436));
 sg13g2_nand2_1 _1761_ (.Y(_0321_),
    .A(net123),
    .B(net362));
 sg13g2_o21ai_1 _1762_ (.B1(_0321_),
    .Y(_0204_),
    .A1(net359),
    .A2(_0320_));
 sg13g2_mux2_1 _1763_ (.A0(net242),
    .A1(\tiny_shader_top_inst.memory_instr[0] ),
    .S(net430),
    .X(_0205_));
 sg13g2_mux2_1 _1764_ (.A0(net247),
    .A1(\tiny_shader_top_inst.memory_instr[1] ),
    .S(net430),
    .X(_0206_));
 sg13g2_mux2_1 _1765_ (.A0(net273),
    .A1(net260),
    .S(net430),
    .X(_0207_));
 sg13g2_mux2_1 _1766_ (.A0(net260),
    .A1(\tiny_shader_top_inst.memory_instr[3] ),
    .S(net430),
    .X(_0208_));
 sg13g2_mux2_1 _1767_ (.A0(net286),
    .A1(net257),
    .S(net430),
    .X(_0209_));
 sg13g2_mux2_1 _1768_ (.A0(net257),
    .A1(net214),
    .S(net430),
    .X(_0210_));
 sg13g2_mux2_1 _1769_ (.A0(net214),
    .A1(\tiny_shader_top_inst.memory_instr[6] ),
    .S(net430),
    .X(_0211_));
 sg13g2_mux2_1 _1770_ (.A0(net271),
    .A1(\tiny_shader_top_inst.memory_instr[7] ),
    .S(net430),
    .X(_0212_));
 sg13g2_nand3b_1 _1771_ (.B(_0018_),
    .C(net30),
    .Y(_0322_),
    .A_N(\tiny_shader_top_inst.spi_receiver_inst.spi_sclk_delayed ));
 sg13g2_mux2_1 _1772_ (.A0(\tiny_shader_top_inst.memory_instr[7] ),
    .A1(net255),
    .S(_0322_),
    .X(_0213_));
 sg13g2_and3_2 _1773_ (.X(_0323_),
    .A(\tiny_shader_top_inst.spi_receiver_inst.spi_cnt[2] ),
    .B(net47),
    .C(_0524_));
 sg13g2_mux2_1 _1774_ (.A0(net201),
    .A1(\tiny_shader_top_inst.spi_receiver_inst.spi_mosi_sync ),
    .S(_0323_),
    .X(_0214_));
 sg13g2_mux2_1 _1775_ (.A0(_0068_),
    .A1(net83),
    .S(_0323_),
    .X(_0215_));
 sg13g2_mux2_1 _1776_ (.A0(net203),
    .A1(\tiny_shader_top_inst.memory_instr[1] ),
    .S(_0323_),
    .X(_0216_));
 sg13g2_mux2_1 _1777_ (.A0(_0069_),
    .A1(net93),
    .S(_0323_),
    .X(_0217_));
 sg13g2_mux2_1 _1778_ (.A0(net228),
    .A1(\tiny_shader_top_inst.memory_instr[3] ),
    .S(_0323_),
    .X(_0218_));
 sg13g2_mux2_1 _1779_ (.A0(_0070_),
    .A1(net91),
    .S(_0323_),
    .X(_0219_));
 sg13g2_nor2_1 _1780_ (.A(net87),
    .B(net431),
    .Y(_0324_));
 sg13g2_a21oi_1 _1781_ (.A1(_0427_),
    .A2(net431),
    .Y(_0220_),
    .B1(_0324_));
 sg13g2_xor2_1 _1782_ (.B(_0522_),
    .A(net134),
    .X(_0221_));
 sg13g2_xnor2_1 _1783_ (.Y(_0222_),
    .A(_0440_),
    .B(_0524_));
 sg13g2_nand2_1 _1784_ (.Y(_0325_),
    .A(net249),
    .B(net294));
 sg13g2_nor4_2 _1785_ (.A(net191),
    .B(net238),
    .C(net378),
    .Y(_0326_),
    .D(_0325_));
 sg13g2_nor2_2 _1786_ (.A(\tiny_shader_top_inst.next_frame ),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_nand2_2 _1787_ (.Y(_0328_),
    .A(net354),
    .B(_0326_));
 sg13g2_inv_1 _1788_ (.Y(_0329_),
    .A(_0328_));
 sg13g2_a22oi_1 _1789_ (.Y(_0330_),
    .B1(_0329_),
    .B2(net79),
    .A2(_0327_),
    .A1(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[0] ));
 sg13g2_inv_1 _1790_ (.Y(_0223_),
    .A(net80));
 sg13g2_a21oi_1 _1791_ (.A1(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[0] ),
    .A2(_0326_),
    .Y(_0331_),
    .B1(net295));
 sg13g2_nand2_1 _1792_ (.Y(_0332_),
    .A(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[0] ),
    .B(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[1] ));
 sg13g2_and3_1 _1793_ (.X(_0333_),
    .A(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[0] ),
    .B(net295),
    .C(_0326_));
 sg13g2_nor3_1 _1794_ (.A(\tiny_shader_top_inst.next_frame ),
    .B(net296),
    .C(_0333_),
    .Y(_0224_));
 sg13g2_nand2_1 _1795_ (.Y(_0334_),
    .A(net143),
    .B(_0327_));
 sg13g2_nor2_1 _1796_ (.A(_0008_),
    .B(_0332_),
    .Y(_0335_));
 sg13g2_xnor2_1 _1797_ (.Y(_0336_),
    .A(_0008_),
    .B(_0332_));
 sg13g2_o21ai_1 _1798_ (.B1(_0334_),
    .Y(_0225_),
    .A1(_0328_),
    .A2(_0336_));
 sg13g2_nand2_1 _1799_ (.Y(_0337_),
    .A(net141),
    .B(_0327_));
 sg13g2_xor2_1 _1800_ (.B(_0335_),
    .A(_0009_),
    .X(_0338_));
 sg13g2_o21ai_1 _1801_ (.B1(_0337_),
    .Y(_0226_),
    .A1(_0328_),
    .A2(_0338_));
 sg13g2_nand2_1 _1802_ (.Y(_0339_),
    .A(net111),
    .B(_0327_));
 sg13g2_nand4_1 _1803_ (.B(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[1] ),
    .C(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[2] ),
    .A(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[0] ),
    .Y(_0340_),
    .D(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[3] ));
 sg13g2_nor2_1 _1804_ (.A(_0010_),
    .B(_0340_),
    .Y(_0341_));
 sg13g2_xnor2_1 _1805_ (.Y(_0342_),
    .A(_0010_),
    .B(_0340_));
 sg13g2_o21ai_1 _1806_ (.B1(_0339_),
    .Y(_0227_),
    .A1(_0328_),
    .A2(_0342_));
 sg13g2_nand2_1 _1807_ (.Y(_0343_),
    .A(net103),
    .B(_0327_));
 sg13g2_xor2_1 _1808_ (.B(_0341_),
    .A(_0012_),
    .X(_0344_));
 sg13g2_o21ai_1 _1809_ (.B1(_0343_),
    .Y(_0228_),
    .A1(_0328_),
    .A2(_0344_));
 sg13g2_a21oi_1 _1810_ (.A1(_0506_),
    .A2(_0285_),
    .Y(_0229_),
    .B1(net274));
 sg13g2_xnor2_1 _1811_ (.Y(_0345_),
    .A(net274),
    .B(net324));
 sg13g2_nor2_1 _1812_ (.A(net263),
    .B(_0345_),
    .Y(_0230_));
 sg13g2_nand3_1 _1813_ (.B(net324),
    .C(net262),
    .A(net274),
    .Y(_0346_));
 sg13g2_a21o_1 _1814_ (.A2(net324),
    .A1(net274),
    .B1(net262),
    .X(_0347_));
 sg13g2_and2_1 _1815_ (.A(_0346_),
    .B(_0347_),
    .X(_0231_));
 sg13g2_nor2_1 _1816_ (.A(_0494_),
    .B(_0231_),
    .Y(_0348_));
 sg13g2_a21oi_1 _1817_ (.A1(_0437_),
    .A2(_0346_),
    .Y(_0232_),
    .B1(_0348_));
 sg13g2_and2_1 _1818_ (.A(net307),
    .B(_0000_),
    .X(_0349_));
 sg13g2_nor2_1 _1819_ (.A(net307),
    .B(net263),
    .Y(_0350_));
 sg13g2_nor3_1 _1820_ (.A(net374),
    .B(_0349_),
    .C(_0350_),
    .Y(_0233_));
 sg13g2_o21ai_1 _1821_ (.B1(net378),
    .Y(_0351_),
    .A1(net314),
    .A2(_0349_));
 sg13g2_a21oi_1 _1822_ (.A1(net314),
    .A2(_0349_),
    .Y(_0234_),
    .B1(_0351_));
 sg13g2_and3_1 _1823_ (.X(_0352_),
    .A(net314),
    .B(net252),
    .C(_0349_));
 sg13g2_a21oi_1 _1824_ (.A1(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[1] ),
    .A2(_0349_),
    .Y(_0353_),
    .B1(net252));
 sg13g2_nor3_1 _1825_ (.A(net374),
    .B(_0352_),
    .C(net253),
    .Y(_0235_));
 sg13g2_and2_1 _1826_ (.A(net325),
    .B(_0352_),
    .X(_0354_));
 sg13g2_nor2_1 _1827_ (.A(net325),
    .B(_0352_),
    .Y(_0355_));
 sg13g2_nor3_1 _1828_ (.A(net374),
    .B(_0354_),
    .C(_0355_),
    .Y(_0236_));
 sg13g2_nand2_1 _1829_ (.Y(_0356_),
    .A(net306),
    .B(_0354_));
 sg13g2_o21ai_1 _1830_ (.B1(net378),
    .Y(_0357_),
    .A1(net306),
    .A2(_0354_));
 sg13g2_nor2b_1 _1831_ (.A(_0357_),
    .B_N(_0356_),
    .Y(_0237_));
 sg13g2_xor2_1 _1832_ (.B(_0356_),
    .A(net322),
    .X(_0358_));
 sg13g2_nor2_1 _1833_ (.A(net374),
    .B(_0358_),
    .Y(_0238_));
 sg13g2_and2_1 _1834_ (.A(net375),
    .B(_0485_),
    .X(_0359_));
 sg13g2_xor2_1 _1835_ (.B(_0359_),
    .A(net249),
    .X(_0239_));
 sg13g2_and3_1 _1836_ (.X(_0360_),
    .A(\tiny_shader_top_inst.y_subpos[0] ),
    .B(net191),
    .C(_0359_));
 sg13g2_and2_1 _1837_ (.A(_0485_),
    .B(_0326_),
    .X(_0361_));
 sg13g2_a21oi_1 _1838_ (.A1(\tiny_shader_top_inst.y_subpos[0] ),
    .A2(_0359_),
    .Y(_0362_),
    .B1(net191));
 sg13g2_nor3_1 _1839_ (.A(_0360_),
    .B(_0361_),
    .C(net192),
    .Y(_0240_));
 sg13g2_nand2_1 _1840_ (.Y(_0363_),
    .A(net238),
    .B(_0360_));
 sg13g2_xor2_1 _1841_ (.B(_0360_),
    .A(net238),
    .X(_0241_));
 sg13g2_xor2_1 _1842_ (.B(_0363_),
    .A(net294),
    .X(_0364_));
 sg13g2_nor2_1 _1843_ (.A(_0361_),
    .B(_0364_),
    .Y(_0242_));
 sg13g2_a21oi_1 _1844_ (.A1(\tiny_shader_top_inst.counter_h[6] ),
    .A2(\tiny_shader_top_inst.counter_h[5] ),
    .Y(_0365_),
    .B1(net435));
 sg13g2_or2_1 _1845_ (.X(_0366_),
    .B(_0365_),
    .A(_0516_));
 sg13g2_or3_1 _1846_ (.A(\tiny_shader_top_inst.counter_v[3] ),
    .B(\tiny_shader_top_inst.counter_v[2] ),
    .C(_0487_),
    .X(_0367_));
 sg13g2_a21oi_1 _1847_ (.A1(\tiny_shader_top_inst.counter_v[4] ),
    .A2(_0367_),
    .Y(_0368_),
    .B1(\tiny_shader_top_inst.counter_v[5] ));
 sg13g2_o21ai_1 _1848_ (.B1(_0366_),
    .Y(_0369_),
    .A1(_0513_),
    .A2(_0368_));
 sg13g2_nor2b_1 _1849_ (.A(net433),
    .B_N(net281),
    .Y(_0370_));
 sg13g2_a21oi_1 _1850_ (.A1(net433),
    .A2(net216),
    .Y(_0371_),
    .B1(net282));
 sg13g2_nor2_1 _1851_ (.A(_0369_),
    .B(net283),
    .Y(_0243_));
 sg13g2_nor2b_1 _1852_ (.A(net434),
    .B_N(net265),
    .Y(_0372_));
 sg13g2_a21oi_1 _1853_ (.A1(net433),
    .A2(net232),
    .Y(_0373_),
    .B1(net266));
 sg13g2_nor2_1 _1854_ (.A(_0369_),
    .B(net267),
    .Y(_0244_));
 sg13g2_nor2b_1 _1855_ (.A(net433),
    .B_N(net209),
    .Y(_0374_));
 sg13g2_a21oi_1 _1856_ (.A1(net433),
    .A2(net175),
    .Y(_0375_),
    .B1(net210));
 sg13g2_nor2_1 _1857_ (.A(_0369_),
    .B(net211),
    .Y(_0245_));
 sg13g2_nor2b_1 _1858_ (.A(net434),
    .B_N(net278),
    .Y(_0376_));
 sg13g2_a21oi_1 _1859_ (.A1(net434),
    .A2(net246),
    .Y(_0377_),
    .B1(net279));
 sg13g2_nor2_1 _1860_ (.A(_0369_),
    .B(net280),
    .Y(_0246_));
 sg13g2_nor2b_1 _1861_ (.A(net433),
    .B_N(net234),
    .Y(_0378_));
 sg13g2_a21oi_1 _1862_ (.A1(net433),
    .A2(net172),
    .Y(_0379_),
    .B1(net235));
 sg13g2_nor2_1 _1863_ (.A(_0369_),
    .B(net236),
    .Y(_0247_));
 sg13g2_nor2b_1 _1864_ (.A(net434),
    .B_N(uo_out[0]),
    .Y(_0380_));
 sg13g2_a21oi_1 _1865_ (.A1(net433),
    .A2(net212),
    .Y(_0381_),
    .B1(_0380_));
 sg13g2_nor2_1 _1866_ (.A(_0369_),
    .B(net213),
    .Y(_0248_));
 sg13g2_mux2_1 _1867_ (.A0(\tiny_shader_top_inst.cur_time[0] ),
    .A1(net162),
    .S(\tiny_shader_top_inst.next_frame ),
    .X(_0249_));
 sg13g2_nor2_1 _1868_ (.A(\tiny_shader_top_inst.cur_time[1] ),
    .B(\tiny_shader_top_inst.time_dir ),
    .Y(_0382_));
 sg13g2_xor2_1 _1869_ (.B(\tiny_shader_top_inst.time_dir ),
    .A(\tiny_shader_top_inst.cur_time[1] ),
    .X(_0383_));
 sg13g2_xnor2_1 _1870_ (.Y(_0384_),
    .A(net162),
    .B(_0383_));
 sg13g2_nor2_1 _1871_ (.A(net355),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_a21oi_1 _1872_ (.A1(_0443_),
    .A2(net355),
    .Y(_0250_),
    .B1(_0385_));
 sg13g2_and2_1 _1873_ (.A(net464),
    .B(\tiny_shader_top_inst.cur_time[2] ),
    .X(_0386_));
 sg13g2_nor2_1 _1874_ (.A(\tiny_shader_top_inst.time_dir ),
    .B(\tiny_shader_top_inst.cur_time[2] ),
    .Y(_0387_));
 sg13g2_nor2_1 _1875_ (.A(_0386_),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_a21oi_1 _1876_ (.A1(\tiny_shader_top_inst.cur_time[1] ),
    .A2(net464),
    .Y(_0389_),
    .B1(\tiny_shader_top_inst.cur_time[0] ));
 sg13g2_nor2_1 _1877_ (.A(_0382_),
    .B(_0389_),
    .Y(_0390_));
 sg13g2_nor4_1 _1878_ (.A(_0382_),
    .B(_0386_),
    .C(_0387_),
    .D(_0389_),
    .Y(_0391_));
 sg13g2_xnor2_1 _1879_ (.Y(_0392_),
    .A(_0388_),
    .B(_0390_));
 sg13g2_nand2_1 _1880_ (.Y(_0393_),
    .A(net250),
    .B(net355));
 sg13g2_o21ai_1 _1881_ (.B1(_0393_),
    .Y(_0251_),
    .A1(net355),
    .A2(_0392_));
 sg13g2_nor2_1 _1882_ (.A(_0386_),
    .B(_0391_),
    .Y(_0394_));
 sg13g2_nor2_1 _1883_ (.A(\tiny_shader_top_inst.cur_time[3] ),
    .B(net464),
    .Y(_0395_));
 sg13g2_and2_1 _1884_ (.A(\tiny_shader_top_inst.cur_time[3] ),
    .B(net464),
    .X(_0396_));
 sg13g2_nor2_1 _1885_ (.A(_0395_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_xor2_1 _1886_ (.B(_0397_),
    .A(_0394_),
    .X(_0398_));
 sg13g2_nand2_1 _1887_ (.Y(_0399_),
    .A(net290),
    .B(net354));
 sg13g2_o21ai_1 _1888_ (.B1(_0399_),
    .Y(_0252_),
    .A1(net354),
    .A2(_0398_));
 sg13g2_nand2_1 _1889_ (.Y(_0400_),
    .A(\tiny_shader_top_inst.cur_time[4] ),
    .B(net464));
 sg13g2_xnor2_1 _1890_ (.Y(_0401_),
    .A(\tiny_shader_top_inst.cur_time[4] ),
    .B(net464));
 sg13g2_nor3_1 _1891_ (.A(_0386_),
    .B(_0391_),
    .C(_0396_),
    .Y(_0402_));
 sg13g2_nor2_1 _1892_ (.A(_0395_),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_or3_1 _1893_ (.A(_0395_),
    .B(_0401_),
    .C(_0402_),
    .X(_0404_));
 sg13g2_xor2_1 _1894_ (.B(_0403_),
    .A(_0401_),
    .X(_0405_));
 sg13g2_nand2_1 _1895_ (.Y(_0406_),
    .A(net309),
    .B(net354));
 sg13g2_o21ai_1 _1896_ (.B1(_0406_),
    .Y(_0253_),
    .A1(net354),
    .A2(_0405_));
 sg13g2_xnor2_1 _1897_ (.Y(_0407_),
    .A(\tiny_shader_top_inst.cur_time[5] ),
    .B(net464));
 sg13g2_nand2_1 _1898_ (.Y(_0408_),
    .A(_0400_),
    .B(_0404_));
 sg13g2_xor2_1 _1899_ (.B(_0408_),
    .A(_0407_),
    .X(_0409_));
 sg13g2_nand2_1 _1900_ (.Y(_0410_),
    .A(net304),
    .B(net354));
 sg13g2_o21ai_1 _1901_ (.B1(_0410_),
    .Y(_0254_),
    .A1(net354),
    .A2(_0409_));
 sg13g2_and2_1 _1902_ (.A(\tiny_shader_top_inst.cur_time[6] ),
    .B(net465),
    .X(_0411_));
 sg13g2_xor2_1 _1903_ (.B(net465),
    .A(\tiny_shader_top_inst.cur_time[6] ),
    .X(_0412_));
 sg13g2_o21ai_1 _1904_ (.B1(net464),
    .Y(_0413_),
    .A1(\tiny_shader_top_inst.cur_time[4] ),
    .A2(\tiny_shader_top_inst.cur_time[5] ));
 sg13g2_nor2_1 _1905_ (.A(_0404_),
    .B(_0407_),
    .Y(_0414_));
 sg13g2_o21ai_1 _1906_ (.B1(_0413_),
    .Y(_0415_),
    .A1(_0404_),
    .A2(_0407_));
 sg13g2_a21oi_1 _1907_ (.A1(_0412_),
    .A2(_0415_),
    .Y(_0416_),
    .B1(net354));
 sg13g2_o21ai_1 _1908_ (.B1(_0416_),
    .Y(_0417_),
    .A1(_0412_),
    .A2(_0415_));
 sg13g2_o21ai_1 _1909_ (.B1(_0417_),
    .Y(_0255_),
    .A1(_0461_),
    .A2(\tiny_shader_top_inst.next_frame ));
 sg13g2_xor2_1 _1910_ (.B(net465),
    .A(\tiny_shader_top_inst.cur_time[7] ),
    .X(_0418_));
 sg13g2_a21oi_1 _1911_ (.A1(_0412_),
    .A2(_0415_),
    .Y(_0419_),
    .B1(_0411_));
 sg13g2_xor2_1 _1912_ (.B(_0419_),
    .A(_0418_),
    .X(_0420_));
 sg13g2_nand2_1 _1913_ (.Y(_0421_),
    .A(net323),
    .B(net356));
 sg13g2_o21ai_1 _1914_ (.B1(_0421_),
    .Y(_0256_),
    .A1(net356),
    .A2(_0420_));
 sg13g2_nand3_1 _1915_ (.B(_0414_),
    .C(_0418_),
    .A(_0412_),
    .Y(_0422_));
 sg13g2_o21ai_1 _1916_ (.B1(net465),
    .Y(_0423_),
    .A1(\tiny_shader_top_inst.cur_time[7] ),
    .A2(\tiny_shader_top_inst.cur_time[6] ));
 sg13g2_nand3_1 _1917_ (.B(_0422_),
    .C(_0423_),
    .A(_0413_),
    .Y(_0424_));
 sg13g2_a21oi_1 _1918_ (.A1(net465),
    .A2(_0424_),
    .Y(_0425_),
    .B1(net356));
 sg13g2_o21ai_1 _1919_ (.B1(_0425_),
    .Y(_0426_),
    .A1(net465),
    .A2(_0424_));
 sg13g2_xnor2_1 _1920_ (.Y(_0257_),
    .A(net136),
    .B(_0426_));
 sg13g2_dfrbp_1 _1921_ (.CLK(net25),
    .RESET_B(net16),
    .D(net1),
    .Q_N(_1040_),
    .Q(rst_n_sync));
 sg13g2_dfrbp_1 _1922_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net404),
    .D(_0082_),
    .Q_N(_1039_),
    .Q(\tiny_shader_top_inst.rgb_o[2] ));
 sg13g2_dfrbp_1 _1923_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net404),
    .D(_0083_),
    .Q_N(_1038_),
    .Q(\tiny_shader_top_inst.rgb_o[3] ));
 sg13g2_dfrbp_1 _1924_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net405),
    .D(_0084_),
    .Q_N(_1037_),
    .Q(\tiny_shader_top_inst.rgb_o[4] ));
 sg13g2_dfrbp_1 _1925_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net417),
    .D(_0085_),
    .Q_N(_1036_),
    .Q(\tiny_shader_top_inst.rgb_o[5] ));
 sg13g2_dfrbp_1 _1926_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net398),
    .D(_0086_),
    .Q_N(_0017_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[0][4] ));
 sg13g2_dfrbp_1 _1927_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net401),
    .D(_0087_),
    .Q_N(\tiny_shader_top_inst.counter_v[0] ),
    .Q(_0042_));
 sg13g2_dfrbp_1 _1928_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net401),
    .D(net118),
    .Q_N(\tiny_shader_top_inst.counter_v[1] ),
    .Q(_0043_));
 sg13g2_dfrbp_1 _1929_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net401),
    .D(_0089_),
    .Q_N(_1035_),
    .Q(\tiny_shader_top_inst.counter_v[2] ));
 sg13g2_dfrbp_1 _1930_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net401),
    .D(net259),
    .Q_N(_1034_),
    .Q(\tiny_shader_top_inst.counter_v[3] ));
 sg13g2_dfrbp_1 _1931_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net401),
    .D(net96),
    .Q_N(\tiny_shader_top_inst.counter_v[4] ),
    .Q(_0044_));
 sg13g2_dfrbp_1 _1932_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net400),
    .D(net327),
    .Q_N(_1033_),
    .Q(\tiny_shader_top_inst.counter_v[5] ));
 sg13g2_dfrbp_1 _1933_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net400),
    .D(net122),
    .Q_N(\tiny_shader_top_inst.counter_v[6] ),
    .Q(_0045_));
 sg13g2_dfrbp_1 _1934_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net400),
    .D(net98),
    .Q_N(\tiny_shader_top_inst.counter_v[7] ),
    .Q(_0046_));
 sg13g2_dfrbp_1 _1935_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net400),
    .D(net146),
    .Q_N(\tiny_shader_top_inst.counter_v[8] ),
    .Q(_0047_));
 sg13g2_dfrbp_1 _1936_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net400),
    .D(net114),
    .Q_N(\tiny_shader_top_inst.counter_v[9] ),
    .Q(_0048_));
 sg13g2_dfrbp_1 _1937_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net400),
    .D(net102),
    .Q_N(\tiny_shader_top_inst.counter_v[10] ),
    .Q(_0049_));
 sg13g2_dfrbp_1 _1938_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net418),
    .D(net339),
    .Q_N(_1032_),
    .Q(\tiny_shader_top_inst.time_dir ));
 sg13g2_dfrbp_1 _1939_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net405),
    .D(_0099_),
    .Q_N(_1031_),
    .Q(\tiny_shader_top_inst.rgb_o[0] ));
 sg13g2_dfrbp_1 _1940_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net405),
    .D(_0100_),
    .Q_N(_1030_),
    .Q(\tiny_shader_top_inst.rgb_o[1] ));
 sg13g2_dfrbp_1 _1941_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net405),
    .D(_0101_),
    .Q_N(_0014_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.skip ));
 sg13g2_dfrbp_1 _1942_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net395),
    .D(_0102_),
    .Q_N(_0021_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[0][0] ));
 sg13g2_dfrbp_1 _1943_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net398),
    .D(_0103_),
    .Q_N(_0023_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[0][1] ));
 sg13g2_dfrbp_1 _1944_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net395),
    .D(net342),
    .Q_N(_0024_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[0][2] ));
 sg13g2_dfrbp_1 _1945_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net398),
    .D(net293),
    .Q_N(_0026_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[0][3] ));
 sg13g2_dfrbp_1 _1946_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net398),
    .D(net226),
    .Q_N(_0027_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[0][5] ));
 sg13g2_dfrbp_1 _1947_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net394),
    .D(_0107_),
    .Q_N(_1029_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[1][0] ));
 sg13g2_dfrbp_1 _1948_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net397),
    .D(_0108_),
    .Q_N(_1028_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[1][1] ));
 sg13g2_dfrbp_1 _1949_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net394),
    .D(_0109_),
    .Q_N(_1027_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[1][2] ));
 sg13g2_dfrbp_1 _1950_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net396),
    .D(_0110_),
    .Q_N(_1026_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[1][3] ));
 sg13g2_dfrbp_1 _1951_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net409),
    .D(_0111_),
    .Q_N(_1025_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[1][4] ));
 sg13g2_dfrbp_1 _1952_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net396),
    .D(net245),
    .Q_N(_1024_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[1][5] ));
 sg13g2_dfrbp_1 _1953_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net394),
    .D(_0113_),
    .Q_N(_1023_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[2][0] ));
 sg13g2_dfrbp_1 _1954_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net397),
    .D(_0114_),
    .Q_N(_1022_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[2][1] ));
 sg13g2_dfrbp_1 _1955_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net394),
    .D(_0115_),
    .Q_N(_1021_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[2][2] ));
 sg13g2_dfrbp_1 _1956_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net398),
    .D(_0116_),
    .Q_N(_1020_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[2][3] ));
 sg13g2_dfrbp_1 _1957_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net409),
    .D(_0117_),
    .Q_N(_1019_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[2][4] ));
 sg13g2_dfrbp_1 _1958_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net396),
    .D(_0118_),
    .Q_N(_1018_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[2][5] ));
 sg13g2_dfrbp_1 _1959_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net423),
    .D(_0119_),
    .Q_N(_1017_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[8][0] ));
 sg13g2_dfrbp_1 _1960_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net411),
    .D(_0120_),
    .Q_N(_1016_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[8][1] ));
 sg13g2_dfrbp_1 _1961_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net396),
    .D(_0121_),
    .Q_N(_1015_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[8][2] ));
 sg13g2_dfrbp_1 _1962_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net415),
    .D(_0122_),
    .Q_N(_1014_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[8][3] ));
 sg13g2_dfrbp_1 _1963_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net407),
    .D(_0123_),
    .Q_N(_1013_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[8][4] ));
 sg13g2_dfrbp_1 _1964_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net414),
    .D(_0124_),
    .Q_N(_1012_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[8][5] ));
 sg13g2_dfrbp_1 _1965_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net421),
    .D(net32),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[8][6] ),
    .Q(_0050_));
 sg13g2_dfrbp_1 _1966_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net410),
    .D(_0126_),
    .Q_N(_1011_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[8][7] ));
 sg13g2_dfrbp_1 _1967_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net394),
    .D(_0127_),
    .Q_N(_0020_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[3][0] ));
 sg13g2_dfrbp_1 _1968_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net394),
    .D(_0128_),
    .Q_N(_0022_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[3][1] ));
 sg13g2_dfrbp_1 _1969_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net394),
    .D(_0129_),
    .Q_N(_0025_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[3][2] ));
 sg13g2_dfrbp_1 _1970_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net396),
    .D(_0130_),
    .Q_N(_1010_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[3][3] ));
 sg13g2_dfrbp_1 _1971_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net409),
    .D(_0131_),
    .Q_N(_1009_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[3][4] ));
 sg13g2_dfrbp_1 _1972_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net408),
    .D(_0132_),
    .Q_N(_1008_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.regs[3][5] ));
 sg13g2_dfrbp_1 _1973_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net425),
    .D(net62),
    .Q_N(_1007_),
    .Q(\tiny_shader_top_inst.instr[0] ));
 sg13g2_dfrbp_1 _1974_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net413),
    .D(net221),
    .Q_N(_1006_),
    .Q(\tiny_shader_top_inst.instr[1] ));
 sg13g2_dfrbp_1 _1975_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net397),
    .D(net50),
    .Q_N(_1005_),
    .Q(\tiny_shader_top_inst.instr[2] ));
 sg13g2_dfrbp_1 _1976_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net412),
    .D(net158),
    .Q_N(_1004_),
    .Q(\tiny_shader_top_inst.instr[3] ));
 sg13g2_dfrbp_1 _1977_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net410),
    .D(net44),
    .Q_N(\tiny_shader_top_inst.instr[4] ),
    .Q(_0051_));
 sg13g2_dfrbp_1 _1978_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net415),
    .D(net171),
    .Q_N(_1003_),
    .Q(\tiny_shader_top_inst.instr[5] ));
 sg13g2_dfrbp_1 _1979_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net414),
    .D(net180),
    .Q_N(_1002_),
    .Q(\tiny_shader_top_inst.instr[6] ));
 sg13g2_dfrbp_1 _1980_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net408),
    .D(net174),
    .Q_N(_1001_),
    .Q(\tiny_shader_top_inst.instr[7] ));
 sg13g2_dfrbp_1 _1981_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net423),
    .D(net160),
    .Q_N(_1000_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[7][0] ));
 sg13g2_dfrbp_1 _1982_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net411),
    .D(net184),
    .Q_N(_0999_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[7][1] ));
 sg13g2_dfrbp_1 _1983_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net396),
    .D(_0143_),
    .Q_N(_0998_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[7][2] ));
 sg13g2_dfrbp_1 _1984_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net413),
    .D(_0144_),
    .Q_N(_0997_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[7][3] ));
 sg13g2_dfrbp_1 _1985_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net412),
    .D(_0145_),
    .Q_N(_0996_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[7][4] ));
 sg13g2_dfrbp_1 _1986_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net416),
    .D(_0146_),
    .Q_N(_0995_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[7][5] ));
 sg13g2_dfrbp_1 _1987_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net421),
    .D(net34),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[7][6] ),
    .Q(_0052_));
 sg13g2_dfrbp_1 _1988_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net407),
    .D(_0148_),
    .Q_N(_0994_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[7][7] ));
 sg13g2_dfrbp_1 _1989_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net421),
    .D(net66),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[1][0] ),
    .Q(_0053_));
 sg13g2_dfrbp_1 _1990_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net411),
    .D(_0150_),
    .Q_N(_0993_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[1][1] ));
 sg13g2_dfrbp_1 _1991_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net397),
    .D(net58),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[1][2] ),
    .Q(_0054_));
 sg13g2_dfrbp_1 _1992_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net412),
    .D(_0152_),
    .Q_N(_0992_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[1][3] ));
 sg13g2_dfrbp_1 _1993_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net410),
    .D(net46),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[1][4] ),
    .Q(_0055_));
 sg13g2_dfrbp_1 _1994_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net415),
    .D(net82),
    .Q_N(_0991_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[1][5] ));
 sg13g2_dfrbp_1 _1995_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net421),
    .D(net72),
    .Q_N(_0990_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[1][6] ));
 sg13g2_dfrbp_1 _1996_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net408),
    .D(_0156_),
    .Q_N(_0989_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[1][7] ));
 sg13g2_dfrbp_1 _1997_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net425),
    .D(net188),
    .Q_N(_0988_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[5][0] ));
 sg13g2_dfrbp_1 _1998_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net411),
    .D(_0158_),
    .Q_N(_0987_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[5][1] ));
 sg13g2_dfrbp_1 _1999_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net396),
    .D(_0159_),
    .Q_N(_0986_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[5][2] ));
 sg13g2_dfrbp_1 _2000_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net412),
    .D(net148),
    .Q_N(_0041_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[5][3] ));
 sg13g2_dfrbp_1 _2001_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net407),
    .D(net156),
    .Q_N(_0040_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[5][4] ));
 sg13g2_dfrbp_1 _2002_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net414),
    .D(net169),
    .Q_N(_0985_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[5][5] ));
 sg13g2_dfrbp_1 _2003_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net425),
    .D(net78),
    .Q_N(_0984_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[5][6] ));
 sg13g2_dfrbp_1 _2004_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net408),
    .D(net195),
    .Q_N(_0039_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[5][7] ));
 sg13g2_dfrbp_1 _2005_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net423),
    .D(net186),
    .Q_N(_0038_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[2][0] ));
 sg13g2_dfrbp_1 _2006_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net411),
    .D(net64),
    .Q_N(_0983_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[2][1] ));
 sg13g2_dfrbp_1 _2007_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net397),
    .D(net74),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[2][2] ),
    .Q(_0056_));
 sg13g2_dfrbp_1 _2008_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net412),
    .D(net52),
    .Q_N(_0982_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[2][3] ));
 sg13g2_dfrbp_1 _2009_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net407),
    .D(net40),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[2][4] ),
    .Q(_0057_));
 sg13g2_dfrbp_1 _2010_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net415),
    .D(net56),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[2][5] ),
    .Q(_0058_));
 sg13g2_dfrbp_1 _2011_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net421),
    .D(net68),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[2][6] ),
    .Q(_0059_));
 sg13g2_dfrbp_1 _2012_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net408),
    .D(net152),
    .Q_N(_0981_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[2][7] ));
 sg13g2_dfrbp_1 _2013_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net423),
    .D(_0173_),
    .Q_N(_0980_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[3][0] ));
 sg13g2_dfrbp_1 _2014_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net411),
    .D(net60),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[3][1] ),
    .Q(_0060_));
 sg13g2_dfrbp_1 _2015_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net397),
    .D(_0175_),
    .Q_N(_0037_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[3][2] ));
 sg13g2_dfrbp_1 _2016_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net412),
    .D(net38),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[3][3] ),
    .Q(_0061_));
 sg13g2_dfrbp_1 _2017_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net407),
    .D(net42),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[3][4] ),
    .Q(_0062_));
 sg13g2_dfrbp_1 _2018_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net414),
    .D(_0178_),
    .Q_N(_0036_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[3][5] ));
 sg13g2_dfrbp_1 _2019_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net421),
    .D(net224),
    .Q_N(_0035_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[3][6] ));
 sg13g2_dfrbp_1 _2020_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net408),
    .D(net70),
    .Q_N(_0979_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[3][7] ));
 sg13g2_dfrbp_1 _2021_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net423),
    .D(_0181_),
    .Q_N(_0978_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[6][0] ));
 sg13g2_dfrbp_1 _2022_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net411),
    .D(_0182_),
    .Q_N(_0977_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[6][1] ));
 sg13g2_dfrbp_1 _2023_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net396),
    .D(_0183_),
    .Q_N(_0976_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[6][2] ));
 sg13g2_dfrbp_1 _2024_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net413),
    .D(_0184_),
    .Q_N(_0975_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[6][3] ));
 sg13g2_dfrbp_1 _2025_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net412),
    .D(_0185_),
    .Q_N(_0974_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[6][4] ));
 sg13g2_dfrbp_1 _2026_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net414),
    .D(net154),
    .Q_N(_0973_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[6][5] ));
 sg13g2_dfrbp_1 _2027_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net421),
    .D(net36),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[6][6] ),
    .Q(_0063_));
 sg13g2_dfrbp_1 _2028_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net407),
    .D(net182),
    .Q_N(_0972_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[6][7] ));
 sg13g2_dfrbp_1 _2029_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net423),
    .D(net190),
    .Q_N(_0971_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[4][0] ));
 sg13g2_dfrbp_1 _2030_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net411),
    .D(net178),
    .Q_N(_0034_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[4][1] ));
 sg13g2_dfrbp_1 _2031_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net397),
    .D(_0191_),
    .Q_N(_0970_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[4][2] ));
 sg13g2_dfrbp_1 _2032_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net412),
    .D(net90),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[4][3] ),
    .Q(_0064_));
 sg13g2_dfrbp_1 _2033_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net407),
    .D(net54),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[4][4] ),
    .Q(_0065_));
 sg13g2_dfrbp_1 _2034_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net414),
    .D(net218),
    .Q_N(_0969_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[4][5] ));
 sg13g2_dfrbp_1 _2035_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net425),
    .D(net165),
    .Q_N(_0968_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[4][6] ));
 sg13g2_dfrbp_1 _2036_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net408),
    .D(net76),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[4][7] ),
    .Q(_0066_));
 sg13g2_dfrbp_1 _2037_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net17),
    .D(net30),
    .Q_N(_0967_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.spi_sclk_delayed ));
 sg13g2_dfrbp_1 _2038_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net422),
    .D(net129),
    .Q_N(_0966_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[9][0] ));
 sg13g2_dfrbp_1 _2039_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net414),
    .D(net106),
    .Q_N(_0965_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[9][1] ));
 sg13g2_dfrbp_1 _2040_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net408),
    .D(net126),
    .Q_N(_0964_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[9][2] ));
 sg13g2_dfrbp_1 _2041_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net415),
    .D(net116),
    .Q_N(_0963_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[9][3] ));
 sg13g2_dfrbp_1 _2042_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net410),
    .D(net138),
    .Q_N(_0962_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[9][4] ));
 sg13g2_dfrbp_1 _2043_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net414),
    .D(net100),
    .Q_N(_0961_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[9][5] ));
 sg13g2_dfrbp_1 _2044_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net421),
    .D(net110),
    .Q_N(\tiny_shader_top_inst.shader_memory_inst.memory[9][6] ),
    .Q(_0067_));
 sg13g2_dfrbp_1 _2045_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net407),
    .D(net124),
    .Q_N(_0960_),
    .Q(\tiny_shader_top_inst.shader_memory_inst.memory[9][7] ));
 sg13g2_dfrbp_1 _2046_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net422),
    .D(net243),
    .Q_N(_0033_),
    .Q(\tiny_shader_top_inst.memory_instr[0] ));
 sg13g2_dfrbp_1 _2047_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net422),
    .D(net248),
    .Q_N(_0959_),
    .Q(\tiny_shader_top_inst.memory_instr[1] ));
 sg13g2_dfrbp_1 _2048_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net409),
    .D(_0207_),
    .Q_N(_0032_),
    .Q(\tiny_shader_top_inst.memory_instr[2] ));
 sg13g2_dfrbp_1 _2049_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net409),
    .D(net261),
    .Q_N(_0958_),
    .Q(\tiny_shader_top_inst.memory_instr[3] ));
 sg13g2_dfrbp_1 _2050_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net409),
    .D(_0209_),
    .Q_N(_0031_),
    .Q(\tiny_shader_top_inst.memory_instr[4] ));
 sg13g2_dfrbp_1 _2051_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net415),
    .D(_0210_),
    .Q_N(_0957_),
    .Q(\tiny_shader_top_inst.memory_instr[5] ));
 sg13g2_dfrbp_1 _2052_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net415),
    .D(net215),
    .Q_N(_0956_),
    .Q(\tiny_shader_top_inst.memory_instr[6] ));
 sg13g2_dfrbp_1 _2053_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net422),
    .D(net272),
    .Q_N(_0955_),
    .Q(\tiny_shader_top_inst.memory_instr[7] ));
 sg13g2_dfrbp_1 _2054_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net419),
    .D(net256),
    .Q_N(_0954_),
    .Q(spi_miso));
 sg13g2_dfrbp_1 _2055_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net422),
    .D(net202),
    .Q_N(_0953_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.user_i[0] ));
 sg13g2_dfrbp_1 _2056_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net422),
    .D(net84),
    .Q_N(\tiny_shader_top_inst.shader_execute_inst.user_i[1] ),
    .Q(_0068_));
 sg13g2_dfrbp_1 _2057_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net422),
    .D(net204),
    .Q_N(_0952_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.user_i[2] ));
 sg13g2_dfrbp_1 _2058_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net409),
    .D(net94),
    .Q_N(\tiny_shader_top_inst.shader_execute_inst.user_i[3] ),
    .Q(_0069_));
 sg13g2_dfrbp_1 _2059_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net417),
    .D(net229),
    .Q_N(_0951_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.user_i[4] ));
 sg13g2_dfrbp_1 _2060_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net409),
    .D(net92),
    .Q_N(\tiny_shader_top_inst.shader_execute_inst.user_i[5] ),
    .Q(_0070_));
 sg13g2_dfrbp_1 _2061_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net424),
    .D(net48),
    .Q_N(_1041_),
    .Q(\tiny_shader_top_inst.memory_load ));
 sg13g2_dfrbp_1 _2062_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net418),
    .D(net6),
    .Q_N(_1042_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.synchronizer_spi_mosi.pipe[0] ));
 sg13g2_dfrbp_1 _2063_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net424),
    .D(net26),
    .Q_N(_1043_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.spi_mosi_sync ));
 sg13g2_dfrbp_1 _2064_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net424),
    .D(net5),
    .Q_N(_1044_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.synchronizer_spi_cs.pipe[0] ));
 sg13g2_dfrbp_1 _2065_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net424),
    .D(net27),
    .Q_N(_0018_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.spi_cs_sync ));
 sg13g2_dfrbp_1 _2066_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net418),
    .D(net7),
    .Q_N(_1045_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.synchronizer_spi_sclk.pipe[0] ));
 sg13g2_dfrbp_1 _2067_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net424),
    .D(net28),
    .Q_N(_1046_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.spi_sclk_sync ));
 sg13g2_dfrbp_1 _2068_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net423),
    .D(net2),
    .Q_N(_1047_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.synchronizer_mode.pipe[0] ));
 sg13g2_dfrbp_1 _2069_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net425),
    .D(net29),
    .Q_N(_0019_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.mode_sync ));
 sg13g2_dfrbp_1 _2070_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net424),
    .D(net88),
    .Q_N(_0030_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.spi_cnt[0] ));
 sg13g2_dfrbp_1 _2071_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net423),
    .D(net135),
    .Q_N(_0950_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.spi_cnt[1] ));
 sg13g2_dfrbp_1 _2072_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net424),
    .D(net277),
    .Q_N(_1048_),
    .Q(\tiny_shader_top_inst.spi_receiver_inst.spi_cnt[2] ));
 sg13g2_dfrbp_1 _2073_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net399),
    .D(_0002_),
    .Q_N(_1049_),
    .Q(\tiny_shader_top_inst.counter_h[0] ));
 sg13g2_dfrbp_1 _2074_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net399),
    .D(_0003_),
    .Q_N(_1050_),
    .Q(\tiny_shader_top_inst.counter_h[1] ));
 sg13g2_dfrbp_1 _2075_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net399),
    .D(_0004_),
    .Q_N(_1051_),
    .Q(\tiny_shader_top_inst.counter_h[2] ));
 sg13g2_dfrbp_1 _2076_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net402),
    .D(_0005_),
    .Q_N(_0016_),
    .Q(\tiny_shader_top_inst.counter_h[3] ));
 sg13g2_dfrbp_1 _2077_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net399),
    .D(_0006_),
    .Q_N(_0015_),
    .Q(\tiny_shader_top_inst.counter_h[4] ));
 sg13g2_dfrbp_1 _2078_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net400),
    .D(_0077_),
    .Q_N(\tiny_shader_top_inst.counter_h[5] ),
    .Q(_0071_));
 sg13g2_dfrbp_1 _2079_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net400),
    .D(net321),
    .Q_N(\tiny_shader_top_inst.counter_h[6] ),
    .Q(_0072_));
 sg13g2_dfrbp_1 _2080_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net399),
    .D(_0007_),
    .Q_N(_0013_),
    .Q(\tiny_shader_top_inst.counter_h[7] ));
 sg13g2_dfrbp_1 _2081_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net399),
    .D(_0079_),
    .Q_N(\tiny_shader_top_inst.counter_h[8] ),
    .Q(_0073_));
 sg13g2_dfrbp_1 _2082_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net402),
    .D(_0080_),
    .Q_N(\tiny_shader_top_inst.counter_h[9] ),
    .Q(_0074_));
 sg13g2_dfrbp_1 _2083_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net401),
    .D(net86),
    .Q_N(\tiny_shader_top_inst.counter_h[10] ),
    .Q(_0075_));
 sg13g2_dfrbp_1 _2084_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net417),
    .D(_0223_),
    .Q_N(_0028_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[0] ));
 sg13g2_dfrbp_1 _2085_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net420),
    .D(net297),
    .Q_N(_0949_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[1] ));
 sg13g2_dfrbp_1 _2086_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net420),
    .D(net144),
    .Q_N(_0008_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[2] ));
 sg13g2_dfrbp_1 _2087_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net417),
    .D(net142),
    .Q_N(_0009_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[3] ));
 sg13g2_dfrbp_1 _2088_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net420),
    .D(net112),
    .Q_N(_0010_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[4] ));
 sg13g2_dfrbp_1 _2089_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net417),
    .D(net104),
    .Q_N(_0012_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[5] ));
 sg13g2_dfrbp_1 _2090_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net403),
    .D(net275),
    .Q_N(_0948_),
    .Q(\tiny_shader_top_inst.x_subpos[0] ));
 sg13g2_dfrbp_1 _2091_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net403),
    .D(_0230_),
    .Q_N(_0947_),
    .Q(\tiny_shader_top_inst.x_subpos[1] ));
 sg13g2_dfrbp_1 _2092_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net403),
    .D(_0231_),
    .Q_N(_0946_),
    .Q(\tiny_shader_top_inst.x_subpos[2] ));
 sg13g2_dfrbp_1 _2093_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net403),
    .D(net206),
    .Q_N(_0945_),
    .Q(\tiny_shader_top_inst.x_subpos[3] ));
 sg13g2_dfrbp_1 _2094_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net399),
    .D(_0233_),
    .Q_N(_0944_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[0] ));
 sg13g2_dfrbp_1 _2095_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net399),
    .D(_0234_),
    .Q_N(_0943_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[1] ));
 sg13g2_dfrbp_1 _2096_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net395),
    .D(net254),
    .Q_N(_0942_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[2] ));
 sg13g2_dfrbp_1 _2097_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net395),
    .D(_0236_),
    .Q_N(_0941_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[3] ));
 sg13g2_dfrbp_1 _2098_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net394),
    .D(_0237_),
    .Q_N(_0940_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[4] ));
 sg13g2_dfrbp_1 _2099_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net395),
    .D(_0238_),
    .Q_N(_0939_),
    .Q(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[5] ));
 sg13g2_dfrbp_1 _2100_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net403),
    .D(_0239_),
    .Q_N(_0938_),
    .Q(\tiny_shader_top_inst.y_subpos[0] ));
 sg13g2_dfrbp_1 _2101_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net403),
    .D(net193),
    .Q_N(_0937_),
    .Q(\tiny_shader_top_inst.y_subpos[1] ));
 sg13g2_dfrbp_1 _2102_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net403),
    .D(net239),
    .Q_N(_0936_),
    .Q(\tiny_shader_top_inst.y_subpos[2] ));
 sg13g2_dfrbp_1 _2103_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net403),
    .D(_0242_),
    .Q_N(_0935_),
    .Q(\tiny_shader_top_inst.y_subpos[3] ));
 sg13g2_dfrbp_1 _2104_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net404),
    .D(_0243_),
    .Q_N(_0934_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _2105_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net418),
    .D(_0244_),
    .Q_N(_0933_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _2106_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net404),
    .D(_0245_),
    .Q_N(_0932_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2107_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net418),
    .D(_0246_),
    .Q_N(_0931_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _2108_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net404),
    .D(_0247_),
    .Q_N(_0930_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2109_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net418),
    .D(_0248_),
    .Q_N(_1052_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _2110_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net404),
    .D(net263),
    .Q_N(_0929_),
    .Q(\tiny_shader_top_inst.capture ));
 sg13g2_dfrbp_1 _2111_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net419),
    .D(net163),
    .Q_N(_0029_),
    .Q(\tiny_shader_top_inst.cur_time[0] ));
 sg13g2_dfrbp_1 _2112_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net419),
    .D(net285),
    .Q_N(_0928_),
    .Q(\tiny_shader_top_inst.cur_time[1] ));
 sg13g2_dfrbp_1 _2113_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net419),
    .D(net251),
    .Q_N(_0927_),
    .Q(\tiny_shader_top_inst.cur_time[2] ));
 sg13g2_dfrbp_1 _2114_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net424),
    .D(_0252_),
    .Q_N(_0926_),
    .Q(\tiny_shader_top_inst.cur_time[3] ));
 sg13g2_dfrbp_1 _2115_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net417),
    .D(_0253_),
    .Q_N(_0925_),
    .Q(\tiny_shader_top_inst.cur_time[4] ));
 sg13g2_dfrbp_1 _2116_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net417),
    .D(_0254_),
    .Q_N(_0924_),
    .Q(\tiny_shader_top_inst.cur_time[5] ));
 sg13g2_dfrbp_1 _2117_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net417),
    .D(_0255_),
    .Q_N(_0923_),
    .Q(\tiny_shader_top_inst.cur_time[6] ));
 sg13g2_dfrbp_1 _2118_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net418),
    .D(_0256_),
    .Q_N(_0922_),
    .Q(\tiny_shader_top_inst.cur_time[7] ));
 sg13g2_dfrbp_1 _2119_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net418),
    .D(_0257_),
    .Q_N(_0011_),
    .Q(\tiny_shader_top_inst.cur_time[8] ));
 sg13g2_dfrbp_1 _2120_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net18),
    .D(\tiny_shader_top_inst.next_frame ),
    .Q_N(_1053_),
    .Q(next_frame));
 sg13g2_dfrbp_1 _2121_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net19),
    .D(net376),
    .Q_N(_1054_),
    .Q(next_vertical));
 sg13g2_dfrbp_1 _2122_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net14),
    .D(net336),
    .Q_N(_1055_),
    .Q(\tiny_shader_top_inst.vsync_o ));
 sg13g2_dfrbp_1 _2123_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net15),
    .D(net317),
    .Q_N(_0921_),
    .Q(hsync));
 sg13g2_tiehi _2123__15 (.L_HI(net15));
 sg13g2_tiehi _1921__16 (.L_HI(net16));
 sg13g2_tiehi _2037__17 (.L_HI(net17));
 sg13g2_tiehi _2120__18 (.L_HI(net18));
 sg13g2_tiehi _2121__19 (.L_HI(net19));
 sg13g2_tiehi tt_um_tiny_shader_mole99_20 (.L_HI(net20));
 sg13g2_tiehi tt_um_tiny_shader_mole99_21 (.L_HI(net21));
 sg13g2_tiehi tt_um_tiny_shader_mole99_22 (.L_HI(net22));
 sg13g2_tiehi tt_um_tiny_shader_mole99_23 (.L_HI(net23));
 sg13g2_tiehi tt_um_tiny_shader_mole99_24 (.L_HI(net24));
 sg13g2_inv_1 _1101__1 (.Y(net25),
    .A(clknet_1_0__leaf_clk));
 sg13g2_tielo tt_um_tiny_shader_mole99_9 (.L_LO(net9));
 sg13g2_tielo tt_um_tiny_shader_mole99_10 (.L_LO(net10));
 sg13g2_tielo tt_um_tiny_shader_mole99_11 (.L_LO(net11));
 sg13g2_tielo tt_um_tiny_shader_mole99_12 (.L_LO(net12));
 sg13g2_tielo tt_um_tiny_shader_mole99_13 (.L_LO(net13));
 sg13g2_tiehi _2122__14 (.L_HI(net14));
 sg13g2_buf_1 _2141_ (.A(spi_miso),
    .X(uio_out[2]));
 sg13g2_buf_1 _2142_ (.A(next_vertical),
    .X(uio_out[4]));
 sg13g2_buf_1 _2143_ (.A(next_frame),
    .X(uio_out[5]));
 sg13g2_buf_1 _2144_ (.A(\tiny_shader_top_inst.vsync_o ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2145_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout352 (.A(_0762_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_0691_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(net356),
    .X(net354));
 sg13g2_buf_1 fanout355 (.A(net356),
    .X(net355));
 sg13g2_buf_1 fanout356 (.A(_0493_),
    .X(net356));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(net359));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(net359));
 sg13g2_buf_2 fanout359 (.A(net373),
    .X(net359));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(net362));
 sg13g2_buf_2 fanout361 (.A(net362),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(net368),
    .X(net362));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(net367));
 sg13g2_buf_2 fanout364 (.A(net367),
    .X(net364));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(net367));
 sg13g2_buf_2 fanout366 (.A(net367),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(net368),
    .X(net367));
 sg13g2_buf_1 fanout368 (.A(net373),
    .X(net368));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(net370));
 sg13g2_buf_2 fanout370 (.A(net373),
    .X(net370));
 sg13g2_buf_4 fanout371 (.X(net371),
    .A(net372));
 sg13g2_buf_2 fanout372 (.A(net373),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_0286_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(net376),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(net376),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(\tiny_shader_top_inst.next_vertical ),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(net378),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_0475_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_0628_),
    .X(net379));
 sg13g2_buf_1 fanout380 (.A(_0628_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_0606_),
    .X(net381));
 sg13g2_buf_1 fanout382 (.A(_0606_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_0600_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_0597_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_0579_),
    .X(net385));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(_0571_));
 sg13g2_buf_4 fanout387 (.X(net387),
    .A(_0565_));
 sg13g2_buf_2 fanout388 (.A(net389),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_0555_),
    .X(net389));
 sg13g2_buf_4 fanout390 (.X(net390),
    .A(net391));
 sg13g2_buf_2 fanout391 (.A(_0551_),
    .X(net391));
 sg13g2_buf_4 fanout392 (.X(net392),
    .A(_0545_));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(_0538_));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(net406));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(net406));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(net397));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(net398));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(net406));
 sg13g2_buf_4 fanout399 (.X(net399),
    .A(net402));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(net402));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(net402));
 sg13g2_buf_2 fanout402 (.A(net406),
    .X(net402));
 sg13g2_buf_4 fanout403 (.X(net403),
    .A(net405));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(net405));
 sg13g2_buf_4 fanout405 (.X(net405),
    .A(net406));
 sg13g2_buf_4 fanout406 (.X(net406),
    .A(rst_n_sync));
 sg13g2_buf_4 fanout407 (.X(net407),
    .A(net410));
 sg13g2_buf_4 fanout408 (.X(net408),
    .A(net410));
 sg13g2_buf_4 fanout409 (.X(net409),
    .A(net410));
 sg13g2_buf_4 fanout410 (.X(net410),
    .A(net426));
 sg13g2_buf_4 fanout411 (.X(net411),
    .A(net413));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(net416));
 sg13g2_buf_2 fanout413 (.A(net416),
    .X(net413));
 sg13g2_buf_4 fanout414 (.X(net414),
    .A(net415));
 sg13g2_buf_4 fanout415 (.X(net415),
    .A(net416));
 sg13g2_buf_2 fanout416 (.A(net426),
    .X(net416));
 sg13g2_buf_4 fanout417 (.X(net417),
    .A(net420));
 sg13g2_buf_4 fanout418 (.X(net418),
    .A(net420));
 sg13g2_buf_2 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(net426),
    .X(net420));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(net422));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(net425));
 sg13g2_buf_4 fanout423 (.X(net423),
    .A(net425));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(net425));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(net426));
 sg13g2_buf_2 fanout426 (.A(rst_n_sync),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_0609_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_0536_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_0536_),
    .X(net429));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(_0521_));
 sg13g2_buf_1 fanout431 (.A(_0521_),
    .X(net431));
 sg13g2_buf_4 fanout432 (.X(net432),
    .A(_0433_));
 sg13g2_buf_2 fanout433 (.A(\tiny_shader_top_inst.capture ),
    .X(net433));
 sg13g2_buf_1 fanout434 (.A(\tiny_shader_top_inst.capture ),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(\tiny_shader_top_inst.counter_h[7] ),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(net438),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(net438),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(\tiny_shader_top_inst.memory_load ),
    .X(net438));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(\tiny_shader_top_inst.instr[7] ));
 sg13g2_buf_2 fanout440 (.A(net441),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(\tiny_shader_top_inst.instr[6] ),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_1 fanout443 (.A(\tiny_shader_top_inst.instr[5] ),
    .X(net443));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(net445));
 sg13g2_buf_1 fanout445 (.A(\tiny_shader_top_inst.instr[4] ),
    .X(net445));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(\tiny_shader_top_inst.instr[3] ));
 sg13g2_buf_4 fanout447 (.X(net447),
    .A(\tiny_shader_top_inst.instr[3] ));
 sg13g2_buf_4 fanout448 (.X(net448),
    .A(net449));
 sg13g2_buf_2 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_4 fanout450 (.X(net450),
    .A(\tiny_shader_top_inst.instr[2] ));
 sg13g2_buf_2 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(net453),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(\tiny_shader_top_inst.instr[1] ),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(net455),
    .X(net454));
 sg13g2_buf_4 fanout455 (.X(net455),
    .A(net456));
 sg13g2_buf_2 fanout456 (.A(\tiny_shader_top_inst.instr[0] ),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[0][3] ),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(net341),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(net460),
    .X(net459));
 sg13g2_buf_1 fanout460 (.A(net461),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(net328),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(net343),
    .X(net462));
 sg13g2_buf_1 fanout463 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[0][0] ),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(net465),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(\tiny_shader_top_inst.time_dir ),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(net340),
    .X(net466));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[0]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[1]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[3]),
    .X(net7));
 sg13g2_tielo tt_um_tiny_shader_mole99_8 (.L_LO(net8));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_leaf_0_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_1_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_2_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_3_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_4_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_5_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_6_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_7_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_8_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_9_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_10_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_11_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_12_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_13_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_14_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_15_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_16_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_17_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_18_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_19_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_20_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_21_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_22_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_23_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_24_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_25_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_26_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_27_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_28_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_3_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_4__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_5__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_6__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_3_7__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_7__leaf_clk_regs));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk_regs));
 sg13g2_buf_2 clkload1 (.A(clknet_3_5__leaf_clk_regs));
 sg13g2_buf_2 clkload2 (.A(clknet_3_7__leaf_clk_regs));
 sg13g2_inv_4 clkload3 (.A(clknet_leaf_0_clk_regs));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_2_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_27_clk_regs));
 sg13g2_inv_8 clkload6 (.A(clknet_leaf_1_clk_regs));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_25_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_4_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_5_clk_regs));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_6_clk_regs));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_10_clk_regs));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_21_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\tiny_shader_top_inst.spi_receiver_inst.synchronizer_spi_mosi.pipe[0] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold2 (.A(\tiny_shader_top_inst.spi_receiver_inst.synchronizer_spi_cs.pipe[0] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold3 (.A(\tiny_shader_top_inst.spi_receiver_inst.synchronizer_spi_sclk.pipe[0] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold4 (.A(\tiny_shader_top_inst.spi_receiver_inst.synchronizer_mode.pipe[0] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold5 (.A(\tiny_shader_top_inst.spi_receiver_inst.spi_sclk_sync ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold6 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[9][6] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0125_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold8 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[8][6] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0147_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold10 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[7][6] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0187_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold12 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[4][3] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0176_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold14 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[3][4] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0169_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold16 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[4][4] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0177_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold18 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[1][4] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0137_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold20 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[2][4] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0153_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0019_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0001_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold24 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[1][2] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0135_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold26 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[3][3] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0168_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0040_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0193_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0036_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0170_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold32 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[2][2] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0151_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0034_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0174_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold36 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[1][0] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0133_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold38 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[3][1] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0166_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0038_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0149_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0035_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0171_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold44 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[4][7] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0180_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold46 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[2][6] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0155_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0037_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0167_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0039_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0196_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold52 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[6][6] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0163_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0028_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0330_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold56 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[2][5] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0154_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0033_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0215_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold60 (.A(\tiny_shader_top_inst.counter_h[10] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0081_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0030_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0220_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0041_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0192_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0031_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0219_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0032_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0217_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0044_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0091_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0046_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0094_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold74 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[9][5] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0202_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0049_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0097_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold78 (.A(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[5] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0228_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold80 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[9][1] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0198_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0016_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0510_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0067_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0203_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold86 (.A(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[4] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0227_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0048_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0096_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold90 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[9][3] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0200_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0043_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0088_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold94 (.A(\tiny_shader_top_inst.counter_v[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0693_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0045_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0093_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold98 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[9][7] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0204_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold100 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[9][2] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0199_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold102 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[8][2] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold103 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[9][0] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0197_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold105 (.A(\tiny_shader_top_inst.counter_h[0] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold106 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[3][1] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold107 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[3][0] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold108 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[3][2] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold109 (.A(\tiny_shader_top_inst.spi_receiver_inst.spi_cnt[1] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0221_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold111 (.A(\tiny_shader_top_inst.cur_time[8] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold112 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[9][4] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0201_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0015_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0511_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold116 (.A(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[3] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0226_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold118 (.A(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[2] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0225_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0047_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0095_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold122 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[6][3] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0160_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold124 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[8][5] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold125 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[8][7] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold126 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[3][7] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0172_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold128 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[7][5] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0186_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold130 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[6][4] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0161_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold132 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[1][3] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0136_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold134 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[8][0] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0141_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold136 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[8][3] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0029_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0249_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold139 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[5][6] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0195_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold141 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[7][2] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold142 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[7][4] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold143 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[6][5] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0162_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold145 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[1][5] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0138_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold147 (.A(\tiny_shader_top_inst.rgb_o[4] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold148 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[1][7] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0140_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold150 (.A(\tiny_shader_top_inst.rgb_o[2] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold151 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[6][2] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold152 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[4][1] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0190_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold154 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[1][6] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0139_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold156 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[7][7] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0188_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold158 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[7][1] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0142_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold160 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[3][0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0165_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold162 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[6][0] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0157_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold164 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[5][0] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0189_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold166 (.A(\tiny_shader_top_inst.y_subpos[1] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0362_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0240_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold169 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[6][7] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0164_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold171 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[7][3] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold172 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[8][4] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold173 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[7][0] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold174 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[6][1] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold175 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[5][2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold176 (.A(\tiny_shader_top_inst.shader_execute_inst.user_i[0] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0214_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold178 (.A(\tiny_shader_top_inst.shader_execute_inst.user_i[2] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0216_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold180 (.A(\tiny_shader_top_inst.x_subpos[3] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0232_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold182 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[4][0] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold183 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[8][1] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold184 (.A(uo_out[5]),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0374_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0375_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold187 (.A(\tiny_shader_top_inst.rgb_o[5] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0381_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold189 (.A(\tiny_shader_top_inst.memory_instr[5] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0211_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold191 (.A(\tiny_shader_top_inst.rgb_o[0] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold192 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[4][5] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0194_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold194 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[5][1] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold195 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[1][1] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0134_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold197 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[2][3] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold198 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[3][6] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0179_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold200 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[0][5] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0106_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold202 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[2][5] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold203 (.A(\tiny_shader_top_inst.shader_execute_inst.user_i[4] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0218_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold205 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[2][7] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold206 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[2][1] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold207 (.A(\tiny_shader_top_inst.rgb_o[1] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold208 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[4][2] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold209 (.A(uo_out[4]),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0378_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0379_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold212 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[3][5] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold213 (.A(\tiny_shader_top_inst.y_subpos[2] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0241_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold215 (.A(\tiny_shader_top_inst.shader_memory_inst.memory[3][2] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold216 (.A(\tiny_shader_top_inst.shader_execute_inst.skip ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold217 (.A(\tiny_shader_top_inst.spi_receiver_inst.spi_mosi_sync ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0205_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold219 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[1][5] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0112_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold221 (.A(\tiny_shader_top_inst.rgb_o[3] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold222 (.A(\tiny_shader_top_inst.memory_instr[0] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0206_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold224 (.A(\tiny_shader_top_inst.y_subpos[0] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold225 (.A(\tiny_shader_top_inst.cur_time[2] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0251_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold227 (.A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[2] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0353_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0235_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold230 (.A(spi_miso),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0213_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold232 (.A(\tiny_shader_top_inst.memory_instr[4] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold233 (.A(\tiny_shader_top_inst.counter_v[3] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0090_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold235 (.A(\tiny_shader_top_inst.memory_instr[2] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0208_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold237 (.A(\tiny_shader_top_inst.x_subpos[2] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0000_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold239 (.A(\tiny_shader_top_inst.counter_h[1] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold240 (.A(uo_out[2]),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0372_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0373_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold243 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[3][5] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0013_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0512_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold246 (.A(\tiny_shader_top_inst.memory_instr[6] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0212_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold248 (.A(\tiny_shader_top_inst.memory_instr[1] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold249 (.A(\tiny_shader_top_inst.x_subpos[0] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0229_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold251 (.A(\tiny_shader_top_inst.spi_receiver_inst.spi_cnt[2] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0222_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold253 (.A(uo_out[1]),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0376_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0377_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold256 (.A(uo_out[6]),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0370_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0371_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold259 (.A(\tiny_shader_top_inst.cur_time[1] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0250_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold261 (.A(\tiny_shader_top_inst.memory_instr[3] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold262 (.A(\tiny_shader_top_inst.counter_v[2] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0697_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold264 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[3][4] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold265 (.A(\tiny_shader_top_inst.cur_time[3] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold266 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[3][3] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold267 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[0][3] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0105_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold269 (.A(\tiny_shader_top_inst.y_subpos[3] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold270 (.A(\tiny_shader_top_inst.shader_execute_inst.y_pos_i[1] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0331_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0224_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold273 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[1][0] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold274 (.A(\tiny_shader_top_inst.counter_h[5] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0482_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold276 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[2][1] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold277 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[2][0] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold278 (.A(\tiny_shader_top_inst.counter_h[2] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold279 (.A(\tiny_shader_top_inst.cur_time[5] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold280 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[2][2] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold281 (.A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[4] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold282 (.A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[0] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold283 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[1][1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold284 (.A(\tiny_shader_top_inst.cur_time[4] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold285 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[1][2] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold286 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[1][4] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold287 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[1][3] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold288 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[2][3] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold289 (.A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[1] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold290 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[2][4] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold291 (.A(\tiny_shader_top_inst.counter_h[6] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold292 (.A(\tiny_shader_top_inst.hsync ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0014_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold294 (.A(\tiny_shader_top_inst.counter_h[4] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0480_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0078_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold297 (.A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[5] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold298 (.A(\tiny_shader_top_inst.cur_time[7] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold299 (.A(\tiny_shader_top_inst.x_subpos[1] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold300 (.A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[3] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold301 (.A(\tiny_shader_top_inst.counter_v[5] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0092_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold303 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[0][1] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold304 (.A(\tiny_shader_top_inst.counter_h[8] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0476_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold306 (.A(\tiny_shader_top_inst.cur_time[6] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold307 (.A(\tiny_shader_top_inst.counter_h[9] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0477_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold309 (.A(\tiny_shader_top_inst.counter_v[4] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0515_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold311 (.A(\tiny_shader_top_inst.timing_ver.sync ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0011_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0719_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0098_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold315 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[0][4] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold316 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[0][2] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0104_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold318 (.A(\tiny_shader_top_inst.shader_execute_inst.regs[0][0] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold319 (.A(\tiny_shader_top_inst.shader_execute_inst.x_pos_i[5] ),
    .X(net344));
 sg13g2_antennanp ANTENNA_1 (.A(net5));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_fill_2 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_4 FILLER_0_171 ();
 sg13g2_fill_1 FILLER_0_175 ();
 sg13g2_fill_1 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_333 ();
 sg13g2_fill_2 FILLER_0_340 ();
 sg13g2_fill_1 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_354 ();
 sg13g2_fill_2 FILLER_0_361 ();
 sg13g2_fill_1 FILLER_0_390 ();
 sg13g2_decap_4 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_4 FILLER_1_91 ();
 sg13g2_decap_4 FILLER_1_184 ();
 sg13g2_fill_2 FILLER_1_188 ();
 sg13g2_decap_4 FILLER_1_252 ();
 sg13g2_fill_2 FILLER_1_338 ();
 sg13g2_fill_2 FILLER_1_344 ();
 sg13g2_fill_2 FILLER_1_375 ();
 sg13g2_fill_1 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_4 FILLER_2_91 ();
 sg13g2_fill_2 FILLER_2_95 ();
 sg13g2_fill_1 FILLER_2_143 ();
 sg13g2_fill_2 FILLER_2_158 ();
 sg13g2_fill_1 FILLER_2_160 ();
 sg13g2_fill_2 FILLER_2_269 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_fill_1 FILLER_3_98 ();
 sg13g2_fill_2 FILLER_3_219 ();
 sg13g2_fill_1 FILLER_3_221 ();
 sg13g2_fill_2 FILLER_3_246 ();
 sg13g2_fill_1 FILLER_3_284 ();
 sg13g2_fill_2 FILLER_3_305 ();
 sg13g2_fill_1 FILLER_3_358 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_fill_2 FILLER_4_70 ();
 sg13g2_fill_1 FILLER_4_72 ();
 sg13g2_decap_8 FILLER_4_83 ();
 sg13g2_fill_1 FILLER_4_90 ();
 sg13g2_fill_2 FILLER_4_119 ();
 sg13g2_fill_1 FILLER_4_139 ();
 sg13g2_decap_8 FILLER_4_150 ();
 sg13g2_fill_2 FILLER_4_175 ();
 sg13g2_fill_2 FILLER_4_203 ();
 sg13g2_fill_2 FILLER_4_266 ();
 sg13g2_fill_1 FILLER_4_268 ();
 sg13g2_fill_2 FILLER_4_349 ();
 sg13g2_fill_1 FILLER_4_351 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_fill_2 FILLER_5_49 ();
 sg13g2_fill_2 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_fill_2 FILLER_5_112 ();
 sg13g2_fill_1 FILLER_5_145 ();
 sg13g2_fill_2 FILLER_5_206 ();
 sg13g2_fill_2 FILLER_5_213 ();
 sg13g2_fill_1 FILLER_5_215 ();
 sg13g2_fill_1 FILLER_5_243 ();
 sg13g2_fill_2 FILLER_5_280 ();
 sg13g2_fill_1 FILLER_5_282 ();
 sg13g2_fill_1 FILLER_5_346 ();
 sg13g2_fill_2 FILLER_5_366 ();
 sg13g2_fill_1 FILLER_5_378 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_4 FILLER_6_35 ();
 sg13g2_fill_2 FILLER_6_39 ();
 sg13g2_decap_4 FILLER_6_45 ();
 sg13g2_fill_1 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_decap_8 FILLER_6_80 ();
 sg13g2_fill_1 FILLER_6_178 ();
 sg13g2_fill_1 FILLER_6_259 ();
 sg13g2_fill_1 FILLER_6_283 ();
 sg13g2_fill_2 FILLER_6_302 ();
 sg13g2_fill_1 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_fill_2 FILLER_7_21 ();
 sg13g2_fill_1 FILLER_7_23 ();
 sg13g2_fill_1 FILLER_7_60 ();
 sg13g2_fill_2 FILLER_7_70 ();
 sg13g2_fill_1 FILLER_7_98 ();
 sg13g2_fill_2 FILLER_7_104 ();
 sg13g2_fill_2 FILLER_7_148 ();
 sg13g2_fill_2 FILLER_7_228 ();
 sg13g2_fill_1 FILLER_7_277 ();
 sg13g2_fill_1 FILLER_7_309 ();
 sg13g2_fill_1 FILLER_7_338 ();
 sg13g2_fill_1 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_4 FILLER_8_21 ();
 sg13g2_fill_1 FILLER_8_25 ();
 sg13g2_decap_4 FILLER_8_80 ();
 sg13g2_fill_2 FILLER_8_84 ();
 sg13g2_fill_2 FILLER_8_159 ();
 sg13g2_fill_2 FILLER_8_184 ();
 sg13g2_fill_1 FILLER_8_225 ();
 sg13g2_fill_2 FILLER_8_236 ();
 sg13g2_fill_1 FILLER_8_238 ();
 sg13g2_fill_2 FILLER_8_291 ();
 sg13g2_fill_1 FILLER_8_293 ();
 sg13g2_fill_1 FILLER_8_389 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_64 ();
 sg13g2_fill_1 FILLER_9_66 ();
 sg13g2_fill_2 FILLER_9_109 ();
 sg13g2_fill_2 FILLER_9_147 ();
 sg13g2_fill_2 FILLER_9_182 ();
 sg13g2_fill_2 FILLER_9_209 ();
 sg13g2_fill_1 FILLER_9_226 ();
 sg13g2_fill_1 FILLER_9_237 ();
 sg13g2_fill_2 FILLER_9_264 ();
 sg13g2_fill_1 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_23 ();
 sg13g2_fill_1 FILLER_10_27 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_fill_2 FILLER_10_91 ();
 sg13g2_fill_1 FILLER_10_93 ();
 sg13g2_decap_8 FILLER_10_100 ();
 sg13g2_decap_8 FILLER_10_107 ();
 sg13g2_decap_8 FILLER_10_117 ();
 sg13g2_decap_8 FILLER_10_124 ();
 sg13g2_decap_8 FILLER_10_131 ();
 sg13g2_fill_2 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_fill_1 FILLER_10_218 ();
 sg13g2_fill_2 FILLER_10_234 ();
 sg13g2_fill_2 FILLER_10_275 ();
 sg13g2_fill_1 FILLER_10_277 ();
 sg13g2_fill_1 FILLER_10_287 ();
 sg13g2_fill_1 FILLER_10_333 ();
 sg13g2_fill_2 FILLER_10_342 ();
 sg13g2_fill_1 FILLER_10_352 ();
 sg13g2_fill_1 FILLER_10_362 ();
 sg13g2_fill_1 FILLER_10_377 ();
 sg13g2_fill_1 FILLER_10_387 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_68 ();
 sg13g2_fill_2 FILLER_11_75 ();
 sg13g2_fill_2 FILLER_11_96 ();
 sg13g2_fill_1 FILLER_11_98 ();
 sg13g2_fill_1 FILLER_11_117 ();
 sg13g2_decap_8 FILLER_11_122 ();
 sg13g2_fill_2 FILLER_11_129 ();
 sg13g2_fill_2 FILLER_11_147 ();
 sg13g2_fill_1 FILLER_11_149 ();
 sg13g2_decap_8 FILLER_11_155 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_176 ();
 sg13g2_fill_2 FILLER_11_187 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_fill_1 FILLER_11_214 ();
 sg13g2_fill_2 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_266 ();
 sg13g2_fill_1 FILLER_11_268 ();
 sg13g2_fill_2 FILLER_11_304 ();
 sg13g2_fill_1 FILLER_11_306 ();
 sg13g2_fill_2 FILLER_11_380 ();
 sg13g2_fill_1 FILLER_11_382 ();
 sg13g2_fill_1 FILLER_12_44 ();
 sg13g2_fill_1 FILLER_12_49 ();
 sg13g2_fill_1 FILLER_12_54 ();
 sg13g2_decap_4 FILLER_12_59 ();
 sg13g2_fill_2 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_fill_2 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_87 ();
 sg13g2_decap_8 FILLER_12_92 ();
 sg13g2_decap_4 FILLER_12_99 ();
 sg13g2_fill_2 FILLER_12_135 ();
 sg13g2_fill_1 FILLER_12_173 ();
 sg13g2_decap_4 FILLER_12_218 ();
 sg13g2_fill_1 FILLER_12_234 ();
 sg13g2_fill_1 FILLER_12_370 ();
 sg13g2_fill_2 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_30 ();
 sg13g2_fill_2 FILLER_13_39 ();
 sg13g2_fill_2 FILLER_13_108 ();
 sg13g2_decap_4 FILLER_13_115 ();
 sg13g2_decap_4 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_150 ();
 sg13g2_fill_2 FILLER_13_156 ();
 sg13g2_fill_1 FILLER_13_185 ();
 sg13g2_fill_1 FILLER_13_200 ();
 sg13g2_fill_2 FILLER_13_209 ();
 sg13g2_fill_1 FILLER_13_222 ();
 sg13g2_fill_2 FILLER_13_244 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_2 FILLER_13_255 ();
 sg13g2_fill_1 FILLER_13_314 ();
 sg13g2_fill_2 FILLER_13_342 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_47 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_80 ();
 sg13g2_fill_2 FILLER_14_107 ();
 sg13g2_fill_1 FILLER_14_109 ();
 sg13g2_fill_2 FILLER_14_141 ();
 sg13g2_fill_2 FILLER_14_173 ();
 sg13g2_fill_2 FILLER_14_223 ();
 sg13g2_fill_1 FILLER_14_239 ();
 sg13g2_fill_2 FILLER_14_266 ();
 sg13g2_fill_1 FILLER_14_268 ();
 sg13g2_fill_1 FILLER_14_292 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_fill_1 FILLER_15_68 ();
 sg13g2_fill_2 FILLER_15_94 ();
 sg13g2_fill_1 FILLER_15_96 ();
 sg13g2_fill_1 FILLER_15_114 ();
 sg13g2_decap_4 FILLER_15_120 ();
 sg13g2_fill_2 FILLER_15_171 ();
 sg13g2_fill_1 FILLER_15_180 ();
 sg13g2_fill_1 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_225 ();
 sg13g2_fill_2 FILLER_15_267 ();
 sg13g2_fill_1 FILLER_15_314 ();
 sg13g2_fill_2 FILLER_15_344 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_1 FILLER_16_26 ();
 sg13g2_fill_2 FILLER_16_97 ();
 sg13g2_decap_4 FILLER_16_124 ();
 sg13g2_fill_2 FILLER_16_179 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_fill_2 FILLER_16_187 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_fill_2 FILLER_16_196 ();
 sg13g2_fill_1 FILLER_16_198 ();
 sg13g2_fill_2 FILLER_16_243 ();
 sg13g2_fill_2 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_1 FILLER_17_54 ();
 sg13g2_fill_2 FILLER_17_77 ();
 sg13g2_fill_1 FILLER_17_90 ();
 sg13g2_fill_2 FILLER_17_95 ();
 sg13g2_fill_2 FILLER_17_102 ();
 sg13g2_fill_1 FILLER_17_104 ();
 sg13g2_fill_1 FILLER_17_109 ();
 sg13g2_fill_2 FILLER_17_134 ();
 sg13g2_fill_1 FILLER_17_145 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_4 FILLER_17_174 ();
 sg13g2_fill_2 FILLER_17_208 ();
 sg13g2_fill_2 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_221 ();
 sg13g2_fill_1 FILLER_17_256 ();
 sg13g2_fill_2 FILLER_17_262 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_fill_1 FILLER_17_278 ();
 sg13g2_fill_2 FILLER_17_393 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_55 ();
 sg13g2_fill_2 FILLER_18_65 ();
 sg13g2_fill_2 FILLER_18_72 ();
 sg13g2_fill_2 FILLER_18_79 ();
 sg13g2_fill_1 FILLER_18_90 ();
 sg13g2_fill_2 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_107 ();
 sg13g2_fill_1 FILLER_18_145 ();
 sg13g2_fill_2 FILLER_18_161 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_fill_2 FILLER_18_197 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_fill_2 FILLER_18_217 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_fill_1 FILLER_18_235 ();
 sg13g2_fill_1 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_284 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_380 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_fill_1 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_74 ();
 sg13g2_fill_2 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_101 ();
 sg13g2_fill_1 FILLER_19_103 ();
 sg13g2_fill_1 FILLER_19_121 ();
 sg13g2_fill_2 FILLER_19_132 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_166 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_fill_2 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_201 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_fill_2 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_259 ();
 sg13g2_fill_1 FILLER_19_364 ();
 sg13g2_fill_2 FILLER_20_46 ();
 sg13g2_fill_1 FILLER_20_48 ();
 sg13g2_fill_2 FILLER_20_92 ();
 sg13g2_fill_1 FILLER_20_94 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_fill_1 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_191 ();
 sg13g2_fill_2 FILLER_20_211 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_268 ();
 sg13g2_fill_1 FILLER_20_321 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_fill_1 FILLER_21_26 ();
 sg13g2_fill_1 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_fill_2 FILLER_21_48 ();
 sg13g2_fill_2 FILLER_21_73 ();
 sg13g2_fill_1 FILLER_21_92 ();
 sg13g2_fill_2 FILLER_21_103 ();
 sg13g2_fill_2 FILLER_21_118 ();
 sg13g2_fill_1 FILLER_21_120 ();
 sg13g2_fill_2 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_190 ();
 sg13g2_fill_2 FILLER_21_215 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_fill_1 FILLER_21_327 ();
 sg13g2_fill_2 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_55 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_2 FILLER_22_162 ();
 sg13g2_fill_1 FILLER_22_164 ();
 sg13g2_fill_2 FILLER_22_222 ();
 sg13g2_fill_1 FILLER_22_224 ();
 sg13g2_fill_1 FILLER_22_296 ();
 sg13g2_fill_2 FILLER_22_316 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_329 ();
 sg13g2_fill_1 FILLER_22_371 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_97 ();
 sg13g2_fill_2 FILLER_23_124 ();
 sg13g2_fill_2 FILLER_23_130 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_fill_2 FILLER_23_157 ();
 sg13g2_fill_1 FILLER_23_164 ();
 sg13g2_fill_2 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_204 ();
 sg13g2_fill_2 FILLER_23_299 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_60 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_fill_2 FILLER_24_164 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_186 ();
 sg13g2_fill_2 FILLER_24_228 ();
 sg13g2_fill_1 FILLER_24_311 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_fill_2 FILLER_25_72 ();
 sg13g2_fill_2 FILLER_25_113 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_26_82 ();
 sg13g2_fill_2 FILLER_26_143 ();
 sg13g2_fill_1 FILLER_26_145 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_2 FILLER_26_244 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_371 ();
 sg13g2_fill_2 FILLER_26_391 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_1 FILLER_28_53 ();
 sg13g2_fill_1 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_153 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_fill_2 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_fill_1 FILLER_29_26 ();
 sg13g2_fill_1 FILLER_29_41 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_165 ();
 sg13g2_fill_2 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_298 ();
 sg13g2_fill_1 FILLER_29_353 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_fill_1 FILLER_30_67 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_371 ();
 sg13g2_fill_1 FILLER_31_46 ();
 sg13g2_fill_1 FILLER_31_187 ();
 sg13g2_fill_1 FILLER_31_289 ();
 sg13g2_fill_2 FILLER_32_17 ();
 sg13g2_fill_2 FILLER_32_37 ();
 sg13g2_fill_2 FILLER_32_288 ();
 sg13g2_fill_1 FILLER_32_325 ();
 sg13g2_fill_2 FILLER_33_83 ();
 sg13g2_fill_2 FILLER_33_139 ();
 sg13g2_fill_2 FILLER_33_172 ();
 sg13g2_fill_1 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_210 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_397 ();
 sg13g2_fill_1 FILLER_33_399 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_54 ();
 sg13g2_fill_2 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_198 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_2 FILLER_35_23 ();
 sg13g2_fill_1 FILLER_35_67 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_fill_1 FILLER_35_185 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_fill_1 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_257 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_36_26 ();
 sg13g2_fill_2 FILLER_36_44 ();
 sg13g2_fill_2 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_130 ();
 sg13g2_fill_2 FILLER_36_225 ();
 sg13g2_fill_2 FILLER_36_241 ();
 sg13g2_fill_1 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_2 FILLER_37_24 ();
 sg13g2_fill_2 FILLER_37_34 ();
 sg13g2_fill_2 FILLER_37_153 ();
 sg13g2_fill_2 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_290 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_39 ();
 sg13g2_fill_1 FILLER_38_46 ();
 sg13g2_fill_1 FILLER_38_56 ();
 sg13g2_fill_1 FILLER_38_69 ();
 sg13g2_fill_2 FILLER_38_110 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_220 ();
 sg13g2_fill_2 FILLER_38_251 ();
 sg13g2_fill_1 FILLER_38_253 ();
 sg13g2_fill_2 FILLER_38_337 ();
 assign uio_oe[0] = net8;
 assign uio_oe[1] = net9;
 assign uio_oe[2] = net20;
 assign uio_oe[3] = net10;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[3] = net13;
endmodule

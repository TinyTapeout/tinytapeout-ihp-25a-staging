module tt_um_two_lif_stdp (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire \lif1.spike ;
 wire \lif1.state[0] ;
 wire \lif1.state[1] ;
 wire \lif1.state[2] ;
 wire \lif1.state[3] ;
 wire \lif1.state[4] ;
 wire \lif1.state[5] ;
 wire \lif1.state[6] ;
 wire \lif1.state[7] ;
 wire \lif2.spike ;
 wire \lif2.weight[0] ;
 wire \lif2.weight[1] ;
 wire \lif2.weight[2] ;
 wire \lif2.weight[3] ;
 wire \lif2.weight[4] ;
 wire \lif2.weight[5] ;
 wire \lif2.weight[6] ;
 wire \lif2.weight[7] ;
 wire \stdp1.post_counter[0] ;
 wire \stdp1.post_counter[1] ;
 wire \stdp1.post_counter[2] ;
 wire \stdp1.post_counter[3] ;
 wire \stdp1.pre_counter[0] ;
 wire \stdp1.pre_counter[1] ;
 wire \stdp1.pre_counter[2] ;
 wire \stdp1.pre_counter[3] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;

 sg13g2_inv_1 _480_ (.Y(_440_),
    .A(uo_out[4]));
 sg13g2_inv_1 _481_ (.Y(_441_),
    .A(net25));
 sg13g2_inv_1 _482_ (.Y(_442_),
    .A(net134));
 sg13g2_inv_1 _483_ (.Y(_443_),
    .A(net23));
 sg13g2_a21oi_1 _484_ (.A1(uo_out[1]),
    .A2(uo_out[2]),
    .Y(_444_),
    .B1(uo_out[3]));
 sg13g2_nor2_1 _485_ (.A(uo_out[5]),
    .B(uo_out[6]),
    .Y(_445_));
 sg13g2_o21ai_1 _486_ (.B1(_445_),
    .Y(_446_),
    .A1(_440_),
    .A2(_444_));
 sg13g2_nand2_1 _487_ (.Y(_447_),
    .A(uo_out[7]),
    .B(_446_));
 sg13g2_inv_2 _488_ (.Y(\lif2.spike ),
    .A(net124));
 sg13g2_a21oi_1 _489_ (.A1(\lif1.state[1] ),
    .A2(net137),
    .Y(_448_),
    .B1(net136));
 sg13g2_nor2_1 _490_ (.A(net132),
    .B(net129),
    .Y(_449_));
 sg13g2_o21ai_1 _491_ (.B1(_449_),
    .Y(_450_),
    .A1(_442_),
    .A2(_448_));
 sg13g2_nand2_2 _492_ (.Y(_451_),
    .A(net50),
    .B(_450_));
 sg13g2_inv_2 _493_ (.Y(\lif1.spike ),
    .A(_451_));
 sg13g2_and2_1 _494_ (.A(net137),
    .B(net1),
    .X(_452_));
 sg13g2_nor2_1 _495_ (.A(net137),
    .B(net1),
    .Y(_453_));
 sg13g2_nor3_1 _496_ (.A(\lif1.spike ),
    .B(_452_),
    .C(_453_),
    .Y(_000_));
 sg13g2_and2_1 _497_ (.A(net136),
    .B(net2),
    .X(_454_));
 sg13g2_xor2_1 _498_ (.B(net2),
    .A(net136),
    .X(_039_));
 sg13g2_and2_1 _499_ (.A(_452_),
    .B(_039_),
    .X(_040_));
 sg13g2_nor2_1 _500_ (.A(_452_),
    .B(_039_),
    .Y(_041_));
 sg13g2_nor3_1 _501_ (.A(\lif1.spike ),
    .B(_040_),
    .C(_041_),
    .Y(_001_));
 sg13g2_nor2_1 _502_ (.A(_454_),
    .B(_040_),
    .Y(_042_));
 sg13g2_nand2_1 _503_ (.Y(_043_),
    .A(net133),
    .B(net3));
 sg13g2_xnor2_1 _504_ (.Y(_044_),
    .A(net133),
    .B(net3));
 sg13g2_or2_1 _505_ (.X(_045_),
    .B(_044_),
    .A(_042_));
 sg13g2_nand2_1 _506_ (.Y(_046_),
    .A(_451_),
    .B(_045_));
 sg13g2_a21oi_1 _507_ (.A1(_042_),
    .A2(_044_),
    .Y(_002_),
    .B1(_046_));
 sg13g2_nand2_1 _508_ (.Y(_047_),
    .A(net131),
    .B(net4));
 sg13g2_xnor2_1 _509_ (.Y(_048_),
    .A(net132),
    .B(net4));
 sg13g2_nand3_1 _510_ (.B(_045_),
    .C(_048_),
    .A(_043_),
    .Y(_049_));
 sg13g2_a21o_1 _511_ (.A2(_045_),
    .A1(_043_),
    .B1(_048_),
    .X(_050_));
 sg13g2_and3_1 _512_ (.X(_003_),
    .A(_451_),
    .B(_049_),
    .C(_050_));
 sg13g2_nand2_1 _513_ (.Y(_051_),
    .A(net129),
    .B(net5));
 sg13g2_xnor2_1 _514_ (.Y(_052_),
    .A(net130),
    .B(net5));
 sg13g2_nand3_1 _515_ (.B(_050_),
    .C(_052_),
    .A(_047_),
    .Y(_053_));
 sg13g2_a21o_1 _516_ (.A2(_050_),
    .A1(_047_),
    .B1(_052_),
    .X(_054_));
 sg13g2_and3_1 _517_ (.X(_004_),
    .A(_451_),
    .B(_053_),
    .C(_054_));
 sg13g2_xnor2_1 _518_ (.Y(_055_),
    .A(net50),
    .B(net6));
 sg13g2_and3_1 _519_ (.X(_056_),
    .A(_051_),
    .B(_054_),
    .C(_055_));
 sg13g2_a21oi_1 _520_ (.A1(_051_),
    .A2(_054_),
    .Y(_057_),
    .B1(_055_));
 sg13g2_nor3_1 _521_ (.A(\lif1.spike ),
    .B(_056_),
    .C(_057_),
    .Y(_005_));
 sg13g2_a21oi_1 _522_ (.A1(net50),
    .A2(net6),
    .Y(_058_),
    .B1(_057_));
 sg13g2_nor2b_1 _523_ (.A(net7),
    .B_N(_058_),
    .Y(_059_));
 sg13g2_nor2b_1 _524_ (.A(_058_),
    .B_N(net7),
    .Y(_060_));
 sg13g2_nor3_1 _525_ (.A(\lif1.spike ),
    .B(_059_),
    .C(_060_),
    .Y(_006_));
 sg13g2_o21ai_1 _526_ (.B1(_451_),
    .Y(_061_),
    .A1(net8),
    .A2(_060_));
 sg13g2_a21oi_1 _527_ (.A1(net8),
    .A2(_060_),
    .Y(_007_),
    .B1(_061_));
 sg13g2_nand2_2 _528_ (.Y(_062_),
    .A(\lif1.state[0] ),
    .B(net148));
 sg13g2_nand2_2 _529_ (.Y(_063_),
    .A(net139),
    .B(net146));
 sg13g2_nor2_1 _530_ (.A(_062_),
    .B(_063_),
    .Y(_064_));
 sg13g2_or2_1 _531_ (.X(_065_),
    .B(_063_),
    .A(_062_));
 sg13g2_and4_1 _532_ (.A(net136),
    .B(net138),
    .C(net152),
    .D(net126),
    .X(_066_));
 sg13g2_nand4_1 _533_ (.B(net137),
    .C(net152),
    .A(net136),
    .Y(_067_),
    .D(net127));
 sg13g2_nand2_1 _534_ (.Y(_068_),
    .A(net139),
    .B(net150));
 sg13g2_a22oi_1 _535_ (.Y(_069_),
    .B1(net126),
    .B2(net136),
    .A2(net152),
    .A1(net137));
 sg13g2_or3_1 _536_ (.A(_066_),
    .B(_068_),
    .C(_069_),
    .X(_070_));
 sg13g2_o21ai_1 _537_ (.B1(_067_),
    .Y(_071_),
    .A1(_068_),
    .A2(_069_));
 sg13g2_nand2_1 _538_ (.Y(_072_),
    .A(net138),
    .B(net150));
 sg13g2_and4_1 _539_ (.A(net135),
    .B(net134),
    .C(net152),
    .D(net126),
    .X(_073_));
 sg13g2_nand4_1 _540_ (.B(net133),
    .C(net151),
    .A(net135),
    .Y(_074_),
    .D(net125));
 sg13g2_a22oi_1 _541_ (.Y(_075_),
    .B1(net125),
    .B2(net134),
    .A2(net151),
    .A1(net135));
 sg13g2_or3_1 _542_ (.A(_072_),
    .B(_073_),
    .C(_075_),
    .X(_076_));
 sg13g2_o21ai_1 _543_ (.B1(_072_),
    .Y(_077_),
    .A1(_073_),
    .A2(_075_));
 sg13g2_and3_1 _544_ (.X(_078_),
    .A(_071_),
    .B(_076_),
    .C(_077_));
 sg13g2_a22oi_1 _545_ (.Y(_079_),
    .B1(net146),
    .B2(\lif1.state[0] ),
    .A2(net148),
    .A1(\lif1.state[1] ));
 sg13g2_nor2_1 _546_ (.A(_064_),
    .B(_079_),
    .Y(_080_));
 sg13g2_a21oi_1 _547_ (.A1(_076_),
    .A2(_077_),
    .Y(_081_),
    .B1(_071_));
 sg13g2_a21o_1 _548_ (.A2(_077_),
    .A1(_076_),
    .B1(_071_),
    .X(_082_));
 sg13g2_a21o_1 _549_ (.A2(_082_),
    .A1(_080_),
    .B1(_078_),
    .X(_083_));
 sg13g2_o21ai_1 _550_ (.B1(_074_),
    .Y(_084_),
    .A1(_072_),
    .A2(_075_));
 sg13g2_nand2_1 _551_ (.Y(_085_),
    .A(net135),
    .B(net150));
 sg13g2_and4_1 _552_ (.A(net131),
    .B(net133),
    .C(net151),
    .D(net125),
    .X(_086_));
 sg13g2_nand4_1 _553_ (.B(net133),
    .C(net151),
    .A(net131),
    .Y(_087_),
    .D(net125));
 sg13g2_a22oi_1 _554_ (.Y(_088_),
    .B1(net125),
    .B2(net131),
    .A2(net151),
    .A1(net133));
 sg13g2_or3_1 _555_ (.A(_085_),
    .B(_086_),
    .C(_088_),
    .X(_089_));
 sg13g2_o21ai_1 _556_ (.B1(_085_),
    .Y(_090_),
    .A1(_086_),
    .A2(_088_));
 sg13g2_and3_1 _557_ (.X(_091_),
    .A(_084_),
    .B(_089_),
    .C(_090_));
 sg13g2_nand3_1 _558_ (.B(_089_),
    .C(_090_),
    .A(_084_),
    .Y(_092_));
 sg13g2_a21oi_1 _559_ (.A1(_089_),
    .A2(_090_),
    .Y(_093_),
    .B1(_084_));
 sg13g2_nand2_1 _560_ (.Y(_094_),
    .A(\lif1.state[0] ),
    .B(net144));
 sg13g2_nand2_1 _561_ (.Y(_095_),
    .A(net138),
    .B(net145));
 sg13g2_nand2_1 _562_ (.Y(_096_),
    .A(net138),
    .B(net148));
 sg13g2_xor2_1 _563_ (.B(_096_),
    .A(_063_),
    .X(_097_));
 sg13g2_nand2b_1 _564_ (.Y(_098_),
    .B(_097_),
    .A_N(_094_));
 sg13g2_xor2_1 _565_ (.B(_097_),
    .A(_094_),
    .X(_099_));
 sg13g2_or3_1 _566_ (.A(_091_),
    .B(_093_),
    .C(_099_),
    .X(_100_));
 sg13g2_o21ai_1 _567_ (.B1(_099_),
    .Y(_101_),
    .A1(_091_),
    .A2(_093_));
 sg13g2_nand3_1 _568_ (.B(_100_),
    .C(_101_),
    .A(_083_),
    .Y(_102_));
 sg13g2_a21oi_1 _569_ (.A1(_100_),
    .A2(_101_),
    .Y(_103_),
    .B1(_083_));
 sg13g2_a21o_1 _570_ (.A2(_101_),
    .A1(_100_),
    .B1(_083_),
    .X(_104_));
 sg13g2_nand2_1 _571_ (.Y(_105_),
    .A(_102_),
    .B(_104_));
 sg13g2_xnor2_1 _572_ (.Y(_106_),
    .A(_064_),
    .B(_105_));
 sg13g2_and4_1 _573_ (.A(net139),
    .B(net137),
    .C(net152),
    .D(net126),
    .X(_107_));
 sg13g2_a22oi_1 _574_ (.Y(_108_),
    .B1(net126),
    .B2(net137),
    .A2(net152),
    .A1(net139));
 sg13g2_nand2_1 _575_ (.Y(_109_),
    .A(\lif1.state[0] ),
    .B(net150));
 sg13g2_nor3_1 _576_ (.A(_107_),
    .B(_108_),
    .C(_109_),
    .Y(_110_));
 sg13g2_or2_1 _577_ (.X(_111_),
    .B(_110_),
    .A(_107_));
 sg13g2_o21ai_1 _578_ (.B1(_068_),
    .Y(_112_),
    .A1(_066_),
    .A2(_069_));
 sg13g2_and3_1 _579_ (.X(_113_),
    .A(_070_),
    .B(_111_),
    .C(_112_));
 sg13g2_nand3_1 _580_ (.B(_111_),
    .C(_112_),
    .A(_070_),
    .Y(_114_));
 sg13g2_a21oi_1 _581_ (.A1(_070_),
    .A2(_112_),
    .Y(_115_),
    .B1(_111_));
 sg13g2_nor2_1 _582_ (.A(_113_),
    .B(_115_),
    .Y(_116_));
 sg13g2_o21ai_1 _583_ (.B1(_114_),
    .Y(_117_),
    .A1(_062_),
    .A2(_115_));
 sg13g2_nor3_1 _584_ (.A(_078_),
    .B(_080_),
    .C(_081_),
    .Y(_118_));
 sg13g2_o21ai_1 _585_ (.B1(_080_),
    .Y(_119_),
    .A1(_078_),
    .A2(_081_));
 sg13g2_nand2b_1 _586_ (.Y(_120_),
    .B(_119_),
    .A_N(_118_));
 sg13g2_nor2_1 _587_ (.A(_117_),
    .B(_120_),
    .Y(_121_));
 sg13g2_and2_1 _588_ (.A(_117_),
    .B(_120_),
    .X(_122_));
 sg13g2_nand2_1 _589_ (.Y(_123_),
    .A(_117_),
    .B(_120_));
 sg13g2_nand4_1 _590_ (.B(\lif1.state[0] ),
    .C(net152),
    .A(net139),
    .Y(_124_),
    .D(net126));
 sg13g2_and3_1 _591_ (.X(_125_),
    .A(net137),
    .B(net126),
    .C(_109_));
 sg13g2_xnor2_1 _592_ (.Y(_126_),
    .A(_062_),
    .B(_116_));
 sg13g2_nor4_1 _593_ (.A(_110_),
    .B(_121_),
    .C(_124_),
    .D(_125_),
    .Y(_127_));
 sg13g2_nand4_1 _594_ (.B(_123_),
    .C(_126_),
    .A(_106_),
    .Y(_128_),
    .D(_127_));
 sg13g2_o21ai_1 _595_ (.B1(_102_),
    .Y(_129_),
    .A1(_065_),
    .A2(_103_));
 sg13g2_o21ai_1 _596_ (.B1(_098_),
    .Y(_130_),
    .A1(_063_),
    .A2(_096_));
 sg13g2_nand2_1 _597_ (.Y(_131_),
    .A(\lif1.state[0] ),
    .B(net142));
 sg13g2_nand2b_1 _598_ (.Y(_132_),
    .B(_130_),
    .A_N(_131_));
 sg13g2_inv_1 _599_ (.Y(_133_),
    .A(_132_));
 sg13g2_xnor2_1 _600_ (.Y(_134_),
    .A(_130_),
    .B(_131_));
 sg13g2_xor2_1 _601_ (.B(_131_),
    .A(_130_),
    .X(_135_));
 sg13g2_o21ai_1 _602_ (.B1(_092_),
    .Y(_136_),
    .A1(_093_),
    .A2(_099_));
 sg13g2_nand2_1 _603_ (.Y(_137_),
    .A(net139),
    .B(net144));
 sg13g2_nand2_1 _604_ (.Y(_138_),
    .A(net135),
    .B(net145));
 sg13g2_nand2_1 _605_ (.Y(_139_),
    .A(net136),
    .B(net148));
 sg13g2_or2_1 _606_ (.X(_140_),
    .B(_138_),
    .A(_096_));
 sg13g2_xnor2_1 _607_ (.Y(_141_),
    .A(_095_),
    .B(_139_));
 sg13g2_xnor2_1 _608_ (.Y(_142_),
    .A(_137_),
    .B(_141_));
 sg13g2_o21ai_1 _609_ (.B1(_087_),
    .Y(_143_),
    .A1(_085_),
    .A2(_088_));
 sg13g2_nand2_1 _610_ (.Y(_144_),
    .A(net133),
    .B(net150));
 sg13g2_nand2_1 _611_ (.Y(_145_),
    .A(net130),
    .B(net153));
 sg13g2_and4_1 _612_ (.A(net131),
    .B(net129),
    .C(net151),
    .D(net125),
    .X(_146_));
 sg13g2_nand4_1 _613_ (.B(net129),
    .C(net151),
    .A(net131),
    .Y(_147_),
    .D(net125));
 sg13g2_a22oi_1 _614_ (.Y(_148_),
    .B1(net125),
    .B2(net129),
    .A2(net151),
    .A1(net131));
 sg13g2_or3_1 _615_ (.A(_144_),
    .B(_146_),
    .C(_148_),
    .X(_149_));
 sg13g2_o21ai_1 _616_ (.B1(_144_),
    .Y(_150_),
    .A1(_146_),
    .A2(_148_));
 sg13g2_and3_1 _617_ (.X(_151_),
    .A(_143_),
    .B(_149_),
    .C(_150_));
 sg13g2_nand3_1 _618_ (.B(_149_),
    .C(_150_),
    .A(_143_),
    .Y(_152_));
 sg13g2_a21oi_1 _619_ (.A1(_149_),
    .A2(_150_),
    .Y(_153_),
    .B1(_143_));
 sg13g2_or3_1 _620_ (.A(_142_),
    .B(_151_),
    .C(_153_),
    .X(_154_));
 sg13g2_o21ai_1 _621_ (.B1(_142_),
    .Y(_155_),
    .A1(_151_),
    .A2(_153_));
 sg13g2_nand3_1 _622_ (.B(_154_),
    .C(_155_),
    .A(_136_),
    .Y(_156_));
 sg13g2_a21oi_1 _623_ (.A1(_154_),
    .A2(_155_),
    .Y(_157_),
    .B1(_136_));
 sg13g2_a21o_1 _624_ (.A2(_155_),
    .A1(_154_),
    .B1(_136_),
    .X(_158_));
 sg13g2_nand3_1 _625_ (.B(_156_),
    .C(_158_),
    .A(_134_),
    .Y(_159_));
 sg13g2_a21o_1 _626_ (.A2(_158_),
    .A1(_156_),
    .B1(_134_),
    .X(_160_));
 sg13g2_nand3_1 _627_ (.B(_159_),
    .C(_160_),
    .A(_129_),
    .Y(_161_));
 sg13g2_a21o_1 _628_ (.A2(_160_),
    .A1(_159_),
    .B1(_129_),
    .X(_162_));
 sg13g2_nand2_1 _629_ (.Y(_163_),
    .A(_161_),
    .B(_162_));
 sg13g2_nand2_1 _630_ (.Y(_164_),
    .A(_106_),
    .B(_122_));
 sg13g2_nand4_1 _631_ (.B(_122_),
    .C(_161_),
    .A(_106_),
    .Y(_165_),
    .D(_162_));
 sg13g2_a22oi_1 _632_ (.Y(_166_),
    .B1(_161_),
    .B2(_162_),
    .A2(_122_),
    .A1(_106_));
 sg13g2_xor2_1 _633_ (.B(_164_),
    .A(_163_),
    .X(_167_));
 sg13g2_xnor2_1 _634_ (.Y(_168_),
    .A(_128_),
    .B(_167_));
 sg13g2_nand2_1 _635_ (.Y(_169_),
    .A(net35),
    .B(_168_));
 sg13g2_o21ai_1 _636_ (.B1(net124),
    .Y(_170_),
    .A1(net35),
    .A2(_168_));
 sg13g2_nor2b_1 _637_ (.A(_170_),
    .B_N(_169_),
    .Y(_008_));
 sg13g2_o21ai_1 _638_ (.B1(_165_),
    .Y(_171_),
    .A1(_128_),
    .A2(_166_));
 sg13g2_o21ai_1 _639_ (.B1(_156_),
    .Y(_172_),
    .A1(_135_),
    .A2(_157_));
 sg13g2_nand2_1 _640_ (.Y(_173_),
    .A(\lif1.state[0] ),
    .B(net140));
 sg13g2_o21ai_1 _641_ (.B1(_140_),
    .Y(_174_),
    .A1(_137_),
    .A2(_141_));
 sg13g2_nand2_1 _642_ (.Y(_175_),
    .A(net139),
    .B(net141));
 sg13g2_nand2b_1 _643_ (.Y(_176_),
    .B(_174_),
    .A_N(_175_));
 sg13g2_xnor2_1 _644_ (.Y(_177_),
    .A(_174_),
    .B(_175_));
 sg13g2_nand2b_1 _645_ (.Y(_178_),
    .B(_177_),
    .A_N(_173_));
 sg13g2_xnor2_1 _646_ (.Y(_179_),
    .A(_173_),
    .B(_177_));
 sg13g2_o21ai_1 _647_ (.B1(_152_),
    .Y(_180_),
    .A1(_142_),
    .A2(_153_));
 sg13g2_nand2_1 _648_ (.Y(_181_),
    .A(net138),
    .B(net144));
 sg13g2_nand2_1 _649_ (.Y(_182_),
    .A(net134),
    .B(net146));
 sg13g2_nand2_1 _650_ (.Y(_183_),
    .A(net133),
    .B(net148));
 sg13g2_xor2_1 _651_ (.B(_183_),
    .A(_138_),
    .X(_184_));
 sg13g2_nand2b_1 _652_ (.Y(_185_),
    .B(_184_),
    .A_N(_181_));
 sg13g2_xnor2_1 _653_ (.Y(_186_),
    .A(_181_),
    .B(_184_));
 sg13g2_o21ai_1 _654_ (.B1(_147_),
    .Y(_187_),
    .A1(_144_),
    .A2(_148_));
 sg13g2_nand2_1 _655_ (.Y(_188_),
    .A(net131),
    .B(net150));
 sg13g2_nand2_1 _656_ (.Y(_189_),
    .A(net128),
    .B(net153));
 sg13g2_and4_1 _657_ (.A(net129),
    .B(net128),
    .C(net153),
    .D(net127),
    .X(_190_));
 sg13g2_a22oi_1 _658_ (.Y(_191_),
    .B1(net127),
    .B2(net128),
    .A2(net153),
    .A1(net129));
 sg13g2_or3_1 _659_ (.A(_188_),
    .B(_190_),
    .C(_191_),
    .X(_192_));
 sg13g2_o21ai_1 _660_ (.B1(_188_),
    .Y(_193_),
    .A1(_190_),
    .A2(_191_));
 sg13g2_nand3_1 _661_ (.B(_192_),
    .C(_193_),
    .A(_187_),
    .Y(_194_));
 sg13g2_a21o_1 _662_ (.A2(_193_),
    .A1(_192_),
    .B1(_187_),
    .X(_195_));
 sg13g2_nand3_1 _663_ (.B(_194_),
    .C(_195_),
    .A(_186_),
    .Y(_196_));
 sg13g2_a21o_1 _664_ (.A2(_195_),
    .A1(_194_),
    .B1(_186_),
    .X(_197_));
 sg13g2_nand3_1 _665_ (.B(_196_),
    .C(_197_),
    .A(_180_),
    .Y(_198_));
 sg13g2_a21o_1 _666_ (.A2(_197_),
    .A1(_196_),
    .B1(_180_),
    .X(_199_));
 sg13g2_nand3_1 _667_ (.B(_198_),
    .C(_199_),
    .A(_179_),
    .Y(_200_));
 sg13g2_a21o_1 _668_ (.A2(_199_),
    .A1(_198_),
    .B1(_179_),
    .X(_201_));
 sg13g2_nand3_1 _669_ (.B(_200_),
    .C(_201_),
    .A(_172_),
    .Y(_202_));
 sg13g2_a21o_1 _670_ (.A2(_201_),
    .A1(_200_),
    .B1(_172_),
    .X(_203_));
 sg13g2_and3_1 _671_ (.X(_204_),
    .A(_133_),
    .B(_202_),
    .C(_203_));
 sg13g2_nand3_1 _672_ (.B(_202_),
    .C(_203_),
    .A(_133_),
    .Y(_205_));
 sg13g2_a21oi_1 _673_ (.A1(_202_),
    .A2(_203_),
    .Y(_206_),
    .B1(_133_));
 sg13g2_nor3_1 _674_ (.A(_161_),
    .B(_204_),
    .C(_206_),
    .Y(_207_));
 sg13g2_or3_1 _675_ (.A(_161_),
    .B(_204_),
    .C(_206_),
    .X(_208_));
 sg13g2_o21ai_1 _676_ (.B1(_161_),
    .Y(_209_),
    .A1(_204_),
    .A2(_206_));
 sg13g2_nand3_1 _677_ (.B(_208_),
    .C(_209_),
    .A(_171_),
    .Y(_210_));
 sg13g2_a21o_1 _678_ (.A2(_209_),
    .A1(_208_),
    .B1(_171_),
    .X(_211_));
 sg13g2_nand3_1 _679_ (.B(_210_),
    .C(_211_),
    .A(uo_out[3]),
    .Y(_212_));
 sg13g2_a21oi_1 _680_ (.A1(_210_),
    .A2(_211_),
    .Y(_213_),
    .B1(uo_out[3]));
 sg13g2_a21o_1 _681_ (.A2(_211_),
    .A1(_210_),
    .B1(net40),
    .X(_214_));
 sg13g2_nand2_1 _682_ (.Y(_215_),
    .A(_212_),
    .B(_214_));
 sg13g2_o21ai_1 _683_ (.B1(net124),
    .Y(_216_),
    .A1(_169_),
    .A2(_215_));
 sg13g2_a21oi_1 _684_ (.A1(_169_),
    .A2(_215_),
    .Y(_009_),
    .B1(_216_));
 sg13g2_o21ai_1 _685_ (.B1(_212_),
    .Y(_217_),
    .A1(_169_),
    .A2(_213_));
 sg13g2_a21oi_1 _686_ (.A1(_171_),
    .A2(_209_),
    .Y(_218_),
    .B1(_207_));
 sg13g2_nand2_1 _687_ (.Y(_219_),
    .A(_202_),
    .B(_205_));
 sg13g2_nand2_1 _688_ (.Y(_220_),
    .A(_176_),
    .B(_178_));
 sg13g2_nand2_1 _689_ (.Y(_221_),
    .A(_198_),
    .B(_200_));
 sg13g2_nand2_1 _690_ (.Y(_222_),
    .A(net139),
    .B(net140));
 sg13g2_o21ai_1 _691_ (.B1(_185_),
    .Y(_223_),
    .A1(_138_),
    .A2(_183_));
 sg13g2_nand2_1 _692_ (.Y(_224_),
    .A(net138),
    .B(net141));
 sg13g2_nand2b_1 _693_ (.Y(_225_),
    .B(_223_),
    .A_N(_224_));
 sg13g2_xnor2_1 _694_ (.Y(_226_),
    .A(_223_),
    .B(_224_));
 sg13g2_nand2b_1 _695_ (.Y(_227_),
    .B(_226_),
    .A_N(_222_));
 sg13g2_xnor2_1 _696_ (.Y(_228_),
    .A(_222_),
    .B(_226_));
 sg13g2_nand2_1 _697_ (.Y(_229_),
    .A(_194_),
    .B(_196_));
 sg13g2_nand2_1 _698_ (.Y(_230_),
    .A(net135),
    .B(net144));
 sg13g2_nand2_1 _699_ (.Y(_231_),
    .A(net132),
    .B(net146));
 sg13g2_nand2_1 _700_ (.Y(_232_),
    .A(net132),
    .B(net148));
 sg13g2_xor2_1 _701_ (.B(_232_),
    .A(_182_),
    .X(_233_));
 sg13g2_nand2b_1 _702_ (.Y(_234_),
    .B(_233_),
    .A_N(_230_));
 sg13g2_xnor2_1 _703_ (.Y(_235_),
    .A(_230_),
    .B(_233_));
 sg13g2_inv_1 _704_ (.Y(_236_),
    .A(_235_));
 sg13g2_nand2b_1 _705_ (.Y(_237_),
    .B(_192_),
    .A_N(_190_));
 sg13g2_nand2_1 _706_ (.Y(_238_),
    .A(net129),
    .B(net150));
 sg13g2_nand2_1 _707_ (.Y(_239_),
    .A(net128),
    .B(net150));
 sg13g2_xor2_1 _708_ (.B(_238_),
    .A(_189_),
    .X(_240_));
 sg13g2_xnor2_1 _709_ (.Y(_241_),
    .A(_237_),
    .B(_240_));
 sg13g2_nor2_1 _710_ (.A(_236_),
    .B(_241_),
    .Y(_242_));
 sg13g2_xnor2_1 _711_ (.Y(_243_),
    .A(_236_),
    .B(_241_));
 sg13g2_nor2b_1 _712_ (.A(_243_),
    .B_N(_229_),
    .Y(_244_));
 sg13g2_nand2b_1 _713_ (.Y(_245_),
    .B(_243_),
    .A_N(_229_));
 sg13g2_xnor2_1 _714_ (.Y(_246_),
    .A(_229_),
    .B(_243_));
 sg13g2_xnor2_1 _715_ (.Y(_247_),
    .A(_228_),
    .B(_246_));
 sg13g2_nor2b_1 _716_ (.A(_247_),
    .B_N(_221_),
    .Y(_248_));
 sg13g2_xor2_1 _717_ (.B(_247_),
    .A(_221_),
    .X(_249_));
 sg13g2_nor2b_1 _718_ (.A(_249_),
    .B_N(_220_),
    .Y(_250_));
 sg13g2_xnor2_1 _719_ (.Y(_251_),
    .A(_220_),
    .B(_249_));
 sg13g2_nand2_1 _720_ (.Y(_252_),
    .A(_219_),
    .B(_251_));
 sg13g2_xnor2_1 _721_ (.Y(_253_),
    .A(_219_),
    .B(_251_));
 sg13g2_xor2_1 _722_ (.B(_253_),
    .A(_218_),
    .X(_254_));
 sg13g2_and2_1 _723_ (.A(net51),
    .B(_254_),
    .X(_255_));
 sg13g2_or2_1 _724_ (.X(_256_),
    .B(_254_),
    .A(uo_out[4]));
 sg13g2_nor2b_1 _725_ (.A(_255_),
    .B_N(_256_),
    .Y(_257_));
 sg13g2_o21ai_1 _726_ (.B1(net124),
    .Y(_258_),
    .A1(_217_),
    .A2(_257_));
 sg13g2_a21oi_1 _727_ (.A1(_217_),
    .A2(_257_),
    .Y(_010_),
    .B1(_258_));
 sg13g2_a21oi_1 _728_ (.A1(_217_),
    .A2(_256_),
    .Y(_259_),
    .B1(_255_));
 sg13g2_o21ai_1 _729_ (.B1(_252_),
    .Y(_260_),
    .A1(_218_),
    .A2(_253_));
 sg13g2_nor2_1 _730_ (.A(_248_),
    .B(_250_),
    .Y(_261_));
 sg13g2_nand2_1 _731_ (.Y(_262_),
    .A(_225_),
    .B(_227_));
 sg13g2_a21o_1 _732_ (.A2(_245_),
    .A1(_228_),
    .B1(_244_),
    .X(_263_));
 sg13g2_nand2_1 _733_ (.Y(_264_),
    .A(net138),
    .B(net140));
 sg13g2_o21ai_1 _734_ (.B1(_234_),
    .Y(_265_),
    .A1(_182_),
    .A2(_232_));
 sg13g2_nand2_1 _735_ (.Y(_266_),
    .A(net135),
    .B(net141));
 sg13g2_nand2b_1 _736_ (.Y(_267_),
    .B(_265_),
    .A_N(_266_));
 sg13g2_xnor2_1 _737_ (.Y(_268_),
    .A(_265_),
    .B(_266_));
 sg13g2_nand2b_1 _738_ (.Y(_269_),
    .B(_268_),
    .A_N(_264_));
 sg13g2_xor2_1 _739_ (.B(_268_),
    .A(_264_),
    .X(_270_));
 sg13g2_a21oi_1 _740_ (.A1(_237_),
    .A2(_240_),
    .Y(_271_),
    .B1(_242_));
 sg13g2_nand2b_1 _741_ (.Y(_272_),
    .B(_145_),
    .A_N(_239_));
 sg13g2_nand2_1 _742_ (.Y(_273_),
    .A(net134),
    .B(net144));
 sg13g2_nand2_2 _743_ (.Y(_274_),
    .A(net130),
    .B(net145));
 sg13g2_nand2_1 _744_ (.Y(_275_),
    .A(net130),
    .B(net148));
 sg13g2_or2_1 _745_ (.X(_276_),
    .B(_274_),
    .A(_232_));
 sg13g2_xnor2_1 _746_ (.Y(_277_),
    .A(_231_),
    .B(_275_));
 sg13g2_xnor2_1 _747_ (.Y(_278_),
    .A(_273_),
    .B(_277_));
 sg13g2_xnor2_1 _748_ (.Y(_279_),
    .A(_272_),
    .B(_278_));
 sg13g2_nor2_1 _749_ (.A(_271_),
    .B(_279_),
    .Y(_280_));
 sg13g2_xnor2_1 _750_ (.Y(_281_),
    .A(_271_),
    .B(_279_));
 sg13g2_nor2_1 _751_ (.A(_270_),
    .B(_281_),
    .Y(_282_));
 sg13g2_xnor2_1 _752_ (.Y(_283_),
    .A(_270_),
    .B(_281_));
 sg13g2_nor2b_1 _753_ (.A(_283_),
    .B_N(_263_),
    .Y(_284_));
 sg13g2_xnor2_1 _754_ (.Y(_285_),
    .A(_263_),
    .B(_283_));
 sg13g2_xnor2_1 _755_ (.Y(_286_),
    .A(_262_),
    .B(_285_));
 sg13g2_nor2_1 _756_ (.A(_261_),
    .B(_286_),
    .Y(_287_));
 sg13g2_xor2_1 _757_ (.B(_286_),
    .A(_261_),
    .X(_288_));
 sg13g2_xnor2_1 _758_ (.Y(_289_),
    .A(_260_),
    .B(_288_));
 sg13g2_or2_1 _759_ (.X(_290_),
    .B(_289_),
    .A(net31));
 sg13g2_xnor2_1 _760_ (.Y(_291_),
    .A(net31),
    .B(_289_));
 sg13g2_o21ai_1 _761_ (.B1(_447_),
    .Y(_292_),
    .A1(_259_),
    .A2(_291_));
 sg13g2_a21oi_1 _762_ (.A1(_259_),
    .A2(_291_),
    .Y(_011_),
    .B1(_292_));
 sg13g2_o21ai_1 _763_ (.B1(_290_),
    .Y(_293_),
    .A1(_259_),
    .A2(_291_));
 sg13g2_a21oi_2 _764_ (.B1(_287_),
    .Y(_294_),
    .A2(_288_),
    .A1(_260_));
 sg13g2_a21o_1 _765_ (.A2(_285_),
    .A1(_262_),
    .B1(_284_),
    .X(_295_));
 sg13g2_nand2_1 _766_ (.Y(_296_),
    .A(_267_),
    .B(_269_));
 sg13g2_nor2_1 _767_ (.A(_280_),
    .B(_282_),
    .Y(_297_));
 sg13g2_a21oi_1 _768_ (.A1(_145_),
    .A2(_278_),
    .Y(_298_),
    .B1(_239_));
 sg13g2_nand2_1 _769_ (.Y(_299_),
    .A(net132),
    .B(net144));
 sg13g2_nand2_1 _770_ (.Y(_300_),
    .A(net128),
    .B(net147));
 sg13g2_or2_1 _771_ (.X(_301_),
    .B(_300_),
    .A(_274_));
 sg13g2_xnor2_1 _772_ (.Y(_302_),
    .A(_274_),
    .B(_300_));
 sg13g2_xor2_1 _773_ (.B(_302_),
    .A(_299_),
    .X(_303_));
 sg13g2_and2_1 _774_ (.A(_298_),
    .B(_303_),
    .X(_304_));
 sg13g2_or2_1 _775_ (.X(_305_),
    .B(_303_),
    .A(_298_));
 sg13g2_nand2b_1 _776_ (.Y(_306_),
    .B(_305_),
    .A_N(_304_));
 sg13g2_nand2_1 _777_ (.Y(_307_),
    .A(net135),
    .B(\lif2.weight[7] ));
 sg13g2_o21ai_1 _778_ (.B1(_276_),
    .Y(_308_),
    .A1(_273_),
    .A2(_277_));
 sg13g2_nand2_1 _779_ (.Y(_309_),
    .A(net134),
    .B(net141));
 sg13g2_nand2b_1 _780_ (.Y(_310_),
    .B(_308_),
    .A_N(_309_));
 sg13g2_xnor2_1 _781_ (.Y(_311_),
    .A(_308_),
    .B(_309_));
 sg13g2_nand2b_1 _782_ (.Y(_312_),
    .B(_311_),
    .A_N(_307_));
 sg13g2_xnor2_1 _783_ (.Y(_313_),
    .A(_307_),
    .B(_311_));
 sg13g2_xnor2_1 _784_ (.Y(_314_),
    .A(_306_),
    .B(_313_));
 sg13g2_nor2b_1 _785_ (.A(_297_),
    .B_N(_314_),
    .Y(_315_));
 sg13g2_xnor2_1 _786_ (.Y(_316_),
    .A(_297_),
    .B(_314_));
 sg13g2_xor2_1 _787_ (.B(_316_),
    .A(_296_),
    .X(_317_));
 sg13g2_nand2_1 _788_ (.Y(_318_),
    .A(_295_),
    .B(_317_));
 sg13g2_xnor2_1 _789_ (.Y(_319_),
    .A(_295_),
    .B(_317_));
 sg13g2_xor2_1 _790_ (.B(_319_),
    .A(_294_),
    .X(_320_));
 sg13g2_nor2b_1 _791_ (.A(_018_),
    .B_N(_320_),
    .Y(_321_));
 sg13g2_xnor2_1 _792_ (.Y(_322_),
    .A(net47),
    .B(_320_));
 sg13g2_a21oi_1 _793_ (.A1(_293_),
    .A2(_322_),
    .Y(_323_),
    .B1(\lif2.spike ));
 sg13g2_o21ai_1 _794_ (.B1(_323_),
    .Y(_324_),
    .A1(_293_),
    .A2(_322_));
 sg13g2_inv_1 _795_ (.Y(_012_),
    .A(_324_));
 sg13g2_a21o_1 _796_ (.A2(_322_),
    .A1(_293_),
    .B1(_321_),
    .X(_325_));
 sg13g2_o21ai_1 _797_ (.B1(_318_),
    .Y(_326_),
    .A1(_294_),
    .A2(_319_));
 sg13g2_a21oi_1 _798_ (.A1(_296_),
    .A2(_316_),
    .Y(_327_),
    .B1(_315_));
 sg13g2_a22oi_1 _799_ (.Y(_328_),
    .B1(net145),
    .B2(net128),
    .A2(net144),
    .A1(net130));
 sg13g2_nand2_1 _800_ (.Y(_329_),
    .A(net128),
    .B(net143));
 sg13g2_or2_1 _801_ (.X(_330_),
    .B(_329_),
    .A(_274_));
 sg13g2_inv_1 _802_ (.Y(_331_),
    .A(_330_));
 sg13g2_nand2b_1 _803_ (.Y(_332_),
    .B(_330_),
    .A_N(_328_));
 sg13g2_nand2_1 _804_ (.Y(_333_),
    .A(net134),
    .B(\lif2.weight[7] ));
 sg13g2_o21ai_1 _805_ (.B1(_301_),
    .Y(_334_),
    .A1(_299_),
    .A2(_302_));
 sg13g2_nand2_1 _806_ (.Y(_335_),
    .A(net132),
    .B(net141));
 sg13g2_nand2b_1 _807_ (.Y(_336_),
    .B(_334_),
    .A_N(_335_));
 sg13g2_xnor2_1 _808_ (.Y(_337_),
    .A(_334_),
    .B(_335_));
 sg13g2_nand2b_1 _809_ (.Y(_338_),
    .B(_337_),
    .A_N(_333_));
 sg13g2_xnor2_1 _810_ (.Y(_339_),
    .A(_333_),
    .B(_337_));
 sg13g2_nand2b_1 _811_ (.Y(_340_),
    .B(_339_),
    .A_N(_332_));
 sg13g2_xnor2_1 _812_ (.Y(_341_),
    .A(_332_),
    .B(_339_));
 sg13g2_a21oi_1 _813_ (.A1(_305_),
    .A2(_313_),
    .Y(_342_),
    .B1(_304_));
 sg13g2_nor2b_1 _814_ (.A(_342_),
    .B_N(_341_),
    .Y(_343_));
 sg13g2_xnor2_1 _815_ (.Y(_344_),
    .A(_341_),
    .B(_342_));
 sg13g2_nand2_1 _816_ (.Y(_345_),
    .A(_310_),
    .B(_312_));
 sg13g2_xnor2_1 _817_ (.Y(_346_),
    .A(_344_),
    .B(_345_));
 sg13g2_nor2_1 _818_ (.A(_327_),
    .B(_346_),
    .Y(_347_));
 sg13g2_xor2_1 _819_ (.B(_346_),
    .A(_327_),
    .X(_348_));
 sg13g2_xnor2_1 _820_ (.Y(_349_),
    .A(_326_),
    .B(_348_));
 sg13g2_nor2_1 _821_ (.A(net42),
    .B(_349_),
    .Y(_350_));
 sg13g2_xor2_1 _822_ (.B(_349_),
    .A(net42),
    .X(_351_));
 sg13g2_o21ai_1 _823_ (.B1(net124),
    .Y(_352_),
    .A1(_325_),
    .A2(_351_));
 sg13g2_a21oi_1 _824_ (.A1(_325_),
    .A2(_351_),
    .Y(_013_),
    .B1(_352_));
 sg13g2_a21o_1 _825_ (.A2(_351_),
    .A1(_325_),
    .B1(_350_),
    .X(_353_));
 sg13g2_a21oi_2 _826_ (.B1(_347_),
    .Y(_354_),
    .A2(_348_),
    .A1(_326_));
 sg13g2_a21oi_2 _827_ (.B1(_343_),
    .Y(_355_),
    .A2(_345_),
    .A1(_344_));
 sg13g2_and2_1 _828_ (.A(net130),
    .B(net141),
    .X(_356_));
 sg13g2_nand2_1 _829_ (.Y(_357_),
    .A(net141),
    .B(_331_));
 sg13g2_o21ai_1 _830_ (.B1(_357_),
    .Y(_358_),
    .A1(_331_),
    .A2(_356_));
 sg13g2_nand2_1 _831_ (.Y(_359_),
    .A(net132),
    .B(\lif2.weight[7] ));
 sg13g2_xor2_1 _832_ (.B(_359_),
    .A(_358_),
    .X(_360_));
 sg13g2_nand2b_1 _833_ (.Y(_361_),
    .B(_360_),
    .A_N(_329_));
 sg13g2_xnor2_1 _834_ (.Y(_362_),
    .A(_329_),
    .B(_360_));
 sg13g2_inv_1 _835_ (.Y(_363_),
    .A(_362_));
 sg13g2_nor2_1 _836_ (.A(_340_),
    .B(_363_),
    .Y(_364_));
 sg13g2_nand2_1 _837_ (.Y(_365_),
    .A(_340_),
    .B(_363_));
 sg13g2_nand2b_1 _838_ (.Y(_366_),
    .B(_365_),
    .A_N(_364_));
 sg13g2_nand2_1 _839_ (.Y(_367_),
    .A(_336_),
    .B(_338_));
 sg13g2_xnor2_1 _840_ (.Y(_368_),
    .A(_366_),
    .B(_367_));
 sg13g2_nand2b_1 _841_ (.Y(_369_),
    .B(_368_),
    .A_N(_355_));
 sg13g2_xnor2_1 _842_ (.Y(_370_),
    .A(_355_),
    .B(_368_));
 sg13g2_inv_1 _843_ (.Y(_371_),
    .A(_370_));
 sg13g2_xnor2_1 _844_ (.Y(_372_),
    .A(_354_),
    .B(_370_));
 sg13g2_or2_1 _845_ (.X(_373_),
    .B(_372_),
    .A(_353_));
 sg13g2_a21oi_1 _846_ (.A1(_353_),
    .A2(_372_),
    .Y(_374_),
    .B1(\lif2.spike ));
 sg13g2_and2_1 _847_ (.A(_373_),
    .B(_374_),
    .X(_014_));
 sg13g2_o21ai_1 _848_ (.B1(_369_),
    .Y(_375_),
    .A1(_354_),
    .A2(_371_));
 sg13g2_a21oi_1 _849_ (.A1(_365_),
    .A2(_367_),
    .Y(_376_),
    .B1(_364_));
 sg13g2_o21ai_1 _850_ (.B1(_357_),
    .Y(_377_),
    .A1(_358_),
    .A2(_359_));
 sg13g2_nand2_1 _851_ (.Y(_378_),
    .A(net128),
    .B(net141));
 sg13g2_nand2_1 _852_ (.Y(_379_),
    .A(net130),
    .B(net140));
 sg13g2_xor2_1 _853_ (.B(_379_),
    .A(_378_),
    .X(_380_));
 sg13g2_xnor2_1 _854_ (.Y(_381_),
    .A(_377_),
    .B(_380_));
 sg13g2_xnor2_1 _855_ (.Y(_382_),
    .A(_361_),
    .B(_381_));
 sg13g2_xnor2_1 _856_ (.Y(_383_),
    .A(_376_),
    .B(_382_));
 sg13g2_xnor2_1 _857_ (.Y(_384_),
    .A(_375_),
    .B(_383_));
 sg13g2_and3_1 _858_ (.X(_385_),
    .A(_353_),
    .B(_372_),
    .C(_384_));
 sg13g2_a21oi_1 _859_ (.A1(_353_),
    .A2(_372_),
    .Y(_386_),
    .B1(_384_));
 sg13g2_nor3_1 _860_ (.A(\lif2.spike ),
    .B(_385_),
    .C(_386_),
    .Y(_015_));
 sg13g2_nor3_1 _861_ (.A(net39),
    .B(net36),
    .C(net21),
    .Y(_387_));
 sg13g2_and2_1 _862_ (.A(_443_),
    .B(_387_),
    .X(_388_));
 sg13g2_nor2_1 _863_ (.A(_451_),
    .B(_388_),
    .Y(_389_));
 sg13g2_nand2b_1 _864_ (.Y(_390_),
    .B(\lif1.spike ),
    .A_N(_388_));
 sg13g2_nor3_1 _865_ (.A(net38),
    .B(net33),
    .C(net19),
    .Y(_391_));
 sg13g2_and2_1 _866_ (.A(_441_),
    .B(_391_),
    .X(_392_));
 sg13g2_nor2_2 _867_ (.A(net124),
    .B(_392_),
    .Y(_393_));
 sg13g2_nor2_2 _868_ (.A(_389_),
    .B(_393_),
    .Y(_394_));
 sg13g2_or2_1 _869_ (.X(_395_),
    .B(_393_),
    .A(net123));
 sg13g2_nand2_1 _870_ (.Y(_396_),
    .A(net147),
    .B(net149));
 sg13g2_a21oi_1 _871_ (.A1(net147),
    .A2(net149),
    .Y(_397_),
    .B1(net145));
 sg13g2_nor2b_1 _872_ (.A(_397_),
    .B_N(net143),
    .Y(_398_));
 sg13g2_and2_1 _873_ (.A(net142),
    .B(_398_),
    .X(_399_));
 sg13g2_and2_2 _874_ (.A(net140),
    .B(_399_),
    .X(_400_));
 sg13g2_o21ai_1 _875_ (.B1(_395_),
    .Y(_401_),
    .A1(_390_),
    .A2(_400_));
 sg13g2_o21ai_1 _876_ (.B1(net147),
    .Y(_402_),
    .A1(net149),
    .A2(net154));
 sg13g2_nand2b_2 _877_ (.Y(_403_),
    .B(_402_),
    .A_N(net145));
 sg13g2_nor2_1 _878_ (.A(net143),
    .B(_403_),
    .Y(_404_));
 sg13g2_nor4_2 _879_ (.A(net142),
    .B(net140),
    .C(net143),
    .Y(_405_),
    .D(_403_));
 sg13g2_o21ai_1 _880_ (.B1(_390_),
    .Y(_406_),
    .A1(net154),
    .A2(_405_));
 sg13g2_mux2_1 _881_ (.A0(_406_),
    .A1(net154),
    .S(_401_),
    .X(_023_));
 sg13g2_nor2_2 _882_ (.A(net123),
    .B(_405_),
    .Y(_407_));
 sg13g2_xnor2_1 _883_ (.Y(_408_),
    .A(net149),
    .B(net154));
 sg13g2_nand2b_1 _884_ (.Y(_409_),
    .B(net149),
    .A_N(_400_));
 sg13g2_a221oi_1 _885_ (.B2(net123),
    .C1(_394_),
    .B1(_409_),
    .A1(_407_),
    .Y(_410_),
    .A2(_408_));
 sg13g2_a21o_1 _886_ (.A2(_394_),
    .A1(net17),
    .B1(_410_),
    .X(_024_));
 sg13g2_xor2_1 _887_ (.B(net149),
    .A(net147),
    .X(_411_));
 sg13g2_o21ai_1 _888_ (.B1(net123),
    .Y(_412_),
    .A1(_400_),
    .A2(_411_));
 sg13g2_nor3_1 _889_ (.A(net147),
    .B(net149),
    .C(net154),
    .Y(_413_));
 sg13g2_and2_1 _890_ (.A(_393_),
    .B(_407_),
    .X(_414_));
 sg13g2_a22oi_1 _891_ (.Y(_415_),
    .B1(_402_),
    .B2(_414_),
    .A2(_394_),
    .A1(net147));
 sg13g2_o21ai_1 _892_ (.B1(_412_),
    .Y(_025_),
    .A1(_413_),
    .A2(_415_));
 sg13g2_a21oi_1 _893_ (.A1(_393_),
    .A2(_402_),
    .Y(_416_),
    .B1(net123));
 sg13g2_nand2_1 _894_ (.Y(_417_),
    .A(net145),
    .B(_416_));
 sg13g2_nand2_1 _895_ (.Y(_418_),
    .A(_016_),
    .B(_396_));
 sg13g2_xnor2_1 _896_ (.Y(_419_),
    .A(net44),
    .B(_396_));
 sg13g2_o21ai_1 _897_ (.B1(net123),
    .Y(_420_),
    .A1(_400_),
    .A2(_419_));
 sg13g2_nand2b_1 _898_ (.Y(_421_),
    .B(_414_),
    .A_N(_403_));
 sg13g2_nand3_1 _899_ (.B(_420_),
    .C(_421_),
    .A(_417_),
    .Y(_026_));
 sg13g2_xnor2_1 _900_ (.Y(_422_),
    .A(net143),
    .B(_403_));
 sg13g2_xor2_1 _901_ (.B(_418_),
    .A(net143),
    .X(_423_));
 sg13g2_o21ai_1 _902_ (.B1(net123),
    .Y(_424_),
    .A1(_400_),
    .A2(_423_));
 sg13g2_o21ai_1 _903_ (.B1(_424_),
    .Y(_425_),
    .A1(net29),
    .A2(_395_));
 sg13g2_a21oi_1 _904_ (.A1(_414_),
    .A2(_422_),
    .Y(_027_),
    .B1(net30));
 sg13g2_xor2_1 _905_ (.B(_404_),
    .A(net142),
    .X(_426_));
 sg13g2_nand2b_1 _906_ (.Y(_427_),
    .B(_399_),
    .A_N(net140));
 sg13g2_o21ai_1 _907_ (.B1(_427_),
    .Y(_428_),
    .A1(net142),
    .A2(_398_));
 sg13g2_o21ai_1 _908_ (.B1(_395_),
    .Y(_429_),
    .A1(_390_),
    .A2(_428_));
 sg13g2_a21oi_1 _909_ (.A1(_407_),
    .A2(_426_),
    .Y(_430_),
    .B1(_429_));
 sg13g2_a21o_1 _910_ (.A2(_394_),
    .A1(net18),
    .B1(_430_),
    .X(_028_));
 sg13g2_a21oi_1 _911_ (.A1(net123),
    .A2(_399_),
    .Y(_431_),
    .B1(net140));
 sg13g2_nor4_1 _912_ (.A(net142),
    .B(net143),
    .C(_401_),
    .D(_403_),
    .Y(_432_));
 sg13g2_nor2_1 _913_ (.A(_431_),
    .B(_432_),
    .Y(_029_));
 sg13g2_nor3_1 _914_ (.A(net21),
    .B(\lif2.spike ),
    .C(_388_),
    .Y(_030_));
 sg13g2_xor2_1 _915_ (.B(net21),
    .A(net36),
    .X(_433_));
 sg13g2_o21ai_1 _916_ (.B1(net124),
    .Y(_031_),
    .A1(_388_),
    .A2(_433_));
 sg13g2_o21ai_1 _917_ (.B1(net39),
    .Y(_434_),
    .A1(net36),
    .A2(net21));
 sg13g2_nor2b_1 _918_ (.A(_387_),
    .B_N(_434_),
    .Y(_435_));
 sg13g2_nor3_1 _919_ (.A(\lif2.spike ),
    .B(_388_),
    .C(_435_),
    .Y(_032_));
 sg13g2_o21ai_1 _920_ (.B1(net124),
    .Y(_033_),
    .A1(_443_),
    .A2(_387_));
 sg13g2_nor3_1 _921_ (.A(net19),
    .B(\lif1.spike ),
    .C(_392_),
    .Y(_034_));
 sg13g2_xor2_1 _922_ (.B(net19),
    .A(net33),
    .X(_436_));
 sg13g2_o21ai_1 _923_ (.B1(_451_),
    .Y(_035_),
    .A1(_392_),
    .A2(_436_));
 sg13g2_o21ai_1 _924_ (.B1(net38),
    .Y(_437_),
    .A1(net33),
    .A2(net19));
 sg13g2_nor2b_1 _925_ (.A(_391_),
    .B_N(_437_),
    .Y(_438_));
 sg13g2_nor3_1 _926_ (.A(\lif1.spike ),
    .B(_392_),
    .C(_438_),
    .Y(_036_));
 sg13g2_o21ai_1 _927_ (.B1(_451_),
    .Y(_037_),
    .A1(_441_),
    .A2(_391_));
 sg13g2_nor2_1 _928_ (.A(_401_),
    .B(_407_),
    .Y(_439_));
 sg13g2_mux2_1 _929_ (.A0(net27),
    .A1(net142),
    .S(_439_),
    .X(_038_));
 sg13g2_dfrbp_1 _930_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net155),
    .D(_023_),
    .Q_N(_465_),
    .Q(\lif2.weight[1] ));
 sg13g2_dfrbp_1 _931_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net155),
    .D(_024_),
    .Q_N(\lif2.weight[2] ),
    .Q(_020_));
 sg13g2_dfrbp_1 _932_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net155),
    .D(net53),
    .Q_N(_464_),
    .Q(\lif2.weight[3] ));
 sg13g2_dfrbp_1 _933_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net155),
    .D(net45),
    .Q_N(_016_),
    .Q(\lif2.weight[4] ));
 sg13g2_dfrbp_1 _934_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net155),
    .D(_027_),
    .Q_N(\lif2.weight[5] ),
    .Q(_021_));
 sg13g2_dfrbp_1 _935_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net155),
    .D(_028_),
    .Q_N(\lif2.weight[6] ),
    .Q(_022_));
 sg13g2_dfrbp_1 _936_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net155),
    .D(net49),
    .Q_N(_466_),
    .Q(\lif2.weight[7] ));
 sg13g2_dfrbp_1 _937_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net160),
    .D(_000_),
    .Q_N(_467_),
    .Q(\lif1.state[0] ));
 sg13g2_dfrbp_1 _938_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net160),
    .D(_001_),
    .Q_N(_468_),
    .Q(\lif1.state[1] ));
 sg13g2_dfrbp_1 _939_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net159),
    .D(_002_),
    .Q_N(_469_),
    .Q(\lif1.state[2] ));
 sg13g2_dfrbp_1 _940_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net159),
    .D(_003_),
    .Q_N(_470_),
    .Q(\lif1.state[3] ));
 sg13g2_dfrbp_1 _941_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net159),
    .D(_004_),
    .Q_N(_471_),
    .Q(\lif1.state[4] ));
 sg13g2_dfrbp_1 _942_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net159),
    .D(_005_),
    .Q_N(_472_),
    .Q(\lif1.state[5] ));
 sg13g2_dfrbp_1 _943_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net159),
    .D(_006_),
    .Q_N(_473_),
    .Q(\lif1.state[6] ));
 sg13g2_dfrbp_1 _944_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net159),
    .D(_007_),
    .Q_N(_463_),
    .Q(\lif1.state[7] ));
 sg13g2_dfrbp_1 _945_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net156),
    .D(net22),
    .Q_N(_462_),
    .Q(\stdp1.post_counter[0] ));
 sg13g2_dfrbp_1 _946_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net156),
    .D(net37),
    .Q_N(_461_),
    .Q(\stdp1.post_counter[1] ));
 sg13g2_dfrbp_1 _947_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net156),
    .D(_032_),
    .Q_N(_460_),
    .Q(\stdp1.post_counter[2] ));
 sg13g2_dfrbp_1 _948_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net156),
    .D(net24),
    .Q_N(_459_),
    .Q(\stdp1.post_counter[3] ));
 sg13g2_dfrbp_1 _949_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net159),
    .D(net20),
    .Q_N(_458_),
    .Q(\stdp1.pre_counter[0] ));
 sg13g2_dfrbp_1 _950_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net157),
    .D(net34),
    .Q_N(_457_),
    .Q(\stdp1.pre_counter[1] ));
 sg13g2_dfrbp_1 _951_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net157),
    .D(_036_),
    .Q_N(_456_),
    .Q(\stdp1.pre_counter[2] ));
 sg13g2_dfrbp_1 _952_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net157),
    .D(net26),
    .Q_N(_455_),
    .Q(\stdp1.pre_counter[3] ));
 sg13g2_dfrbp_1 _953_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net155),
    .D(net28),
    .Q_N(_474_),
    .Q(\lif2.weight[0] ));
 sg13g2_dfrbp_1 _954_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net159),
    .D(_008_),
    .Q_N(_475_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _955_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net157),
    .D(net41),
    .Q_N(_476_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _956_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net157),
    .D(_010_),
    .Q_N(_477_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _957_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net157),
    .D(net32),
    .Q_N(_478_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _958_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net158),
    .D(_012_),
    .Q_N(_479_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _959_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net158),
    .D(net43),
    .Q_N(_017_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _960_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net157),
    .D(_014_),
    .Q_N(_018_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _961_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net157),
    .D(_015_),
    .Q_N(_019_),
    .Q(uo_out[7]));
 sg13g2_tiehi tt_um_two_lif_stdp_10 (.L_HI(net10));
 sg13g2_tiehi tt_um_two_lif_stdp_11 (.L_HI(net11));
 sg13g2_tiehi tt_um_two_lif_stdp_12 (.L_HI(net12));
 sg13g2_tiehi tt_um_two_lif_stdp_13 (.L_HI(net13));
 sg13g2_tiehi tt_um_two_lif_stdp_14 (.L_HI(net14));
 sg13g2_tiehi tt_um_two_lif_stdp_15 (.L_HI(net15));
 sg13g2_tiehi tt_um_two_lif_stdp_16 (.L_HI(net16));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _970_ (.A(\lif2.weight[0] ),
    .X(uio_out[0]));
 sg13g2_buf_1 _971_ (.A(net154),
    .X(uio_out[1]));
 sg13g2_buf_1 _972_ (.A(net149),
    .X(uio_out[2]));
 sg13g2_buf_1 _973_ (.A(net147),
    .X(uio_out[3]));
 sg13g2_buf_1 _974_ (.A(net145),
    .X(uio_out[4]));
 sg13g2_buf_1 _975_ (.A(net143),
    .X(uio_out[5]));
 sg13g2_buf_1 _976_ (.A(\lif2.spike ),
    .X(uio_out[6]));
 sg13g2_buf_1 _977_ (.A(\lif1.spike ),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout123 (.A(_389_),
    .X(net123));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(_447_));
 sg13g2_buf_2 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(net127),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(\lif2.weight[0] ),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(\lif1.state[7] ),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(\lif1.state[6] ),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(\lif1.state[5] ),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(\lif1.state[4] ));
 sg13g2_buf_2 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(\lif1.state[3] ),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(net138),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(\lif1.state[2] ),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(\lif1.state[1] ),
    .X(net139));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(\lif2.weight[7] ));
 sg13g2_buf_2 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net48));
 sg13g2_buf_2 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(\lif2.weight[5] ));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(\lif2.weight[4] ));
 sg13g2_buf_2 fanout146 (.A(\lif2.weight[4] ),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(\lif2.weight[3] ),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(\lif2.weight[3] ));
 sg13g2_buf_2 fanout149 (.A(net52),
    .X(net149));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(\lif2.weight[2] ));
 sg13g2_buf_2 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net46),
    .X(net154));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(net158));
 sg13g2_buf_2 fanout156 (.A(net158),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(net158));
 sg13g2_buf_2 fanout158 (.A(net160),
    .X(net158));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(net160));
 sg13g2_buf_2 fanout160 (.A(rst_n),
    .X(net160));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tiehi tt_um_two_lif_stdp_9 (.L_HI(net9));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_020_),
    .X(net17));
 sg13g2_dlygate4sd3_1 hold2 (.A(_022_),
    .X(net18));
 sg13g2_dlygate4sd3_1 hold3 (.A(\stdp1.pre_counter[0] ),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold4 (.A(_034_),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold5 (.A(\stdp1.post_counter[0] ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold6 (.A(_030_),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold7 (.A(\stdp1.post_counter[3] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold8 (.A(_033_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold9 (.A(\stdp1.pre_counter[3] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold10 (.A(_037_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold11 (.A(\lif2.weight[0] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold12 (.A(_038_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold13 (.A(_021_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold14 (.A(_425_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold15 (.A(_017_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold16 (.A(_011_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold17 (.A(\stdp1.pre_counter[1] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold18 (.A(_035_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold19 (.A(uo_out[2]),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold20 (.A(\stdp1.post_counter[1] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold21 (.A(_031_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold22 (.A(\stdp1.pre_counter[2] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold23 (.A(\stdp1.post_counter[2] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold24 (.A(uo_out[3]),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold25 (.A(_009_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold26 (.A(_019_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold27 (.A(_013_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold28 (.A(_016_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold29 (.A(_026_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold30 (.A(\lif2.weight[1] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold31 (.A(_018_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold32 (.A(\lif2.weight[6] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold33 (.A(_029_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold34 (.A(\lif1.state[7] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold35 (.A(uo_out[4]),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold36 (.A(\lif2.weight[2] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold37 (.A(_025_),
    .X(net53));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_fill_1 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_decap_4 FILLER_21_237 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_fill_2 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_276 ();
 sg13g2_fill_1 FILLER_21_283 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_4 FILLER_21_298 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_fill_1 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_269 ();
 sg13g2_decap_4 FILLER_22_300 ();
 sg13g2_decap_4 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_4 FILLER_23_175 ();
 sg13g2_fill_2 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_230 ();
 sg13g2_decap_4 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_267 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_decap_4 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_168 ();
 sg13g2_fill_2 FILLER_24_178 ();
 sg13g2_decap_4 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_220 ();
 sg13g2_decap_8 FILLER_24_239 ();
 sg13g2_decap_8 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_253 ();
 sg13g2_fill_2 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_fill_2 FILLER_24_302 ();
 sg13g2_fill_1 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_344 ();
 sg13g2_fill_2 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_4 FILLER_24_383 ();
 sg13g2_fill_1 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_decap_4 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_decap_8 FILLER_25_129 ();
 sg13g2_decap_4 FILLER_25_136 ();
 sg13g2_fill_1 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_149 ();
 sg13g2_fill_2 FILLER_25_156 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_decap_8 FILLER_25_216 ();
 sg13g2_fill_2 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_253 ();
 sg13g2_decap_8 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_289 ();
 sg13g2_decap_4 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_300 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_322 ();
 sg13g2_decap_4 FILLER_25_344 ();
 sg13g2_fill_2 FILLER_25_348 ();
 sg13g2_fill_2 FILLER_25_358 ();
 sg13g2_fill_1 FILLER_25_360 ();
 sg13g2_fill_2 FILLER_25_377 ();
 sg13g2_fill_1 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_fill_1 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_139 ();
 sg13g2_decap_8 FILLER_26_146 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_172 ();
 sg13g2_decap_4 FILLER_26_187 ();
 sg13g2_fill_2 FILLER_26_195 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_209 ();
 sg13g2_decap_4 FILLER_26_226 ();
 sg13g2_fill_2 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_fill_1 FILLER_26_279 ();
 sg13g2_fill_1 FILLER_26_292 ();
 sg13g2_fill_2 FILLER_26_305 ();
 sg13g2_fill_1 FILLER_26_307 ();
 sg13g2_decap_4 FILLER_26_311 ();
 sg13g2_fill_1 FILLER_26_331 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_353 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_fill_2 FILLER_26_383 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_84 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_1 FILLER_27_111 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_fill_2 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_2 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_decap_8 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_274 ();
 sg13g2_fill_1 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_290 ();
 sg13g2_decap_4 FILLER_27_296 ();
 sg13g2_fill_2 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_324 ();
 sg13g2_decap_4 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_4 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_351 ();
 sg13g2_decap_4 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_4 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_67 ();
 sg13g2_fill_2 FILLER_28_103 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_decap_4 FILLER_28_186 ();
 sg13g2_fill_1 FILLER_28_190 ();
 sg13g2_decap_4 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_decap_8 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_232 ();
 sg13g2_decap_4 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_4 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_333 ();
 sg13g2_fill_1 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_387 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_4 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_81 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_decap_8 FILLER_29_176 ();
 sg13g2_decap_4 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_decap_8 FILLER_29_204 ();
 sg13g2_decap_4 FILLER_29_223 ();
 sg13g2_fill_1 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_254 ();
 sg13g2_decap_4 FILLER_29_261 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_decap_4 FILLER_29_278 ();
 sg13g2_decap_4 FILLER_29_287 ();
 sg13g2_fill_1 FILLER_29_291 ();
 sg13g2_decap_4 FILLER_29_309 ();
 sg13g2_fill_2 FILLER_29_313 ();
 sg13g2_decap_4 FILLER_29_334 ();
 sg13g2_decap_4 FILLER_29_358 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_128 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_decap_4 FILLER_30_202 ();
 sg13g2_decap_8 FILLER_30_215 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_262 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_decap_4 FILLER_30_333 ();
 sg13g2_fill_1 FILLER_30_337 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_4 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_decap_4 FILLER_31_110 ();
 sg13g2_decap_4 FILLER_31_125 ();
 sg13g2_fill_2 FILLER_31_179 ();
 sg13g2_fill_1 FILLER_31_181 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_224 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_fill_2 FILLER_31_270 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_287 ();
 sg13g2_decap_4 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_298 ();
 sg13g2_decap_4 FILLER_31_304 ();
 sg13g2_fill_2 FILLER_31_308 ();
 sg13g2_fill_1 FILLER_31_344 ();
 sg13g2_decap_4 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_decap_4 FILLER_31_383 ();
 sg13g2_fill_1 FILLER_31_387 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_4 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_81 ();
 sg13g2_fill_1 FILLER_32_113 ();
 sg13g2_decap_4 FILLER_32_132 ();
 sg13g2_decap_4 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_fill_2 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_265 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_310 ();
 sg13g2_decap_4 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_decap_4 FILLER_32_354 ();
 sg13g2_decap_4 FILLER_32_382 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_fill_1 FILLER_32_393 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_4 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_100 ();
 sg13g2_fill_1 FILLER_33_172 ();
 sg13g2_fill_2 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_decap_8 FILLER_33_278 ();
 sg13g2_fill_2 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_292 ();
 sg13g2_fill_2 FILLER_33_297 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_decap_4 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_359 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_fill_2 FILLER_33_379 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_4 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_95 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_fill_1 FILLER_34_220 ();
 sg13g2_decap_4 FILLER_34_240 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_2 FILLER_34_290 ();
 sg13g2_decap_4 FILLER_34_309 ();
 sg13g2_fill_1 FILLER_34_313 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_340 ();
 sg13g2_fill_2 FILLER_34_347 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_4 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_124 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_1 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_160 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_fill_1 FILLER_35_168 ();
 sg13g2_fill_2 FILLER_35_178 ();
 sg13g2_decap_4 FILLER_35_258 ();
 sg13g2_decap_4 FILLER_35_276 ();
 sg13g2_fill_1 FILLER_35_352 ();
 sg13g2_fill_1 FILLER_35_361 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_133 ();
 sg13g2_fill_1 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_193 ();
 sg13g2_fill_1 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_fill_1 FILLER_36_262 ();
 sg13g2_fill_1 FILLER_36_289 ();
 sg13g2_fill_2 FILLER_36_319 ();
 sg13g2_fill_2 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_343 ();
 sg13g2_fill_1 FILLER_36_345 ();
 sg13g2_decap_4 FILLER_36_354 ();
 sg13g2_decap_4 FILLER_36_364 ();
 sg13g2_decap_4 FILLER_36_383 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_1 FILLER_37_322 ();
 sg13g2_fill_1 FILLER_37_354 ();
 sg13g2_fill_1 FILLER_37_384 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_149 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_361 ();
 sg13g2_fill_2 FILLER_38_382 ();
 sg13g2_fill_1 FILLER_38_384 ();
 sg13g2_fill_2 FILLER_38_389 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
endmodule

module tt_um_wokwi_group_3 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire net237;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire \proj_10.net10 ;
 wire \proj_10.net11 ;
 wire \proj_10.net12 ;
 wire \proj_10.net13 ;
 wire \proj_10.net9 ;
 wire \proj_12.net10 ;
 wire \proj_12.net11 ;
 wire \proj_12.net12 ;
 wire \proj_12.net13 ;
 wire \proj_12.net18 ;
 wire \proj_12.net19 ;
 wire \proj_12.net20 ;
 wire \proj_12.net21 ;
 wire \proj_12.net22 ;
 wire \proj_12.net23 ;
 wire \proj_12.net24 ;
 wire \proj_12.net25 ;
 wire \proj_12.net26 ;
 wire \proj_12.net27 ;
 wire \proj_12.net28 ;
 wire \proj_12.net29 ;
 wire \proj_12.net9 ;
 wire \proj_13.net12 ;
 wire \proj_13.net13 ;
 wire \proj_13.net7 ;
 wire \proj_13.net8 ;
 wire \proj_14.net100 ;
 wire \proj_14.net101 ;
 wire \proj_14.net102 ;
 wire \proj_14.net104 ;
 wire \proj_14.net105 ;
 wire \proj_14.net106 ;
 wire \proj_14.net108 ;
 wire \proj_14.net11 ;
 wire \proj_14.net110 ;
 wire \proj_14.net111 ;
 wire \proj_14.net112 ;
 wire \proj_14.net114 ;
 wire \proj_14.net115 ;
 wire \proj_14.net116 ;
 wire \proj_14.net117 ;
 wire \proj_14.net119 ;
 wire \proj_14.net12 ;
 wire \proj_14.net120 ;
 wire \proj_14.net121 ;
 wire \proj_14.net122 ;
 wire \proj_14.net124 ;
 wire \proj_14.net125 ;
 wire \proj_14.net126 ;
 wire \proj_14.net127 ;
 wire \proj_14.net129 ;
 wire \proj_14.net13 ;
 wire \proj_14.net130 ;
 wire \proj_14.net131 ;
 wire \proj_14.net132 ;
 wire \proj_14.net133 ;
 wire \proj_14.net135 ;
 wire \proj_14.net136 ;
 wire \proj_14.net137 ;
 wire \proj_14.net138 ;
 wire \proj_14.net14 ;
 wire \proj_14.net140 ;
 wire \proj_14.net141 ;
 wire \proj_14.net142 ;
 wire \proj_14.net143 ;
 wire \proj_14.net145 ;
 wire \proj_14.net146 ;
 wire \proj_14.net147 ;
 wire \proj_14.net148 ;
 wire \proj_14.net15 ;
 wire \proj_14.net150 ;
 wire \proj_14.net151 ;
 wire \proj_14.net152 ;
 wire \proj_14.net153 ;
 wire \proj_14.net155 ;
 wire \proj_14.net156 ;
 wire \proj_14.net157 ;
 wire \proj_14.net158 ;
 wire \proj_14.net16 ;
 wire \proj_14.net160 ;
 wire \proj_14.net161 ;
 wire \proj_14.net162 ;
 wire \proj_14.net163 ;
 wire \proj_14.net165 ;
 wire \proj_14.net166 ;
 wire \proj_14.net167 ;
 wire \proj_14.net168 ;
 wire \proj_14.net17 ;
 wire \proj_14.net170 ;
 wire \proj_14.net171 ;
 wire \proj_14.net172 ;
 wire \proj_14.net173 ;
 wire \proj_14.net175 ;
 wire \proj_14.net176 ;
 wire \proj_14.net177 ;
 wire \proj_14.net178 ;
 wire \proj_14.net180 ;
 wire \proj_14.net181 ;
 wire \proj_14.net182 ;
 wire \proj_14.net183 ;
 wire \proj_14.net184 ;
 wire \proj_14.net185 ;
 wire \proj_14.net186 ;
 wire \proj_14.net187 ;
 wire \proj_14.net188 ;
 wire \proj_14.net189 ;
 wire \proj_14.net190 ;
 wire \proj_14.net191 ;
 wire \proj_14.net192 ;
 wire \proj_14.net193 ;
 wire \proj_14.net194 ;
 wire \proj_14.net195 ;
 wire \proj_14.net196 ;
 wire \proj_14.net197 ;
 wire \proj_14.net198 ;
 wire \proj_14.net199 ;
 wire \proj_14.net200 ;
 wire \proj_14.net201 ;
 wire \proj_14.net202 ;
 wire \proj_14.net203 ;
 wire \proj_14.net204 ;
 wire \proj_14.net205 ;
 wire \proj_14.net206 ;
 wire \proj_14.net207 ;
 wire \proj_14.net209 ;
 wire \proj_14.net210 ;
 wire \proj_14.net211 ;
 wire \proj_14.net212 ;
 wire \proj_14.net214 ;
 wire \proj_14.net215 ;
 wire \proj_14.net216 ;
 wire \proj_14.net217 ;
 wire \proj_14.net218 ;
 wire \proj_14.net219 ;
 wire \proj_14.net220 ;
 wire \proj_14.net221 ;
 wire \proj_14.net222 ;
 wire \proj_14.net223 ;
 wire \proj_14.net224 ;
 wire \proj_14.net226 ;
 wire \proj_14.net227 ;
 wire \proj_14.net228 ;
 wire \proj_14.net229 ;
 wire \proj_14.net23 ;
 wire \proj_14.net231 ;
 wire \proj_14.net232 ;
 wire \proj_14.net233 ;
 wire \proj_14.net234 ;
 wire \proj_14.net235 ;
 wire \proj_14.net236 ;
 wire \proj_14.net237 ;
 wire \proj_14.net238 ;
 wire \proj_14.net239 ;
 wire \proj_14.net240 ;
 wire \proj_14.net241 ;
 wire \proj_14.net242 ;
 wire \proj_14.net243 ;
 wire \proj_14.net244 ;
 wire \proj_14.net245 ;
 wire \proj_14.net246 ;
 wire \proj_14.net247 ;
 wire \proj_14.net248 ;
 wire \proj_14.net249 ;
 wire \proj_14.net25 ;
 wire \proj_14.net250 ;
 wire \proj_14.net251 ;
 wire \proj_14.net252 ;
 wire \proj_14.net253 ;
 wire \proj_14.net254 ;
 wire \proj_14.net255 ;
 wire \proj_14.net256 ;
 wire \proj_14.net257 ;
 wire \proj_14.net258 ;
 wire \proj_14.net259 ;
 wire \proj_14.net26 ;
 wire \proj_14.net260 ;
 wire \proj_14.net261 ;
 wire \proj_14.net262 ;
 wire \proj_14.net263 ;
 wire \proj_14.net264 ;
 wire \proj_14.net265 ;
 wire \proj_14.net266 ;
 wire \proj_14.net267 ;
 wire \proj_14.net268 ;
 wire \proj_14.net269 ;
 wire \proj_14.net27 ;
 wire \proj_14.net270 ;
 wire \proj_14.net271 ;
 wire \proj_14.net272 ;
 wire \proj_14.net273 ;
 wire \proj_14.net274 ;
 wire \proj_14.net275 ;
 wire \proj_14.net276 ;
 wire \proj_14.net277 ;
 wire \proj_14.net278 ;
 wire \proj_14.net279 ;
 wire \proj_14.net28 ;
 wire \proj_14.net280 ;
 wire \proj_14.net281 ;
 wire \proj_14.net282 ;
 wire \proj_14.net283 ;
 wire \proj_14.net284 ;
 wire \proj_14.net285 ;
 wire \proj_14.net286 ;
 wire \proj_14.net287 ;
 wire \proj_14.net288 ;
 wire \proj_14.net289 ;
 wire \proj_14.net29 ;
 wire \proj_14.net30 ;
 wire \proj_14.net31 ;
 wire \proj_14.net32 ;
 wire \proj_14.net33 ;
 wire \proj_14.net34 ;
 wire \proj_14.net36 ;
 wire \proj_14.net37 ;
 wire \proj_14.net38 ;
 wire \proj_14.net39 ;
 wire \proj_14.net40 ;
 wire \proj_14.net41 ;
 wire \proj_14.net42 ;
 wire \proj_14.net43 ;
 wire \proj_14.net44 ;
 wire \proj_14.net45 ;
 wire \proj_14.net46 ;
 wire \proj_14.net47 ;
 wire \proj_14.net48 ;
 wire \proj_14.net50 ;
 wire \proj_14.net51 ;
 wire \proj_14.net52 ;
 wire \proj_14.net53 ;
 wire \proj_14.net54 ;
 wire \proj_14.net55 ;
 wire \proj_14.net56 ;
 wire \proj_14.net57 ;
 wire \proj_14.net58 ;
 wire \proj_14.net59 ;
 wire \proj_14.net60 ;
 wire \proj_14.net61 ;
 wire \proj_14.net62 ;
 wire \proj_14.net63 ;
 wire \proj_14.net64 ;
 wire \proj_14.net65 ;
 wire \proj_14.net66 ;
 wire \proj_14.net67 ;
 wire \proj_14.net68 ;
 wire \proj_14.net69 ;
 wire \proj_14.net70 ;
 wire \proj_14.net71 ;
 wire \proj_14.net72 ;
 wire \proj_14.net73 ;
 wire \proj_14.net74 ;
 wire \proj_14.net75 ;
 wire \proj_14.net76 ;
 wire \proj_14.net77 ;
 wire \proj_14.net78 ;
 wire \proj_14.net79 ;
 wire \proj_14.net80 ;
 wire \proj_14.net81 ;
 wire \proj_14.net82 ;
 wire \proj_14.net83 ;
 wire \proj_14.net84 ;
 wire \proj_14.net85 ;
 wire \proj_14.net86 ;
 wire \proj_14.net87 ;
 wire \proj_14.net88 ;
 wire \proj_14.net89 ;
 wire \proj_14.net90 ;
 wire \proj_14.net91 ;
 wire \proj_14.net92 ;
 wire \proj_14.net93 ;
 wire \proj_14.net94 ;
 wire \proj_14.net95 ;
 wire \proj_14.net96 ;
 wire \proj_14.net97 ;
 wire \proj_14.net98 ;
 wire \proj_14.net99 ;
 wire \proj__0.net10 ;
 wire \proj__0.net11 ;
 wire \proj__0.net9 ;
 wire \proj__1.net10 ;
 wire \proj__1.net16 ;
 wire \proj__1.net17 ;
 wire \proj__1.net18 ;
 wire \proj__1.net19 ;
 wire \proj__1.net20 ;
 wire \proj__1.net21 ;
 wire \proj__1.net22 ;
 wire \proj__1.net23 ;
 wire \proj__1.net24 ;
 wire \proj__1.net9 ;
 wire \proj__2.net10 ;
 wire \proj__2.net11 ;
 wire \proj__2.net12 ;
 wire \proj__2.net9 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net13 ;
 wire \proj__3.net3 ;
 wire \proj__3.net4 ;
 wire \proj__3.net5 ;
 wire \proj__4.net11 ;
 wire \proj__4.net12 ;
 wire \proj__4.net13 ;
 wire \proj__4.net14 ;
 wire \proj__4.net15 ;
 wire \proj__4.net16 ;
 wire \proj__4.net17 ;
 wire \proj__4.net18 ;
 wire \proj__5.net10 ;
 wire \proj__5.net11 ;
 wire \proj__5.net12 ;
 wire \proj__5.net9 ;
 wire \proj__6.net10 ;
 wire \proj__6.net9 ;
 wire \proj__7.net14 ;
 wire \proj__7.net15 ;
 wire \proj__7.net5 ;
 wire \proj__7.net6 ;
 wire \proj__7.net7 ;
 wire \proj__7.net8 ;
 wire \proj__8.net7 ;
 wire \proj__9.net11 ;
 wire \proj__9.net12 ;
 wire \proj__9.net13 ;
 wire \proj__9.net14 ;
 wire \proj__9.net15 ;
 wire \proj__9.net17 ;
 wire \proj__9.net5 ;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire \proj_10.nand1/b ;
 wire net238;
 wire \proj_13.flop1/notq ;
 wire net239;
 wire \proj_13.flop2/notq ;
 wire net240;
 wire \proj_13.flop3/notq ;
 wire \proj_14.flop1/_0_ ;
 wire \proj_14.flop1/_1_ ;
 wire net147;
 wire net148;
 wire \proj_14.flop10/_0_ ;
 wire \proj_14.flop10/_1_ ;
 wire net149;
 wire net150;
 wire \proj_14.flop11/_0_ ;
 wire \proj_14.flop11/_1_ ;
 wire net151;
 wire net152;
 wire \proj_14.flop12/_0_ ;
 wire \proj_14.flop12/_1_ ;
 wire net153;
 wire net154;
 wire \proj_14.flop13/_0_ ;
 wire \proj_14.flop13/_1_ ;
 wire net155;
 wire net156;
 wire \proj_14.flop14/_0_ ;
 wire \proj_14.flop14/_1_ ;
 wire net157;
 wire net158;
 wire \proj_14.flop15/_0_ ;
 wire \proj_14.flop15/_1_ ;
 wire net159;
 wire net160;
 wire \proj_14.flop16/_0_ ;
 wire \proj_14.flop16/_1_ ;
 wire net161;
 wire net162;
 wire \proj_14.flop17/_0_ ;
 wire \proj_14.flop17/_1_ ;
 wire net163;
 wire net164;
 wire \proj_14.flop18/_0_ ;
 wire \proj_14.flop18/_1_ ;
 wire net165;
 wire net166;
 wire \proj_14.flop19/_0_ ;
 wire \proj_14.flop19/_1_ ;
 wire net167;
 wire net168;
 wire \proj_14.flop2/_0_ ;
 wire \proj_14.flop2/_1_ ;
 wire net169;
 wire net170;
 wire \proj_14.flop20/_0_ ;
 wire \proj_14.flop20/_1_ ;
 wire net171;
 wire net172;
 wire \proj_14.flop21/_0_ ;
 wire \proj_14.flop21/_1_ ;
 wire net173;
 wire net174;
 wire \proj_14.flop22/_0_ ;
 wire \proj_14.flop22/_1_ ;
 wire net175;
 wire net176;
 wire \proj_14.flop23/_0_ ;
 wire \proj_14.flop23/_1_ ;
 wire net177;
 wire net178;
 wire \proj_14.flop24/_0_ ;
 wire \proj_14.flop24/_1_ ;
 wire net179;
 wire net180;
 wire \proj_14.flop25/_0_ ;
 wire \proj_14.flop25/_1_ ;
 wire net181;
 wire net182;
 wire \proj_14.flop25/notq ;
 wire \proj_14.flop26/_0_ ;
 wire \proj_14.flop26/_1_ ;
 wire net183;
 wire net184;
 wire \proj_14.flop26/notq ;
 wire \proj_14.flop27/_0_ ;
 wire \proj_14.flop27/_1_ ;
 wire net185;
 wire net186;
 wire \proj_14.flop27/q ;
 wire net241;
 wire \proj_14.flop28/notq ;
 wire \proj_14.flop29/_0_ ;
 wire \proj_14.flop29/_1_ ;
 wire net187;
 wire net188;
 wire \proj_14.flop3/_0_ ;
 wire \proj_14.flop3/_1_ ;
 wire net189;
 wire net190;
 wire \proj_14.flop30/_0_ ;
 wire \proj_14.flop30/_1_ ;
 wire net191;
 wire net192;
 wire \proj_14.flop31/_0_ ;
 wire \proj_14.flop31/_1_ ;
 wire net193;
 wire net194;
 wire \proj_14.flop31/notq ;
 wire \proj_14.flop32/_0_ ;
 wire \proj_14.flop32/_1_ ;
 wire net195;
 wire net196;
 wire \proj_14.flop32/notq ;
 wire \proj_14.flop33/_0_ ;
 wire \proj_14.flop33/_1_ ;
 wire net197;
 wire net198;
 wire \proj_14.flop33/notq ;
 wire \proj_14.flop34/_0_ ;
 wire \proj_14.flop34/_1_ ;
 wire net199;
 wire net200;
 wire \proj_14.flop34/notq ;
 wire \proj_14.flop35/_0_ ;
 wire \proj_14.flop35/_1_ ;
 wire net201;
 wire net202;
 wire \proj_14.flop35/notq ;
 wire \proj_14.flop36/_0_ ;
 wire \proj_14.flop36/_1_ ;
 wire net203;
 wire net204;
 wire \proj_14.flop36/notq ;
 wire \proj_14.flop37/_0_ ;
 wire \proj_14.flop37/_1_ ;
 wire net205;
 wire net206;
 wire \proj_14.flop37/notq ;
 wire \proj_14.flop4/_0_ ;
 wire \proj_14.flop4/_1_ ;
 wire net207;
 wire net208;
 wire net242;
 wire \proj_14.flop46/notq ;
 wire net243;
 wire \proj_14.flop47/notq ;
 wire net244;
 wire \proj_14.flop48/notq ;
 wire net245;
 wire \proj_14.flop49/notq ;
 wire \proj_14.flop5/_0_ ;
 wire \proj_14.flop5/_1_ ;
 wire net209;
 wire net210;
 wire net246;
 wire \proj_14.flop50/notq ;
 wire net247;
 wire \proj_14.flop51/notq ;
 wire net248;
 wire \proj_14.flop52/notq ;
 wire net249;
 wire \proj_14.flop53/notq ;
 wire net250;
 wire \proj_14.flop54/notq ;
 wire net251;
 wire \proj_14.flop55/notq ;
 wire net252;
 wire \proj_14.flop56/notq ;
 wire \proj_14.flop6/_0_ ;
 wire \proj_14.flop6/_1_ ;
 wire net211;
 wire net212;
 wire \proj_14.flop7/_0_ ;
 wire \proj_14.flop7/_1_ ;
 wire net213;
 wire net214;
 wire \proj_14.flop8/_0_ ;
 wire \proj_14.flop8/_1_ ;
 wire net215;
 wire net216;
 wire \proj_14.flop9/_0_ ;
 wire \proj_14.flop9/_1_ ;
 wire net217;
 wire net218;
 wire \proj__4.flop1/_0_ ;
 wire \proj__4.flop1/_1_ ;
 wire net219;
 wire net220;
 wire \proj__4.flop1/q ;
 wire \proj__4.flop1/s ;
 wire \proj__4.flop2/_0_ ;
 wire \proj__4.flop2/_1_ ;
 wire net221;
 wire net222;
 wire \proj__4.flop2/q ;
 wire \proj__4.flop2/s ;
 wire \proj__4.flop3/_0_ ;
 wire \proj__4.flop3/_1_ ;
 wire net223;
 wire net224;
 wire \proj__4.flop3/q ;
 wire \proj__4.flop3/s ;
 wire \proj__4.flop4/_0_ ;
 wire \proj__4.flop4/_1_ ;
 wire net225;
 wire net226;
 wire \proj__4.flop4/q ;
 wire \proj__4.flop4/s ;
 wire \proj__4.flop5/_0_ ;
 wire \proj__4.flop5/_1_ ;
 wire net227;
 wire net228;
 wire \proj__4.flop5/notq ;
 wire \proj__4.flop5/s ;
 wire \proj__4.flop6/_0_ ;
 wire \proj__4.flop6/_1_ ;
 wire net229;
 wire net230;
 wire \proj__4.flop6/notq ;
 wire \proj__4.flop6/s ;
 wire \proj__4.flop8/_0_ ;
 wire \proj__4.flop8/_1_ ;
 wire net231;
 wire net232;
 wire \proj__4.flop8/notq ;
 wire \proj__4.flop8/s ;
 wire \proj__4.flop9/_0_ ;
 wire \proj__4.flop9/_1_ ;
 wire net233;
 wire net234;
 wire \proj__4.flop9/notq ;
 wire \proj__4.flop9/s ;
 wire net253;
 wire net254;
 wire \proj__9.flop1/_0_ ;
 wire \proj__9.flop1/_1_ ;
 wire net235;
 wire net236;
 wire \proj__9.flop1/notq ;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;

 sg13g2_inv_1 _181_ (.Y(_041_),
    .A(net11));
 sg13g2_nor2_2 _182_ (.A(net8),
    .B(net9),
    .Y(_042_));
 sg13g2_nor3_1 _183_ (.A(net8),
    .B(net9),
    .C(net10),
    .Y(_043_));
 sg13g2_nor2_2 _184_ (.A(net11),
    .B(net10),
    .Y(_044_));
 sg13g2_nand2_1 _185_ (.Y(_045_),
    .A(_042_),
    .B(_044_));
 sg13g2_nor2_1 _186_ (.A(\proj__0.net9 ),
    .B(_045_),
    .Y(_046_));
 sg13g2_nand2_1 _187_ (.Y(_047_),
    .A(net8),
    .B(net9));
 sg13g2_nor3_2 _188_ (.A(net11),
    .B(net10),
    .C(_047_),
    .Y(_048_));
 sg13g2_nor2b_2 _189_ (.A(net8),
    .B_N(net9),
    .Y(_049_));
 sg13g2_nand2b_2 _190_ (.Y(_050_),
    .B(net10),
    .A_N(net11));
 sg13g2_and3_1 _191_ (.X(_051_),
    .A(_041_),
    .B(net10),
    .C(_049_));
 sg13g2_o21ai_1 _192_ (.B1(net40),
    .Y(_052_),
    .A1(_048_),
    .A2(_051_));
 sg13g2_nor2b_2 _193_ (.A(net9),
    .B_N(net8),
    .Y(_053_));
 sg13g2_nor2b_1 _194_ (.A(net10),
    .B_N(net11),
    .Y(_054_));
 sg13g2_and2_1 _195_ (.A(\proj__9.net5 ),
    .B(_054_),
    .X(_055_));
 sg13g2_nor2b_2 _196_ (.A(_050_),
    .B_N(_053_),
    .Y(_056_));
 sg13g2_a22oi_1 _197_ (.Y(_057_),
    .B1(_056_),
    .B2(\proj__5.net9 ),
    .A2(_055_),
    .A1(_053_));
 sg13g2_and2_1 _198_ (.A(_044_),
    .B(_049_),
    .X(_058_));
 sg13g2_nor3_2 _199_ (.A(net8),
    .B(net9),
    .C(_050_),
    .Y(_059_));
 sg13g2_and2_1 _200_ (.A(net11),
    .B(net10),
    .X(_060_));
 sg13g2_and2_1 _201_ (.A(_053_),
    .B(_060_),
    .X(_061_));
 sg13g2_and3_1 _202_ (.X(_062_),
    .A(\proj__8.net7 ),
    .B(_042_),
    .C(_054_));
 sg13g2_and2_2 _203_ (.A(_049_),
    .B(_060_),
    .X(_063_));
 sg13g2_and2_2 _204_ (.A(_042_),
    .B(_060_),
    .X(_064_));
 sg13g2_nand2_1 _205_ (.Y(_065_),
    .A(\proj_12.net9 ),
    .B(_064_));
 sg13g2_nor2_2 _206_ (.A(_047_),
    .B(_050_),
    .Y(_066_));
 sg13g2_nand3_1 _207_ (.B(_044_),
    .C(_053_),
    .A(\proj__1.net9 ),
    .Y(_067_));
 sg13g2_and2_2 _208_ (.A(_049_),
    .B(_054_),
    .X(_068_));
 sg13g2_a22oi_1 _209_ (.Y(_069_),
    .B1(_066_),
    .B2(\proj__7.net5 ),
    .A2(_058_),
    .A1(\proj__2.net9 ));
 sg13g2_a21oi_1 _210_ (.A1(_042_),
    .A2(_044_),
    .Y(_070_),
    .B1(_062_));
 sg13g2_and4_1 _211_ (.A(_052_),
    .B(_065_),
    .C(_067_),
    .D(_070_),
    .X(_000_));
 sg13g2_a22oi_1 _212_ (.Y(_001_),
    .B1(_063_),
    .B2(\proj_14.net11 ),
    .A2(_059_),
    .A1(\proj__4.net11 ));
 sg13g2_a22oi_1 _213_ (.Y(_002_),
    .B1(_068_),
    .B2(\proj_10.net9 ),
    .A2(_061_),
    .A1(\proj_13.net7 ));
 sg13g2_and4_1 _214_ (.A(_057_),
    .B(_069_),
    .C(_001_),
    .D(_002_),
    .X(_003_));
 sg13g2_a21oi_2 _215_ (.B1(_046_),
    .Y(uo_out[0]),
    .A2(_003_),
    .A1(_000_));
 sg13g2_o21ai_1 _216_ (.B1(net38),
    .Y(_004_),
    .A1(_048_),
    .A2(_051_));
 sg13g2_a21oi_1 _217_ (.A1(\proj_13.net8 ),
    .A2(_061_),
    .Y(_005_),
    .B1(_062_));
 sg13g2_a22oi_1 _218_ (.Y(_006_),
    .B1(_064_),
    .B2(\proj_12.net10 ),
    .A2(_063_),
    .A1(\proj_14.net12 ));
 sg13g2_a22oi_1 _219_ (.Y(_007_),
    .B1(_066_),
    .B2(\proj__7.net6 ),
    .A2(_059_),
    .A1(\proj__4.net12 ));
 sg13g2_a22oi_1 _220_ (.Y(_008_),
    .B1(_068_),
    .B2(net37),
    .A2(_058_),
    .A1(\proj__2.net10 ));
 sg13g2_and3_1 _221_ (.X(_009_),
    .A(_004_),
    .B(_007_),
    .C(_008_));
 sg13g2_nand3_1 _222_ (.B(_006_),
    .C(_009_),
    .A(_005_),
    .Y(uo_out[1]));
 sg13g2_nor2_1 _223_ (.A(\proj__0.net10 ),
    .B(_045_),
    .Y(_010_));
 sg13g2_a22oi_1 _224_ (.Y(_011_),
    .B1(_063_),
    .B2(\proj_14.net13 ),
    .A2(_051_),
    .A1(\proj__6.net9 ));
 sg13g2_a22oi_1 _225_ (.Y(_012_),
    .B1(_064_),
    .B2(\proj_12.net11 ),
    .A2(_058_),
    .A1(\proj__2.net11 ));
 sg13g2_a21oi_1 _226_ (.A1(net35),
    .A2(_068_),
    .Y(_013_),
    .B1(_062_));
 sg13g2_a22oi_1 _227_ (.Y(_014_),
    .B1(_059_),
    .B2(\proj__4.net13 ),
    .A2(_044_),
    .A1(_042_));
 sg13g2_nand4_1 _228_ (.B(_012_),
    .C(_013_),
    .A(_011_),
    .Y(_015_),
    .D(_014_));
 sg13g2_nor2b_2 _229_ (.A(_010_),
    .B_N(_015_),
    .Y(uo_out[2]));
 sg13g2_nor2_1 _230_ (.A(\proj__0.net11 ),
    .B(_045_),
    .Y(_016_));
 sg13g2_a22oi_1 _231_ (.Y(_017_),
    .B1(_064_),
    .B2(\proj_12.net12 ),
    .A2(_051_),
    .A1(\proj__6.net10 ));
 sg13g2_a22oi_1 _232_ (.Y(_018_),
    .B1(_063_),
    .B2(\proj_14.net14 ),
    .A2(_059_),
    .A1(\proj__4.net14 ));
 sg13g2_a22oi_1 _233_ (.Y(_019_),
    .B1(_058_),
    .B2(\proj__2.net12 ),
    .A2(_044_),
    .A1(_042_));
 sg13g2_nand4_1 _234_ (.B(_017_),
    .C(_018_),
    .A(_013_),
    .Y(_020_),
    .D(_019_));
 sg13g2_nor2b_2 _235_ (.A(_016_),
    .B_N(_020_),
    .Y(uo_out[3]));
 sg13g2_a221oi_1 _236_ (.B2(_060_),
    .C1(_043_),
    .B1(_053_),
    .A1(_041_),
    .Y(_021_),
    .A2(_049_));
 sg13g2_inv_1 _237_ (.Y(_022_),
    .A(_021_));
 sg13g2_nand2b_1 _238_ (.Y(_023_),
    .B(_021_),
    .A_N(_066_));
 sg13g2_nand2_1 _239_ (.Y(_024_),
    .A(net4),
    .B(_023_));
 sg13g2_nand2_1 _240_ (.Y(_025_),
    .A(\proj_12.net13 ),
    .B(_064_));
 sg13g2_nand2_1 _241_ (.Y(_026_),
    .A(\proj_10.net10 ),
    .B(_068_));
 sg13g2_a22oi_1 _242_ (.Y(_027_),
    .B1(_063_),
    .B2(\proj_14.net15 ),
    .A2(_056_),
    .A1(\proj__5.net10 ));
 sg13g2_a22oi_1 _243_ (.Y(_028_),
    .B1(_059_),
    .B2(\proj__4.net15 ),
    .A2(_048_),
    .A1(\proj__3.net3 ));
 sg13g2_and4_1 _244_ (.A(_067_),
    .B(_025_),
    .C(_026_),
    .D(_028_),
    .X(_029_));
 sg13g2_nand3_1 _245_ (.B(_027_),
    .C(_029_),
    .A(_024_),
    .Y(uo_out[4]));
 sg13g2_nand2_1 _246_ (.Y(_030_),
    .A(\proj__5.net11 ),
    .B(_056_));
 sg13g2_a22oi_1 _247_ (.Y(_031_),
    .B1(_063_),
    .B2(\proj_14.net16 ),
    .A2(_059_),
    .A1(\proj__4.net16 ));
 sg13g2_a22oi_1 _248_ (.Y(_032_),
    .B1(_068_),
    .B2(\proj_10.net11 ),
    .A2(_048_),
    .A1(\proj__3.net4 ));
 sg13g2_nand4_1 _249_ (.B(_030_),
    .C(_031_),
    .A(_067_),
    .Y(_033_),
    .D(_032_));
 sg13g2_a21o_1 _250_ (.A2(_023_),
    .A1(net35),
    .B1(_033_),
    .X(uo_out[5]));
 sg13g2_nand2_1 _251_ (.Y(_034_),
    .A(net6),
    .B(_022_));
 sg13g2_a22oi_1 _252_ (.Y(_035_),
    .B1(_066_),
    .B2(\proj__7.net7 ),
    .A2(_056_),
    .A1(\proj__5.net12 ));
 sg13g2_a22oi_1 _253_ (.Y(_036_),
    .B1(_063_),
    .B2(\proj_14.net17 ),
    .A2(_059_),
    .A1(\proj__4.net17 ));
 sg13g2_a22oi_1 _254_ (.Y(_037_),
    .B1(_068_),
    .B2(\proj_10.net12 ),
    .A2(_048_),
    .A1(\proj__3.net5 ));
 sg13g2_nand4_1 _255_ (.B(_035_),
    .C(_036_),
    .A(_034_),
    .Y(uo_out[6]),
    .D(_037_));
 sg13g2_o21ai_1 _256_ (.B1(net7),
    .Y(_038_),
    .A1(_056_),
    .A2(_022_));
 sg13g2_nand2_1 _257_ (.Y(_039_),
    .A(\proj__4.net18 ),
    .B(_059_));
 sg13g2_a22oi_1 _258_ (.Y(_040_),
    .B1(_068_),
    .B2(\proj_10.net13 ),
    .A2(_066_),
    .A1(\proj__7.net8 ));
 sg13g2_nand3_1 _259_ (.B(_039_),
    .C(_040_),
    .A(_038_),
    .Y(uo_out[7]));
 sg13g2_tiehi \proj_13.flop1/_1__228  (.L_HI(net237));
 sg13g2_tielo \proj_13.flop2/_1__13  (.L_LO(net13));
 sg13g2_tielo \proj_13.flop3/_1__14  (.L_LO(net14));
 sg13g2_tielo \proj_14.flop1/dffsr_15  (.L_LO(net15));
 sg13g2_tielo \proj_14.flop1/_4__16  (.L_LO(net16));
 sg13g2_tielo \proj_14.flop10/dffsr_17  (.L_LO(net17));
 sg13g2_tielo \proj_14.flop10/_4__18  (.L_LO(net18));
 sg13g2_tielo \proj_14.flop11/dffsr_19  (.L_LO(net19));
 sg13g2_tielo \proj_14.flop11/_4__20  (.L_LO(net20));
 sg13g2_tielo \proj_14.flop12/dffsr_21  (.L_LO(net21));
 sg13g2_tielo \proj_14.flop12/_4__22  (.L_LO(net22));
 sg13g2_tielo \proj_14.flop13/dffsr_23  (.L_LO(net23));
 sg13g2_tielo \proj_14.flop13/_4__24  (.L_LO(net24));
 sg13g2_tielo \proj_14.flop14/dffsr_25  (.L_LO(net25));
 sg13g2_tielo \proj_14.flop14/_4__26  (.L_LO(net26));
 sg13g2_tielo \proj_14.flop15/dffsr_27  (.L_LO(net27));
 sg13g2_tielo \proj_14.flop15/_4__28  (.L_LO(net28));
 sg13g2_tielo \proj_14.flop16/dffsr_29  (.L_LO(net29));
 sg13g2_tielo \proj_14.flop16/_4__30  (.L_LO(net30));
 sg13g2_tielo \proj_14.flop17/dffsr_31  (.L_LO(net31));
 sg13g2_tielo \proj_14.flop17/_4__32  (.L_LO(net32));
 sg13g2_tielo \proj_14.flop18/dffsr_33  (.L_LO(net33));
 sg13g2_tielo \proj_14.flop18/_4__34  (.L_LO(net34));
 sg13g2_tielo \proj_14.flop19/dffsr_35  (.L_LO(net44));
 sg13g2_tielo \proj_14.flop19/_4__36  (.L_LO(net45));
 sg13g2_tielo \proj_14.flop2/dffsr_37  (.L_LO(net46));
 sg13g2_tielo \proj_14.flop2/_4__38  (.L_LO(net47));
 sg13g2_tielo \proj_14.flop20/dffsr_39  (.L_LO(net48));
 sg13g2_tielo \proj_14.flop20/_4__40  (.L_LO(net49));
 sg13g2_tielo \proj_14.flop21/dffsr_41  (.L_LO(net50));
 sg13g2_tielo \proj_14.flop21/_4__42  (.L_LO(net51));
 sg13g2_tielo \proj_14.flop22/dffsr_43  (.L_LO(net52));
 sg13g2_tielo \proj_14.flop22/_4__44  (.L_LO(net53));
 sg13g2_tielo \proj_14.flop23/dffsr_45  (.L_LO(net54));
 sg13g2_tielo \proj_14.flop23/_4__46  (.L_LO(net55));
 sg13g2_tielo \proj_14.flop24/dffsr_47  (.L_LO(net56));
 sg13g2_tielo \proj_14.flop24/_4__48  (.L_LO(net57));
 sg13g2_tielo \proj_14.flop25/dffsr_49  (.L_LO(net58));
 sg13g2_tielo \proj_14.flop25/_4__50  (.L_LO(net59));
 sg13g2_tielo \proj_14.flop26/dffsr_51  (.L_LO(net60));
 sg13g2_tielo \proj_14.flop26/_4__52  (.L_LO(net61));
 sg13g2_tielo \proj_14.flop27/dffsr_53  (.L_LO(net62));
 sg13g2_tielo \proj_14.flop27/_4__54  (.L_LO(net63));
 sg13g2_tielo \proj_14.flop28/_1__55  (.L_LO(net64));
 sg13g2_tielo \proj_14.flop29/dffsr_56  (.L_LO(net65));
 sg13g2_tielo \proj_14.flop29/_4__57  (.L_LO(net66));
 sg13g2_tielo \proj_14.flop3/dffsr_58  (.L_LO(net67));
 sg13g2_tielo \proj_14.flop3/_4__59  (.L_LO(net68));
 sg13g2_tielo \proj_14.flop30/dffsr_60  (.L_LO(net69));
 sg13g2_tielo \proj_14.flop30/_4__61  (.L_LO(net70));
 sg13g2_tielo \proj_14.flop31/dffsr_62  (.L_LO(net71));
 sg13g2_tielo \proj_14.flop32/dffsr_63  (.L_LO(net72));
 sg13g2_tielo \proj_14.flop32/_4__64  (.L_LO(net73));
 sg13g2_tielo \proj_14.flop33/dffsr_65  (.L_LO(net74));
 sg13g2_tielo \proj_14.flop33/_4__66  (.L_LO(net75));
 sg13g2_tielo \proj_14.flop34/dffsr_67  (.L_LO(net76));
 sg13g2_tielo \proj_14.flop34/_4__68  (.L_LO(net77));
 sg13g2_tielo \proj_14.flop35/dffsr_69  (.L_LO(net78));
 sg13g2_tielo \proj_14.flop35/_5__70  (.L_LO(net79));
 sg13g2_tielo \proj_14.flop36/dffsr_71  (.L_LO(net80));
 sg13g2_tielo \proj_14.flop36/_4__72  (.L_LO(net81));
 sg13g2_tielo \proj_14.flop37/dffsr_73  (.L_LO(net82));
 sg13g2_tielo \proj_14.flop37/_5__74  (.L_LO(net83));
 sg13g2_tielo \proj_14.flop4/dffsr_75  (.L_LO(net84));
 sg13g2_tielo \proj_14.flop4/_5__76  (.L_LO(net85));
 sg13g2_tielo \proj_14.flop46/_1__77  (.L_LO(net86));
 sg13g2_tielo \proj_14.flop47/_1__78  (.L_LO(net87));
 sg13g2_tielo \proj_14.flop48/_1__79  (.L_LO(net88));
 sg13g2_tielo \proj_14.flop49/_1__80  (.L_LO(net89));
 sg13g2_tielo \proj_14.flop5/dffsr_81  (.L_LO(net90));
 sg13g2_tielo \proj_14.flop5/_4__82  (.L_LO(net91));
 sg13g2_tielo \proj_14.flop50/_1__83  (.L_LO(net92));
 sg13g2_tielo \proj_14.flop51/_1__84  (.L_LO(net93));
 sg13g2_tielo \proj_14.flop52/_1__85  (.L_LO(net94));
 sg13g2_tielo \proj_14.flop53/_1__86  (.L_LO(net95));
 sg13g2_tielo \proj_14.flop54/_1__87  (.L_LO(net96));
 sg13g2_tielo \proj_14.flop55/_1__88  (.L_LO(net97));
 sg13g2_tielo \proj_14.flop56/_1__89  (.L_LO(net98));
 sg13g2_tielo \proj_14.flop6/dffsr_90  (.L_LO(net99));
 sg13g2_tielo \proj_14.flop6/_5__91  (.L_LO(net100));
 sg13g2_tielo \proj_14.flop7/dffsr_92  (.L_LO(net101));
 sg13g2_tielo \proj_14.flop7/_4__93  (.L_LO(net102));
 sg13g2_tielo \proj_14.flop8/dffsr_94  (.L_LO(net103));
 sg13g2_tielo \proj_14.flop8/_4__95  (.L_LO(net104));
 sg13g2_tielo \proj_14.flop9/dffsr_96  (.L_LO(net105));
 sg13g2_tielo \proj_14.flop9/_5__97  (.L_LO(net106));
 sg13g2_tielo \proj_14.not1/_0__98  (.L_LO(net107));
 sg13g2_tielo \proj_14.not5/_0__99  (.L_LO(net108));
 sg13g2_tielo \proj__4.flop1/dffsr_100  (.L_LO(net109));
 sg13g2_tielo \proj__4.flop1/_5__101  (.L_LO(net110));
 sg13g2_tielo \proj__4.flop2/dffsr_102  (.L_LO(net111));
 sg13g2_tielo \proj__4.flop2/_5__103  (.L_LO(net112));
 sg13g2_tielo \proj__4.flop3/dffsr_104  (.L_LO(net113));
 sg13g2_tielo \proj__4.flop3/_5__105  (.L_LO(net114));
 sg13g2_tielo \proj__4.flop4/dffsr_106  (.L_LO(net115));
 sg13g2_tielo \proj__4.flop4/_5__107  (.L_LO(net116));
 sg13g2_tielo \proj__4.flop5/dffsr_108  (.L_LO(net117));
 sg13g2_tielo \proj__4.flop5/_5__109  (.L_LO(net118));
 sg13g2_tielo \proj__4.flop6/dffsr_110  (.L_LO(net119));
 sg13g2_tielo \proj__4.flop6/_5__111  (.L_LO(net120));
 sg13g2_tielo \proj__4.flop8/dffsr_112  (.L_LO(net121));
 sg13g2_tielo \proj__4.flop8/_5__113  (.L_LO(net122));
 sg13g2_tielo \proj__4.flop9/dffsr_114  (.L_LO(net123));
 sg13g2_tielo \proj__4.flop9/_5__115  (.L_LO(net124));
 sg13g2_tielo \proj__7.flop1/_1__116  (.L_LO(net125));
 sg13g2_tielo \proj__7.flop2/_1__117  (.L_LO(net126));
 sg13g2_tielo \proj__9.flop1/dffsr_118  (.L_LO(net127));
 sg13g2_tielo \proj__9.flop1/_4__119  (.L_LO(net128));
 sg13g2_tielo \proj__9.not3/_0__120  (.L_LO(net129));
 sg13g2_tielo tt_um_wokwi_group_3_121 (.L_LO(net130));
 sg13g2_tielo tt_um_wokwi_group_3_122 (.L_LO(net131));
 sg13g2_tielo tt_um_wokwi_group_3_123 (.L_LO(net132));
 sg13g2_tielo tt_um_wokwi_group_3_124 (.L_LO(net133));
 sg13g2_tielo tt_um_wokwi_group_3_125 (.L_LO(net134));
 sg13g2_tielo tt_um_wokwi_group_3_126 (.L_LO(net135));
 sg13g2_tielo tt_um_wokwi_group_3_127 (.L_LO(net136));
 sg13g2_tielo tt_um_wokwi_group_3_128 (.L_LO(net137));
 sg13g2_tielo tt_um_wokwi_group_3_129 (.L_LO(net138));
 sg13g2_tielo tt_um_wokwi_group_3_130 (.L_LO(net139));
 sg13g2_tielo tt_um_wokwi_group_3_131 (.L_LO(net140));
 sg13g2_tielo tt_um_wokwi_group_3_132 (.L_LO(net141));
 sg13g2_tielo tt_um_wokwi_group_3_133 (.L_LO(net142));
 sg13g2_tielo tt_um_wokwi_group_3_134 (.L_LO(net143));
 sg13g2_tielo tt_um_wokwi_group_3_135 (.L_LO(net144));
 sg13g2_tielo tt_um_wokwi_group_3_136 (.L_LO(net145));
 sg13g2_tielo \proj_14.flop1/dffsr_137  (.L_LO(net146));
 sg13g2_mux2_1 \proj_10.mux2/_0_  (.A0(net41),
    .A1(net39),
    .S(net37),
    .X(\proj_10.net9 ));
 sg13g2_nand2_1 \proj_10.nand1/_0_  (.Y(\proj_10.net10 ),
    .A(\proj_10.nand1/b ),
    .B(net36));
 sg13g2_inv_1 \proj_10.not1/_0_  (.Y(\proj_10.net12 ),
    .A(net6));
 sg13g2_inv_1 \proj_10.not2/_0_  (.Y(\proj_10.net13 ),
    .A(net7));
 sg13g2_xor2_1 \proj_10.xor1/_0_  (.B(net4),
    .A(net35),
    .X(\proj_10.net11 ));
 sg13g2_and2_1 \proj_12.and1/_0_  (.A(net38),
    .B(net40),
    .X(\proj_12.net18 ));
 sg13g2_and2_1 \proj_12.and2/_0_  (.A(net36),
    .B(net37),
    .X(\proj_12.net20 ));
 sg13g2_and2_1 \proj_12.and4/_0_  (.A(\proj_12.net19 ),
    .B(\proj_12.net18 ),
    .X(\proj_12.net21 ));
 sg13g2_and2_1 \proj_12.and5/_0_  (.A(net35),
    .B(net4),
    .X(\proj_12.net24 ));
 sg13g2_and2_1 \proj_12.and6/_0_  (.A(\proj_12.net23 ),
    .B(\proj_12.net22 ),
    .X(\proj_12.net25 ));
 sg13g2_and2_1 \proj_12.and7/_0_  (.A(net7),
    .B(net6),
    .X(\proj_12.net28 ));
 sg13g2_and2_1 \proj_12.and8/_0_  (.A(\proj_12.net27 ),
    .B(\proj_12.net26 ),
    .X(\proj_12.net29 ));
 sg13g2_or2_1 \proj_12.or1/_0_  (.X(\proj_12.net22 ),
    .B(\proj_12.net21 ),
    .A(\proj_12.net20 ));
 sg13g2_or2_1 \proj_12.or2/_0_  (.X(\proj_12.net26 ),
    .B(\proj_12.net25 ),
    .A(\proj_12.net24 ));
 sg13g2_or2_1 \proj_12.or3/_0_  (.X(\proj_12.net13 ),
    .B(\proj_12.net29 ),
    .A(\proj_12.net28 ));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(net40),
    .A(net38),
    .X(\proj_12.net9 ));
 sg13g2_xor2_1 \proj_12.xor2/_0_  (.B(net37),
    .A(net36),
    .X(\proj_12.net19 ));
 sg13g2_xor2_1 \proj_12.xor3/_0_  (.B(\proj_12.net19 ),
    .A(\proj_12.net18 ),
    .X(\proj_12.net10 ));
 sg13g2_xor2_1 \proj_12.xor4/_0_  (.B(net4),
    .A(net35),
    .X(\proj_12.net23 ));
 sg13g2_xor2_1 \proj_12.xor5/_0_  (.B(\proj_12.net23 ),
    .A(\proj_12.net22 ),
    .X(\proj_12.net11 ));
 sg13g2_xor2_1 \proj_12.xor6/_0_  (.B(net6),
    .A(net7),
    .X(\proj_12.net27 ));
 sg13g2_xor2_1 \proj_12.xor7/_0_  (.B(\proj_12.net27 ),
    .A(\proj_12.net26 ),
    .X(\proj_12.net12 ));
 sg13g2_dfrbp_1 \proj_13.flop1/_1_  (.CLK(net12),
    .RESET_B(net237),
    .D(net41),
    .Q_N(\proj_13.flop1/notq ),
    .Q(\proj_13.net12 ));
 sg13g2_tiehi \proj_13.flop2/_1__229  (.L_HI(net238));
 sg13g2_dfrbp_1 \proj_13.flop2/_1_  (.CLK(net13),
    .RESET_B(net238),
    .D(\proj_13.net12 ),
    .Q_N(\proj_13.flop2/notq ),
    .Q(\proj_13.net13 ));
 sg13g2_tiehi \proj_13.flop3/_1__230  (.L_HI(net239));
 sg13g2_dfrbp_1 \proj_13.flop3/_1_  (.CLK(net14),
    .RESET_B(net239),
    .D(\proj_13.net13 ),
    .Q_N(\proj_13.flop3/notq ),
    .Q(\proj_13.net8 ));
 sg13g2_tiehi \proj_14.flop28/_1__231  (.L_HI(net240));
 sg13g2_inv_1 \proj_13.not5/_0_  (.Y(\proj_13.net7 ),
    .A(\proj_13.net13 ));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(\proj_14.net30 ),
    .B(\proj_14.net33 ),
    .X(\proj_14.net58 ));
 sg13g2_and2_1 \proj_14.and10/_0_  (.A(\proj_14.net32 ),
    .B(\proj_14.net30 ),
    .X(\proj_14.net64 ));
 sg13g2_and2_1 \proj_14.and11/_0_  (.A(\proj_14.net40 ),
    .B(\proj_14.net43 ),
    .X(\proj_14.net68 ));
 sg13g2_and2_1 \proj_14.and12/_0_  (.A(\proj_14.net68 ),
    .B(\proj_14.net37 ),
    .X(\proj_14.net69 ));
 sg13g2_and2_1 \proj_14.and13/_0_  (.A(\proj_14.net68 ),
    .B(\proj_14.net36 ),
    .X(\proj_14.net70 ));
 sg13g2_and2_1 \proj_14.and14/_0_  (.A(\proj_14.net39 ),
    .B(\proj_14.net43 ),
    .X(\proj_14.net71 ));
 sg13g2_and2_1 \proj_14.and15/_0_  (.A(\proj_14.net71 ),
    .B(\proj_14.net37 ),
    .X(\proj_14.net72 ));
 sg13g2_and2_1 \proj_14.and16/_0_  (.A(\proj_14.net71 ),
    .B(\proj_14.net36 ),
    .X(\proj_14.net73 ));
 sg13g2_and2_1 \proj_14.and17/_0_  (.A(\proj_14.net74 ),
    .B(\proj_14.net37 ),
    .X(\proj_14.net75 ));
 sg13g2_and2_1 \proj_14.and18/_0_  (.A(\proj_14.net74 ),
    .B(\proj_14.net36 ),
    .X(\proj_14.net76 ));
 sg13g2_and2_1 \proj_14.and19/_0_  (.A(\proj_14.net42 ),
    .B(\proj_14.net39 ),
    .X(\proj_14.net77 ));
 sg13g2_and2_1 \proj_14.and2/_0_  (.A(\proj_14.net58 ),
    .B(\proj_14.net27 ),
    .X(\proj_14.net59 ));
 sg13g2_and2_1 \proj_14.and20/_0_  (.A(\proj_14.net42 ),
    .B(\proj_14.net40 ),
    .X(\proj_14.net74 ));
 sg13g2_and2_1 \proj_14.and21/_0_  (.A(\proj_14.net54 ),
    .B(\proj_14.net57 ),
    .X(\proj_14.net78 ));
 sg13g2_and2_1 \proj_14.and22/_0_  (.A(\proj_14.net78 ),
    .B(\proj_14.net51 ),
    .X(\proj_14.net79 ));
 sg13g2_and2_1 \proj_14.and23/_0_  (.A(\proj_14.net78 ),
    .B(\proj_14.net50 ),
    .X(\proj_14.net80 ));
 sg13g2_and2_1 \proj_14.and24/_0_  (.A(\proj_14.net53 ),
    .B(\proj_14.net57 ),
    .X(\proj_14.net81 ));
 sg13g2_and2_1 \proj_14.and25/_0_  (.A(\proj_14.net81 ),
    .B(\proj_14.net51 ),
    .X(\proj_14.net82 ));
 sg13g2_and2_1 \proj_14.and26/_0_  (.A(\proj_14.net81 ),
    .B(\proj_14.net50 ),
    .X(\proj_14.net83 ));
 sg13g2_and2_1 \proj_14.and27/_0_  (.A(\proj_14.net84 ),
    .B(\proj_14.net51 ),
    .X(\proj_14.net85 ));
 sg13g2_and2_1 \proj_14.and28/_0_  (.A(\proj_14.net84 ),
    .B(\proj_14.net50 ),
    .X(\proj_14.net86 ));
 sg13g2_and2_1 \proj_14.and29/_0_  (.A(\proj_14.net56 ),
    .B(\proj_14.net53 ),
    .X(\proj_14.net87 ));
 sg13g2_and2_1 \proj_14.and3/_0_  (.A(\proj_14.net58 ),
    .B(\proj_14.net26 ),
    .X(\proj_14.net60 ));
 sg13g2_and2_1 \proj_14.and30/_0_  (.A(\proj_14.net56 ),
    .B(\proj_14.net54 ),
    .X(\proj_14.net84 ));
 sg13g2_and2_1 \proj_14.and31/_0_  (.A(\proj_14.net105 ),
    .B(\proj_14.net110 ),
    .X(\proj_14.net116 ));
 sg13g2_and2_1 \proj_14.and32/_0_  (.A(\proj_14.net116 ),
    .B(\proj_14.net114 ),
    .X(\proj_14.net121 ));
 sg13g2_and2_1 \proj_14.and33/_0_  (.A(\proj_14.net121 ),
    .B(\proj_14.net119 ),
    .X(\proj_14.net126 ));
 sg13g2_and2_1 \proj_14.and34/_0_  (.A(\proj_14.net126 ),
    .B(\proj_14.net124 ),
    .X(\proj_14.net131 ));
 sg13g2_and2_1 \proj_14.and35/_0_  (.A(\proj_14.net137 ),
    .B(\proj_14.net135 ),
    .X(\proj_14.net142 ));
 sg13g2_and2_1 \proj_14.and36/_0_  (.A(\proj_14.net142 ),
    .B(\proj_14.net140 ),
    .X(\proj_14.net147 ));
 sg13g2_and2_1 \proj_14.and37/_0_  (.A(\proj_14.net147 ),
    .B(\proj_14.net145 ),
    .X(\proj_14.net152 ));
 sg13g2_and2_1 \proj_14.and38/_0_  (.A(\proj_14.net152 ),
    .B(\proj_14.net150 ),
    .X(\proj_14.net157 ));
 sg13g2_and2_1 \proj_14.and39/_0_  (.A(\proj_14.net131 ),
    .B(\proj_14.net129 ),
    .X(\proj_14.net137 ));
 sg13g2_and2_1 \proj_14.and4/_0_  (.A(\proj_14.net29 ),
    .B(\proj_14.net33 ),
    .X(\proj_14.net61 ));
 sg13g2_and2_1 \proj_14.and40/_0_  (.A(\proj_14.net157 ),
    .B(\proj_14.net155 ),
    .X(\proj_14.net162 ));
 sg13g2_and2_1 \proj_14.and41/_0_  (.A(\proj_14.net162 ),
    .B(\proj_14.net160 ),
    .X(\proj_14.net167 ));
 sg13g2_and2_1 \proj_14.and42/_0_  (.A(\proj_14.net167 ),
    .B(\proj_14.net165 ),
    .X(\proj_14.net172 ));
 sg13g2_and2_1 \proj_14.and43/_0_  (.A(\proj_14.net172 ),
    .B(\proj_14.net170 ),
    .X(\proj_14.net177 ));
 sg13g2_and2_1 \proj_14.and44/_0_  (.A(\proj_14.net193 ),
    .B(\proj_14.net192 ),
    .X(\proj_14.net194 ));
 sg13g2_and2_1 \proj_14.and45/_0_  (.A(\proj_14.net196 ),
    .B(\proj_14.net195 ),
    .X(\proj_14.net197 ));
 sg13g2_and2_1 \proj_14.and46/_0_  (.A(\proj_14.net199 ),
    .B(\proj_14.net198 ),
    .X(\proj_14.net200 ));
 sg13g2_and2_1 \proj_14.and47/_0_  (.A(\proj_14.net202 ),
    .B(\proj_14.net201 ),
    .X(\proj_14.net203 ));
 sg13g2_and2_1 \proj_14.and48/_0_  (.A(\proj_14.net203 ),
    .B(\proj_14.net200 ),
    .X(\proj_14.net204 ));
 sg13g2_and2_1 \proj_14.and49/_0_  (.A(\proj_14.net197 ),
    .B(\proj_14.net205 ),
    .X(\proj_14.net206 ));
 sg13g2_and2_1 \proj_14.and5/_0_  (.A(\proj_14.net61 ),
    .B(\proj_14.net27 ),
    .X(\proj_14.net62 ));
 sg13g2_and2_1 \proj_14.and50/_0_  (.A(\proj_14.net204 ),
    .B(\proj_14.net206 ),
    .X(\proj_14.net178 ));
 sg13g2_and2_1 \proj_14.and51/_0_  (.A(\proj_14.net59 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net234 ));
 sg13g2_and2_1 \proj_14.and52/_0_  (.A(\proj_14.net60 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net235 ));
 sg13g2_and2_1 \proj_14.and53/_0_  (.A(\proj_14.net62 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net236 ));
 sg13g2_and2_1 \proj_14.and54/_0_  (.A(\proj_14.net63 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net237 ));
 sg13g2_and2_1 \proj_14.and55/_0_  (.A(\proj_14.net65 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net238 ));
 sg13g2_and2_1 \proj_14.and57/_0_  (.A(\proj_14.net67 ),
    .B(\proj_14.net210 ),
    .X(\proj_14.net239 ));
 sg13g2_and2_1 \proj_14.and58/_0_  (.A(\proj_14.net59 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net240 ));
 sg13g2_and2_1 \proj_14.and59/_0_  (.A(\proj_14.net60 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net241 ));
 sg13g2_and2_1 \proj_14.and6/_0_  (.A(\proj_14.net61 ),
    .B(\proj_14.net26 ),
    .X(\proj_14.net63 ));
 sg13g2_and2_1 \proj_14.and60/_0_  (.A(\proj_14.net62 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net242 ));
 sg13g2_and2_1 \proj_14.and61/_0_  (.A(\proj_14.net63 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net243 ));
 sg13g2_and2_1 \proj_14.and62/_0_  (.A(\proj_14.net65 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net244 ));
 sg13g2_and2_1 \proj_14.and63/_0_  (.A(\proj_14.net66 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net245 ));
 sg13g2_and2_1 \proj_14.and64/_0_  (.A(\proj_14.net182 ),
    .B(\proj_14.net181 ),
    .X(\proj_14.net183 ));
 sg13g2_and2_1 \proj_14.and65/_0_  (.A(\proj_14.net67 ),
    .B(\proj_14.net209 ),
    .X(\proj_14.net246 ));
 sg13g2_and2_1 \proj_14.and66/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net235 ),
    .X(\proj_14.net249 ));
 sg13g2_and2_1 \proj_14.and67/_0_  (.A(\proj_14.net235 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net248 ));
 sg13g2_and2_1 \proj_14.and68/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net238 ),
    .X(\proj_14.net252 ));
 sg13g2_and2_1 \proj_14.and69/_0_  (.A(\proj_14.net238 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net254 ));
 sg13g2_and2_1 \proj_14.and7/_0_  (.A(\proj_14.net64 ),
    .B(\proj_14.net27 ),
    .X(\proj_14.net65 ));
 sg13g2_and2_1 \proj_14.and70/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net239 ),
    .X(\proj_14.net258 ));
 sg13g2_and2_1 \proj_14.and71/_0_  (.A(\proj_14.net239 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net256 ));
 sg13g2_and2_1 \proj_14.and72/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net242 ),
    .X(\proj_14.net265 ));
 sg13g2_and2_1 \proj_14.and73/_0_  (.A(\proj_14.net242 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net261 ));
 sg13g2_and2_1 \proj_14.and74/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net245 ),
    .X(\proj_14.net267 ));
 sg13g2_and2_1 \proj_14.and75/_0_  (.A(\proj_14.net214 ),
    .B(\proj_14.net246 ),
    .X(\proj_14.net259 ));
 sg13g2_and2_1 \proj_14.and76/_0_  (.A(\proj_14.net246 ),
    .B(\proj_14.net215 ),
    .X(\proj_14.net269 ));
 sg13g2_and2_1 \proj_14.and77/_0_  (.A(\proj_14.net194 ),
    .B(\proj_14.net135 ),
    .X(\proj_14.net205 ));
 sg13g2_and2_1 \proj_14.and8/_0_  (.A(\proj_14.net64 ),
    .B(\proj_14.net26 ),
    .X(\proj_14.net66 ));
 sg13g2_and2_1 \proj_14.and9/_0_  (.A(\proj_14.net32 ),
    .B(\proj_14.net29 ),
    .X(\proj_14.net67 ));
 sg13g2_inv_1 \proj_14.flop1/_4_  (.Y(\proj_14.flop1/_1_ ),
    .A(net16));
 sg13g2_inv_1 \proj_14.flop1/_5_  (.Y(\proj_14.flop1/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop1/dffsr_138  (.L_LO(net147));
 sg13g2_tielo \proj_14.flop10/dffsr_139  (.L_LO(net148));
 sg13g2_sdfbbp_1 \proj_14.flop1/dffsr  (.Q(\proj_14.net26 ),
    .Q_N(\proj_14.net27 ),
    .RESET_B(\proj_14.flop1/_0_ ),
    .SET_B(\proj_14.flop1/_1_ ),
    .D(\proj_14.net23 ),
    .SCE(net147),
    .SCD(net146),
    .CLK(net15));
 sg13g2_inv_1 \proj_14.flop10/_4_  (.Y(\proj_14.flop10/_1_ ),
    .A(net18));
 sg13g2_inv_1 \proj_14.flop10/_5_  (.Y(\proj_14.flop10/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop10/dffsr_140  (.L_LO(net149));
 sg13g2_tielo \proj_14.flop11/dffsr_141  (.L_LO(net150));
 sg13g2_sdfbbp_1 \proj_14.flop10/dffsr  (.Q(\proj_14.net105 ),
    .Q_N(\proj_14.net106 ),
    .RESET_B(\proj_14.flop10/_0_ ),
    .SET_B(\proj_14.flop10/_1_ ),
    .D(\proj_14.net102 ),
    .SCE(net149),
    .SCD(net148),
    .CLK(net17));
 sg13g2_inv_1 \proj_14.flop11/_4_  (.Y(\proj_14.flop11/_1_ ),
    .A(net20));
 sg13g2_inv_1 \proj_14.flop11/_5_  (.Y(\proj_14.flop11/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop11/dffsr_142  (.L_LO(net151));
 sg13g2_tielo \proj_14.flop12/dffsr_143  (.L_LO(net152));
 sg13g2_sdfbbp_1 \proj_14.flop11/dffsr  (.Q(\proj_14.net110 ),
    .Q_N(\proj_14.net111 ),
    .RESET_B(\proj_14.flop11/_0_ ),
    .SET_B(\proj_14.flop11/_1_ ),
    .D(\proj_14.net108 ),
    .SCE(net151),
    .SCD(net150),
    .CLK(net19));
 sg13g2_inv_1 \proj_14.flop12/_4_  (.Y(\proj_14.flop12/_1_ ),
    .A(net22));
 sg13g2_inv_1 \proj_14.flop12/_5_  (.Y(\proj_14.flop12/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop12/dffsr_144  (.L_LO(net153));
 sg13g2_tielo \proj_14.flop13/dffsr_145  (.L_LO(net154));
 sg13g2_sdfbbp_1 \proj_14.flop12/dffsr  (.Q(\proj_14.net114 ),
    .Q_N(\proj_14.net115 ),
    .RESET_B(\proj_14.flop12/_0_ ),
    .SET_B(\proj_14.flop12/_1_ ),
    .D(\proj_14.net112 ),
    .SCE(net153),
    .SCD(net152),
    .CLK(net21));
 sg13g2_inv_1 \proj_14.flop13/_4_  (.Y(\proj_14.flop13/_1_ ),
    .A(net24));
 sg13g2_inv_1 \proj_14.flop13/_5_  (.Y(\proj_14.flop13/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop13/dffsr_146  (.L_LO(net155));
 sg13g2_tielo \proj_14.flop14/dffsr_147  (.L_LO(net156));
 sg13g2_sdfbbp_1 \proj_14.flop13/dffsr  (.Q(\proj_14.net119 ),
    .Q_N(\proj_14.net120 ),
    .RESET_B(\proj_14.flop13/_0_ ),
    .SET_B(\proj_14.flop13/_1_ ),
    .D(\proj_14.net117 ),
    .SCE(net155),
    .SCD(net154),
    .CLK(net23));
 sg13g2_inv_1 \proj_14.flop14/_4_  (.Y(\proj_14.flop14/_1_ ),
    .A(net26));
 sg13g2_inv_1 \proj_14.flop14/_5_  (.Y(\proj_14.flop14/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop14/dffsr_148  (.L_LO(net157));
 sg13g2_tielo \proj_14.flop15/dffsr_149  (.L_LO(net158));
 sg13g2_sdfbbp_1 \proj_14.flop14/dffsr  (.Q(\proj_14.net124 ),
    .Q_N(\proj_14.net125 ),
    .RESET_B(\proj_14.flop14/_0_ ),
    .SET_B(\proj_14.flop14/_1_ ),
    .D(\proj_14.net122 ),
    .SCE(net157),
    .SCD(net156),
    .CLK(net25));
 sg13g2_inv_1 \proj_14.flop15/_4_  (.Y(\proj_14.flop15/_1_ ),
    .A(net28));
 sg13g2_inv_1 \proj_14.flop15/_5_  (.Y(\proj_14.flop15/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop15/dffsr_150  (.L_LO(net159));
 sg13g2_tielo \proj_14.flop16/dffsr_151  (.L_LO(net160));
 sg13g2_sdfbbp_1 \proj_14.flop15/dffsr  (.Q(\proj_14.net129 ),
    .Q_N(\proj_14.net130 ),
    .RESET_B(\proj_14.flop15/_0_ ),
    .SET_B(\proj_14.flop15/_1_ ),
    .D(\proj_14.net127 ),
    .SCE(net159),
    .SCD(net158),
    .CLK(net27));
 sg13g2_inv_1 \proj_14.flop16/_4_  (.Y(\proj_14.flop16/_1_ ),
    .A(net30));
 sg13g2_inv_1 \proj_14.flop16/_5_  (.Y(\proj_14.flop16/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop16/dffsr_152  (.L_LO(net161));
 sg13g2_tielo \proj_14.flop17/dffsr_153  (.L_LO(net162));
 sg13g2_sdfbbp_1 \proj_14.flop16/dffsr  (.Q(\proj_14.net135 ),
    .Q_N(\proj_14.net136 ),
    .RESET_B(\proj_14.flop16/_0_ ),
    .SET_B(\proj_14.flop16/_1_ ),
    .D(\proj_14.net133 ),
    .SCE(net161),
    .SCD(net160),
    .CLK(net29));
 sg13g2_inv_1 \proj_14.flop17/_4_  (.Y(\proj_14.flop17/_1_ ),
    .A(net32));
 sg13g2_inv_1 \proj_14.flop17/_5_  (.Y(\proj_14.flop17/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop17/dffsr_154  (.L_LO(net163));
 sg13g2_tielo \proj_14.flop18/dffsr_155  (.L_LO(net164));
 sg13g2_sdfbbp_1 \proj_14.flop17/dffsr  (.Q(\proj_14.net140 ),
    .Q_N(\proj_14.net141 ),
    .RESET_B(\proj_14.flop17/_0_ ),
    .SET_B(\proj_14.flop17/_1_ ),
    .D(\proj_14.net138 ),
    .SCE(net163),
    .SCD(net162),
    .CLK(net31));
 sg13g2_inv_1 \proj_14.flop18/_4_  (.Y(\proj_14.flop18/_1_ ),
    .A(net34));
 sg13g2_inv_1 \proj_14.flop18/_5_  (.Y(\proj_14.flop18/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop18/dffsr_156  (.L_LO(net165));
 sg13g2_tielo \proj_14.flop19/dffsr_157  (.L_LO(net166));
 sg13g2_sdfbbp_1 \proj_14.flop18/dffsr  (.Q(\proj_14.net145 ),
    .Q_N(\proj_14.net146 ),
    .RESET_B(\proj_14.flop18/_0_ ),
    .SET_B(\proj_14.flop18/_1_ ),
    .D(\proj_14.net143 ),
    .SCE(net165),
    .SCD(net164),
    .CLK(net33));
 sg13g2_inv_1 \proj_14.flop19/_4_  (.Y(\proj_14.flop19/_1_ ),
    .A(net45));
 sg13g2_inv_1 \proj_14.flop19/_5_  (.Y(\proj_14.flop19/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop19/dffsr_158  (.L_LO(net167));
 sg13g2_tielo \proj_14.flop2/dffsr_159  (.L_LO(net168));
 sg13g2_sdfbbp_1 \proj_14.flop19/dffsr  (.Q(\proj_14.net150 ),
    .Q_N(\proj_14.net151 ),
    .RESET_B(\proj_14.flop19/_0_ ),
    .SET_B(\proj_14.flop19/_1_ ),
    .D(\proj_14.net148 ),
    .SCE(net167),
    .SCD(net166),
    .CLK(net44));
 sg13g2_inv_1 \proj_14.flop2/_4_  (.Y(\proj_14.flop2/_1_ ),
    .A(net47));
 sg13g2_inv_1 \proj_14.flop2/_5_  (.Y(\proj_14.flop2/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop2/dffsr_160  (.L_LO(net169));
 sg13g2_tielo \proj_14.flop20/dffsr_161  (.L_LO(net170));
 sg13g2_sdfbbp_1 \proj_14.flop2/dffsr  (.Q(\proj_14.net29 ),
    .Q_N(\proj_14.net30 ),
    .RESET_B(\proj_14.flop2/_0_ ),
    .SET_B(\proj_14.flop2/_1_ ),
    .D(\proj_14.net28 ),
    .SCE(net169),
    .SCD(net168),
    .CLK(net46));
 sg13g2_inv_1 \proj_14.flop20/_4_  (.Y(\proj_14.flop20/_1_ ),
    .A(net49));
 sg13g2_inv_1 \proj_14.flop20/_5_  (.Y(\proj_14.flop20/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop20/dffsr_162  (.L_LO(net171));
 sg13g2_tielo \proj_14.flop21/dffsr_163  (.L_LO(net172));
 sg13g2_sdfbbp_1 \proj_14.flop20/dffsr  (.Q(\proj_14.net155 ),
    .Q_N(\proj_14.net156 ),
    .RESET_B(\proj_14.flop20/_0_ ),
    .SET_B(\proj_14.flop20/_1_ ),
    .D(\proj_14.net153 ),
    .SCE(net171),
    .SCD(net170),
    .CLK(net48));
 sg13g2_inv_1 \proj_14.flop21/_4_  (.Y(\proj_14.flop21/_1_ ),
    .A(net51));
 sg13g2_inv_1 \proj_14.flop21/_5_  (.Y(\proj_14.flop21/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop21/dffsr_164  (.L_LO(net173));
 sg13g2_tielo \proj_14.flop22/dffsr_165  (.L_LO(net174));
 sg13g2_sdfbbp_1 \proj_14.flop21/dffsr  (.Q(\proj_14.net160 ),
    .Q_N(\proj_14.net161 ),
    .RESET_B(\proj_14.flop21/_0_ ),
    .SET_B(\proj_14.flop21/_1_ ),
    .D(\proj_14.net158 ),
    .SCE(net173),
    .SCD(net172),
    .CLK(net50));
 sg13g2_inv_1 \proj_14.flop22/_4_  (.Y(\proj_14.flop22/_1_ ),
    .A(net53));
 sg13g2_inv_1 \proj_14.flop22/_5_  (.Y(\proj_14.flop22/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop22/dffsr_166  (.L_LO(net175));
 sg13g2_tielo \proj_14.flop23/dffsr_167  (.L_LO(net176));
 sg13g2_sdfbbp_1 \proj_14.flop22/dffsr  (.Q(\proj_14.net165 ),
    .Q_N(\proj_14.net166 ),
    .RESET_B(\proj_14.flop22/_0_ ),
    .SET_B(\proj_14.flop22/_1_ ),
    .D(\proj_14.net163 ),
    .SCE(net175),
    .SCD(net174),
    .CLK(net52));
 sg13g2_inv_1 \proj_14.flop23/_4_  (.Y(\proj_14.flop23/_1_ ),
    .A(net55));
 sg13g2_inv_1 \proj_14.flop23/_5_  (.Y(\proj_14.flop23/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop23/dffsr_168  (.L_LO(net177));
 sg13g2_tielo \proj_14.flop24/dffsr_169  (.L_LO(net178));
 sg13g2_sdfbbp_1 \proj_14.flop23/dffsr  (.Q(\proj_14.net170 ),
    .Q_N(\proj_14.net171 ),
    .RESET_B(\proj_14.flop23/_0_ ),
    .SET_B(\proj_14.flop23/_1_ ),
    .D(\proj_14.net168 ),
    .SCE(net177),
    .SCD(net176),
    .CLK(net54));
 sg13g2_inv_1 \proj_14.flop24/_4_  (.Y(\proj_14.flop24/_1_ ),
    .A(net57));
 sg13g2_inv_1 \proj_14.flop24/_5_  (.Y(\proj_14.flop24/_0_ ),
    .A(\proj_14.net104 ));
 sg13g2_tielo \proj_14.flop24/dffsr_170  (.L_LO(net179));
 sg13g2_tielo \proj_14.flop25/dffsr_171  (.L_LO(net180));
 sg13g2_sdfbbp_1 \proj_14.flop24/dffsr  (.Q(\proj_14.net175 ),
    .Q_N(\proj_14.net176 ),
    .RESET_B(\proj_14.flop24/_0_ ),
    .SET_B(\proj_14.flop24/_1_ ),
    .D(\proj_14.net173 ),
    .SCE(net179),
    .SCD(net178),
    .CLK(net56));
 sg13g2_inv_1 \proj_14.flop25/_4_  (.Y(\proj_14.flop25/_1_ ),
    .A(net59));
 sg13g2_inv_1 \proj_14.flop25/_5_  (.Y(\proj_14.flop25/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop25/dffsr_172  (.L_LO(net181));
 sg13g2_tielo \proj_14.flop26/dffsr_173  (.L_LO(net182));
 sg13g2_sdfbbp_1 \proj_14.flop25/dffsr  (.Q(\proj_14.net180 ),
    .Q_N(\proj_14.flop25/notq ),
    .RESET_B(\proj_14.flop25/_0_ ),
    .SET_B(\proj_14.flop25/_1_ ),
    .D(\proj_14.net178 ),
    .SCE(net181),
    .SCD(net180),
    .CLK(net58));
 sg13g2_inv_1 \proj_14.flop26/_4_  (.Y(\proj_14.flop26/_1_ ),
    .A(net61));
 sg13g2_inv_1 \proj_14.flop26/_5_  (.Y(\proj_14.flop26/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop26/dffsr_174  (.L_LO(net183));
 sg13g2_tielo \proj_14.flop27/dffsr_175  (.L_LO(net184));
 sg13g2_sdfbbp_1 \proj_14.flop26/dffsr  (.Q(\proj_14.net181 ),
    .Q_N(\proj_14.flop26/notq ),
    .RESET_B(\proj_14.flop26/_0_ ),
    .SET_B(\proj_14.flop26/_1_ ),
    .D(\proj_14.net180 ),
    .SCE(net183),
    .SCD(net182),
    .CLK(net60));
 sg13g2_inv_1 \proj_14.flop27/_4_  (.Y(\proj_14.flop27/_1_ ),
    .A(net63));
 sg13g2_inv_1 \proj_14.flop27/_5_  (.Y(\proj_14.flop27/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop27/dffsr_176  (.L_LO(net185));
 sg13g2_tielo \proj_14.flop29/dffsr_177  (.L_LO(net186));
 sg13g2_sdfbbp_1 \proj_14.flop27/dffsr  (.Q(\proj_14.flop27/q ),
    .Q_N(\proj_14.net182 ),
    .RESET_B(\proj_14.flop27/_0_ ),
    .SET_B(\proj_14.flop27/_1_ ),
    .D(\proj_14.net181 ),
    .SCE(net185),
    .SCD(net184),
    .CLK(net62));
 sg13g2_dfrbp_1 \proj_14.flop28/_1_  (.CLK(net64),
    .RESET_B(net240),
    .D(\proj_14.net95 ),
    .Q_N(\proj_14.flop28/notq ),
    .Q(\proj_14.net11 ));
 sg13g2_tiehi \proj_14.flop46/_1__232  (.L_HI(net241));
 sg13g2_inv_1 \proj_14.flop29/_4_  (.Y(\proj_14.flop29/_1_ ),
    .A(net66));
 sg13g2_inv_1 \proj_14.flop29/_5_  (.Y(\proj_14.flop29/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop29/dffsr_178  (.L_LO(net187));
 sg13g2_tielo \proj_14.flop3/dffsr_179  (.L_LO(net188));
 sg13g2_sdfbbp_1 \proj_14.flop29/dffsr  (.Q(\proj_14.net209 ),
    .Q_N(\proj_14.net210 ),
    .RESET_B(\proj_14.flop29/_0_ ),
    .SET_B(\proj_14.flop29/_1_ ),
    .D(\proj_14.net207 ),
    .SCE(net187),
    .SCD(net186),
    .CLK(net65));
 sg13g2_inv_1 \proj_14.flop3/_4_  (.Y(\proj_14.flop3/_1_ ),
    .A(net68));
 sg13g2_inv_1 \proj_14.flop3/_5_  (.Y(\proj_14.flop3/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop3/dffsr_180  (.L_LO(net189));
 sg13g2_tielo \proj_14.flop30/dffsr_181  (.L_LO(net190));
 sg13g2_sdfbbp_1 \proj_14.flop3/dffsr  (.Q(\proj_14.net32 ),
    .Q_N(\proj_14.net33 ),
    .RESET_B(\proj_14.flop3/_0_ ),
    .SET_B(\proj_14.flop3/_1_ ),
    .D(\proj_14.net31 ),
    .SCE(net189),
    .SCD(net188),
    .CLK(net67));
 sg13g2_inv_1 \proj_14.flop30/_4_  (.Y(\proj_14.flop30/_1_ ),
    .A(net70));
 sg13g2_inv_1 \proj_14.flop30/_5_  (.Y(\proj_14.flop30/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop30/dffsr_182  (.L_LO(net191));
 sg13g2_tielo \proj_14.flop31/dffsr_183  (.L_LO(net192));
 sg13g2_sdfbbp_1 \proj_14.flop30/dffsr  (.Q(\proj_14.net214 ),
    .Q_N(\proj_14.net215 ),
    .RESET_B(\proj_14.flop30/_0_ ),
    .SET_B(\proj_14.flop30/_1_ ),
    .D(\proj_14.net212 ),
    .SCE(net191),
    .SCD(net190),
    .CLK(net69));
 sg13g2_inv_1 \proj_14.flop31/_4_  (.Y(\proj_14.flop31/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop31/_5_  (.Y(\proj_14.flop31/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop31/dffsr_184  (.L_LO(net193));
 sg13g2_tielo \proj_14.flop32/dffsr_185  (.L_LO(net194));
 sg13g2_sdfbbp_1 \proj_14.flop31/dffsr  (.Q(\proj_14.net217 ),
    .Q_N(\proj_14.flop31/notq ),
    .RESET_B(\proj_14.flop31/_0_ ),
    .SET_B(\proj_14.flop31/_1_ ),
    .D(\proj_14.net216 ),
    .SCE(net193),
    .SCD(net192),
    .CLK(net71));
 sg13g2_inv_1 \proj_14.flop32/_4_  (.Y(\proj_14.flop32/_1_ ),
    .A(net73));
 sg13g2_inv_1 \proj_14.flop32/_5_  (.Y(\proj_14.flop32/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop32/dffsr_186  (.L_LO(net195));
 sg13g2_tielo \proj_14.flop33/dffsr_187  (.L_LO(net196));
 sg13g2_sdfbbp_1 \proj_14.flop32/dffsr  (.Q(\proj_14.net219 ),
    .Q_N(\proj_14.flop32/notq ),
    .RESET_B(\proj_14.flop32/_0_ ),
    .SET_B(\proj_14.flop32/_1_ ),
    .D(\proj_14.net218 ),
    .SCE(net195),
    .SCD(net194),
    .CLK(net72));
 sg13g2_inv_1 \proj_14.flop33/_4_  (.Y(\proj_14.flop33/_1_ ),
    .A(net75));
 sg13g2_inv_1 \proj_14.flop33/_5_  (.Y(\proj_14.flop33/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop33/dffsr_188  (.L_LO(net197));
 sg13g2_tielo \proj_14.flop34/dffsr_189  (.L_LO(net198));
 sg13g2_sdfbbp_1 \proj_14.flop33/dffsr  (.Q(\proj_14.net221 ),
    .Q_N(\proj_14.flop33/notq ),
    .RESET_B(\proj_14.flop33/_0_ ),
    .SET_B(\proj_14.flop33/_1_ ),
    .D(\proj_14.net220 ),
    .SCE(net197),
    .SCD(net196),
    .CLK(net74));
 sg13g2_inv_1 \proj_14.flop34/_4_  (.Y(\proj_14.flop34/_1_ ),
    .A(net77));
 sg13g2_inv_1 \proj_14.flop34/_5_  (.Y(\proj_14.flop34/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop34/dffsr_190  (.L_LO(net199));
 sg13g2_tielo \proj_14.flop35/dffsr_191  (.L_LO(net200));
 sg13g2_sdfbbp_1 \proj_14.flop34/dffsr  (.Q(\proj_14.net223 ),
    .Q_N(\proj_14.flop34/notq ),
    .RESET_B(\proj_14.flop34/_0_ ),
    .SET_B(\proj_14.flop34/_1_ ),
    .D(\proj_14.net222 ),
    .SCE(net199),
    .SCD(net198),
    .CLK(net76));
 sg13g2_inv_1 \proj_14.flop35/_4_  (.Y(\proj_14.flop35/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop35/_5_  (.Y(\proj_14.flop35/_0_ ),
    .A(net79));
 sg13g2_tielo \proj_14.flop35/dffsr_192  (.L_LO(net201));
 sg13g2_tielo \proj_14.flop36/dffsr_193  (.L_LO(net202));
 sg13g2_sdfbbp_1 \proj_14.flop35/dffsr  (.Q(\proj_14.net226 ),
    .Q_N(\proj_14.flop35/notq ),
    .RESET_B(\proj_14.flop35/_0_ ),
    .SET_B(\proj_14.flop35/_1_ ),
    .D(\proj_14.net224 ),
    .SCE(net201),
    .SCD(net200),
    .CLK(net78));
 sg13g2_inv_1 \proj_14.flop36/_4_  (.Y(\proj_14.flop36/_1_ ),
    .A(net81));
 sg13g2_inv_1 \proj_14.flop36/_5_  (.Y(\proj_14.flop36/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop36/dffsr_194  (.L_LO(net203));
 sg13g2_tielo \proj_14.flop37/dffsr_195  (.L_LO(net204));
 sg13g2_sdfbbp_1 \proj_14.flop36/dffsr  (.Q(\proj_14.net228 ),
    .Q_N(\proj_14.flop36/notq ),
    .RESET_B(\proj_14.flop36/_0_ ),
    .SET_B(\proj_14.flop36/_1_ ),
    .D(\proj_14.net227 ),
    .SCE(net203),
    .SCD(net202),
    .CLK(net80));
 sg13g2_inv_1 \proj_14.flop37/_4_  (.Y(\proj_14.flop37/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop37/_5_  (.Y(\proj_14.flop37/_0_ ),
    .A(net83));
 sg13g2_tielo \proj_14.flop37/dffsr_196  (.L_LO(net205));
 sg13g2_tielo \proj_14.flop4/dffsr_197  (.L_LO(net206));
 sg13g2_sdfbbp_1 \proj_14.flop37/dffsr  (.Q(\proj_14.net231 ),
    .Q_N(\proj_14.flop37/notq ),
    .RESET_B(\proj_14.flop37/_0_ ),
    .SET_B(\proj_14.flop37/_1_ ),
    .D(\proj_14.net229 ),
    .SCE(net205),
    .SCD(net204),
    .CLK(net82));
 sg13g2_inv_1 \proj_14.flop4/_4_  (.Y(\proj_14.flop4/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop4/_5_  (.Y(\proj_14.flop4/_0_ ),
    .A(net85));
 sg13g2_tielo \proj_14.flop4/dffsr_198  (.L_LO(net207));
 sg13g2_tielo \proj_14.flop5/dffsr_199  (.L_LO(net208));
 sg13g2_sdfbbp_1 \proj_14.flop4/dffsr  (.Q(\proj_14.net36 ),
    .Q_N(\proj_14.net37 ),
    .RESET_B(\proj_14.flop4/_0_ ),
    .SET_B(\proj_14.flop4/_1_ ),
    .D(\proj_14.net34 ),
    .SCE(net207),
    .SCD(net206),
    .CLK(net84));
 sg13g2_dfrbp_1 \proj_14.flop46/_1_  (.CLK(net86),
    .RESET_B(net241),
    .D(\proj_14.net96 ),
    .Q_N(\proj_14.flop46/notq ),
    .Q(\proj_14.net12 ));
 sg13g2_tiehi \proj_14.flop47/_1__233  (.L_HI(net242));
 sg13g2_dfrbp_1 \proj_14.flop47/_1_  (.CLK(net87),
    .RESET_B(net242),
    .D(\proj_14.net97 ),
    .Q_N(\proj_14.flop47/notq ),
    .Q(\proj_14.net13 ));
 sg13g2_tiehi \proj_14.flop48/_1__234  (.L_HI(net243));
 sg13g2_dfrbp_1 \proj_14.flop48/_1_  (.CLK(net88),
    .RESET_B(net243),
    .D(\proj_14.net98 ),
    .Q_N(\proj_14.flop48/notq ),
    .Q(\proj_14.net14 ));
 sg13g2_tiehi \proj_14.flop49/_1__235  (.L_HI(net244));
 sg13g2_dfrbp_1 \proj_14.flop49/_1_  (.CLK(net89),
    .RESET_B(net244),
    .D(\proj_14.net99 ),
    .Q_N(\proj_14.flop49/notq ),
    .Q(\proj_14.net15 ));
 sg13g2_tiehi \proj_14.flop50/_1__236  (.L_HI(net245));
 sg13g2_inv_1 \proj_14.flop5/_4_  (.Y(\proj_14.flop5/_1_ ),
    .A(net91));
 sg13g2_inv_1 \proj_14.flop5/_5_  (.Y(\proj_14.flop5/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop5/dffsr_200  (.L_LO(net209));
 sg13g2_tielo \proj_14.flop6/dffsr_201  (.L_LO(net210));
 sg13g2_sdfbbp_1 \proj_14.flop5/dffsr  (.Q(\proj_14.net39 ),
    .Q_N(\proj_14.net40 ),
    .RESET_B(\proj_14.flop5/_0_ ),
    .SET_B(\proj_14.flop5/_1_ ),
    .D(\proj_14.net38 ),
    .SCE(net209),
    .SCD(net208),
    .CLK(net90));
 sg13g2_dfrbp_1 \proj_14.flop50/_1_  (.CLK(net92),
    .RESET_B(net245),
    .D(\proj_14.net100 ),
    .Q_N(\proj_14.flop50/notq ),
    .Q(\proj_14.net16 ));
 sg13g2_tiehi \proj_14.flop51/_1__237  (.L_HI(net246));
 sg13g2_dfrbp_1 \proj_14.flop51/_1_  (.CLK(net93),
    .RESET_B(net246),
    .D(\proj_14.net101 ),
    .Q_N(\proj_14.flop51/notq ),
    .Q(\proj_14.net17 ));
 sg13g2_tiehi \proj_14.flop52/_1__238  (.L_HI(net247));
 sg13g2_dfrbp_1 \proj_14.flop52/_1_  (.CLK(net94),
    .RESET_B(net247),
    .D(\proj_14.net183 ),
    .Q_N(\proj_14.flop52/notq ),
    .Q(\proj_14.net45 ));
 sg13g2_tiehi \proj_14.flop53/_1__239  (.L_HI(net248));
 sg13g2_dfrbp_1 \proj_14.flop53/_1_  (.CLK(net95),
    .RESET_B(net248),
    .D(\proj_14.net275 ),
    .Q_N(\proj_14.flop53/notq ),
    .Q(\proj_14.net44 ));
 sg13g2_tiehi \proj_14.flop54/_1__240  (.L_HI(net249));
 sg13g2_dfrbp_1 \proj_14.flop54/_1_  (.CLK(net96),
    .RESET_B(net249),
    .D(\proj_14.net277 ),
    .Q_N(\proj_14.flop54/notq ),
    .Q(\proj_14.net46 ));
 sg13g2_tiehi \proj_14.flop55/_1__241  (.L_HI(net250));
 sg13g2_dfrbp_1 \proj_14.flop55/_1_  (.CLK(net97),
    .RESET_B(net250),
    .D(\proj_14.net280 ),
    .Q_N(\proj_14.flop55/notq ),
    .Q(\proj_14.net47 ));
 sg13g2_tiehi \proj_14.flop56/_1__242  (.L_HI(net251));
 sg13g2_dfrbp_1 \proj_14.flop56/_1_  (.CLK(net98),
    .RESET_B(net251),
    .D(\proj_14.net281 ),
    .Q_N(\proj_14.flop56/notq ),
    .Q(\proj_14.net211 ));
 sg13g2_tiehi \proj__7.flop1/_1__243  (.L_HI(net252));
 sg13g2_inv_1 \proj_14.flop6/_4_  (.Y(\proj_14.flop6/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop6/_5_  (.Y(\proj_14.flop6/_0_ ),
    .A(net100));
 sg13g2_tielo \proj_14.flop6/dffsr_202  (.L_LO(net211));
 sg13g2_tielo \proj_14.flop7/dffsr_203  (.L_LO(net212));
 sg13g2_sdfbbp_1 \proj_14.flop6/dffsr  (.Q(\proj_14.net42 ),
    .Q_N(\proj_14.net43 ),
    .RESET_B(\proj_14.flop6/_0_ ),
    .SET_B(\proj_14.flop6/_1_ ),
    .D(\proj_14.net41 ),
    .SCE(net211),
    .SCD(net210),
    .CLK(net99));
 sg13g2_inv_1 \proj_14.flop7/_4_  (.Y(\proj_14.flop7/_1_ ),
    .A(net102));
 sg13g2_inv_1 \proj_14.flop7/_5_  (.Y(\proj_14.flop7/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop7/dffsr_204  (.L_LO(net213));
 sg13g2_tielo \proj_14.flop8/dffsr_205  (.L_LO(net214));
 sg13g2_sdfbbp_1 \proj_14.flop7/dffsr  (.Q(\proj_14.net50 ),
    .Q_N(\proj_14.net51 ),
    .RESET_B(\proj_14.flop7/_0_ ),
    .SET_B(\proj_14.flop7/_1_ ),
    .D(\proj_14.net48 ),
    .SCE(net213),
    .SCD(net212),
    .CLK(net101));
 sg13g2_inv_1 \proj_14.flop8/_4_  (.Y(\proj_14.flop8/_1_ ),
    .A(net104));
 sg13g2_inv_1 \proj_14.flop8/_5_  (.Y(\proj_14.flop8/_0_ ),
    .A(\proj_14.net25 ));
 sg13g2_tielo \proj_14.flop8/dffsr_206  (.L_LO(net215));
 sg13g2_tielo \proj_14.flop9/dffsr_207  (.L_LO(net216));
 sg13g2_sdfbbp_1 \proj_14.flop8/dffsr  (.Q(\proj_14.net53 ),
    .Q_N(\proj_14.net54 ),
    .RESET_B(\proj_14.flop8/_0_ ),
    .SET_B(\proj_14.flop8/_1_ ),
    .D(\proj_14.net52 ),
    .SCE(net215),
    .SCD(net214),
    .CLK(net103));
 sg13g2_inv_1 \proj_14.flop9/_4_  (.Y(\proj_14.flop9/_1_ ),
    .A(\proj_14.net25 ));
 sg13g2_inv_1 \proj_14.flop9/_5_  (.Y(\proj_14.flop9/_0_ ),
    .A(net106));
 sg13g2_tielo \proj_14.flop9/dffsr_208  (.L_LO(net217));
 sg13g2_tielo \proj__4.flop1/dffsr_209  (.L_LO(net218));
 sg13g2_sdfbbp_1 \proj_14.flop9/dffsr  (.Q(\proj_14.net56 ),
    .Q_N(\proj_14.net57 ),
    .RESET_B(\proj_14.flop9/_0_ ),
    .SET_B(\proj_14.flop9/_1_ ),
    .D(\proj_14.net55 ),
    .SCE(net217),
    .SCD(net216),
    .CLK(net105));
 sg13g2_mux2_1 \proj_14.mux1/_0_  (.A0(\proj_14.net23 ),
    .A1(\proj_14.net44 ),
    .S(net43),
    .X(\proj_14.net23 ));
 sg13g2_mux2_1 \proj_14.mux10/_0_  (.A0(\proj_14.net105 ),
    .A1(\proj_14.net106 ),
    .S(net236),
    .X(\proj_14.net102 ));
 sg13g2_mux2_1 \proj_14.mux11/_0_  (.A0(\proj_14.net110 ),
    .A1(\proj_14.net111 ),
    .S(\proj_14.net105 ),
    .X(\proj_14.net108 ));
 sg13g2_mux2_1 \proj_14.mux12/_0_  (.A0(\proj_14.net114 ),
    .A1(\proj_14.net115 ),
    .S(\proj_14.net116 ),
    .X(\proj_14.net112 ));
 sg13g2_mux2_1 \proj_14.mux13/_0_  (.A0(\proj_14.net119 ),
    .A1(\proj_14.net120 ),
    .S(\proj_14.net121 ),
    .X(\proj_14.net117 ));
 sg13g2_mux2_1 \proj_14.mux14/_0_  (.A0(\proj_14.net124 ),
    .A1(\proj_14.net125 ),
    .S(\proj_14.net126 ),
    .X(\proj_14.net122 ));
 sg13g2_mux2_1 \proj_14.mux15/_0_  (.A0(\proj_14.net129 ),
    .A1(\proj_14.net130 ),
    .S(\proj_14.net131 ),
    .X(\proj_14.net127 ));
 sg13g2_mux2_1 \proj_14.mux16/_0_  (.A0(\proj_14.net135 ),
    .A1(\proj_14.net136 ),
    .S(\proj_14.net137 ),
    .X(\proj_14.net133 ));
 sg13g2_mux2_1 \proj_14.mux17/_0_  (.A0(\proj_14.net140 ),
    .A1(\proj_14.net141 ),
    .S(\proj_14.net142 ),
    .X(\proj_14.net138 ));
 sg13g2_mux2_1 \proj_14.mux18/_0_  (.A0(\proj_14.net145 ),
    .A1(\proj_14.net146 ),
    .S(\proj_14.net147 ),
    .X(\proj_14.net143 ));
 sg13g2_mux2_1 \proj_14.mux19/_0_  (.A0(\proj_14.net150 ),
    .A1(\proj_14.net151 ),
    .S(\proj_14.net152 ),
    .X(\proj_14.net148 ));
 sg13g2_mux2_1 \proj_14.mux2/_0_  (.A0(\proj_14.net28 ),
    .A1(\proj_14.net46 ),
    .S(net43),
    .X(\proj_14.net28 ));
 sg13g2_mux2_1 \proj_14.mux20/_0_  (.A0(\proj_14.net155 ),
    .A1(\proj_14.net156 ),
    .S(\proj_14.net157 ),
    .X(\proj_14.net153 ));
 sg13g2_mux2_1 \proj_14.mux21/_0_  (.A0(\proj_14.net160 ),
    .A1(\proj_14.net161 ),
    .S(\proj_14.net162 ),
    .X(\proj_14.net158 ));
 sg13g2_mux2_1 \proj_14.mux22/_0_  (.A0(\proj_14.net165 ),
    .A1(\proj_14.net166 ),
    .S(\proj_14.net167 ),
    .X(\proj_14.net163 ));
 sg13g2_mux2_1 \proj_14.mux23/_0_  (.A0(\proj_14.net170 ),
    .A1(\proj_14.net171 ),
    .S(\proj_14.net172 ),
    .X(\proj_14.net168 ));
 sg13g2_mux2_1 \proj_14.mux24/_0_  (.A0(\proj_14.net175 ),
    .A1(\proj_14.net176 ),
    .S(\proj_14.net177 ),
    .X(\proj_14.net173 ));
 sg13g2_mux2_1 \proj_14.mux25/_0_  (.A0(\proj_14.net209 ),
    .A1(\proj_14.net211 ),
    .S(net43),
    .X(\proj_14.net207 ));
 sg13g2_mux2_1 \proj_14.mux26/_0_  (.A0(\proj_14.net214 ),
    .A1(\proj_14.net233 ),
    .S(net42),
    .X(\proj_14.net212 ));
 sg13g2_mux2_1 \proj_14.mux27/_0_  (.A0(\proj_14.net217 ),
    .A1(\proj_14.net214 ),
    .S(net42),
    .X(\proj_14.net216 ));
 sg13g2_mux2_1 \proj_14.mux28/_0_  (.A0(\proj_14.net219 ),
    .A1(\proj_14.net217 ),
    .S(net42),
    .X(\proj_14.net218 ));
 sg13g2_mux2_1 \proj_14.mux29/_0_  (.A0(\proj_14.net221 ),
    .A1(\proj_14.net219 ),
    .S(net42),
    .X(\proj_14.net220 ));
 sg13g2_mux2_1 \proj_14.mux3/_0_  (.A0(\proj_14.net31 ),
    .A1(\proj_14.net47 ),
    .S(net43),
    .X(\proj_14.net31 ));
 sg13g2_mux2_1 \proj_14.mux30/_0_  (.A0(\proj_14.net223 ),
    .A1(\proj_14.net221 ),
    .S(net42),
    .X(\proj_14.net222 ));
 sg13g2_mux2_1 \proj_14.mux31/_0_  (.A0(\proj_14.net226 ),
    .A1(\proj_14.net223 ),
    .S(net42),
    .X(\proj_14.net224 ));
 sg13g2_mux2_1 \proj_14.mux32/_0_  (.A0(\proj_14.net228 ),
    .A1(\proj_14.net226 ),
    .S(net42),
    .X(\proj_14.net227 ));
 sg13g2_mux2_1 \proj_14.mux33/_0_  (.A0(\proj_14.net231 ),
    .A1(\proj_14.net228 ),
    .S(net42),
    .X(\proj_14.net229 ));
 sg13g2_mux2_1 \proj_14.mux4/_0_  (.A0(\proj_14.net34 ),
    .A1(\proj_14.net26 ),
    .S(net43),
    .X(\proj_14.net34 ));
 sg13g2_mux2_1 \proj_14.mux5/_0_  (.A0(\proj_14.net38 ),
    .A1(\proj_14.net29 ),
    .S(\proj_14.net45 ),
    .X(\proj_14.net38 ));
 sg13g2_mux2_1 \proj_14.mux6/_0_  (.A0(\proj_14.net41 ),
    .A1(\proj_14.net32 ),
    .S(net43),
    .X(\proj_14.net41 ));
 sg13g2_mux2_1 \proj_14.mux7/_0_  (.A0(\proj_14.net48 ),
    .A1(\proj_14.net36 ),
    .S(net43),
    .X(\proj_14.net48 ));
 sg13g2_mux2_1 \proj_14.mux8/_0_  (.A0(\proj_14.net52 ),
    .A1(\proj_14.net39 ),
    .S(\proj_14.net45 ),
    .X(\proj_14.net52 ));
 sg13g2_mux2_1 \proj_14.mux9/_0_  (.A0(\proj_14.net55 ),
    .A1(\proj_14.net42 ),
    .S(\proj_14.net45 ),
    .X(\proj_14.net55 ));
 sg13g2_inv_1 \proj_14.not1/_0_  (.Y(\proj_14.net132 ),
    .A(net107));
 sg13g2_inv_1 \proj_14.not10/_0_  (.Y(\proj_14.net193 ),
    .A(\proj_14.net190 ));
 sg13g2_inv_1 \proj_14.not2/_0_  (.Y(\proj_14.net202 ),
    .A(\proj_14.net184 ));
 sg13g2_inv_1 \proj_14.not3/_0_  (.Y(\proj_14.net201 ),
    .A(\proj_14.net185 ));
 sg13g2_inv_1 \proj_14.not4/_0_  (.Y(\proj_14.net198 ),
    .A(\proj_14.net187 ));
 sg13g2_inv_1 \proj_14.not5/_0_  (.Y(\proj_14.net25 ),
    .A(net108));
 sg13g2_inv_1 \proj_14.not6/_0_  (.Y(\proj_14.net199 ),
    .A(\proj_14.net186 ));
 sg13g2_inv_1 \proj_14.not7/_0_  (.Y(\proj_14.net195 ),
    .A(\proj_14.net189 ));
 sg13g2_inv_1 \proj_14.not8/_0_  (.Y(\proj_14.net196 ),
    .A(\proj_14.net188 ));
 sg13g2_inv_1 \proj_14.not9/_0_  (.Y(\proj_14.net192 ),
    .A(\proj_14.net191 ));
 sg13g2_or2_1 \proj_14.or1/_0_  (.X(\proj_14.net104 ),
    .B(\proj_14.net132 ),
    .A(\proj_14.net183 ));
 sg13g2_or2_1 \proj_14.or10/_0_  (.X(\proj_14.net96 ),
    .B(\proj_14.net60 ),
    .A(\proj_14.net89 ));
 sg13g2_or2_1 \proj_14.or11/_0_  (.X(\proj_14.net97 ),
    .B(\proj_14.net62 ),
    .A(\proj_14.net90 ));
 sg13g2_or2_1 \proj_14.or12/_0_  (.X(\proj_14.net98 ),
    .B(\proj_14.net63 ),
    .A(\proj_14.net91 ));
 sg13g2_or2_1 \proj_14.or13/_0_  (.X(\proj_14.net99 ),
    .B(\proj_14.net65 ),
    .A(\proj_14.net92 ));
 sg13g2_or2_1 \proj_14.or14/_0_  (.X(\proj_14.net100 ),
    .B(\proj_14.net66 ),
    .A(\proj_14.net93 ));
 sg13g2_or2_1 \proj_14.or15/_0_  (.X(\proj_14.net101 ),
    .B(\proj_14.net67 ),
    .A(\proj_14.net94 ));
 sg13g2_or2_1 \proj_14.or16/_0_  (.X(\proj_14.net247 ),
    .B(\proj_14.net236 ),
    .A(\proj_14.net234 ));
 sg13g2_or2_1 \proj_14.or17/_0_  (.X(\proj_14.net250 ),
    .B(\proj_14.net248 ),
    .A(\proj_14.net249 ));
 sg13g2_or2_1 \proj_14.or18/_0_  (.X(\proj_14.net255 ),
    .B(\proj_14.net254 ),
    .A(\proj_14.net252 ));
 sg13g2_or2_1 \proj_14.or19/_0_  (.X(\proj_14.net251 ),
    .B(\proj_14.net237 ),
    .A(\proj_14.net248 ));
 sg13g2_or2_1 \proj_14.or2/_0_  (.X(\proj_14.net95 ),
    .B(\proj_14.net59 ),
    .A(\proj_14.net88 ));
 sg13g2_or2_1 \proj_14.or20/_0_  (.X(\proj_14.net253 ),
    .B(\proj_14.net252 ),
    .A(\proj_14.net236 ));
 sg13g2_or2_1 \proj_14.or21/_0_  (.X(\proj_14.net257 ),
    .B(\proj_14.net254 ),
    .A(\proj_14.net256 ));
 sg13g2_or2_1 \proj_14.or22/_0_  (.X(\proj_14.net272 ),
    .B(\proj_14.net253 ),
    .A(\proj_14.net250 ));
 sg13g2_or2_1 \proj_14.or23/_0_  (.X(\proj_14.net287 ),
    .B(\proj_14.net285 ),
    .A(\proj_14.net286 ));
 sg13g2_or2_1 \proj_14.or24/_0_  (.X(\proj_14.net260 ),
    .B(\proj_14.net259 ),
    .A(\proj_14.net240 ));
 sg13g2_or2_1 \proj_14.or25/_0_  (.X(\proj_14.net262 ),
    .B(\proj_14.net261 ),
    .A(\proj_14.net240 ));
 sg13g2_or2_1 \proj_14.or26/_0_  (.X(\proj_14.net263 ),
    .B(\proj_14.net243 ),
    .A(\proj_14.net261 ));
 sg13g2_or2_1 \proj_14.or27/_0_  (.X(\proj_14.net264 ),
    .B(\proj_14.net251 ),
    .A(\proj_14.net245 ));
 sg13g2_or2_1 \proj_14.or28/_0_  (.X(\proj_14.net266 ),
    .B(\proj_14.net244 ),
    .A(\proj_14.net265 ));
 sg13g2_or2_1 \proj_14.or29/_0_  (.X(\proj_14.net268 ),
    .B(\proj_14.net244 ),
    .A(\proj_14.net267 ));
 sg13g2_or2_1 \proj_14.or3/_0_  (.X(\proj_14.net88 ),
    .B(\proj_14.net69 ),
    .A(\proj_14.net79 ));
 sg13g2_or2_1 \proj_14.or30/_0_  (.X(\proj_14.net273 ),
    .B(\proj_14.net266 ),
    .A(\proj_14.net260 ));
 sg13g2_or2_1 \proj_14.or31/_0_  (.X(\proj_14.net270 ),
    .B(\proj_14.net269 ),
    .A(\proj_14.net268 ));
 sg13g2_or2_1 \proj_14.or32/_0_  (.X(\proj_14.net271 ),
    .B(\proj_14.net256 ),
    .A(\proj_14.net258 ));
 sg13g2_or2_1 \proj_14.or33/_0_  (.X(\proj_14.net274 ),
    .B(\proj_14.net257 ),
    .A(\proj_14.net247 ));
 sg13g2_or2_1 \proj_14.or34/_0_  (.X(\proj_14.net275 ),
    .B(\proj_14.net273 ),
    .A(\proj_14.net274 ));
 sg13g2_or2_1 \proj_14.or35/_0_  (.X(\proj_14.net276 ),
    .B(\proj_14.net263 ),
    .A(\proj_14.net272 ));
 sg13g2_or2_1 \proj_14.or36/_0_  (.X(\proj_14.net277 ),
    .B(\proj_14.net270 ),
    .A(\proj_14.net276 ));
 sg13g2_or2_1 \proj_14.or37/_0_  (.X(\proj_14.net278 ),
    .B(\proj_14.net271 ),
    .A(\proj_14.net262 ));
 sg13g2_or2_1 \proj_14.or38/_0_  (.X(\proj_14.net279 ),
    .B(\proj_14.net255 ),
    .A(\proj_14.net264 ));
 sg13g2_or2_1 \proj_14.or39/_0_  (.X(\proj_14.net280 ),
    .B(\proj_14.net278 ),
    .A(\proj_14.net279 ));
 sg13g2_or2_1 \proj_14.or4/_0_  (.X(\proj_14.net89 ),
    .B(\proj_14.net70 ),
    .A(\proj_14.net80 ));
 sg13g2_or2_1 \proj_14.or40/_0_  (.X(\proj_14.net283 ),
    .B(\proj_14.net240 ),
    .A(\proj_14.net241 ));
 sg13g2_or2_1 \proj_14.or41/_0_  (.X(\proj_14.net284 ),
    .B(\proj_14.net243 ),
    .A(\proj_14.net244 ));
 sg13g2_or2_1 \proj_14.or42/_0_  (.X(\proj_14.net285 ),
    .B(\proj_14.net283 ),
    .A(\proj_14.net284 ));
 sg13g2_or2_1 \proj_14.or43/_0_  (.X(\proj_14.net286 ),
    .B(\proj_14.net259 ),
    .A(\proj_14.net258 ));
 sg13g2_or2_1 \proj_14.or44/_0_  (.X(\proj_14.net288 ),
    .B(\proj_14.net265 ),
    .A(\proj_14.net252 ));
 sg13g2_or2_1 \proj_14.or45/_0_  (.X(\proj_14.net281 ),
    .B(\proj_14.net287 ),
    .A(\proj_14.net289 ));
 sg13g2_or2_1 \proj_14.or46/_0_  (.X(\proj_14.net289 ),
    .B(\proj_14.net245 ),
    .A(\proj_14.net288 ));
 sg13g2_or2_1 \proj_14.or5/_0_  (.X(\proj_14.net90 ),
    .B(\proj_14.net72 ),
    .A(\proj_14.net82 ));
 sg13g2_or2_1 \proj_14.or6/_0_  (.X(\proj_14.net91 ),
    .B(\proj_14.net73 ),
    .A(\proj_14.net83 ));
 sg13g2_or2_1 \proj_14.or7/_0_  (.X(\proj_14.net92 ),
    .B(\proj_14.net75 ),
    .A(\proj_14.net85 ));
 sg13g2_or2_1 \proj_14.or8/_0_  (.X(\proj_14.net93 ),
    .B(\proj_14.net76 ),
    .A(\proj_14.net86 ));
 sg13g2_or2_1 \proj_14.or9/_0_  (.X(\proj_14.net94 ),
    .B(\proj_14.net77 ),
    .A(\proj_14.net87 ));
 sg13g2_xor2_1 \proj_14.xor1/_0_  (.B(net7),
    .A(\proj_14.net175 ),
    .X(\proj_14.net184 ));
 sg13g2_xor2_1 \proj_14.xor10/_0_  (.B(\proj_14.net226 ),
    .A(\proj_14.net231 ),
    .X(\proj_14.net282 ));
 sg13g2_xor2_1 \proj_14.xor11/_0_  (.B(\proj_14.net221 ),
    .A(\proj_14.net232 ),
    .X(\proj_14.net233 ));
 sg13g2_xor2_1 \proj_14.xor2/_0_  (.B(net6),
    .A(\proj_14.net170 ),
    .X(\proj_14.net185 ));
 sg13g2_xor2_1 \proj_14.xor3/_0_  (.B(net5),
    .A(\proj_14.net165 ),
    .X(\proj_14.net186 ));
 sg13g2_xor2_1 \proj_14.xor4/_0_  (.B(net4),
    .A(\proj_14.net160 ),
    .X(\proj_14.net187 ));
 sg13g2_xor2_1 \proj_14.xor5/_0_  (.B(net3),
    .A(\proj_14.net155 ),
    .X(\proj_14.net188 ));
 sg13g2_xor2_1 \proj_14.xor6/_0_  (.B(net2),
    .A(\proj_14.net150 ),
    .X(\proj_14.net189 ));
 sg13g2_xor2_1 \proj_14.xor7/_0_  (.B(net39),
    .A(\proj_14.net145 ),
    .X(\proj_14.net190 ));
 sg13g2_xor2_1 \proj_14.xor8/_0_  (.B(net41),
    .A(\proj_14.net140 ),
    .X(\proj_14.net191 ));
 sg13g2_xor2_1 \proj_14.xor9/_0_  (.B(\proj_14.net223 ),
    .A(\proj_14.net282 ),
    .X(\proj_14.net232 ));
 sg13g2_inv_1 \proj__0.not3/_0_  (.Y(\proj__0.net10 ),
    .A(net37));
 sg13g2_inv_1 \proj__0.not4/_0_  (.Y(\proj__0.net11 ),
    .A(net36));
 sg13g2_xor2_1 \proj__0.xor1/_0_  (.B(net40),
    .A(net38),
    .X(\proj__0.net9 ));
 sg13g2_and2_1 \proj__1.and1/_0_  (.A(\proj__1.net18 ),
    .B(net41),
    .X(\proj__1.net19 ));
 sg13g2_and2_1 \proj__1.and2/_0_  (.A(\proj__1.net16 ),
    .B(net2),
    .X(\proj__1.net20 ));
 sg13g2_and2_1 \proj__1.and3/_0_  (.A(\proj__1.net10 ),
    .B(net4),
    .X(\proj__1.net21 ));
 sg13g2_and2_1 \proj__1.and4/_0_  (.A(\proj__1.net17 ),
    .B(net6),
    .X(\proj__1.net22 ));
 sg13g2_and2_1 \proj__1.and5/_0_  (.A(\proj__1.net20 ),
    .B(\proj__1.net19 ),
    .X(\proj__1.net23 ));
 sg13g2_and2_1 \proj__1.and6/_0_  (.A(\proj__1.net22 ),
    .B(\proj__1.net21 ),
    .X(\proj__1.net24 ));
 sg13g2_and2_1 \proj__1.and7/_0_  (.A(\proj__1.net24 ),
    .B(\proj__1.net23 ),
    .X(\proj__1.net9 ));
 sg13g2_inv_1 \proj__1.not1/_0_  (.Y(\proj__1.net16 ),
    .A(net3));
 sg13g2_inv_1 \proj__1.not2/_0_  (.Y(\proj__1.net17 ),
    .A(net7));
 sg13g2_inv_1 \proj__1.not3/_0_  (.Y(\proj__1.net18 ),
    .A(net39));
 sg13g2_inv_1 \proj__1.not4/_0_  (.Y(\proj__1.net10 ),
    .A(net35));
 sg13g2_inv_1 \proj__2.not1/_0_  (.Y(\proj__2.net9 ),
    .A(net40));
 sg13g2_inv_1 \proj__2.not2/_0_  (.Y(\proj__2.net10 ),
    .A(net38));
 sg13g2_inv_1 \proj__2.not3/_0_  (.Y(\proj__2.net11 ),
    .A(net37));
 sg13g2_inv_1 \proj__2.not4/_0_  (.Y(\proj__2.net12 ),
    .A(net36));
 sg13g2_and2_1 \proj__3.and3/_0_  (.A(\proj__3.net11 ),
    .B(net40),
    .X(\proj__3.net4 ));
 sg13g2_and2_1 \proj__3.and4/_0_  (.A(net38),
    .B(\proj__3.net12 ),
    .X(\proj__3.net3 ));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net11 ),
    .A(net38));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net12 ),
    .A(net40));
 sg13g2_inv_1 \proj__3.not6/_0_  (.Y(\proj__3.net5 ),
    .A(\proj__3.net13 ));
 sg13g2_or2_1 \proj__3.or4/_0_  (.X(\proj__3.net13 ),
    .B(\proj__3.net4 ),
    .A(\proj__3.net3 ));
 sg13g2_inv_1 \proj__4.flop1/_4_  (.Y(\proj__4.flop1/_1_ ),
    .A(\proj__4.flop1/s ));
 sg13g2_inv_1 \proj__4.flop1/_5_  (.Y(\proj__4.flop1/_0_ ),
    .A(net110));
 sg13g2_tielo \proj__4.flop1/dffsr_210  (.L_LO(net219));
 sg13g2_tielo \proj__4.flop2/dffsr_211  (.L_LO(net220));
 sg13g2_sdfbbp_1 \proj__4.flop1/dffsr  (.Q(\proj__4.flop1/q ),
    .Q_N(\proj__4.net11 ),
    .RESET_B(\proj__4.flop1/_0_ ),
    .SET_B(\proj__4.flop1/_1_ ),
    .D(net41),
    .SCE(net219),
    .SCD(net218),
    .CLK(net109));
 sg13g2_inv_1 \proj__4.flop2/_4_  (.Y(\proj__4.flop2/_1_ ),
    .A(\proj__4.flop2/s ));
 sg13g2_inv_1 \proj__4.flop2/_5_  (.Y(\proj__4.flop2/_0_ ),
    .A(net112));
 sg13g2_tielo \proj__4.flop2/dffsr_212  (.L_LO(net221));
 sg13g2_tielo \proj__4.flop3/dffsr_213  (.L_LO(net222));
 sg13g2_sdfbbp_1 \proj__4.flop2/dffsr  (.Q(\proj__4.flop2/q ),
    .Q_N(\proj__4.net12 ),
    .RESET_B(\proj__4.flop2/_0_ ),
    .SET_B(\proj__4.flop2/_1_ ),
    .D(net39),
    .SCE(net221),
    .SCD(net220),
    .CLK(net111));
 sg13g2_inv_1 \proj__4.flop3/_4_  (.Y(\proj__4.flop3/_1_ ),
    .A(\proj__4.flop3/s ));
 sg13g2_inv_1 \proj__4.flop3/_5_  (.Y(\proj__4.flop3/_0_ ),
    .A(net114));
 sg13g2_tielo \proj__4.flop3/dffsr_214  (.L_LO(net223));
 sg13g2_tielo \proj__4.flop4/dffsr_215  (.L_LO(net224));
 sg13g2_sdfbbp_1 \proj__4.flop3/dffsr  (.Q(\proj__4.flop3/q ),
    .Q_N(\proj__4.net13 ),
    .RESET_B(\proj__4.flop3/_0_ ),
    .SET_B(\proj__4.flop3/_1_ ),
    .D(net2),
    .SCE(net223),
    .SCD(net222),
    .CLK(net113));
 sg13g2_inv_1 \proj__4.flop4/_4_  (.Y(\proj__4.flop4/_1_ ),
    .A(\proj__4.flop4/s ));
 sg13g2_inv_1 \proj__4.flop4/_5_  (.Y(\proj__4.flop4/_0_ ),
    .A(net116));
 sg13g2_tielo \proj__4.flop4/dffsr_216  (.L_LO(net225));
 sg13g2_tielo \proj__4.flop5/dffsr_217  (.L_LO(net226));
 sg13g2_sdfbbp_1 \proj__4.flop4/dffsr  (.Q(\proj__4.flop4/q ),
    .Q_N(\proj__4.net14 ),
    .RESET_B(\proj__4.flop4/_0_ ),
    .SET_B(\proj__4.flop4/_1_ ),
    .D(net36),
    .SCE(net225),
    .SCD(net224),
    .CLK(net115));
 sg13g2_inv_1 \proj__4.flop5/_4_  (.Y(\proj__4.flop5/_1_ ),
    .A(\proj__4.flop5/s ));
 sg13g2_inv_1 \proj__4.flop5/_5_  (.Y(\proj__4.flop5/_0_ ),
    .A(net118));
 sg13g2_tielo \proj__4.flop5/dffsr_218  (.L_LO(net227));
 sg13g2_tielo \proj__4.flop6/dffsr_219  (.L_LO(net228));
 sg13g2_sdfbbp_1 \proj__4.flop5/dffsr  (.Q(\proj__4.net15 ),
    .Q_N(\proj__4.flop5/notq ),
    .RESET_B(\proj__4.flop5/_0_ ),
    .SET_B(\proj__4.flop5/_1_ ),
    .D(net4),
    .SCE(net227),
    .SCD(net226),
    .CLK(net117));
 sg13g2_inv_1 \proj__4.flop6/_4_  (.Y(\proj__4.flop6/_1_ ),
    .A(\proj__4.flop6/s ));
 sg13g2_inv_1 \proj__4.flop6/_5_  (.Y(\proj__4.flop6/_0_ ),
    .A(net120));
 sg13g2_tielo \proj__4.flop6/dffsr_220  (.L_LO(net229));
 sg13g2_tielo \proj__4.flop8/dffsr_221  (.L_LO(net230));
 sg13g2_sdfbbp_1 \proj__4.flop6/dffsr  (.Q(\proj__4.net16 ),
    .Q_N(\proj__4.flop6/notq ),
    .RESET_B(\proj__4.flop6/_0_ ),
    .SET_B(\proj__4.flop6/_1_ ),
    .D(net35),
    .SCE(net229),
    .SCD(net228),
    .CLK(net119));
 sg13g2_inv_1 \proj__4.flop8/_4_  (.Y(\proj__4.flop8/_1_ ),
    .A(\proj__4.flop8/s ));
 sg13g2_inv_1 \proj__4.flop8/_5_  (.Y(\proj__4.flop8/_0_ ),
    .A(net122));
 sg13g2_tielo \proj__4.flop8/dffsr_222  (.L_LO(net231));
 sg13g2_tielo \proj__4.flop9/dffsr_223  (.L_LO(net232));
 sg13g2_sdfbbp_1 \proj__4.flop8/dffsr  (.Q(\proj__4.net17 ),
    .Q_N(\proj__4.flop8/notq ),
    .RESET_B(\proj__4.flop8/_0_ ),
    .SET_B(\proj__4.flop8/_1_ ),
    .D(net6),
    .SCE(net231),
    .SCD(net230),
    .CLK(net121));
 sg13g2_inv_1 \proj__4.flop9/_4_  (.Y(\proj__4.flop9/_1_ ),
    .A(\proj__4.flop9/s ));
 sg13g2_inv_1 \proj__4.flop9/_5_  (.Y(\proj__4.flop9/_0_ ),
    .A(net124));
 sg13g2_tielo \proj__4.flop9/dffsr_224  (.L_LO(net233));
 sg13g2_tielo \proj__9.flop1/dffsr_225  (.L_LO(net234));
 sg13g2_sdfbbp_1 \proj__4.flop9/dffsr  (.Q(\proj__4.net18 ),
    .Q_N(\proj__4.flop9/notq ),
    .RESET_B(\proj__4.flop9/_0_ ),
    .SET_B(\proj__4.flop9/_1_ ),
    .D(net7),
    .SCE(net233),
    .SCD(net232),
    .CLK(net123));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net39),
    .B(net41),
    .X(\proj__5.net9 ));
 sg13g2_and2_1 \proj__5.and2/_0_  (.A(net36),
    .B(net37),
    .X(\proj__5.net12 ));
 sg13g2_inv_1 \proj__5.not1/_0_  (.Y(\proj__5.net10 ),
    .A(net6));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net11 ),
    .B(net4),
    .A(net35));
 sg13g2_inv_1 \proj__6.not3/_0_  (.Y(\proj__6.net9 ),
    .A(net37));
 sg13g2_inv_1 \proj__6.not4/_0_  (.Y(\proj__6.net10 ),
    .A(net36));
 sg13g2_dfrbp_1 \proj__7.flop1/_1_  (.CLK(net125),
    .RESET_B(net252),
    .D(net7),
    .Q_N(\proj__7.net6 ),
    .Q(\proj__7.net5 ));
 sg13g2_tiehi \proj__7.flop2/_1__244  (.L_HI(net253));
 sg13g2_dfrbp_1 \proj__7.flop2/_1_  (.CLK(net126),
    .RESET_B(net253),
    .D(\proj__7.net14 ),
    .Q_N(\proj__7.net14 ),
    .Q(\proj__7.net8 ));
 sg13g2_tiehi \proj__7.flop3/_1__245  (.L_HI(net254));
 sg13g2_dfrbp_1 \proj__7.flop3/_1_  (.CLK(\proj__7.net14 ),
    .RESET_B(net254),
    .D(\proj__7.net15 ),
    .Q_N(\proj__7.net15 ),
    .Q(\proj__7.net7 ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_and2_1 \proj__8.and1/_0_  (.A(net38),
    .B(net40),
    .X(\proj__8.net7 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(\proj__9.net11 ),
    .B(net1),
    .X(\proj__9.net12 ));
 sg13g2_and2_1 \proj__9.and2/_0_  (.A(net39),
    .B(\proj__9.net13 ),
    .X(\proj__9.net14 ));
 sg13g2_inv_1 \proj__9.flop1/_4_  (.Y(\proj__9.flop1/_1_ ),
    .A(net128));
 sg13g2_inv_1 \proj__9.flop1/_5_  (.Y(\proj__9.flop1/_0_ ),
    .A(\proj__9.net17 ));
 sg13g2_tielo \proj__9.flop1/dffsr_226  (.L_LO(net235));
 sg13g2_tiehi \proj_14.mux10/_0__227  (.L_HI(net236));
 sg13g2_sdfbbp_1 \proj__9.flop1/dffsr  (.Q(\proj__9.net5 ),
    .Q_N(\proj__9.flop1/notq ),
    .RESET_B(\proj__9.flop1/_0_ ),
    .SET_B(\proj__9.flop1/_1_ ),
    .D(\proj__9.net15 ),
    .SCE(net235),
    .SCD(net234),
    .CLK(net127));
 sg13g2_inv_1 \proj__9.not1/_0_  (.Y(\proj__9.net11 ),
    .A(net39));
 sg13g2_inv_1 \proj__9.not2/_0_  (.Y(\proj__9.net13 ),
    .A(net41));
 sg13g2_inv_1 \proj__9.not3/_0_  (.Y(\proj__9.net17 ),
    .A(net129));
 sg13g2_or2_1 \proj__9.or1/_0_  (.X(\proj__9.net15 ),
    .B(\proj__9.net12 ),
    .A(\proj__9.net14 ));
 sg13g2_buf_4 fanout35 (.X(net35),
    .A(net5));
 sg13g2_buf_2 fanout36 (.A(net3),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(net2),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(net39),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(ui_in[1]),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(net41),
    .X(net40));
 sg13g2_buf_4 fanout41 (.X(net41),
    .A(net1));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(net43));
 sg13g2_buf_4 fanout43 (.X(net43),
    .A(\proj_14.net45 ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[4]));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_4 input6 (.X(net6),
    .A(ui_in[6]));
 sg13g2_buf_2 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_tielo \proj_13.flop1/_1__12  (.L_LO(net12));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_4 FILLER_14_336 ();
 sg13g2_fill_2 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_4 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_4 FILLER_16_294 ();
 sg13g2_fill_2 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_303 ();
 sg13g2_fill_2 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_4 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_fill_2 FILLER_16_340 ();
 sg13g2_fill_1 FILLER_16_342 ();
 sg13g2_decap_4 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_32 ();
 sg13g2_decap_8 FILLER_17_39 ();
 sg13g2_decap_8 FILLER_17_46 ();
 sg13g2_decap_8 FILLER_17_53 ();
 sg13g2_decap_8 FILLER_17_60 ();
 sg13g2_fill_2 FILLER_17_67 ();
 sg13g2_decap_4 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_76 ();
 sg13g2_decap_8 FILLER_17_81 ();
 sg13g2_decap_8 FILLER_17_88 ();
 sg13g2_decap_8 FILLER_17_95 ();
 sg13g2_decap_8 FILLER_17_102 ();
 sg13g2_decap_8 FILLER_17_109 ();
 sg13g2_decap_8 FILLER_17_116 ();
 sg13g2_decap_8 FILLER_17_123 ();
 sg13g2_decap_8 FILLER_17_130 ();
 sg13g2_decap_8 FILLER_17_137 ();
 sg13g2_decap_8 FILLER_17_144 ();
 sg13g2_decap_8 FILLER_17_151 ();
 sg13g2_decap_8 FILLER_17_158 ();
 sg13g2_decap_8 FILLER_17_165 ();
 sg13g2_decap_8 FILLER_17_172 ();
 sg13g2_decap_8 FILLER_17_179 ();
 sg13g2_decap_8 FILLER_17_186 ();
 sg13g2_decap_8 FILLER_17_193 ();
 sg13g2_decap_8 FILLER_17_200 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_221 ();
 sg13g2_decap_8 FILLER_17_228 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_decap_8 FILLER_17_242 ();
 sg13g2_decap_8 FILLER_17_249 ();
 sg13g2_decap_8 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_263 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_fill_1 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_339 ();
 sg13g2_fill_2 FILLER_17_344 ();
 sg13g2_decap_4 FILLER_17_350 ();
 sg13g2_decap_4 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_9 ();
 sg13g2_fill_2 FILLER_18_48 ();
 sg13g2_fill_1 FILLER_18_50 ();
 sg13g2_decap_4 FILLER_18_90 ();
 sg13g2_fill_2 FILLER_18_98 ();
 sg13g2_fill_1 FILLER_18_100 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_decap_8 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_186 ();
 sg13g2_decap_8 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_fill_2 FILLER_18_284 ();
 sg13g2_fill_2 FILLER_18_298 ();
 sg13g2_fill_1 FILLER_18_300 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_312 ();
 sg13g2_fill_1 FILLER_18_314 ();
 sg13g2_decap_4 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_323 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_1 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_17 ();
 sg13g2_decap_8 FILLER_19_23 ();
 sg13g2_decap_8 FILLER_19_34 ();
 sg13g2_fill_2 FILLER_19_41 ();
 sg13g2_fill_1 FILLER_19_43 ();
 sg13g2_fill_1 FILLER_19_58 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_fill_2 FILLER_19_74 ();
 sg13g2_fill_1 FILLER_19_76 ();
 sg13g2_fill_2 FILLER_19_87 ();
 sg13g2_decap_8 FILLER_19_131 ();
 sg13g2_fill_2 FILLER_19_138 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_148 ();
 sg13g2_decap_8 FILLER_19_155 ();
 sg13g2_decap_8 FILLER_19_162 ();
 sg13g2_decap_8 FILLER_19_169 ();
 sg13g2_decap_8 FILLER_19_176 ();
 sg13g2_decap_8 FILLER_19_183 ();
 sg13g2_decap_8 FILLER_19_190 ();
 sg13g2_decap_4 FILLER_19_197 ();
 sg13g2_decap_8 FILLER_19_204 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_225 ();
 sg13g2_decap_8 FILLER_19_232 ();
 sg13g2_decap_8 FILLER_19_239 ();
 sg13g2_decap_8 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_253 ();
 sg13g2_decap_8 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_267 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_352 ();
 sg13g2_decap_4 FILLER_19_358 ();
 sg13g2_fill_2 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_11 ();
 sg13g2_fill_1 FILLER_20_13 ();
 sg13g2_decap_4 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_26 ();
 sg13g2_fill_2 FILLER_20_36 ();
 sg13g2_fill_1 FILLER_20_38 ();
 sg13g2_decap_4 FILLER_20_49 ();
 sg13g2_fill_1 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_62 ();
 sg13g2_fill_2 FILLER_20_69 ();
 sg13g2_fill_2 FILLER_20_81 ();
 sg13g2_decap_4 FILLER_20_87 ();
 sg13g2_fill_2 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_96 ();
 sg13g2_decap_4 FILLER_20_106 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_114 ();
 sg13g2_decap_8 FILLER_20_121 ();
 sg13g2_fill_2 FILLER_20_132 ();
 sg13g2_decap_8 FILLER_20_138 ();
 sg13g2_decap_8 FILLER_20_145 ();
 sg13g2_decap_8 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_decap_8 FILLER_20_173 ();
 sg13g2_decap_4 FILLER_20_180 ();
 sg13g2_decap_4 FILLER_20_222 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_4 FILLER_20_294 ();
 sg13g2_decap_4 FILLER_20_310 ();
 sg13g2_fill_1 FILLER_20_314 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_fill_2 FILLER_20_336 ();
 sg13g2_decap_4 FILLER_20_385 ();
 sg13g2_fill_2 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_114 ();
 sg13g2_fill_2 FILLER_21_121 ();
 sg13g2_decap_8 FILLER_21_149 ();
 sg13g2_decap_8 FILLER_21_156 ();
 sg13g2_decap_8 FILLER_21_163 ();
 sg13g2_fill_1 FILLER_21_170 ();
 sg13g2_decap_8 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_fill_2 FILLER_21_191 ();
 sg13g2_decap_4 FILLER_21_197 ();
 sg13g2_fill_1 FILLER_21_201 ();
 sg13g2_decap_8 FILLER_21_206 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_decap_8 FILLER_21_220 ();
 sg13g2_decap_8 FILLER_21_234 ();
 sg13g2_decap_8 FILLER_21_241 ();
 sg13g2_fill_2 FILLER_21_248 ();
 sg13g2_decap_8 FILLER_21_253 ();
 sg13g2_decap_8 FILLER_21_260 ();
 sg13g2_decap_8 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_fill_1 FILLER_21_364 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_4 ();
 sg13g2_decap_4 FILLER_22_10 ();
 sg13g2_fill_2 FILLER_22_18 ();
 sg13g2_decap_4 FILLER_22_27 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_decap_8 FILLER_22_36 ();
 sg13g2_decap_8 FILLER_22_43 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_decap_4 FILLER_22_61 ();
 sg13g2_decap_8 FILLER_22_69 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_111 ();
 sg13g2_decap_8 FILLER_22_117 ();
 sg13g2_fill_2 FILLER_22_128 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_4 FILLER_22_188 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_197 ();
 sg13g2_fill_1 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_22_204 ();
 sg13g2_fill_1 FILLER_22_211 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_decap_4 FILLER_22_229 ();
 sg13g2_fill_2 FILLER_22_233 ();
 sg13g2_fill_2 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_decap_4 FILLER_22_288 ();
 sg13g2_fill_1 FILLER_22_299 ();
 sg13g2_fill_1 FILLER_22_310 ();
 sg13g2_decap_4 FILLER_22_316 ();
 sg13g2_decap_4 FILLER_22_332 ();
 sg13g2_fill_2 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_352 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_decap_4 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_fill_2 FILLER_22_390 ();
 sg13g2_fill_1 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_50 ();
 sg13g2_decap_8 FILLER_23_139 ();
 sg13g2_fill_2 FILLER_23_146 ();
 sg13g2_fill_1 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_157 ();
 sg13g2_decap_4 FILLER_23_163 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_176 ();
 sg13g2_decap_4 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_fill_2 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_250 ();
 sg13g2_decap_8 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_262 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_4 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_fill_1 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_4 FILLER_23_312 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_321 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_decap_4 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_332 ();
 sg13g2_decap_4 FILLER_23_337 ();
 sg13g2_fill_2 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_decap_8 FILLER_23_355 ();
 sg13g2_decap_4 FILLER_23_362 ();
 sg13g2_fill_2 FILLER_23_366 ();
 sg13g2_fill_2 FILLER_23_372 ();
 sg13g2_decap_4 FILLER_23_378 ();
 sg13g2_decap_4 FILLER_23_386 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_9 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_16 ();
 sg13g2_decap_4 FILLER_24_24 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_32 ();
 sg13g2_fill_2 FILLER_24_39 ();
 sg13g2_decap_4 FILLER_24_51 ();
 sg13g2_fill_2 FILLER_24_55 ();
 sg13g2_decap_8 FILLER_24_61 ();
 sg13g2_decap_4 FILLER_24_68 ();
 sg13g2_fill_2 FILLER_24_72 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_decap_4 FILLER_24_92 ();
 sg13g2_fill_1 FILLER_24_96 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_fill_2 FILLER_24_110 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_decap_4 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_148 ();
 sg13g2_decap_4 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_195 ();
 sg13g2_fill_2 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_decap_4 FILLER_24_207 ();
 sg13g2_fill_2 FILLER_24_211 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_2 FILLER_24_240 ();
 sg13g2_decap_4 FILLER_24_246 ();
 sg13g2_decap_4 FILLER_24_254 ();
 sg13g2_fill_2 FILLER_24_258 ();
 sg13g2_fill_2 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_298 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_decap_4 FILLER_25_47 ();
 sg13g2_fill_2 FILLER_25_51 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_138 ();
 sg13g2_fill_2 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_152 ();
 sg13g2_fill_2 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_188 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_312 ();
 sg13g2_fill_1 FILLER_25_314 ();
 sg13g2_fill_2 FILLER_25_322 ();
 sg13g2_fill_1 FILLER_25_324 ();
 sg13g2_decap_4 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_fill_1 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_decap_4 FILLER_25_356 ();
 sg13g2_fill_2 FILLER_25_360 ();
 sg13g2_fill_2 FILLER_25_366 ();
 sg13g2_fill_2 FILLER_25_372 ();
 sg13g2_fill_1 FILLER_25_374 ();
 sg13g2_fill_2 FILLER_25_378 ();
 sg13g2_fill_1 FILLER_25_380 ();
 sg13g2_fill_2 FILLER_25_384 ();
 sg13g2_fill_2 FILLER_25_389 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_fill_2 FILLER_26_28 ();
 sg13g2_decap_4 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_60 ();
 sg13g2_fill_2 FILLER_26_69 ();
 sg13g2_fill_2 FILLER_26_75 ();
 sg13g2_fill_2 FILLER_26_80 ();
 sg13g2_decap_8 FILLER_26_86 ();
 sg13g2_fill_2 FILLER_26_93 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_110 ();
 sg13g2_fill_1 FILLER_26_117 ();
 sg13g2_decap_4 FILLER_26_131 ();
 sg13g2_fill_2 FILLER_26_135 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_157 ();
 sg13g2_fill_1 FILLER_26_159 ();
 sg13g2_fill_1 FILLER_26_165 ();
 sg13g2_decap_4 FILLER_26_171 ();
 sg13g2_fill_2 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_4 FILLER_26_196 ();
 sg13g2_fill_2 FILLER_26_204 ();
 sg13g2_fill_1 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_215 ();
 sg13g2_decap_4 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_223 ();
 sg13g2_decap_8 FILLER_26_229 ();
 sg13g2_fill_1 FILLER_26_236 ();
 sg13g2_fill_2 FILLER_26_241 ();
 sg13g2_fill_1 FILLER_26_243 ();
 sg13g2_fill_1 FILLER_26_248 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_263 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_decap_8 FILLER_26_274 ();
 sg13g2_decap_8 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_30 ();
 sg13g2_fill_2 FILLER_27_39 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_108 ();
 sg13g2_decap_4 FILLER_27_115 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_180 ();
 sg13g2_decap_4 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_decap_4 FILLER_27_274 ();
 sg13g2_fill_2 FILLER_27_278 ();
 sg13g2_decap_4 FILLER_27_295 ();
 sg13g2_decap_4 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_315 ();
 sg13g2_fill_2 FILLER_27_321 ();
 sg13g2_decap_4 FILLER_27_327 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_decap_4 FILLER_27_335 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_4 FILLER_27_370 ();
 sg13g2_fill_2 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_25 ();
 sg13g2_fill_1 FILLER_28_62 ();
 sg13g2_fill_2 FILLER_28_67 ();
 sg13g2_decap_4 FILLER_28_73 ();
 sg13g2_fill_1 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_82 ();
 sg13g2_decap_8 FILLER_28_89 ();
 sg13g2_fill_1 FILLER_28_96 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_127 ();
 sg13g2_decap_4 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_decap_4 FILLER_28_142 ();
 sg13g2_decap_8 FILLER_28_149 ();
 sg13g2_decap_4 FILLER_28_156 ();
 sg13g2_fill_2 FILLER_28_160 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_fill_1 FILLER_28_201 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_212 ();
 sg13g2_decap_4 FILLER_28_219 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_decap_8 FILLER_28_227 ();
 sg13g2_decap_4 FILLER_28_234 ();
 sg13g2_decap_4 FILLER_28_245 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_decap_4 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_257 ();
 sg13g2_decap_4 FILLER_28_284 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_309 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_decap_8 FILLER_29_65 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_decap_8 FILLER_29_88 ();
 sg13g2_decap_4 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_164 ();
 sg13g2_fill_1 FILLER_29_166 ();
 sg13g2_fill_1 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_fill_2 FILLER_29_195 ();
 sg13g2_fill_1 FILLER_29_223 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_fill_2 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_283 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_decap_4 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_344 ();
 sg13g2_decap_8 FILLER_29_361 ();
 sg13g2_decap_4 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_384 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_31 ();
 sg13g2_decap_4 FILLER_30_37 ();
 sg13g2_fill_2 FILLER_30_48 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_fill_2 FILLER_30_54 ();
 sg13g2_fill_1 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_67 ();
 sg13g2_decap_4 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_107 ();
 sg13g2_decap_8 FILLER_30_118 ();
 sg13g2_fill_2 FILLER_30_125 ();
 sg13g2_fill_1 FILLER_30_127 ();
 sg13g2_fill_2 FILLER_30_136 ();
 sg13g2_decap_4 FILLER_30_142 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_decap_8 FILLER_30_151 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_decap_4 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_180 ();
 sg13g2_decap_8 FILLER_30_187 ();
 sg13g2_decap_4 FILLER_30_194 ();
 sg13g2_fill_2 FILLER_30_198 ();
 sg13g2_fill_2 FILLER_30_204 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_fill_1 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_fill_1 FILLER_30_250 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_fill_2 FILLER_30_281 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_decap_8 FILLER_30_307 ();
 sg13g2_fill_2 FILLER_30_314 ();
 sg13g2_fill_1 FILLER_30_316 ();
 sg13g2_fill_2 FILLER_30_330 ();
 sg13g2_fill_1 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_fill_1 FILLER_30_347 ();
 sg13g2_decap_4 FILLER_30_361 ();
 sg13g2_decap_4 FILLER_30_369 ();
 sg13g2_fill_2 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_4 FILLER_30_385 ();
 sg13g2_fill_1 FILLER_30_389 ();
 sg13g2_decap_4 FILLER_30_393 ();
 sg13g2_fill_1 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_11 ();
 sg13g2_fill_2 FILLER_31_16 ();
 sg13g2_decap_4 FILLER_31_22 ();
 sg13g2_fill_1 FILLER_31_26 ();
 sg13g2_decap_8 FILLER_31_37 ();
 sg13g2_decap_8 FILLER_31_44 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_decap_4 FILLER_31_62 ();
 sg13g2_fill_2 FILLER_31_71 ();
 sg13g2_decap_4 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_92 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_4 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_130 ();
 sg13g2_fill_2 FILLER_31_135 ();
 sg13g2_decap_8 FILLER_31_141 ();
 sg13g2_fill_2 FILLER_31_148 ();
 sg13g2_decap_8 FILLER_31_162 ();
 sg13g2_decap_8 FILLER_31_221 ();
 sg13g2_decap_4 FILLER_31_228 ();
 sg13g2_decap_4 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_248 ();
 sg13g2_decap_4 FILLER_31_255 ();
 sg13g2_fill_2 FILLER_31_259 ();
 sg13g2_fill_2 FILLER_31_270 ();
 sg13g2_fill_1 FILLER_31_277 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_335 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_2 FILLER_31_396 ();
 sg13g2_fill_1 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_33 ();
 sg13g2_fill_2 FILLER_32_37 ();
 sg13g2_fill_1 FILLER_32_64 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_117 ();
 sg13g2_decap_4 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_173 ();
 sg13g2_decap_8 FILLER_32_187 ();
 sg13g2_decap_4 FILLER_32_194 ();
 sg13g2_fill_1 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_275 ();
 sg13g2_fill_2 FILLER_32_282 ();
 sg13g2_decap_8 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_299 ();
 sg13g2_fill_2 FILLER_32_303 ();
 sg13g2_fill_1 FILLER_32_305 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_fill_1 FILLER_32_348 ();
 sg13g2_decap_4 FILLER_32_354 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_363 ();
 sg13g2_decap_4 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_95 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_decap_8 FILLER_33_121 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_decap_8 FILLER_33_134 ();
 sg13g2_decap_8 FILLER_33_141 ();
 sg13g2_fill_1 FILLER_33_148 ();
 sg13g2_decap_8 FILLER_33_152 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_4 FILLER_33_196 ();
 sg13g2_fill_2 FILLER_33_208 ();
 sg13g2_decap_4 FILLER_33_214 ();
 sg13g2_fill_1 FILLER_33_218 ();
 sg13g2_decap_4 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_232 ();
 sg13g2_decap_4 FILLER_33_243 ();
 sg13g2_fill_2 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_decap_4 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_decap_4 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_333 ();
 sg13g2_fill_2 FILLER_33_372 ();
 sg13g2_fill_1 FILLER_33_374 ();
 sg13g2_decap_4 FILLER_33_387 ();
 sg13g2_fill_2 FILLER_33_391 ();
 sg13g2_fill_2 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_4 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_58 ();
 sg13g2_fill_1 FILLER_34_62 ();
 sg13g2_decap_8 FILLER_34_68 ();
 sg13g2_decap_4 FILLER_34_75 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_4 FILLER_34_91 ();
 sg13g2_fill_1 FILLER_34_95 ();
 sg13g2_fill_2 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_108 ();
 sg13g2_fill_2 FILLER_34_113 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_fill_2 FILLER_34_168 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_decap_4 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_314 ();
 sg13g2_decap_4 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_325 ();
 sg13g2_decap_4 FILLER_34_331 ();
 sg13g2_fill_2 FILLER_34_346 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_decap_8 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_4 FILLER_34_389 ();
 sg13g2_fill_2 FILLER_34_393 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_4 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_102 ();
 sg13g2_decap_8 FILLER_35_130 ();
 sg13g2_decap_8 FILLER_35_137 ();
 sg13g2_decap_8 FILLER_35_144 ();
 sg13g2_decap_8 FILLER_35_151 ();
 sg13g2_decap_8 FILLER_35_158 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_decap_8 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_183 ();
 sg13g2_decap_8 FILLER_35_190 ();
 sg13g2_decap_8 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_decap_4 FILLER_35_221 ();
 sg13g2_fill_2 FILLER_35_225 ();
 sg13g2_decap_8 FILLER_35_230 ();
 sg13g2_decap_8 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_decap_8 FILLER_35_278 ();
 sg13g2_decap_8 FILLER_35_285 ();
 sg13g2_decap_4 FILLER_35_292 ();
 sg13g2_fill_1 FILLER_35_310 ();
 sg13g2_decap_4 FILLER_35_317 ();
 sg13g2_fill_2 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_4 FILLER_35_364 ();
 sg13g2_fill_1 FILLER_35_368 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_4 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_200 ();
 sg13g2_fill_2 FILLER_36_268 ();
 sg13g2_decap_8 FILLER_36_283 ();
 sg13g2_fill_2 FILLER_36_290 ();
 sg13g2_fill_2 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_decap_4 FILLER_36_349 ();
 sg13g2_fill_2 FILLER_36_353 ();
 sg13g2_fill_2 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_365 ();
 sg13g2_fill_2 FILLER_36_372 ();
 sg13g2_fill_1 FILLER_36_374 ();
 sg13g2_fill_2 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_4 FILLER_37_203 ();
 sg13g2_fill_2 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_fill_1 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_236 ();
 sg13g2_decap_8 FILLER_37_243 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_fill_2 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_250 ();
 sg13g2_decap_4 FILLER_38_263 ();
 sg13g2_fill_1 FILLER_38_267 ();
 sg13g2_decap_4 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net130;
 assign uio_oe[1] = net131;
 assign uio_oe[2] = net132;
 assign uio_oe[3] = net133;
 assign uio_oe[4] = net134;
 assign uio_oe[5] = net135;
 assign uio_oe[6] = net136;
 assign uio_oe[7] = net137;
 assign uio_out[0] = net138;
 assign uio_out[1] = net139;
 assign uio_out[2] = net140;
 assign uio_out[3] = net141;
 assign uio_out[4] = net142;
 assign uio_out[5] = net143;
 assign uio_out[6] = net144;
 assign uio_out[7] = net145;
endmodule

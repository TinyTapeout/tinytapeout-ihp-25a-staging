module tt_um_rtfb_collatz (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire clknet_0_clk;
 wire \collatz.busy ;
 wire \collatz.comp ;
 wire \collatz.iter[0] ;
 wire \collatz.iter[100] ;
 wire \collatz.iter[101] ;
 wire \collatz.iter[102] ;
 wire \collatz.iter[103] ;
 wire \collatz.iter[104] ;
 wire \collatz.iter[105] ;
 wire \collatz.iter[106] ;
 wire \collatz.iter[107] ;
 wire \collatz.iter[108] ;
 wire \collatz.iter[109] ;
 wire \collatz.iter[10] ;
 wire \collatz.iter[110] ;
 wire \collatz.iter[111] ;
 wire \collatz.iter[112] ;
 wire \collatz.iter[113] ;
 wire \collatz.iter[114] ;
 wire \collatz.iter[115] ;
 wire \collatz.iter[116] ;
 wire \collatz.iter[117] ;
 wire \collatz.iter[118] ;
 wire \collatz.iter[119] ;
 wire \collatz.iter[11] ;
 wire \collatz.iter[120] ;
 wire \collatz.iter[121] ;
 wire \collatz.iter[122] ;
 wire \collatz.iter[123] ;
 wire \collatz.iter[124] ;
 wire \collatz.iter[125] ;
 wire \collatz.iter[126] ;
 wire \collatz.iter[127] ;
 wire \collatz.iter[128] ;
 wire \collatz.iter[129] ;
 wire \collatz.iter[12] ;
 wire \collatz.iter[130] ;
 wire \collatz.iter[131] ;
 wire \collatz.iter[132] ;
 wire \collatz.iter[133] ;
 wire \collatz.iter[134] ;
 wire \collatz.iter[135] ;
 wire \collatz.iter[136] ;
 wire \collatz.iter[137] ;
 wire \collatz.iter[138] ;
 wire \collatz.iter[139] ;
 wire \collatz.iter[13] ;
 wire \collatz.iter[140] ;
 wire \collatz.iter[141] ;
 wire \collatz.iter[142] ;
 wire \collatz.iter[143] ;
 wire \collatz.iter[14] ;
 wire \collatz.iter[15] ;
 wire \collatz.iter[16] ;
 wire \collatz.iter[17] ;
 wire \collatz.iter[18] ;
 wire \collatz.iter[19] ;
 wire \collatz.iter[1] ;
 wire \collatz.iter[20] ;
 wire \collatz.iter[21] ;
 wire \collatz.iter[22] ;
 wire \collatz.iter[23] ;
 wire \collatz.iter[24] ;
 wire \collatz.iter[25] ;
 wire \collatz.iter[26] ;
 wire \collatz.iter[27] ;
 wire \collatz.iter[28] ;
 wire \collatz.iter[29] ;
 wire \collatz.iter[2] ;
 wire \collatz.iter[30] ;
 wire \collatz.iter[31] ;
 wire \collatz.iter[32] ;
 wire \collatz.iter[33] ;
 wire \collatz.iter[34] ;
 wire \collatz.iter[35] ;
 wire \collatz.iter[36] ;
 wire \collatz.iter[37] ;
 wire \collatz.iter[38] ;
 wire \collatz.iter[39] ;
 wire \collatz.iter[3] ;
 wire \collatz.iter[40] ;
 wire \collatz.iter[41] ;
 wire \collatz.iter[42] ;
 wire \collatz.iter[43] ;
 wire \collatz.iter[44] ;
 wire \collatz.iter[45] ;
 wire \collatz.iter[46] ;
 wire \collatz.iter[47] ;
 wire \collatz.iter[48] ;
 wire \collatz.iter[49] ;
 wire \collatz.iter[4] ;
 wire \collatz.iter[50] ;
 wire \collatz.iter[51] ;
 wire \collatz.iter[52] ;
 wire \collatz.iter[53] ;
 wire \collatz.iter[54] ;
 wire \collatz.iter[55] ;
 wire \collatz.iter[56] ;
 wire \collatz.iter[57] ;
 wire \collatz.iter[58] ;
 wire \collatz.iter[59] ;
 wire \collatz.iter[5] ;
 wire \collatz.iter[60] ;
 wire \collatz.iter[61] ;
 wire \collatz.iter[62] ;
 wire \collatz.iter[63] ;
 wire \collatz.iter[64] ;
 wire \collatz.iter[65] ;
 wire \collatz.iter[66] ;
 wire \collatz.iter[67] ;
 wire \collatz.iter[68] ;
 wire \collatz.iter[69] ;
 wire \collatz.iter[6] ;
 wire \collatz.iter[70] ;
 wire \collatz.iter[71] ;
 wire \collatz.iter[72] ;
 wire \collatz.iter[73] ;
 wire \collatz.iter[74] ;
 wire \collatz.iter[75] ;
 wire \collatz.iter[76] ;
 wire \collatz.iter[77] ;
 wire \collatz.iter[78] ;
 wire \collatz.iter[79] ;
 wire \collatz.iter[7] ;
 wire \collatz.iter[80] ;
 wire \collatz.iter[81] ;
 wire \collatz.iter[82] ;
 wire \collatz.iter[83] ;
 wire \collatz.iter[84] ;
 wire \collatz.iter[85] ;
 wire \collatz.iter[86] ;
 wire \collatz.iter[87] ;
 wire \collatz.iter[88] ;
 wire \collatz.iter[89] ;
 wire \collatz.iter[8] ;
 wire \collatz.iter[90] ;
 wire \collatz.iter[91] ;
 wire \collatz.iter[92] ;
 wire \collatz.iter[93] ;
 wire \collatz.iter[94] ;
 wire \collatz.iter[95] ;
 wire \collatz.iter[96] ;
 wire \collatz.iter[97] ;
 wire \collatz.iter[98] ;
 wire \collatz.iter[99] ;
 wire \collatz.iter[9] ;
 wire \collatz.orbit_len[0] ;
 wire \collatz.orbit_len[10] ;
 wire \collatz.orbit_len[11] ;
 wire \collatz.orbit_len[12] ;
 wire \collatz.orbit_len[13] ;
 wire \collatz.orbit_len[14] ;
 wire \collatz.orbit_len[15] ;
 wire \collatz.orbit_len[1] ;
 wire \collatz.orbit_len[2] ;
 wire \collatz.orbit_len[3] ;
 wire \collatz.orbit_len[4] ;
 wire \collatz.orbit_len[5] ;
 wire \collatz.orbit_len[6] ;
 wire \collatz.orbit_len[7] ;
 wire \collatz.orbit_len[8] ;
 wire \collatz.orbit_len[9] ;
 wire \collatz.path_record_h16[0] ;
 wire \collatz.path_record_h16[10] ;
 wire \collatz.path_record_h16[11] ;
 wire \collatz.path_record_h16[12] ;
 wire \collatz.path_record_h16[13] ;
 wire \collatz.path_record_h16[14] ;
 wire \collatz.path_record_h16[15] ;
 wire \collatz.path_record_h16[1] ;
 wire \collatz.path_record_h16[2] ;
 wire \collatz.path_record_h16[3] ;
 wire \collatz.path_record_h16[4] ;
 wire \collatz.path_record_h16[5] ;
 wire \collatz.path_record_h16[6] ;
 wire \collatz.path_record_h16[7] ;
 wire \collatz.path_record_h16[8] ;
 wire \collatz.path_record_h16[9] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;

 sg13g2_inv_1 _2328_ (.Y(_1375_),
    .A(net213));
 sg13g2_inv_1 _2329_ (.Y(_1376_),
    .A(net234));
 sg13g2_inv_1 _2330_ (.Y(_1377_),
    .A(net248));
 sg13g2_inv_1 _2331_ (.Y(_1378_),
    .A(net228));
 sg13g2_inv_1 _2332_ (.Y(_1379_),
    .A(net256));
 sg13g2_inv_1 _2333_ (.Y(_1380_),
    .A(net262));
 sg13g2_inv_1 _2334_ (.Y(_1381_),
    .A(net214));
 sg13g2_inv_1 _2335_ (.Y(_1382_),
    .A(net218));
 sg13g2_inv_1 _2336_ (.Y(_1383_),
    .A(net217));
 sg13g2_inv_1 _2337_ (.Y(_1384_),
    .A(net247));
 sg13g2_inv_1 _2338_ (.Y(_1385_),
    .A(net260));
 sg13g2_inv_1 _2339_ (.Y(_1386_),
    .A(net258));
 sg13g2_inv_1 _2340_ (.Y(_1387_),
    .A(net257));
 sg13g2_inv_1 _2341_ (.Y(_1388_),
    .A(net249));
 sg13g2_inv_1 _2342_ (.Y(_1389_),
    .A(net236));
 sg13g2_inv_1 _2343_ (.Y(_1390_),
    .A(net229));
 sg13g2_inv_1 _2344_ (.Y(_1391_),
    .A(net785));
 sg13g2_inv_1 _2345_ (.Y(_1392_),
    .A(net853));
 sg13g2_inv_1 _2346_ (.Y(_1393_),
    .A(\collatz.iter[142] ));
 sg13g2_inv_1 _2347_ (.Y(_1394_),
    .A(\collatz.iter[141] ));
 sg13g2_inv_1 _2348_ (.Y(_1395_),
    .A(\collatz.iter[140] ));
 sg13g2_inv_1 _2349_ (.Y(_1396_),
    .A(\collatz.iter[139] ));
 sg13g2_inv_1 _2350_ (.Y(_1397_),
    .A(\collatz.iter[137] ));
 sg13g2_inv_1 _2351_ (.Y(_1398_),
    .A(\collatz.iter[136] ));
 sg13g2_inv_1 _2352_ (.Y(_1399_),
    .A(\collatz.iter[135] ));
 sg13g2_inv_1 _2353_ (.Y(_1400_),
    .A(\collatz.iter[133] ));
 sg13g2_inv_1 _2354_ (.Y(_1401_),
    .A(\collatz.iter[132] ));
 sg13g2_inv_1 _2355_ (.Y(_1402_),
    .A(\collatz.iter[98] ));
 sg13g2_inv_1 _2356_ (.Y(_1403_),
    .A(\collatz.iter[86] ));
 sg13g2_inv_1 _2357_ (.Y(_1404_),
    .A(\collatz.iter[30] ));
 sg13g2_inv_1 _2358_ (.Y(_1405_),
    .A(\collatz.iter[26] ));
 sg13g2_inv_1 _2359_ (.Y(_1406_),
    .A(\collatz.iter[17] ));
 sg13g2_inv_1 _2360_ (.Y(_1407_),
    .A(\collatz.iter[16] ));
 sg13g2_inv_1 _2361_ (.Y(_1408_),
    .A(\collatz.iter[15] ));
 sg13g2_inv_1 _2362_ (.Y(_1409_),
    .A(\collatz.iter[14] ));
 sg13g2_inv_1 _2363_ (.Y(_1410_),
    .A(\collatz.iter[13] ));
 sg13g2_inv_1 _2364_ (.Y(_1411_),
    .A(\collatz.iter[12] ));
 sg13g2_inv_1 _2365_ (.Y(_1412_),
    .A(\collatz.iter[11] ));
 sg13g2_inv_1 _2366_ (.Y(_1413_),
    .A(net713));
 sg13g2_inv_1 _2367_ (.Y(_1414_),
    .A(_0008_));
 sg13g2_inv_1 _2368_ (.Y(_1415_),
    .A(_0005_));
 sg13g2_inv_1 _2369_ (.Y(_1416_),
    .A(_0007_));
 sg13g2_inv_2 _2370_ (.Y(_1417_),
    .A(net7));
 sg13g2_inv_1 _2371_ (.Y(_1418_),
    .A(net1));
 sg13g2_inv_4 _2372_ (.A(net829),
    .Y(_1419_));
 sg13g2_and2_1 _2373_ (.A(\collatz.orbit_len[13] ),
    .B(\collatz.orbit_len[12] ),
    .X(_1420_));
 sg13g2_nand4_1 _2374_ (.B(\collatz.orbit_len[10] ),
    .C(\collatz.orbit_len[9] ),
    .A(net219),
    .Y(_1421_),
    .D(_1420_));
 sg13g2_nand3_1 _2375_ (.B(net238),
    .C(net246),
    .A(net224),
    .Y(_1422_));
 sg13g2_nand3_1 _2376_ (.B(net210),
    .C(net336),
    .A(net226),
    .Y(_1423_));
 sg13g2_nand4_1 _2377_ (.B(\collatz.orbit_len[8] ),
    .C(\collatz.orbit_len[7] ),
    .A(\collatz.orbit_len[14] ),
    .Y(_1424_),
    .D(\collatz.orbit_len[3] ));
 sg13g2_or4_1 _2378_ (.A(_1421_),
    .B(_1422_),
    .C(_1423_),
    .D(_1424_),
    .X(_1425_));
 sg13g2_o21ai_1 _2379_ (.B1(net787),
    .Y(_1426_),
    .A1(_1390_),
    .A2(_1425_));
 sg13g2_nor2_1 _2380_ (.A(net702),
    .B(\collatz.iter[60] ),
    .Y(_1427_));
 sg13g2_nor2_2 _2381_ (.A(\collatz.iter[21] ),
    .B(\collatz.iter[20] ),
    .Y(_1428_));
 sg13g2_nor2_2 _2382_ (.A(net711),
    .B(\collatz.iter[2] ),
    .Y(_1429_));
 sg13g2_nor2_1 _2383_ (.A(\collatz.iter[65] ),
    .B(\collatz.iter[64] ),
    .Y(_1430_));
 sg13g2_nor2_1 _2384_ (.A(\collatz.iter[73] ),
    .B(\collatz.iter[72] ),
    .Y(_1431_));
 sg13g2_nor2_1 _2385_ (.A(net709),
    .B(\collatz.iter[32] ),
    .Y(_1432_));
 sg13g2_nor2_1 _2386_ (.A(\collatz.iter[77] ),
    .B(\collatz.iter[76] ),
    .Y(_1433_));
 sg13g2_nor2_1 _2387_ (.A(net803),
    .B(\collatz.iter[124] ),
    .Y(_1434_));
 sg13g2_nor2_2 _2388_ (.A(\collatz.iter[139] ),
    .B(\collatz.iter[138] ),
    .Y(_1435_));
 sg13g2_nor2_2 _2389_ (.A(\collatz.iter[49] ),
    .B(\collatz.iter[48] ),
    .Y(_1436_));
 sg13g2_nor2_1 _2390_ (.A(\collatz.iter[93] ),
    .B(\collatz.iter[92] ),
    .Y(_1437_));
 sg13g2_nor2_2 _2391_ (.A(net697),
    .B(\collatz.iter[114] ),
    .Y(_1438_));
 sg13g2_nor2_1 _2392_ (.A(net706),
    .B(\collatz.iter[44] ),
    .Y(_1439_));
 sg13g2_nor2_1 _2393_ (.A(\collatz.iter[67] ),
    .B(\collatz.iter[66] ),
    .Y(_1440_));
 sg13g2_nor2_2 _2394_ (.A(\collatz.iter[5] ),
    .B(\collatz.iter[4] ),
    .Y(_1441_));
 sg13g2_nor2_1 _2395_ (.A(\collatz.iter[129] ),
    .B(\collatz.iter[128] ),
    .Y(_1442_));
 sg13g2_nor2_1 _2396_ (.A(net707),
    .B(\collatz.iter[40] ),
    .Y(_1443_));
 sg13g2_nor2_1 _2397_ (.A(net703),
    .B(net704),
    .Y(_1444_));
 sg13g2_nor2_1 _2398_ (.A(\collatz.iter[101] ),
    .B(\collatz.iter[100] ),
    .Y(_1445_));
 sg13g2_nor2_1 _2399_ (.A(\collatz.iter[133] ),
    .B(\collatz.iter[132] ),
    .Y(_1446_));
 sg13g2_nor2_1 _2400_ (.A(\collatz.iter[9] ),
    .B(\collatz.iter[8] ),
    .Y(_1447_));
 sg13g2_nor2_1 _2401_ (.A(\collatz.iter[89] ),
    .B(\collatz.iter[88] ),
    .Y(_1448_));
 sg13g2_nor2_1 _2402_ (.A(net708),
    .B(\collatz.iter[36] ),
    .Y(_1449_));
 sg13g2_nor2_2 _2403_ (.A(\collatz.iter[121] ),
    .B(\collatz.iter[120] ),
    .Y(_1450_));
 sg13g2_nand2_1 _2404_ (.Y(_1451_),
    .A(net305),
    .B(net682));
 sg13g2_nor2_1 _2405_ (.A(net710),
    .B(\collatz.iter[24] ),
    .Y(_1452_));
 sg13g2_nor2_1 _2406_ (.A(net699),
    .B(\collatz.iter[96] ),
    .Y(_1453_));
 sg13g2_nor2_2 _2407_ (.A(\collatz.iter[117] ),
    .B(\collatz.iter[116] ),
    .Y(_1454_));
 sg13g2_nor2_2 _2408_ (.A(\collatz.iter[105] ),
    .B(\collatz.iter[104] ),
    .Y(_1455_));
 sg13g2_nor2_1 _2409_ (.A(\collatz.iter[29] ),
    .B(\collatz.iter[28] ),
    .Y(_1456_));
 sg13g2_nor2_2 _2410_ (.A(\collatz.iter[57] ),
    .B(\collatz.iter[56] ),
    .Y(_1457_));
 sg13g2_nor2_1 _2411_ (.A(\collatz.iter[69] ),
    .B(\collatz.iter[68] ),
    .Y(_1458_));
 sg13g2_or2_1 _2412_ (.X(_1459_),
    .B(\collatz.iter[130] ),
    .A(\collatz.iter[131] ));
 sg13g2_nor2_1 _2413_ (.A(\collatz.iter[109] ),
    .B(\collatz.iter[108] ),
    .Y(_1460_));
 sg13g2_nor2_1 _2414_ (.A(\collatz.iter[81] ),
    .B(\collatz.iter[80] ),
    .Y(_1461_));
 sg13g2_nor2_1 _2415_ (.A(\collatz.iter[85] ),
    .B(\collatz.iter[84] ),
    .Y(_1462_));
 sg13g2_nor4_1 _2416_ (.A(\collatz.iter[113] ),
    .B(\collatz.iter[112] ),
    .C(\collatz.iter[11] ),
    .D(\collatz.iter[10] ),
    .Y(_1463_));
 sg13g2_nor4_2 _2417_ (.A(net803),
    .B(\collatz.iter[124] ),
    .C(\collatz.iter[123] ),
    .Y(_1464_),
    .D(\collatz.iter[122] ));
 sg13g2_nor4_1 _2418_ (.A(\collatz.iter[91] ),
    .B(\collatz.iter[90] ),
    .C(\collatz.iter[75] ),
    .D(\collatz.iter[74] ),
    .Y(_1465_));
 sg13g2_nor4_1 _2419_ (.A(\collatz.iter[103] ),
    .B(\collatz.iter[102] ),
    .C(\collatz.iter[87] ),
    .D(\collatz.iter[86] ),
    .Y(_1466_));
 sg13g2_nand4_1 _2420_ (.B(_1464_),
    .C(_1465_),
    .A(_1463_),
    .Y(_1467_),
    .D(_1466_));
 sg13g2_nor4_2 _2421_ (.A(\collatz.iter[141] ),
    .B(\collatz.iter[140] ),
    .C(\collatz.iter[13] ),
    .Y(_1468_),
    .D(\collatz.iter[12] ));
 sg13g2_and2_1 _2422_ (.A(_1445_),
    .B(_1453_),
    .X(_1469_));
 sg13g2_nor4_1 _2423_ (.A(\collatz.iter[79] ),
    .B(\collatz.iter[78] ),
    .C(\collatz.iter[51] ),
    .D(\collatz.iter[50] ),
    .Y(_1470_));
 sg13g2_and2_1 _2424_ (.A(_1437_),
    .B(_1450_),
    .X(_1471_));
 sg13g2_nand4_1 _2425_ (.B(_1469_),
    .C(_1470_),
    .A(_1468_),
    .Y(_1472_),
    .D(_1471_));
 sg13g2_nor3_2 _2426_ (.A(\collatz.iter[15] ),
    .B(\collatz.iter[14] ),
    .C(_1451_),
    .Y(_1473_));
 sg13g2_and4_1 _2427_ (.A(_1397_),
    .B(_1398_),
    .C(_1454_),
    .D(_1473_),
    .X(_1474_));
 sg13g2_nor4_2 _2428_ (.A(\collatz.iter[127] ),
    .B(\collatz.iter[126] ),
    .C(\collatz.iter[63] ),
    .Y(_1475_),
    .D(\collatz.iter[62] ));
 sg13g2_nand4_1 _2429_ (.B(_1455_),
    .C(_1474_),
    .A(_1438_),
    .Y(_1476_),
    .D(_1475_));
 sg13g2_nor4_2 _2430_ (.A(\collatz.iter[95] ),
    .B(\collatz.iter[94] ),
    .C(net700),
    .Y(_1477_),
    .D(\collatz.iter[84] ));
 sg13g2_nor4_1 _2431_ (.A(\collatz.iter[135] ),
    .B(\collatz.iter[134] ),
    .C(\collatz.iter[71] ),
    .D(\collatz.iter[70] ),
    .Y(_1478_));
 sg13g2_nor4_2 _2432_ (.A(\collatz.iter[119] ),
    .B(\collatz.iter[118] ),
    .C(net703),
    .Y(_1479_),
    .D(net704));
 sg13g2_and2_1 _2433_ (.A(_1478_),
    .B(_1479_),
    .X(_1480_));
 sg13g2_nand4_1 _2434_ (.B(_1458_),
    .C(_1477_),
    .A(_1436_),
    .Y(_1481_),
    .D(_1480_));
 sg13g2_nor4_2 _2435_ (.A(_1467_),
    .B(_1472_),
    .C(_1476_),
    .Y(_1482_),
    .D(_1481_));
 sg13g2_nor4_2 _2436_ (.A(net707),
    .B(\collatz.iter[40] ),
    .C(\collatz.iter[35] ),
    .Y(_1483_),
    .D(\collatz.iter[34] ));
 sg13g2_nor4_1 _2437_ (.A(\collatz.iter[45] ),
    .B(\collatz.iter[44] ),
    .C(\collatz.iter[17] ),
    .D(\collatz.iter[16] ),
    .Y(_1484_));
 sg13g2_nor4_2 _2438_ (.A(\collatz.iter[55] ),
    .B(\collatz.iter[54] ),
    .C(\collatz.iter[39] ),
    .Y(_1485_),
    .D(\collatz.iter[38] ));
 sg13g2_nor4_2 _2439_ (.A(\collatz.iter[25] ),
    .B(\collatz.iter[24] ),
    .C(\collatz.iter[19] ),
    .Y(_1486_),
    .D(\collatz.iter[18] ));
 sg13g2_nand4_1 _2440_ (.B(_1484_),
    .C(_1485_),
    .A(_1483_),
    .Y(_1487_),
    .D(_1486_));
 sg13g2_nor4_2 _2441_ (.A(\collatz.iter[47] ),
    .B(\collatz.iter[46] ),
    .C(\collatz.iter[31] ),
    .Y(_1488_),
    .D(\collatz.iter[30] ));
 sg13g2_nor4_2 _2442_ (.A(\collatz.iter[107] ),
    .B(\collatz.iter[106] ),
    .C(net701),
    .Y(_1489_),
    .D(\collatz.iter[80] ));
 sg13g2_and2_1 _2443_ (.A(_1488_),
    .B(_1489_),
    .X(_1490_));
 sg13g2_nor4_1 _2444_ (.A(\collatz.iter[33] ),
    .B(\collatz.iter[32] ),
    .C(\collatz.iter[27] ),
    .D(\collatz.iter[26] ),
    .Y(_1491_));
 sg13g2_nand4_1 _2445_ (.B(_1460_),
    .C(_1490_),
    .A(_1429_),
    .Y(_1492_),
    .D(_1491_));
 sg13g2_nor4_2 _2446_ (.A(\collatz.iter[23] ),
    .B(\collatz.iter[22] ),
    .C(\collatz.iter[7] ),
    .Y(_1493_),
    .D(\collatz.iter[6] ));
 sg13g2_nor4_2 _2447_ (.A(\collatz.iter[59] ),
    .B(\collatz.iter[58] ),
    .C(\collatz.iter[37] ),
    .Y(_1494_),
    .D(\collatz.iter[36] ));
 sg13g2_and2_1 _2448_ (.A(_1493_),
    .B(_1494_),
    .X(_1495_));
 sg13g2_nor4_2 _2449_ (.A(\collatz.iter[61] ),
    .B(\collatz.iter[60] ),
    .C(\collatz.iter[43] ),
    .Y(_1496_),
    .D(\collatz.iter[42] ));
 sg13g2_nand4_1 _2450_ (.B(_1456_),
    .C(_1495_),
    .A(_1428_),
    .Y(_1497_),
    .D(_1496_));
 sg13g2_or3_2 _2451_ (.A(_1487_),
    .B(_1492_),
    .C(_1497_),
    .X(_1498_));
 sg13g2_nand2_1 _2452_ (.Y(_1499_),
    .A(_1446_),
    .B(_1457_));
 sg13g2_nor4_1 _2453_ (.A(\collatz.iter[9] ),
    .B(\collatz.iter[8] ),
    .C(_1459_),
    .D(_1499_),
    .Y(_1500_));
 sg13g2_nor4_2 _2454_ (.A(\collatz.iter[111] ),
    .B(\collatz.iter[110] ),
    .C(\collatz.iter[99] ),
    .Y(_1501_),
    .D(\collatz.iter[98] ));
 sg13g2_nor4_2 _2455_ (.A(\collatz.iter[143] ),
    .B(\collatz.iter[142] ),
    .C(\collatz.iter[83] ),
    .Y(_1502_),
    .D(\collatz.iter[82] ));
 sg13g2_nand3_1 _2456_ (.B(_1501_),
    .C(_1502_),
    .A(_1500_),
    .Y(_1503_));
 sg13g2_nand4_1 _2457_ (.B(_1440_),
    .C(_1441_),
    .A(_1433_),
    .Y(_1504_),
    .D(_1448_));
 sg13g2_nand4_1 _2458_ (.B(_1431_),
    .C(_1435_),
    .A(_1430_),
    .Y(_1505_),
    .D(_1442_));
 sg13g2_nor4_2 _2459_ (.A(_1498_),
    .B(_1503_),
    .C(_1504_),
    .Y(_1506_),
    .D(_1505_));
 sg13g2_a21oi_2 _2460_ (.B1(_1426_),
    .Y(\collatz.busy ),
    .A2(_1506_),
    .A1(_1482_));
 sg13g2_nor2_1 _2461_ (.A(net692),
    .B(\collatz.busy ),
    .Y(_1507_));
 sg13g2_nor3_2 _2462_ (.A(net691),
    .B(net816),
    .C(\collatz.busy ),
    .Y(_1508_));
 sg13g2_and3_2 _2463_ (.X(_1509_),
    .A(net1),
    .B(net826),
    .C(_1419_));
 sg13g2_nor2_1 _2464_ (.A(net1),
    .B(net826),
    .Y(_1510_));
 sg13g2_nor3_2 _2465_ (.A(net1),
    .B(net826),
    .C(net828),
    .Y(_1511_));
 sg13g2_nor2b_2 _2466_ (.A(net3),
    .B_N(_1511_),
    .Y(_1512_));
 sg13g2_xnor2_1 _2467_ (.Y(_1513_),
    .A(net3),
    .B(_1511_));
 sg13g2_xnor2_1 _2468_ (.Y(_1514_),
    .A(net4),
    .B(_1512_));
 sg13g2_and2_1 _2469_ (.A(net7),
    .B(_1514_),
    .X(_1515_));
 sg13g2_nor2b_2 _2470_ (.A(_1513_),
    .B_N(net662),
    .Y(_1516_));
 sg13g2_a21oi_2 _2471_ (.B1(net650),
    .Y(_1517_),
    .A2(net655),
    .A1(net679));
 sg13g2_and2_1 _2472_ (.A(net830),
    .B(net679),
    .X(_1518_));
 sg13g2_a22oi_1 _2473_ (.Y(_1519_),
    .B1(_1518_),
    .B2(net654),
    .A2(_1517_),
    .A1(\collatz.iter[119] ));
 sg13g2_or2_1 _2474_ (.X(_1520_),
    .B(_1519_),
    .A(net760));
 sg13g2_xor2_1 _2475_ (.B(\collatz.iter[118] ),
    .A(\collatz.iter[119] ),
    .X(_1521_));
 sg13g2_and2_1 _2476_ (.A(\collatz.iter[118] ),
    .B(\collatz.iter[117] ),
    .X(_1522_));
 sg13g2_xor2_1 _2477_ (.B(\collatz.iter[117] ),
    .A(\collatz.iter[118] ),
    .X(_1523_));
 sg13g2_nand2_1 _2478_ (.Y(_1524_),
    .A(\collatz.iter[116] ),
    .B(net697));
 sg13g2_o21ai_1 _2479_ (.B1(\collatz.iter[116] ),
    .Y(_1525_),
    .A1(\collatz.iter[117] ),
    .A2(net697));
 sg13g2_inv_1 _2480_ (.Y(_1526_),
    .A(_1525_));
 sg13g2_xnor2_1 _2481_ (.Y(_1527_),
    .A(\collatz.iter[116] ),
    .B(net697));
 sg13g2_nand2_1 _2482_ (.Y(_1528_),
    .A(\collatz.iter[114] ),
    .B(net698));
 sg13g2_nand2_1 _2483_ (.Y(_1529_),
    .A(net697),
    .B(\collatz.iter[114] ));
 sg13g2_o21ai_1 _2484_ (.B1(\collatz.iter[114] ),
    .Y(_1530_),
    .A1(net697),
    .A2(net698));
 sg13g2_nand2_1 _2485_ (.Y(_1531_),
    .A(_1528_),
    .B(_1529_));
 sg13g2_nand2_1 _2486_ (.Y(_1532_),
    .A(\collatz.iter[112] ),
    .B(\collatz.iter[111] ));
 sg13g2_xnor2_1 _2487_ (.Y(_1533_),
    .A(\collatz.iter[112] ),
    .B(\collatz.iter[111] ));
 sg13g2_and2_1 _2488_ (.A(\collatz.iter[110] ),
    .B(\collatz.iter[109] ),
    .X(_1534_));
 sg13g2_xor2_1 _2489_ (.B(\collatz.iter[109] ),
    .A(\collatz.iter[110] ),
    .X(_1535_));
 sg13g2_xor2_1 _2490_ (.B(\collatz.iter[110] ),
    .A(\collatz.iter[111] ),
    .X(_1536_));
 sg13g2_and2_1 _2491_ (.A(_1535_),
    .B(_1536_),
    .X(_1537_));
 sg13g2_nand2_1 _2492_ (.Y(_1538_),
    .A(_1535_),
    .B(_1536_));
 sg13g2_nand2_1 _2493_ (.Y(_1539_),
    .A(\collatz.iter[108] ),
    .B(\collatz.iter[107] ));
 sg13g2_o21ai_1 _2494_ (.B1(\collatz.iter[108] ),
    .Y(_1540_),
    .A1(\collatz.iter[109] ),
    .A2(\collatz.iter[107] ));
 sg13g2_xor2_1 _2495_ (.B(\collatz.iter[107] ),
    .A(\collatz.iter[108] ),
    .X(_1541_));
 sg13g2_xor2_1 _2496_ (.B(\collatz.iter[108] ),
    .A(\collatz.iter[109] ),
    .X(_1542_));
 sg13g2_nand2_1 _2497_ (.Y(_1543_),
    .A(_1541_),
    .B(_1542_));
 sg13g2_and2_1 _2498_ (.A(\collatz.iter[106] ),
    .B(\collatz.iter[105] ),
    .X(_1544_));
 sg13g2_xor2_1 _2499_ (.B(\collatz.iter[105] ),
    .A(\collatz.iter[106] ),
    .X(_1545_));
 sg13g2_xor2_1 _2500_ (.B(\collatz.iter[106] ),
    .A(\collatz.iter[107] ),
    .X(_1546_));
 sg13g2_nand2_1 _2501_ (.Y(_1547_),
    .A(\collatz.iter[104] ),
    .B(\collatz.iter[103] ));
 sg13g2_o21ai_1 _2502_ (.B1(\collatz.iter[104] ),
    .Y(_1548_),
    .A1(\collatz.iter[105] ),
    .A2(\collatz.iter[103] ));
 sg13g2_nand3b_1 _2503_ (.B(_1546_),
    .C(_1545_),
    .Y(_1549_),
    .A_N(_1548_));
 sg13g2_o21ai_1 _2504_ (.B1(\collatz.iter[106] ),
    .Y(_1550_),
    .A1(\collatz.iter[107] ),
    .A2(\collatz.iter[105] ));
 sg13g2_and2_1 _2505_ (.A(_1549_),
    .B(_1550_),
    .X(_1551_));
 sg13g2_o21ai_1 _2506_ (.B1(_1540_),
    .Y(_1552_),
    .A1(_1543_),
    .A2(_1551_));
 sg13g2_xor2_1 _2507_ (.B(\collatz.iter[104] ),
    .A(\collatz.iter[105] ),
    .X(_1553_));
 sg13g2_xor2_1 _2508_ (.B(\collatz.iter[103] ),
    .A(\collatz.iter[104] ),
    .X(_1554_));
 sg13g2_nand4_1 _2509_ (.B(_1546_),
    .C(_1553_),
    .A(_1545_),
    .Y(_1555_),
    .D(_1554_));
 sg13g2_nor3_2 _2510_ (.A(_1538_),
    .B(_1543_),
    .C(_1555_),
    .Y(_1556_));
 sg13g2_and2_1 _2511_ (.A(\collatz.iter[102] ),
    .B(\collatz.iter[101] ),
    .X(_1557_));
 sg13g2_xor2_1 _2512_ (.B(\collatz.iter[101] ),
    .A(\collatz.iter[102] ),
    .X(_1558_));
 sg13g2_xnor2_1 _2513_ (.Y(_1559_),
    .A(\collatz.iter[102] ),
    .B(\collatz.iter[101] ));
 sg13g2_nand2_1 _2514_ (.Y(_1560_),
    .A(\collatz.iter[103] ),
    .B(\collatz.iter[102] ));
 sg13g2_xnor2_1 _2515_ (.Y(_1561_),
    .A(\collatz.iter[103] ),
    .B(\collatz.iter[102] ));
 sg13g2_xnor2_1 _2516_ (.Y(_1562_),
    .A(\collatz.iter[101] ),
    .B(\collatz.iter[100] ));
 sg13g2_nand2_1 _2517_ (.Y(_1563_),
    .A(\collatz.iter[100] ),
    .B(\collatz.iter[99] ));
 sg13g2_xnor2_1 _2518_ (.Y(_1564_),
    .A(\collatz.iter[100] ),
    .B(\collatz.iter[99] ));
 sg13g2_nor4_2 _2519_ (.A(_1559_),
    .B(_1561_),
    .C(_1562_),
    .Y(_1565_),
    .D(_1564_));
 sg13g2_and2_1 _2520_ (.A(\collatz.iter[98] ),
    .B(net699),
    .X(_1566_));
 sg13g2_xor2_1 _2521_ (.B(net699),
    .A(\collatz.iter[98] ),
    .X(_1567_));
 sg13g2_xnor2_1 _2522_ (.Y(_1568_),
    .A(\collatz.iter[98] ),
    .B(net699));
 sg13g2_xnor2_1 _2523_ (.Y(_1569_),
    .A(\collatz.iter[99] ),
    .B(\collatz.iter[98] ));
 sg13g2_nand2_1 _2524_ (.Y(_1570_),
    .A(\collatz.iter[96] ),
    .B(\collatz.iter[95] ));
 sg13g2_o21ai_1 _2525_ (.B1(\collatz.iter[96] ),
    .Y(_1571_),
    .A1(net699),
    .A2(\collatz.iter[95] ));
 sg13g2_nor3_1 _2526_ (.A(_1568_),
    .B(_1569_),
    .C(_1571_),
    .Y(_1572_));
 sg13g2_o21ai_1 _2527_ (.B1(\collatz.iter[98] ),
    .Y(_1573_),
    .A1(\collatz.iter[99] ),
    .A2(net699));
 sg13g2_inv_1 _2528_ (.Y(_1574_),
    .A(_1573_));
 sg13g2_nand2b_1 _2529_ (.Y(_1575_),
    .B(_1573_),
    .A_N(_1572_));
 sg13g2_o21ai_1 _2530_ (.B1(_1565_),
    .Y(_1576_),
    .A1(_1572_),
    .A2(_1574_));
 sg13g2_o21ai_1 _2531_ (.B1(\collatz.iter[100] ),
    .Y(_1577_),
    .A1(\collatz.iter[101] ),
    .A2(\collatz.iter[99] ));
 sg13g2_nor3_1 _2532_ (.A(_1559_),
    .B(_1561_),
    .C(_1577_),
    .Y(_1578_));
 sg13g2_nor2_1 _2533_ (.A(_1557_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_nand3_1 _2534_ (.B(_1576_),
    .C(_1579_),
    .A(_1560_),
    .Y(_1580_));
 sg13g2_o21ai_1 _2535_ (.B1(\collatz.iter[110] ),
    .Y(_1581_),
    .A1(\collatz.iter[111] ),
    .A2(\collatz.iter[109] ));
 sg13g2_inv_1 _2536_ (.Y(_1582_),
    .A(_1581_));
 sg13g2_a21o_1 _2537_ (.A2(_1552_),
    .A1(_1537_),
    .B1(_1582_),
    .X(_1583_));
 sg13g2_a221oi_1 _2538_ (.B2(_1580_),
    .C1(_1582_),
    .B1(_1556_),
    .A1(_1537_),
    .Y(_1584_),
    .A2(_1552_));
 sg13g2_xor2_1 _2539_ (.B(\collatz.iter[95] ),
    .A(\collatz.iter[96] ),
    .X(_1585_));
 sg13g2_xnor2_1 _2540_ (.Y(_1586_),
    .A(\collatz.iter[97] ),
    .B(\collatz.iter[96] ));
 sg13g2_nor3_1 _2541_ (.A(_1568_),
    .B(_1569_),
    .C(_1586_),
    .Y(_1587_));
 sg13g2_and2_1 _2542_ (.A(_1585_),
    .B(_1587_),
    .X(_1588_));
 sg13g2_and2_1 _2543_ (.A(_1565_),
    .B(_1588_),
    .X(_1589_));
 sg13g2_and2_1 _2544_ (.A(_1556_),
    .B(_1589_),
    .X(_1590_));
 sg13g2_and2_1 _2545_ (.A(\collatz.iter[94] ),
    .B(\collatz.iter[93] ),
    .X(_1591_));
 sg13g2_xor2_1 _2546_ (.B(\collatz.iter[93] ),
    .A(\collatz.iter[94] ),
    .X(_1592_));
 sg13g2_xor2_1 _2547_ (.B(\collatz.iter[94] ),
    .A(\collatz.iter[95] ),
    .X(_1593_));
 sg13g2_nand2_1 _2548_ (.Y(_1594_),
    .A(_1592_),
    .B(_1593_));
 sg13g2_inv_1 _2549_ (.Y(_1595_),
    .A(_1594_));
 sg13g2_nand2_1 _2550_ (.Y(_1596_),
    .A(\collatz.iter[92] ),
    .B(\collatz.iter[91] ));
 sg13g2_o21ai_1 _2551_ (.B1(\collatz.iter[92] ),
    .Y(_1597_),
    .A1(\collatz.iter[93] ),
    .A2(\collatz.iter[91] ));
 sg13g2_xor2_1 _2552_ (.B(\collatz.iter[91] ),
    .A(\collatz.iter[92] ),
    .X(_1598_));
 sg13g2_xor2_1 _2553_ (.B(\collatz.iter[92] ),
    .A(\collatz.iter[93] ),
    .X(_1599_));
 sg13g2_nand2_1 _2554_ (.Y(_1600_),
    .A(_1598_),
    .B(_1599_));
 sg13g2_xnor2_1 _2555_ (.Y(_1601_),
    .A(\collatz.iter[90] ),
    .B(\collatz.iter[89] ));
 sg13g2_xnor2_1 _2556_ (.Y(_1602_),
    .A(\collatz.iter[91] ),
    .B(\collatz.iter[90] ));
 sg13g2_nand2_1 _2557_ (.Y(_1603_),
    .A(\collatz.iter[88] ),
    .B(\collatz.iter[87] ));
 sg13g2_o21ai_1 _2558_ (.B1(\collatz.iter[88] ),
    .Y(_1604_),
    .A1(\collatz.iter[89] ),
    .A2(\collatz.iter[87] ));
 sg13g2_nor3_1 _2559_ (.A(_1601_),
    .B(_1602_),
    .C(_1604_),
    .Y(_1605_));
 sg13g2_o21ai_1 _2560_ (.B1(\collatz.iter[90] ),
    .Y(_1606_),
    .A1(\collatz.iter[91] ),
    .A2(\collatz.iter[89] ));
 sg13g2_nor2b_1 _2561_ (.A(_1605_),
    .B_N(_1606_),
    .Y(_1607_));
 sg13g2_o21ai_1 _2562_ (.B1(_1597_),
    .Y(_1608_),
    .A1(_1600_),
    .A2(_1607_));
 sg13g2_o21ai_1 _2563_ (.B1(\collatz.iter[94] ),
    .Y(_1609_),
    .A1(\collatz.iter[95] ),
    .A2(\collatz.iter[93] ));
 sg13g2_inv_1 _2564_ (.Y(_1610_),
    .A(_1609_));
 sg13g2_xor2_1 _2565_ (.B(\collatz.iter[88] ),
    .A(\collatz.iter[89] ),
    .X(_1611_));
 sg13g2_xnor2_1 _2566_ (.Y(_1612_),
    .A(\collatz.iter[88] ),
    .B(\collatz.iter[87] ));
 sg13g2_nor3_1 _2567_ (.A(_1601_),
    .B(_1602_),
    .C(_1612_),
    .Y(_1613_));
 sg13g2_nand2_1 _2568_ (.Y(_1614_),
    .A(_1611_),
    .B(_1613_));
 sg13g2_nor3_2 _2569_ (.A(_1594_),
    .B(_1600_),
    .C(_1614_),
    .Y(_1615_));
 sg13g2_xnor2_1 _2570_ (.Y(_1616_),
    .A(\collatz.iter[86] ),
    .B(net700));
 sg13g2_xnor2_1 _2571_ (.Y(_1617_),
    .A(\collatz.iter[87] ),
    .B(\collatz.iter[86] ));
 sg13g2_xnor2_1 _2572_ (.Y(_1618_),
    .A(net700),
    .B(\collatz.iter[84] ));
 sg13g2_nand2_1 _2573_ (.Y(_1619_),
    .A(\collatz.iter[84] ),
    .B(\collatz.iter[83] ));
 sg13g2_xnor2_1 _2574_ (.Y(_1620_),
    .A(\collatz.iter[84] ),
    .B(\collatz.iter[83] ));
 sg13g2_nor4_1 _2575_ (.A(_1616_),
    .B(_1617_),
    .C(_1618_),
    .D(_1620_),
    .Y(_1621_));
 sg13g2_and2_1 _2576_ (.A(\collatz.iter[82] ),
    .B(net701),
    .X(_1622_));
 sg13g2_xor2_1 _2577_ (.B(net701),
    .A(\collatz.iter[82] ),
    .X(_1623_));
 sg13g2_xor2_1 _2578_ (.B(\collatz.iter[82] ),
    .A(\collatz.iter[83] ),
    .X(_1624_));
 sg13g2_nand2_1 _2579_ (.Y(_1625_),
    .A(_1623_),
    .B(_1624_));
 sg13g2_nand2_1 _2580_ (.Y(_1626_),
    .A(\collatz.iter[80] ),
    .B(\collatz.iter[79] ));
 sg13g2_o21ai_1 _2581_ (.B1(\collatz.iter[80] ),
    .Y(_1627_),
    .A1(net701),
    .A2(\collatz.iter[79] ));
 sg13g2_o21ai_1 _2582_ (.B1(\collatz.iter[82] ),
    .Y(_1628_),
    .A1(\collatz.iter[83] ),
    .A2(net701));
 sg13g2_o21ai_1 _2583_ (.B1(_1628_),
    .Y(_1629_),
    .A1(_1625_),
    .A2(_1627_));
 sg13g2_o21ai_1 _2584_ (.B1(\collatz.iter[86] ),
    .Y(_1630_),
    .A1(\collatz.iter[87] ),
    .A2(net700));
 sg13g2_o21ai_1 _2585_ (.B1(\collatz.iter[84] ),
    .Y(_1631_),
    .A1(net700),
    .A2(\collatz.iter[83] ));
 sg13g2_nor3_1 _2586_ (.A(_1616_),
    .B(_1617_),
    .C(_1631_),
    .Y(_1632_));
 sg13g2_nand2b_1 _2587_ (.Y(_1633_),
    .B(_1630_),
    .A_N(_1632_));
 sg13g2_a21o_1 _2588_ (.A2(_1629_),
    .A1(_1621_),
    .B1(_1633_),
    .X(_1634_));
 sg13g2_a221oi_1 _2589_ (.B2(_1634_),
    .C1(_1610_),
    .B1(_1615_),
    .A1(_1595_),
    .Y(_1635_),
    .A2(_1608_));
 sg13g2_and2_1 _2590_ (.A(\collatz.iter[78] ),
    .B(\collatz.iter[77] ),
    .X(_1636_));
 sg13g2_xor2_1 _2591_ (.B(\collatz.iter[77] ),
    .A(\collatz.iter[78] ),
    .X(_1637_));
 sg13g2_xor2_1 _2592_ (.B(\collatz.iter[78] ),
    .A(\collatz.iter[79] ),
    .X(_1638_));
 sg13g2_nand2_1 _2593_ (.Y(_1639_),
    .A(_1637_),
    .B(_1638_));
 sg13g2_xor2_1 _2594_ (.B(\collatz.iter[76] ),
    .A(\collatz.iter[77] ),
    .X(_1640_));
 sg13g2_nand2_1 _2595_ (.Y(_1641_),
    .A(\collatz.iter[76] ),
    .B(\collatz.iter[75] ));
 sg13g2_xor2_1 _2596_ (.B(\collatz.iter[75] ),
    .A(\collatz.iter[76] ),
    .X(_1642_));
 sg13g2_nand4_1 _2597_ (.B(_1638_),
    .C(_1640_),
    .A(_1637_),
    .Y(_1643_),
    .D(_1642_));
 sg13g2_inv_1 _2598_ (.Y(_1644_),
    .A(_1643_));
 sg13g2_and2_1 _2599_ (.A(\collatz.iter[74] ),
    .B(\collatz.iter[73] ),
    .X(_1645_));
 sg13g2_xor2_1 _2600_ (.B(\collatz.iter[73] ),
    .A(\collatz.iter[74] ),
    .X(_1646_));
 sg13g2_xor2_1 _2601_ (.B(\collatz.iter[74] ),
    .A(\collatz.iter[75] ),
    .X(_1647_));
 sg13g2_nand2_2 _2602_ (.Y(_1648_),
    .A(_1646_),
    .B(_1647_));
 sg13g2_nand2_1 _2603_ (.Y(_1649_),
    .A(\collatz.iter[72] ),
    .B(\collatz.iter[71] ));
 sg13g2_xor2_1 _2604_ (.B(\collatz.iter[71] ),
    .A(\collatz.iter[72] ),
    .X(_1650_));
 sg13g2_inv_1 _2605_ (.Y(_1651_),
    .A(_1650_));
 sg13g2_xnor2_1 _2606_ (.Y(_1652_),
    .A(\collatz.iter[73] ),
    .B(\collatz.iter[72] ));
 sg13g2_nor4_2 _2607_ (.A(_1643_),
    .B(_1648_),
    .C(_1651_),
    .Y(_1653_),
    .D(_1652_));
 sg13g2_and2_1 _2608_ (.A(\collatz.iter[70] ),
    .B(\collatz.iter[69] ),
    .X(_1654_));
 sg13g2_xor2_1 _2609_ (.B(\collatz.iter[69] ),
    .A(\collatz.iter[70] ),
    .X(_1655_));
 sg13g2_xor2_1 _2610_ (.B(\collatz.iter[70] ),
    .A(\collatz.iter[71] ),
    .X(_1656_));
 sg13g2_nand2_1 _2611_ (.Y(_1657_),
    .A(\collatz.iter[68] ),
    .B(\collatz.iter[67] ));
 sg13g2_xor2_1 _2612_ (.B(\collatz.iter[67] ),
    .A(\collatz.iter[68] ),
    .X(_1658_));
 sg13g2_xor2_1 _2613_ (.B(\collatz.iter[68] ),
    .A(\collatz.iter[69] ),
    .X(_1659_));
 sg13g2_nand4_1 _2614_ (.B(_1656_),
    .C(_1658_),
    .A(_1655_),
    .Y(_1660_),
    .D(_1659_));
 sg13g2_and2_1 _2615_ (.A(\collatz.iter[66] ),
    .B(\collatz.iter[65] ),
    .X(_1661_));
 sg13g2_xor2_1 _2616_ (.B(\collatz.iter[65] ),
    .A(\collatz.iter[66] ),
    .X(_1662_));
 sg13g2_xor2_1 _2617_ (.B(\collatz.iter[66] ),
    .A(\collatz.iter[67] ),
    .X(_1663_));
 sg13g2_nand2_1 _2618_ (.Y(_1664_),
    .A(\collatz.iter[64] ),
    .B(\collatz.iter[63] ));
 sg13g2_o21ai_1 _2619_ (.B1(\collatz.iter[64] ),
    .Y(_1665_),
    .A1(\collatz.iter[65] ),
    .A2(\collatz.iter[63] ));
 sg13g2_nand3b_1 _2620_ (.B(_1663_),
    .C(_1662_),
    .Y(_1666_),
    .A_N(_1665_));
 sg13g2_o21ai_1 _2621_ (.B1(\collatz.iter[66] ),
    .Y(_1667_),
    .A1(\collatz.iter[67] ),
    .A2(\collatz.iter[65] ));
 sg13g2_and2_1 _2622_ (.A(_1666_),
    .B(_1667_),
    .X(_1668_));
 sg13g2_o21ai_1 _2623_ (.B1(\collatz.iter[70] ),
    .Y(_1669_),
    .A1(\collatz.iter[71] ),
    .A2(\collatz.iter[69] ));
 sg13g2_o21ai_1 _2624_ (.B1(\collatz.iter[68] ),
    .Y(_1670_),
    .A1(\collatz.iter[69] ),
    .A2(\collatz.iter[67] ));
 sg13g2_nand3b_1 _2625_ (.B(_1656_),
    .C(_1655_),
    .Y(_1671_),
    .A_N(_1670_));
 sg13g2_and2_1 _2626_ (.A(_1669_),
    .B(_1671_),
    .X(_1672_));
 sg13g2_o21ai_1 _2627_ (.B1(_1672_),
    .Y(_1673_),
    .A1(_1660_),
    .A2(_1668_));
 sg13g2_o21ai_1 _2628_ (.B1(\collatz.iter[76] ),
    .Y(_1674_),
    .A1(\collatz.iter[77] ),
    .A2(\collatz.iter[75] ));
 sg13g2_o21ai_1 _2629_ (.B1(\collatz.iter[78] ),
    .Y(_1675_),
    .A1(\collatz.iter[79] ),
    .A2(\collatz.iter[77] ));
 sg13g2_o21ai_1 _2630_ (.B1(_1675_),
    .Y(_1676_),
    .A1(_1639_),
    .A2(_1674_));
 sg13g2_o21ai_1 _2631_ (.B1(\collatz.iter[72] ),
    .Y(_1677_),
    .A1(\collatz.iter[73] ),
    .A2(\collatz.iter[71] ));
 sg13g2_o21ai_1 _2632_ (.B1(\collatz.iter[74] ),
    .Y(_1678_),
    .A1(\collatz.iter[75] ),
    .A2(\collatz.iter[73] ));
 sg13g2_o21ai_1 _2633_ (.B1(_1678_),
    .Y(_1679_),
    .A1(_1648_),
    .A2(_1677_));
 sg13g2_a221oi_1 _2634_ (.B2(_1644_),
    .C1(_1676_),
    .B1(_1679_),
    .A1(_1653_),
    .Y(_1680_),
    .A2(_1673_));
 sg13g2_xor2_1 _2635_ (.B(\collatz.iter[79] ),
    .A(\collatz.iter[80] ),
    .X(_1681_));
 sg13g2_xor2_1 _2636_ (.B(\collatz.iter[80] ),
    .A(net701),
    .X(_1682_));
 sg13g2_and4_1 _2637_ (.A(_1623_),
    .B(_1624_),
    .C(_1681_),
    .D(_1682_),
    .X(_1683_));
 sg13g2_and2_2 _2638_ (.A(_1621_),
    .B(_1683_),
    .X(_1684_));
 sg13g2_nand2_1 _2639_ (.Y(_1685_),
    .A(_1615_),
    .B(_1684_));
 sg13g2_o21ai_1 _2640_ (.B1(_1635_),
    .Y(_1686_),
    .A1(_1680_),
    .A2(_1685_));
 sg13g2_xnor2_1 _2641_ (.Y(_1687_),
    .A(\collatz.iter[30] ),
    .B(\collatz.iter[29] ));
 sg13g2_xnor2_1 _2642_ (.Y(_1688_),
    .A(\collatz.iter[31] ),
    .B(\collatz.iter[30] ));
 sg13g2_xnor2_1 _2643_ (.Y(_1689_),
    .A(\collatz.iter[29] ),
    .B(\collatz.iter[28] ));
 sg13g2_nand2_1 _2644_ (.Y(_1690_),
    .A(\collatz.iter[28] ),
    .B(\collatz.iter[27] ));
 sg13g2_xnor2_1 _2645_ (.Y(_1691_),
    .A(\collatz.iter[28] ),
    .B(\collatz.iter[27] ));
 sg13g2_nor4_2 _2646_ (.A(_1687_),
    .B(_1688_),
    .C(_1689_),
    .Y(_1692_),
    .D(_1691_));
 sg13g2_and2_1 _2647_ (.A(\collatz.iter[26] ),
    .B(net710),
    .X(_1693_));
 sg13g2_xor2_1 _2648_ (.B(net710),
    .A(\collatz.iter[26] ),
    .X(_1694_));
 sg13g2_xnor2_1 _2649_ (.Y(_1695_),
    .A(\collatz.iter[26] ),
    .B(net710));
 sg13g2_xnor2_1 _2650_ (.Y(_1696_),
    .A(\collatz.iter[27] ),
    .B(\collatz.iter[26] ));
 sg13g2_nand2_1 _2651_ (.Y(_1697_),
    .A(\collatz.iter[24] ),
    .B(\collatz.iter[23] ));
 sg13g2_xor2_1 _2652_ (.B(\collatz.iter[23] ),
    .A(\collatz.iter[24] ),
    .X(_1698_));
 sg13g2_xnor2_1 _2653_ (.Y(_1699_),
    .A(net710),
    .B(\collatz.iter[24] ));
 sg13g2_nor3_1 _2654_ (.A(_1695_),
    .B(_1696_),
    .C(_1699_),
    .Y(_1700_));
 sg13g2_and2_1 _2655_ (.A(_1698_),
    .B(_1700_),
    .X(_1701_));
 sg13g2_and2_1 _2656_ (.A(_1692_),
    .B(_1701_),
    .X(_1702_));
 sg13g2_o21ai_1 _2657_ (.B1(\collatz.iter[28] ),
    .Y(_1703_),
    .A1(\collatz.iter[29] ),
    .A2(\collatz.iter[27] ));
 sg13g2_nor3_1 _2658_ (.A(_1687_),
    .B(_1688_),
    .C(_1703_),
    .Y(_1704_));
 sg13g2_o21ai_1 _2659_ (.B1(\collatz.iter[30] ),
    .Y(_1705_),
    .A1(\collatz.iter[31] ),
    .A2(\collatz.iter[29] ));
 sg13g2_nand2b_2 _2660_ (.Y(_1706_),
    .B(_1705_),
    .A_N(_1704_));
 sg13g2_o21ai_1 _2661_ (.B1(\collatz.iter[24] ),
    .Y(_1707_),
    .A1(\collatz.iter[25] ),
    .A2(\collatz.iter[23] ));
 sg13g2_nor3_1 _2662_ (.A(_1695_),
    .B(_1696_),
    .C(_1707_),
    .Y(_1708_));
 sg13g2_o21ai_1 _2663_ (.B1(\collatz.iter[26] ),
    .Y(_1709_),
    .A1(\collatz.iter[27] ),
    .A2(net710));
 sg13g2_nand2b_1 _2664_ (.Y(_1710_),
    .B(_1709_),
    .A_N(_1708_));
 sg13g2_xnor2_1 _2665_ (.Y(_1711_),
    .A(\collatz.iter[14] ),
    .B(\collatz.iter[13] ));
 sg13g2_xnor2_1 _2666_ (.Y(_1712_),
    .A(\collatz.iter[15] ),
    .B(\collatz.iter[14] ));
 sg13g2_nor2_1 _2667_ (.A(_1711_),
    .B(_1712_),
    .Y(_1713_));
 sg13g2_xor2_1 _2668_ (.B(\collatz.iter[11] ),
    .A(\collatz.iter[12] ),
    .X(_1714_));
 sg13g2_xor2_1 _2669_ (.B(\collatz.iter[12] ),
    .A(\collatz.iter[13] ),
    .X(_1715_));
 sg13g2_nand3_1 _2670_ (.B(_1714_),
    .C(_1715_),
    .A(_1713_),
    .Y(_1716_));
 sg13g2_a21oi_1 _2671_ (.A1(_1408_),
    .A2(_1410_),
    .Y(_1717_),
    .B1(_1409_));
 sg13g2_o21ai_1 _2672_ (.B1(\collatz.iter[12] ),
    .Y(_1718_),
    .A1(\collatz.iter[13] ),
    .A2(\collatz.iter[11] ));
 sg13g2_nor3_1 _2673_ (.A(_1711_),
    .B(_1712_),
    .C(_1718_),
    .Y(_1719_));
 sg13g2_nor2_1 _2674_ (.A(_1717_),
    .B(_1719_),
    .Y(_1720_));
 sg13g2_nand2_2 _2675_ (.Y(_1721_),
    .A(_1716_),
    .B(_1720_));
 sg13g2_o21ai_1 _2676_ (.B1(net756),
    .Y(_1722_),
    .A1(\collatz.iter[1] ),
    .A2(\collatz.iter[2] ));
 sg13g2_o21ai_1 _2677_ (.B1(\collatz.iter[2] ),
    .Y(_1723_),
    .A1(\collatz.iter[1] ),
    .A2(net711));
 sg13g2_o21ai_1 _2678_ (.B1(_1723_),
    .Y(_1724_),
    .A1(_1429_),
    .A2(_1722_));
 sg13g2_xnor2_1 _2679_ (.Y(_1725_),
    .A(\collatz.iter[6] ),
    .B(\collatz.iter[5] ));
 sg13g2_xnor2_1 _2680_ (.Y(_1726_),
    .A(\collatz.iter[7] ),
    .B(\collatz.iter[6] ));
 sg13g2_nor2_1 _2681_ (.A(_1725_),
    .B(_1726_),
    .Y(_1727_));
 sg13g2_xnor2_1 _2682_ (.Y(_1728_),
    .A(\collatz.iter[5] ),
    .B(\collatz.iter[4] ));
 sg13g2_xnor2_1 _2683_ (.Y(_1729_),
    .A(\collatz.iter[4] ),
    .B(\collatz.iter[3] ));
 sg13g2_nor4_1 _2684_ (.A(_1725_),
    .B(_1726_),
    .C(_1728_),
    .D(_1729_),
    .Y(_1730_));
 sg13g2_o21ai_1 _2685_ (.B1(\collatz.iter[4] ),
    .Y(_1731_),
    .A1(\collatz.iter[5] ),
    .A2(net711));
 sg13g2_inv_1 _2686_ (.Y(_1732_),
    .A(_1731_));
 sg13g2_o21ai_1 _2687_ (.B1(\collatz.iter[6] ),
    .Y(_1733_),
    .A1(\collatz.iter[7] ),
    .A2(\collatz.iter[5] ));
 sg13g2_inv_1 _2688_ (.Y(_1734_),
    .A(_1733_));
 sg13g2_a221oi_1 _2689_ (.B2(_1727_),
    .C1(_1734_),
    .B1(_1732_),
    .A1(_1724_),
    .Y(_1735_),
    .A2(_1730_));
 sg13g2_and2_1 _2690_ (.A(\collatz.iter[10] ),
    .B(\collatz.iter[9] ),
    .X(_1736_));
 sg13g2_xnor2_1 _2691_ (.Y(_1737_),
    .A(\collatz.iter[10] ),
    .B(\collatz.iter[9] ));
 sg13g2_xnor2_1 _2692_ (.Y(_1738_),
    .A(\collatz.iter[11] ),
    .B(\collatz.iter[10] ));
 sg13g2_nor2_1 _2693_ (.A(_1737_),
    .B(_1738_),
    .Y(_1739_));
 sg13g2_xnor2_1 _2694_ (.Y(_1740_),
    .A(\collatz.iter[8] ),
    .B(\collatz.iter[7] ));
 sg13g2_inv_1 _2695_ (.Y(_1741_),
    .A(_1740_));
 sg13g2_xor2_1 _2696_ (.B(\collatz.iter[8] ),
    .A(\collatz.iter[9] ),
    .X(_1742_));
 sg13g2_nand3_1 _2697_ (.B(_1741_),
    .C(_1742_),
    .A(_1739_),
    .Y(_1743_));
 sg13g2_nor2_1 _2698_ (.A(_1735_),
    .B(_1743_),
    .Y(_1744_));
 sg13g2_o21ai_1 _2699_ (.B1(\collatz.iter[8] ),
    .Y(_1745_),
    .A1(\collatz.iter[9] ),
    .A2(\collatz.iter[7] ));
 sg13g2_nor3_1 _2700_ (.A(_1737_),
    .B(_1738_),
    .C(_1745_),
    .Y(_1746_));
 sg13g2_a21o_1 _2701_ (.A2(\collatz.iter[10] ),
    .A1(\collatz.iter[11] ),
    .B1(_1736_),
    .X(_1747_));
 sg13g2_or2_1 _2702_ (.X(_1748_),
    .B(_1747_),
    .A(_1746_));
 sg13g2_nor4_1 _2703_ (.A(_1717_),
    .B(_1719_),
    .C(_1746_),
    .D(_1747_),
    .Y(_1749_));
 sg13g2_o21ai_1 _2704_ (.B1(_1749_),
    .Y(_1750_),
    .A1(_1735_),
    .A2(_1743_));
 sg13g2_and2_1 _2705_ (.A(_1721_),
    .B(_1750_),
    .X(_1751_));
 sg13g2_nand2_1 _2706_ (.Y(_1752_),
    .A(_1721_),
    .B(_1750_));
 sg13g2_and2_1 _2707_ (.A(\collatz.iter[22] ),
    .B(\collatz.iter[21] ),
    .X(_1753_));
 sg13g2_xor2_1 _2708_ (.B(\collatz.iter[21] ),
    .A(\collatz.iter[22] ),
    .X(_1754_));
 sg13g2_xor2_1 _2709_ (.B(\collatz.iter[22] ),
    .A(\collatz.iter[23] ),
    .X(_1755_));
 sg13g2_nand2_1 _2710_ (.Y(_1756_),
    .A(_1754_),
    .B(_1755_));
 sg13g2_nand2_1 _2711_ (.Y(_1757_),
    .A(\collatz.iter[20] ),
    .B(\collatz.iter[19] ));
 sg13g2_xor2_1 _2712_ (.B(\collatz.iter[19] ),
    .A(\collatz.iter[20] ),
    .X(_1758_));
 sg13g2_xor2_1 _2713_ (.B(\collatz.iter[20] ),
    .A(\collatz.iter[21] ),
    .X(_1759_));
 sg13g2_nand4_1 _2714_ (.B(_1755_),
    .C(_1758_),
    .A(_1754_),
    .Y(_1760_),
    .D(_1759_));
 sg13g2_and2_1 _2715_ (.A(\collatz.iter[18] ),
    .B(\collatz.iter[17] ),
    .X(_1761_));
 sg13g2_xor2_1 _2716_ (.B(\collatz.iter[17] ),
    .A(\collatz.iter[18] ),
    .X(_1762_));
 sg13g2_xor2_1 _2717_ (.B(\collatz.iter[18] ),
    .A(\collatz.iter[19] ),
    .X(_1763_));
 sg13g2_xor2_1 _2718_ (.B(\collatz.iter[15] ),
    .A(\collatz.iter[16] ),
    .X(_1764_));
 sg13g2_xor2_1 _2719_ (.B(\collatz.iter[16] ),
    .A(\collatz.iter[17] ),
    .X(_1765_));
 sg13g2_nand4_1 _2720_ (.B(_1763_),
    .C(_1764_),
    .A(_1762_),
    .Y(_1766_),
    .D(_1765_));
 sg13g2_nor2_1 _2721_ (.A(_1760_),
    .B(_1766_),
    .Y(_1767_));
 sg13g2_o21ai_1 _2722_ (.B1(\collatz.iter[16] ),
    .Y(_1768_),
    .A1(\collatz.iter[17] ),
    .A2(\collatz.iter[15] ));
 sg13g2_nand3b_1 _2723_ (.B(_1763_),
    .C(_1762_),
    .Y(_1769_),
    .A_N(_1768_));
 sg13g2_o21ai_1 _2724_ (.B1(\collatz.iter[18] ),
    .Y(_1770_),
    .A1(\collatz.iter[19] ),
    .A2(\collatz.iter[17] ));
 sg13g2_a21oi_1 _2725_ (.A1(_1769_),
    .A2(_1770_),
    .Y(_1771_),
    .B1(_1760_));
 sg13g2_o21ai_1 _2726_ (.B1(\collatz.iter[22] ),
    .Y(_1772_),
    .A1(\collatz.iter[23] ),
    .A2(\collatz.iter[21] ));
 sg13g2_o21ai_1 _2727_ (.B1(\collatz.iter[20] ),
    .Y(_1773_),
    .A1(\collatz.iter[21] ),
    .A2(\collatz.iter[19] ));
 sg13g2_o21ai_1 _2728_ (.B1(_1772_),
    .Y(_1774_),
    .A1(_1756_),
    .A2(_1773_));
 sg13g2_or2_1 _2729_ (.X(_1775_),
    .B(_1774_),
    .A(_1771_));
 sg13g2_a221oi_1 _2730_ (.B2(_1702_),
    .C1(_1706_),
    .B1(_1775_),
    .A1(_1692_),
    .Y(_1776_),
    .A2(_1710_));
 sg13g2_nand4_1 _2731_ (.B(_1721_),
    .C(_1750_),
    .A(_1702_),
    .Y(_1777_),
    .D(_1767_));
 sg13g2_nand2_2 _2732_ (.Y(_1778_),
    .A(_1776_),
    .B(_1777_));
 sg13g2_and2_1 _2733_ (.A(\collatz.iter[58] ),
    .B(\collatz.iter[57] ),
    .X(_1779_));
 sg13g2_xor2_1 _2734_ (.B(\collatz.iter[57] ),
    .A(\collatz.iter[58] ),
    .X(_1780_));
 sg13g2_xor2_1 _2735_ (.B(\collatz.iter[58] ),
    .A(\collatz.iter[59] ),
    .X(_1781_));
 sg13g2_nand2_1 _2736_ (.Y(_1782_),
    .A(_1780_),
    .B(_1781_));
 sg13g2_xor2_1 _2737_ (.B(\collatz.iter[56] ),
    .A(\collatz.iter[57] ),
    .X(_1783_));
 sg13g2_nand2_1 _2738_ (.Y(_1784_),
    .A(\collatz.iter[56] ),
    .B(\collatz.iter[55] ));
 sg13g2_xor2_1 _2739_ (.B(\collatz.iter[55] ),
    .A(\collatz.iter[56] ),
    .X(_1785_));
 sg13g2_and4_1 _2740_ (.A(_1780_),
    .B(_1781_),
    .C(_1783_),
    .D(_1785_),
    .X(_1786_));
 sg13g2_nand2_1 _2741_ (.Y(_1787_),
    .A(\collatz.iter[60] ),
    .B(\collatz.iter[59] ));
 sg13g2_xnor2_1 _2742_ (.Y(_1788_),
    .A(\collatz.iter[60] ),
    .B(\collatz.iter[59] ));
 sg13g2_xnor2_1 _2743_ (.Y(_1789_),
    .A(net702),
    .B(\collatz.iter[60] ));
 sg13g2_nor2_1 _2744_ (.A(_1788_),
    .B(_1789_),
    .Y(_1790_));
 sg13g2_and2_1 _2745_ (.A(\collatz.iter[62] ),
    .B(net702),
    .X(_1791_));
 sg13g2_xor2_1 _2746_ (.B(net702),
    .A(\collatz.iter[62] ),
    .X(_1792_));
 sg13g2_xor2_1 _2747_ (.B(\collatz.iter[62] ),
    .A(\collatz.iter[63] ),
    .X(_1793_));
 sg13g2_nand2_1 _2748_ (.Y(_1794_),
    .A(_1792_),
    .B(_1793_));
 sg13g2_nand4_1 _2749_ (.B(_1790_),
    .C(_1792_),
    .A(_1786_),
    .Y(_1795_),
    .D(_1793_));
 sg13g2_and2_1 _2750_ (.A(\collatz.iter[54] ),
    .B(net703),
    .X(_1796_));
 sg13g2_xor2_1 _2751_ (.B(net703),
    .A(\collatz.iter[54] ),
    .X(_1797_));
 sg13g2_xor2_1 _2752_ (.B(\collatz.iter[54] ),
    .A(\collatz.iter[55] ),
    .X(_1798_));
 sg13g2_nand2_1 _2753_ (.Y(_1799_),
    .A(_1797_),
    .B(_1798_));
 sg13g2_xor2_1 _2754_ (.B(net704),
    .A(net703),
    .X(_1800_));
 sg13g2_nand2_1 _2755_ (.Y(_1801_),
    .A(net704),
    .B(net705));
 sg13g2_xor2_1 _2756_ (.B(net705),
    .A(net704),
    .X(_1802_));
 sg13g2_xnor2_1 _2757_ (.Y(_1803_),
    .A(net704),
    .B(net705));
 sg13g2_nand4_1 _2758_ (.B(_1798_),
    .C(_1800_),
    .A(_1797_),
    .Y(_1804_),
    .D(_1802_));
 sg13g2_and2_1 _2759_ (.A(\collatz.iter[50] ),
    .B(\collatz.iter[49] ),
    .X(_1805_));
 sg13g2_xor2_1 _2760_ (.B(\collatz.iter[49] ),
    .A(\collatz.iter[50] ),
    .X(_1806_));
 sg13g2_xor2_1 _2761_ (.B(\collatz.iter[50] ),
    .A(net705),
    .X(_1807_));
 sg13g2_nand2_1 _2762_ (.Y(_1808_),
    .A(\collatz.iter[48] ),
    .B(\collatz.iter[47] ));
 sg13g2_xor2_1 _2763_ (.B(\collatz.iter[47] ),
    .A(\collatz.iter[48] ),
    .X(_1809_));
 sg13g2_xor2_1 _2764_ (.B(\collatz.iter[48] ),
    .A(\collatz.iter[49] ),
    .X(_1810_));
 sg13g2_nand4_1 _2765_ (.B(_1807_),
    .C(_1809_),
    .A(_1806_),
    .Y(_1811_),
    .D(_1810_));
 sg13g2_or2_1 _2766_ (.X(_1812_),
    .B(_1811_),
    .A(_1804_));
 sg13g2_or2_1 _2767_ (.X(_1813_),
    .B(_1812_),
    .A(_1795_));
 sg13g2_and2_1 _2768_ (.A(\collatz.iter[46] ),
    .B(net706),
    .X(_1814_));
 sg13g2_xor2_1 _2769_ (.B(net706),
    .A(\collatz.iter[46] ),
    .X(_1815_));
 sg13g2_xor2_1 _2770_ (.B(\collatz.iter[46] ),
    .A(\collatz.iter[47] ),
    .X(_1816_));
 sg13g2_nand2_1 _2771_ (.Y(_1817_),
    .A(_1815_),
    .B(_1816_));
 sg13g2_xor2_1 _2772_ (.B(\collatz.iter[44] ),
    .A(net706),
    .X(_1818_));
 sg13g2_nand2_1 _2773_ (.Y(_1819_),
    .A(\collatz.iter[44] ),
    .B(\collatz.iter[43] ));
 sg13g2_xor2_1 _2774_ (.B(\collatz.iter[43] ),
    .A(\collatz.iter[44] ),
    .X(_1820_));
 sg13g2_nand4_1 _2775_ (.B(_1816_),
    .C(_1818_),
    .A(_1815_),
    .Y(_1821_),
    .D(_1820_));
 sg13g2_and2_1 _2776_ (.A(\collatz.iter[42] ),
    .B(\collatz.iter[41] ),
    .X(_1822_));
 sg13g2_xor2_1 _2777_ (.B(net707),
    .A(\collatz.iter[42] ),
    .X(_1823_));
 sg13g2_xor2_1 _2778_ (.B(\collatz.iter[42] ),
    .A(\collatz.iter[43] ),
    .X(_1824_));
 sg13g2_nand2_1 _2779_ (.Y(_1825_),
    .A(\collatz.iter[40] ),
    .B(\collatz.iter[39] ));
 sg13g2_xor2_1 _2780_ (.B(\collatz.iter[39] ),
    .A(\collatz.iter[40] ),
    .X(_1826_));
 sg13g2_xor2_1 _2781_ (.B(\collatz.iter[40] ),
    .A(net707),
    .X(_1827_));
 sg13g2_nand4_1 _2782_ (.B(_1824_),
    .C(_1826_),
    .A(_1823_),
    .Y(_1828_),
    .D(_1827_));
 sg13g2_nor2_1 _2783_ (.A(_1821_),
    .B(_1828_),
    .Y(_1829_));
 sg13g2_and2_1 _2784_ (.A(\collatz.iter[38] ),
    .B(net708),
    .X(_1830_));
 sg13g2_xor2_1 _2785_ (.B(net708),
    .A(\collatz.iter[38] ),
    .X(_1831_));
 sg13g2_xor2_1 _2786_ (.B(\collatz.iter[38] ),
    .A(\collatz.iter[39] ),
    .X(_1832_));
 sg13g2_nand2_1 _2787_ (.Y(_1833_),
    .A(_1831_),
    .B(_1832_));
 sg13g2_nand2_1 _2788_ (.Y(_1834_),
    .A(\collatz.iter[36] ),
    .B(\collatz.iter[35] ));
 sg13g2_xor2_1 _2789_ (.B(\collatz.iter[35] ),
    .A(\collatz.iter[36] ),
    .X(_1835_));
 sg13g2_xor2_1 _2790_ (.B(\collatz.iter[36] ),
    .A(net708),
    .X(_1836_));
 sg13g2_nand4_1 _2791_ (.B(_1832_),
    .C(_1835_),
    .A(_1831_),
    .Y(_1837_),
    .D(_1836_));
 sg13g2_and2_1 _2792_ (.A(\collatz.iter[34] ),
    .B(net709),
    .X(_1838_));
 sg13g2_xor2_1 _2793_ (.B(net709),
    .A(\collatz.iter[34] ),
    .X(_1839_));
 sg13g2_xor2_1 _2794_ (.B(\collatz.iter[34] ),
    .A(\collatz.iter[35] ),
    .X(_1840_));
 sg13g2_nand2_1 _2795_ (.Y(_1841_),
    .A(_1839_),
    .B(_1840_));
 sg13g2_nand2_1 _2796_ (.Y(_1842_),
    .A(\collatz.iter[32] ),
    .B(\collatz.iter[31] ));
 sg13g2_xnor2_1 _2797_ (.Y(_1843_),
    .A(\collatz.iter[32] ),
    .B(\collatz.iter[31] ));
 sg13g2_xnor2_1 _2798_ (.Y(_1844_),
    .A(net709),
    .B(\collatz.iter[32] ));
 sg13g2_nor3_1 _2799_ (.A(_1841_),
    .B(_1843_),
    .C(_1844_),
    .Y(_1845_));
 sg13g2_nor4_1 _2800_ (.A(_1837_),
    .B(_1841_),
    .C(_1843_),
    .D(_1844_),
    .Y(_1846_));
 sg13g2_and2_1 _2801_ (.A(_1829_),
    .B(_1846_),
    .X(_1847_));
 sg13g2_nand2b_1 _2802_ (.Y(_1848_),
    .B(_1847_),
    .A_N(_1813_));
 sg13g2_a21oi_2 _2803_ (.B1(_1848_),
    .Y(_1849_),
    .A2(_1777_),
    .A1(_1776_));
 sg13g2_o21ai_1 _2804_ (.B1(\collatz.iter[32] ),
    .Y(_1850_),
    .A1(net709),
    .A2(\collatz.iter[31] ));
 sg13g2_nand3b_1 _2805_ (.B(_1840_),
    .C(_1839_),
    .Y(_1851_),
    .A_N(_1850_));
 sg13g2_o21ai_1 _2806_ (.B1(\collatz.iter[34] ),
    .Y(_1852_),
    .A1(\collatz.iter[35] ),
    .A2(net709));
 sg13g2_nand2_1 _2807_ (.Y(_1853_),
    .A(_1851_),
    .B(_1852_));
 sg13g2_a21oi_1 _2808_ (.A1(_1851_),
    .A2(_1852_),
    .Y(_1854_),
    .B1(_1837_));
 sg13g2_o21ai_1 _2809_ (.B1(\collatz.iter[38] ),
    .Y(_1855_),
    .A1(\collatz.iter[39] ),
    .A2(net708));
 sg13g2_o21ai_1 _2810_ (.B1(\collatz.iter[36] ),
    .Y(_1856_),
    .A1(net708),
    .A2(\collatz.iter[35] ));
 sg13g2_o21ai_1 _2811_ (.B1(_1855_),
    .Y(_1857_),
    .A1(_1833_),
    .A2(_1856_));
 sg13g2_o21ai_1 _2812_ (.B1(_1829_),
    .Y(_1858_),
    .A1(_1854_),
    .A2(_1857_));
 sg13g2_o21ai_1 _2813_ (.B1(\collatz.iter[44] ),
    .Y(_1859_),
    .A1(net706),
    .A2(\collatz.iter[43] ));
 sg13g2_o21ai_1 _2814_ (.B1(\collatz.iter[46] ),
    .Y(_1860_),
    .A1(\collatz.iter[47] ),
    .A2(net706));
 sg13g2_o21ai_1 _2815_ (.B1(_1860_),
    .Y(_1861_),
    .A1(_1817_),
    .A2(_1859_));
 sg13g2_o21ai_1 _2816_ (.B1(\collatz.iter[40] ),
    .Y(_1862_),
    .A1(net707),
    .A2(\collatz.iter[39] ));
 sg13g2_nand3b_1 _2817_ (.B(_1824_),
    .C(_1823_),
    .Y(_1863_),
    .A_N(_1862_));
 sg13g2_o21ai_1 _2818_ (.B1(\collatz.iter[42] ),
    .Y(_1864_),
    .A1(\collatz.iter[43] ),
    .A2(net707));
 sg13g2_and2_1 _2819_ (.A(_1863_),
    .B(_1864_),
    .X(_1865_));
 sg13g2_a21oi_1 _2820_ (.A1(_1863_),
    .A2(_1864_),
    .Y(_1866_),
    .B1(_1821_));
 sg13g2_nor2_1 _2821_ (.A(_1861_),
    .B(_1866_),
    .Y(_1867_));
 sg13g2_nand2_1 _2822_ (.Y(_1868_),
    .A(_1858_),
    .B(_1867_));
 sg13g2_a21oi_2 _2823_ (.B1(_1813_),
    .Y(_1869_),
    .A2(_1867_),
    .A1(_1858_));
 sg13g2_o21ai_1 _2824_ (.B1(\collatz.iter[48] ),
    .Y(_1870_),
    .A1(\collatz.iter[49] ),
    .A2(\collatz.iter[47] ));
 sg13g2_nand3b_1 _2825_ (.B(_1807_),
    .C(_1806_),
    .Y(_1871_),
    .A_N(_1870_));
 sg13g2_o21ai_1 _2826_ (.B1(\collatz.iter[50] ),
    .Y(_1872_),
    .A1(net705),
    .A2(\collatz.iter[49] ));
 sg13g2_and2_1 _2827_ (.A(_1871_),
    .B(_1872_),
    .X(_1873_));
 sg13g2_a21oi_1 _2828_ (.A1(_1871_),
    .A2(_1872_),
    .Y(_1874_),
    .B1(_1804_));
 sg13g2_o21ai_1 _2829_ (.B1(\collatz.iter[54] ),
    .Y(_1875_),
    .A1(\collatz.iter[55] ),
    .A2(net703));
 sg13g2_o21ai_1 _2830_ (.B1(net704),
    .Y(_1876_),
    .A1(net703),
    .A2(net705));
 sg13g2_o21ai_1 _2831_ (.B1(_1875_),
    .Y(_1877_),
    .A1(_1799_),
    .A2(_1876_));
 sg13g2_nor2_2 _2832_ (.A(_1874_),
    .B(_1877_),
    .Y(_1878_));
 sg13g2_o21ai_1 _2833_ (.B1(\collatz.iter[62] ),
    .Y(_1879_),
    .A1(\collatz.iter[63] ),
    .A2(net702));
 sg13g2_o21ai_1 _2834_ (.B1(\collatz.iter[60] ),
    .Y(_1880_),
    .A1(net702),
    .A2(\collatz.iter[59] ));
 sg13g2_o21ai_1 _2835_ (.B1(\collatz.iter[56] ),
    .Y(_1881_),
    .A1(\collatz.iter[57] ),
    .A2(\collatz.iter[55] ));
 sg13g2_o21ai_1 _2836_ (.B1(\collatz.iter[58] ),
    .Y(_1882_),
    .A1(\collatz.iter[59] ),
    .A2(\collatz.iter[57] ));
 sg13g2_o21ai_1 _2837_ (.B1(_1882_),
    .Y(_1883_),
    .A1(_1782_),
    .A2(_1881_));
 sg13g2_nand2_1 _2838_ (.Y(_1884_),
    .A(_1790_),
    .B(_1883_));
 sg13g2_a21oi_1 _2839_ (.A1(_1880_),
    .A2(_1884_),
    .Y(_1885_),
    .B1(_1794_));
 sg13g2_o21ai_1 _2840_ (.B1(_1879_),
    .Y(_1886_),
    .A1(_1795_),
    .A2(_1878_));
 sg13g2_or3_2 _2841_ (.A(_1869_),
    .B(_1885_),
    .C(_1886_),
    .X(_1887_));
 sg13g2_nor2_2 _2842_ (.A(_1849_),
    .B(_1887_),
    .Y(_1888_));
 sg13g2_xor2_1 _2843_ (.B(\collatz.iter[63] ),
    .A(\collatz.iter[64] ),
    .X(_1889_));
 sg13g2_xor2_1 _2844_ (.B(\collatz.iter[64] ),
    .A(\collatz.iter[65] ),
    .X(_1890_));
 sg13g2_nand4_1 _2845_ (.B(_1663_),
    .C(_1889_),
    .A(_1662_),
    .Y(_1891_),
    .D(_1890_));
 sg13g2_nor2_1 _2846_ (.A(_1660_),
    .B(_1891_),
    .Y(_1892_));
 sg13g2_nand2_1 _2847_ (.Y(_1893_),
    .A(_1653_),
    .B(_1892_));
 sg13g2_and4_2 _2848_ (.A(_1615_),
    .B(_1653_),
    .C(_1684_),
    .D(_1892_),
    .X(_1894_));
 sg13g2_o21ai_1 _2849_ (.B1(_1894_),
    .Y(_1895_),
    .A1(_1849_),
    .A2(_1887_));
 sg13g2_nand2b_2 _2850_ (.Y(_1896_),
    .B(_1895_),
    .A_N(_1686_));
 sg13g2_a221oi_1 _2851_ (.B2(_1896_),
    .C1(_1583_),
    .B1(_1590_),
    .A1(_1556_),
    .Y(_1897_),
    .A2(_1580_));
 sg13g2_o21ai_1 _2852_ (.B1(\collatz.iter[112] ),
    .Y(_1898_),
    .A1(net698),
    .A2(\collatz.iter[111] ));
 sg13g2_inv_1 _2853_ (.Y(_1899_),
    .A(_1898_));
 sg13g2_o21ai_1 _2854_ (.B1(_1898_),
    .Y(_1900_),
    .A1(_1533_),
    .A2(_1897_));
 sg13g2_o21ai_1 _2855_ (.B1(_1532_),
    .Y(_1901_),
    .A1(_1533_),
    .A2(_1897_));
 sg13g2_o21ai_1 _2856_ (.B1(_1900_),
    .Y(_1902_),
    .A1(net698),
    .A2(\collatz.iter[112] ));
 sg13g2_xnor2_1 _2857_ (.Y(_1903_),
    .A(\collatz.iter[114] ),
    .B(net698));
 sg13g2_or2_1 _2858_ (.X(_1904_),
    .B(_1903_),
    .A(_1902_));
 sg13g2_nand2_1 _2859_ (.Y(_1905_),
    .A(_1528_),
    .B(_1904_));
 sg13g2_xnor2_1 _2860_ (.Y(_1906_),
    .A(\collatz.iter[115] ),
    .B(\collatz.iter[114] ));
 sg13g2_a21oi_1 _2861_ (.A1(_1530_),
    .A2(_1904_),
    .Y(_1907_),
    .B1(_1438_));
 sg13g2_nand2b_1 _2862_ (.Y(_1908_),
    .B(_1907_),
    .A_N(_1527_));
 sg13g2_a21oi_1 _2863_ (.A1(_1525_),
    .A2(_1908_),
    .Y(_1909_),
    .B1(_1454_));
 sg13g2_a21oi_1 _2864_ (.A1(_1523_),
    .A2(_1909_),
    .Y(_1910_),
    .B1(_1522_));
 sg13g2_xor2_1 _2865_ (.B(_1910_),
    .A(_1521_),
    .X(_1911_));
 sg13g2_o21ai_1 _2866_ (.B1(net760),
    .Y(_1912_),
    .A1(\collatz.iter[120] ),
    .A2(net717));
 sg13g2_a21o_1 _2867_ (.A2(_1911_),
    .A1(net713),
    .B1(_1912_),
    .X(_1913_));
 sg13g2_a21oi_1 _2868_ (.A1(_1520_),
    .A2(_1913_),
    .Y(_0011_),
    .B1(net805));
 sg13g2_and3_1 _2869_ (.X(_1914_),
    .A(net1),
    .B(net826),
    .C(net829));
 sg13g2_a21oi_2 _2870_ (.B1(net650),
    .Y(_1915_),
    .A2(net804),
    .A1(net657));
 sg13g2_and2_1 _2871_ (.A(net844),
    .B(net804),
    .X(_1916_));
 sg13g2_a22oi_1 _2872_ (.Y(_1917_),
    .B1(_1916_),
    .B2(net655),
    .A2(_1915_),
    .A1(\collatz.iter[120] ));
 sg13g2_or2_1 _2873_ (.X(_1918_),
    .B(_1917_),
    .A(net761));
 sg13g2_nand2_1 _2874_ (.Y(_1919_),
    .A(\collatz.iter[120] ),
    .B(\collatz.iter[119] ));
 sg13g2_xor2_1 _2875_ (.B(\collatz.iter[119] ),
    .A(\collatz.iter[120] ),
    .X(_1920_));
 sg13g2_nand2_1 _2876_ (.Y(_1921_),
    .A(_1521_),
    .B(_1523_));
 sg13g2_xnor2_1 _2877_ (.Y(_1922_),
    .A(\collatz.iter[117] ),
    .B(\collatz.iter[116] ));
 sg13g2_nor2_1 _2878_ (.A(_1527_),
    .B(_1922_),
    .Y(_1923_));
 sg13g2_nor4_2 _2879_ (.A(_1527_),
    .B(_1903_),
    .C(_1906_),
    .Y(_1924_),
    .D(_1922_));
 sg13g2_inv_1 _2880_ (.Y(_1925_),
    .A(_1924_));
 sg13g2_a221oi_1 _2881_ (.B2(_1899_),
    .C1(_1526_),
    .B1(_1924_),
    .A1(_1531_),
    .Y(_1926_),
    .A2(_1923_));
 sg13g2_o21ai_1 _2882_ (.B1(\collatz.iter[118] ),
    .Y(_1927_),
    .A1(\collatz.iter[119] ),
    .A2(\collatz.iter[117] ));
 sg13g2_o21ai_1 _2883_ (.B1(_1927_),
    .Y(_1928_),
    .A1(_1921_),
    .A2(_1926_));
 sg13g2_inv_1 _2884_ (.Y(_1929_),
    .A(_1928_));
 sg13g2_xor2_1 _2885_ (.B(\collatz.iter[112] ),
    .A(net698),
    .X(_1930_));
 sg13g2_nand2b_1 _2886_ (.Y(_1931_),
    .B(_1930_),
    .A_N(_1533_));
 sg13g2_nor3_2 _2887_ (.A(_1921_),
    .B(_1925_),
    .C(_1931_),
    .Y(_1932_));
 sg13g2_inv_1 _2888_ (.Y(_1933_),
    .A(_1932_));
 sg13g2_o21ai_1 _2889_ (.B1(_1929_),
    .Y(_1934_),
    .A1(_1897_),
    .A2(_1933_));
 sg13g2_nand2_1 _2890_ (.Y(_1935_),
    .A(_1920_),
    .B(_1934_));
 sg13g2_xnor2_1 _2891_ (.Y(_1936_),
    .A(_1920_),
    .B(_1934_));
 sg13g2_o21ai_1 _2892_ (.B1(net761),
    .Y(_1937_),
    .A1(\collatz.iter[121] ),
    .A2(net719));
 sg13g2_a21o_1 _2893_ (.A2(_1936_),
    .A1(net719),
    .B1(_1937_),
    .X(_1938_));
 sg13g2_a21oi_1 _2894_ (.A1(_1918_),
    .A2(_1938_),
    .Y(_0012_),
    .B1(net807));
 sg13g2_and2_1 _2895_ (.A(net842),
    .B(net804),
    .X(_1939_));
 sg13g2_a22oi_1 _2896_ (.Y(_1940_),
    .B1(_1939_),
    .B2(net655),
    .A2(_1915_),
    .A1(\collatz.iter[121] ));
 sg13g2_or2_1 _2897_ (.X(_1941_),
    .B(_1940_),
    .A(net761));
 sg13g2_xor2_1 _2898_ (.B(\collatz.iter[120] ),
    .A(\collatz.iter[121] ),
    .X(_1942_));
 sg13g2_nand2_1 _2899_ (.Y(_1943_),
    .A(_1919_),
    .B(_1935_));
 sg13g2_xnor2_1 _2900_ (.Y(_1944_),
    .A(_1942_),
    .B(_1943_));
 sg13g2_a21oi_1 _2901_ (.A1(net719),
    .A2(_1944_),
    .Y(_1945_),
    .B1(net685));
 sg13g2_o21ai_1 _2902_ (.B1(_1945_),
    .Y(_1946_),
    .A1(net309),
    .A2(net717));
 sg13g2_a21oi_1 _2903_ (.A1(_1941_),
    .A2(_1946_),
    .Y(_0013_),
    .B1(net807));
 sg13g2_and2_1 _2904_ (.A(net840),
    .B(net804),
    .X(_1947_));
 sg13g2_a22oi_1 _2905_ (.Y(_1948_),
    .B1(_1947_),
    .B2(net655),
    .A2(_1915_),
    .A1(net335));
 sg13g2_or2_1 _2906_ (.X(_1949_),
    .B(_1948_),
    .A(net761));
 sg13g2_and2_1 _2907_ (.A(\collatz.iter[122] ),
    .B(\collatz.iter[121] ),
    .X(_1950_));
 sg13g2_xor2_1 _2908_ (.B(\collatz.iter[121] ),
    .A(\collatz.iter[122] ),
    .X(_1951_));
 sg13g2_o21ai_1 _2909_ (.B1(\collatz.iter[120] ),
    .Y(_1952_),
    .A1(\collatz.iter[121] ),
    .A2(\collatz.iter[119] ));
 sg13g2_a21oi_1 _2910_ (.A1(_1935_),
    .A2(_1952_),
    .Y(_1953_),
    .B1(_1450_));
 sg13g2_xnor2_1 _2911_ (.Y(_1954_),
    .A(_1951_),
    .B(_1953_));
 sg13g2_o21ai_1 _2912_ (.B1(net761),
    .Y(_1955_),
    .A1(\collatz.iter[123] ),
    .A2(net717));
 sg13g2_a21o_1 _2913_ (.A2(_1954_),
    .A1(net717),
    .B1(_1955_),
    .X(_1956_));
 sg13g2_a21oi_1 _2914_ (.A1(_1949_),
    .A2(_1956_),
    .Y(_0014_),
    .B1(net807));
 sg13g2_and2_1 _2915_ (.A(net838),
    .B(net804),
    .X(_1957_));
 sg13g2_a22oi_1 _2916_ (.Y(_1958_),
    .B1(_1957_),
    .B2(net655),
    .A2(_1915_),
    .A1(\collatz.iter[123] ));
 sg13g2_or2_1 _2917_ (.X(_1959_),
    .B(_1958_),
    .A(net761));
 sg13g2_xor2_1 _2918_ (.B(\collatz.iter[122] ),
    .A(\collatz.iter[123] ),
    .X(_1960_));
 sg13g2_a21oi_1 _2919_ (.A1(_1951_),
    .A2(_1953_),
    .Y(_1961_),
    .B1(_1950_));
 sg13g2_xor2_1 _2920_ (.B(_1961_),
    .A(_1960_),
    .X(_1962_));
 sg13g2_a21oi_1 _2921_ (.A1(net717),
    .A2(_1962_),
    .Y(_1963_),
    .B1(net685));
 sg13g2_o21ai_1 _2922_ (.B1(_1963_),
    .Y(_1964_),
    .A1(net304),
    .A2(net729));
 sg13g2_a21oi_1 _2923_ (.A1(_1959_),
    .A2(_1964_),
    .Y(_0015_),
    .B1(net807));
 sg13g2_and2_1 _2924_ (.A(net836),
    .B(_1914_),
    .X(_1965_));
 sg13g2_a22oi_1 _2925_ (.Y(_1966_),
    .B1(_1965_),
    .B2(_1516_),
    .A2(_1915_),
    .A1(net337));
 sg13g2_or2_1 _2926_ (.X(_1967_),
    .B(_1966_),
    .A(net760));
 sg13g2_nand2_1 _2927_ (.Y(_1968_),
    .A(\collatz.iter[124] ),
    .B(\collatz.iter[123] ));
 sg13g2_xnor2_1 _2928_ (.Y(_0196_),
    .A(\collatz.iter[124] ),
    .B(\collatz.iter[123] ));
 sg13g2_nand3b_1 _2929_ (.B(_1960_),
    .C(_1951_),
    .Y(_0197_),
    .A_N(_1952_));
 sg13g2_o21ai_1 _2930_ (.B1(\collatz.iter[122] ),
    .Y(_0198_),
    .A1(\collatz.iter[123] ),
    .A2(\collatz.iter[121] ));
 sg13g2_nand4_1 _2931_ (.B(_1942_),
    .C(_1951_),
    .A(_1920_),
    .Y(_0199_),
    .D(_1960_));
 sg13g2_nand2b_1 _2932_ (.Y(_0200_),
    .B(_1934_),
    .A_N(_0199_));
 sg13g2_and3_1 _2933_ (.X(_0201_),
    .A(_0197_),
    .B(_0198_),
    .C(_0200_));
 sg13g2_or2_1 _2934_ (.X(_0202_),
    .B(_0201_),
    .A(_0196_));
 sg13g2_xnor2_1 _2935_ (.Y(_0203_),
    .A(_0196_),
    .B(_0201_));
 sg13g2_o21ai_1 _2936_ (.B1(net768),
    .Y(_0204_),
    .A1(net803),
    .A2(net729));
 sg13g2_a21o_1 _2937_ (.A2(_0203_),
    .A1(net729),
    .B1(_0204_),
    .X(_0205_));
 sg13g2_a21oi_1 _2938_ (.A1(_1967_),
    .A2(_0205_),
    .Y(_0016_),
    .B1(net811));
 sg13g2_and2_1 _2939_ (.A(net834),
    .B(_1914_),
    .X(_0206_));
 sg13g2_a22oi_1 _2940_ (.Y(_0207_),
    .B1(_0206_),
    .B2(net657),
    .A2(_1915_),
    .A1(net803));
 sg13g2_or2_1 _2941_ (.X(_0208_),
    .B(_0207_),
    .A(net768));
 sg13g2_xnor2_1 _2942_ (.Y(_0209_),
    .A(net803),
    .B(\collatz.iter[124] ));
 sg13g2_nand2_1 _2943_ (.Y(_0210_),
    .A(_1968_),
    .B(_0202_));
 sg13g2_xor2_1 _2944_ (.B(_0210_),
    .A(_0209_),
    .X(_0211_));
 sg13g2_a21oi_1 _2945_ (.A1(net729),
    .A2(_0211_),
    .Y(_0212_),
    .B1(net688));
 sg13g2_o21ai_1 _2946_ (.B1(_0212_),
    .Y(_0213_),
    .A1(net298),
    .A2(net729));
 sg13g2_a21oi_1 _2947_ (.A1(_0208_),
    .A2(_0213_),
    .Y(_0017_),
    .B1(net811));
 sg13g2_and2_1 _2948_ (.A(net832),
    .B(net804),
    .X(_0214_));
 sg13g2_a22oi_1 _2949_ (.Y(_0215_),
    .B1(_0214_),
    .B2(net657),
    .A2(_1915_),
    .A1(net298));
 sg13g2_or2_1 _2950_ (.X(_0216_),
    .B(_0215_),
    .A(net768));
 sg13g2_and2_1 _2951_ (.A(\collatz.iter[126] ),
    .B(net803),
    .X(_0217_));
 sg13g2_xor2_1 _2952_ (.B(\collatz.iter[125] ),
    .A(\collatz.iter[126] ),
    .X(_0218_));
 sg13g2_o21ai_1 _2953_ (.B1(\collatz.iter[124] ),
    .Y(_0219_),
    .A1(net803),
    .A2(\collatz.iter[123] ));
 sg13g2_a21oi_1 _2954_ (.A1(_0202_),
    .A2(_0219_),
    .Y(_0220_),
    .B1(_1434_));
 sg13g2_xnor2_1 _2955_ (.Y(_0221_),
    .A(_0218_),
    .B(_0220_));
 sg13g2_o21ai_1 _2956_ (.B1(net768),
    .Y(_0222_),
    .A1(\collatz.iter[127] ),
    .A2(net731));
 sg13g2_a21o_1 _2957_ (.A2(_0221_),
    .A1(net729),
    .B1(_0222_),
    .X(_0223_));
 sg13g2_a21oi_1 _2958_ (.A1(_0216_),
    .A2(_0223_),
    .Y(_0018_),
    .B1(net811));
 sg13g2_and2_1 _2959_ (.A(net830),
    .B(net804),
    .X(_0224_));
 sg13g2_a22oi_1 _2960_ (.Y(_0225_),
    .B1(_0224_),
    .B2(net657),
    .A2(_1915_),
    .A1(\collatz.iter[127] ));
 sg13g2_or2_1 _2961_ (.X(_0226_),
    .B(_0225_),
    .A(net768));
 sg13g2_xor2_1 _2962_ (.B(\collatz.iter[126] ),
    .A(\collatz.iter[127] ),
    .X(_0227_));
 sg13g2_a21oi_1 _2963_ (.A1(_0218_),
    .A2(_0220_),
    .Y(_0228_),
    .B1(_0217_));
 sg13g2_xor2_1 _2964_ (.B(_0228_),
    .A(_0227_),
    .X(_0229_));
 sg13g2_a21oi_1 _2965_ (.A1(net729),
    .A2(_0229_),
    .Y(_0230_),
    .B1(net688));
 sg13g2_o21ai_1 _2966_ (.B1(_0230_),
    .Y(_0231_),
    .A1(net317),
    .A2(net732));
 sg13g2_a21oi_1 _2967_ (.A1(_0226_),
    .A2(_0231_),
    .Y(_0019_),
    .B1(net811));
 sg13g2_and2_1 _2968_ (.A(net7),
    .B(net4),
    .X(_0232_));
 sg13g2_and2_2 _2969_ (.A(_1512_),
    .B(_0232_),
    .X(_0233_));
 sg13g2_and2_2 _2970_ (.A(net691),
    .B(_0233_),
    .X(_0234_));
 sg13g2_nand2_1 _2971_ (.Y(_0235_),
    .A(_0218_),
    .B(_0227_));
 sg13g2_inv_1 _2972_ (.Y(_0236_),
    .A(_0235_));
 sg13g2_or2_1 _2973_ (.X(_0237_),
    .B(_0209_),
    .A(_0196_));
 sg13g2_nor3_2 _2974_ (.A(_0199_),
    .B(_0235_),
    .C(_0237_),
    .Y(_0238_));
 sg13g2_a21oi_1 _2975_ (.A1(_0197_),
    .A2(_0198_),
    .Y(_0239_),
    .B1(_0237_));
 sg13g2_nand2b_1 _2976_ (.Y(_0240_),
    .B(_0219_),
    .A_N(_0239_));
 sg13g2_o21ai_1 _2977_ (.B1(\collatz.iter[126] ),
    .Y(_0241_),
    .A1(\collatz.iter[127] ),
    .A2(net803));
 sg13g2_inv_1 _2978_ (.Y(_0242_),
    .A(_0241_));
 sg13g2_a221oi_1 _2979_ (.B2(_0236_),
    .C1(_0242_),
    .B1(_0240_),
    .A1(_1928_),
    .Y(_0243_),
    .A2(_0238_));
 sg13g2_nand2_1 _2980_ (.Y(_0244_),
    .A(_1932_),
    .B(_0238_));
 sg13g2_o21ai_1 _2981_ (.B1(_0243_),
    .Y(_0245_),
    .A1(_1584_),
    .A2(_0244_));
 sg13g2_and3_1 _2982_ (.X(_0246_),
    .A(_1590_),
    .B(_1932_),
    .C(_0238_));
 sg13g2_a21oi_2 _2983_ (.B1(_0245_),
    .Y(_0247_),
    .A2(_0246_),
    .A1(_1686_));
 sg13g2_and4_1 _2984_ (.A(_1590_),
    .B(_1894_),
    .C(_1932_),
    .D(_0238_),
    .X(_0248_));
 sg13g2_o21ai_1 _2985_ (.B1(_0248_),
    .Y(_0249_),
    .A1(_1849_),
    .A2(_1887_));
 sg13g2_and2_1 _2986_ (.A(\collatz.iter[128] ),
    .B(\collatz.iter[127] ),
    .X(_0250_));
 sg13g2_xnor2_1 _2987_ (.Y(_0251_),
    .A(\collatz.iter[128] ),
    .B(\collatz.iter[127] ));
 sg13g2_nand3_1 _2988_ (.B(_0249_),
    .C(_0251_),
    .A(_0247_),
    .Y(_0252_));
 sg13g2_a21oi_2 _2989_ (.B1(_0251_),
    .Y(_0253_),
    .A2(_0249_),
    .A1(_0247_));
 sg13g2_nor2_1 _2990_ (.A(net683),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_a22oi_1 _2991_ (.Y(_0255_),
    .B1(_0252_),
    .B2(_0254_),
    .A2(_1416_),
    .A1(net680));
 sg13g2_nor2_1 _2992_ (.A(net691),
    .B(_0255_),
    .Y(_0256_));
 sg13g2_nor2b_1 _2993_ (.A(net768),
    .B_N(\collatz.iter[128] ),
    .Y(_0257_));
 sg13g2_nor2_2 _2994_ (.A(_1508_),
    .B(_0233_),
    .Y(_0258_));
 sg13g2_a221oi_1 _2995_ (.B2(_0258_),
    .C1(_0256_),
    .B1(_0257_),
    .A1(net844),
    .Y(_0259_),
    .A2(_0234_));
 sg13g2_nor2_1 _2996_ (.A(net812),
    .B(_0259_),
    .Y(_0020_));
 sg13g2_xor2_1 _2997_ (.B(\collatz.iter[128] ),
    .A(\collatz.iter[129] ),
    .X(_0260_));
 sg13g2_xnor2_1 _2998_ (.Y(_0261_),
    .A(\collatz.iter[129] ),
    .B(\collatz.iter[128] ));
 sg13g2_o21ai_1 _2999_ (.B1(_0261_),
    .Y(_0262_),
    .A1(_0250_),
    .A2(_0253_));
 sg13g2_nor3_1 _3000_ (.A(_0250_),
    .B(_0253_),
    .C(_0261_),
    .Y(_0263_));
 sg13g2_nor2_1 _3001_ (.A(net680),
    .B(_0263_),
    .Y(_0264_));
 sg13g2_a22oi_1 _3002_ (.Y(_0265_),
    .B1(_0262_),
    .B2(_0264_),
    .A2(net261),
    .A1(net680));
 sg13g2_nand2_1 _3003_ (.Y(_0266_),
    .A(net768),
    .B(_0265_));
 sg13g2_nor2b_1 _3004_ (.A(net768),
    .B_N(\collatz.iter[129] ),
    .Y(_0267_));
 sg13g2_a22oi_1 _3005_ (.Y(_0268_),
    .B1(_0258_),
    .B2(_0267_),
    .A2(_0234_),
    .A1(net842));
 sg13g2_a21oi_1 _3006_ (.A1(_0266_),
    .A2(_0268_),
    .Y(_0021_),
    .B1(net812));
 sg13g2_nor2_1 _3007_ (.A(\collatz.iter[131] ),
    .B(net740),
    .Y(_0269_));
 sg13g2_and2_1 _3008_ (.A(\collatz.iter[130] ),
    .B(\collatz.iter[129] ),
    .X(_0270_));
 sg13g2_xor2_1 _3009_ (.B(\collatz.iter[129] ),
    .A(\collatz.iter[130] ),
    .X(_0271_));
 sg13g2_o21ai_1 _3010_ (.B1(\collatz.iter[128] ),
    .Y(_0272_),
    .A1(\collatz.iter[129] ),
    .A2(\collatz.iter[127] ));
 sg13g2_inv_1 _3011_ (.Y(_0273_),
    .A(_0272_));
 sg13g2_a21o_1 _3012_ (.A2(_0260_),
    .A1(_0253_),
    .B1(_0273_),
    .X(_0274_));
 sg13g2_xnor2_1 _3013_ (.Y(_0275_),
    .A(_0271_),
    .B(_0274_));
 sg13g2_a21oi_2 _3014_ (.B1(_0269_),
    .Y(_0276_),
    .A2(_0275_),
    .A1(net740));
 sg13g2_nand2_1 _3015_ (.Y(_0277_),
    .A(net781),
    .B(_0276_));
 sg13g2_nor2b_1 _3016_ (.A(net781),
    .B_N(net302),
    .Y(_0278_));
 sg13g2_a22oi_1 _3017_ (.Y(_0279_),
    .B1(_0258_),
    .B2(_0278_),
    .A2(_0234_),
    .A1(net840));
 sg13g2_a21oi_1 _3018_ (.A1(_0277_),
    .A2(_0279_),
    .Y(_0022_),
    .B1(net816));
 sg13g2_nor2_1 _3019_ (.A(net740),
    .B(net271),
    .Y(_0280_));
 sg13g2_nand2_1 _3020_ (.Y(_0281_),
    .A(\collatz.iter[131] ),
    .B(\collatz.iter[130] ));
 sg13g2_and2_1 _3021_ (.A(_1459_),
    .B(_0281_),
    .X(_0282_));
 sg13g2_a21oi_1 _3022_ (.A1(_0271_),
    .A2(_0274_),
    .Y(_0283_),
    .B1(_0270_));
 sg13g2_nand2b_1 _3023_ (.Y(_0284_),
    .B(_0282_),
    .A_N(_0283_));
 sg13g2_a221oi_1 _3024_ (.B2(_1459_),
    .C1(_0270_),
    .B1(_0281_),
    .A1(_0271_),
    .Y(_0285_),
    .A2(_0274_));
 sg13g2_nor2_1 _3025_ (.A(net681),
    .B(_0285_),
    .Y(_0286_));
 sg13g2_a21o_1 _3026_ (.A2(_0286_),
    .A1(_0284_),
    .B1(_0280_),
    .X(_0287_));
 sg13g2_nand2_1 _3027_ (.Y(_0288_),
    .A(net781),
    .B(_0287_));
 sg13g2_nor2b_1 _3028_ (.A(net782),
    .B_N(\collatz.iter[131] ),
    .Y(_0289_));
 sg13g2_a22oi_1 _3029_ (.Y(_0290_),
    .B1(_0258_),
    .B2(_0289_),
    .A2(_0234_),
    .A1(net839));
 sg13g2_a21oi_1 _3030_ (.A1(_0288_),
    .A2(_0290_),
    .Y(_0023_),
    .B1(net816));
 sg13g2_nand3_1 _3031_ (.B(_0273_),
    .C(_0282_),
    .A(_0271_),
    .Y(_0291_));
 sg13g2_nand3b_1 _3032_ (.B(_0281_),
    .C(_0291_),
    .Y(_0292_),
    .A_N(_0270_));
 sg13g2_nor2_1 _3033_ (.A(_0251_),
    .B(_0261_),
    .Y(_0293_));
 sg13g2_nand3_1 _3034_ (.B(_0282_),
    .C(_0293_),
    .A(_0271_),
    .Y(_0294_));
 sg13g2_a21oi_1 _3035_ (.A1(_0247_),
    .A2(_0249_),
    .Y(_0295_),
    .B1(_0294_));
 sg13g2_nand2_1 _3036_ (.Y(_0296_),
    .A(\collatz.iter[132] ),
    .B(\collatz.iter[131] ));
 sg13g2_xor2_1 _3037_ (.B(\collatz.iter[131] ),
    .A(\collatz.iter[132] ),
    .X(_0297_));
 sg13g2_o21ai_1 _3038_ (.B1(_0297_),
    .Y(_0298_),
    .A1(_0292_),
    .A2(_0295_));
 sg13g2_or3_1 _3039_ (.A(_0292_),
    .B(_0295_),
    .C(_0297_),
    .X(_0299_));
 sg13g2_nand3_1 _3040_ (.B(_0298_),
    .C(_0299_),
    .A(net740),
    .Y(_0300_));
 sg13g2_o21ai_1 _3041_ (.B1(_0300_),
    .Y(_0301_),
    .A1(_1400_),
    .A2(net741));
 sg13g2_nand2_1 _3042_ (.Y(_0302_),
    .A(net781),
    .B(_0301_));
 sg13g2_o21ai_1 _3043_ (.B1(_0302_),
    .Y(_0303_),
    .A1(net781),
    .A2(_1401_));
 sg13g2_nor3_1 _3044_ (.A(net782),
    .B(_1401_),
    .C(_0233_),
    .Y(_0304_));
 sg13g2_a21oi_1 _3045_ (.A1(net837),
    .A2(_0234_),
    .Y(_0305_),
    .B1(_0304_));
 sg13g2_a21oi_1 _3046_ (.A1(_0302_),
    .A2(_0305_),
    .Y(_0024_),
    .B1(net816));
 sg13g2_xor2_1 _3047_ (.B(\collatz.iter[132] ),
    .A(\collatz.iter[133] ),
    .X(_0306_));
 sg13g2_a21oi_1 _3048_ (.A1(_0296_),
    .A2(_0298_),
    .Y(_0307_),
    .B1(_0306_));
 sg13g2_and3_1 _3049_ (.X(_0308_),
    .A(_0296_),
    .B(_0298_),
    .C(_0306_));
 sg13g2_o21ai_1 _3050_ (.B1(net741),
    .Y(_0309_),
    .A1(_0307_),
    .A2(_0308_));
 sg13g2_o21ai_1 _3051_ (.B1(_0309_),
    .Y(_0310_),
    .A1(net741),
    .A2(net266));
 sg13g2_nand2_1 _3052_ (.Y(_0311_),
    .A(net782),
    .B(_0310_));
 sg13g2_nor3_1 _3053_ (.A(net783),
    .B(_1400_),
    .C(_0233_),
    .Y(_0312_));
 sg13g2_a21oi_1 _3054_ (.A1(net835),
    .A2(_0234_),
    .Y(_0313_),
    .B1(_0312_));
 sg13g2_a21oi_1 _3055_ (.A1(_0311_),
    .A2(_0313_),
    .Y(_0025_),
    .B1(net817));
 sg13g2_xnor2_1 _3056_ (.Y(_0314_),
    .A(\collatz.iter[134] ),
    .B(\collatz.iter[133] ));
 sg13g2_o21ai_1 _3057_ (.B1(\collatz.iter[132] ),
    .Y(_0315_),
    .A1(\collatz.iter[133] ),
    .A2(\collatz.iter[131] ));
 sg13g2_a21oi_1 _3058_ (.A1(_0298_),
    .A2(_0315_),
    .Y(_0316_),
    .B1(_1446_));
 sg13g2_a221oi_1 _3059_ (.B2(_0315_),
    .C1(_0314_),
    .B1(_0298_),
    .A1(_1400_),
    .Y(_0317_),
    .A2(_1401_));
 sg13g2_xor2_1 _3060_ (.B(_0316_),
    .A(_0314_),
    .X(_0318_));
 sg13g2_nor2_1 _3061_ (.A(\collatz.iter[135] ),
    .B(net741),
    .Y(_0319_));
 sg13g2_a21oi_2 _3062_ (.B1(_0319_),
    .Y(_0320_),
    .A2(_0318_),
    .A1(net741));
 sg13g2_nand2_1 _3063_ (.Y(_0321_),
    .A(net782),
    .B(_0320_));
 sg13g2_nor2b_1 _3064_ (.A(net783),
    .B_N(net324),
    .Y(_0322_));
 sg13g2_a22oi_1 _3065_ (.Y(_0323_),
    .B1(_0258_),
    .B2(_0322_),
    .A2(_0234_),
    .A1(net833));
 sg13g2_a21oi_1 _3066_ (.A1(_0321_),
    .A2(_0323_),
    .Y(_0026_),
    .B1(net817));
 sg13g2_xnor2_1 _3067_ (.Y(_0324_),
    .A(\collatz.iter[135] ),
    .B(\collatz.iter[134] ));
 sg13g2_a21oi_1 _3068_ (.A1(\collatz.iter[134] ),
    .A2(\collatz.iter[133] ),
    .Y(_0325_),
    .B1(_0317_));
 sg13g2_xnor2_1 _3069_ (.Y(_0326_),
    .A(_0324_),
    .B(_0325_));
 sg13g2_mux2_1 _3070_ (.A0(net268),
    .A1(_0326_),
    .S(net741),
    .X(_0327_));
 sg13g2_nand2b_1 _3071_ (.Y(_0328_),
    .B(net784),
    .A_N(_0327_));
 sg13g2_nor3_1 _3072_ (.A(net784),
    .B(_1399_),
    .C(_0233_),
    .Y(_0329_));
 sg13g2_a21oi_1 _3073_ (.A1(net831),
    .A2(_0234_),
    .Y(_0330_),
    .B1(_0329_));
 sg13g2_a21oi_1 _3074_ (.A1(_0328_),
    .A2(_0330_),
    .Y(_0027_),
    .B1(net817));
 sg13g2_nor2_1 _3075_ (.A(\collatz.iter[137] ),
    .B(net741),
    .Y(_0331_));
 sg13g2_nand2_1 _3076_ (.Y(_0332_),
    .A(_0297_),
    .B(_0306_));
 sg13g2_or2_1 _3077_ (.X(_0333_),
    .B(_0324_),
    .A(_0314_));
 sg13g2_nor3_1 _3078_ (.A(_0294_),
    .B(_0332_),
    .C(_0333_),
    .Y(_0334_));
 sg13g2_inv_1 _3079_ (.Y(_0335_),
    .A(_0334_));
 sg13g2_a21oi_2 _3080_ (.B1(_0335_),
    .Y(_0336_),
    .A2(_0249_),
    .A1(_0247_));
 sg13g2_nand2b_1 _3081_ (.Y(_0337_),
    .B(_0292_),
    .A_N(_0332_));
 sg13g2_a21oi_1 _3082_ (.A1(_0315_),
    .A2(_0337_),
    .Y(_0338_),
    .B1(_0333_));
 sg13g2_o21ai_1 _3083_ (.B1(\collatz.iter[134] ),
    .Y(_0339_),
    .A1(\collatz.iter[135] ),
    .A2(\collatz.iter[133] ));
 sg13g2_nand2b_2 _3084_ (.Y(_0340_),
    .B(_0339_),
    .A_N(_0338_));
 sg13g2_nor2_1 _3085_ (.A(_0336_),
    .B(_0340_),
    .Y(_0341_));
 sg13g2_nand2_1 _3086_ (.Y(_0342_),
    .A(\collatz.iter[136] ),
    .B(\collatz.iter[135] ));
 sg13g2_xnor2_1 _3087_ (.Y(_0343_),
    .A(\collatz.iter[136] ),
    .B(\collatz.iter[135] ));
 sg13g2_xnor2_1 _3088_ (.Y(_0344_),
    .A(_0341_),
    .B(_0343_));
 sg13g2_a21oi_1 _3089_ (.A1(net749),
    .A2(_0344_),
    .Y(_0345_),
    .B1(_0331_));
 sg13g2_nand2_1 _3090_ (.Y(_0346_),
    .A(net784),
    .B(_0345_));
 sg13g2_nor3_2 _3091_ (.A(net796),
    .B(_1417_),
    .C(_1514_),
    .Y(_0347_));
 sg13g2_nor4_2 _3092_ (.A(net3),
    .B(net1),
    .C(net2),
    .Y(_0348_),
    .D(_1419_));
 sg13g2_and2_1 _3093_ (.A(net845),
    .B(net678),
    .X(_0349_));
 sg13g2_nor2_1 _3094_ (.A(net784),
    .B(_1398_),
    .Y(_0350_));
 sg13g2_a21oi_2 _3095_ (.B1(_1508_),
    .Y(_0351_),
    .A2(net677),
    .A1(_0232_));
 sg13g2_a22oi_1 _3096_ (.Y(_0352_),
    .B1(_0350_),
    .B2(_0351_),
    .A2(_0349_),
    .A1(_0347_));
 sg13g2_a21oi_1 _3097_ (.A1(_0346_),
    .A2(_0352_),
    .Y(_0028_),
    .B1(net817));
 sg13g2_xnor2_1 _3098_ (.Y(_0353_),
    .A(\collatz.iter[137] ),
    .B(\collatz.iter[136] ));
 sg13g2_o21ai_1 _3099_ (.B1(_0342_),
    .Y(_0354_),
    .A1(_0341_),
    .A2(_0343_));
 sg13g2_nor2_1 _3100_ (.A(net750),
    .B(net301),
    .Y(_0355_));
 sg13g2_xnor2_1 _3101_ (.Y(_0356_),
    .A(_0353_),
    .B(_0354_));
 sg13g2_a21oi_1 _3102_ (.A1(net749),
    .A2(_0356_),
    .Y(_0357_),
    .B1(_0355_));
 sg13g2_or2_1 _3103_ (.X(_0358_),
    .B(_0357_),
    .A(net692));
 sg13g2_and2_1 _3104_ (.A(net843),
    .B(net678),
    .X(_0359_));
 sg13g2_nor2_1 _3105_ (.A(net784),
    .B(_1397_),
    .Y(_0360_));
 sg13g2_a22oi_1 _3106_ (.Y(_0361_),
    .B1(_0360_),
    .B2(_0351_),
    .A2(_0359_),
    .A1(_0347_));
 sg13g2_a21oi_1 _3107_ (.A1(_0358_),
    .A2(_0361_),
    .Y(_0029_),
    .B1(net817));
 sg13g2_and2_1 _3108_ (.A(\collatz.iter[138] ),
    .B(\collatz.iter[137] ),
    .X(_0362_));
 sg13g2_xnor2_1 _3109_ (.Y(_0363_),
    .A(\collatz.iter[138] ),
    .B(\collatz.iter[137] ));
 sg13g2_o21ai_1 _3110_ (.B1(\collatz.iter[136] ),
    .Y(_0364_),
    .A1(\collatz.iter[137] ),
    .A2(\collatz.iter[135] ));
 sg13g2_nor2_1 _3111_ (.A(_0343_),
    .B(_0353_),
    .Y(_0365_));
 sg13g2_o21ai_1 _3112_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_0336_),
    .A2(_0340_));
 sg13g2_a21oi_1 _3113_ (.A1(_0364_),
    .A2(_0366_),
    .Y(_0367_),
    .B1(_0363_));
 sg13g2_nand3_1 _3114_ (.B(_0364_),
    .C(_0366_),
    .A(_0363_),
    .Y(_0368_));
 sg13g2_nand3b_1 _3115_ (.B(_0368_),
    .C(net749),
    .Y(_0369_),
    .A_N(_0367_));
 sg13g2_o21ai_1 _3116_ (.B1(_0369_),
    .Y(_0370_),
    .A1(_1396_),
    .A2(net749));
 sg13g2_nand3_1 _3117_ (.B(_0347_),
    .C(net678),
    .A(net841),
    .Y(_0371_));
 sg13g2_nor2b_1 _3118_ (.A(net784),
    .B_N(\collatz.iter[138] ),
    .Y(_0372_));
 sg13g2_a22oi_1 _3119_ (.Y(_0373_),
    .B1(_0372_),
    .B2(_0351_),
    .A2(_0370_),
    .A1(net786));
 sg13g2_a21oi_1 _3120_ (.A1(_0371_),
    .A2(_0373_),
    .Y(_0030_),
    .B1(net823));
 sg13g2_xor2_1 _3121_ (.B(\collatz.iter[138] ),
    .A(\collatz.iter[139] ),
    .X(_0374_));
 sg13g2_xnor2_1 _3122_ (.Y(_0375_),
    .A(\collatz.iter[139] ),
    .B(\collatz.iter[138] ));
 sg13g2_or2_1 _3123_ (.X(_0376_),
    .B(net277),
    .A(net749));
 sg13g2_or3_1 _3124_ (.A(_0362_),
    .B(_0367_),
    .C(_0374_),
    .X(_0377_));
 sg13g2_o21ai_1 _3125_ (.B1(_0374_),
    .Y(_0378_),
    .A1(_0362_),
    .A2(_0367_));
 sg13g2_nand3_1 _3126_ (.B(_0377_),
    .C(_0378_),
    .A(net749),
    .Y(_0379_));
 sg13g2_a21o_1 _3127_ (.A2(_0379_),
    .A1(_0376_),
    .B1(net692),
    .X(_0380_));
 sg13g2_nor2_1 _3128_ (.A(net786),
    .B(_1396_),
    .Y(_0381_));
 sg13g2_and2_1 _3129_ (.A(net839),
    .B(net678),
    .X(_0382_));
 sg13g2_a22oi_1 _3130_ (.Y(_0383_),
    .B1(_0382_),
    .B2(_0347_),
    .A2(_0381_),
    .A1(_0351_));
 sg13g2_a21oi_1 _3131_ (.A1(_0380_),
    .A2(_0383_),
    .Y(_0031_),
    .B1(net823));
 sg13g2_nand3b_1 _3132_ (.B(_0365_),
    .C(_0374_),
    .Y(_0384_),
    .A_N(_0363_));
 sg13g2_inv_1 _3133_ (.Y(_0385_),
    .A(_0384_));
 sg13g2_o21ai_1 _3134_ (.B1(_0385_),
    .Y(_0386_),
    .A1(_0336_),
    .A2(_0340_));
 sg13g2_nor3_1 _3135_ (.A(_0363_),
    .B(_0364_),
    .C(_0375_),
    .Y(_0387_));
 sg13g2_o21ai_1 _3136_ (.B1(\collatz.iter[138] ),
    .Y(_0388_),
    .A1(\collatz.iter[139] ),
    .A2(\collatz.iter[137] ));
 sg13g2_nor2b_2 _3137_ (.A(_0387_),
    .B_N(_0388_),
    .Y(_0389_));
 sg13g2_xnor2_1 _3138_ (.Y(_0390_),
    .A(\collatz.iter[140] ),
    .B(\collatz.iter[139] ));
 sg13g2_a21oi_1 _3139_ (.A1(_0386_),
    .A2(_0389_),
    .Y(_0391_),
    .B1(_0390_));
 sg13g2_nand3_1 _3140_ (.B(_0389_),
    .C(_0390_),
    .A(_0386_),
    .Y(_0392_));
 sg13g2_nand3b_1 _3141_ (.B(_0392_),
    .C(net749),
    .Y(_0393_),
    .A_N(_0391_));
 sg13g2_o21ai_1 _3142_ (.B1(_0393_),
    .Y(_0394_),
    .A1(_1394_),
    .A2(net749));
 sg13g2_nand2_1 _3143_ (.Y(_0395_),
    .A(net787),
    .B(_0394_));
 sg13g2_and2_1 _3144_ (.A(net837),
    .B(net678),
    .X(_0396_));
 sg13g2_nor2_1 _3145_ (.A(net786),
    .B(_1395_),
    .Y(_0397_));
 sg13g2_a22oi_1 _3146_ (.Y(_0398_),
    .B1(_0397_),
    .B2(_0351_),
    .A2(_0396_),
    .A1(_0347_));
 sg13g2_a21oi_1 _3147_ (.A1(_0395_),
    .A2(_0398_),
    .Y(_0032_),
    .B1(net823));
 sg13g2_xor2_1 _3148_ (.B(\collatz.iter[140] ),
    .A(\collatz.iter[141] ),
    .X(_0399_));
 sg13g2_a21oi_1 _3149_ (.A1(\collatz.iter[140] ),
    .A2(\collatz.iter[139] ),
    .Y(_0400_),
    .B1(_0391_));
 sg13g2_or2_1 _3150_ (.X(_0401_),
    .B(_0000_),
    .A(net750));
 sg13g2_xor2_1 _3151_ (.B(_0400_),
    .A(_0399_),
    .X(_0402_));
 sg13g2_o21ai_1 _3152_ (.B1(_0401_),
    .Y(_0403_),
    .A1(net682),
    .A2(_0402_));
 sg13g2_nand2_1 _3153_ (.Y(_0404_),
    .A(net787),
    .B(_0403_));
 sg13g2_nor2_1 _3154_ (.A(net786),
    .B(_1394_),
    .Y(_0405_));
 sg13g2_and2_1 _3155_ (.A(net835),
    .B(net677),
    .X(_0406_));
 sg13g2_a22oi_1 _3156_ (.Y(_0407_),
    .B1(_0406_),
    .B2(_0347_),
    .A2(_0405_),
    .A1(_0351_));
 sg13g2_a21oi_1 _3157_ (.A1(_0404_),
    .A2(_0407_),
    .Y(_0033_),
    .B1(net823));
 sg13g2_nand2_1 _3158_ (.Y(_0408_),
    .A(\collatz.iter[142] ),
    .B(\collatz.iter[141] ));
 sg13g2_xnor2_1 _3159_ (.Y(_0409_),
    .A(\collatz.iter[142] ),
    .B(\collatz.iter[141] ));
 sg13g2_inv_1 _3160_ (.Y(_0410_),
    .A(_0409_));
 sg13g2_nor2b_1 _3161_ (.A(_0390_),
    .B_N(_0399_),
    .Y(_0411_));
 sg13g2_inv_1 _3162_ (.Y(_0412_),
    .A(_0411_));
 sg13g2_a21oi_1 _3163_ (.A1(_0386_),
    .A2(_0389_),
    .Y(_0413_),
    .B1(_0412_));
 sg13g2_a21oi_1 _3164_ (.A1(_1394_),
    .A2(_1396_),
    .Y(_0414_),
    .B1(_1395_));
 sg13g2_o21ai_1 _3165_ (.B1(_0410_),
    .Y(_0415_),
    .A1(_0413_),
    .A2(_0414_));
 sg13g2_nor3_1 _3166_ (.A(_0410_),
    .B(_0413_),
    .C(_0414_),
    .Y(_0416_));
 sg13g2_nor2_1 _3167_ (.A(net682),
    .B(_0416_),
    .Y(_0417_));
 sg13g2_a22oi_1 _3168_ (.Y(_0418_),
    .B1(_0415_),
    .B2(_0417_),
    .A2(net682),
    .A1(\collatz.iter[143] ));
 sg13g2_or2_1 _3169_ (.X(_0419_),
    .B(_0418_),
    .A(net692));
 sg13g2_and2_1 _3170_ (.A(net833),
    .B(net677),
    .X(_0420_));
 sg13g2_nor2_1 _3171_ (.A(net786),
    .B(_1393_),
    .Y(_0421_));
 sg13g2_a22oi_1 _3172_ (.Y(_0422_),
    .B1(_0421_),
    .B2(_0351_),
    .A2(_0420_),
    .A1(_0347_));
 sg13g2_a21oi_1 _3173_ (.A1(_0419_),
    .A2(_0422_),
    .Y(_0034_),
    .B1(net823));
 sg13g2_xnor2_1 _3174_ (.Y(_0423_),
    .A(\collatz.iter[143] ),
    .B(\collatz.iter[142] ));
 sg13g2_nand3_1 _3175_ (.B(_0415_),
    .C(_0423_),
    .A(_0408_),
    .Y(_0424_));
 sg13g2_a21o_1 _3176_ (.A2(_0415_),
    .A1(_0408_),
    .B1(_0423_),
    .X(_0425_));
 sg13g2_and3_1 _3177_ (.X(_0426_),
    .A(net750),
    .B(_0424_),
    .C(_0425_));
 sg13g2_nand3_1 _3178_ (.B(_0424_),
    .C(_0425_),
    .A(net750),
    .Y(_0427_));
 sg13g2_nand2_1 _3179_ (.Y(_0428_),
    .A(net796),
    .B(_0426_));
 sg13g2_and2_1 _3180_ (.A(net831),
    .B(_0348_),
    .X(_0429_));
 sg13g2_nor2b_1 _3181_ (.A(net796),
    .B_N(\collatz.iter[143] ),
    .Y(_0430_));
 sg13g2_a22oi_1 _3182_ (.Y(_0431_),
    .B1(_0430_),
    .B2(_0351_),
    .A2(_0429_),
    .A1(_0347_));
 sg13g2_a21oi_1 _3183_ (.A1(_0428_),
    .A2(_0431_),
    .Y(_0035_),
    .B1(net822));
 sg13g2_nand2_1 _3184_ (.Y(_0432_),
    .A(net6),
    .B(net850));
 sg13g2_o21ai_1 _3185_ (.B1(net850),
    .Y(_0433_),
    .A1(net796),
    .A2(net6));
 sg13g2_nor2_1 _3186_ (.A(_1507_),
    .B(_0433_),
    .Y(_0036_));
 sg13g2_nand2b_1 _3187_ (.Y(_0434_),
    .B(net692),
    .A_N(_0432_));
 sg13g2_inv_1 _3188_ (.Y(_0435_),
    .A(_0434_));
 sg13g2_nand2_2 _3189_ (.Y(_0436_),
    .A(net853),
    .B(net673));
 sg13g2_xnor2_1 _3190_ (.Y(_0437_),
    .A(net253),
    .B(net788));
 sg13g2_nor2_1 _3191_ (.A(_0436_),
    .B(_0437_),
    .Y(_0037_));
 sg13g2_and3_1 _3192_ (.X(_0438_),
    .A(net210),
    .B(\collatz.orbit_len[0] ),
    .C(net788));
 sg13g2_a21oi_1 _3193_ (.A1(\collatz.orbit_len[0] ),
    .A2(net788),
    .Y(_0439_),
    .B1(net210));
 sg13g2_nor3_1 _3194_ (.A(_0436_),
    .B(_0438_),
    .C(net211),
    .Y(_0038_));
 sg13g2_nor2_1 _3195_ (.A(net226),
    .B(_0438_),
    .Y(_0440_));
 sg13g2_nor2_1 _3196_ (.A(net692),
    .B(_1423_),
    .Y(_0441_));
 sg13g2_nor3_1 _3197_ (.A(_0436_),
    .B(net227),
    .C(_0441_),
    .Y(_0039_));
 sg13g2_nor2_1 _3198_ (.A(net231),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_and2_1 _3199_ (.A(net231),
    .B(_0441_),
    .X(_0443_));
 sg13g2_nor3_1 _3200_ (.A(_0436_),
    .B(net232),
    .C(_0443_),
    .Y(_0040_));
 sg13g2_a21oi_1 _3201_ (.A1(net246),
    .A2(net673),
    .Y(_0444_),
    .B1(_0443_));
 sg13g2_and2_1 _3202_ (.A(net246),
    .B(_0443_),
    .X(_0445_));
 sg13g2_nor3_1 _3203_ (.A(net821),
    .B(_0444_),
    .C(_0445_),
    .Y(_0041_));
 sg13g2_a21oi_1 _3204_ (.A1(net238),
    .A2(net673),
    .Y(_0446_),
    .B1(_0445_));
 sg13g2_and2_1 _3205_ (.A(net238),
    .B(_0445_),
    .X(_0447_));
 sg13g2_nor3_1 _3206_ (.A(net821),
    .B(net239),
    .C(_0447_),
    .Y(_0042_));
 sg13g2_nor2_1 _3207_ (.A(net224),
    .B(_0447_),
    .Y(_0448_));
 sg13g2_nor2b_2 _3208_ (.A(_1422_),
    .B_N(_0443_),
    .Y(_0449_));
 sg13g2_nor3_1 _3209_ (.A(_0436_),
    .B(net225),
    .C(_0449_),
    .Y(_0043_));
 sg13g2_a21oi_1 _3210_ (.A1(net254),
    .A2(net673),
    .Y(_0450_),
    .B1(_0449_));
 sg13g2_a21oi_1 _3211_ (.A1(net254),
    .A2(_0449_),
    .Y(_0451_),
    .B1(net821));
 sg13g2_nor2b_1 _3212_ (.A(_0450_),
    .B_N(_0451_),
    .Y(_0044_));
 sg13g2_a22oi_1 _3213_ (.Y(_0452_),
    .B1(_0449_),
    .B2(\collatz.orbit_len[7] ),
    .A2(net673),
    .A1(net243));
 sg13g2_and3_1 _3214_ (.X(_0453_),
    .A(net243),
    .B(net254),
    .C(_0449_));
 sg13g2_nor3_1 _3215_ (.A(net821),
    .B(net244),
    .C(_0453_),
    .Y(_0045_));
 sg13g2_nor2_1 _3216_ (.A(net255),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_and2_1 _3217_ (.A(net255),
    .B(_0453_),
    .X(_0455_));
 sg13g2_nor3_1 _3218_ (.A(_0436_),
    .B(_0454_),
    .C(_0455_),
    .Y(_0046_));
 sg13g2_a21oi_1 _3219_ (.A1(net251),
    .A2(net673),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_a21oi_1 _3220_ (.A1(net251),
    .A2(_0455_),
    .Y(_0457_),
    .B1(net823));
 sg13g2_nor2b_1 _3221_ (.A(net252),
    .B_N(_0457_),
    .Y(_0047_));
 sg13g2_a22oi_1 _3222_ (.Y(_0458_),
    .B1(_0455_),
    .B2(\collatz.orbit_len[10] ),
    .A2(net673),
    .A1(net219));
 sg13g2_nand3_1 _3223_ (.B(\collatz.orbit_len[10] ),
    .C(_0455_),
    .A(net219),
    .Y(_0459_));
 sg13g2_inv_1 _3224_ (.Y(_0460_),
    .A(_0459_));
 sg13g2_nor3_1 _3225_ (.A(net821),
    .B(net220),
    .C(_0460_),
    .Y(_0048_));
 sg13g2_xor2_1 _3226_ (.B(_0459_),
    .A(net241),
    .X(_0461_));
 sg13g2_nor2_1 _3227_ (.A(_0436_),
    .B(net242),
    .Y(_0049_));
 sg13g2_a22oi_1 _3228_ (.Y(_0462_),
    .B1(_0460_),
    .B2(\collatz.orbit_len[12] ),
    .A2(net673),
    .A1(net215));
 sg13g2_nand2b_1 _3229_ (.Y(_0463_),
    .B(_0453_),
    .A_N(_1421_));
 sg13g2_nand2_1 _3230_ (.Y(_0464_),
    .A(net853),
    .B(_0463_));
 sg13g2_nor2_1 _3231_ (.A(net216),
    .B(_0464_),
    .Y(_0050_));
 sg13g2_xor2_1 _3232_ (.B(_0463_),
    .A(net259),
    .X(_0465_));
 sg13g2_nor2_1 _3233_ (.A(_0436_),
    .B(_0465_),
    .Y(_0051_));
 sg13g2_nand3_1 _3234_ (.B(net692),
    .C(_0432_),
    .A(net229),
    .Y(_0466_));
 sg13g2_a221oi_1 _3235_ (.B2(_0466_),
    .C1(net821),
    .B1(_1426_),
    .A1(_1390_),
    .Y(_0052_),
    .A2(_1425_));
 sg13g2_a221oi_1 _3236_ (.B2(_0417_),
    .C1(_1376_),
    .B1(_0415_),
    .A1(\collatz.iter[143] ),
    .Y(_0467_),
    .A2(net682));
 sg13g2_a21o_1 _3237_ (.A2(_0427_),
    .A1(_1414_),
    .B1(_0467_),
    .X(_0468_));
 sg13g2_nand4_1 _3238_ (.B(_0008_),
    .C(_0424_),
    .A(net750),
    .Y(_0469_),
    .D(_0425_));
 sg13g2_o21ai_1 _3239_ (.B1(_0469_),
    .Y(_0470_),
    .A1(\collatz.path_record_h16[14] ),
    .A2(_0418_));
 sg13g2_nor2_1 _3240_ (.A(_0468_),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_nand2b_1 _3241_ (.Y(_0472_),
    .B(\collatz.path_record_h16[13] ),
    .A_N(_0403_));
 sg13g2_nand2b_1 _3242_ (.Y(_0473_),
    .B(\collatz.path_record_h16[12] ),
    .A_N(_0394_));
 sg13g2_xnor2_1 _3243_ (.Y(_0474_),
    .A(_1378_),
    .B(_0394_));
 sg13g2_and2_1 _3244_ (.A(_1377_),
    .B(_0403_),
    .X(_0475_));
 sg13g2_xnor2_1 _3245_ (.Y(_0476_),
    .A(_1377_),
    .B(_0403_));
 sg13g2_nor4_2 _3246_ (.A(_0468_),
    .B(_0470_),
    .C(_0474_),
    .Y(_0477_),
    .D(_0476_));
 sg13g2_and3_1 _3247_ (.X(_0478_),
    .A(\collatz.path_record_h16[11] ),
    .B(_0376_),
    .C(_0379_));
 sg13g2_nand3_1 _3248_ (.B(_0376_),
    .C(_0379_),
    .A(\collatz.path_record_h16[11] ),
    .Y(_0479_));
 sg13g2_a21oi_1 _3249_ (.A1(_0376_),
    .A2(_0379_),
    .Y(_0480_),
    .B1(\collatz.path_record_h16[11] ));
 sg13g2_nand2b_1 _3250_ (.Y(_0481_),
    .B(\collatz.path_record_h16[10] ),
    .A_N(_0370_));
 sg13g2_xnor2_1 _3251_ (.Y(_0482_),
    .A(_1380_),
    .B(_0370_));
 sg13g2_nor3_1 _3252_ (.A(_0478_),
    .B(_0480_),
    .C(_0482_),
    .Y(_0483_));
 sg13g2_nand2_1 _3253_ (.Y(_0484_),
    .A(\collatz.path_record_h16[9] ),
    .B(_0357_));
 sg13g2_nor2_1 _3254_ (.A(\collatz.path_record_h16[9] ),
    .B(_0357_),
    .Y(_0485_));
 sg13g2_nand2b_1 _3255_ (.Y(_0486_),
    .B(\collatz.path_record_h16[8] ),
    .A_N(_0345_));
 sg13g2_o21ai_1 _3256_ (.B1(_0484_),
    .Y(_0487_),
    .A1(_0485_),
    .A2(_0486_));
 sg13g2_o21ai_1 _3257_ (.B1(_0479_),
    .Y(_0488_),
    .A1(_0480_),
    .A2(_0481_));
 sg13g2_a21o_1 _3258_ (.A2(_0487_),
    .A1(_0483_),
    .B1(_0488_),
    .X(_0489_));
 sg13g2_a21o_1 _3259_ (.A2(_0469_),
    .A1(_0468_),
    .B1(net694),
    .X(_0490_));
 sg13g2_o21ai_1 _3260_ (.B1(_0472_),
    .Y(_0491_),
    .A1(_0473_),
    .A2(_0475_));
 sg13g2_a221oi_1 _3261_ (.B2(_0471_),
    .C1(_0490_),
    .B1(_0491_),
    .A1(_0477_),
    .Y(_0492_),
    .A2(_0489_));
 sg13g2_and2_1 _3262_ (.A(_1384_),
    .B(_0320_),
    .X(_0493_));
 sg13g2_nand2_1 _3263_ (.Y(_0494_),
    .A(_1385_),
    .B(_0310_));
 sg13g2_nand2b_1 _3264_ (.Y(_0495_),
    .B(\collatz.path_record_h16[4] ),
    .A_N(_0301_));
 sg13g2_o21ai_1 _3265_ (.B1(_0495_),
    .Y(_0496_),
    .A1(_1385_),
    .A2(_0310_));
 sg13g2_a221oi_1 _3266_ (.B2(_0286_),
    .C1(_1387_),
    .B1(_0284_),
    .A1(net681),
    .Y(_0497_),
    .A2(_1415_));
 sg13g2_nor2_1 _3267_ (.A(_1388_),
    .B(_0276_),
    .Y(_0498_));
 sg13g2_o21ai_1 _3268_ (.B1(\collatz.path_record_h16[1] ),
    .Y(_0499_),
    .A1(\collatz.path_record_h16[0] ),
    .A2(_0255_));
 sg13g2_nor3_1 _3269_ (.A(\collatz.path_record_h16[1] ),
    .B(\collatz.path_record_h16[0] ),
    .C(_0255_),
    .Y(_0500_));
 sg13g2_a221oi_1 _3270_ (.B2(_0265_),
    .C1(_0500_),
    .B1(_0499_),
    .A1(_1388_),
    .Y(_0501_),
    .A2(_0276_));
 sg13g2_or3_1 _3271_ (.A(_0497_),
    .B(_0498_),
    .C(_0501_),
    .X(_0502_));
 sg13g2_xnor2_1 _3272_ (.Y(_0503_),
    .A(_1386_),
    .B(_0301_));
 sg13g2_a221oi_1 _3273_ (.B2(_1385_),
    .C1(_0503_),
    .B1(_0310_),
    .A1(_1387_),
    .Y(_0504_),
    .A2(_0287_));
 sg13g2_nand2_1 _3274_ (.Y(_0505_),
    .A(\collatz.path_record_h16[7] ),
    .B(_0327_));
 sg13g2_nor2_1 _3275_ (.A(_1384_),
    .B(_0320_),
    .Y(_0506_));
 sg13g2_a221oi_1 _3276_ (.B2(_0504_),
    .C1(_0506_),
    .B1(_0502_),
    .A1(_0494_),
    .Y(_0507_),
    .A2(_0496_));
 sg13g2_o21ai_1 _3277_ (.B1(_0505_),
    .Y(_0508_),
    .A1(_0493_),
    .A2(_0507_));
 sg13g2_nor2_1 _3278_ (.A(\collatz.path_record_h16[7] ),
    .B(_0327_),
    .Y(_0509_));
 sg13g2_nand2_1 _3279_ (.Y(_0510_),
    .A(_1382_),
    .B(_0345_));
 sg13g2_nand3_1 _3280_ (.B(_0486_),
    .C(_0510_),
    .A(_0484_),
    .Y(_0511_));
 sg13g2_nor3_1 _3281_ (.A(_0485_),
    .B(_0509_),
    .C(_0511_),
    .Y(_0512_));
 sg13g2_nand4_1 _3282_ (.B(_0483_),
    .C(_0508_),
    .A(_0477_),
    .Y(_0513_),
    .D(_0512_));
 sg13g2_a21oi_1 _3283_ (.A1(_0492_),
    .A2(_0513_),
    .Y(_0514_),
    .B1(_0435_));
 sg13g2_nand2b_1 _3284_ (.Y(_0515_),
    .B(net645),
    .A_N(net273));
 sg13g2_or3_1 _3285_ (.A(_0256_),
    .B(_0257_),
    .C(net645),
    .X(_0516_));
 sg13g2_and3_1 _3286_ (.X(_0053_),
    .A(net847),
    .B(_0515_),
    .C(_0516_));
 sg13g2_a21o_1 _3287_ (.A2(_0265_),
    .A1(net781),
    .B1(_0267_),
    .X(_0517_));
 sg13g2_o21ai_1 _3288_ (.B1(net848),
    .Y(_0518_),
    .A1(net645),
    .A2(_0517_));
 sg13g2_a21oi_1 _3289_ (.A1(_1389_),
    .A2(net645),
    .Y(_0054_),
    .B1(_0518_));
 sg13g2_a21o_1 _3290_ (.A2(_0276_),
    .A1(net781),
    .B1(_0278_),
    .X(_0519_));
 sg13g2_o21ai_1 _3291_ (.B1(net848),
    .Y(_0520_),
    .A1(net645),
    .A2(_0519_));
 sg13g2_a21oi_1 _3292_ (.A1(_1388_),
    .A2(net645),
    .Y(_0055_),
    .B1(_0520_));
 sg13g2_a21o_1 _3293_ (.A2(_0287_),
    .A1(net781),
    .B1(_0289_),
    .X(_0521_));
 sg13g2_o21ai_1 _3294_ (.B1(net848),
    .Y(_0522_),
    .A1(net646),
    .A2(_0521_));
 sg13g2_a21oi_1 _3295_ (.A1(_1387_),
    .A2(net646),
    .Y(_0056_),
    .B1(_0522_));
 sg13g2_o21ai_1 _3296_ (.B1(net848),
    .Y(_0523_),
    .A1(_0303_),
    .A2(net646));
 sg13g2_a21oi_1 _3297_ (.A1(_1386_),
    .A2(net646),
    .Y(_0057_),
    .B1(_0523_));
 sg13g2_o21ai_1 _3298_ (.B1(_0311_),
    .Y(_0524_),
    .A1(net782),
    .A2(_1400_));
 sg13g2_o21ai_1 _3299_ (.B1(net848),
    .Y(_0525_),
    .A1(net645),
    .A2(_0524_));
 sg13g2_a21oi_1 _3300_ (.A1(_1385_),
    .A2(net646),
    .Y(_0058_),
    .B1(_0525_));
 sg13g2_a21o_1 _3301_ (.A2(_0320_),
    .A1(net782),
    .B1(_0322_),
    .X(_0526_));
 sg13g2_o21ai_1 _3302_ (.B1(net848),
    .Y(_0527_),
    .A1(net646),
    .A2(_0526_));
 sg13g2_a21oi_1 _3303_ (.A1(_1384_),
    .A2(net645),
    .Y(_0059_),
    .B1(_0527_));
 sg13g2_o21ai_1 _3304_ (.B1(_0328_),
    .Y(_0528_),
    .A1(net782),
    .A2(_1399_));
 sg13g2_o21ai_1 _3305_ (.B1(net848),
    .Y(_0529_),
    .A1(net648),
    .A2(_0528_));
 sg13g2_a21oi_1 _3306_ (.A1(_1383_),
    .A2(net648),
    .Y(_0060_),
    .B1(_0529_));
 sg13g2_o21ai_1 _3307_ (.B1(_0346_),
    .Y(_0530_),
    .A1(net784),
    .A2(_1398_));
 sg13g2_o21ai_1 _3308_ (.B1(net850),
    .Y(_0531_),
    .A1(net648),
    .A2(_0530_));
 sg13g2_a21oi_1 _3309_ (.A1(_1382_),
    .A2(net648),
    .Y(_0061_),
    .B1(_0531_));
 sg13g2_o21ai_1 _3310_ (.B1(_0358_),
    .Y(_0532_),
    .A1(net784),
    .A2(_1397_));
 sg13g2_o21ai_1 _3311_ (.B1(net850),
    .Y(_0533_),
    .A1(net648),
    .A2(_0532_));
 sg13g2_a21oi_1 _3312_ (.A1(_1381_),
    .A2(net648),
    .Y(_0062_),
    .B1(_0533_));
 sg13g2_a21oi_1 _3313_ (.A1(net787),
    .A2(_0370_),
    .Y(_0534_),
    .B1(_0372_));
 sg13g2_mux2_1 _3314_ (.A0(_0534_),
    .A1(_1380_),
    .S(net648),
    .X(_0535_));
 sg13g2_nor2_1 _3315_ (.A(net823),
    .B(_0535_),
    .Y(_0063_));
 sg13g2_o21ai_1 _3316_ (.B1(_0380_),
    .Y(_0536_),
    .A1(net786),
    .A2(_1396_));
 sg13g2_o21ai_1 _3317_ (.B1(net850),
    .Y(_0537_),
    .A1(net647),
    .A2(_0536_));
 sg13g2_a21oi_1 _3318_ (.A1(_1379_),
    .A2(net647),
    .Y(_0064_),
    .B1(_0537_));
 sg13g2_o21ai_1 _3319_ (.B1(_0395_),
    .Y(_0538_),
    .A1(net786),
    .A2(_1395_));
 sg13g2_o21ai_1 _3320_ (.B1(net850),
    .Y(_0539_),
    .A1(net649),
    .A2(_0538_));
 sg13g2_a21oi_1 _3321_ (.A1(_1378_),
    .A2(net648),
    .Y(_0065_),
    .B1(_0539_));
 sg13g2_o21ai_1 _3322_ (.B1(_0404_),
    .Y(_0540_),
    .A1(net787),
    .A2(_1394_));
 sg13g2_o21ai_1 _3323_ (.B1(net853),
    .Y(_0541_),
    .A1(net647),
    .A2(_0540_));
 sg13g2_a21oi_1 _3324_ (.A1(_1377_),
    .A2(net647),
    .Y(_0066_),
    .B1(_0541_));
 sg13g2_o21ai_1 _3325_ (.B1(_0419_),
    .Y(_0542_),
    .A1(net786),
    .A2(_1393_));
 sg13g2_o21ai_1 _3326_ (.B1(net850),
    .Y(_0543_),
    .A1(net647),
    .A2(_0542_));
 sg13g2_a21oi_1 _3327_ (.A1(_1376_),
    .A2(net647),
    .Y(_0067_),
    .B1(_0543_));
 sg13g2_a21o_1 _3328_ (.A2(_0426_),
    .A1(net788),
    .B1(_0430_),
    .X(_0544_));
 sg13g2_o21ai_1 _3329_ (.B1(net850),
    .Y(_0545_),
    .A1(net647),
    .A2(_0544_));
 sg13g2_a21oi_1 _3330_ (.A1(_1375_),
    .A2(net647),
    .Y(_0068_),
    .B1(_0545_));
 sg13g2_nand2_1 _3331_ (.Y(_0546_),
    .A(net692),
    .B(_1417_));
 sg13g2_nor3_2 _3332_ (.A(net1),
    .B(net826),
    .C(net672),
    .Y(_0547_));
 sg13g2_mux4_1 _3333_ (.S0(net827),
    .A0(\collatz.orbit_len[0] ),
    .A1(\collatz.orbit_len[8] ),
    .A2(\collatz.path_record_h16[0] ),
    .A3(\collatz.path_record_h16[8] ),
    .S1(net5),
    .X(_0548_));
 sg13g2_a22oi_1 _3334_ (.Y(_0549_),
    .B1(_0547_),
    .B2(_0548_),
    .A2(_0546_),
    .A1(net240));
 sg13g2_nor2_1 _3335_ (.A(net822),
    .B(_0549_),
    .Y(_0069_));
 sg13g2_mux4_1 _3336_ (.S0(net827),
    .A0(\collatz.orbit_len[1] ),
    .A1(\collatz.orbit_len[9] ),
    .A2(\collatz.path_record_h16[1] ),
    .A3(\collatz.path_record_h16[9] ),
    .S1(net5),
    .X(_0550_));
 sg13g2_a22oi_1 _3337_ (.Y(_0551_),
    .B1(_0547_),
    .B2(_0550_),
    .A2(net672),
    .A1(net245));
 sg13g2_nor2_1 _3338_ (.A(net822),
    .B(_0551_),
    .Y(_0070_));
 sg13g2_mux4_1 _3339_ (.S0(net827),
    .A0(\collatz.orbit_len[2] ),
    .A1(\collatz.orbit_len[10] ),
    .A2(\collatz.path_record_h16[2] ),
    .A3(\collatz.path_record_h16[10] ),
    .S1(net5),
    .X(_0552_));
 sg13g2_a22oi_1 _3340_ (.Y(_0553_),
    .B1(_0547_),
    .B2(_0552_),
    .A2(net672),
    .A1(net250));
 sg13g2_nor2_1 _3341_ (.A(net822),
    .B(_0553_),
    .Y(_0071_));
 sg13g2_mux4_1 _3342_ (.S0(net827),
    .A0(\collatz.orbit_len[3] ),
    .A1(\collatz.orbit_len[11] ),
    .A2(\collatz.path_record_h16[3] ),
    .A3(\collatz.path_record_h16[11] ),
    .S1(net5),
    .X(_0554_));
 sg13g2_a22oi_1 _3343_ (.Y(_0555_),
    .B1(_0547_),
    .B2(_0554_),
    .A2(net672),
    .A1(net235));
 sg13g2_nor2_1 _3344_ (.A(net822),
    .B(_0555_),
    .Y(_0072_));
 sg13g2_mux4_1 _3345_ (.S0(net827),
    .A0(net342),
    .A1(\collatz.orbit_len[12] ),
    .A2(\collatz.path_record_h16[4] ),
    .A3(\collatz.path_record_h16[12] ),
    .S1(net5),
    .X(_0556_));
 sg13g2_a22oi_1 _3346_ (.Y(_0557_),
    .B1(_0547_),
    .B2(_0556_),
    .A2(net672),
    .A1(net223));
 sg13g2_nor2_1 _3347_ (.A(net822),
    .B(_0557_),
    .Y(_0073_));
 sg13g2_mux4_1 _3348_ (.S0(net827),
    .A0(net331),
    .A1(net215),
    .A2(\collatz.path_record_h16[5] ),
    .A3(\collatz.path_record_h16[13] ),
    .S1(net5),
    .X(_0558_));
 sg13g2_a22oi_1 _3349_ (.Y(_0559_),
    .B1(_0547_),
    .B2(_0558_),
    .A2(net672),
    .A1(net237));
 sg13g2_nor2_1 _3350_ (.A(net821),
    .B(_0559_),
    .Y(_0074_));
 sg13g2_mux4_1 _3351_ (.S0(net827),
    .A0(net224),
    .A1(net338),
    .A2(\collatz.path_record_h16[6] ),
    .A3(\collatz.path_record_h16[14] ),
    .S1(net5),
    .X(_0560_));
 sg13g2_a22oi_1 _3352_ (.Y(_0561_),
    .B1(_0547_),
    .B2(_0560_),
    .A2(net672),
    .A1(net233));
 sg13g2_nor2_1 _3353_ (.A(net821),
    .B(_0561_),
    .Y(_0075_));
 sg13g2_mux4_1 _3354_ (.S0(net827),
    .A0(\collatz.orbit_len[7] ),
    .A1(\collatz.orbit_len[15] ),
    .A2(\collatz.path_record_h16[7] ),
    .A3(\collatz.path_record_h16[15] ),
    .S1(net5),
    .X(_0562_));
 sg13g2_a22oi_1 _3355_ (.Y(_0563_),
    .B1(_0547_),
    .B2(_0562_),
    .A2(net672),
    .A1(net222));
 sg13g2_nor2_1 _3356_ (.A(net822),
    .B(_0563_),
    .Y(_0076_));
 sg13g2_nor2_2 _3357_ (.A(_1417_),
    .B(net4),
    .Y(_0564_));
 sg13g2_and2_1 _3358_ (.A(_1512_),
    .B(_0564_),
    .X(_0565_));
 sg13g2_nor2_2 _3359_ (.A(net651),
    .B(net671),
    .Y(_0566_));
 sg13g2_a22oi_1 _3360_ (.Y(_0567_),
    .B1(_0566_),
    .B2(\collatz.iter[1] ),
    .A2(_0565_),
    .A1(net843));
 sg13g2_nor2_1 _3361_ (.A(net798),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_nand3_1 _3362_ (.B(\collatz.iter[2] ),
    .C(net681),
    .A(net798),
    .Y(_0569_));
 sg13g2_o21ai_1 _3363_ (.B1(_0569_),
    .Y(_0570_),
    .A1(_0009_),
    .A2(net207));
 sg13g2_nor2_1 _3364_ (.A(_0568_),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_nor3_1 _3365_ (.A(\collatz.iter[1] ),
    .B(_0009_),
    .C(net207),
    .Y(_0572_));
 sg13g2_nor3_1 _3366_ (.A(net824),
    .B(_0571_),
    .C(net208),
    .Y(_0077_));
 sg13g2_nand2_1 _3367_ (.Y(_0573_),
    .A(net756),
    .B(_0566_));
 sg13g2_a21oi_1 _3368_ (.A1(net845),
    .A2(net671),
    .Y(_0574_),
    .B1(net798));
 sg13g2_a221oi_1 _3369_ (.B2(_0574_),
    .C1(net824),
    .B1(_0573_),
    .A1(net798),
    .Y(_0078_),
    .A2(_1451_));
 sg13g2_a22oi_1 _3370_ (.Y(_0575_),
    .B1(_0566_),
    .B2(net323),
    .A2(net671),
    .A1(net841));
 sg13g2_a21oi_1 _3371_ (.A1(\collatz.iter[1] ),
    .A2(\collatz.iter[2] ),
    .Y(_0576_),
    .B1(_1722_));
 sg13g2_o21ai_1 _3372_ (.B1(net798),
    .Y(_0577_),
    .A1(net711),
    .A2(net757));
 sg13g2_or2_1 _3373_ (.X(_0578_),
    .B(_0577_),
    .A(_0576_));
 sg13g2_o21ai_1 _3374_ (.B1(_0578_),
    .Y(_0579_),
    .A1(net798),
    .A2(_0575_));
 sg13g2_and2_1 _3375_ (.A(net853),
    .B(_0579_),
    .X(_0079_));
 sg13g2_nand2_1 _3376_ (.Y(_0580_),
    .A(net711),
    .B(_0566_));
 sg13g2_a21oi_1 _3377_ (.A1(net839),
    .A2(net671),
    .Y(_0581_),
    .B1(net799));
 sg13g2_xor2_1 _3378_ (.B(\collatz.iter[2] ),
    .A(net711),
    .X(_0582_));
 sg13g2_o21ai_1 _3379_ (.B1(net757),
    .Y(_0583_),
    .A1(\collatz.iter[1] ),
    .A2(net711));
 sg13g2_a21oi_1 _3380_ (.A1(\collatz.iter[1] ),
    .A2(_0582_),
    .Y(_0584_),
    .B1(_0583_));
 sg13g2_a21oi_1 _3381_ (.A1(net291),
    .A2(net682),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_a221oi_1 _3382_ (.B2(net799),
    .C1(net824),
    .B1(_0585_),
    .A1(_0580_),
    .Y(_0080_),
    .A2(_0581_));
 sg13g2_nor2b_1 _3383_ (.A(_1729_),
    .B_N(_1724_),
    .Y(_0586_));
 sg13g2_a22oi_1 _3384_ (.Y(_0587_),
    .B1(_0566_),
    .B2(\collatz.iter[4] ),
    .A2(net671),
    .A1(net837));
 sg13g2_xor2_1 _3385_ (.B(_1729_),
    .A(_1724_),
    .X(_0588_));
 sg13g2_o21ai_1 _3386_ (.B1(net799),
    .Y(_0589_),
    .A1(\collatz.iter[5] ),
    .A2(net756));
 sg13g2_a21o_1 _3387_ (.A2(_0588_),
    .A1(net756),
    .B1(_0589_),
    .X(_0590_));
 sg13g2_o21ai_1 _3388_ (.B1(_0590_),
    .Y(_0591_),
    .A1(net799),
    .A2(_0587_));
 sg13g2_and2_1 _3389_ (.A(net851),
    .B(_0591_),
    .X(_0081_));
 sg13g2_a22oi_1 _3390_ (.Y(_0592_),
    .B1(_0566_),
    .B2(\collatz.iter[5] ),
    .A2(net671),
    .A1(net835));
 sg13g2_a21oi_1 _3391_ (.A1(\collatz.iter[4] ),
    .A2(net711),
    .Y(_0593_),
    .B1(_0586_));
 sg13g2_xnor2_1 _3392_ (.Y(_0594_),
    .A(_1728_),
    .B(_0593_));
 sg13g2_a21oi_1 _3393_ (.A1(net756),
    .A2(_0594_),
    .Y(_0595_),
    .B1(net694));
 sg13g2_o21ai_1 _3394_ (.B1(_0595_),
    .Y(_0596_),
    .A1(\collatz.iter[6] ),
    .A2(net756));
 sg13g2_o21ai_1 _3395_ (.B1(_0596_),
    .Y(_0597_),
    .A1(net798),
    .A2(_0592_));
 sg13g2_and2_1 _3396_ (.A(net851),
    .B(_0597_),
    .X(_0082_));
 sg13g2_a22oi_1 _3397_ (.Y(_0598_),
    .B1(_0566_),
    .B2(\collatz.iter[6] ),
    .A2(net671),
    .A1(net833));
 sg13g2_nor2_1 _3398_ (.A(_1732_),
    .B(_0586_),
    .Y(_0599_));
 sg13g2_nor3_1 _3399_ (.A(_1441_),
    .B(_1725_),
    .C(_0599_),
    .Y(_0600_));
 sg13g2_o21ai_1 _3400_ (.B1(_1725_),
    .Y(_0601_),
    .A1(_1441_),
    .A2(_0599_));
 sg13g2_nor2b_1 _3401_ (.A(_0600_),
    .B_N(_0601_),
    .Y(_0602_));
 sg13g2_nand2_1 _3402_ (.Y(_0603_),
    .A(net284),
    .B(net682));
 sg13g2_a21oi_1 _3403_ (.A1(net756),
    .A2(_0602_),
    .Y(_0604_),
    .B1(net693));
 sg13g2_a221oi_1 _3404_ (.B2(_0604_),
    .C1(net824),
    .B1(_0603_),
    .A1(net693),
    .Y(_0083_),
    .A2(_0598_));
 sg13g2_a22oi_1 _3405_ (.Y(_0605_),
    .B1(_0566_),
    .B2(\collatz.iter[7] ),
    .A2(net671),
    .A1(net831));
 sg13g2_a21oi_1 _3406_ (.A1(\collatz.iter[6] ),
    .A2(\collatz.iter[5] ),
    .Y(_0606_),
    .B1(_0600_));
 sg13g2_xnor2_1 _3407_ (.Y(_0607_),
    .A(_1726_),
    .B(_0606_));
 sg13g2_a21oi_1 _3408_ (.A1(net756),
    .A2(_0607_),
    .Y(_0608_),
    .B1(net693));
 sg13g2_o21ai_1 _3409_ (.B1(_0608_),
    .Y(_0609_),
    .A1(\collatz.iter[8] ),
    .A2(net757));
 sg13g2_o21ai_1 _3410_ (.B1(_0609_),
    .Y(_0610_),
    .A1(net798),
    .A2(_0605_));
 sg13g2_and2_1 _3411_ (.A(net851),
    .B(_0610_),
    .X(_0084_));
 sg13g2_a21oi_2 _3412_ (.B1(net651),
    .Y(_0611_),
    .A2(_0564_),
    .A1(_0348_));
 sg13g2_nand2_1 _3413_ (.Y(_0612_),
    .A(\collatz.iter[8] ),
    .B(_0611_));
 sg13g2_nand3_1 _3414_ (.B(net662),
    .C(net677),
    .A(net845),
    .Y(_0613_));
 sg13g2_a21oi_1 _3415_ (.A1(_0612_),
    .A2(_0613_),
    .Y(_0614_),
    .B1(net795));
 sg13g2_nor2_1 _3416_ (.A(_1735_),
    .B(_1740_),
    .Y(_0615_));
 sg13g2_xnor2_1 _3417_ (.Y(_0616_),
    .A(_1735_),
    .B(_1740_));
 sg13g2_o21ai_1 _3418_ (.B1(net795),
    .Y(_0617_),
    .A1(\collatz.iter[9] ),
    .A2(net754));
 sg13g2_a21oi_1 _3419_ (.A1(net754),
    .A2(_0616_),
    .Y(_0618_),
    .B1(_0617_));
 sg13g2_o21ai_1 _3420_ (.B1(net852),
    .Y(_0619_),
    .A1(_0614_),
    .A2(_0618_));
 sg13g2_inv_1 _3421_ (.Y(_0085_),
    .A(_0619_));
 sg13g2_nand2_1 _3422_ (.Y(_0620_),
    .A(\collatz.iter[9] ),
    .B(_0611_));
 sg13g2_nand3_1 _3423_ (.B(net662),
    .C(net678),
    .A(net843),
    .Y(_0621_));
 sg13g2_a21oi_1 _3424_ (.A1(_0620_),
    .A2(_0621_),
    .Y(_0622_),
    .B1(net795));
 sg13g2_a21oi_1 _3425_ (.A1(\collatz.iter[8] ),
    .A2(\collatz.iter[7] ),
    .Y(_0623_),
    .B1(_0615_));
 sg13g2_xor2_1 _3426_ (.B(_0623_),
    .A(_1742_),
    .X(_0624_));
 sg13g2_o21ai_1 _3427_ (.B1(net797),
    .Y(_0625_),
    .A1(\collatz.iter[10] ),
    .A2(net753));
 sg13g2_a21oi_1 _3428_ (.A1(net753),
    .A2(_0624_),
    .Y(_0626_),
    .B1(_0625_));
 sg13g2_o21ai_1 _3429_ (.B1(net852),
    .Y(_0627_),
    .A1(_0622_),
    .A2(_0626_));
 sg13g2_inv_1 _3430_ (.Y(_0086_),
    .A(_0627_));
 sg13g2_nand2_1 _3431_ (.Y(_0628_),
    .A(\collatz.iter[10] ),
    .B(_0611_));
 sg13g2_nand3_1 _3432_ (.B(net662),
    .C(net678),
    .A(net841),
    .Y(_0629_));
 sg13g2_a21oi_1 _3433_ (.A1(_0628_),
    .A2(_0629_),
    .Y(_0630_),
    .B1(net795));
 sg13g2_nor2b_1 _3434_ (.A(_0615_),
    .B_N(_1745_),
    .Y(_0631_));
 sg13g2_nor3_1 _3435_ (.A(_1447_),
    .B(_1737_),
    .C(_0631_),
    .Y(_0632_));
 sg13g2_o21ai_1 _3436_ (.B1(_1737_),
    .Y(_0633_),
    .A1(_1447_),
    .A2(_0631_));
 sg13g2_nand2b_1 _3437_ (.Y(_0634_),
    .B(_0633_),
    .A_N(_0632_));
 sg13g2_o21ai_1 _3438_ (.B1(net795),
    .Y(_0635_),
    .A1(\collatz.iter[11] ),
    .A2(net753));
 sg13g2_a21oi_1 _3439_ (.A1(net753),
    .A2(_0634_),
    .Y(_0636_),
    .B1(_0635_));
 sg13g2_o21ai_1 _3440_ (.B1(net852),
    .Y(_0637_),
    .A1(_0630_),
    .A2(_0636_));
 sg13g2_inv_1 _3441_ (.Y(_0087_),
    .A(_0637_));
 sg13g2_nand2_1 _3442_ (.Y(_0638_),
    .A(\collatz.iter[11] ),
    .B(_0611_));
 sg13g2_nand3_1 _3443_ (.B(net662),
    .C(net677),
    .A(net839),
    .Y(_0639_));
 sg13g2_a21oi_1 _3444_ (.A1(_0638_),
    .A2(_0639_),
    .Y(_0640_),
    .B1(net795));
 sg13g2_nor2_1 _3445_ (.A(_1736_),
    .B(_0632_),
    .Y(_0641_));
 sg13g2_xnor2_1 _3446_ (.Y(_0642_),
    .A(_1738_),
    .B(_0641_));
 sg13g2_o21ai_1 _3447_ (.B1(net795),
    .Y(_0643_),
    .A1(\collatz.iter[12] ),
    .A2(net754));
 sg13g2_a21oi_1 _3448_ (.A1(net754),
    .A2(_0642_),
    .Y(_0644_),
    .B1(_0643_));
 sg13g2_o21ai_1 _3449_ (.B1(net851),
    .Y(_0645_),
    .A1(_0640_),
    .A2(_0644_));
 sg13g2_inv_1 _3450_ (.Y(_0088_),
    .A(_0645_));
 sg13g2_nand2_1 _3451_ (.Y(_0646_),
    .A(\collatz.iter[12] ),
    .B(_0611_));
 sg13g2_nand3_1 _3452_ (.B(net662),
    .C(net677),
    .A(net837),
    .Y(_0647_));
 sg13g2_a21oi_1 _3453_ (.A1(_0646_),
    .A2(_0647_),
    .Y(_0648_),
    .B1(net796));
 sg13g2_nor3_1 _3454_ (.A(_1714_),
    .B(_1744_),
    .C(_1748_),
    .Y(_0649_));
 sg13g2_o21ai_1 _3455_ (.B1(_1714_),
    .Y(_0650_),
    .A1(_1744_),
    .A2(_1748_));
 sg13g2_nand2b_1 _3456_ (.Y(_0651_),
    .B(_0650_),
    .A_N(_0649_));
 sg13g2_o21ai_1 _3457_ (.B1(net796),
    .Y(_0652_),
    .A1(\collatz.iter[13] ),
    .A2(net754));
 sg13g2_a21oi_1 _3458_ (.A1(net755),
    .A2(_0651_),
    .Y(_0653_),
    .B1(_0652_));
 sg13g2_o21ai_1 _3459_ (.B1(net851),
    .Y(_0654_),
    .A1(_0648_),
    .A2(_0653_));
 sg13g2_inv_1 _3460_ (.Y(_0089_),
    .A(_0654_));
 sg13g2_nand2_1 _3461_ (.Y(_0655_),
    .A(\collatz.iter[13] ),
    .B(_0611_));
 sg13g2_nand3_1 _3462_ (.B(net662),
    .C(net677),
    .A(net835),
    .Y(_0656_));
 sg13g2_a21oi_1 _3463_ (.A1(_0655_),
    .A2(_0656_),
    .Y(_0657_),
    .B1(net796));
 sg13g2_o21ai_1 _3464_ (.B1(_0650_),
    .Y(_0658_),
    .A1(_1411_),
    .A2(_1412_));
 sg13g2_xnor2_1 _3465_ (.Y(_0659_),
    .A(_1715_),
    .B(_0658_));
 sg13g2_o21ai_1 _3466_ (.B1(net796),
    .Y(_0660_),
    .A1(\collatz.iter[14] ),
    .A2(net755));
 sg13g2_a21oi_1 _3467_ (.A1(net755),
    .A2(_0659_),
    .Y(_0661_),
    .B1(_0660_));
 sg13g2_o21ai_1 _3468_ (.B1(net851),
    .Y(_0662_),
    .A1(_0657_),
    .A2(_0661_));
 sg13g2_inv_1 _3469_ (.Y(_0090_),
    .A(_0662_));
 sg13g2_nand2_1 _3470_ (.Y(_0663_),
    .A(\collatz.iter[14] ),
    .B(_0611_));
 sg13g2_nand3_1 _3471_ (.B(net662),
    .C(net677),
    .A(net833),
    .Y(_0664_));
 sg13g2_a21oi_1 _3472_ (.A1(_0663_),
    .A2(_0664_),
    .Y(_0665_),
    .B1(net797));
 sg13g2_a22oi_1 _3473_ (.Y(_0666_),
    .B1(_1718_),
    .B2(_0650_),
    .A2(_1411_),
    .A1(_1410_));
 sg13g2_nor2b_1 _3474_ (.A(_1711_),
    .B_N(_0666_),
    .Y(_0667_));
 sg13g2_xor2_1 _3475_ (.B(_0666_),
    .A(_1711_),
    .X(_0668_));
 sg13g2_o21ai_1 _3476_ (.B1(net797),
    .Y(_0669_),
    .A1(\collatz.iter[15] ),
    .A2(net754));
 sg13g2_a21oi_1 _3477_ (.A1(net755),
    .A2(_0668_),
    .Y(_0670_),
    .B1(_0669_));
 sg13g2_o21ai_1 _3478_ (.B1(net851),
    .Y(_0671_),
    .A1(_0665_),
    .A2(_0670_));
 sg13g2_inv_1 _3479_ (.Y(_0091_),
    .A(_0671_));
 sg13g2_a22oi_1 _3480_ (.Y(_0672_),
    .B1(_0611_),
    .B2(\collatz.iter[15] ),
    .A2(_0429_),
    .A1(_1515_));
 sg13g2_a21oi_1 _3481_ (.A1(\collatz.iter[14] ),
    .A2(\collatz.iter[13] ),
    .Y(_0673_),
    .B1(_0667_));
 sg13g2_xnor2_1 _3482_ (.Y(_0674_),
    .A(_1712_),
    .B(_0673_));
 sg13g2_a21oi_1 _3483_ (.A1(net754),
    .A2(_0674_),
    .Y(_0675_),
    .B1(net693));
 sg13g2_o21ai_1 _3484_ (.B1(_0675_),
    .Y(_0676_),
    .A1(\collatz.iter[16] ),
    .A2(net754));
 sg13g2_o21ai_1 _3485_ (.B1(_0676_),
    .Y(_0677_),
    .A1(net795),
    .A2(_0672_));
 sg13g2_and2_1 _3486_ (.A(net851),
    .B(_0677_),
    .X(_0092_));
 sg13g2_nand2_1 _3487_ (.Y(_0678_),
    .A(_1751_),
    .B(_1764_));
 sg13g2_nor2_1 _3488_ (.A(_1751_),
    .B(_1764_),
    .Y(_0679_));
 sg13g2_nand2_1 _3489_ (.Y(_0680_),
    .A(net751),
    .B(_0678_));
 sg13g2_nor2_1 _3490_ (.A(_0679_),
    .B(_0680_),
    .Y(_0681_));
 sg13g2_o21ai_1 _3491_ (.B1(net800),
    .Y(_0682_),
    .A1(_1406_),
    .A2(net752));
 sg13g2_and2_1 _3492_ (.A(_1513_),
    .B(_0564_),
    .X(_0683_));
 sg13g2_nor3_2 _3493_ (.A(_1418_),
    .B(net826),
    .C(net828),
    .Y(_0684_));
 sg13g2_nand2_1 _3494_ (.Y(_0685_),
    .A(net669),
    .B(_0684_));
 sg13g2_and2_1 _3495_ (.A(net845),
    .B(net676),
    .X(_0686_));
 sg13g2_a22oi_1 _3496_ (.Y(_0687_),
    .B1(_0686_),
    .B2(net668),
    .A2(_0685_),
    .A1(\collatz.iter[16] ));
 sg13g2_o21ai_1 _3497_ (.B1(net852),
    .Y(_0688_),
    .A1(_0681_),
    .A2(_0682_));
 sg13g2_a21oi_1 _3498_ (.A1(net693),
    .A2(_0687_),
    .Y(_0093_),
    .B1(_0688_));
 sg13g2_nor2b_2 _3499_ (.A(net651),
    .B_N(_0685_),
    .Y(_0689_));
 sg13g2_and2_1 _3500_ (.A(net843),
    .B(net676),
    .X(_0690_));
 sg13g2_a22oi_1 _3501_ (.Y(_0691_),
    .B1(_0690_),
    .B2(net668),
    .A2(_0689_),
    .A1(\collatz.iter[17] ));
 sg13g2_o21ai_1 _3502_ (.B1(_0678_),
    .Y(_0692_),
    .A1(_1407_),
    .A2(_1408_));
 sg13g2_xnor2_1 _3503_ (.Y(_0693_),
    .A(_1765_),
    .B(_0692_));
 sg13g2_a21oi_1 _3504_ (.A1(net751),
    .A2(_0693_),
    .Y(_0694_),
    .B1(net693));
 sg13g2_o21ai_1 _3505_ (.B1(_0694_),
    .Y(_0695_),
    .A1(\collatz.iter[18] ),
    .A2(net752));
 sg13g2_o21ai_1 _3506_ (.B1(_0695_),
    .Y(_0696_),
    .A1(net800),
    .A2(_0691_));
 sg13g2_and2_1 _3507_ (.A(net852),
    .B(_0696_),
    .X(_0094_));
 sg13g2_and2_1 _3508_ (.A(net841),
    .B(net676),
    .X(_0697_));
 sg13g2_a22oi_1 _3509_ (.Y(_0698_),
    .B1(_0697_),
    .B2(net668),
    .A2(_0689_),
    .A1(\collatz.iter[18] ));
 sg13g2_a22oi_1 _3510_ (.Y(_0699_),
    .B1(_1768_),
    .B2(_0678_),
    .A2(_1407_),
    .A1(_1406_));
 sg13g2_xnor2_1 _3511_ (.Y(_0700_),
    .A(_1762_),
    .B(_0699_));
 sg13g2_o21ai_1 _3512_ (.B1(net800),
    .Y(_0701_),
    .A1(\collatz.iter[19] ),
    .A2(net752));
 sg13g2_a21o_1 _3513_ (.A2(_0700_),
    .A1(net751),
    .B1(_0701_),
    .X(_0702_));
 sg13g2_o21ai_1 _3514_ (.B1(_0702_),
    .Y(_0703_),
    .A1(net800),
    .A2(_0698_));
 sg13g2_and2_1 _3515_ (.A(net852),
    .B(_0703_),
    .X(_0095_));
 sg13g2_and2_1 _3516_ (.A(net839),
    .B(net676),
    .X(_0704_));
 sg13g2_a22oi_1 _3517_ (.Y(_0705_),
    .B1(_0704_),
    .B2(net668),
    .A2(_0689_),
    .A1(\collatz.iter[19] ));
 sg13g2_a21oi_1 _3518_ (.A1(_1762_),
    .A2(_0699_),
    .Y(_0706_),
    .B1(_1761_));
 sg13g2_xor2_1 _3519_ (.B(_0706_),
    .A(_1763_),
    .X(_0707_));
 sg13g2_a21oi_1 _3520_ (.A1(net752),
    .A2(_0707_),
    .Y(_0708_),
    .B1(net693));
 sg13g2_o21ai_1 _3521_ (.B1(_0708_),
    .Y(_0709_),
    .A1(\collatz.iter[20] ),
    .A2(net751));
 sg13g2_o21ai_1 _3522_ (.B1(_0709_),
    .Y(_0710_),
    .A1(net800),
    .A2(_0705_));
 sg13g2_and2_1 _3523_ (.A(net852),
    .B(_0710_),
    .X(_0096_));
 sg13g2_and2_1 _3524_ (.A(net837),
    .B(net676),
    .X(_0711_));
 sg13g2_a22oi_1 _3525_ (.Y(_0712_),
    .B1(_0711_),
    .B2(net668),
    .A2(_0689_),
    .A1(\collatz.iter[20] ));
 sg13g2_or2_1 _3526_ (.X(_0713_),
    .B(_1766_),
    .A(_1752_));
 sg13g2_nand3_1 _3527_ (.B(_1770_),
    .C(_0713_),
    .A(_1769_),
    .Y(_0714_));
 sg13g2_nand2_1 _3528_ (.Y(_0715_),
    .A(_1758_),
    .B(_0714_));
 sg13g2_xnor2_1 _3529_ (.Y(_0716_),
    .A(_1758_),
    .B(_0714_));
 sg13g2_o21ai_1 _3530_ (.B1(net793),
    .Y(_0717_),
    .A1(\collatz.iter[21] ),
    .A2(net751));
 sg13g2_a21o_1 _3531_ (.A2(_0716_),
    .A1(net751),
    .B1(_0717_),
    .X(_0718_));
 sg13g2_o21ai_1 _3532_ (.B1(_0718_),
    .Y(_0719_),
    .A1(net800),
    .A2(_0712_));
 sg13g2_and2_1 _3533_ (.A(net852),
    .B(_0719_),
    .X(_0097_));
 sg13g2_and2_1 _3534_ (.A(net835),
    .B(net676),
    .X(_0720_));
 sg13g2_a22oi_1 _3535_ (.Y(_0721_),
    .B1(_0720_),
    .B2(net668),
    .A2(_0689_),
    .A1(\collatz.iter[21] ));
 sg13g2_nand2_1 _3536_ (.Y(_0722_),
    .A(_1757_),
    .B(_0715_));
 sg13g2_xnor2_1 _3537_ (.Y(_0723_),
    .A(_1759_),
    .B(_0722_));
 sg13g2_a21oi_1 _3538_ (.A1(net751),
    .A2(_0723_),
    .Y(_0724_),
    .B1(net693));
 sg13g2_o21ai_1 _3539_ (.B1(_0724_),
    .Y(_0725_),
    .A1(\collatz.iter[22] ),
    .A2(net751));
 sg13g2_o21ai_1 _3540_ (.B1(_0725_),
    .Y(_0726_),
    .A1(net793),
    .A2(_0721_));
 sg13g2_and2_1 _3541_ (.A(net849),
    .B(_0726_),
    .X(_0098_));
 sg13g2_and2_1 _3542_ (.A(net833),
    .B(net676),
    .X(_0727_));
 sg13g2_a22oi_1 _3543_ (.Y(_0728_),
    .B1(_0727_),
    .B2(net668),
    .A2(_0689_),
    .A1(\collatz.iter[22] ));
 sg13g2_a21oi_1 _3544_ (.A1(_1773_),
    .A2(_0715_),
    .Y(_0729_),
    .B1(_1428_));
 sg13g2_xnor2_1 _3545_ (.Y(_0730_),
    .A(_1754_),
    .B(_0729_));
 sg13g2_o21ai_1 _3546_ (.B1(net793),
    .Y(_0731_),
    .A1(\collatz.iter[23] ),
    .A2(net747));
 sg13g2_a21o_1 _3547_ (.A2(_0730_),
    .A1(net747),
    .B1(_0731_),
    .X(_0732_));
 sg13g2_o21ai_1 _3548_ (.B1(_0732_),
    .Y(_0733_),
    .A1(net792),
    .A2(_0728_));
 sg13g2_and2_1 _3549_ (.A(net849),
    .B(_0733_),
    .X(_0099_));
 sg13g2_and2_1 _3550_ (.A(net830),
    .B(net676),
    .X(_0734_));
 sg13g2_a22oi_1 _3551_ (.Y(_0735_),
    .B1(_0734_),
    .B2(net668),
    .A2(_0689_),
    .A1(\collatz.iter[23] ));
 sg13g2_or2_1 _3552_ (.X(_0736_),
    .B(_0735_),
    .A(net793));
 sg13g2_a21oi_1 _3553_ (.A1(_1754_),
    .A2(_0729_),
    .Y(_0737_),
    .B1(_1753_));
 sg13g2_xor2_1 _3554_ (.B(_0737_),
    .A(_1755_),
    .X(_0738_));
 sg13g2_a21oi_1 _3555_ (.A1(net746),
    .A2(_0738_),
    .Y(_0739_),
    .B1(net690));
 sg13g2_o21ai_1 _3556_ (.B1(_0739_),
    .Y(_0740_),
    .A1(net308),
    .A2(net746));
 sg13g2_a21oi_1 _3557_ (.A1(_0736_),
    .A2(_0740_),
    .Y(_0100_),
    .B1(net819));
 sg13g2_nor3_2 _3558_ (.A(_1418_),
    .B(net826),
    .C(_1419_),
    .Y(_0741_));
 sg13g2_a21oi_2 _3559_ (.B1(net651),
    .Y(_0742_),
    .A2(net675),
    .A1(net669));
 sg13g2_and2_1 _3560_ (.A(net845),
    .B(_0741_),
    .X(_0743_));
 sg13g2_a22oi_1 _3561_ (.Y(_0744_),
    .B1(_0743_),
    .B2(net669),
    .A2(_0742_),
    .A1(\collatz.iter[24] ));
 sg13g2_a21o_2 _3562_ (.A2(_1767_),
    .A1(_1751_),
    .B1(_1775_),
    .X(_0745_));
 sg13g2_nand2_1 _3563_ (.Y(_0746_),
    .A(_1698_),
    .B(_0745_));
 sg13g2_xnor2_1 _3564_ (.Y(_0747_),
    .A(_1698_),
    .B(_0745_));
 sg13g2_o21ai_1 _3565_ (.B1(net791),
    .Y(_0748_),
    .A1(net710),
    .A2(net743));
 sg13g2_a21o_1 _3566_ (.A2(_0747_),
    .A1(net744),
    .B1(_0748_),
    .X(_0749_));
 sg13g2_o21ai_1 _3567_ (.B1(_0749_),
    .Y(_0750_),
    .A1(net791),
    .A2(_0744_));
 sg13g2_and2_1 _3568_ (.A(net849),
    .B(_0750_),
    .X(_0101_));
 sg13g2_and2_1 _3569_ (.A(net843),
    .B(net675),
    .X(_0751_));
 sg13g2_a22oi_1 _3570_ (.Y(_0752_),
    .B1(_0751_),
    .B2(net669),
    .A2(_0742_),
    .A1(net710));
 sg13g2_or2_1 _3571_ (.X(_0753_),
    .B(_0752_),
    .A(net794));
 sg13g2_nand2_1 _3572_ (.Y(_0754_),
    .A(_1697_),
    .B(_0746_));
 sg13g2_xnor2_1 _3573_ (.Y(_0755_),
    .A(_1699_),
    .B(_0754_));
 sg13g2_a21oi_1 _3574_ (.A1(_1405_),
    .A2(net681),
    .Y(_0756_),
    .B1(net690));
 sg13g2_o21ai_1 _3575_ (.B1(_0756_),
    .Y(_0757_),
    .A1(net681),
    .A2(_0755_));
 sg13g2_a21oi_1 _3576_ (.A1(_0753_),
    .A2(_0757_),
    .Y(_0102_),
    .B1(net818));
 sg13g2_and2_1 _3577_ (.A(net840),
    .B(_0741_),
    .X(_0758_));
 sg13g2_a22oi_1 _3578_ (.Y(_0759_),
    .B1(_0758_),
    .B2(net669),
    .A2(_0742_),
    .A1(\collatz.iter[26] ));
 sg13g2_a21oi_1 _3579_ (.A1(_1707_),
    .A2(_0746_),
    .Y(_0760_),
    .B1(_1452_));
 sg13g2_xnor2_1 _3580_ (.Y(_0761_),
    .A(_1694_),
    .B(_0760_));
 sg13g2_o21ai_1 _3581_ (.B1(net791),
    .Y(_0762_),
    .A1(\collatz.iter[27] ),
    .A2(net743));
 sg13g2_a21o_1 _3582_ (.A2(_0761_),
    .A1(net743),
    .B1(_0762_),
    .X(_0763_));
 sg13g2_o21ai_1 _3583_ (.B1(_0763_),
    .Y(_0764_),
    .A1(net791),
    .A2(_0759_));
 sg13g2_and2_1 _3584_ (.A(net849),
    .B(_0764_),
    .X(_0103_));
 sg13g2_and2_1 _3585_ (.A(net838),
    .B(net675),
    .X(_0765_));
 sg13g2_a22oi_1 _3586_ (.Y(_0766_),
    .B1(_0765_),
    .B2(net669),
    .A2(_0742_),
    .A1(\collatz.iter[27] ));
 sg13g2_or2_1 _3587_ (.X(_0767_),
    .B(_0766_),
    .A(net779));
 sg13g2_a21oi_1 _3588_ (.A1(_1694_),
    .A2(_0760_),
    .Y(_0768_),
    .B1(_1693_));
 sg13g2_xnor2_1 _3589_ (.Y(_0769_),
    .A(_1696_),
    .B(_0768_));
 sg13g2_a21oi_1 _3590_ (.A1(net743),
    .A2(_0769_),
    .Y(_0770_),
    .B1(net690));
 sg13g2_o21ai_1 _3591_ (.B1(_0770_),
    .Y(_0771_),
    .A1(net297),
    .A2(net735));
 sg13g2_a21oi_1 _3592_ (.A1(_0767_),
    .A2(_0771_),
    .Y(_0104_),
    .B1(net813));
 sg13g2_and2_1 _3593_ (.A(net836),
    .B(net675),
    .X(_0772_));
 sg13g2_a22oi_1 _3594_ (.Y(_0773_),
    .B1(_0772_),
    .B2(net669),
    .A2(_0742_),
    .A1(net340));
 sg13g2_a21oi_2 _3595_ (.B1(_1710_),
    .Y(_0774_),
    .A2(_0745_),
    .A1(_1701_));
 sg13g2_or2_1 _3596_ (.X(_0775_),
    .B(_0774_),
    .A(_1691_));
 sg13g2_xnor2_1 _3597_ (.Y(_0776_),
    .A(_1691_),
    .B(_0774_));
 sg13g2_o21ai_1 _3598_ (.B1(net779),
    .Y(_0777_),
    .A1(\collatz.iter[29] ),
    .A2(net735));
 sg13g2_a21o_1 _3599_ (.A2(_0776_),
    .A1(net735),
    .B1(_0777_),
    .X(_0778_));
 sg13g2_o21ai_1 _3600_ (.B1(_0778_),
    .Y(_0779_),
    .A1(net778),
    .A2(_0773_));
 sg13g2_and2_1 _3601_ (.A(net847),
    .B(_0779_),
    .X(_0105_));
 sg13g2_and2_1 _3602_ (.A(net834),
    .B(net675),
    .X(_0780_));
 sg13g2_a22oi_1 _3603_ (.Y(_0781_),
    .B1(_0780_),
    .B2(net669),
    .A2(_0742_),
    .A1(net326));
 sg13g2_or2_1 _3604_ (.X(_0782_),
    .B(_0781_),
    .A(net778));
 sg13g2_nand2_1 _3605_ (.Y(_0783_),
    .A(_1690_),
    .B(_0775_));
 sg13g2_xnor2_1 _3606_ (.Y(_0784_),
    .A(_1689_),
    .B(_0783_));
 sg13g2_a21oi_1 _3607_ (.A1(_1404_),
    .A2(net683),
    .Y(_0785_),
    .B1(net689));
 sg13g2_o21ai_1 _3608_ (.B1(_0785_),
    .Y(_0786_),
    .A1(net683),
    .A2(_0784_));
 sg13g2_a21oi_1 _3609_ (.A1(_0782_),
    .A2(_0786_),
    .Y(_0106_),
    .B1(net813));
 sg13g2_and2_1 _3610_ (.A(net832),
    .B(net675),
    .X(_0787_));
 sg13g2_a22oi_1 _3611_ (.Y(_0788_),
    .B1(_0787_),
    .B2(net667),
    .A2(_0742_),
    .A1(\collatz.iter[30] ));
 sg13g2_or2_1 _3612_ (.X(_0789_),
    .B(_0788_),
    .A(net779));
 sg13g2_a21oi_1 _3613_ (.A1(_1703_),
    .A2(_0775_),
    .Y(_0790_),
    .B1(_1456_));
 sg13g2_nor2b_1 _3614_ (.A(_1687_),
    .B_N(_0790_),
    .Y(_0791_));
 sg13g2_xor2_1 _3615_ (.B(_0790_),
    .A(_1687_),
    .X(_0792_));
 sg13g2_o21ai_1 _3616_ (.B1(net779),
    .Y(_0793_),
    .A1(\collatz.iter[31] ),
    .A2(net735));
 sg13g2_a21o_1 _3617_ (.A2(_0792_),
    .A1(net735),
    .B1(_0793_),
    .X(_0794_));
 sg13g2_a21oi_1 _3618_ (.A1(_0789_),
    .A2(_0794_),
    .Y(_0107_),
    .B1(net814));
 sg13g2_and2_1 _3619_ (.A(net830),
    .B(net675),
    .X(_0795_));
 sg13g2_a22oi_1 _3620_ (.Y(_0796_),
    .B1(_0795_),
    .B2(net667),
    .A2(_0742_),
    .A1(\collatz.iter[31] ));
 sg13g2_or2_1 _3621_ (.X(_0797_),
    .B(_0796_),
    .A(net779));
 sg13g2_a21oi_1 _3622_ (.A1(\collatz.iter[30] ),
    .A2(\collatz.iter[29] ),
    .Y(_0798_),
    .B1(_0791_));
 sg13g2_xnor2_1 _3623_ (.Y(_0799_),
    .A(_1688_),
    .B(_0798_));
 sg13g2_a21oi_1 _3624_ (.A1(net735),
    .A2(_0799_),
    .Y(_0800_),
    .B1(net688));
 sg13g2_o21ai_1 _3625_ (.B1(_0800_),
    .Y(_0801_),
    .A1(\collatz.iter[32] ),
    .A2(net737));
 sg13g2_a21oi_1 _3626_ (.A1(_0797_),
    .A2(_0801_),
    .Y(_0108_),
    .B1(net814));
 sg13g2_nor2b_1 _3627_ (.A(_1778_),
    .B_N(_1843_),
    .Y(_0802_));
 sg13g2_a21o_1 _3628_ (.A2(_1777_),
    .A1(_1776_),
    .B1(_1843_),
    .X(_0803_));
 sg13g2_nor2_1 _3629_ (.A(net680),
    .B(_0802_),
    .Y(_0804_));
 sg13g2_a22oi_1 _3630_ (.Y(_0805_),
    .B1(_0803_),
    .B2(_0804_),
    .A2(net680),
    .A1(net709));
 sg13g2_nor2b_1 _3631_ (.A(net1),
    .B_N(net826),
    .Y(_0806_));
 sg13g2_and2_1 _3632_ (.A(_1419_),
    .B(_0806_),
    .X(_0807_));
 sg13g2_nand2_1 _3633_ (.Y(_0808_),
    .A(net667),
    .B(_0807_));
 sg13g2_mux2_1 _3634_ (.A0(net844),
    .A1(\collatz.iter[32] ),
    .S(_0808_),
    .X(_0809_));
 sg13g2_o21ai_1 _3635_ (.B1(net846),
    .Y(_0810_),
    .A1(net773),
    .A2(_0809_));
 sg13g2_a21oi_1 _3636_ (.A1(net773),
    .A2(_0805_),
    .Y(_0109_),
    .B1(_0810_));
 sg13g2_nor2b_2 _3637_ (.A(net650),
    .B_N(_0808_),
    .Y(_0811_));
 sg13g2_and2_1 _3638_ (.A(net842),
    .B(net674),
    .X(_0812_));
 sg13g2_a22oi_1 _3639_ (.Y(_0813_),
    .B1(_0812_),
    .B2(net666),
    .A2(_0811_),
    .A1(net709));
 sg13g2_nand2_1 _3640_ (.Y(_0814_),
    .A(_1842_),
    .B(_0803_));
 sg13g2_xor2_1 _3641_ (.B(_0814_),
    .A(_1844_),
    .X(_0815_));
 sg13g2_a21oi_1 _3642_ (.A1(net726),
    .A2(_0815_),
    .Y(_0816_),
    .B1(net686));
 sg13g2_o21ai_1 _3643_ (.B1(_0816_),
    .Y(_0817_),
    .A1(\collatz.iter[34] ),
    .A2(net726));
 sg13g2_o21ai_1 _3644_ (.B1(_0817_),
    .Y(_0818_),
    .A1(net773),
    .A2(_0813_));
 sg13g2_and2_1 _3645_ (.A(net846),
    .B(_0818_),
    .X(_0110_));
 sg13g2_and2_1 _3646_ (.A(net840),
    .B(net674),
    .X(_0819_));
 sg13g2_a22oi_1 _3647_ (.Y(_0820_),
    .B1(_0819_),
    .B2(net666),
    .A2(_0811_),
    .A1(\collatz.iter[34] ));
 sg13g2_a21oi_1 _3648_ (.A1(_1850_),
    .A2(_0803_),
    .Y(_0821_),
    .B1(_1432_));
 sg13g2_xnor2_1 _3649_ (.Y(_0822_),
    .A(_1839_),
    .B(_0821_));
 sg13g2_o21ai_1 _3650_ (.B1(net773),
    .Y(_0823_),
    .A1(\collatz.iter[35] ),
    .A2(net725));
 sg13g2_a21o_1 _3651_ (.A2(_0822_),
    .A1(net725),
    .B1(_0823_),
    .X(_0824_));
 sg13g2_o21ai_1 _3652_ (.B1(_0824_),
    .Y(_0825_),
    .A1(net773),
    .A2(_0820_));
 sg13g2_and2_1 _3653_ (.A(net846),
    .B(_0825_),
    .X(_0111_));
 sg13g2_and2_1 _3654_ (.A(net838),
    .B(net674),
    .X(_0826_));
 sg13g2_a22oi_1 _3655_ (.Y(_0827_),
    .B1(_0826_),
    .B2(net666),
    .A2(_0811_),
    .A1(\collatz.iter[35] ));
 sg13g2_or2_1 _3656_ (.X(_0828_),
    .B(_0827_),
    .A(net772));
 sg13g2_a21oi_1 _3657_ (.A1(_1839_),
    .A2(_0821_),
    .Y(_0829_),
    .B1(_1838_));
 sg13g2_xor2_1 _3658_ (.B(_0829_),
    .A(_1840_),
    .X(_0830_));
 sg13g2_a21oi_1 _3659_ (.A1(net721),
    .A2(_0830_),
    .Y(_0831_),
    .B1(net686));
 sg13g2_o21ai_1 _3660_ (.B1(_0831_),
    .Y(_0832_),
    .A1(\collatz.iter[36] ),
    .A2(net728));
 sg13g2_a21oi_1 _3661_ (.A1(_0828_),
    .A2(_0832_),
    .Y(_0112_),
    .B1(net810));
 sg13g2_and2_1 _3662_ (.A(net836),
    .B(net674),
    .X(_0833_));
 sg13g2_a22oi_1 _3663_ (.Y(_0834_),
    .B1(_0833_),
    .B2(net666),
    .A2(_0811_),
    .A1(\collatz.iter[36] ));
 sg13g2_a21oi_2 _3664_ (.B1(_1853_),
    .Y(_0835_),
    .A2(_1845_),
    .A1(_1778_));
 sg13g2_nand2b_1 _3665_ (.Y(_0836_),
    .B(_1835_),
    .A_N(_0835_));
 sg13g2_xor2_1 _3666_ (.B(_0835_),
    .A(_1835_),
    .X(_0837_));
 sg13g2_o21ai_1 _3667_ (.B1(net772),
    .Y(_0838_),
    .A1(net708),
    .A2(net722));
 sg13g2_a21o_1 _3668_ (.A2(_0837_),
    .A1(net722),
    .B1(_0838_),
    .X(_0839_));
 sg13g2_o21ai_1 _3669_ (.B1(_0839_),
    .Y(_0840_),
    .A1(net770),
    .A2(_0834_));
 sg13g2_and2_1 _3670_ (.A(net846),
    .B(_0840_),
    .X(_0113_));
 sg13g2_and2_1 _3671_ (.A(net834),
    .B(net674),
    .X(_0841_));
 sg13g2_a22oi_1 _3672_ (.Y(_0842_),
    .B1(_0841_),
    .B2(net666),
    .A2(_0811_),
    .A1(net708));
 sg13g2_or2_1 _3673_ (.X(_0843_),
    .B(_0842_),
    .A(net770));
 sg13g2_nand2_1 _3674_ (.Y(_0844_),
    .A(_1834_),
    .B(_0836_));
 sg13g2_xnor2_1 _3675_ (.Y(_0845_),
    .A(_1836_),
    .B(_0844_));
 sg13g2_a21oi_1 _3676_ (.A1(net722),
    .A2(_0845_),
    .Y(_0846_),
    .B1(net686));
 sg13g2_o21ai_1 _3677_ (.B1(_0846_),
    .Y(_0847_),
    .A1(net288),
    .A2(net722));
 sg13g2_a21oi_1 _3678_ (.A1(_0843_),
    .A2(_0847_),
    .Y(_0114_),
    .B1(net809));
 sg13g2_and2_1 _3679_ (.A(net832),
    .B(net674),
    .X(_0848_));
 sg13g2_a22oi_1 _3680_ (.Y(_0849_),
    .B1(_0848_),
    .B2(net666),
    .A2(_0811_),
    .A1(net341));
 sg13g2_or2_1 _3681_ (.X(_0850_),
    .B(_0849_),
    .A(net770));
 sg13g2_a21oi_1 _3682_ (.A1(_1856_),
    .A2(_0836_),
    .Y(_0851_),
    .B1(_1449_));
 sg13g2_xnor2_1 _3683_ (.Y(_0852_),
    .A(_1831_),
    .B(_0851_));
 sg13g2_o21ai_1 _3684_ (.B1(net772),
    .Y(_0853_),
    .A1(\collatz.iter[39] ),
    .A2(net722));
 sg13g2_a21o_1 _3685_ (.A2(_0852_),
    .A1(net722),
    .B1(_0853_),
    .X(_0854_));
 sg13g2_a21oi_1 _3686_ (.A1(_0850_),
    .A2(_0854_),
    .Y(_0115_),
    .B1(net809));
 sg13g2_and2_1 _3687_ (.A(net830),
    .B(net674),
    .X(_0855_));
 sg13g2_a22oi_1 _3688_ (.Y(_0856_),
    .B1(_0855_),
    .B2(net666),
    .A2(_0811_),
    .A1(\collatz.iter[39] ));
 sg13g2_or2_1 _3689_ (.X(_0857_),
    .B(_0856_),
    .A(net772));
 sg13g2_a21oi_1 _3690_ (.A1(_1831_),
    .A2(_0851_),
    .Y(_0858_),
    .B1(_1830_));
 sg13g2_xor2_1 _3691_ (.B(_0858_),
    .A(_1832_),
    .X(_0859_));
 sg13g2_a21oi_1 _3692_ (.A1(net721),
    .A2(_0859_),
    .Y(_0860_),
    .B1(net686));
 sg13g2_o21ai_1 _3693_ (.B1(_0860_),
    .Y(_0861_),
    .A1(net328),
    .A2(net721));
 sg13g2_a21oi_1 _3694_ (.A1(_0857_),
    .A2(_0861_),
    .Y(_0116_),
    .B1(net809));
 sg13g2_and3_1 _3695_ (.X(_0862_),
    .A(net829),
    .B(net667),
    .C(_0806_));
 sg13g2_nor2_2 _3696_ (.A(net650),
    .B(net661),
    .Y(_0863_));
 sg13g2_a22oi_1 _3697_ (.Y(_0864_),
    .B1(_0863_),
    .B2(\collatz.iter[40] ),
    .A2(net661),
    .A1(net844));
 sg13g2_and2_1 _3698_ (.A(_1778_),
    .B(_1846_),
    .X(_0865_));
 sg13g2_nor3_2 _3699_ (.A(_1854_),
    .B(_1857_),
    .C(_0865_),
    .Y(_0866_));
 sg13g2_nand2b_1 _3700_ (.Y(_0867_),
    .B(_1826_),
    .A_N(_0866_));
 sg13g2_xor2_1 _3701_ (.B(_0866_),
    .A(_1826_),
    .X(_0868_));
 sg13g2_o21ai_1 _3702_ (.B1(net775),
    .Y(_0869_),
    .A1(net707),
    .A2(net721));
 sg13g2_a21o_1 _3703_ (.A2(_0868_),
    .A1(net721),
    .B1(_0869_),
    .X(_0870_));
 sg13g2_o21ai_1 _3704_ (.B1(_0870_),
    .Y(_0871_),
    .A1(net775),
    .A2(_0864_));
 sg13g2_and2_1 _3705_ (.A(net846),
    .B(_0871_),
    .X(_0117_));
 sg13g2_a22oi_1 _3706_ (.Y(_0872_),
    .B1(_0863_),
    .B2(net707),
    .A2(net661),
    .A1(net842));
 sg13g2_or2_1 _3707_ (.X(_0873_),
    .B(_0872_),
    .A(net772));
 sg13g2_nand2_1 _3708_ (.Y(_0874_),
    .A(_1825_),
    .B(_0867_));
 sg13g2_xnor2_1 _3709_ (.Y(_0875_),
    .A(_1827_),
    .B(_0874_));
 sg13g2_a21oi_1 _3710_ (.A1(net721),
    .A2(_0875_),
    .Y(_0876_),
    .B1(net686));
 sg13g2_o21ai_1 _3711_ (.B1(_0876_),
    .Y(_0877_),
    .A1(net322),
    .A2(net721));
 sg13g2_a21oi_1 _3712_ (.A1(_0873_),
    .A2(_0877_),
    .Y(_0118_),
    .B1(net809));
 sg13g2_a22oi_1 _3713_ (.Y(_0878_),
    .B1(_0863_),
    .B2(\collatz.iter[42] ),
    .A2(net661),
    .A1(net840));
 sg13g2_or2_1 _3714_ (.X(_0879_),
    .B(_0878_),
    .A(net772));
 sg13g2_a21oi_1 _3715_ (.A1(_1862_),
    .A2(_0867_),
    .Y(_0880_),
    .B1(_1443_));
 sg13g2_xnor2_1 _3716_ (.Y(_0881_),
    .A(_1823_),
    .B(_0880_));
 sg13g2_o21ai_1 _3717_ (.B1(net772),
    .Y(_0882_),
    .A1(\collatz.iter[43] ),
    .A2(net725));
 sg13g2_a21o_1 _3718_ (.A2(_0881_),
    .A1(net725),
    .B1(_0882_),
    .X(_0883_));
 sg13g2_a21oi_1 _3719_ (.A1(_0879_),
    .A2(_0883_),
    .Y(_0119_),
    .B1(net809));
 sg13g2_a22oi_1 _3720_ (.Y(_0884_),
    .B1(_0863_),
    .B2(\collatz.iter[43] ),
    .A2(net661),
    .A1(net838));
 sg13g2_or2_1 _3721_ (.X(_0885_),
    .B(_0884_),
    .A(net774));
 sg13g2_a21oi_1 _3722_ (.A1(_1823_),
    .A2(_0880_),
    .Y(_0886_),
    .B1(_1822_));
 sg13g2_xor2_1 _3723_ (.B(_0886_),
    .A(_1824_),
    .X(_0887_));
 sg13g2_a21oi_1 _3724_ (.A1(net725),
    .A2(_0887_),
    .Y(_0888_),
    .B1(net686));
 sg13g2_o21ai_1 _3725_ (.B1(_0888_),
    .Y(_0889_),
    .A1(net318),
    .A2(net725));
 sg13g2_a21oi_1 _3726_ (.A1(_0885_),
    .A2(_0889_),
    .Y(_0120_),
    .B1(net810));
 sg13g2_a22oi_1 _3727_ (.Y(_0890_),
    .B1(_0863_),
    .B2(net332),
    .A2(_0862_),
    .A1(net836));
 sg13g2_or2_1 _3728_ (.X(_0891_),
    .B(_0890_),
    .A(net773));
 sg13g2_o21ai_1 _3729_ (.B1(_1865_),
    .Y(_0892_),
    .A1(_1828_),
    .A2(_0866_));
 sg13g2_nand2_1 _3730_ (.Y(_0893_),
    .A(_1820_),
    .B(_0892_));
 sg13g2_xnor2_1 _3731_ (.Y(_0894_),
    .A(_1820_),
    .B(_0892_));
 sg13g2_o21ai_1 _3732_ (.B1(net774),
    .Y(_0895_),
    .A1(net706),
    .A2(net726));
 sg13g2_a21o_1 _3733_ (.A2(_0894_),
    .A1(net725),
    .B1(_0895_),
    .X(_0896_));
 sg13g2_a21oi_1 _3734_ (.A1(_0891_),
    .A2(_0896_),
    .Y(_0121_),
    .B1(net810));
 sg13g2_a22oi_1 _3735_ (.Y(_0897_),
    .B1(_0863_),
    .B2(net706),
    .A2(net661),
    .A1(net834));
 sg13g2_or2_1 _3736_ (.X(_0898_),
    .B(_0897_),
    .A(net773));
 sg13g2_nand2_1 _3737_ (.Y(_0899_),
    .A(_1819_),
    .B(_0893_));
 sg13g2_xnor2_1 _3738_ (.Y(_0900_),
    .A(_1818_),
    .B(_0899_));
 sg13g2_a21oi_1 _3739_ (.A1(net725),
    .A2(_0900_),
    .Y(_0901_),
    .B1(net686));
 sg13g2_o21ai_1 _3740_ (.B1(_0901_),
    .Y(_0902_),
    .A1(net321),
    .A2(net737));
 sg13g2_a21oi_1 _3741_ (.A1(_0898_),
    .A2(_0902_),
    .Y(_0122_),
    .B1(net814));
 sg13g2_a22oi_1 _3742_ (.Y(_0903_),
    .B1(_0863_),
    .B2(net321),
    .A2(net661),
    .A1(net832));
 sg13g2_or2_1 _3743_ (.X(_0904_),
    .B(_0903_),
    .A(net774));
 sg13g2_a21oi_1 _3744_ (.A1(_1859_),
    .A2(_0893_),
    .Y(_0905_),
    .B1(_1439_));
 sg13g2_xnor2_1 _3745_ (.Y(_0906_),
    .A(_1815_),
    .B(_0905_));
 sg13g2_o21ai_1 _3746_ (.B1(net774),
    .Y(_0907_),
    .A1(\collatz.iter[47] ),
    .A2(net737));
 sg13g2_a21o_1 _3747_ (.A2(_0906_),
    .A1(net726),
    .B1(_0907_),
    .X(_0908_));
 sg13g2_a21oi_1 _3748_ (.A1(_0904_),
    .A2(_0908_),
    .Y(_0123_),
    .B1(net814));
 sg13g2_a22oi_1 _3749_ (.Y(_0909_),
    .B1(_0863_),
    .B2(\collatz.iter[47] ),
    .A2(net661),
    .A1(net830));
 sg13g2_or2_1 _3750_ (.X(_0910_),
    .B(_0909_),
    .A(net772));
 sg13g2_a21oi_1 _3751_ (.A1(_1815_),
    .A2(_0905_),
    .Y(_0911_),
    .B1(_1814_));
 sg13g2_xor2_1 _3752_ (.B(_0911_),
    .A(_1816_),
    .X(_0912_));
 sg13g2_a21oi_1 _3753_ (.A1(net721),
    .A2(_0912_),
    .Y(_0913_),
    .B1(net686));
 sg13g2_o21ai_1 _3754_ (.B1(_0913_),
    .Y(_0914_),
    .A1(net320),
    .A2(net722));
 sg13g2_a21oi_1 _3755_ (.A1(_0910_),
    .A2(_0914_),
    .Y(_0124_),
    .B1(net809));
 sg13g2_a21oi_2 _3756_ (.B1(net650),
    .Y(_0915_),
    .A2(net665),
    .A1(_1509_));
 sg13g2_and2_1 _3757_ (.A(net844),
    .B(net679),
    .X(_0916_));
 sg13g2_a22oi_1 _3758_ (.Y(_0917_),
    .B1(_0916_),
    .B2(net664),
    .A2(_0915_),
    .A1(\collatz.iter[48] ));
 sg13g2_a21oi_2 _3759_ (.B1(_1868_),
    .Y(_0918_),
    .A2(_1847_),
    .A1(_1778_));
 sg13g2_nand2b_1 _3760_ (.Y(_0919_),
    .B(_1809_),
    .A_N(_0918_));
 sg13g2_xor2_1 _3761_ (.B(_0918_),
    .A(_1809_),
    .X(_0920_));
 sg13g2_o21ai_1 _3762_ (.B1(net770),
    .Y(_0921_),
    .A1(\collatz.iter[49] ),
    .A2(net714));
 sg13g2_a21o_1 _3763_ (.A2(_0920_),
    .A1(net714),
    .B1(_0921_),
    .X(_0922_));
 sg13g2_o21ai_1 _3764_ (.B1(_0922_),
    .Y(_0923_),
    .A1(net770),
    .A2(_0917_));
 sg13g2_and2_1 _3765_ (.A(net846),
    .B(_0923_),
    .X(_0125_));
 sg13g2_and2_1 _3766_ (.A(net842),
    .B(_1509_),
    .X(_0924_));
 sg13g2_a22oi_1 _3767_ (.Y(_0925_),
    .B1(_0924_),
    .B2(net664),
    .A2(_0915_),
    .A1(\collatz.iter[49] ));
 sg13g2_or2_1 _3768_ (.X(_0926_),
    .B(_0925_),
    .A(net763));
 sg13g2_nand2_1 _3769_ (.Y(_0927_),
    .A(_1808_),
    .B(_0919_));
 sg13g2_xnor2_1 _3770_ (.Y(_0928_),
    .A(_1810_),
    .B(_0927_));
 sg13g2_a21oi_1 _3771_ (.A1(net715),
    .A2(_0928_),
    .Y(_0929_),
    .B1(net684));
 sg13g2_o21ai_1 _3772_ (.B1(_0929_),
    .Y(_0930_),
    .A1(\collatz.iter[50] ),
    .A2(net715));
 sg13g2_a21oi_1 _3773_ (.A1(_0926_),
    .A2(_0930_),
    .Y(_0126_),
    .B1(net806));
 sg13g2_and2_1 _3774_ (.A(net840),
    .B(net679),
    .X(_0931_));
 sg13g2_a22oi_1 _3775_ (.Y(_0932_),
    .B1(_0931_),
    .B2(net664),
    .A2(_0915_),
    .A1(\collatz.iter[50] ));
 sg13g2_or2_1 _3776_ (.X(_0933_),
    .B(_0932_),
    .A(net763));
 sg13g2_a21oi_1 _3777_ (.A1(_1870_),
    .A2(_0919_),
    .Y(_0934_),
    .B1(_1436_));
 sg13g2_xnor2_1 _3778_ (.Y(_0935_),
    .A(_1806_),
    .B(_0934_));
 sg13g2_o21ai_1 _3779_ (.B1(net770),
    .Y(_0936_),
    .A1(net705),
    .A2(net715));
 sg13g2_a21o_1 _3780_ (.A2(_0935_),
    .A1(net715),
    .B1(_0936_),
    .X(_0937_));
 sg13g2_a21oi_1 _3781_ (.A1(_0933_),
    .A2(_0937_),
    .Y(_0127_),
    .B1(net806));
 sg13g2_and2_1 _3782_ (.A(net838),
    .B(net679),
    .X(_0938_));
 sg13g2_a22oi_1 _3783_ (.Y(_0939_),
    .B1(_0938_),
    .B2(net664),
    .A2(_0915_),
    .A1(net705));
 sg13g2_or2_1 _3784_ (.X(_0940_),
    .B(_0939_),
    .A(net763));
 sg13g2_a21oi_1 _3785_ (.A1(_1806_),
    .A2(_0934_),
    .Y(_0941_),
    .B1(_1805_));
 sg13g2_xor2_1 _3786_ (.B(_0941_),
    .A(_1807_),
    .X(_0942_));
 sg13g2_a21oi_1 _3787_ (.A1(net715),
    .A2(_0942_),
    .Y(_0943_),
    .B1(net684));
 sg13g2_o21ai_1 _3788_ (.B1(_0943_),
    .Y(_0944_),
    .A1(net704),
    .A2(net714));
 sg13g2_a21oi_1 _3789_ (.A1(_0940_),
    .A2(_0944_),
    .Y(_0128_),
    .B1(net806));
 sg13g2_and2_1 _3790_ (.A(net836),
    .B(net679),
    .X(_0945_));
 sg13g2_a22oi_1 _3791_ (.Y(_0946_),
    .B1(_0945_),
    .B2(net664),
    .A2(_0915_),
    .A1(net263));
 sg13g2_or2_1 _3792_ (.X(_0947_),
    .B(_0946_),
    .A(net762));
 sg13g2_or2_1 _3793_ (.X(_0948_),
    .B(_0918_),
    .A(_1811_));
 sg13g2_nand3_1 _3794_ (.B(_1873_),
    .C(_0948_),
    .A(_1803_),
    .Y(_0949_));
 sg13g2_a21o_1 _3795_ (.A2(_0948_),
    .A1(_1873_),
    .B1(_1803_),
    .X(_0950_));
 sg13g2_a21oi_1 _3796_ (.A1(_0949_),
    .A2(_0950_),
    .Y(_0951_),
    .B1(net680));
 sg13g2_o21ai_1 _3797_ (.B1(net763),
    .Y(_0952_),
    .A1(net703),
    .A2(net712));
 sg13g2_or2_1 _3798_ (.X(_0953_),
    .B(_0952_),
    .A(_0951_));
 sg13g2_a21oi_1 _3799_ (.A1(_0947_),
    .A2(_0953_),
    .Y(_0129_),
    .B1(net806));
 sg13g2_and2_1 _3800_ (.A(net834),
    .B(net679),
    .X(_0954_));
 sg13g2_a22oi_1 _3801_ (.Y(_0955_),
    .B1(_0954_),
    .B2(net664),
    .A2(_0915_),
    .A1(net264));
 sg13g2_or2_1 _3802_ (.X(_0956_),
    .B(_0955_),
    .A(net762));
 sg13g2_nand2_1 _3803_ (.Y(_0957_),
    .A(_1801_),
    .B(_0950_));
 sg13g2_xnor2_1 _3804_ (.Y(_0958_),
    .A(_1800_),
    .B(_0957_));
 sg13g2_a21oi_1 _3805_ (.A1(net714),
    .A2(_0958_),
    .Y(_0959_),
    .B1(net684));
 sg13g2_o21ai_1 _3806_ (.B1(_0959_),
    .Y(_0960_),
    .A1(\collatz.iter[54] ),
    .A2(net712));
 sg13g2_a21oi_1 _3807_ (.A1(_0956_),
    .A2(_0960_),
    .Y(_0130_),
    .B1(net806));
 sg13g2_and2_1 _3808_ (.A(net832),
    .B(net679),
    .X(_0961_));
 sg13g2_a22oi_1 _3809_ (.Y(_0962_),
    .B1(_0961_),
    .B2(net664),
    .A2(_0915_),
    .A1(\collatz.iter[54] ));
 sg13g2_or2_1 _3810_ (.X(_0963_),
    .B(_0962_),
    .A(net763));
 sg13g2_a21oi_1 _3811_ (.A1(_1876_),
    .A2(_0950_),
    .Y(_0964_),
    .B1(_1444_));
 sg13g2_xnor2_1 _3812_ (.Y(_0965_),
    .A(_1797_),
    .B(_0964_));
 sg13g2_o21ai_1 _3813_ (.B1(net763),
    .Y(_0966_),
    .A1(\collatz.iter[55] ),
    .A2(net714));
 sg13g2_a21o_1 _3814_ (.A2(_0965_),
    .A1(net714),
    .B1(_0966_),
    .X(_0967_));
 sg13g2_a21oi_1 _3815_ (.A1(_0963_),
    .A2(_0967_),
    .Y(_0131_),
    .B1(net805));
 sg13g2_a22oi_1 _3816_ (.Y(_0968_),
    .B1(_0915_),
    .B2(\collatz.iter[55] ),
    .A2(net664),
    .A1(_1518_));
 sg13g2_or2_1 _3817_ (.X(_0969_),
    .B(_0968_),
    .A(net762));
 sg13g2_a21oi_1 _3818_ (.A1(_1797_),
    .A2(_0964_),
    .Y(_0970_),
    .B1(_1796_));
 sg13g2_xor2_1 _3819_ (.B(_0970_),
    .A(_1798_),
    .X(_0971_));
 sg13g2_a21oi_1 _3820_ (.A1(net714),
    .A2(_0971_),
    .Y(_0972_),
    .B1(net684));
 sg13g2_o21ai_1 _3821_ (.B1(_0972_),
    .Y(_0973_),
    .A1(\collatz.iter[56] ),
    .A2(net714));
 sg13g2_a21oi_1 _3822_ (.A1(_0969_),
    .A2(_0973_),
    .Y(_0132_),
    .B1(net806));
 sg13g2_a21oi_2 _3823_ (.B1(net650),
    .Y(_0974_),
    .A2(net667),
    .A1(net804));
 sg13g2_a22oi_1 _3824_ (.Y(_0975_),
    .B1(_0974_),
    .B2(\collatz.iter[56] ),
    .A2(net665),
    .A1(_1916_));
 sg13g2_o21ai_1 _3825_ (.B1(_1878_),
    .Y(_0976_),
    .A1(_1812_),
    .A2(_0918_));
 sg13g2_nand2_1 _3826_ (.Y(_0977_),
    .A(_1785_),
    .B(_0976_));
 sg13g2_xnor2_1 _3827_ (.Y(_0978_),
    .A(_1785_),
    .B(_0976_));
 sg13g2_o21ai_1 _3828_ (.B1(net763),
    .Y(_0979_),
    .A1(\collatz.iter[57] ),
    .A2(net716));
 sg13g2_a21o_1 _3829_ (.A2(_0978_),
    .A1(net716),
    .B1(_0979_),
    .X(_0980_));
 sg13g2_o21ai_1 _3830_ (.B1(_0980_),
    .Y(_0981_),
    .A1(net762),
    .A2(_0975_));
 sg13g2_and2_1 _3831_ (.A(net846),
    .B(_0981_),
    .X(_0133_));
 sg13g2_a22oi_1 _3832_ (.Y(_0982_),
    .B1(_0974_),
    .B2(net327),
    .A2(net665),
    .A1(_1939_));
 sg13g2_or2_1 _3833_ (.X(_0983_),
    .B(_0982_),
    .A(net765));
 sg13g2_nand2_1 _3834_ (.Y(_0984_),
    .A(_1784_),
    .B(_0977_));
 sg13g2_xnor2_1 _3835_ (.Y(_0985_),
    .A(_1783_),
    .B(_0984_));
 sg13g2_a21oi_1 _3836_ (.A1(net716),
    .A2(_0985_),
    .Y(_0986_),
    .B1(net684));
 sg13g2_o21ai_1 _3837_ (.B1(_0986_),
    .Y(_0987_),
    .A1(net316),
    .A2(net718));
 sg13g2_a21oi_1 _3838_ (.A1(_0983_),
    .A2(_0987_),
    .Y(_0134_),
    .B1(net808));
 sg13g2_a22oi_1 _3839_ (.Y(_0988_),
    .B1(_0974_),
    .B2(net316),
    .A2(net665),
    .A1(_1947_));
 sg13g2_or2_1 _3840_ (.X(_0989_),
    .B(_0988_),
    .A(net764));
 sg13g2_a21oi_1 _3841_ (.A1(_1881_),
    .A2(_0977_),
    .Y(_0990_),
    .B1(_1457_));
 sg13g2_xnor2_1 _3842_ (.Y(_0991_),
    .A(_1780_),
    .B(_0990_));
 sg13g2_o21ai_1 _3843_ (.B1(net765),
    .Y(_0992_),
    .A1(\collatz.iter[59] ),
    .A2(net718));
 sg13g2_a21o_1 _3844_ (.A2(_0991_),
    .A1(net718),
    .B1(_0992_),
    .X(_0993_));
 sg13g2_a21oi_1 _3845_ (.A1(_0989_),
    .A2(_0993_),
    .Y(_0135_),
    .B1(net808));
 sg13g2_a22oi_1 _3846_ (.Y(_0994_),
    .B1(_0974_),
    .B2(\collatz.iter[59] ),
    .A2(net665),
    .A1(_1957_));
 sg13g2_or2_1 _3847_ (.X(_0995_),
    .B(_0994_),
    .A(net765));
 sg13g2_a21oi_1 _3848_ (.A1(_1780_),
    .A2(_0990_),
    .Y(_0996_),
    .B1(_1779_));
 sg13g2_xor2_1 _3849_ (.B(_0996_),
    .A(_1781_),
    .X(_0997_));
 sg13g2_a21oi_1 _3850_ (.A1(net718),
    .A2(_0997_),
    .Y(_0998_),
    .B1(net684));
 sg13g2_o21ai_1 _3851_ (.B1(_0998_),
    .Y(_0999_),
    .A1(net315),
    .A2(net718));
 sg13g2_a21oi_1 _3852_ (.A1(_0995_),
    .A2(_0999_),
    .Y(_0136_),
    .B1(net807));
 sg13g2_a22oi_1 _3853_ (.Y(_1000_),
    .B1(_0974_),
    .B2(net339),
    .A2(net665),
    .A1(_1965_));
 sg13g2_or2_1 _3854_ (.X(_1001_),
    .B(_1000_),
    .A(net764));
 sg13g2_a21oi_1 _3855_ (.A1(_1786_),
    .A2(_0976_),
    .Y(_1002_),
    .B1(_1883_));
 sg13g2_or2_1 _3856_ (.X(_1003_),
    .B(_1002_),
    .A(_1788_));
 sg13g2_xnor2_1 _3857_ (.Y(_1004_),
    .A(_1788_),
    .B(_1002_));
 sg13g2_o21ai_1 _3858_ (.B1(net764),
    .Y(_1005_),
    .A1(net702),
    .A2(net718));
 sg13g2_a21o_1 _3859_ (.A2(_1004_),
    .A1(net719),
    .B1(_1005_),
    .X(_1006_));
 sg13g2_a21oi_1 _3860_ (.A1(_1001_),
    .A2(_1006_),
    .Y(_0137_),
    .B1(net807));
 sg13g2_a22oi_1 _3861_ (.Y(_1007_),
    .B1(_0974_),
    .B2(net702),
    .A2(net667),
    .A1(_0206_));
 sg13g2_or2_1 _3862_ (.X(_1008_),
    .B(_1007_),
    .A(net764));
 sg13g2_nand2_1 _3863_ (.Y(_1009_),
    .A(_1787_),
    .B(_1003_));
 sg13g2_xor2_1 _3864_ (.B(_1009_),
    .A(_1789_),
    .X(_1010_));
 sg13g2_a21oi_1 _3865_ (.A1(net718),
    .A2(_1010_),
    .Y(_1011_),
    .B1(net685));
 sg13g2_o21ai_1 _3866_ (.B1(_1011_),
    .Y(_1012_),
    .A1(net289),
    .A2(net718));
 sg13g2_a21oi_1 _3867_ (.A1(_1008_),
    .A2(_1012_),
    .Y(_0138_),
    .B1(net807));
 sg13g2_a22oi_1 _3868_ (.Y(_1013_),
    .B1(_0974_),
    .B2(net289),
    .A2(net670),
    .A1(_0214_));
 sg13g2_or2_1 _3869_ (.X(_1014_),
    .B(_1013_),
    .A(net764));
 sg13g2_a21oi_1 _3870_ (.A1(_1880_),
    .A2(_1003_),
    .Y(_1015_),
    .B1(_1427_));
 sg13g2_xnor2_1 _3871_ (.Y(_1016_),
    .A(_1792_),
    .B(_1015_));
 sg13g2_o21ai_1 _3872_ (.B1(net764),
    .Y(_1017_),
    .A1(\collatz.iter[63] ),
    .A2(net730));
 sg13g2_a21o_1 _3873_ (.A2(_1016_),
    .A1(net730),
    .B1(_1017_),
    .X(_1018_));
 sg13g2_a21oi_1 _3874_ (.A1(_1014_),
    .A2(_1018_),
    .Y(_0139_),
    .B1(net812));
 sg13g2_a22oi_1 _3875_ (.Y(_1019_),
    .B1(_0974_),
    .B2(\collatz.iter[63] ),
    .A2(net667),
    .A1(_0224_));
 sg13g2_or2_1 _3876_ (.X(_1020_),
    .B(_1019_),
    .A(net767));
 sg13g2_a21oi_1 _3877_ (.A1(_1792_),
    .A2(_1015_),
    .Y(_1021_),
    .B1(_1791_));
 sg13g2_xor2_1 _3878_ (.B(_1021_),
    .A(_1793_),
    .X(_1022_));
 sg13g2_a21oi_1 _3879_ (.A1(net730),
    .A2(_1022_),
    .Y(_1023_),
    .B1(net688));
 sg13g2_o21ai_1 _3880_ (.B1(_1023_),
    .Y(_1024_),
    .A1(net267),
    .A2(net729));
 sg13g2_a21oi_1 _3881_ (.A1(_1020_),
    .A2(_1024_),
    .Y(_0140_),
    .B1(net811));
 sg13g2_and3_1 _3882_ (.X(_1025_),
    .A(net3),
    .B(_1511_),
    .C(_0564_));
 sg13g2_nor2_2 _3883_ (.A(net650),
    .B(net663),
    .Y(_1026_));
 sg13g2_a22oi_1 _3884_ (.Y(_1027_),
    .B1(_1026_),
    .B2(net267),
    .A2(net663),
    .A1(net844));
 sg13g2_o21ai_1 _3885_ (.B1(_1889_),
    .Y(_1028_),
    .A1(_1849_),
    .A2(_1887_));
 sg13g2_xor2_1 _3886_ (.B(_1889_),
    .A(_1888_),
    .X(_1029_));
 sg13g2_o21ai_1 _3887_ (.B1(net767),
    .Y(_1030_),
    .A1(\collatz.iter[65] ),
    .A2(net733));
 sg13g2_a21o_1 _3888_ (.A2(_1029_),
    .A1(net733),
    .B1(_1030_),
    .X(_1031_));
 sg13g2_o21ai_1 _3889_ (.B1(_1031_),
    .Y(_1032_),
    .A1(net766),
    .A2(_1027_));
 sg13g2_and2_1 _3890_ (.A(net847),
    .B(_1032_),
    .X(_0141_));
 sg13g2_a22oi_1 _3891_ (.Y(_1033_),
    .B1(_1026_),
    .B2(\collatz.iter[65] ),
    .A2(net663),
    .A1(net842));
 sg13g2_or2_1 _3892_ (.X(_1034_),
    .B(_1033_),
    .A(net766));
 sg13g2_nand2_1 _3893_ (.Y(_1035_),
    .A(_1664_),
    .B(_1028_));
 sg13g2_xnor2_1 _3894_ (.Y(_1036_),
    .A(_1890_),
    .B(_1035_));
 sg13g2_a21oi_1 _3895_ (.A1(net732),
    .A2(_1036_),
    .Y(_1037_),
    .B1(net688));
 sg13g2_o21ai_1 _3896_ (.B1(_1037_),
    .Y(_1038_),
    .A1(net278),
    .A2(net732));
 sg13g2_a21oi_1 _3897_ (.A1(_1034_),
    .A2(_1038_),
    .Y(_0142_),
    .B1(net812));
 sg13g2_a22oi_1 _3898_ (.Y(_1039_),
    .B1(_1026_),
    .B2(net278),
    .A2(net663),
    .A1(net840));
 sg13g2_or2_1 _3899_ (.X(_1040_),
    .B(_1039_),
    .A(net766));
 sg13g2_a21oi_1 _3900_ (.A1(_1665_),
    .A2(_1028_),
    .Y(_1041_),
    .B1(_1430_));
 sg13g2_xnor2_1 _3901_ (.Y(_1042_),
    .A(_1662_),
    .B(_1041_));
 sg13g2_o21ai_1 _3902_ (.B1(net766),
    .Y(_1043_),
    .A1(\collatz.iter[67] ),
    .A2(net732));
 sg13g2_a21o_1 _3903_ (.A2(_1042_),
    .A1(net732),
    .B1(_1043_),
    .X(_1044_));
 sg13g2_a21oi_1 _3904_ (.A1(_1040_),
    .A2(_1044_),
    .Y(_0143_),
    .B1(net812));
 sg13g2_a22oi_1 _3905_ (.Y(_1045_),
    .B1(_1026_),
    .B2(\collatz.iter[67] ),
    .A2(net663),
    .A1(net838));
 sg13g2_or2_1 _3906_ (.X(_1046_),
    .B(_1045_),
    .A(net766));
 sg13g2_a21oi_1 _3907_ (.A1(_1662_),
    .A2(_1041_),
    .Y(_1047_),
    .B1(_1661_));
 sg13g2_xor2_1 _3908_ (.B(_1047_),
    .A(_1663_),
    .X(_1048_));
 sg13g2_a21oi_1 _3909_ (.A1(net732),
    .A2(_1048_),
    .Y(_1049_),
    .B1(net688));
 sg13g2_o21ai_1 _3910_ (.B1(_1049_),
    .Y(_1050_),
    .A1(net280),
    .A2(net732));
 sg13g2_a21oi_1 _3911_ (.A1(_1046_),
    .A2(_1050_),
    .Y(_0144_),
    .B1(net812));
 sg13g2_a22oi_1 _3912_ (.Y(_1051_),
    .B1(_1026_),
    .B2(net280),
    .A2(net663),
    .A1(net836));
 sg13g2_o21ai_1 _3913_ (.B1(_1668_),
    .Y(_1052_),
    .A1(_1888_),
    .A2(_1891_));
 sg13g2_nand2_1 _3914_ (.Y(_1053_),
    .A(_1658_),
    .B(_1052_));
 sg13g2_xnor2_1 _3915_ (.Y(_1054_),
    .A(_1658_),
    .B(_1052_));
 sg13g2_o21ai_1 _3916_ (.B1(net766),
    .Y(_1055_),
    .A1(\collatz.iter[69] ),
    .A2(net732));
 sg13g2_a21o_1 _3917_ (.A2(_1054_),
    .A1(net733),
    .B1(_1055_),
    .X(_1056_));
 sg13g2_o21ai_1 _3918_ (.B1(_1056_),
    .Y(_1057_),
    .A1(net766),
    .A2(_1051_));
 sg13g2_and2_1 _3919_ (.A(net846),
    .B(_1057_),
    .X(_0145_));
 sg13g2_a22oi_1 _3920_ (.Y(_1058_),
    .B1(_1026_),
    .B2(\collatz.iter[69] ),
    .A2(_1025_),
    .A1(net834));
 sg13g2_or2_1 _3921_ (.X(_1059_),
    .B(_1058_),
    .A(net766));
 sg13g2_nand2_1 _3922_ (.Y(_1060_),
    .A(_1657_),
    .B(_1053_));
 sg13g2_xnor2_1 _3923_ (.Y(_1061_),
    .A(_1659_),
    .B(_1060_));
 sg13g2_a21oi_1 _3924_ (.A1(net739),
    .A2(_1061_),
    .Y(_1062_),
    .B1(net691));
 sg13g2_o21ai_1 _3925_ (.B1(_1062_),
    .Y(_1063_),
    .A1(net282),
    .A2(net740));
 sg13g2_a21oi_1 _3926_ (.A1(_1059_),
    .A2(_1063_),
    .Y(_0146_),
    .B1(net816));
 sg13g2_a22oi_1 _3927_ (.Y(_1064_),
    .B1(_1026_),
    .B2(net282),
    .A2(net663),
    .A1(net832));
 sg13g2_or2_1 _3928_ (.X(_1065_),
    .B(_1064_),
    .A(net783));
 sg13g2_a21oi_1 _3929_ (.A1(_1670_),
    .A2(_1053_),
    .Y(_1066_),
    .B1(_1458_));
 sg13g2_xnor2_1 _3930_ (.Y(_1067_),
    .A(_1655_),
    .B(_1066_));
 sg13g2_o21ai_1 _3931_ (.B1(net783),
    .Y(_1068_),
    .A1(\collatz.iter[71] ),
    .A2(net739));
 sg13g2_a21o_1 _3932_ (.A2(_1067_),
    .A1(net739),
    .B1(_1068_),
    .X(_1069_));
 sg13g2_a21oi_1 _3933_ (.A1(_1065_),
    .A2(_1069_),
    .Y(_0147_),
    .B1(net816));
 sg13g2_a22oi_1 _3934_ (.Y(_1070_),
    .B1(_1026_),
    .B2(\collatz.iter[71] ),
    .A2(net663),
    .A1(net831));
 sg13g2_or2_1 _3935_ (.X(_1071_),
    .B(_1070_),
    .A(net783));
 sg13g2_a21oi_1 _3936_ (.A1(_1655_),
    .A2(_1066_),
    .Y(_1072_),
    .B1(_1654_));
 sg13g2_xor2_1 _3937_ (.B(_1072_),
    .A(_1656_),
    .X(_1073_));
 sg13g2_a21oi_1 _3938_ (.A1(net739),
    .A2(_1073_),
    .Y(_1074_),
    .B1(net691));
 sg13g2_o21ai_1 _3939_ (.B1(_1074_),
    .Y(_1075_),
    .A1(net269),
    .A2(net740));
 sg13g2_a21oi_1 _3940_ (.A1(_1071_),
    .A2(_1075_),
    .Y(_0148_),
    .B1(net816));
 sg13g2_and3_1 _3941_ (.X(_1076_),
    .A(net828),
    .B(_1510_),
    .C(net660));
 sg13g2_nor2_2 _3942_ (.A(_1508_),
    .B(net653),
    .Y(_1077_));
 sg13g2_a22oi_1 _3943_ (.Y(_1078_),
    .B1(_1077_),
    .B2(net269),
    .A2(net653),
    .A1(net845));
 sg13g2_o21ai_1 _3944_ (.B1(_1892_),
    .Y(_1079_),
    .A1(_1849_),
    .A2(_1887_));
 sg13g2_nand2b_1 _3945_ (.Y(_1080_),
    .B(_1079_),
    .A_N(_1673_));
 sg13g2_nand2_1 _3946_ (.Y(_1081_),
    .A(_1650_),
    .B(_1080_));
 sg13g2_xnor2_1 _3947_ (.Y(_1082_),
    .A(_1650_),
    .B(_1080_));
 sg13g2_o21ai_1 _3948_ (.B1(net783),
    .Y(_1083_),
    .A1(\collatz.iter[73] ),
    .A2(net739));
 sg13g2_a21o_1 _3949_ (.A2(_1082_),
    .A1(net739),
    .B1(_1083_),
    .X(_1084_));
 sg13g2_o21ai_1 _3950_ (.B1(_1084_),
    .Y(_1085_),
    .A1(net783),
    .A2(_1078_));
 sg13g2_and2_1 _3951_ (.A(net848),
    .B(_1085_),
    .X(_0149_));
 sg13g2_a22oi_1 _3952_ (.Y(_1086_),
    .B1(_1077_),
    .B2(\collatz.iter[73] ),
    .A2(net653),
    .A1(net842));
 sg13g2_or2_1 _3953_ (.X(_1087_),
    .B(_1086_),
    .A(net783));
 sg13g2_nand2_1 _3954_ (.Y(_1088_),
    .A(_1649_),
    .B(_1081_));
 sg13g2_xor2_1 _3955_ (.B(_1088_),
    .A(_1652_),
    .X(_1089_));
 sg13g2_a21oi_1 _3956_ (.A1(net739),
    .A2(_1089_),
    .Y(_1090_),
    .B1(net691));
 sg13g2_o21ai_1 _3957_ (.B1(_1090_),
    .Y(_1091_),
    .A1(net286),
    .A2(net739));
 sg13g2_a21oi_1 _3958_ (.A1(_1087_),
    .A2(_1091_),
    .Y(_0150_),
    .B1(net816));
 sg13g2_a22oi_1 _3959_ (.Y(_1092_),
    .B1(_1077_),
    .B2(net286),
    .A2(net653),
    .A1(net841));
 sg13g2_or2_1 _3960_ (.X(_1093_),
    .B(_1092_),
    .A(net789));
 sg13g2_a21oi_1 _3961_ (.A1(_1677_),
    .A2(_1081_),
    .Y(_1094_),
    .B1(_1431_));
 sg13g2_xnor2_1 _3962_ (.Y(_1095_),
    .A(_1646_),
    .B(_1094_));
 sg13g2_o21ai_1 _3963_ (.B1(net789),
    .Y(_1096_),
    .A1(\collatz.iter[75] ),
    .A2(net742));
 sg13g2_a21o_1 _3964_ (.A2(_1095_),
    .A1(net741),
    .B1(_1096_),
    .X(_1097_));
 sg13g2_a21oi_1 _3965_ (.A1(_1093_),
    .A2(_1097_),
    .Y(_0151_),
    .B1(net817));
 sg13g2_a22oi_1 _3966_ (.Y(_1098_),
    .B1(_1077_),
    .B2(\collatz.iter[75] ),
    .A2(net653),
    .A1(net838));
 sg13g2_or2_1 _3967_ (.X(_1099_),
    .B(_1098_),
    .A(net789));
 sg13g2_a21oi_1 _3968_ (.A1(_1646_),
    .A2(_1094_),
    .Y(_1100_),
    .B1(_1645_));
 sg13g2_xor2_1 _3969_ (.B(_1100_),
    .A(_1647_),
    .X(_1101_));
 sg13g2_a21oi_1 _3970_ (.A1(net742),
    .A2(_1101_),
    .Y(_1102_),
    .B1(net691));
 sg13g2_o21ai_1 _3971_ (.B1(_1102_),
    .Y(_1103_),
    .A1(net295),
    .A2(net742));
 sg13g2_a21oi_1 _3972_ (.A1(_1099_),
    .A2(_1103_),
    .Y(_0152_),
    .B1(net819));
 sg13g2_a22oi_1 _3973_ (.Y(_1104_),
    .B1(_1077_),
    .B2(net295),
    .A2(net653),
    .A1(net836));
 sg13g2_or2_1 _3974_ (.X(_1105_),
    .B(_1104_),
    .A(net789));
 sg13g2_nor3_1 _3975_ (.A(_1648_),
    .B(_1652_),
    .C(_1081_),
    .Y(_1106_));
 sg13g2_nor3_1 _3976_ (.A(_1642_),
    .B(_1679_),
    .C(_1106_),
    .Y(_1107_));
 sg13g2_o21ai_1 _3977_ (.B1(_1642_),
    .Y(_1108_),
    .A1(_1679_),
    .A2(_1106_));
 sg13g2_nand2b_1 _3978_ (.Y(_1109_),
    .B(_1108_),
    .A_N(_1107_));
 sg13g2_o21ai_1 _3979_ (.B1(net789),
    .Y(_1110_),
    .A1(\collatz.iter[77] ),
    .A2(net745));
 sg13g2_a21o_1 _3980_ (.A2(_1109_),
    .A1(net745),
    .B1(_1110_),
    .X(_1111_));
 sg13g2_a21oi_1 _3981_ (.A1(_1105_),
    .A2(_1111_),
    .Y(_0153_),
    .B1(net818));
 sg13g2_a22oi_1 _3982_ (.Y(_1112_),
    .B1(_1077_),
    .B2(\collatz.iter[77] ),
    .A2(net653),
    .A1(net834));
 sg13g2_or2_1 _3983_ (.X(_1113_),
    .B(_1112_),
    .A(net789));
 sg13g2_nand2_1 _3984_ (.Y(_1114_),
    .A(_1641_),
    .B(_1108_));
 sg13g2_xnor2_1 _3985_ (.Y(_1115_),
    .A(_1640_),
    .B(_1114_));
 sg13g2_a21oi_1 _3986_ (.A1(net745),
    .A2(_1115_),
    .Y(_1116_),
    .B1(net690));
 sg13g2_o21ai_1 _3987_ (.B1(_1116_),
    .Y(_1117_),
    .A1(net293),
    .A2(net745));
 sg13g2_a21oi_1 _3988_ (.A1(_1113_),
    .A2(_1117_),
    .Y(_0154_),
    .B1(net818));
 sg13g2_a22oi_1 _3989_ (.Y(_1118_),
    .B1(_1077_),
    .B2(net293),
    .A2(_1076_),
    .A1(net832));
 sg13g2_or2_1 _3990_ (.X(_1119_),
    .B(_1118_),
    .A(net789));
 sg13g2_a21oi_1 _3991_ (.A1(_1674_),
    .A2(_1108_),
    .Y(_1120_),
    .B1(_1433_));
 sg13g2_xnor2_1 _3992_ (.Y(_1121_),
    .A(_1637_),
    .B(_1120_));
 sg13g2_o21ai_1 _3993_ (.B1(net790),
    .Y(_1122_),
    .A1(\collatz.iter[79] ),
    .A2(net745));
 sg13g2_a21o_1 _3994_ (.A2(_1121_),
    .A1(net745),
    .B1(_1122_),
    .X(_1123_));
 sg13g2_a21oi_1 _3995_ (.A1(_1119_),
    .A2(_1123_),
    .Y(_0155_),
    .B1(net818));
 sg13g2_a22oi_1 _3996_ (.Y(_1124_),
    .B1(_1077_),
    .B2(\collatz.iter[79] ),
    .A2(net653),
    .A1(net830));
 sg13g2_or2_1 _3997_ (.X(_1125_),
    .B(_1124_),
    .A(net789));
 sg13g2_a21oi_1 _3998_ (.A1(_1637_),
    .A2(_1120_),
    .Y(_1126_),
    .B1(_1636_));
 sg13g2_xor2_1 _3999_ (.B(_1126_),
    .A(_1638_),
    .X(_1127_));
 sg13g2_a21oi_1 _4000_ (.A1(net745),
    .A2(_1127_),
    .Y(_1128_),
    .B1(net690));
 sg13g2_o21ai_1 _4001_ (.B1(_1128_),
    .Y(_1129_),
    .A1(\collatz.iter[80] ),
    .A2(net745));
 sg13g2_a21oi_1 _4002_ (.A1(_1125_),
    .A2(_1129_),
    .Y(_0156_),
    .B1(net818));
 sg13g2_a21oi_2 _4003_ (.B1(net651),
    .Y(_1130_),
    .A2(_0684_),
    .A1(net659));
 sg13g2_a22oi_1 _4004_ (.Y(_1131_),
    .B1(_1130_),
    .B2(\collatz.iter[80] ),
    .A2(_0686_),
    .A1(net659));
 sg13g2_o21ai_1 _4005_ (.B1(_1680_),
    .Y(_1132_),
    .A1(_1888_),
    .A2(_1893_));
 sg13g2_nand2_1 _4006_ (.Y(_1133_),
    .A(_1681_),
    .B(_1132_));
 sg13g2_xnor2_1 _4007_ (.Y(_1134_),
    .A(_1681_),
    .B(_1132_));
 sg13g2_o21ai_1 _4008_ (.B1(net790),
    .Y(_1135_),
    .A1(net701),
    .A2(net746));
 sg13g2_a21o_1 _4009_ (.A2(_1134_),
    .A1(net746),
    .B1(_1135_),
    .X(_1136_));
 sg13g2_o21ai_1 _4010_ (.B1(_1136_),
    .Y(_1137_),
    .A1(net790),
    .A2(_1131_));
 sg13g2_and2_1 _4011_ (.A(net849),
    .B(_1137_),
    .X(_0157_));
 sg13g2_a22oi_1 _4012_ (.Y(_1138_),
    .B1(_1130_),
    .B2(net701),
    .A2(_0690_),
    .A1(net659));
 sg13g2_or2_1 _4013_ (.X(_1139_),
    .B(_1138_),
    .A(net790));
 sg13g2_nand3_1 _4014_ (.B(_1682_),
    .C(_1133_),
    .A(_1626_),
    .Y(_1140_));
 sg13g2_a21oi_1 _4015_ (.A1(_1626_),
    .A2(_1133_),
    .Y(_1141_),
    .B1(_1682_));
 sg13g2_nor2_1 _4016_ (.A(net681),
    .B(_1141_),
    .Y(_1142_));
 sg13g2_a21oi_1 _4017_ (.A1(_1140_),
    .A2(_1142_),
    .Y(_1143_),
    .B1(net695));
 sg13g2_o21ai_1 _4018_ (.B1(_1143_),
    .Y(_1144_),
    .A1(net325),
    .A2(net746));
 sg13g2_a21oi_1 _4019_ (.A1(_1139_),
    .A2(_1144_),
    .Y(_0158_),
    .B1(net819));
 sg13g2_a22oi_1 _4020_ (.Y(_1145_),
    .B1(_1130_),
    .B2(net325),
    .A2(_0697_),
    .A1(net659));
 sg13g2_or2_1 _4021_ (.X(_1146_),
    .B(_1145_),
    .A(net790));
 sg13g2_a21oi_1 _4022_ (.A1(_1627_),
    .A2(_1133_),
    .Y(_1147_),
    .B1(_1461_));
 sg13g2_xnor2_1 _4023_ (.Y(_1148_),
    .A(_1623_),
    .B(_1147_));
 sg13g2_o21ai_1 _4024_ (.B1(net790),
    .Y(_1149_),
    .A1(\collatz.iter[83] ),
    .A2(net753));
 sg13g2_a21o_1 _4025_ (.A2(_1148_),
    .A1(net753),
    .B1(_1149_),
    .X(_1150_));
 sg13g2_a21oi_1 _4026_ (.A1(_1146_),
    .A2(_1150_),
    .Y(_0159_),
    .B1(net819));
 sg13g2_a22oi_1 _4027_ (.Y(_1151_),
    .B1(_1130_),
    .B2(\collatz.iter[83] ),
    .A2(_0704_),
    .A1(net660));
 sg13g2_or2_1 _4028_ (.X(_1152_),
    .B(_1151_),
    .A(net792));
 sg13g2_a21oi_1 _4029_ (.A1(_1623_),
    .A2(_1147_),
    .Y(_1153_),
    .B1(_1622_));
 sg13g2_xor2_1 _4030_ (.B(_1153_),
    .A(_1624_),
    .X(_1154_));
 sg13g2_a21oi_1 _4031_ (.A1(net746),
    .A2(_1154_),
    .Y(_1155_),
    .B1(net695));
 sg13g2_o21ai_1 _4032_ (.B1(_1155_),
    .Y(_1156_),
    .A1(\collatz.iter[84] ),
    .A2(net753));
 sg13g2_a21oi_1 _4033_ (.A1(_1152_),
    .A2(_1156_),
    .Y(_0160_),
    .B1(net824));
 sg13g2_a22oi_1 _4034_ (.Y(_1157_),
    .B1(_1130_),
    .B2(\collatz.iter[84] ),
    .A2(_0711_),
    .A1(net659));
 sg13g2_or2_1 _4035_ (.X(_1158_),
    .B(_1157_),
    .A(net792));
 sg13g2_a21oi_1 _4036_ (.A1(_1683_),
    .A2(_1132_),
    .Y(_1159_),
    .B1(_1629_));
 sg13g2_or2_1 _4037_ (.X(_1160_),
    .B(_1159_),
    .A(_1620_));
 sg13g2_xnor2_1 _4038_ (.Y(_1161_),
    .A(_1620_),
    .B(_1159_));
 sg13g2_o21ai_1 _4039_ (.B1(net792),
    .Y(_1162_),
    .A1(net700),
    .A2(net746));
 sg13g2_a21o_1 _4040_ (.A2(_1161_),
    .A1(net746),
    .B1(_1162_),
    .X(_1163_));
 sg13g2_a21oi_1 _4041_ (.A1(_1158_),
    .A2(_1163_),
    .Y(_0161_),
    .B1(net819));
 sg13g2_a22oi_1 _4042_ (.Y(_1164_),
    .B1(_1130_),
    .B2(net700),
    .A2(_0720_),
    .A1(net659));
 sg13g2_or2_1 _4043_ (.X(_1165_),
    .B(_1164_),
    .A(net792));
 sg13g2_nand2_1 _4044_ (.Y(_1166_),
    .A(_1619_),
    .B(_1160_));
 sg13g2_xnor2_1 _4045_ (.Y(_1167_),
    .A(_1618_),
    .B(_1166_));
 sg13g2_a21oi_1 _4046_ (.A1(_1403_),
    .A2(net681),
    .Y(_1168_),
    .B1(net695));
 sg13g2_o21ai_1 _4047_ (.B1(_1168_),
    .Y(_1169_),
    .A1(net681),
    .A2(_1167_));
 sg13g2_a21oi_1 _4048_ (.A1(_1165_),
    .A2(_1169_),
    .Y(_0162_),
    .B1(net819));
 sg13g2_a22oi_1 _4049_ (.Y(_1170_),
    .B1(_1130_),
    .B2(\collatz.iter[86] ),
    .A2(_0727_),
    .A1(net659));
 sg13g2_or2_1 _4050_ (.X(_1171_),
    .B(_1170_),
    .A(net792));
 sg13g2_a21oi_1 _4051_ (.A1(_1631_),
    .A2(_1160_),
    .Y(_1172_),
    .B1(_1462_));
 sg13g2_nor2b_1 _4052_ (.A(_1616_),
    .B_N(_1172_),
    .Y(_1173_));
 sg13g2_xor2_1 _4053_ (.B(_1172_),
    .A(_1616_),
    .X(_1174_));
 sg13g2_o21ai_1 _4054_ (.B1(net792),
    .Y(_1175_),
    .A1(\collatz.iter[87] ),
    .A2(net747));
 sg13g2_a21o_1 _4055_ (.A2(_1174_),
    .A1(net747),
    .B1(_1175_),
    .X(_1176_));
 sg13g2_a21oi_1 _4056_ (.A1(_1171_),
    .A2(_1176_),
    .Y(_0163_),
    .B1(net819));
 sg13g2_a22oi_1 _4057_ (.Y(_1177_),
    .B1(_1130_),
    .B2(\collatz.iter[87] ),
    .A2(_0734_),
    .A1(net659));
 sg13g2_or2_1 _4058_ (.X(_1178_),
    .B(_1177_),
    .A(net792));
 sg13g2_a21oi_1 _4059_ (.A1(\collatz.iter[86] ),
    .A2(net700),
    .Y(_1179_),
    .B1(_1173_));
 sg13g2_xnor2_1 _4060_ (.Y(_1180_),
    .A(_1617_),
    .B(_1179_));
 sg13g2_a21oi_1 _4061_ (.A1(net747),
    .A2(_1180_),
    .Y(_1181_),
    .B1(net690));
 sg13g2_o21ai_1 _4062_ (.B1(_1181_),
    .Y(_1182_),
    .A1(net299),
    .A2(net747));
 sg13g2_a21oi_1 _4063_ (.A1(_1178_),
    .A2(_1182_),
    .Y(_0164_),
    .B1(net819));
 sg13g2_a21oi_2 _4064_ (.B1(net651),
    .Y(_1183_),
    .A2(net675),
    .A1(net658));
 sg13g2_a22oi_1 _4065_ (.Y(_1184_),
    .B1(_1183_),
    .B2(net299),
    .A2(_0743_),
    .A1(net660));
 sg13g2_or2_1 _4066_ (.X(_1185_),
    .B(_1184_),
    .A(net791));
 sg13g2_a21oi_2 _4067_ (.B1(_1634_),
    .Y(_1186_),
    .A2(_1132_),
    .A1(_1684_));
 sg13g2_or2_1 _4068_ (.X(_1187_),
    .B(_1186_),
    .A(_1612_));
 sg13g2_xnor2_1 _4069_ (.Y(_1188_),
    .A(_1612_),
    .B(_1186_));
 sg13g2_o21ai_1 _4070_ (.B1(net791),
    .Y(_1189_),
    .A1(\collatz.iter[89] ),
    .A2(net744));
 sg13g2_a21o_1 _4071_ (.A2(_1188_),
    .A1(net744),
    .B1(_1189_),
    .X(_1190_));
 sg13g2_a21oi_1 _4072_ (.A1(_1185_),
    .A2(_1190_),
    .Y(_0165_),
    .B1(net818));
 sg13g2_a22oi_1 _4073_ (.Y(_1191_),
    .B1(_1183_),
    .B2(\collatz.iter[89] ),
    .A2(_0751_),
    .A1(net658));
 sg13g2_or2_1 _4074_ (.X(_1192_),
    .B(_1191_),
    .A(net794));
 sg13g2_nand2_1 _4075_ (.Y(_1193_),
    .A(_1603_),
    .B(_1187_));
 sg13g2_xnor2_1 _4076_ (.Y(_1194_),
    .A(_1611_),
    .B(_1193_));
 sg13g2_a21oi_1 _4077_ (.A1(net744),
    .A2(_1194_),
    .Y(_1195_),
    .B1(net690));
 sg13g2_o21ai_1 _4078_ (.B1(_1195_),
    .Y(_1196_),
    .A1(net319),
    .A2(net744));
 sg13g2_a21oi_1 _4079_ (.A1(_1192_),
    .A2(_1196_),
    .Y(_0166_),
    .B1(net818));
 sg13g2_a22oi_1 _4080_ (.Y(_1197_),
    .B1(_1183_),
    .B2(net319),
    .A2(_0758_),
    .A1(net658));
 sg13g2_or2_1 _4081_ (.X(_1198_),
    .B(_1197_),
    .A(net791));
 sg13g2_a21oi_1 _4082_ (.A1(_1604_),
    .A2(_1187_),
    .Y(_1199_),
    .B1(_1448_));
 sg13g2_nor2b_1 _4083_ (.A(_1601_),
    .B_N(_1199_),
    .Y(_1200_));
 sg13g2_xor2_1 _4084_ (.B(_1199_),
    .A(_1601_),
    .X(_1201_));
 sg13g2_o21ai_1 _4085_ (.B1(net791),
    .Y(_1202_),
    .A1(\collatz.iter[91] ),
    .A2(net743));
 sg13g2_a21o_1 _4086_ (.A2(_1201_),
    .A1(net743),
    .B1(_1202_),
    .X(_1203_));
 sg13g2_a21oi_1 _4087_ (.A1(_1198_),
    .A2(_1203_),
    .Y(_0167_),
    .B1(net818));
 sg13g2_a22oi_1 _4088_ (.Y(_1204_),
    .B1(_1183_),
    .B2(\collatz.iter[91] ),
    .A2(_0765_),
    .A1(net658));
 sg13g2_or2_1 _4089_ (.X(_1205_),
    .B(_1204_),
    .A(net778));
 sg13g2_a21oi_1 _4090_ (.A1(\collatz.iter[90] ),
    .A2(\collatz.iter[89] ),
    .Y(_1206_),
    .B1(_1200_));
 sg13g2_xnor2_1 _4091_ (.Y(_1207_),
    .A(_1602_),
    .B(_1206_));
 sg13g2_a21oi_1 _4092_ (.A1(net743),
    .A2(_1207_),
    .Y(_1208_),
    .B1(net690));
 sg13g2_o21ai_1 _4093_ (.B1(_1208_),
    .Y(_1209_),
    .A1(net274),
    .A2(net743));
 sg13g2_a21oi_1 _4094_ (.A1(_1205_),
    .A2(_1209_),
    .Y(_0168_),
    .B1(net815));
 sg13g2_a22oi_1 _4095_ (.Y(_1210_),
    .B1(_1183_),
    .B2(net274),
    .A2(_0772_),
    .A1(net658));
 sg13g2_or2_1 _4096_ (.X(_1211_),
    .B(_1210_),
    .A(net778));
 sg13g2_o21ai_1 _4097_ (.B1(_1607_),
    .Y(_1212_),
    .A1(_1614_),
    .A2(_1186_));
 sg13g2_nand2_1 _4098_ (.Y(_1213_),
    .A(_1598_),
    .B(_1212_));
 sg13g2_xnor2_1 _4099_ (.Y(_1214_),
    .A(_1598_),
    .B(_1212_));
 sg13g2_o21ai_1 _4100_ (.B1(net778),
    .Y(_1215_),
    .A1(\collatz.iter[93] ),
    .A2(net736));
 sg13g2_a21o_1 _4101_ (.A2(_1214_),
    .A1(net735),
    .B1(_1215_),
    .X(_1216_));
 sg13g2_a21oi_1 _4102_ (.A1(_1211_),
    .A2(_1216_),
    .Y(_0169_),
    .B1(net815));
 sg13g2_a22oi_1 _4103_ (.Y(_1217_),
    .B1(_1183_),
    .B2(net290),
    .A2(_0780_),
    .A1(net658));
 sg13g2_or2_1 _4104_ (.X(_1218_),
    .B(_1217_),
    .A(net778));
 sg13g2_nand2_1 _4105_ (.Y(_1219_),
    .A(_1596_),
    .B(_1213_));
 sg13g2_xnor2_1 _4106_ (.Y(_1220_),
    .A(_1599_),
    .B(_1219_));
 sg13g2_a21oi_1 _4107_ (.A1(net736),
    .A2(_1220_),
    .Y(_1221_),
    .B1(net689));
 sg13g2_o21ai_1 _4108_ (.B1(_1221_),
    .Y(_1222_),
    .A1(net313),
    .A2(net735));
 sg13g2_a21oi_1 _4109_ (.A1(_1218_),
    .A2(_1222_),
    .Y(_0170_),
    .B1(net813));
 sg13g2_a22oi_1 _4110_ (.Y(_1223_),
    .B1(_1183_),
    .B2(net313),
    .A2(_0787_),
    .A1(net658));
 sg13g2_or2_1 _4111_ (.X(_1224_),
    .B(_1223_),
    .A(net778));
 sg13g2_a21oi_1 _4112_ (.A1(_1597_),
    .A2(_1213_),
    .Y(_1225_),
    .B1(_1437_));
 sg13g2_xnor2_1 _4113_ (.Y(_1226_),
    .A(_1592_),
    .B(_1225_));
 sg13g2_o21ai_1 _4114_ (.B1(net778),
    .Y(_1227_),
    .A1(\collatz.iter[95] ),
    .A2(net736));
 sg13g2_a21o_1 _4115_ (.A2(_1226_),
    .A1(net734),
    .B1(_1227_),
    .X(_1228_));
 sg13g2_a21oi_1 _4116_ (.A1(_1224_),
    .A2(_1228_),
    .Y(_0171_),
    .B1(net813));
 sg13g2_a22oi_1 _4117_ (.Y(_1229_),
    .B1(_1183_),
    .B2(\collatz.iter[95] ),
    .A2(_0795_),
    .A1(net658));
 sg13g2_or2_1 _4118_ (.X(_1230_),
    .B(_1229_),
    .A(net779));
 sg13g2_a21oi_1 _4119_ (.A1(_1592_),
    .A2(_1225_),
    .Y(_1231_),
    .B1(_1591_));
 sg13g2_xor2_1 _4120_ (.B(_1231_),
    .A(_1593_),
    .X(_1232_));
 sg13g2_a21oi_1 _4121_ (.A1(net734),
    .A2(_1232_),
    .Y(_1233_),
    .B1(net689));
 sg13g2_o21ai_1 _4122_ (.B1(_1233_),
    .Y(_1234_),
    .A1(net311),
    .A2(net737));
 sg13g2_a21oi_1 _4123_ (.A1(_1230_),
    .A2(_1234_),
    .Y(_0172_),
    .B1(net814));
 sg13g2_a21oi_2 _4124_ (.B1(net650),
    .Y(_1235_),
    .A2(net674),
    .A1(net656));
 sg13g2_nand2_1 _4125_ (.Y(_1236_),
    .A(\collatz.iter[96] ),
    .B(_1235_));
 sg13g2_nand3_1 _4126_ (.B(net657),
    .C(_0807_),
    .A(net844),
    .Y(_1237_));
 sg13g2_a21oi_1 _4127_ (.A1(_1236_),
    .A2(_1237_),
    .Y(_1238_),
    .B1(net776));
 sg13g2_nand2_1 _4128_ (.Y(_1239_),
    .A(_1585_),
    .B(_1896_));
 sg13g2_xnor2_1 _4129_ (.Y(_1240_),
    .A(_1585_),
    .B(_1896_));
 sg13g2_o21ai_1 _4130_ (.B1(net777),
    .Y(_1241_),
    .A1(net699),
    .A2(net737));
 sg13g2_a21oi_1 _4131_ (.A1(net737),
    .A2(_1240_),
    .Y(_1242_),
    .B1(_1241_));
 sg13g2_o21ai_1 _4132_ (.B1(net847),
    .Y(_1243_),
    .A1(_1238_),
    .A2(_1242_));
 sg13g2_inv_1 _4133_ (.Y(_0173_),
    .A(_1243_));
 sg13g2_a22oi_1 _4134_ (.Y(_1244_),
    .B1(_1235_),
    .B2(net699),
    .A2(_0812_),
    .A1(net657));
 sg13g2_or2_1 _4135_ (.X(_1245_),
    .B(_1244_),
    .A(net773));
 sg13g2_nand2_1 _4136_ (.Y(_1246_),
    .A(_1570_),
    .B(_1239_));
 sg13g2_xnor2_1 _4137_ (.Y(_1247_),
    .A(_1586_),
    .B(_1246_));
 sg13g2_a21oi_1 _4138_ (.A1(_1402_),
    .A2(net680),
    .Y(_1248_),
    .B1(net689));
 sg13g2_o21ai_1 _4139_ (.B1(_1248_),
    .Y(_1249_),
    .A1(net680),
    .A2(_1247_));
 sg13g2_a21oi_1 _4140_ (.A1(_1245_),
    .A2(_1249_),
    .Y(_0174_),
    .B1(net814));
 sg13g2_a22oi_1 _4141_ (.Y(_1250_),
    .B1(_1235_),
    .B2(\collatz.iter[98] ),
    .A2(_0819_),
    .A1(net656));
 sg13g2_or2_1 _4142_ (.X(_1251_),
    .B(_1250_),
    .A(net771));
 sg13g2_a21oi_1 _4143_ (.A1(_1571_),
    .A2(_1239_),
    .Y(_1252_),
    .B1(_1453_));
 sg13g2_xnor2_1 _4144_ (.Y(_1253_),
    .A(_1567_),
    .B(_1252_));
 sg13g2_o21ai_1 _4145_ (.B1(net771),
    .Y(_1254_),
    .A1(\collatz.iter[99] ),
    .A2(net724));
 sg13g2_a21o_1 _4146_ (.A2(_1253_),
    .A1(net724),
    .B1(_1254_),
    .X(_1255_));
 sg13g2_a21oi_1 _4147_ (.A1(_1251_),
    .A2(_1255_),
    .Y(_0175_),
    .B1(net810));
 sg13g2_a22oi_1 _4148_ (.Y(_1256_),
    .B1(_1235_),
    .B2(\collatz.iter[99] ),
    .A2(_0826_),
    .A1(net656));
 sg13g2_or2_1 _4149_ (.X(_1257_),
    .B(_1256_),
    .A(net771));
 sg13g2_a21oi_1 _4150_ (.A1(_1567_),
    .A2(_1252_),
    .Y(_1258_),
    .B1(_1566_));
 sg13g2_xnor2_1 _4151_ (.Y(_1259_),
    .A(_1569_),
    .B(_1258_));
 sg13g2_a21oi_1 _4152_ (.A1(net724),
    .A2(_1259_),
    .Y(_1260_),
    .B1(net687));
 sg13g2_o21ai_1 _4153_ (.B1(_1260_),
    .Y(_1261_),
    .A1(net312),
    .A2(net723));
 sg13g2_a21oi_1 _4154_ (.A1(_1257_),
    .A2(_1261_),
    .Y(_0176_),
    .B1(net810));
 sg13g2_a22oi_1 _4155_ (.Y(_1262_),
    .B1(_1235_),
    .B2(net312),
    .A2(_0833_),
    .A1(net656));
 sg13g2_or2_1 _4156_ (.X(_1263_),
    .B(_1262_),
    .A(net771));
 sg13g2_a21oi_2 _4157_ (.B1(_1575_),
    .Y(_1264_),
    .A2(_1896_),
    .A1(_1588_));
 sg13g2_or2_1 _4158_ (.X(_1265_),
    .B(_1264_),
    .A(_1564_));
 sg13g2_xnor2_1 _4159_ (.Y(_1266_),
    .A(_1564_),
    .B(_1264_));
 sg13g2_o21ai_1 _4160_ (.B1(net770),
    .Y(_1267_),
    .A1(\collatz.iter[101] ),
    .A2(net723));
 sg13g2_a21o_1 _4161_ (.A2(_1266_),
    .A1(net723),
    .B1(_1267_),
    .X(_1268_));
 sg13g2_a21oi_1 _4162_ (.A1(_1263_),
    .A2(_1268_),
    .Y(_0177_),
    .B1(net809));
 sg13g2_a22oi_1 _4163_ (.Y(_1269_),
    .B1(_1235_),
    .B2(\collatz.iter[101] ),
    .A2(_0841_),
    .A1(net656));
 sg13g2_or2_1 _4164_ (.X(_1270_),
    .B(_1269_),
    .A(net771));
 sg13g2_nand2_1 _4165_ (.Y(_1271_),
    .A(_1563_),
    .B(_1265_));
 sg13g2_xor2_1 _4166_ (.B(_1271_),
    .A(_1562_),
    .X(_1272_));
 sg13g2_a21oi_1 _4167_ (.A1(net723),
    .A2(_1272_),
    .Y(_1273_),
    .B1(net687));
 sg13g2_o21ai_1 _4168_ (.B1(_1273_),
    .Y(_1274_),
    .A1(\collatz.iter[102] ),
    .A2(net723));
 sg13g2_a21oi_1 _4169_ (.A1(_1270_),
    .A2(_1274_),
    .Y(_0178_),
    .B1(net809));
 sg13g2_a22oi_1 _4170_ (.Y(_1275_),
    .B1(_1235_),
    .B2(\collatz.iter[102] ),
    .A2(_0848_),
    .A1(net656));
 sg13g2_or2_1 _4171_ (.X(_1276_),
    .B(_1275_),
    .A(net770));
 sg13g2_a21oi_1 _4172_ (.A1(_1577_),
    .A2(_1265_),
    .Y(_1277_),
    .B1(_1445_));
 sg13g2_xnor2_1 _4173_ (.Y(_1278_),
    .A(_1558_),
    .B(_1277_));
 sg13g2_o21ai_1 _4174_ (.B1(net771),
    .Y(_1279_),
    .A1(\collatz.iter[103] ),
    .A2(net723));
 sg13g2_a21o_1 _4175_ (.A2(_1278_),
    .A1(net723),
    .B1(_1279_),
    .X(_1280_));
 sg13g2_a21oi_1 _4176_ (.A1(_1276_),
    .A2(_1280_),
    .Y(_0179_),
    .B1(net810));
 sg13g2_a22oi_1 _4177_ (.Y(_1281_),
    .B1(_1235_),
    .B2(\collatz.iter[103] ),
    .A2(_0855_),
    .A1(net656));
 sg13g2_or2_1 _4178_ (.X(_1282_),
    .B(_1281_),
    .A(net771));
 sg13g2_a21oi_1 _4179_ (.A1(_1558_),
    .A2(_1277_),
    .Y(_1283_),
    .B1(_1557_));
 sg13g2_xnor2_1 _4180_ (.Y(_1284_),
    .A(_1561_),
    .B(_1283_));
 sg13g2_a21oi_1 _4181_ (.A1(net724),
    .A2(_1284_),
    .Y(_1285_),
    .B1(net687));
 sg13g2_o21ai_1 _4182_ (.B1(_1285_),
    .Y(_1286_),
    .A1(net329),
    .A2(net723));
 sg13g2_a21oi_1 _4183_ (.A1(_1282_),
    .A2(_1286_),
    .Y(_0180_),
    .B1(net810));
 sg13g2_and3_1 _4184_ (.X(_1287_),
    .A(net829),
    .B(net657),
    .C(_0806_));
 sg13g2_nor2_2 _4185_ (.A(net651),
    .B(net652),
    .Y(_1288_));
 sg13g2_a22oi_1 _4186_ (.Y(_1289_),
    .B1(_1288_),
    .B2(net334),
    .A2(net652),
    .A1(net844));
 sg13g2_or2_1 _4187_ (.X(_1290_),
    .B(_1289_),
    .A(net776));
 sg13g2_a21oi_2 _4188_ (.B1(_1580_),
    .Y(_1291_),
    .A2(_1896_),
    .A1(_1589_));
 sg13g2_nand2b_1 _4189_ (.Y(_1292_),
    .B(_1554_),
    .A_N(_1291_));
 sg13g2_xor2_1 _4190_ (.B(_1291_),
    .A(_1554_),
    .X(_1293_));
 sg13g2_o21ai_1 _4191_ (.B1(net776),
    .Y(_1294_),
    .A1(\collatz.iter[105] ),
    .A2(net737));
 sg13g2_a21o_1 _4192_ (.A2(_1293_),
    .A1(net737),
    .B1(_1294_),
    .X(_1295_));
 sg13g2_a21oi_1 _4193_ (.A1(_1290_),
    .A2(_1295_),
    .Y(_0181_),
    .B1(net814));
 sg13g2_a22oi_1 _4194_ (.Y(_1296_),
    .B1(_1288_),
    .B2(\collatz.iter[105] ),
    .A2(_1287_),
    .A1(net842));
 sg13g2_or2_1 _4195_ (.X(_1297_),
    .B(_1296_),
    .A(net777));
 sg13g2_nand2_1 _4196_ (.Y(_1298_),
    .A(_1547_),
    .B(_1292_));
 sg13g2_xnor2_1 _4197_ (.Y(_1299_),
    .A(_1553_),
    .B(_1298_));
 sg13g2_a21oi_1 _4198_ (.A1(net734),
    .A2(_1299_),
    .Y(_1300_),
    .B1(net689));
 sg13g2_o21ai_1 _4199_ (.B1(_1300_),
    .Y(_1301_),
    .A1(net300),
    .A2(net734));
 sg13g2_a21oi_1 _4200_ (.A1(_1297_),
    .A2(_1301_),
    .Y(_0182_),
    .B1(net813));
 sg13g2_a22oi_1 _4201_ (.Y(_1302_),
    .B1(_1288_),
    .B2(net300),
    .A2(net652),
    .A1(net840));
 sg13g2_or2_1 _4202_ (.X(_1303_),
    .B(_1302_),
    .A(net777));
 sg13g2_a21oi_1 _4203_ (.A1(_1548_),
    .A2(_1292_),
    .Y(_1304_),
    .B1(_1455_));
 sg13g2_xnor2_1 _4204_ (.Y(_1305_),
    .A(_1545_),
    .B(_1304_));
 sg13g2_o21ai_1 _4205_ (.B1(net777),
    .Y(_1306_),
    .A1(\collatz.iter[107] ),
    .A2(net734));
 sg13g2_a21o_1 _4206_ (.A2(_1305_),
    .A1(net734),
    .B1(_1306_),
    .X(_1307_));
 sg13g2_a21oi_1 _4207_ (.A1(_1303_),
    .A2(_1307_),
    .Y(_0183_),
    .B1(net813));
 sg13g2_a22oi_1 _4208_ (.Y(_1308_),
    .B1(_1288_),
    .B2(\collatz.iter[107] ),
    .A2(net652),
    .A1(net838));
 sg13g2_or2_1 _4209_ (.X(_1309_),
    .B(_1308_),
    .A(net777));
 sg13g2_a21oi_1 _4210_ (.A1(_1545_),
    .A2(_1304_),
    .Y(_1310_),
    .B1(_1544_));
 sg13g2_xor2_1 _4211_ (.B(_1310_),
    .A(_1546_),
    .X(_1311_));
 sg13g2_a21oi_1 _4212_ (.A1(net734),
    .A2(_1311_),
    .Y(_1312_),
    .B1(net689));
 sg13g2_o21ai_1 _4213_ (.B1(_1312_),
    .Y(_1313_),
    .A1(net314),
    .A2(net734));
 sg13g2_a21oi_1 _4214_ (.A1(_1309_),
    .A2(_1313_),
    .Y(_0184_),
    .B1(net813));
 sg13g2_a22oi_1 _4215_ (.Y(_1314_),
    .B1(_1288_),
    .B2(net314),
    .A2(net652),
    .A1(net836));
 sg13g2_or2_1 _4216_ (.X(_1315_),
    .B(_1314_),
    .A(net776));
 sg13g2_o21ai_1 _4217_ (.B1(_1551_),
    .Y(_1316_),
    .A1(_1555_),
    .A2(_1291_));
 sg13g2_nand2_1 _4218_ (.Y(_1317_),
    .A(_1541_),
    .B(_1316_));
 sg13g2_xnor2_1 _4219_ (.Y(_1318_),
    .A(_1541_),
    .B(_1316_));
 sg13g2_o21ai_1 _4220_ (.B1(net776),
    .Y(_1319_),
    .A1(\collatz.iter[109] ),
    .A2(net733));
 sg13g2_a21o_1 _4221_ (.A2(_1318_),
    .A1(net733),
    .B1(_1319_),
    .X(_1320_));
 sg13g2_a21oi_1 _4222_ (.A1(_1315_),
    .A2(_1320_),
    .Y(_0185_),
    .B1(net813));
 sg13g2_a22oi_1 _4223_ (.Y(_1321_),
    .B1(_1288_),
    .B2(\collatz.iter[109] ),
    .A2(net652),
    .A1(net834));
 sg13g2_or2_1 _4224_ (.X(_1322_),
    .B(_1321_),
    .A(net776));
 sg13g2_nand2_1 _4225_ (.Y(_1323_),
    .A(_1539_),
    .B(_1317_));
 sg13g2_xnor2_1 _4226_ (.Y(_1324_),
    .A(_1542_),
    .B(_1323_));
 sg13g2_a21oi_1 _4227_ (.A1(net730),
    .A2(_1324_),
    .Y(_1325_),
    .B1(net688));
 sg13g2_o21ai_1 _4228_ (.B1(_1325_),
    .Y(_1326_),
    .A1(net306),
    .A2(net730));
 sg13g2_a21oi_1 _4229_ (.A1(_1322_),
    .A2(_1326_),
    .Y(_0186_),
    .B1(net811));
 sg13g2_a22oi_1 _4230_ (.Y(_1327_),
    .B1(_1288_),
    .B2(net306),
    .A2(net652),
    .A1(net832));
 sg13g2_or2_1 _4231_ (.X(_1328_),
    .B(_1327_),
    .A(net776));
 sg13g2_a21oi_1 _4232_ (.A1(_1540_),
    .A2(_1317_),
    .Y(_1329_),
    .B1(_1460_));
 sg13g2_xnor2_1 _4233_ (.Y(_1330_),
    .A(_1535_),
    .B(_1329_));
 sg13g2_o21ai_1 _4234_ (.B1(net776),
    .Y(_1331_),
    .A1(\collatz.iter[111] ),
    .A2(net730));
 sg13g2_a21o_1 _4235_ (.A2(_1330_),
    .A1(net730),
    .B1(_1331_),
    .X(_1332_));
 sg13g2_a21oi_1 _4236_ (.A1(_1328_),
    .A2(_1332_),
    .Y(_0187_),
    .B1(net811));
 sg13g2_a22oi_1 _4237_ (.Y(_1333_),
    .B1(_1288_),
    .B2(\collatz.iter[111] ),
    .A2(net652),
    .A1(net830));
 sg13g2_or2_1 _4238_ (.X(_1334_),
    .B(_1333_),
    .A(net767));
 sg13g2_a21oi_1 _4239_ (.A1(_1535_),
    .A2(_1329_),
    .Y(_1335_),
    .B1(_1534_));
 sg13g2_xor2_1 _4240_ (.B(_1335_),
    .A(_1536_),
    .X(_1336_));
 sg13g2_a21oi_1 _4241_ (.A1(net730),
    .A2(_1336_),
    .Y(_1337_),
    .B1(net688));
 sg13g2_o21ai_1 _4242_ (.B1(_1337_),
    .Y(_1338_),
    .A1(\collatz.iter[112] ),
    .A2(net731));
 sg13g2_a21oi_1 _4243_ (.A1(_1334_),
    .A2(_1338_),
    .Y(_0188_),
    .B1(net811));
 sg13g2_a22oi_1 _4244_ (.Y(_1339_),
    .B1(_0916_),
    .B2(net654),
    .A2(_1517_),
    .A1(\collatz.iter[112] ));
 sg13g2_or2_1 _4245_ (.X(_1340_),
    .B(_1339_),
    .A(net764));
 sg13g2_xnor2_1 _4246_ (.Y(_1341_),
    .A(_1533_),
    .B(_1897_));
 sg13g2_o21ai_1 _4247_ (.B1(net764),
    .Y(_1342_),
    .A1(net698),
    .A2(net717));
 sg13g2_a21o_1 _4248_ (.A2(_1341_),
    .A1(net717),
    .B1(_1342_),
    .X(_1343_));
 sg13g2_a21oi_1 _4249_ (.A1(_1340_),
    .A2(_1343_),
    .Y(_0189_),
    .B1(net807));
 sg13g2_a22oi_1 _4250_ (.Y(_1344_),
    .B1(_0924_),
    .B2(net654),
    .A2(_1517_),
    .A1(net698));
 sg13g2_or2_1 _4251_ (.X(_1345_),
    .B(_1344_),
    .A(net762));
 sg13g2_xnor2_1 _4252_ (.Y(_1346_),
    .A(_1901_),
    .B(_1930_));
 sg13g2_a21oi_1 _4253_ (.A1(net717),
    .A2(_1346_),
    .Y(_1347_),
    .B1(net685));
 sg13g2_o21ai_1 _4254_ (.B1(_1347_),
    .Y(_1348_),
    .A1(net330),
    .A2(net713));
 sg13g2_a21oi_1 _4255_ (.A1(_1345_),
    .A2(_1348_),
    .Y(_0190_),
    .B1(net805));
 sg13g2_a22oi_1 _4256_ (.Y(_1349_),
    .B1(_0931_),
    .B2(net654),
    .A2(_1517_),
    .A1(\collatz.iter[114] ));
 sg13g2_or2_1 _4257_ (.X(_1350_),
    .B(_1349_),
    .A(net762));
 sg13g2_xnor2_1 _4258_ (.Y(_1351_),
    .A(_1902_),
    .B(_1903_));
 sg13g2_o21ai_1 _4259_ (.B1(net762),
    .Y(_1352_),
    .A1(net697),
    .A2(net713));
 sg13g2_a21o_1 _4260_ (.A2(_1351_),
    .A1(net713),
    .B1(_1352_),
    .X(_1353_));
 sg13g2_a21oi_1 _4261_ (.A1(_1350_),
    .A2(_1353_),
    .Y(_0191_),
    .B1(net805));
 sg13g2_a22oi_1 _4262_ (.Y(_1354_),
    .B1(_0938_),
    .B2(net654),
    .A2(_1517_),
    .A1(net697));
 sg13g2_or2_1 _4263_ (.X(_1355_),
    .B(_1354_),
    .A(net762));
 sg13g2_xor2_1 _4264_ (.B(_1906_),
    .A(_1905_),
    .X(_1356_));
 sg13g2_a21oi_1 _4265_ (.A1(net712),
    .A2(_1356_),
    .Y(_1357_),
    .B1(net684));
 sg13g2_o21ai_1 _4266_ (.B1(_1357_),
    .Y(_1358_),
    .A1(net310),
    .A2(net712));
 sg13g2_a21oi_1 _4267_ (.A1(_1355_),
    .A2(_1358_),
    .Y(_0192_),
    .B1(net805));
 sg13g2_a22oi_1 _4268_ (.Y(_1359_),
    .B1(_0945_),
    .B2(net654),
    .A2(_1517_),
    .A1(net333));
 sg13g2_or2_1 _4269_ (.X(_1360_),
    .B(_1359_),
    .A(net760));
 sg13g2_xor2_1 _4270_ (.B(_1907_),
    .A(_1527_),
    .X(_1361_));
 sg13g2_o21ai_1 _4271_ (.B1(net760),
    .Y(_1362_),
    .A1(\collatz.iter[117] ),
    .A2(net712));
 sg13g2_a21o_1 _4272_ (.A2(_1361_),
    .A1(net712),
    .B1(_1362_),
    .X(_1363_));
 sg13g2_a21oi_1 _4273_ (.A1(_1360_),
    .A2(_1363_),
    .Y(_0193_),
    .B1(net805));
 sg13g2_a22oi_1 _4274_ (.Y(_1364_),
    .B1(_0954_),
    .B2(net654),
    .A2(_1517_),
    .A1(\collatz.iter[117] ));
 sg13g2_or2_1 _4275_ (.X(_1365_),
    .B(_1364_),
    .A(net760));
 sg13g2_and2_1 _4276_ (.A(_1524_),
    .B(_1908_),
    .X(_1366_));
 sg13g2_xnor2_1 _4277_ (.Y(_1367_),
    .A(_1922_),
    .B(_1366_));
 sg13g2_a21oi_1 _4278_ (.A1(net712),
    .A2(_1367_),
    .Y(_1368_),
    .B1(net684));
 sg13g2_o21ai_1 _4279_ (.B1(_1368_),
    .Y(_1369_),
    .A1(net303),
    .A2(net712));
 sg13g2_a21oi_1 _4280_ (.A1(_1365_),
    .A2(_1369_),
    .Y(_0194_),
    .B1(net805));
 sg13g2_a22oi_1 _4281_ (.Y(_1370_),
    .B1(_0961_),
    .B2(net654),
    .A2(_1517_),
    .A1(\collatz.iter[118] ));
 sg13g2_or2_1 _4282_ (.X(_1371_),
    .B(_1370_),
    .A(net760));
 sg13g2_xnor2_1 _4283_ (.Y(_1372_),
    .A(_1523_),
    .B(_1909_));
 sg13g2_o21ai_1 _4284_ (.B1(net760),
    .Y(_1373_),
    .A1(\collatz.iter[119] ),
    .A2(net713));
 sg13g2_a21o_1 _4285_ (.A2(_1372_),
    .A1(net713),
    .B1(_1373_),
    .X(_1374_));
 sg13g2_a21oi_1 _4286_ (.A1(_1371_),
    .A2(_1374_),
    .Y(_0195_),
    .B1(net805));
 sg13g2_dfrbp_1 _4287_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net63),
    .D(_0011_),
    .Q_N(_2142_),
    .Q(\collatz.iter[119] ));
 sg13g2_dfrbp_1 _4288_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net170),
    .D(_0012_),
    .Q_N(_2141_),
    .Q(\collatz.iter[120] ));
 sg13g2_dfrbp_1 _4289_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net169),
    .D(_0013_),
    .Q_N(_2140_),
    .Q(\collatz.iter[121] ));
 sg13g2_dfrbp_1 _4290_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net168),
    .D(_0014_),
    .Q_N(_2139_),
    .Q(\collatz.iter[122] ));
 sg13g2_dfrbp_1 _4291_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net167),
    .D(_0015_),
    .Q_N(_2138_),
    .Q(\collatz.iter[123] ));
 sg13g2_dfrbp_1 _4292_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net166),
    .D(_0016_),
    .Q_N(_2137_),
    .Q(\collatz.iter[124] ));
 sg13g2_dfrbp_1 _4293_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net165),
    .D(_0017_),
    .Q_N(_2136_),
    .Q(\collatz.iter[125] ));
 sg13g2_dfrbp_1 _4294_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net164),
    .D(_0018_),
    .Q_N(_2135_),
    .Q(\collatz.iter[126] ));
 sg13g2_dfrbp_1 _4295_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net163),
    .D(_0019_),
    .Q_N(_2134_),
    .Q(\collatz.iter[127] ));
 sg13g2_dfrbp_1 _4296_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net162),
    .D(_0020_),
    .Q_N(_2133_),
    .Q(\collatz.iter[128] ));
 sg13g2_dfrbp_1 _4297_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net161),
    .D(_0021_),
    .Q_N(_0007_),
    .Q(\collatz.iter[129] ));
 sg13g2_dfrbp_1 _4298_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net160),
    .D(_0022_),
    .Q_N(_0006_),
    .Q(\collatz.iter[130] ));
 sg13g2_dfrbp_1 _4299_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net159),
    .D(net272),
    .Q_N(_2132_),
    .Q(\collatz.iter[131] ));
 sg13g2_dfrbp_1 _4300_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net158),
    .D(_0024_),
    .Q_N(_0005_),
    .Q(\collatz.iter[132] ));
 sg13g2_dfrbp_1 _4301_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net157),
    .D(_0025_),
    .Q_N(_2131_),
    .Q(\collatz.iter[133] ));
 sg13g2_dfrbp_1 _4302_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net156),
    .D(_0026_),
    .Q_N(_0004_),
    .Q(\collatz.iter[134] ));
 sg13g2_dfrbp_1 _4303_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net155),
    .D(_0027_),
    .Q_N(_2130_),
    .Q(\collatz.iter[135] ));
 sg13g2_dfrbp_1 _4304_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net154),
    .D(_0028_),
    .Q_N(_0003_),
    .Q(\collatz.iter[136] ));
 sg13g2_dfrbp_1 _4305_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net153),
    .D(_0029_),
    .Q_N(_2129_),
    .Q(\collatz.iter[137] ));
 sg13g2_dfrbp_1 _4306_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net152),
    .D(_0030_),
    .Q_N(_0002_),
    .Q(\collatz.iter[138] ));
 sg13g2_dfrbp_1 _4307_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net151),
    .D(_0031_),
    .Q_N(_2128_),
    .Q(\collatz.iter[139] ));
 sg13g2_dfrbp_1 _4308_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net150),
    .D(_0032_),
    .Q_N(_0001_),
    .Q(\collatz.iter[140] ));
 sg13g2_dfrbp_1 _4309_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net149),
    .D(_0033_),
    .Q_N(_2127_),
    .Q(\collatz.iter[141] ));
 sg13g2_dfrbp_1 _4310_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net148),
    .D(_0034_),
    .Q_N(_0000_),
    .Q(\collatz.iter[142] ));
 sg13g2_dfrbp_1 _4311_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net147),
    .D(_0035_),
    .Q_N(_2126_),
    .Q(\collatz.iter[143] ));
 sg13g2_dfrbp_1 _4312_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net146),
    .D(_0036_),
    .Q_N(_0010_),
    .Q(\collatz.comp ));
 sg13g2_dfrbp_1 _4313_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net144),
    .D(_0037_),
    .Q_N(_2125_),
    .Q(\collatz.orbit_len[0] ));
 sg13g2_dfrbp_1 _4314_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net142),
    .D(net212),
    .Q_N(_2124_),
    .Q(\collatz.orbit_len[1] ));
 sg13g2_dfrbp_1 _4315_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net140),
    .D(_0039_),
    .Q_N(_2123_),
    .Q(\collatz.orbit_len[2] ));
 sg13g2_dfrbp_1 _4316_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net138),
    .D(_0040_),
    .Q_N(_2122_),
    .Q(\collatz.orbit_len[3] ));
 sg13g2_dfrbp_1 _4317_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net136),
    .D(_0041_),
    .Q_N(_2121_),
    .Q(\collatz.orbit_len[4] ));
 sg13g2_dfrbp_1 _4318_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net134),
    .D(_0042_),
    .Q_N(_2120_),
    .Q(\collatz.orbit_len[5] ));
 sg13g2_dfrbp_1 _4319_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net132),
    .D(_0043_),
    .Q_N(_2119_),
    .Q(\collatz.orbit_len[6] ));
 sg13g2_dfrbp_1 _4320_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net130),
    .D(_0044_),
    .Q_N(_2118_),
    .Q(\collatz.orbit_len[7] ));
 sg13g2_dfrbp_1 _4321_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net128),
    .D(_0045_),
    .Q_N(_2117_),
    .Q(\collatz.orbit_len[8] ));
 sg13g2_dfrbp_1 _4322_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net126),
    .D(_0046_),
    .Q_N(_2116_),
    .Q(\collatz.orbit_len[9] ));
 sg13g2_dfrbp_1 _4323_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net124),
    .D(_0047_),
    .Q_N(_2115_),
    .Q(\collatz.orbit_len[10] ));
 sg13g2_dfrbp_1 _4324_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net122),
    .D(net221),
    .Q_N(_2114_),
    .Q(\collatz.orbit_len[11] ));
 sg13g2_dfrbp_1 _4325_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net120),
    .D(_0049_),
    .Q_N(_2113_),
    .Q(\collatz.orbit_len[12] ));
 sg13g2_dfrbp_1 _4326_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net118),
    .D(_0050_),
    .Q_N(_2112_),
    .Q(\collatz.orbit_len[13] ));
 sg13g2_dfrbp_1 _4327_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net116),
    .D(_0051_),
    .Q_N(_2111_),
    .Q(\collatz.orbit_len[14] ));
 sg13g2_dfrbp_1 _4328_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net114),
    .D(net230),
    .Q_N(_2110_),
    .Q(\collatz.orbit_len[15] ));
 sg13g2_dfrbp_1 _4329_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net112),
    .D(_0053_),
    .Q_N(_2109_),
    .Q(\collatz.path_record_h16[0] ));
 sg13g2_dfrbp_1 _4330_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net110),
    .D(_0054_),
    .Q_N(_2108_),
    .Q(\collatz.path_record_h16[1] ));
 sg13g2_dfrbp_1 _4331_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net108),
    .D(_0055_),
    .Q_N(_2107_),
    .Q(\collatz.path_record_h16[2] ));
 sg13g2_dfrbp_1 _4332_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net106),
    .D(_0056_),
    .Q_N(_2106_),
    .Q(\collatz.path_record_h16[3] ));
 sg13g2_dfrbp_1 _4333_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net104),
    .D(_0057_),
    .Q_N(_2105_),
    .Q(\collatz.path_record_h16[4] ));
 sg13g2_dfrbp_1 _4334_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net102),
    .D(_0058_),
    .Q_N(_2104_),
    .Q(\collatz.path_record_h16[5] ));
 sg13g2_dfrbp_1 _4335_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net100),
    .D(_0059_),
    .Q_N(_2103_),
    .Q(\collatz.path_record_h16[6] ));
 sg13g2_dfrbp_1 _4336_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net98),
    .D(_0060_),
    .Q_N(_2102_),
    .Q(\collatz.path_record_h16[7] ));
 sg13g2_dfrbp_1 _4337_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net96),
    .D(_0061_),
    .Q_N(_2101_),
    .Q(\collatz.path_record_h16[8] ));
 sg13g2_dfrbp_1 _4338_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net94),
    .D(_0062_),
    .Q_N(_2100_),
    .Q(\collatz.path_record_h16[9] ));
 sg13g2_dfrbp_1 _4339_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net92),
    .D(_0063_),
    .Q_N(_2099_),
    .Q(\collatz.path_record_h16[10] ));
 sg13g2_dfrbp_1 _4340_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net90),
    .D(_0064_),
    .Q_N(_2098_),
    .Q(\collatz.path_record_h16[11] ));
 sg13g2_dfrbp_1 _4341_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net88),
    .D(_0065_),
    .Q_N(_2097_),
    .Q(\collatz.path_record_h16[12] ));
 sg13g2_dfrbp_1 _4342_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net86),
    .D(_0066_),
    .Q_N(_2096_),
    .Q(\collatz.path_record_h16[13] ));
 sg13g2_dfrbp_1 _4343_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net84),
    .D(_0067_),
    .Q_N(_2095_),
    .Q(\collatz.path_record_h16[14] ));
 sg13g2_dfrbp_1 _4344_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net82),
    .D(_0068_),
    .Q_N(_0008_),
    .Q(\collatz.path_record_h16[15] ));
 sg13g2_dfrbp_1 _4345_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net80),
    .D(_0069_),
    .Q_N(_2094_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _4346_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net78),
    .D(_0070_),
    .Q_N(_2093_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _4347_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net76),
    .D(_0071_),
    .Q_N(_2092_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _4348_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net74),
    .D(_0072_),
    .Q_N(_2091_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _4349_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net72),
    .D(_0073_),
    .Q_N(_2090_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _4350_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net70),
    .D(_0074_),
    .Q_N(_2089_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _4351_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net68),
    .D(_0075_),
    .Q_N(_2088_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _4352_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net66),
    .D(_0076_),
    .Q_N(_2087_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _4353_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net64),
    .D(net209),
    .Q_N(_2086_),
    .Q(\collatz.iter[1] ));
 sg13g2_dfrbp_1 _4354_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net62),
    .D(_0078_),
    .Q_N(_0009_),
    .Q(\collatz.iter[0] ));
 sg13g2_dfrbp_1 _4355_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net61),
    .D(_0079_),
    .Q_N(_2085_),
    .Q(\collatz.iter[2] ));
 sg13g2_dfrbp_1 _4356_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net60),
    .D(net292),
    .Q_N(_2084_),
    .Q(\collatz.iter[3] ));
 sg13g2_dfrbp_1 _4357_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net59),
    .D(_0081_),
    .Q_N(_2083_),
    .Q(\collatz.iter[4] ));
 sg13g2_dfrbp_1 _4358_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net58),
    .D(_0082_),
    .Q_N(_2082_),
    .Q(\collatz.iter[5] ));
 sg13g2_dfrbp_1 _4359_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net57),
    .D(net285),
    .Q_N(_2081_),
    .Q(\collatz.iter[6] ));
 sg13g2_dfrbp_1 _4360_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net56),
    .D(_0084_),
    .Q_N(_2080_),
    .Q(\collatz.iter[7] ));
 sg13g2_dfrbp_1 _4361_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net55),
    .D(_0085_),
    .Q_N(_2079_),
    .Q(\collatz.iter[8] ));
 sg13g2_dfrbp_1 _4362_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net54),
    .D(_0086_),
    .Q_N(_2078_),
    .Q(\collatz.iter[9] ));
 sg13g2_dfrbp_1 _4363_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net53),
    .D(_0087_),
    .Q_N(_2077_),
    .Q(\collatz.iter[10] ));
 sg13g2_dfrbp_1 _4364_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net52),
    .D(_0088_),
    .Q_N(_2076_),
    .Q(\collatz.iter[11] ));
 sg13g2_dfrbp_1 _4365_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net51),
    .D(_0089_),
    .Q_N(_2075_),
    .Q(\collatz.iter[12] ));
 sg13g2_dfrbp_1 _4366_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net50),
    .D(_0090_),
    .Q_N(_2074_),
    .Q(\collatz.iter[13] ));
 sg13g2_dfrbp_1 _4367_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net49),
    .D(_0091_),
    .Q_N(_2073_),
    .Q(\collatz.iter[14] ));
 sg13g2_dfrbp_1 _4368_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net48),
    .D(_0092_),
    .Q_N(_2072_),
    .Q(\collatz.iter[15] ));
 sg13g2_dfrbp_1 _4369_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net47),
    .D(_0093_),
    .Q_N(_2071_),
    .Q(\collatz.iter[16] ));
 sg13g2_dfrbp_1 _4370_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net46),
    .D(_0094_),
    .Q_N(_2070_),
    .Q(\collatz.iter[17] ));
 sg13g2_dfrbp_1 _4371_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net45),
    .D(_0095_),
    .Q_N(_2069_),
    .Q(\collatz.iter[18] ));
 sg13g2_dfrbp_1 _4372_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net44),
    .D(_0096_),
    .Q_N(_2068_),
    .Q(\collatz.iter[19] ));
 sg13g2_dfrbp_1 _4373_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net43),
    .D(_0097_),
    .Q_N(_2067_),
    .Q(\collatz.iter[20] ));
 sg13g2_dfrbp_1 _4374_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net42),
    .D(_0098_),
    .Q_N(_2066_),
    .Q(\collatz.iter[21] ));
 sg13g2_dfrbp_1 _4375_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net41),
    .D(_0099_),
    .Q_N(_2065_),
    .Q(\collatz.iter[22] ));
 sg13g2_dfrbp_1 _4376_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net40),
    .D(_0100_),
    .Q_N(_2064_),
    .Q(\collatz.iter[23] ));
 sg13g2_dfrbp_1 _4377_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net39),
    .D(_0101_),
    .Q_N(_2063_),
    .Q(\collatz.iter[24] ));
 sg13g2_dfrbp_1 _4378_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net38),
    .D(_0102_),
    .Q_N(_2062_),
    .Q(\collatz.iter[25] ));
 sg13g2_dfrbp_1 _4379_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net37),
    .D(_0103_),
    .Q_N(_2061_),
    .Q(\collatz.iter[26] ));
 sg13g2_dfrbp_1 _4380_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net36),
    .D(_0104_),
    .Q_N(_2060_),
    .Q(\collatz.iter[27] ));
 sg13g2_dfrbp_1 _4381_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net35),
    .D(_0105_),
    .Q_N(_2059_),
    .Q(\collatz.iter[28] ));
 sg13g2_dfrbp_1 _4382_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net34),
    .D(_0106_),
    .Q_N(_2058_),
    .Q(\collatz.iter[29] ));
 sg13g2_dfrbp_1 _4383_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net33),
    .D(_0107_),
    .Q_N(_2057_),
    .Q(\collatz.iter[30] ));
 sg13g2_dfrbp_1 _4384_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net32),
    .D(_0108_),
    .Q_N(_2056_),
    .Q(\collatz.iter[31] ));
 sg13g2_dfrbp_1 _4385_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net31),
    .D(_0109_),
    .Q_N(_2055_),
    .Q(\collatz.iter[32] ));
 sg13g2_dfrbp_1 _4386_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net30),
    .D(_0110_),
    .Q_N(_2054_),
    .Q(\collatz.iter[33] ));
 sg13g2_dfrbp_1 _4387_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net29),
    .D(_0111_),
    .Q_N(_2053_),
    .Q(\collatz.iter[34] ));
 sg13g2_dfrbp_1 _4388_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net28),
    .D(_0112_),
    .Q_N(_2052_),
    .Q(\collatz.iter[35] ));
 sg13g2_dfrbp_1 _4389_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net27),
    .D(_0113_),
    .Q_N(_2051_),
    .Q(\collatz.iter[36] ));
 sg13g2_dfrbp_1 _4390_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net26),
    .D(_0114_),
    .Q_N(_2050_),
    .Q(\collatz.iter[37] ));
 sg13g2_dfrbp_1 _4391_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net25),
    .D(_0115_),
    .Q_N(_2049_),
    .Q(\collatz.iter[38] ));
 sg13g2_dfrbp_1 _4392_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net24),
    .D(_0116_),
    .Q_N(_2048_),
    .Q(\collatz.iter[39] ));
 sg13g2_dfrbp_1 _4393_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net23),
    .D(_0117_),
    .Q_N(_2047_),
    .Q(\collatz.iter[40] ));
 sg13g2_dfrbp_1 _4394_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net22),
    .D(_0118_),
    .Q_N(_2046_),
    .Q(\collatz.iter[41] ));
 sg13g2_dfrbp_1 _4395_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net206),
    .D(_0119_),
    .Q_N(_2045_),
    .Q(\collatz.iter[42] ));
 sg13g2_dfrbp_1 _4396_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net205),
    .D(_0120_),
    .Q_N(_2044_),
    .Q(\collatz.iter[43] ));
 sg13g2_dfrbp_1 _4397_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net204),
    .D(_0121_),
    .Q_N(_2043_),
    .Q(\collatz.iter[44] ));
 sg13g2_dfrbp_1 _4398_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net203),
    .D(_0122_),
    .Q_N(_2042_),
    .Q(\collatz.iter[45] ));
 sg13g2_dfrbp_1 _4399_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net202),
    .D(_0123_),
    .Q_N(_2041_),
    .Q(\collatz.iter[46] ));
 sg13g2_dfrbp_1 _4400_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net201),
    .D(_0124_),
    .Q_N(_2040_),
    .Q(\collatz.iter[47] ));
 sg13g2_dfrbp_1 _4401_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net200),
    .D(_0125_),
    .Q_N(_2039_),
    .Q(\collatz.iter[48] ));
 sg13g2_dfrbp_1 _4402_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net199),
    .D(_0126_),
    .Q_N(_2038_),
    .Q(\collatz.iter[49] ));
 sg13g2_dfrbp_1 _4403_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net198),
    .D(_0127_),
    .Q_N(_2037_),
    .Q(\collatz.iter[50] ));
 sg13g2_dfrbp_1 _4404_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net197),
    .D(_0128_),
    .Q_N(_2036_),
    .Q(\collatz.iter[51] ));
 sg13g2_dfrbp_1 _4405_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net196),
    .D(_0129_),
    .Q_N(_2035_),
    .Q(\collatz.iter[52] ));
 sg13g2_dfrbp_1 _4406_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net195),
    .D(net265),
    .Q_N(_2034_),
    .Q(\collatz.iter[53] ));
 sg13g2_dfrbp_1 _4407_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net194),
    .D(_0131_),
    .Q_N(_2033_),
    .Q(\collatz.iter[54] ));
 sg13g2_dfrbp_1 _4408_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net193),
    .D(_0132_),
    .Q_N(_2032_),
    .Q(\collatz.iter[55] ));
 sg13g2_dfrbp_1 _4409_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net192),
    .D(_0133_),
    .Q_N(_2031_),
    .Q(\collatz.iter[56] ));
 sg13g2_dfrbp_1 _4410_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net191),
    .D(_0134_),
    .Q_N(_2030_),
    .Q(\collatz.iter[57] ));
 sg13g2_dfrbp_1 _4411_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net190),
    .D(_0135_),
    .Q_N(_2029_),
    .Q(\collatz.iter[58] ));
 sg13g2_dfrbp_1 _4412_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net189),
    .D(_0136_),
    .Q_N(_2028_),
    .Q(\collatz.iter[59] ));
 sg13g2_dfrbp_1 _4413_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net188),
    .D(_0137_),
    .Q_N(_2027_),
    .Q(\collatz.iter[60] ));
 sg13g2_dfrbp_1 _4414_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net187),
    .D(_0138_),
    .Q_N(_2026_),
    .Q(\collatz.iter[61] ));
 sg13g2_dfrbp_1 _4415_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net186),
    .D(_0139_),
    .Q_N(_2025_),
    .Q(\collatz.iter[62] ));
 sg13g2_dfrbp_1 _4416_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net185),
    .D(_0140_),
    .Q_N(_2024_),
    .Q(\collatz.iter[63] ));
 sg13g2_dfrbp_1 _4417_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net184),
    .D(_0141_),
    .Q_N(_2023_),
    .Q(\collatz.iter[64] ));
 sg13g2_dfrbp_1 _4418_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net183),
    .D(net279),
    .Q_N(_2022_),
    .Q(\collatz.iter[65] ));
 sg13g2_dfrbp_1 _4419_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net182),
    .D(_0143_),
    .Q_N(_2021_),
    .Q(\collatz.iter[66] ));
 sg13g2_dfrbp_1 _4420_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net181),
    .D(net281),
    .Q_N(_2020_),
    .Q(\collatz.iter[67] ));
 sg13g2_dfrbp_1 _4421_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net180),
    .D(_0145_),
    .Q_N(_2019_),
    .Q(\collatz.iter[68] ));
 sg13g2_dfrbp_1 _4422_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net179),
    .D(net283),
    .Q_N(_2018_),
    .Q(\collatz.iter[69] ));
 sg13g2_dfrbp_1 _4423_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net178),
    .D(_0147_),
    .Q_N(_2017_),
    .Q(\collatz.iter[70] ));
 sg13g2_dfrbp_1 _4424_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net177),
    .D(net270),
    .Q_N(_2016_),
    .Q(\collatz.iter[71] ));
 sg13g2_dfrbp_1 _4425_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net176),
    .D(_0149_),
    .Q_N(_2015_),
    .Q(\collatz.iter[72] ));
 sg13g2_dfrbp_1 _4426_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net175),
    .D(net287),
    .Q_N(_2014_),
    .Q(\collatz.iter[73] ));
 sg13g2_dfrbp_1 _4427_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net174),
    .D(_0151_),
    .Q_N(_2013_),
    .Q(\collatz.iter[74] ));
 sg13g2_dfrbp_1 _4428_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net173),
    .D(net296),
    .Q_N(_2012_),
    .Q(\collatz.iter[75] ));
 sg13g2_dfrbp_1 _4429_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net172),
    .D(_0153_),
    .Q_N(_2011_),
    .Q(\collatz.iter[76] ));
 sg13g2_dfrbp_1 _4430_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net171),
    .D(net294),
    .Q_N(_2010_),
    .Q(\collatz.iter[77] ));
 sg13g2_dfrbp_1 _4431_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net145),
    .D(_0155_),
    .Q_N(_2009_),
    .Q(\collatz.iter[78] ));
 sg13g2_dfrbp_1 _4432_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net143),
    .D(_0156_),
    .Q_N(_2008_),
    .Q(\collatz.iter[79] ));
 sg13g2_dfrbp_1 _4433_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net141),
    .D(_0157_),
    .Q_N(_2007_),
    .Q(\collatz.iter[80] ));
 sg13g2_dfrbp_1 _4434_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net139),
    .D(_0158_),
    .Q_N(_2006_),
    .Q(\collatz.iter[81] ));
 sg13g2_dfrbp_1 _4435_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net137),
    .D(_0159_),
    .Q_N(_2005_),
    .Q(\collatz.iter[82] ));
 sg13g2_dfrbp_1 _4436_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net135),
    .D(_0160_),
    .Q_N(_2004_),
    .Q(\collatz.iter[83] ));
 sg13g2_dfrbp_1 _4437_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net133),
    .D(_0161_),
    .Q_N(_2003_),
    .Q(\collatz.iter[84] ));
 sg13g2_dfrbp_1 _4438_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net131),
    .D(_0162_),
    .Q_N(_2002_),
    .Q(\collatz.iter[85] ));
 sg13g2_dfrbp_1 _4439_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net129),
    .D(_0163_),
    .Q_N(_2001_),
    .Q(\collatz.iter[86] ));
 sg13g2_dfrbp_1 _4440_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net127),
    .D(_0164_),
    .Q_N(_2000_),
    .Q(\collatz.iter[87] ));
 sg13g2_dfrbp_1 _4441_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net125),
    .D(_0165_),
    .Q_N(_1999_),
    .Q(\collatz.iter[88] ));
 sg13g2_dfrbp_1 _4442_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net123),
    .D(_0166_),
    .Q_N(_1998_),
    .Q(\collatz.iter[89] ));
 sg13g2_dfrbp_1 _4443_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net121),
    .D(_0167_),
    .Q_N(_1997_),
    .Q(\collatz.iter[90] ));
 sg13g2_dfrbp_1 _4444_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net119),
    .D(net275),
    .Q_N(_1996_),
    .Q(\collatz.iter[91] ));
 sg13g2_dfrbp_1 _4445_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net117),
    .D(_0169_),
    .Q_N(_1995_),
    .Q(\collatz.iter[92] ));
 sg13g2_dfrbp_1 _4446_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net115),
    .D(_0170_),
    .Q_N(_1994_),
    .Q(\collatz.iter[93] ));
 sg13g2_dfrbp_1 _4447_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net113),
    .D(_0171_),
    .Q_N(_1993_),
    .Q(\collatz.iter[94] ));
 sg13g2_dfrbp_1 _4448_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net111),
    .D(_0172_),
    .Q_N(_1992_),
    .Q(\collatz.iter[95] ));
 sg13g2_dfrbp_1 _4449_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net109),
    .D(_0173_),
    .Q_N(_1991_),
    .Q(\collatz.iter[96] ));
 sg13g2_dfrbp_1 _4450_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net107),
    .D(_0174_),
    .Q_N(_1990_),
    .Q(\collatz.iter[97] ));
 sg13g2_dfrbp_1 _4451_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net105),
    .D(_0175_),
    .Q_N(_1989_),
    .Q(\collatz.iter[98] ));
 sg13g2_dfrbp_1 _4452_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net103),
    .D(_0176_),
    .Q_N(_1988_),
    .Q(\collatz.iter[99] ));
 sg13g2_dfrbp_1 _4453_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net101),
    .D(_0177_),
    .Q_N(_1987_),
    .Q(\collatz.iter[100] ));
 sg13g2_dfrbp_1 _4454_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net99),
    .D(_0178_),
    .Q_N(_1986_),
    .Q(\collatz.iter[101] ));
 sg13g2_dfrbp_1 _4455_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net97),
    .D(_0179_),
    .Q_N(_1985_),
    .Q(\collatz.iter[102] ));
 sg13g2_dfrbp_1 _4456_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net95),
    .D(_0180_),
    .Q_N(_1984_),
    .Q(\collatz.iter[103] ));
 sg13g2_dfrbp_1 _4457_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net93),
    .D(_0181_),
    .Q_N(_1983_),
    .Q(\collatz.iter[104] ));
 sg13g2_dfrbp_1 _4458_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net91),
    .D(_0182_),
    .Q_N(_1982_),
    .Q(\collatz.iter[105] ));
 sg13g2_dfrbp_1 _4459_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net89),
    .D(_0183_),
    .Q_N(_1981_),
    .Q(\collatz.iter[106] ));
 sg13g2_dfrbp_1 _4460_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net87),
    .D(_0184_),
    .Q_N(_1980_),
    .Q(\collatz.iter[107] ));
 sg13g2_dfrbp_1 _4461_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net85),
    .D(_0185_),
    .Q_N(_1979_),
    .Q(\collatz.iter[108] ));
 sg13g2_dfrbp_1 _4462_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net83),
    .D(net307),
    .Q_N(_1978_),
    .Q(\collatz.iter[109] ));
 sg13g2_dfrbp_1 _4463_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net81),
    .D(_0187_),
    .Q_N(_1977_),
    .Q(\collatz.iter[110] ));
 sg13g2_dfrbp_1 _4464_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net79),
    .D(_0188_),
    .Q_N(_1976_),
    .Q(\collatz.iter[111] ));
 sg13g2_dfrbp_1 _4465_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net77),
    .D(_0189_),
    .Q_N(_1975_),
    .Q(\collatz.iter[112] ));
 sg13g2_dfrbp_1 _4466_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net75),
    .D(_0190_),
    .Q_N(_1974_),
    .Q(\collatz.iter[113] ));
 sg13g2_dfrbp_1 _4467_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net73),
    .D(_0191_),
    .Q_N(_1973_),
    .Q(\collatz.iter[114] ));
 sg13g2_dfrbp_1 _4468_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net71),
    .D(_0192_),
    .Q_N(_1972_),
    .Q(\collatz.iter[115] ));
 sg13g2_dfrbp_1 _4469_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net69),
    .D(_0193_),
    .Q_N(_1971_),
    .Q(\collatz.iter[116] ));
 sg13g2_dfrbp_1 _4470_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net67),
    .D(_0194_),
    .Q_N(_1970_),
    .Q(\collatz.iter[117] ));
 sg13g2_dfrbp_1 _4471_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net65),
    .D(_0195_),
    .Q_N(_1969_),
    .Q(\collatz.iter[118] ));
 sg13g2_tiehi _4393__23 (.L_HI(net23));
 sg13g2_tiehi _4392__24 (.L_HI(net24));
 sg13g2_tiehi _4391__25 (.L_HI(net25));
 sg13g2_tiehi _4390__26 (.L_HI(net26));
 sg13g2_tiehi _4389__27 (.L_HI(net27));
 sg13g2_tiehi _4388__28 (.L_HI(net28));
 sg13g2_tiehi _4387__29 (.L_HI(net29));
 sg13g2_tiehi _4386__30 (.L_HI(net30));
 sg13g2_tiehi _4385__31 (.L_HI(net31));
 sg13g2_tiehi _4384__32 (.L_HI(net32));
 sg13g2_tiehi _4383__33 (.L_HI(net33));
 sg13g2_tiehi _4382__34 (.L_HI(net34));
 sg13g2_tiehi _4381__35 (.L_HI(net35));
 sg13g2_tiehi _4380__36 (.L_HI(net36));
 sg13g2_tiehi _4379__37 (.L_HI(net37));
 sg13g2_tiehi _4378__38 (.L_HI(net38));
 sg13g2_tiehi _4377__39 (.L_HI(net39));
 sg13g2_tiehi _4376__40 (.L_HI(net40));
 sg13g2_tiehi _4375__41 (.L_HI(net41));
 sg13g2_tiehi _4374__42 (.L_HI(net42));
 sg13g2_tiehi _4373__43 (.L_HI(net43));
 sg13g2_tiehi _4372__44 (.L_HI(net44));
 sg13g2_tiehi _4371__45 (.L_HI(net45));
 sg13g2_tiehi _4370__46 (.L_HI(net46));
 sg13g2_tiehi _4369__47 (.L_HI(net47));
 sg13g2_tiehi _4368__48 (.L_HI(net48));
 sg13g2_tiehi _4367__49 (.L_HI(net49));
 sg13g2_tiehi _4366__50 (.L_HI(net50));
 sg13g2_tiehi _4365__51 (.L_HI(net51));
 sg13g2_tiehi _4364__52 (.L_HI(net52));
 sg13g2_tiehi _4363__53 (.L_HI(net53));
 sg13g2_tiehi _4362__54 (.L_HI(net54));
 sg13g2_tiehi _4361__55 (.L_HI(net55));
 sg13g2_tiehi _4360__56 (.L_HI(net56));
 sg13g2_tiehi _4359__57 (.L_HI(net57));
 sg13g2_tiehi _4358__58 (.L_HI(net58));
 sg13g2_tiehi _4357__59 (.L_HI(net59));
 sg13g2_tiehi _4356__60 (.L_HI(net60));
 sg13g2_tiehi _4355__61 (.L_HI(net61));
 sg13g2_tiehi _4354__62 (.L_HI(net62));
 sg13g2_tiehi _4287__63 (.L_HI(net63));
 sg13g2_tiehi _4353__64 (.L_HI(net64));
 sg13g2_tiehi _4471__65 (.L_HI(net65));
 sg13g2_tiehi _4352__66 (.L_HI(net66));
 sg13g2_tiehi _4470__67 (.L_HI(net67));
 sg13g2_tiehi _4351__68 (.L_HI(net68));
 sg13g2_tiehi _4469__69 (.L_HI(net69));
 sg13g2_tiehi _4350__70 (.L_HI(net70));
 sg13g2_tiehi _4468__71 (.L_HI(net71));
 sg13g2_tiehi _4349__72 (.L_HI(net72));
 sg13g2_tiehi _4467__73 (.L_HI(net73));
 sg13g2_tiehi _4348__74 (.L_HI(net74));
 sg13g2_tiehi _4466__75 (.L_HI(net75));
 sg13g2_tiehi _4347__76 (.L_HI(net76));
 sg13g2_tiehi _4465__77 (.L_HI(net77));
 sg13g2_tiehi _4346__78 (.L_HI(net78));
 sg13g2_tiehi _4464__79 (.L_HI(net79));
 sg13g2_tiehi _4345__80 (.L_HI(net80));
 sg13g2_tiehi _4463__81 (.L_HI(net81));
 sg13g2_tiehi _4344__82 (.L_HI(net82));
 sg13g2_tiehi _4462__83 (.L_HI(net83));
 sg13g2_tiehi _4343__84 (.L_HI(net84));
 sg13g2_tiehi _4461__85 (.L_HI(net85));
 sg13g2_tiehi _4342__86 (.L_HI(net86));
 sg13g2_tiehi _4460__87 (.L_HI(net87));
 sg13g2_tiehi _4341__88 (.L_HI(net88));
 sg13g2_tiehi _4459__89 (.L_HI(net89));
 sg13g2_tiehi _4340__90 (.L_HI(net90));
 sg13g2_tiehi _4458__91 (.L_HI(net91));
 sg13g2_tiehi _4339__92 (.L_HI(net92));
 sg13g2_tiehi _4457__93 (.L_HI(net93));
 sg13g2_tiehi _4338__94 (.L_HI(net94));
 sg13g2_tiehi _4456__95 (.L_HI(net95));
 sg13g2_tiehi _4337__96 (.L_HI(net96));
 sg13g2_tiehi _4455__97 (.L_HI(net97));
 sg13g2_tiehi _4336__98 (.L_HI(net98));
 sg13g2_tiehi _4454__99 (.L_HI(net99));
 sg13g2_tiehi _4335__100 (.L_HI(net100));
 sg13g2_tiehi _4453__101 (.L_HI(net101));
 sg13g2_tiehi _4334__102 (.L_HI(net102));
 sg13g2_tiehi _4452__103 (.L_HI(net103));
 sg13g2_tiehi _4333__104 (.L_HI(net104));
 sg13g2_tiehi _4451__105 (.L_HI(net105));
 sg13g2_tiehi _4332__106 (.L_HI(net106));
 sg13g2_tiehi _4450__107 (.L_HI(net107));
 sg13g2_tiehi _4331__108 (.L_HI(net108));
 sg13g2_tiehi _4449__109 (.L_HI(net109));
 sg13g2_tiehi _4330__110 (.L_HI(net110));
 sg13g2_tiehi _4448__111 (.L_HI(net111));
 sg13g2_tiehi _4329__112 (.L_HI(net112));
 sg13g2_tiehi _4447__113 (.L_HI(net113));
 sg13g2_tiehi _4328__114 (.L_HI(net114));
 sg13g2_tiehi _4446__115 (.L_HI(net115));
 sg13g2_tiehi _4327__116 (.L_HI(net116));
 sg13g2_tiehi _4445__117 (.L_HI(net117));
 sg13g2_tiehi _4326__118 (.L_HI(net118));
 sg13g2_tiehi _4444__119 (.L_HI(net119));
 sg13g2_tiehi _4325__120 (.L_HI(net120));
 sg13g2_tiehi _4443__121 (.L_HI(net121));
 sg13g2_tiehi _4324__122 (.L_HI(net122));
 sg13g2_tiehi _4442__123 (.L_HI(net123));
 sg13g2_tiehi _4323__124 (.L_HI(net124));
 sg13g2_tiehi _4441__125 (.L_HI(net125));
 sg13g2_tiehi _4322__126 (.L_HI(net126));
 sg13g2_tiehi _4440__127 (.L_HI(net127));
 sg13g2_tiehi _4321__128 (.L_HI(net128));
 sg13g2_tiehi _4439__129 (.L_HI(net129));
 sg13g2_tiehi _4320__130 (.L_HI(net130));
 sg13g2_tiehi _4438__131 (.L_HI(net131));
 sg13g2_tiehi _4319__132 (.L_HI(net132));
 sg13g2_tiehi _4437__133 (.L_HI(net133));
 sg13g2_tiehi _4318__134 (.L_HI(net134));
 sg13g2_tiehi _4436__135 (.L_HI(net135));
 sg13g2_tiehi _4317__136 (.L_HI(net136));
 sg13g2_tiehi _4435__137 (.L_HI(net137));
 sg13g2_tiehi _4316__138 (.L_HI(net138));
 sg13g2_tiehi _4434__139 (.L_HI(net139));
 sg13g2_tiehi _4315__140 (.L_HI(net140));
 sg13g2_tiehi _4433__141 (.L_HI(net141));
 sg13g2_tiehi _4314__142 (.L_HI(net142));
 sg13g2_tiehi _4432__143 (.L_HI(net143));
 sg13g2_tiehi _4313__144 (.L_HI(net144));
 sg13g2_tiehi _4431__145 (.L_HI(net145));
 sg13g2_tiehi _4312__146 (.L_HI(net146));
 sg13g2_tiehi _4311__147 (.L_HI(net147));
 sg13g2_tiehi _4310__148 (.L_HI(net148));
 sg13g2_tiehi _4309__149 (.L_HI(net149));
 sg13g2_tiehi _4308__150 (.L_HI(net150));
 sg13g2_tiehi _4307__151 (.L_HI(net151));
 sg13g2_tiehi _4306__152 (.L_HI(net152));
 sg13g2_tiehi _4305__153 (.L_HI(net153));
 sg13g2_tiehi _4304__154 (.L_HI(net154));
 sg13g2_tiehi _4303__155 (.L_HI(net155));
 sg13g2_tiehi _4302__156 (.L_HI(net156));
 sg13g2_tiehi _4301__157 (.L_HI(net157));
 sg13g2_tiehi _4300__158 (.L_HI(net158));
 sg13g2_tiehi _4299__159 (.L_HI(net159));
 sg13g2_tiehi _4298__160 (.L_HI(net160));
 sg13g2_tiehi _4297__161 (.L_HI(net161));
 sg13g2_tiehi _4296__162 (.L_HI(net162));
 sg13g2_tiehi _4295__163 (.L_HI(net163));
 sg13g2_tiehi _4294__164 (.L_HI(net164));
 sg13g2_tiehi _4293__165 (.L_HI(net165));
 sg13g2_tiehi _4292__166 (.L_HI(net166));
 sg13g2_tiehi _4291__167 (.L_HI(net167));
 sg13g2_tiehi _4290__168 (.L_HI(net168));
 sg13g2_tiehi _4289__169 (.L_HI(net169));
 sg13g2_tiehi _4288__170 (.L_HI(net170));
 sg13g2_tiehi _4430__171 (.L_HI(net171));
 sg13g2_tiehi _4429__172 (.L_HI(net172));
 sg13g2_tiehi _4428__173 (.L_HI(net173));
 sg13g2_tiehi _4427__174 (.L_HI(net174));
 sg13g2_tiehi _4426__175 (.L_HI(net175));
 sg13g2_tiehi _4425__176 (.L_HI(net176));
 sg13g2_tiehi _4424__177 (.L_HI(net177));
 sg13g2_tiehi _4423__178 (.L_HI(net178));
 sg13g2_tiehi _4422__179 (.L_HI(net179));
 sg13g2_tiehi _4421__180 (.L_HI(net180));
 sg13g2_tiehi _4420__181 (.L_HI(net181));
 sg13g2_tiehi _4419__182 (.L_HI(net182));
 sg13g2_tiehi _4418__183 (.L_HI(net183));
 sg13g2_tiehi _4417__184 (.L_HI(net184));
 sg13g2_tiehi _4416__185 (.L_HI(net185));
 sg13g2_tiehi _4415__186 (.L_HI(net186));
 sg13g2_tiehi _4414__187 (.L_HI(net187));
 sg13g2_tiehi _4413__188 (.L_HI(net188));
 sg13g2_tiehi _4412__189 (.L_HI(net189));
 sg13g2_tiehi _4411__190 (.L_HI(net190));
 sg13g2_tiehi _4410__191 (.L_HI(net191));
 sg13g2_tiehi _4409__192 (.L_HI(net192));
 sg13g2_tiehi _4408__193 (.L_HI(net193));
 sg13g2_tiehi _4407__194 (.L_HI(net194));
 sg13g2_tiehi _4406__195 (.L_HI(net195));
 sg13g2_tiehi _4405__196 (.L_HI(net196));
 sg13g2_tiehi _4404__197 (.L_HI(net197));
 sg13g2_tiehi _4403__198 (.L_HI(net198));
 sg13g2_tiehi _4402__199 (.L_HI(net199));
 sg13g2_tiehi _4401__200 (.L_HI(net200));
 sg13g2_tiehi _4400__201 (.L_HI(net201));
 sg13g2_tiehi _4399__202 (.L_HI(net202));
 sg13g2_tiehi _4398__203 (.L_HI(net203));
 sg13g2_tiehi _4397__204 (.L_HI(net204));
 sg13g2_tiehi _4396__205 (.L_HI(net205));
 sg13g2_tiehi _4395__206 (.L_HI(net206));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_rtfb_collatz_9 (.L_LO(net9));
 sg13g2_tielo tt_um_rtfb_collatz_10 (.L_LO(net10));
 sg13g2_tielo tt_um_rtfb_collatz_11 (.L_LO(net11));
 sg13g2_tielo tt_um_rtfb_collatz_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rtfb_collatz_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rtfb_collatz_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rtfb_collatz_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rtfb_collatz_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rtfb_collatz_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rtfb_collatz_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rtfb_collatz_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rtfb_collatz_20 (.L_LO(net20));
 sg13g2_tielo tt_um_rtfb_collatz_21 (.L_LO(net21));
 sg13g2_tiehi _4394__22 (.L_HI(net22));
 sg13g2_buf_1 _4671_ (.A(net788),
    .X(uio_oe[7]));
 sg13g2_buf_2 _4672_ (.A(\collatz.busy ),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout645 (.A(net649),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(net649),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(net649),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(net649),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_0514_),
    .X(net649));
 sg13g2_buf_8 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_8 fanout651 (.A(_1508_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_1287_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_1076_),
    .X(net653));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(net655));
 sg13g2_buf_2 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(net657));
 sg13g2_buf_4 fanout657 (.X(net657),
    .A(_1516_));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(net660));
 sg13g2_buf_2 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_1516_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_0862_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_1515_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_1025_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(net666),
    .X(net665));
 sg13g2_buf_4 fanout666 (.X(net666),
    .A(net667));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(net670));
 sg13g2_buf_2 fanout668 (.A(net670),
    .X(net668));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(net670));
 sg13g2_buf_4 fanout670 (.X(net670),
    .A(_0683_));
 sg13g2_buf_2 fanout671 (.A(_0565_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_0546_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_0434_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_0807_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_0741_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_0684_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_0348_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_1509_),
    .X(net679));
 sg13g2_buf_4 fanout680 (.X(net680),
    .A(net683));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(net683));
 sg13g2_buf_2 fanout682 (.A(net683),
    .X(net682));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(_1413_));
 sg13g2_buf_2 fanout684 (.A(net687),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(net687),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(net696),
    .X(net687));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(net696));
 sg13g2_buf_2 fanout689 (.A(net696),
    .X(net689));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(net691));
 sg13g2_buf_4 fanout691 (.X(net691),
    .A(net695));
 sg13g2_buf_4 fanout692 (.X(net692),
    .A(net694));
 sg13g2_buf_2 fanout693 (.A(net694),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_4 fanout696 (.X(net696),
    .A(_1391_));
 sg13g2_buf_2 fanout697 (.A(\collatz.iter[115] ),
    .X(net697));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(\collatz.iter[113] ));
 sg13g2_buf_2 fanout699 (.A(\collatz.iter[97] ),
    .X(net699));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(\collatz.iter[85] ));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(\collatz.iter[81] ));
 sg13g2_buf_2 fanout702 (.A(\collatz.iter[61] ),
    .X(net702));
 sg13g2_buf_4 fanout703 (.X(net703),
    .A(\collatz.iter[53] ));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(net263));
 sg13g2_buf_4 fanout705 (.X(net705),
    .A(\collatz.iter[51] ));
 sg13g2_buf_2 fanout706 (.A(\collatz.iter[45] ),
    .X(net706));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(\collatz.iter[41] ));
 sg13g2_buf_2 fanout708 (.A(\collatz.iter[37] ),
    .X(net708));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(net276));
 sg13g2_buf_2 fanout710 (.A(\collatz.iter[25] ),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(\collatz.iter[3] ),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(net720),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(net720));
 sg13g2_buf_2 fanout714 (.A(net716),
    .X(net714));
 sg13g2_buf_1 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(net720),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(net719),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(net719),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(net720),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(net728),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(net722),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(net728),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(net727),
    .X(net723));
 sg13g2_buf_1 fanout724 (.A(net727),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(net727),
    .X(net725));
 sg13g2_buf_1 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_1 fanout727 (.A(net728),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(\collatz.iter[0] ),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(net731),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(net731),
    .X(net730));
 sg13g2_buf_1 fanout731 (.A(net738),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(net738),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(net738),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(net736),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(net736),
    .X(net735));
 sg13g2_buf_1 fanout736 (.A(net738),
    .X(net736));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(net738));
 sg13g2_buf_2 fanout738 (.A(\collatz.iter[0] ),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(net740),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(net742),
    .X(net740));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(net742));
 sg13g2_buf_2 fanout742 (.A(net759),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(net748),
    .X(net743));
 sg13g2_buf_1 fanout744 (.A(net748),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(net748),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(net748),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(net748),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(net759),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(net750),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(net759),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(net758),
    .X(net751));
 sg13g2_buf_1 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(net758),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(net758),
    .X(net754));
 sg13g2_buf_1 fanout755 (.A(net758),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(net757),
    .X(net756));
 sg13g2_buf_1 fanout757 (.A(net758),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(\collatz.iter[0] ),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(net769),
    .X(net760));
 sg13g2_buf_1 fanout761 (.A(net769),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(net765),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(net765),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(net769),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(net767),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(net769),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(net769),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(net802),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(net771),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(net780),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(net775),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(net775),
    .X(net773));
 sg13g2_buf_1 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(net780),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(net780),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(net779),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(net780),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(net802),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(net782),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(net785),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(net785),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_1 fanout785 (.A(net802),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(net788),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(net802),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(net790),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(net801),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(net794),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(net794),
    .X(net792));
 sg13g2_buf_1 fanout793 (.A(net794),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(net801),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(net797),
    .X(net795));
 sg13g2_buf_4 fanout796 (.X(net796),
    .A(net797));
 sg13g2_buf_2 fanout797 (.A(net801),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(net800),
    .X(net798));
 sg13g2_buf_1 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(net801),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(net802),
    .X(net801));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(\collatz.comp ));
 sg13g2_buf_2 fanout803 (.A(\collatz.iter[125] ),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(_1914_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(net808),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(net808),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(net808),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(net825),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(net810),
    .X(net809));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(net825));
 sg13g2_buf_2 fanout811 (.A(net812),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(net815),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(net814),
    .X(net813));
 sg13g2_buf_4 fanout814 (.X(net814),
    .A(net815));
 sg13g2_buf_2 fanout815 (.A(net825),
    .X(net815));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(net820));
 sg13g2_buf_2 fanout817 (.A(net820),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(net820),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(net820),
    .X(net819));
 sg13g2_buf_1 fanout820 (.A(net825),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(net822),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(net823),
    .X(net822));
 sg13g2_buf_4 fanout823 (.X(net823),
    .A(net824));
 sg13g2_buf_2 fanout824 (.A(net825),
    .X(net824));
 sg13g2_buf_4 fanout825 (.X(net825),
    .A(_1392_));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(net2));
 sg13g2_buf_8 fanout827 (.A(net828),
    .X(net827));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(net829));
 sg13g2_buf_2 fanout829 (.A(uio_in[0]),
    .X(net829));
 sg13g2_buf_4 fanout830 (.X(net830),
    .A(ui_in[7]));
 sg13g2_buf_2 fanout831 (.A(ui_in[7]),
    .X(net831));
 sg13g2_buf_8 fanout832 (.A(ui_in[6]),
    .X(net832));
 sg13g2_buf_4 fanout833 (.X(net833),
    .A(ui_in[6]));
 sg13g2_buf_8 fanout834 (.A(ui_in[5]),
    .X(net834));
 sg13g2_buf_4 fanout835 (.X(net835),
    .A(ui_in[5]));
 sg13g2_buf_8 fanout836 (.A(ui_in[4]),
    .X(net836));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(ui_in[4]));
 sg13g2_buf_8 fanout838 (.A(ui_in[3]),
    .X(net838));
 sg13g2_buf_4 fanout839 (.X(net839),
    .A(ui_in[3]));
 sg13g2_buf_4 fanout840 (.X(net840),
    .A(ui_in[2]));
 sg13g2_buf_2 fanout841 (.A(ui_in[2]),
    .X(net841));
 sg13g2_buf_8 fanout842 (.A(ui_in[1]),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(ui_in[1]),
    .X(net843));
 sg13g2_buf_4 fanout844 (.X(net844),
    .A(ui_in[0]));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(ui_in[0]));
 sg13g2_buf_4 fanout846 (.X(net846),
    .A(net854));
 sg13g2_buf_2 fanout847 (.A(net854),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(net854),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net854),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net853),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(net853),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_4 fanout853 (.X(net853),
    .A(net854));
 sg13g2_buf_2 fanout854 (.A(rst_n),
    .X(net854));
 sg13g2_buf_4 input1 (.X(net1),
    .A(uio_in[1]));
 sg13g2_buf_2 input2 (.A(uio_in[2]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(uio_in[3]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(uio_in[4]),
    .X(net4));
 sg13g2_buf_4 input5 (.X(net5),
    .A(uio_in[5]));
 sg13g2_buf_2 input6 (.A(uio_in[6]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[7]),
    .X(net7));
 sg13g2_tielo tt_um_rtfb_collatz_8 (.L_LO(net8));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0010_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0572_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0077_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold4 (.A(\collatz.orbit_len[1] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0439_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0038_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold7 (.A(\collatz.path_record_h16[15] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold8 (.A(\collatz.path_record_h16[9] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold9 (.A(\collatz.orbit_len[13] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0462_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold11 (.A(\collatz.path_record_h16[7] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold12 (.A(\collatz.path_record_h16[8] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold13 (.A(\collatz.orbit_len[11] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0458_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0048_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold16 (.A(uo_out[7]),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold17 (.A(uo_out[4]),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold18 (.A(\collatz.orbit_len[6] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0448_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold20 (.A(\collatz.orbit_len[2] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0440_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold22 (.A(\collatz.path_record_h16[12] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold23 (.A(\collatz.orbit_len[15] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0052_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold25 (.A(\collatz.orbit_len[3] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0442_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold27 (.A(uo_out[6]),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold28 (.A(\collatz.path_record_h16[14] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold29 (.A(uo_out[3]),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold30 (.A(\collatz.path_record_h16[1] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold31 (.A(uo_out[5]),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold32 (.A(\collatz.orbit_len[5] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0446_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold34 (.A(uo_out[0]),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold35 (.A(\collatz.orbit_len[12] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0461_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold37 (.A(\collatz.orbit_len[8] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0452_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold39 (.A(uo_out[1]),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold40 (.A(\collatz.orbit_len[4] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold41 (.A(\collatz.path_record_h16[6] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold42 (.A(\collatz.path_record_h16[13] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold43 (.A(\collatz.path_record_h16[2] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold44 (.A(uo_out[2]),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold45 (.A(\collatz.orbit_len[10] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0456_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold47 (.A(\collatz.orbit_len[0] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold48 (.A(\collatz.orbit_len[7] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold49 (.A(\collatz.orbit_len[9] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold50 (.A(\collatz.path_record_h16[11] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold51 (.A(\collatz.path_record_h16[3] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold52 (.A(\collatz.path_record_h16[4] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold53 (.A(\collatz.orbit_len[14] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold54 (.A(\collatz.path_record_h16[5] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0006_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold56 (.A(\collatz.path_record_h16[10] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold57 (.A(\collatz.iter[52] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold58 (.A(\collatz.iter[53] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0130_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0004_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold61 (.A(\collatz.iter[64] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0003_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold63 (.A(\collatz.iter[72] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0148_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0005_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0023_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold67 (.A(\collatz.path_record_h16[0] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold68 (.A(\collatz.iter[92] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0168_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold70 (.A(\collatz.iter[33] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0001_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold72 (.A(\collatz.iter[66] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0142_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold74 (.A(\collatz.iter[68] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0144_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold76 (.A(\collatz.iter[70] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0146_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold78 (.A(\collatz.iter[7] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0083_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold80 (.A(\collatz.iter[74] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0150_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold82 (.A(\collatz.iter[38] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold83 (.A(\collatz.iter[62] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold84 (.A(\collatz.iter[93] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold85 (.A(\collatz.iter[4] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0080_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold87 (.A(\collatz.iter[78] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0154_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold89 (.A(\collatz.iter[76] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0152_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold91 (.A(\collatz.iter[28] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold92 (.A(\collatz.iter[126] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold93 (.A(\collatz.iter[88] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold94 (.A(\collatz.iter[106] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0002_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold96 (.A(\collatz.iter[130] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold97 (.A(\collatz.iter[118] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold98 (.A(\collatz.iter[124] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold99 (.A(\collatz.iter[1] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold100 (.A(\collatz.iter[110] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0186_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold102 (.A(\collatz.iter[24] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold103 (.A(\collatz.iter[122] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold104 (.A(\collatz.iter[116] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold105 (.A(\collatz.iter[96] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold106 (.A(\collatz.iter[100] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold107 (.A(\collatz.iter[94] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold108 (.A(\collatz.iter[108] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold109 (.A(\collatz.iter[60] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold110 (.A(\collatz.iter[58] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold111 (.A(\collatz.iter[128] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold112 (.A(\collatz.iter[44] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold113 (.A(\collatz.iter[90] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold114 (.A(\collatz.iter[48] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold115 (.A(\collatz.iter[46] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold116 (.A(\collatz.iter[42] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold117 (.A(\collatz.iter[2] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold118 (.A(\collatz.iter[134] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold119 (.A(\collatz.iter[82] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold120 (.A(\collatz.iter[29] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold121 (.A(\collatz.iter[57] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold122 (.A(\collatz.iter[40] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold123 (.A(\collatz.iter[104] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold124 (.A(\collatz.iter[114] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold125 (.A(\collatz.orbit_len[5] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold126 (.A(\collatz.iter[44] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold127 (.A(\collatz.iter[116] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold128 (.A(\collatz.iter[104] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold129 (.A(\collatz.iter[122] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold130 (.A(\collatz.orbit_len[0] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold131 (.A(\collatz.iter[124] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold132 (.A(\collatz.orbit_len[14] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold133 (.A(\collatz.iter[60] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold134 (.A(\collatz.iter[28] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold135 (.A(\collatz.iter[38] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold136 (.A(\collatz.orbit_len[4] ),
    .X(net342));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_decap_8 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_fill_1 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_311 ();
 sg13g2_decap_8 FILLER_0_318 ();
 sg13g2_decap_8 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_4 FILLER_1_193 ();
 sg13g2_fill_2 FILLER_1_197 ();
 sg13g2_fill_2 FILLER_1_225 ();
 sg13g2_decap_4 FILLER_1_239 ();
 sg13g2_fill_2 FILLER_1_243 ();
 sg13g2_decap_8 FILLER_1_271 ();
 sg13g2_fill_2 FILLER_1_278 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_decap_8 FILLER_1_298 ();
 sg13g2_decap_4 FILLER_1_305 ();
 sg13g2_fill_1 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_314 ();
 sg13g2_decap_8 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_354 ();
 sg13g2_decap_8 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_368 ();
 sg13g2_decap_8 FILLER_1_375 ();
 sg13g2_decap_8 FILLER_1_382 ();
 sg13g2_decap_8 FILLER_1_389 ();
 sg13g2_decap_8 FILLER_1_396 ();
 sg13g2_decap_4 FILLER_1_403 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_fill_1 FILLER_2_161 ();
 sg13g2_fill_2 FILLER_2_214 ();
 sg13g2_fill_1 FILLER_2_216 ();
 sg13g2_fill_2 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_259 ();
 sg13g2_decap_4 FILLER_2_264 ();
 sg13g2_fill_1 FILLER_2_268 ();
 sg13g2_decap_4 FILLER_2_295 ();
 sg13g2_fill_2 FILLER_2_325 ();
 sg13g2_decap_4 FILLER_2_336 ();
 sg13g2_fill_2 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_fill_2 FILLER_3_175 ();
 sg13g2_fill_1 FILLER_3_177 ();
 sg13g2_fill_2 FILLER_3_204 ();
 sg13g2_fill_1 FILLER_3_206 ();
 sg13g2_fill_2 FILLER_3_215 ();
 sg13g2_fill_1 FILLER_3_217 ();
 sg13g2_decap_4 FILLER_3_257 ();
 sg13g2_fill_1 FILLER_3_261 ();
 sg13g2_fill_2 FILLER_3_270 ();
 sg13g2_fill_1 FILLER_3_272 ();
 sg13g2_decap_8 FILLER_3_278 ();
 sg13g2_decap_8 FILLER_3_285 ();
 sg13g2_decap_4 FILLER_3_292 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_4 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_172 ();
 sg13g2_fill_1 FILLER_4_237 ();
 sg13g2_fill_2 FILLER_4_272 ();
 sg13g2_fill_1 FILLER_4_274 ();
 sg13g2_decap_8 FILLER_4_283 ();
 sg13g2_fill_2 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_fill_1 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_fill_1 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_188 ();
 sg13g2_fill_2 FILLER_5_195 ();
 sg13g2_decap_4 FILLER_5_218 ();
 sg13g2_fill_1 FILLER_5_222 ();
 sg13g2_fill_2 FILLER_5_238 ();
 sg13g2_fill_1 FILLER_5_257 ();
 sg13g2_fill_1 FILLER_5_280 ();
 sg13g2_fill_2 FILLER_5_307 ();
 sg13g2_decap_4 FILLER_5_353 ();
 sg13g2_fill_2 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_4 FILLER_6_179 ();
 sg13g2_decap_4 FILLER_6_196 ();
 sg13g2_fill_1 FILLER_6_200 ();
 sg13g2_fill_2 FILLER_6_243 ();
 sg13g2_fill_2 FILLER_6_289 ();
 sg13g2_fill_2 FILLER_6_332 ();
 sg13g2_decap_4 FILLER_6_339 ();
 sg13g2_fill_2 FILLER_6_343 ();
 sg13g2_fill_2 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_4 FILLER_7_140 ();
 sg13g2_fill_1 FILLER_7_144 ();
 sg13g2_fill_1 FILLER_7_171 ();
 sg13g2_fill_2 FILLER_7_193 ();
 sg13g2_fill_2 FILLER_7_221 ();
 sg13g2_decap_8 FILLER_7_240 ();
 sg13g2_fill_2 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_270 ();
 sg13g2_fill_1 FILLER_7_294 ();
 sg13g2_fill_1 FILLER_7_319 ();
 sg13g2_decap_4 FILLER_7_327 ();
 sg13g2_fill_2 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_fill_1 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_170 ();
 sg13g2_fill_2 FILLER_8_207 ();
 sg13g2_fill_1 FILLER_8_209 ();
 sg13g2_fill_2 FILLER_8_232 ();
 sg13g2_fill_1 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_256 ();
 sg13g2_fill_2 FILLER_8_269 ();
 sg13g2_fill_1 FILLER_8_271 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_8 FILLER_8_291 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_fill_2 FILLER_8_357 ();
 sg13g2_fill_1 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_177 ();
 sg13g2_fill_1 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_220 ();
 sg13g2_fill_1 FILLER_9_227 ();
 sg13g2_fill_2 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_4 FILLER_9_273 ();
 sg13g2_fill_2 FILLER_9_277 ();
 sg13g2_fill_1 FILLER_9_305 ();
 sg13g2_fill_2 FILLER_9_329 ();
 sg13g2_fill_1 FILLER_9_346 ();
 sg13g2_fill_2 FILLER_9_352 ();
 sg13g2_fill_2 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_4 FILLER_10_133 ();
 sg13g2_fill_2 FILLER_10_137 ();
 sg13g2_fill_1 FILLER_10_175 ();
 sg13g2_fill_2 FILLER_10_188 ();
 sg13g2_fill_2 FILLER_10_211 ();
 sg13g2_fill_1 FILLER_10_213 ();
 sg13g2_decap_8 FILLER_10_219 ();
 sg13g2_decap_4 FILLER_10_231 ();
 sg13g2_fill_1 FILLER_10_235 ();
 sg13g2_fill_1 FILLER_10_252 ();
 sg13g2_decap_4 FILLER_10_257 ();
 sg13g2_fill_1 FILLER_10_261 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_fill_1 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_fill_2 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_fill_1 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_fill_1 FILLER_10_338 ();
 sg13g2_fill_2 FILLER_10_344 ();
 sg13g2_fill_1 FILLER_10_346 ();
 sg13g2_fill_1 FILLER_10_357 ();
 sg13g2_fill_1 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_fill_2 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_156 ();
 sg13g2_decap_8 FILLER_11_162 ();
 sg13g2_fill_2 FILLER_11_169 ();
 sg13g2_fill_1 FILLER_11_171 ();
 sg13g2_fill_2 FILLER_11_186 ();
 sg13g2_fill_2 FILLER_11_200 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_fill_2 FILLER_11_213 ();
 sg13g2_decap_8 FILLER_11_236 ();
 sg13g2_decap_4 FILLER_11_243 ();
 sg13g2_fill_2 FILLER_11_309 ();
 sg13g2_fill_1 FILLER_11_311 ();
 sg13g2_decap_4 FILLER_11_318 ();
 sg13g2_fill_1 FILLER_11_337 ();
 sg13g2_fill_2 FILLER_11_348 ();
 sg13g2_fill_2 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_fill_2 FILLER_12_147 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_fill_1 FILLER_12_180 ();
 sg13g2_decap_4 FILLER_12_190 ();
 sg13g2_fill_1 FILLER_12_194 ();
 sg13g2_fill_1 FILLER_12_205 ();
 sg13g2_fill_2 FILLER_12_211 ();
 sg13g2_decap_4 FILLER_12_218 ();
 sg13g2_fill_2 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_fill_1 FILLER_12_257 ();
 sg13g2_fill_2 FILLER_12_262 ();
 sg13g2_decap_8 FILLER_12_269 ();
 sg13g2_decap_8 FILLER_12_276 ();
 sg13g2_fill_1 FILLER_12_283 ();
 sg13g2_fill_1 FILLER_12_338 ();
 sg13g2_fill_2 FILLER_12_357 ();
 sg13g2_fill_1 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_fill_2 FILLER_13_133 ();
 sg13g2_fill_2 FILLER_13_186 ();
 sg13g2_fill_1 FILLER_13_200 ();
 sg13g2_fill_2 FILLER_13_207 ();
 sg13g2_fill_1 FILLER_13_209 ();
 sg13g2_fill_1 FILLER_13_220 ();
 sg13g2_decap_8 FILLER_13_255 ();
 sg13g2_decap_8 FILLER_13_262 ();
 sg13g2_decap_8 FILLER_13_269 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_fill_2 FILLER_13_283 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_fill_1 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_fill_2 FILLER_13_333 ();
 sg13g2_decap_4 FILLER_13_341 ();
 sg13g2_fill_2 FILLER_13_351 ();
 sg13g2_fill_1 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_4 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_4 FILLER_14_133 ();
 sg13g2_fill_2 FILLER_14_137 ();
 sg13g2_fill_2 FILLER_14_176 ();
 sg13g2_fill_1 FILLER_14_178 ();
 sg13g2_fill_1 FILLER_14_193 ();
 sg13g2_decap_4 FILLER_14_213 ();
 sg13g2_fill_2 FILLER_14_217 ();
 sg13g2_fill_2 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_226 ();
 sg13g2_fill_2 FILLER_14_237 ();
 sg13g2_fill_1 FILLER_14_239 ();
 sg13g2_decap_4 FILLER_14_244 ();
 sg13g2_decap_4 FILLER_14_257 ();
 sg13g2_fill_2 FILLER_14_261 ();
 sg13g2_decap_4 FILLER_14_289 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_fill_1 FILLER_14_339 ();
 sg13g2_fill_1 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_358 ();
 sg13g2_fill_2 FILLER_14_365 ();
 sg13g2_decap_8 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_133 ();
 sg13g2_fill_1 FILLER_15_135 ();
 sg13g2_fill_1 FILLER_15_162 ();
 sg13g2_fill_2 FILLER_15_171 ();
 sg13g2_fill_1 FILLER_15_173 ();
 sg13g2_fill_2 FILLER_15_179 ();
 sg13g2_fill_1 FILLER_15_181 ();
 sg13g2_decap_4 FILLER_15_190 ();
 sg13g2_fill_1 FILLER_15_194 ();
 sg13g2_decap_8 FILLER_15_208 ();
 sg13g2_decap_4 FILLER_15_215 ();
 sg13g2_fill_1 FILLER_15_229 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_fill_1 FILLER_15_307 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_fill_2 FILLER_15_325 ();
 sg13g2_fill_2 FILLER_15_341 ();
 sg13g2_fill_1 FILLER_15_343 ();
 sg13g2_fill_2 FILLER_15_368 ();
 sg13g2_fill_1 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_fill_1 FILLER_16_164 ();
 sg13g2_decap_8 FILLER_16_172 ();
 sg13g2_decap_4 FILLER_16_179 ();
 sg13g2_fill_1 FILLER_16_183 ();
 sg13g2_fill_2 FILLER_16_198 ();
 sg13g2_fill_1 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_214 ();
 sg13g2_fill_1 FILLER_16_221 ();
 sg13g2_decap_4 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_240 ();
 sg13g2_fill_1 FILLER_16_242 ();
 sg13g2_fill_1 FILLER_16_264 ();
 sg13g2_decap_4 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_282 ();
 sg13g2_fill_2 FILLER_16_289 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_4 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_172 ();
 sg13g2_decap_8 FILLER_17_179 ();
 sg13g2_fill_1 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_200 ();
 sg13g2_decap_8 FILLER_17_271 ();
 sg13g2_fill_2 FILLER_17_300 ();
 sg13g2_fill_1 FILLER_17_302 ();
 sg13g2_fill_2 FILLER_17_308 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_fill_2 FILLER_17_320 ();
 sg13g2_fill_1 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_fill_1 FILLER_18_178 ();
 sg13g2_decap_4 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_188 ();
 sg13g2_fill_1 FILLER_18_218 ();
 sg13g2_fill_2 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_fill_2 FILLER_18_269 ();
 sg13g2_fill_1 FILLER_18_271 ();
 sg13g2_decap_4 FILLER_18_323 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_decap_4 FILLER_18_350 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_4 FILLER_18_366 ();
 sg13g2_fill_1 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_159 ();
 sg13g2_fill_2 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_170 ();
 sg13g2_fill_2 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_183 ();
 sg13g2_fill_2 FILLER_19_229 ();
 sg13g2_fill_1 FILLER_19_231 ();
 sg13g2_fill_1 FILLER_19_271 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_decap_8 FILLER_19_332 ();
 sg13g2_decap_8 FILLER_19_339 ();
 sg13g2_decap_4 FILLER_19_358 ();
 sg13g2_fill_2 FILLER_19_362 ();
 sg13g2_fill_2 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_4 FILLER_20_126 ();
 sg13g2_fill_1 FILLER_20_130 ();
 sg13g2_fill_2 FILLER_20_202 ();
 sg13g2_fill_1 FILLER_20_204 ();
 sg13g2_fill_2 FILLER_20_233 ();
 sg13g2_fill_1 FILLER_20_235 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_312 ();
 sg13g2_fill_2 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_fill_2 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_fill_2 FILLER_21_192 ();
 sg13g2_fill_1 FILLER_21_194 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_decap_8 FILLER_21_211 ();
 sg13g2_decap_4 FILLER_21_218 ();
 sg13g2_fill_2 FILLER_21_222 ();
 sg13g2_decap_4 FILLER_21_235 ();
 sg13g2_decap_4 FILLER_21_248 ();
 sg13g2_decap_4 FILLER_21_270 ();
 sg13g2_fill_2 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_282 ();
 sg13g2_fill_2 FILLER_21_291 ();
 sg13g2_fill_1 FILLER_21_359 ();
 sg13g2_decap_4 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_160 ();
 sg13g2_fill_2 FILLER_22_175 ();
 sg13g2_fill_2 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_191 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_fill_2 FILLER_22_213 ();
 sg13g2_fill_1 FILLER_22_215 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_decap_4 FILLER_22_242 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_258 ();
 sg13g2_decap_4 FILLER_22_265 ();
 sg13g2_fill_2 FILLER_22_269 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_4 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_295 ();
 sg13g2_decap_4 FILLER_22_314 ();
 sg13g2_fill_2 FILLER_22_318 ();
 sg13g2_fill_2 FILLER_22_325 ();
 sg13g2_fill_1 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_350 ();
 sg13g2_fill_1 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_4 FILLER_23_133 ();
 sg13g2_fill_2 FILLER_23_137 ();
 sg13g2_fill_2 FILLER_23_143 ();
 sg13g2_fill_1 FILLER_23_168 ();
 sg13g2_fill_2 FILLER_23_184 ();
 sg13g2_fill_1 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_218 ();
 sg13g2_decap_4 FILLER_23_250 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_294 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_fill_2 FILLER_23_337 ();
 sg13g2_fill_1 FILLER_23_339 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_decap_4 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_126 ();
 sg13g2_decap_4 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_170 ();
 sg13g2_fill_2 FILLER_24_182 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_decap_4 FILLER_24_196 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_decap_4 FILLER_24_220 ();
 sg13g2_fill_1 FILLER_24_274 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_decap_4 FILLER_24_304 ();
 sg13g2_fill_2 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_314 ();
 sg13g2_fill_2 FILLER_24_320 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_fill_1 FILLER_24_349 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_153 ();
 sg13g2_fill_1 FILLER_25_155 ();
 sg13g2_fill_2 FILLER_25_160 ();
 sg13g2_fill_2 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_284 ();
 sg13g2_decap_4 FILLER_25_317 ();
 sg13g2_fill_2 FILLER_25_336 ();
 sg13g2_fill_1 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_fill_2 FILLER_25_358 ();
 sg13g2_fill_1 FILLER_25_360 ();
 sg13g2_decap_4 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_4 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_142 ();
 sg13g2_fill_2 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_fill_2 FILLER_26_157 ();
 sg13g2_fill_1 FILLER_26_159 ();
 sg13g2_fill_2 FILLER_26_177 ();
 sg13g2_fill_1 FILLER_26_187 ();
 sg13g2_fill_2 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_198 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_225 ();
 sg13g2_fill_2 FILLER_26_240 ();
 sg13g2_decap_8 FILLER_26_282 ();
 sg13g2_decap_8 FILLER_26_302 ();
 sg13g2_fill_1 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_318 ();
 sg13g2_fill_2 FILLER_26_345 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_4 FILLER_27_133 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_180 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_195 ();
 sg13g2_decap_8 FILLER_27_202 ();
 sg13g2_decap_4 FILLER_27_209 ();
 sg13g2_fill_1 FILLER_27_213 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_fill_2 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_decap_8 FILLER_27_260 ();
 sg13g2_decap_8 FILLER_27_271 ();
 sg13g2_fill_1 FILLER_27_278 ();
 sg13g2_fill_1 FILLER_27_306 ();
 sg13g2_decap_4 FILLER_27_332 ();
 sg13g2_fill_1 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_4 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_194 ();
 sg13g2_fill_1 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_fill_2 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_228 ();
 sg13g2_fill_1 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_257 ();
 sg13g2_decap_8 FILLER_28_264 ();
 sg13g2_decap_4 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_decap_4 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_4 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_141 ();
 sg13g2_fill_2 FILLER_29_174 ();
 sg13g2_fill_1 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_236 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_290 ();
 sg13g2_fill_1 FILLER_29_292 ();
 sg13g2_fill_2 FILLER_29_302 ();
 sg13g2_fill_1 FILLER_29_304 ();
 sg13g2_decap_4 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_29_367 ();
 sg13g2_fill_1 FILLER_29_374 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_4 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_decap_4 FILLER_30_206 ();
 sg13g2_decap_8 FILLER_30_225 ();
 sg13g2_decap_8 FILLER_30_232 ();
 sg13g2_decap_8 FILLER_30_239 ();
 sg13g2_decap_4 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_decap_4 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_279 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_fill_2 FILLER_30_294 ();
 sg13g2_fill_1 FILLER_30_316 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_fill_1 FILLER_30_333 ();
 sg13g2_decap_4 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_fill_2 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_fill_1 FILLER_31_180 ();
 sg13g2_decap_4 FILLER_31_186 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_211 ();
 sg13g2_decap_8 FILLER_31_244 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_decap_8 FILLER_31_256 ();
 sg13g2_decap_8 FILLER_31_278 ();
 sg13g2_decap_8 FILLER_31_285 ();
 sg13g2_fill_2 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_327 ();
 sg13g2_decap_4 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_338 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_fill_2 FILLER_32_194 ();
 sg13g2_fill_1 FILLER_32_196 ();
 sg13g2_decap_4 FILLER_32_209 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_287 ();
 sg13g2_decap_4 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_349 ();
 sg13g2_decap_8 FILLER_32_356 ();
 sg13g2_decap_8 FILLER_32_363 ();
 sg13g2_fill_2 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_152 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_170 ();
 sg13g2_decap_8 FILLER_33_183 ();
 sg13g2_decap_8 FILLER_33_190 ();
 sg13g2_decap_4 FILLER_33_197 ();
 sg13g2_fill_2 FILLER_33_201 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_decap_4 FILLER_33_248 ();
 sg13g2_decap_4 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_390 ();
 sg13g2_decap_8 FILLER_33_397 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_4 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_142 ();
 sg13g2_decap_8 FILLER_34_152 ();
 sg13g2_fill_1 FILLER_34_159 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_decap_8 FILLER_34_219 ();
 sg13g2_fill_2 FILLER_34_226 ();
 sg13g2_fill_1 FILLER_34_228 ();
 sg13g2_decap_8 FILLER_34_233 ();
 sg13g2_decap_8 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_267 ();
 sg13g2_fill_1 FILLER_34_269 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_decap_4 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_fill_2 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_146 ();
 sg13g2_decap_8 FILLER_35_152 ();
 sg13g2_decap_8 FILLER_35_159 ();
 sg13g2_decap_8 FILLER_35_169 ();
 sg13g2_decap_8 FILLER_35_176 ();
 sg13g2_decap_4 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_194 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_226 ();
 sg13g2_fill_2 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_268 ();
 sg13g2_fill_2 FILLER_35_273 ();
 sg13g2_decap_4 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_311 ();
 sg13g2_fill_1 FILLER_35_313 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_fill_2 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_335 ();
 sg13g2_fill_2 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_165 ();
 sg13g2_decap_4 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_268 ();
 sg13g2_fill_2 FILLER_36_304 ();
 sg13g2_fill_1 FILLER_36_306 ();
 sg13g2_fill_2 FILLER_36_329 ();
 sg13g2_fill_2 FILLER_36_339 ();
 sg13g2_fill_1 FILLER_36_341 ();
 sg13g2_fill_2 FILLER_36_356 ();
 sg13g2_fill_2 FILLER_36_384 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_132 ();
 sg13g2_fill_1 FILLER_37_138 ();
 sg13g2_decap_4 FILLER_37_227 ();
 sg13g2_fill_2 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_241 ();
 sg13g2_decap_4 FILLER_37_246 ();
 sg13g2_decap_4 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_259 ();
 sg13g2_fill_2 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_fill_2 FILLER_37_343 ();
 sg13g2_fill_1 FILLER_37_361 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_4 FILLER_38_105 ();
 sg13g2_fill_2 FILLER_38_109 ();
 sg13g2_fill_2 FILLER_38_147 ();
 sg13g2_fill_1 FILLER_38_166 ();
 sg13g2_fill_2 FILLER_38_193 ();
 sg13g2_fill_2 FILLER_38_219 ();
 sg13g2_decap_4 FILLER_38_243 ();
 sg13g2_fill_2 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_decap_4 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_fill_2 FILLER_38_354 ();
 sg13g2_fill_1 FILLER_38_356 ();
 sg13g2_fill_2 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_fill_2 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_104 ();
 sg13g2_fill_2 FILLER_39_111 ();
 sg13g2_fill_2 FILLER_39_120 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_fill_2 FILLER_39_135 ();
 sg13g2_fill_2 FILLER_39_146 ();
 sg13g2_fill_1 FILLER_39_148 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_fill_1 FILLER_39_175 ();
 sg13g2_decap_4 FILLER_39_231 ();
 sg13g2_fill_2 FILLER_39_235 ();
 sg13g2_fill_2 FILLER_39_242 ();
 sg13g2_fill_1 FILLER_39_244 ();
 sg13g2_fill_2 FILLER_39_276 ();
 sg13g2_fill_1 FILLER_39_278 ();
 sg13g2_fill_2 FILLER_39_283 ();
 sg13g2_fill_1 FILLER_39_285 ();
 sg13g2_fill_2 FILLER_39_291 ();
 sg13g2_decap_8 FILLER_39_313 ();
 sg13g2_decap_8 FILLER_39_320 ();
 sg13g2_fill_1 FILLER_39_327 ();
 sg13g2_fill_2 FILLER_39_337 ();
 sg13g2_decap_4 FILLER_39_344 ();
 sg13g2_fill_1 FILLER_39_348 ();
 sg13g2_decap_8 FILLER_39_396 ();
 sg13g2_decap_4 FILLER_39_403 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_4 FILLER_40_84 ();
 sg13g2_fill_1 FILLER_40_88 ();
 sg13g2_decap_4 FILLER_40_115 ();
 sg13g2_decap_4 FILLER_40_126 ();
 sg13g2_fill_2 FILLER_40_141 ();
 sg13g2_fill_1 FILLER_40_143 ();
 sg13g2_fill_1 FILLER_40_158 ();
 sg13g2_decap_8 FILLER_40_163 ();
 sg13g2_fill_2 FILLER_40_170 ();
 sg13g2_decap_4 FILLER_40_197 ();
 sg13g2_fill_2 FILLER_40_201 ();
 sg13g2_fill_2 FILLER_40_211 ();
 sg13g2_fill_1 FILLER_40_219 ();
 sg13g2_fill_1 FILLER_40_241 ();
 sg13g2_fill_1 FILLER_40_255 ();
 sg13g2_decap_8 FILLER_40_260 ();
 sg13g2_fill_1 FILLER_40_267 ();
 sg13g2_fill_1 FILLER_40_275 ();
 sg13g2_fill_2 FILLER_40_286 ();
 sg13g2_decap_8 FILLER_40_316 ();
 sg13g2_decap_4 FILLER_40_323 ();
 sg13g2_decap_8 FILLER_40_332 ();
 sg13g2_decap_4 FILLER_40_339 ();
 sg13g2_fill_2 FILLER_40_343 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_fill_1 FILLER_41_91 ();
 sg13g2_fill_1 FILLER_41_109 ();
 sg13g2_decap_8 FILLER_41_115 ();
 sg13g2_fill_1 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_155 ();
 sg13g2_fill_2 FILLER_41_162 ();
 sg13g2_fill_2 FILLER_41_197 ();
 sg13g2_fill_2 FILLER_41_209 ();
 sg13g2_fill_1 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_225 ();
 sg13g2_decap_8 FILLER_41_253 ();
 sg13g2_fill_1 FILLER_41_260 ();
 sg13g2_fill_1 FILLER_41_267 ();
 sg13g2_decap_4 FILLER_41_289 ();
 sg13g2_fill_1 FILLER_41_293 ();
 sg13g2_fill_2 FILLER_41_363 ();
 sg13g2_fill_1 FILLER_41_365 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_fill_2 FILLER_42_84 ();
 sg13g2_fill_2 FILLER_42_104 ();
 sg13g2_fill_1 FILLER_42_106 ();
 sg13g2_fill_2 FILLER_42_124 ();
 sg13g2_fill_2 FILLER_42_155 ();
 sg13g2_fill_1 FILLER_42_157 ();
 sg13g2_decap_4 FILLER_42_163 ();
 sg13g2_fill_2 FILLER_42_193 ();
 sg13g2_fill_1 FILLER_42_195 ();
 sg13g2_decap_4 FILLER_42_211 ();
 sg13g2_fill_1 FILLER_42_227 ();
 sg13g2_fill_2 FILLER_42_237 ();
 sg13g2_fill_1 FILLER_42_239 ();
 sg13g2_fill_2 FILLER_42_246 ();
 sg13g2_fill_1 FILLER_42_248 ();
 sg13g2_fill_2 FILLER_42_259 ();
 sg13g2_fill_2 FILLER_42_287 ();
 sg13g2_fill_2 FILLER_42_362 ();
 sg13g2_fill_2 FILLER_42_385 ();
 sg13g2_fill_1 FILLER_42_387 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_fill_1 FILLER_43_84 ();
 sg13g2_fill_2 FILLER_43_138 ();
 sg13g2_fill_1 FILLER_43_140 ();
 sg13g2_fill_2 FILLER_43_151 ();
 sg13g2_fill_1 FILLER_43_153 ();
 sg13g2_fill_2 FILLER_43_159 ();
 sg13g2_fill_1 FILLER_43_161 ();
 sg13g2_fill_2 FILLER_43_173 ();
 sg13g2_decap_4 FILLER_43_183 ();
 sg13g2_fill_2 FILLER_43_187 ();
 sg13g2_fill_1 FILLER_43_210 ();
 sg13g2_decap_4 FILLER_43_215 ();
 sg13g2_fill_2 FILLER_43_219 ();
 sg13g2_fill_1 FILLER_43_234 ();
 sg13g2_decap_8 FILLER_43_244 ();
 sg13g2_decap_8 FILLER_43_251 ();
 sg13g2_fill_2 FILLER_43_258 ();
 sg13g2_decap_4 FILLER_43_265 ();
 sg13g2_fill_2 FILLER_43_269 ();
 sg13g2_fill_2 FILLER_43_305 ();
 sg13g2_fill_1 FILLER_43_307 ();
 sg13g2_decap_4 FILLER_43_317 ();
 sg13g2_decap_4 FILLER_43_325 ();
 sg13g2_fill_2 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_4 FILLER_43_385 ();
 sg13g2_fill_2 FILLER_43_389 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_fill_2 FILLER_44_77 ();
 sg13g2_fill_1 FILLER_44_79 ();
 sg13g2_fill_2 FILLER_44_106 ();
 sg13g2_fill_2 FILLER_44_124 ();
 sg13g2_fill_2 FILLER_44_131 ();
 sg13g2_fill_1 FILLER_44_133 ();
 sg13g2_fill_2 FILLER_44_144 ();
 sg13g2_decap_8 FILLER_44_163 ();
 sg13g2_decap_8 FILLER_44_170 ();
 sg13g2_decap_4 FILLER_44_177 ();
 sg13g2_fill_2 FILLER_44_181 ();
 sg13g2_decap_4 FILLER_44_188 ();
 sg13g2_fill_1 FILLER_44_192 ();
 sg13g2_fill_1 FILLER_44_201 ();
 sg13g2_fill_1 FILLER_44_226 ();
 sg13g2_decap_8 FILLER_44_239 ();
 sg13g2_fill_2 FILLER_44_246 ();
 sg13g2_fill_1 FILLER_44_248 ();
 sg13g2_decap_8 FILLER_44_264 ();
 sg13g2_decap_8 FILLER_44_271 ();
 sg13g2_decap_8 FILLER_44_278 ();
 sg13g2_fill_2 FILLER_44_285 ();
 sg13g2_fill_1 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_293 ();
 sg13g2_decap_4 FILLER_44_300 ();
 sg13g2_fill_2 FILLER_44_304 ();
 sg13g2_decap_8 FILLER_44_316 ();
 sg13g2_fill_1 FILLER_44_323 ();
 sg13g2_decap_8 FILLER_44_341 ();
 sg13g2_decap_8 FILLER_44_348 ();
 sg13g2_decap_8 FILLER_44_387 ();
 sg13g2_decap_8 FILLER_44_394 ();
 sg13g2_decap_8 FILLER_44_401 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_118 ();
 sg13g2_fill_1 FILLER_45_125 ();
 sg13g2_fill_1 FILLER_45_157 ();
 sg13g2_decap_8 FILLER_45_171 ();
 sg13g2_fill_1 FILLER_45_178 ();
 sg13g2_fill_2 FILLER_45_193 ();
 sg13g2_fill_1 FILLER_45_195 ();
 sg13g2_fill_1 FILLER_45_224 ();
 sg13g2_fill_2 FILLER_45_236 ();
 sg13g2_decap_8 FILLER_45_269 ();
 sg13g2_decap_8 FILLER_45_276 ();
 sg13g2_fill_2 FILLER_45_283 ();
 sg13g2_decap_8 FILLER_45_311 ();
 sg13g2_fill_1 FILLER_45_342 ();
 sg13g2_decap_4 FILLER_45_355 ();
 sg13g2_fill_2 FILLER_45_359 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_fill_2 FILLER_46_98 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_decap_4 FILLER_46_104 ();
 sg13g2_fill_2 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_114 ();
 sg13g2_fill_1 FILLER_46_140 ();
 sg13g2_fill_2 FILLER_46_170 ();
 sg13g2_fill_1 FILLER_46_172 ();
 sg13g2_decap_4 FILLER_46_204 ();
 sg13g2_fill_1 FILLER_46_246 ();
 sg13g2_fill_2 FILLER_46_251 ();
 sg13g2_decap_4 FILLER_46_279 ();
 sg13g2_fill_2 FILLER_46_283 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_4 FILLER_47_84 ();
 sg13g2_fill_2 FILLER_47_88 ();
 sg13g2_fill_1 FILLER_47_142 ();
 sg13g2_fill_2 FILLER_47_164 ();
 sg13g2_fill_1 FILLER_47_179 ();
 sg13g2_fill_1 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_196 ();
 sg13g2_decap_4 FILLER_47_213 ();
 sg13g2_fill_2 FILLER_47_222 ();
 sg13g2_fill_1 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_fill_2 FILLER_47_245 ();
 sg13g2_fill_2 FILLER_47_255 ();
 sg13g2_fill_1 FILLER_47_257 ();
 sg13g2_fill_2 FILLER_47_269 ();
 sg13g2_fill_1 FILLER_47_279 ();
 sg13g2_decap_4 FILLER_47_288 ();
 sg13g2_fill_2 FILLER_47_300 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_fill_1 FILLER_47_315 ();
 sg13g2_fill_2 FILLER_47_331 ();
 sg13g2_fill_1 FILLER_47_362 ();
 sg13g2_fill_2 FILLER_47_372 ();
 sg13g2_decap_8 FILLER_47_389 ();
 sg13g2_decap_8 FILLER_47_396 ();
 sg13g2_decap_4 FILLER_47_403 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_fill_1 FILLER_48_127 ();
 sg13g2_fill_2 FILLER_48_153 ();
 sg13g2_decap_8 FILLER_48_176 ();
 sg13g2_decap_8 FILLER_48_183 ();
 sg13g2_decap_4 FILLER_48_190 ();
 sg13g2_fill_1 FILLER_48_194 ();
 sg13g2_decap_8 FILLER_48_229 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_decap_8 FILLER_48_297 ();
 sg13g2_decap_8 FILLER_48_312 ();
 sg13g2_decap_8 FILLER_48_319 ();
 sg13g2_fill_1 FILLER_48_329 ();
 sg13g2_fill_2 FILLER_48_350 ();
 sg13g2_fill_1 FILLER_48_352 ();
 sg13g2_fill_2 FILLER_48_376 ();
 sg13g2_fill_1 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_4 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_139 ();
 sg13g2_decap_8 FILLER_49_151 ();
 sg13g2_fill_2 FILLER_49_158 ();
 sg13g2_decap_8 FILLER_49_165 ();
 sg13g2_fill_1 FILLER_49_172 ();
 sg13g2_fill_1 FILLER_49_208 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_fill_2 FILLER_49_271 ();
 sg13g2_fill_1 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_290 ();
 sg13g2_decap_8 FILLER_49_297 ();
 sg13g2_decap_8 FILLER_49_312 ();
 sg13g2_fill_1 FILLER_49_319 ();
 sg13g2_decap_8 FILLER_49_328 ();
 sg13g2_decap_8 FILLER_49_335 ();
 sg13g2_decap_8 FILLER_49_342 ();
 sg13g2_fill_1 FILLER_49_349 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_4 FILLER_50_77 ();
 sg13g2_fill_1 FILLER_50_81 ();
 sg13g2_fill_1 FILLER_50_113 ();
 sg13g2_fill_1 FILLER_50_122 ();
 sg13g2_decap_8 FILLER_50_128 ();
 sg13g2_decap_4 FILLER_50_135 ();
 sg13g2_fill_2 FILLER_50_143 ();
 sg13g2_fill_1 FILLER_50_145 ();
 sg13g2_fill_1 FILLER_50_151 ();
 sg13g2_decap_4 FILLER_50_159 ();
 sg13g2_decap_8 FILLER_50_173 ();
 sg13g2_fill_1 FILLER_50_217 ();
 sg13g2_fill_1 FILLER_50_284 ();
 sg13g2_fill_1 FILLER_50_295 ();
 sg13g2_fill_2 FILLER_50_300 ();
 sg13g2_fill_2 FILLER_50_323 ();
 sg13g2_decap_8 FILLER_50_338 ();
 sg13g2_decap_8 FILLER_50_345 ();
 sg13g2_fill_2 FILLER_50_352 ();
 sg13g2_fill_1 FILLER_50_354 ();
 sg13g2_decap_8 FILLER_50_393 ();
 sg13g2_decap_8 FILLER_50_400 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_4 FILLER_51_84 ();
 sg13g2_fill_1 FILLER_51_113 ();
 sg13g2_decap_4 FILLER_51_127 ();
 sg13g2_decap_4 FILLER_51_173 ();
 sg13g2_fill_2 FILLER_51_177 ();
 sg13g2_fill_2 FILLER_51_204 ();
 sg13g2_fill_2 FILLER_51_216 ();
 sg13g2_fill_1 FILLER_51_218 ();
 sg13g2_fill_2 FILLER_51_231 ();
 sg13g2_decap_8 FILLER_51_251 ();
 sg13g2_decap_4 FILLER_51_258 ();
 sg13g2_fill_1 FILLER_51_262 ();
 sg13g2_decap_4 FILLER_51_273 ();
 sg13g2_fill_2 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_284 ();
 sg13g2_decap_8 FILLER_51_311 ();
 sg13g2_decap_4 FILLER_51_326 ();
 sg13g2_decap_4 FILLER_51_343 ();
 sg13g2_decap_8 FILLER_51_352 ();
 sg13g2_decap_4 FILLER_51_359 ();
 sg13g2_fill_1 FILLER_51_363 ();
 sg13g2_decap_4 FILLER_51_369 ();
 sg13g2_fill_1 FILLER_51_373 ();
 sg13g2_decap_4 FILLER_51_404 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_fill_1 FILLER_52_103 ();
 sg13g2_decap_4 FILLER_52_127 ();
 sg13g2_fill_2 FILLER_52_138 ();
 sg13g2_fill_1 FILLER_52_140 ();
 sg13g2_fill_2 FILLER_52_147 ();
 sg13g2_fill_1 FILLER_52_149 ();
 sg13g2_decap_8 FILLER_52_172 ();
 sg13g2_fill_2 FILLER_52_179 ();
 sg13g2_decap_4 FILLER_52_212 ();
 sg13g2_fill_2 FILLER_52_216 ();
 sg13g2_fill_1 FILLER_52_234 ();
 sg13g2_decap_8 FILLER_52_239 ();
 sg13g2_decap_4 FILLER_52_246 ();
 sg13g2_fill_2 FILLER_52_250 ();
 sg13g2_fill_2 FILLER_52_258 ();
 sg13g2_fill_1 FILLER_52_273 ();
 sg13g2_decap_4 FILLER_52_300 ();
 sg13g2_fill_1 FILLER_52_304 ();
 sg13g2_decap_4 FILLER_52_318 ();
 sg13g2_fill_1 FILLER_52_330 ();
 sg13g2_fill_1 FILLER_52_336 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_fill_2 FILLER_53_84 ();
 sg13g2_fill_1 FILLER_53_86 ();
 sg13g2_fill_1 FILLER_53_95 ();
 sg13g2_fill_2 FILLER_53_105 ();
 sg13g2_fill_2 FILLER_53_127 ();
 sg13g2_fill_1 FILLER_53_165 ();
 sg13g2_decap_4 FILLER_53_176 ();
 sg13g2_decap_8 FILLER_53_185 ();
 sg13g2_decap_4 FILLER_53_196 ();
 sg13g2_fill_2 FILLER_53_200 ();
 sg13g2_decap_8 FILLER_53_242 ();
 sg13g2_decap_4 FILLER_53_249 ();
 sg13g2_fill_1 FILLER_53_263 ();
 sg13g2_fill_1 FILLER_53_290 ();
 sg13g2_decap_8 FILLER_53_300 ();
 sg13g2_decap_8 FILLER_53_307 ();
 sg13g2_decap_8 FILLER_53_314 ();
 sg13g2_decap_4 FILLER_53_321 ();
 sg13g2_fill_2 FILLER_53_325 ();
 sg13g2_decap_4 FILLER_53_348 ();
 sg13g2_fill_1 FILLER_53_365 ();
 sg13g2_fill_2 FILLER_53_392 ();
 sg13g2_decap_8 FILLER_53_398 ();
 sg13g2_decap_4 FILLER_53_405 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_fill_2 FILLER_54_81 ();
 sg13g2_fill_1 FILLER_54_152 ();
 sg13g2_decap_4 FILLER_54_204 ();
 sg13g2_fill_1 FILLER_54_234 ();
 sg13g2_fill_1 FILLER_54_243 ();
 sg13g2_decap_4 FILLER_54_258 ();
 sg13g2_decap_4 FILLER_54_295 ();
 sg13g2_fill_1 FILLER_54_317 ();
 sg13g2_decap_4 FILLER_54_323 ();
 sg13g2_decap_8 FILLER_54_332 ();
 sg13g2_fill_1 FILLER_54_357 ();
 sg13g2_fill_2 FILLER_54_393 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_fill_2 FILLER_55_63 ();
 sg13g2_fill_1 FILLER_55_65 ();
 sg13g2_fill_1 FILLER_55_132 ();
 sg13g2_fill_2 FILLER_55_137 ();
 sg13g2_fill_1 FILLER_55_139 ();
 sg13g2_fill_1 FILLER_55_152 ();
 sg13g2_fill_1 FILLER_55_171 ();
 sg13g2_decap_8 FILLER_55_176 ();
 sg13g2_decap_4 FILLER_55_193 ();
 sg13g2_fill_2 FILLER_55_197 ();
 sg13g2_fill_2 FILLER_55_234 ();
 sg13g2_fill_2 FILLER_55_244 ();
 sg13g2_fill_1 FILLER_55_246 ();
 sg13g2_decap_4 FILLER_55_256 ();
 sg13g2_fill_1 FILLER_55_260 ();
 sg13g2_decap_4 FILLER_55_338 ();
 sg13g2_fill_2 FILLER_55_347 ();
 sg13g2_fill_1 FILLER_55_349 ();
 sg13g2_decap_4 FILLER_55_371 ();
 sg13g2_decap_4 FILLER_55_387 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_4 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_60 ();
 sg13g2_decap_4 FILLER_56_128 ();
 sg13g2_decap_8 FILLER_56_136 ();
 sg13g2_decap_4 FILLER_56_143 ();
 sg13g2_fill_1 FILLER_56_147 ();
 sg13g2_fill_1 FILLER_56_153 ();
 sg13g2_decap_8 FILLER_56_172 ();
 sg13g2_decap_4 FILLER_56_179 ();
 sg13g2_fill_2 FILLER_56_183 ();
 sg13g2_decap_8 FILLER_56_189 ();
 sg13g2_decap_8 FILLER_56_196 ();
 sg13g2_decap_4 FILLER_56_203 ();
 sg13g2_fill_2 FILLER_56_207 ();
 sg13g2_fill_2 FILLER_56_213 ();
 sg13g2_fill_1 FILLER_56_215 ();
 sg13g2_fill_1 FILLER_56_222 ();
 sg13g2_decap_4 FILLER_56_238 ();
 sg13g2_fill_2 FILLER_56_250 ();
 sg13g2_fill_1 FILLER_56_258 ();
 sg13g2_fill_1 FILLER_56_284 ();
 sg13g2_fill_1 FILLER_56_290 ();
 sg13g2_fill_2 FILLER_56_335 ();
 sg13g2_fill_1 FILLER_56_337 ();
 sg13g2_decap_8 FILLER_56_346 ();
 sg13g2_decap_4 FILLER_56_353 ();
 sg13g2_fill_2 FILLER_56_357 ();
 sg13g2_fill_1 FILLER_56_364 ();
 sg13g2_fill_1 FILLER_56_369 ();
 sg13g2_fill_1 FILLER_56_373 ();
 sg13g2_decap_8 FILLER_56_379 ();
 sg13g2_fill_2 FILLER_56_386 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_4 FILLER_57_49 ();
 sg13g2_fill_2 FILLER_57_53 ();
 sg13g2_fill_1 FILLER_57_83 ();
 sg13g2_fill_2 FILLER_57_101 ();
 sg13g2_fill_1 FILLER_57_116 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_fill_2 FILLER_57_165 ();
 sg13g2_fill_2 FILLER_57_177 ();
 sg13g2_fill_1 FILLER_57_179 ();
 sg13g2_decap_8 FILLER_57_200 ();
 sg13g2_decap_4 FILLER_57_207 ();
 sg13g2_fill_1 FILLER_57_211 ();
 sg13g2_fill_1 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_258 ();
 sg13g2_decap_8 FILLER_57_265 ();
 sg13g2_fill_2 FILLER_57_289 ();
 sg13g2_fill_1 FILLER_57_291 ();
 sg13g2_fill_1 FILLER_57_321 ();
 sg13g2_fill_2 FILLER_57_346 ();
 sg13g2_fill_1 FILLER_57_348 ();
 sg13g2_fill_1 FILLER_57_380 ();
 sg13g2_decap_4 FILLER_57_389 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_fill_2 FILLER_58_49 ();
 sg13g2_fill_1 FILLER_58_138 ();
 sg13g2_fill_1 FILLER_58_144 ();
 sg13g2_fill_1 FILLER_58_222 ();
 sg13g2_fill_2 FILLER_58_249 ();
 sg13g2_decap_4 FILLER_58_277 ();
 sg13g2_decap_8 FILLER_58_286 ();
 sg13g2_decap_4 FILLER_58_293 ();
 sg13g2_fill_2 FILLER_58_297 ();
 sg13g2_decap_4 FILLER_58_317 ();
 sg13g2_fill_2 FILLER_58_360 ();
 sg13g2_fill_2 FILLER_58_380 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_4 FILLER_59_35 ();
 sg13g2_fill_1 FILLER_59_69 ();
 sg13g2_fill_2 FILLER_59_88 ();
 sg13g2_fill_1 FILLER_59_90 ();
 sg13g2_fill_2 FILLER_59_148 ();
 sg13g2_fill_1 FILLER_59_171 ();
 sg13g2_fill_2 FILLER_59_187 ();
 sg13g2_fill_1 FILLER_59_201 ();
 sg13g2_fill_1 FILLER_59_216 ();
 sg13g2_fill_2 FILLER_59_233 ();
 sg13g2_fill_1 FILLER_59_235 ();
 sg13g2_decap_8 FILLER_59_275 ();
 sg13g2_decap_8 FILLER_59_282 ();
 sg13g2_fill_2 FILLER_59_289 ();
 sg13g2_decap_4 FILLER_59_295 ();
 sg13g2_fill_1 FILLER_59_299 ();
 sg13g2_decap_4 FILLER_59_309 ();
 sg13g2_fill_1 FILLER_59_313 ();
 sg13g2_fill_2 FILLER_59_317 ();
 sg13g2_fill_1 FILLER_59_319 ();
 sg13g2_fill_2 FILLER_59_325 ();
 sg13g2_fill_1 FILLER_59_355 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_fill_1 FILLER_60_42 ();
 sg13g2_fill_2 FILLER_60_125 ();
 sg13g2_fill_2 FILLER_60_146 ();
 sg13g2_fill_1 FILLER_60_148 ();
 sg13g2_decap_8 FILLER_60_153 ();
 sg13g2_fill_1 FILLER_60_160 ();
 sg13g2_decap_4 FILLER_60_165 ();
 sg13g2_fill_1 FILLER_60_169 ();
 sg13g2_decap_8 FILLER_60_179 ();
 sg13g2_decap_8 FILLER_60_186 ();
 sg13g2_decap_8 FILLER_60_197 ();
 sg13g2_decap_8 FILLER_60_204 ();
 sg13g2_decap_8 FILLER_60_211 ();
 sg13g2_fill_2 FILLER_60_218 ();
 sg13g2_fill_1 FILLER_60_220 ();
 sg13g2_fill_2 FILLER_60_231 ();
 sg13g2_fill_1 FILLER_60_233 ();
 sg13g2_fill_2 FILLER_60_238 ();
 sg13g2_fill_1 FILLER_60_240 ();
 sg13g2_fill_1 FILLER_60_255 ();
 sg13g2_fill_2 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_370 ();
 sg13g2_fill_1 FILLER_60_377 ();
 sg13g2_fill_2 FILLER_60_390 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_100 ();
 sg13g2_decap_4 FILLER_61_107 ();
 sg13g2_fill_2 FILLER_61_120 ();
 sg13g2_fill_2 FILLER_61_154 ();
 sg13g2_fill_1 FILLER_61_156 ();
 sg13g2_fill_2 FILLER_61_185 ();
 sg13g2_decap_8 FILLER_61_192 ();
 sg13g2_decap_8 FILLER_61_199 ();
 sg13g2_decap_8 FILLER_61_206 ();
 sg13g2_decap_8 FILLER_61_213 ();
 sg13g2_decap_4 FILLER_61_220 ();
 sg13g2_decap_8 FILLER_61_228 ();
 sg13g2_decap_8 FILLER_61_235 ();
 sg13g2_fill_2 FILLER_61_242 ();
 sg13g2_decap_8 FILLER_61_248 ();
 sg13g2_decap_8 FILLER_61_260 ();
 sg13g2_fill_1 FILLER_61_317 ();
 sg13g2_decap_4 FILLER_61_344 ();
 sg13g2_fill_1 FILLER_61_348 ();
 sg13g2_fill_2 FILLER_61_354 ();
 sg13g2_fill_1 FILLER_61_356 ();
 sg13g2_decap_8 FILLER_61_365 ();
 sg13g2_decap_8 FILLER_61_372 ();
 sg13g2_decap_4 FILLER_61_379 ();
 sg13g2_fill_1 FILLER_61_383 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_4 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_83 ();
 sg13g2_fill_2 FILLER_62_99 ();
 sg13g2_fill_1 FILLER_62_101 ();
 sg13g2_fill_2 FILLER_62_119 ();
 sg13g2_fill_2 FILLER_62_172 ();
 sg13g2_fill_2 FILLER_62_192 ();
 sg13g2_decap_4 FILLER_62_200 ();
 sg13g2_fill_2 FILLER_62_260 ();
 sg13g2_fill_2 FILLER_62_267 ();
 sg13g2_fill_1 FILLER_62_281 ();
 sg13g2_fill_2 FILLER_62_287 ();
 sg13g2_fill_1 FILLER_62_309 ();
 sg13g2_decap_4 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_401 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_4 FILLER_63_35 ();
 sg13g2_fill_1 FILLER_63_39 ();
 sg13g2_decap_4 FILLER_63_92 ();
 sg13g2_decap_4 FILLER_63_170 ();
 sg13g2_fill_1 FILLER_63_221 ();
 sg13g2_fill_2 FILLER_63_253 ();
 sg13g2_decap_4 FILLER_63_286 ();
 sg13g2_fill_2 FILLER_63_290 ();
 sg13g2_decap_8 FILLER_63_296 ();
 sg13g2_decap_4 FILLER_63_303 ();
 sg13g2_fill_2 FILLER_63_321 ();
 sg13g2_fill_1 FILLER_63_323 ();
 sg13g2_decap_4 FILLER_63_334 ();
 sg13g2_fill_2 FILLER_63_338 ();
 sg13g2_decap_8 FILLER_63_363 ();
 sg13g2_decap_4 FILLER_63_389 ();
 sg13g2_decap_4 FILLER_63_405 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_fill_1 FILLER_64_35 ();
 sg13g2_fill_1 FILLER_64_71 ();
 sg13g2_fill_1 FILLER_64_142 ();
 sg13g2_fill_2 FILLER_64_166 ();
 sg13g2_fill_1 FILLER_64_173 ();
 sg13g2_decap_4 FILLER_64_202 ();
 sg13g2_fill_1 FILLER_64_206 ();
 sg13g2_fill_2 FILLER_64_223 ();
 sg13g2_decap_8 FILLER_64_251 ();
 sg13g2_fill_2 FILLER_64_278 ();
 sg13g2_fill_1 FILLER_64_280 ();
 sg13g2_decap_4 FILLER_64_290 ();
 sg13g2_fill_2 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_303 ();
 sg13g2_decap_8 FILLER_64_310 ();
 sg13g2_decap_8 FILLER_64_317 ();
 sg13g2_decap_8 FILLER_64_324 ();
 sg13g2_fill_1 FILLER_64_331 ();
 sg13g2_decap_8 FILLER_64_353 ();
 sg13g2_fill_2 FILLER_64_377 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_fill_2 FILLER_65_35 ();
 sg13g2_fill_1 FILLER_65_81 ();
 sg13g2_fill_1 FILLER_65_134 ();
 sg13g2_fill_2 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_143 ();
 sg13g2_fill_2 FILLER_65_149 ();
 sg13g2_decap_8 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_fill_2 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_219 ();
 sg13g2_decap_4 FILLER_65_229 ();
 sg13g2_decap_8 FILLER_65_241 ();
 sg13g2_fill_2 FILLER_65_248 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_fill_2 FILLER_66_35 ();
 sg13g2_fill_1 FILLER_66_63 ();
 sg13g2_fill_2 FILLER_66_73 ();
 sg13g2_fill_1 FILLER_66_95 ();
 sg13g2_fill_1 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_135 ();
 sg13g2_fill_1 FILLER_66_142 ();
 sg13g2_decap_4 FILLER_66_148 ();
 sg13g2_decap_8 FILLER_66_159 ();
 sg13g2_decap_8 FILLER_66_184 ();
 sg13g2_decap_8 FILLER_66_191 ();
 sg13g2_decap_8 FILLER_66_198 ();
 sg13g2_fill_1 FILLER_66_205 ();
 sg13g2_fill_2 FILLER_66_211 ();
 sg13g2_fill_1 FILLER_66_213 ();
 sg13g2_decap_4 FILLER_66_219 ();
 sg13g2_decap_4 FILLER_66_230 ();
 sg13g2_fill_2 FILLER_66_234 ();
 sg13g2_fill_2 FILLER_66_262 ();
 sg13g2_fill_1 FILLER_66_264 ();
 sg13g2_fill_2 FILLER_66_293 ();
 sg13g2_fill_2 FILLER_66_305 ();
 sg13g2_fill_2 FILLER_66_333 ();
 sg13g2_decap_4 FILLER_66_378 ();
 sg13g2_fill_1 FILLER_66_382 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_4 FILLER_67_42 ();
 sg13g2_fill_1 FILLER_67_46 ();
 sg13g2_fill_2 FILLER_67_89 ();
 sg13g2_fill_2 FILLER_67_100 ();
 sg13g2_fill_1 FILLER_67_102 ();
 sg13g2_fill_2 FILLER_67_112 ();
 sg13g2_fill_1 FILLER_67_114 ();
 sg13g2_decap_8 FILLER_67_137 ();
 sg13g2_fill_2 FILLER_67_144 ();
 sg13g2_fill_1 FILLER_67_146 ();
 sg13g2_fill_1 FILLER_67_208 ();
 sg13g2_decap_8 FILLER_67_240 ();
 sg13g2_decap_8 FILLER_67_251 ();
 sg13g2_fill_1 FILLER_67_258 ();
 sg13g2_fill_1 FILLER_67_299 ();
 sg13g2_fill_1 FILLER_67_304 ();
 sg13g2_fill_1 FILLER_67_325 ();
 sg13g2_fill_1 FILLER_67_331 ();
 sg13g2_fill_2 FILLER_67_342 ();
 sg13g2_fill_2 FILLER_67_348 ();
 sg13g2_fill_2 FILLER_67_356 ();
 sg13g2_fill_2 FILLER_67_370 ();
 sg13g2_decap_8 FILLER_67_398 ();
 sg13g2_decap_4 FILLER_67_405 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_fill_2 FILLER_68_42 ();
 sg13g2_fill_1 FILLER_68_70 ();
 sg13g2_fill_1 FILLER_68_86 ();
 sg13g2_decap_4 FILLER_68_139 ();
 sg13g2_fill_1 FILLER_68_143 ();
 sg13g2_decap_8 FILLER_68_181 ();
 sg13g2_fill_2 FILLER_68_188 ();
 sg13g2_decap_4 FILLER_68_252 ();
 sg13g2_fill_2 FILLER_68_256 ();
 sg13g2_fill_1 FILLER_68_274 ();
 sg13g2_decap_8 FILLER_68_307 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_decap_4 FILLER_68_336 ();
 sg13g2_fill_1 FILLER_68_346 ();
 sg13g2_decap_8 FILLER_68_373 ();
 sg13g2_fill_2 FILLER_68_380 ();
 sg13g2_decap_8 FILLER_68_386 ();
 sg13g2_fill_1 FILLER_68_393 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_fill_1 FILLER_69_180 ();
 sg13g2_fill_2 FILLER_69_186 ();
 sg13g2_fill_1 FILLER_69_206 ();
 sg13g2_decap_8 FILLER_69_217 ();
 sg13g2_fill_1 FILLER_69_224 ();
 sg13g2_fill_2 FILLER_69_233 ();
 sg13g2_decap_8 FILLER_69_245 ();
 sg13g2_decap_8 FILLER_69_252 ();
 sg13g2_fill_2 FILLER_69_271 ();
 sg13g2_fill_1 FILLER_69_282 ();
 sg13g2_fill_2 FILLER_69_306 ();
 sg13g2_decap_8 FILLER_69_319 ();
 sg13g2_decap_4 FILLER_69_326 ();
 sg13g2_fill_1 FILLER_69_330 ();
 sg13g2_decap_8 FILLER_69_341 ();
 sg13g2_fill_1 FILLER_69_348 ();
 sg13g2_fill_2 FILLER_69_355 ();
 sg13g2_fill_1 FILLER_69_357 ();
 sg13g2_decap_8 FILLER_69_370 ();
 sg13g2_decap_8 FILLER_69_377 ();
 sg13g2_decap_4 FILLER_69_405 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_fill_1 FILLER_70_109 ();
 sg13g2_decap_4 FILLER_70_158 ();
 sg13g2_fill_1 FILLER_70_166 ();
 sg13g2_fill_2 FILLER_70_172 ();
 sg13g2_fill_2 FILLER_70_194 ();
 sg13g2_decap_4 FILLER_70_201 ();
 sg13g2_fill_2 FILLER_70_205 ();
 sg13g2_decap_8 FILLER_70_212 ();
 sg13g2_fill_2 FILLER_70_219 ();
 sg13g2_fill_1 FILLER_70_221 ();
 sg13g2_fill_2 FILLER_70_227 ();
 sg13g2_fill_1 FILLER_70_229 ();
 sg13g2_fill_2 FILLER_70_235 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_fill_1 FILLER_70_257 ();
 sg13g2_fill_2 FILLER_70_275 ();
 sg13g2_fill_1 FILLER_70_277 ();
 sg13g2_fill_2 FILLER_70_298 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_4 FILLER_70_322 ();
 sg13g2_decap_8 FILLER_70_352 ();
 sg13g2_fill_1 FILLER_70_359 ();
 sg13g2_decap_4 FILLER_70_366 ();
 sg13g2_decap_4 FILLER_70_376 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_4 FILLER_71_35 ();
 sg13g2_fill_1 FILLER_71_39 ();
 sg13g2_fill_2 FILLER_71_108 ();
 sg13g2_fill_2 FILLER_71_146 ();
 sg13g2_fill_1 FILLER_71_148 ();
 sg13g2_decap_4 FILLER_71_163 ();
 sg13g2_fill_1 FILLER_71_171 ();
 sg13g2_fill_1 FILLER_71_183 ();
 sg13g2_decap_8 FILLER_71_194 ();
 sg13g2_decap_4 FILLER_71_201 ();
 sg13g2_fill_2 FILLER_71_205 ();
 sg13g2_fill_1 FILLER_71_212 ();
 sg13g2_fill_2 FILLER_71_283 ();
 sg13g2_fill_1 FILLER_71_285 ();
 sg13g2_fill_1 FILLER_71_311 ();
 sg13g2_decap_4 FILLER_71_327 ();
 sg13g2_fill_2 FILLER_71_331 ();
 sg13g2_decap_8 FILLER_71_349 ();
 sg13g2_decap_8 FILLER_71_356 ();
 sg13g2_fill_2 FILLER_71_379 ();
 sg13g2_fill_1 FILLER_71_381 ();
 sg13g2_fill_1 FILLER_71_387 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_fill_2 FILLER_72_42 ();
 sg13g2_fill_2 FILLER_72_73 ();
 sg13g2_fill_2 FILLER_72_101 ();
 sg13g2_fill_2 FILLER_72_127 ();
 sg13g2_fill_2 FILLER_72_134 ();
 sg13g2_fill_2 FILLER_72_141 ();
 sg13g2_fill_1 FILLER_72_143 ();
 sg13g2_fill_2 FILLER_72_159 ();
 sg13g2_fill_1 FILLER_72_166 ();
 sg13g2_fill_2 FILLER_72_173 ();
 sg13g2_fill_1 FILLER_72_201 ();
 sg13g2_fill_1 FILLER_72_225 ();
 sg13g2_fill_2 FILLER_72_285 ();
 sg13g2_fill_1 FILLER_72_287 ();
 sg13g2_decap_8 FILLER_72_338 ();
 sg13g2_fill_1 FILLER_72_350 ();
 sg13g2_fill_1 FILLER_72_380 ();
 sg13g2_fill_2 FILLER_72_389 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_fill_1 FILLER_73_75 ();
 sg13g2_fill_2 FILLER_73_191 ();
 sg13g2_fill_2 FILLER_73_266 ();
 sg13g2_fill_2 FILLER_73_287 ();
 sg13g2_fill_1 FILLER_73_289 ();
 sg13g2_decap_8 FILLER_73_343 ();
 sg13g2_decap_8 FILLER_73_350 ();
 sg13g2_decap_4 FILLER_73_357 ();
 sg13g2_fill_2 FILLER_73_365 ();
 sg13g2_fill_2 FILLER_73_377 ();
 sg13g2_fill_2 FILLER_73_389 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_42 ();
 sg13g2_fill_2 FILLER_74_74 ();
 sg13g2_fill_1 FILLER_74_76 ();
 sg13g2_fill_2 FILLER_74_160 ();
 sg13g2_fill_1 FILLER_74_162 ();
 sg13g2_decap_8 FILLER_74_181 ();
 sg13g2_decap_8 FILLER_74_188 ();
 sg13g2_decap_8 FILLER_74_195 ();
 sg13g2_fill_2 FILLER_74_221 ();
 sg13g2_decap_8 FILLER_74_232 ();
 sg13g2_decap_4 FILLER_74_239 ();
 sg13g2_fill_2 FILLER_74_243 ();
 sg13g2_decap_8 FILLER_74_259 ();
 sg13g2_fill_2 FILLER_74_266 ();
 sg13g2_fill_1 FILLER_74_268 ();
 sg13g2_fill_2 FILLER_74_274 ();
 sg13g2_fill_1 FILLER_74_276 ();
 sg13g2_fill_1 FILLER_74_282 ();
 sg13g2_fill_1 FILLER_74_301 ();
 sg13g2_fill_2 FILLER_74_314 ();
 sg13g2_decap_8 FILLER_74_358 ();
 sg13g2_fill_1 FILLER_74_365 ();
 sg13g2_fill_1 FILLER_74_371 ();
 sg13g2_fill_1 FILLER_74_377 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_4 FILLER_75_42 ();
 sg13g2_fill_1 FILLER_75_46 ();
 sg13g2_fill_1 FILLER_75_100 ();
 sg13g2_fill_2 FILLER_75_144 ();
 sg13g2_fill_1 FILLER_75_171 ();
 sg13g2_decap_4 FILLER_75_182 ();
 sg13g2_fill_2 FILLER_75_186 ();
 sg13g2_decap_8 FILLER_75_193 ();
 sg13g2_decap_8 FILLER_75_200 ();
 sg13g2_decap_8 FILLER_75_207 ();
 sg13g2_decap_8 FILLER_75_214 ();
 sg13g2_fill_1 FILLER_75_221 ();
 sg13g2_fill_1 FILLER_75_227 ();
 sg13g2_decap_4 FILLER_75_233 ();
 sg13g2_fill_1 FILLER_75_237 ();
 sg13g2_fill_1 FILLER_75_247 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_4 FILLER_75_287 ();
 sg13g2_fill_1 FILLER_75_345 ();
 sg13g2_decap_8 FILLER_75_382 ();
 sg13g2_decap_4 FILLER_75_389 ();
 sg13g2_fill_1 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_398 ();
 sg13g2_decap_4 FILLER_75_405 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_fill_2 FILLER_76_56 ();
 sg13g2_fill_2 FILLER_76_80 ();
 sg13g2_fill_1 FILLER_76_82 ();
 sg13g2_fill_2 FILLER_76_92 ();
 sg13g2_fill_1 FILLER_76_94 ();
 sg13g2_fill_1 FILLER_76_157 ();
 sg13g2_fill_1 FILLER_76_198 ();
 sg13g2_decap_4 FILLER_76_202 ();
 sg13g2_fill_2 FILLER_76_206 ();
 sg13g2_fill_1 FILLER_76_253 ();
 sg13g2_fill_1 FILLER_76_265 ();
 sg13g2_fill_2 FILLER_76_297 ();
 sg13g2_fill_1 FILLER_76_333 ();
 sg13g2_fill_1 FILLER_76_347 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_fill_2 FILLER_77_63 ();
 sg13g2_fill_1 FILLER_77_129 ();
 sg13g2_fill_1 FILLER_77_174 ();
 sg13g2_fill_1 FILLER_77_187 ();
 sg13g2_fill_1 FILLER_77_220 ();
 sg13g2_fill_2 FILLER_77_234 ();
 sg13g2_fill_1 FILLER_77_255 ();
 sg13g2_decap_4 FILLER_77_302 ();
 sg13g2_fill_2 FILLER_77_364 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_4 FILLER_78_56 ();
 sg13g2_fill_1 FILLER_78_172 ();
 sg13g2_decap_8 FILLER_78_184 ();
 sg13g2_decap_4 FILLER_78_191 ();
 sg13g2_fill_1 FILLER_78_195 ();
 sg13g2_fill_1 FILLER_78_255 ();
 sg13g2_fill_1 FILLER_78_264 ();
 sg13g2_fill_2 FILLER_78_321 ();
 sg13g2_fill_2 FILLER_78_331 ();
 sg13g2_fill_1 FILLER_78_333 ();
 sg13g2_fill_1 FILLER_78_340 ();
 sg13g2_fill_1 FILLER_78_345 ();
 sg13g2_fill_2 FILLER_78_356 ();
 sg13g2_fill_1 FILLER_78_358 ();
 sg13g2_fill_2 FILLER_78_378 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_4 FILLER_79_63 ();
 sg13g2_fill_1 FILLER_79_67 ();
 sg13g2_fill_2 FILLER_79_138 ();
 sg13g2_fill_1 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_145 ();
 sg13g2_decap_4 FILLER_79_152 ();
 sg13g2_fill_1 FILLER_79_156 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_fill_2 FILLER_79_224 ();
 sg13g2_fill_1 FILLER_79_226 ();
 sg13g2_fill_2 FILLER_79_280 ();
 sg13g2_fill_1 FILLER_79_282 ();
 sg13g2_decap_4 FILLER_79_361 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_56 ();
 sg13g2_fill_2 FILLER_80_115 ();
 sg13g2_fill_1 FILLER_80_117 ();
 sg13g2_fill_2 FILLER_80_130 ();
 sg13g2_fill_1 FILLER_80_132 ();
 sg13g2_fill_2 FILLER_80_141 ();
 sg13g2_fill_1 FILLER_80_143 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_fill_1 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_206 ();
 sg13g2_decap_8 FILLER_80_213 ();
 sg13g2_decap_8 FILLER_80_220 ();
 sg13g2_decap_8 FILLER_80_227 ();
 sg13g2_decap_4 FILLER_80_234 ();
 sg13g2_fill_1 FILLER_80_238 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_fill_1 FILLER_80_249 ();
 sg13g2_decap_4 FILLER_80_260 ();
 sg13g2_fill_1 FILLER_80_287 ();
 sg13g2_fill_2 FILLER_80_293 ();
 sg13g2_fill_1 FILLER_80_295 ();
 sg13g2_decap_4 FILLER_80_312 ();
 sg13g2_fill_1 FILLER_80_316 ();
 sg13g2_decap_8 FILLER_80_321 ();
 sg13g2_decap_8 FILLER_80_328 ();
 sg13g2_decap_8 FILLER_80_335 ();
 sg13g2_decap_8 FILLER_80_342 ();
 sg13g2_decap_8 FILLER_80_349 ();
 sg13g2_decap_8 FILLER_80_356 ();
 sg13g2_fill_2 FILLER_80_363 ();
 sg13g2_fill_1 FILLER_80_365 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net8;
 assign uio_oe[1] = net9;
 assign uio_oe[2] = net10;
 assign uio_oe[3] = net11;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
endmodule

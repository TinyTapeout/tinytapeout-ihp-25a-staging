module tt_um_pdm_correlator_arghunter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire \u_top_module.addr[0] ;
 wire \u_top_module.addr[1] ;
 wire \u_top_module.addr[2] ;
 wire \u_top_module.addr[3] ;
 wire \u_top_module.addr[4] ;
 wire \u_top_module.addr[5] ;
 wire \u_top_module.addr[6] ;
 wire \u_top_module.addr[7] ;
 wire \u_top_module.capture_reg[0] ;
 wire \u_top_module.capture_reg[1] ;
 wire \u_top_module.capture_reg[2] ;
 wire \u_top_module.capture_reg[3] ;
 wire \u_top_module.capture_reg[4] ;
 wire \u_top_module.capture_reg[5] ;
 wire \u_top_module.capture_reg[6] ;
 wire \u_top_module.capture_reg[7] ;
 wire \u_top_module.corr_dec_clk ;
 wire \u_top_module.dec_clk ;
 wire \u_top_module.dec_data_1 ;
 wire \u_top_module.dec_data_2 ;
 wire \u_top_module.decimation_ratio[0] ;
 wire \u_top_module.decimation_ratio[1] ;
 wire \u_top_module.decimation_ratio[2] ;
 wire \u_top_module.decimation_ratio[3] ;
 wire \u_top_module.decimation_ratio[4] ;
 wire \u_top_module.decimation_ratio[5] ;
 wire \u_top_module.decimation_ratio[6] ;
 wire \u_top_module.decimation_ratio[7] ;
 wire \u_top_module.filter_length[1] ;
 wire \u_top_module.filter_length[2] ;
 wire \u_top_module.filter_length[3] ;
 wire \u_top_module.filter_length[4] ;
 wire \u_top_module.filter_length[5] ;
 wire \u_top_module.filter_length[6] ;
 wire \u_top_module.filter_length[7] ;
 wire \u_top_module.mem_out[0] ;
 wire \u_top_module.mem_out[1] ;
 wire \u_top_module.mem_out[2] ;
 wire \u_top_module.mem_out[3] ;
 wire \u_top_module.mem_out[4] ;
 wire \u_top_module.mem_out[5] ;
 wire \u_top_module.mem_out[6] ;
 wire \u_top_module.mem_out[7] ;
 wire \u_top_module.neg ;
 wire \u_top_module.pos ;
 wire \u_top_module.u_buffer.corr_neg[0] ;
 wire \u_top_module.u_buffer.corr_neg[1] ;
 wire \u_top_module.u_buffer.corr_neg[2] ;
 wire \u_top_module.u_buffer.corr_neg[3] ;
 wire \u_top_module.u_buffer.corr_neg[4] ;
 wire \u_top_module.u_buffer.corr_neg[5] ;
 wire \u_top_module.u_buffer.corr_neg[6] ;
 wire \u_top_module.u_buffer.corr_neg[7] ;
 wire \u_top_module.u_buffer.corr_pos[0] ;
 wire \u_top_module.u_buffer.corr_pos[1] ;
 wire \u_top_module.u_buffer.corr_pos[2] ;
 wire \u_top_module.u_buffer.corr_pos[3] ;
 wire \u_top_module.u_buffer.corr_pos[4] ;
 wire \u_top_module.u_buffer.corr_pos[5] ;
 wire \u_top_module.u_buffer.corr_pos[6] ;
 wire \u_top_module.u_buffer.corr_pos[7] ;
 wire \u_top_module.u_buffer.shift_reg_1[0] ;
 wire \u_top_module.u_buffer.shift_reg_1[100] ;
 wire \u_top_module.u_buffer.shift_reg_1[101] ;
 wire \u_top_module.u_buffer.shift_reg_1[102] ;
 wire \u_top_module.u_buffer.shift_reg_1[103] ;
 wire \u_top_module.u_buffer.shift_reg_1[104] ;
 wire \u_top_module.u_buffer.shift_reg_1[105] ;
 wire \u_top_module.u_buffer.shift_reg_1[106] ;
 wire \u_top_module.u_buffer.shift_reg_1[107] ;
 wire \u_top_module.u_buffer.shift_reg_1[108] ;
 wire \u_top_module.u_buffer.shift_reg_1[109] ;
 wire \u_top_module.u_buffer.shift_reg_1[10] ;
 wire \u_top_module.u_buffer.shift_reg_1[110] ;
 wire \u_top_module.u_buffer.shift_reg_1[111] ;
 wire \u_top_module.u_buffer.shift_reg_1[112] ;
 wire \u_top_module.u_buffer.shift_reg_1[113] ;
 wire \u_top_module.u_buffer.shift_reg_1[114] ;
 wire \u_top_module.u_buffer.shift_reg_1[115] ;
 wire \u_top_module.u_buffer.shift_reg_1[116] ;
 wire \u_top_module.u_buffer.shift_reg_1[117] ;
 wire \u_top_module.u_buffer.shift_reg_1[118] ;
 wire \u_top_module.u_buffer.shift_reg_1[119] ;
 wire \u_top_module.u_buffer.shift_reg_1[11] ;
 wire \u_top_module.u_buffer.shift_reg_1[120] ;
 wire \u_top_module.u_buffer.shift_reg_1[121] ;
 wire \u_top_module.u_buffer.shift_reg_1[122] ;
 wire \u_top_module.u_buffer.shift_reg_1[123] ;
 wire \u_top_module.u_buffer.shift_reg_1[124] ;
 wire \u_top_module.u_buffer.shift_reg_1[125] ;
 wire \u_top_module.u_buffer.shift_reg_1[126] ;
 wire \u_top_module.u_buffer.shift_reg_1[127] ;
 wire \u_top_module.u_buffer.shift_reg_1[128] ;
 wire \u_top_module.u_buffer.shift_reg_1[129] ;
 wire \u_top_module.u_buffer.shift_reg_1[12] ;
 wire \u_top_module.u_buffer.shift_reg_1[130] ;
 wire \u_top_module.u_buffer.shift_reg_1[131] ;
 wire \u_top_module.u_buffer.shift_reg_1[132] ;
 wire \u_top_module.u_buffer.shift_reg_1[133] ;
 wire \u_top_module.u_buffer.shift_reg_1[134] ;
 wire \u_top_module.u_buffer.shift_reg_1[135] ;
 wire \u_top_module.u_buffer.shift_reg_1[136] ;
 wire \u_top_module.u_buffer.shift_reg_1[137] ;
 wire \u_top_module.u_buffer.shift_reg_1[138] ;
 wire \u_top_module.u_buffer.shift_reg_1[139] ;
 wire \u_top_module.u_buffer.shift_reg_1[13] ;
 wire \u_top_module.u_buffer.shift_reg_1[140] ;
 wire \u_top_module.u_buffer.shift_reg_1[141] ;
 wire \u_top_module.u_buffer.shift_reg_1[142] ;
 wire \u_top_module.u_buffer.shift_reg_1[143] ;
 wire \u_top_module.u_buffer.shift_reg_1[144] ;
 wire \u_top_module.u_buffer.shift_reg_1[145] ;
 wire \u_top_module.u_buffer.shift_reg_1[146] ;
 wire \u_top_module.u_buffer.shift_reg_1[147] ;
 wire \u_top_module.u_buffer.shift_reg_1[148] ;
 wire \u_top_module.u_buffer.shift_reg_1[149] ;
 wire \u_top_module.u_buffer.shift_reg_1[14] ;
 wire \u_top_module.u_buffer.shift_reg_1[150] ;
 wire \u_top_module.u_buffer.shift_reg_1[151] ;
 wire \u_top_module.u_buffer.shift_reg_1[152] ;
 wire \u_top_module.u_buffer.shift_reg_1[153] ;
 wire \u_top_module.u_buffer.shift_reg_1[154] ;
 wire \u_top_module.u_buffer.shift_reg_1[155] ;
 wire \u_top_module.u_buffer.shift_reg_1[156] ;
 wire \u_top_module.u_buffer.shift_reg_1[157] ;
 wire \u_top_module.u_buffer.shift_reg_1[158] ;
 wire \u_top_module.u_buffer.shift_reg_1[159] ;
 wire \u_top_module.u_buffer.shift_reg_1[15] ;
 wire \u_top_module.u_buffer.shift_reg_1[160] ;
 wire \u_top_module.u_buffer.shift_reg_1[161] ;
 wire \u_top_module.u_buffer.shift_reg_1[162] ;
 wire \u_top_module.u_buffer.shift_reg_1[163] ;
 wire \u_top_module.u_buffer.shift_reg_1[164] ;
 wire \u_top_module.u_buffer.shift_reg_1[165] ;
 wire \u_top_module.u_buffer.shift_reg_1[166] ;
 wire \u_top_module.u_buffer.shift_reg_1[167] ;
 wire \u_top_module.u_buffer.shift_reg_1[168] ;
 wire \u_top_module.u_buffer.shift_reg_1[169] ;
 wire \u_top_module.u_buffer.shift_reg_1[16] ;
 wire \u_top_module.u_buffer.shift_reg_1[170] ;
 wire \u_top_module.u_buffer.shift_reg_1[171] ;
 wire \u_top_module.u_buffer.shift_reg_1[172] ;
 wire \u_top_module.u_buffer.shift_reg_1[173] ;
 wire \u_top_module.u_buffer.shift_reg_1[174] ;
 wire \u_top_module.u_buffer.shift_reg_1[175] ;
 wire \u_top_module.u_buffer.shift_reg_1[176] ;
 wire \u_top_module.u_buffer.shift_reg_1[177] ;
 wire \u_top_module.u_buffer.shift_reg_1[178] ;
 wire \u_top_module.u_buffer.shift_reg_1[179] ;
 wire \u_top_module.u_buffer.shift_reg_1[17] ;
 wire \u_top_module.u_buffer.shift_reg_1[180] ;
 wire \u_top_module.u_buffer.shift_reg_1[181] ;
 wire \u_top_module.u_buffer.shift_reg_1[182] ;
 wire \u_top_module.u_buffer.shift_reg_1[183] ;
 wire \u_top_module.u_buffer.shift_reg_1[184] ;
 wire \u_top_module.u_buffer.shift_reg_1[185] ;
 wire \u_top_module.u_buffer.shift_reg_1[186] ;
 wire \u_top_module.u_buffer.shift_reg_1[187] ;
 wire \u_top_module.u_buffer.shift_reg_1[188] ;
 wire \u_top_module.u_buffer.shift_reg_1[189] ;
 wire \u_top_module.u_buffer.shift_reg_1[18] ;
 wire \u_top_module.u_buffer.shift_reg_1[190] ;
 wire \u_top_module.u_buffer.shift_reg_1[191] ;
 wire \u_top_module.u_buffer.shift_reg_1[192] ;
 wire \u_top_module.u_buffer.shift_reg_1[193] ;
 wire \u_top_module.u_buffer.shift_reg_1[194] ;
 wire \u_top_module.u_buffer.shift_reg_1[195] ;
 wire \u_top_module.u_buffer.shift_reg_1[196] ;
 wire \u_top_module.u_buffer.shift_reg_1[197] ;
 wire \u_top_module.u_buffer.shift_reg_1[198] ;
 wire \u_top_module.u_buffer.shift_reg_1[199] ;
 wire \u_top_module.u_buffer.shift_reg_1[19] ;
 wire \u_top_module.u_buffer.shift_reg_1[1] ;
 wire \u_top_module.u_buffer.shift_reg_1[200] ;
 wire \u_top_module.u_buffer.shift_reg_1[201] ;
 wire \u_top_module.u_buffer.shift_reg_1[202] ;
 wire \u_top_module.u_buffer.shift_reg_1[203] ;
 wire \u_top_module.u_buffer.shift_reg_1[204] ;
 wire \u_top_module.u_buffer.shift_reg_1[205] ;
 wire \u_top_module.u_buffer.shift_reg_1[206] ;
 wire \u_top_module.u_buffer.shift_reg_1[207] ;
 wire \u_top_module.u_buffer.shift_reg_1[208] ;
 wire \u_top_module.u_buffer.shift_reg_1[209] ;
 wire \u_top_module.u_buffer.shift_reg_1[20] ;
 wire \u_top_module.u_buffer.shift_reg_1[210] ;
 wire \u_top_module.u_buffer.shift_reg_1[211] ;
 wire \u_top_module.u_buffer.shift_reg_1[212] ;
 wire \u_top_module.u_buffer.shift_reg_1[213] ;
 wire \u_top_module.u_buffer.shift_reg_1[214] ;
 wire \u_top_module.u_buffer.shift_reg_1[215] ;
 wire \u_top_module.u_buffer.shift_reg_1[216] ;
 wire \u_top_module.u_buffer.shift_reg_1[217] ;
 wire \u_top_module.u_buffer.shift_reg_1[218] ;
 wire \u_top_module.u_buffer.shift_reg_1[219] ;
 wire \u_top_module.u_buffer.shift_reg_1[21] ;
 wire \u_top_module.u_buffer.shift_reg_1[220] ;
 wire \u_top_module.u_buffer.shift_reg_1[221] ;
 wire \u_top_module.u_buffer.shift_reg_1[222] ;
 wire \u_top_module.u_buffer.shift_reg_1[223] ;
 wire \u_top_module.u_buffer.shift_reg_1[224] ;
 wire \u_top_module.u_buffer.shift_reg_1[225] ;
 wire \u_top_module.u_buffer.shift_reg_1[226] ;
 wire \u_top_module.u_buffer.shift_reg_1[227] ;
 wire \u_top_module.u_buffer.shift_reg_1[228] ;
 wire \u_top_module.u_buffer.shift_reg_1[229] ;
 wire \u_top_module.u_buffer.shift_reg_1[22] ;
 wire \u_top_module.u_buffer.shift_reg_1[230] ;
 wire \u_top_module.u_buffer.shift_reg_1[231] ;
 wire \u_top_module.u_buffer.shift_reg_1[232] ;
 wire \u_top_module.u_buffer.shift_reg_1[233] ;
 wire \u_top_module.u_buffer.shift_reg_1[234] ;
 wire \u_top_module.u_buffer.shift_reg_1[235] ;
 wire \u_top_module.u_buffer.shift_reg_1[236] ;
 wire \u_top_module.u_buffer.shift_reg_1[237] ;
 wire \u_top_module.u_buffer.shift_reg_1[238] ;
 wire \u_top_module.u_buffer.shift_reg_1[239] ;
 wire \u_top_module.u_buffer.shift_reg_1[23] ;
 wire \u_top_module.u_buffer.shift_reg_1[240] ;
 wire \u_top_module.u_buffer.shift_reg_1[241] ;
 wire \u_top_module.u_buffer.shift_reg_1[242] ;
 wire \u_top_module.u_buffer.shift_reg_1[243] ;
 wire \u_top_module.u_buffer.shift_reg_1[244] ;
 wire \u_top_module.u_buffer.shift_reg_1[245] ;
 wire \u_top_module.u_buffer.shift_reg_1[246] ;
 wire \u_top_module.u_buffer.shift_reg_1[247] ;
 wire \u_top_module.u_buffer.shift_reg_1[248] ;
 wire \u_top_module.u_buffer.shift_reg_1[249] ;
 wire \u_top_module.u_buffer.shift_reg_1[24] ;
 wire \u_top_module.u_buffer.shift_reg_1[250] ;
 wire \u_top_module.u_buffer.shift_reg_1[251] ;
 wire \u_top_module.u_buffer.shift_reg_1[252] ;
 wire \u_top_module.u_buffer.shift_reg_1[253] ;
 wire \u_top_module.u_buffer.shift_reg_1[254] ;
 wire \u_top_module.u_buffer.shift_reg_1[255] ;
 wire \u_top_module.u_buffer.shift_reg_1[25] ;
 wire \u_top_module.u_buffer.shift_reg_1[26] ;
 wire \u_top_module.u_buffer.shift_reg_1[27] ;
 wire \u_top_module.u_buffer.shift_reg_1[28] ;
 wire \u_top_module.u_buffer.shift_reg_1[29] ;
 wire \u_top_module.u_buffer.shift_reg_1[2] ;
 wire \u_top_module.u_buffer.shift_reg_1[30] ;
 wire \u_top_module.u_buffer.shift_reg_1[31] ;
 wire \u_top_module.u_buffer.shift_reg_1[32] ;
 wire \u_top_module.u_buffer.shift_reg_1[33] ;
 wire \u_top_module.u_buffer.shift_reg_1[34] ;
 wire \u_top_module.u_buffer.shift_reg_1[35] ;
 wire \u_top_module.u_buffer.shift_reg_1[36] ;
 wire \u_top_module.u_buffer.shift_reg_1[37] ;
 wire \u_top_module.u_buffer.shift_reg_1[38] ;
 wire \u_top_module.u_buffer.shift_reg_1[39] ;
 wire \u_top_module.u_buffer.shift_reg_1[3] ;
 wire \u_top_module.u_buffer.shift_reg_1[40] ;
 wire \u_top_module.u_buffer.shift_reg_1[41] ;
 wire \u_top_module.u_buffer.shift_reg_1[42] ;
 wire \u_top_module.u_buffer.shift_reg_1[43] ;
 wire \u_top_module.u_buffer.shift_reg_1[44] ;
 wire \u_top_module.u_buffer.shift_reg_1[45] ;
 wire \u_top_module.u_buffer.shift_reg_1[46] ;
 wire \u_top_module.u_buffer.shift_reg_1[47] ;
 wire \u_top_module.u_buffer.shift_reg_1[48] ;
 wire \u_top_module.u_buffer.shift_reg_1[49] ;
 wire \u_top_module.u_buffer.shift_reg_1[4] ;
 wire \u_top_module.u_buffer.shift_reg_1[50] ;
 wire \u_top_module.u_buffer.shift_reg_1[51] ;
 wire \u_top_module.u_buffer.shift_reg_1[52] ;
 wire \u_top_module.u_buffer.shift_reg_1[53] ;
 wire \u_top_module.u_buffer.shift_reg_1[54] ;
 wire \u_top_module.u_buffer.shift_reg_1[55] ;
 wire \u_top_module.u_buffer.shift_reg_1[56] ;
 wire \u_top_module.u_buffer.shift_reg_1[57] ;
 wire \u_top_module.u_buffer.shift_reg_1[58] ;
 wire \u_top_module.u_buffer.shift_reg_1[59] ;
 wire \u_top_module.u_buffer.shift_reg_1[5] ;
 wire \u_top_module.u_buffer.shift_reg_1[60] ;
 wire \u_top_module.u_buffer.shift_reg_1[61] ;
 wire \u_top_module.u_buffer.shift_reg_1[62] ;
 wire \u_top_module.u_buffer.shift_reg_1[63] ;
 wire \u_top_module.u_buffer.shift_reg_1[64] ;
 wire \u_top_module.u_buffer.shift_reg_1[65] ;
 wire \u_top_module.u_buffer.shift_reg_1[66] ;
 wire \u_top_module.u_buffer.shift_reg_1[67] ;
 wire \u_top_module.u_buffer.shift_reg_1[68] ;
 wire \u_top_module.u_buffer.shift_reg_1[69] ;
 wire \u_top_module.u_buffer.shift_reg_1[6] ;
 wire \u_top_module.u_buffer.shift_reg_1[70] ;
 wire \u_top_module.u_buffer.shift_reg_1[71] ;
 wire \u_top_module.u_buffer.shift_reg_1[72] ;
 wire \u_top_module.u_buffer.shift_reg_1[73] ;
 wire \u_top_module.u_buffer.shift_reg_1[74] ;
 wire \u_top_module.u_buffer.shift_reg_1[75] ;
 wire \u_top_module.u_buffer.shift_reg_1[76] ;
 wire \u_top_module.u_buffer.shift_reg_1[77] ;
 wire \u_top_module.u_buffer.shift_reg_1[78] ;
 wire \u_top_module.u_buffer.shift_reg_1[79] ;
 wire \u_top_module.u_buffer.shift_reg_1[7] ;
 wire \u_top_module.u_buffer.shift_reg_1[80] ;
 wire \u_top_module.u_buffer.shift_reg_1[81] ;
 wire \u_top_module.u_buffer.shift_reg_1[82] ;
 wire \u_top_module.u_buffer.shift_reg_1[83] ;
 wire \u_top_module.u_buffer.shift_reg_1[84] ;
 wire \u_top_module.u_buffer.shift_reg_1[85] ;
 wire \u_top_module.u_buffer.shift_reg_1[86] ;
 wire \u_top_module.u_buffer.shift_reg_1[87] ;
 wire \u_top_module.u_buffer.shift_reg_1[88] ;
 wire \u_top_module.u_buffer.shift_reg_1[89] ;
 wire \u_top_module.u_buffer.shift_reg_1[8] ;
 wire \u_top_module.u_buffer.shift_reg_1[90] ;
 wire \u_top_module.u_buffer.shift_reg_1[91] ;
 wire \u_top_module.u_buffer.shift_reg_1[92] ;
 wire \u_top_module.u_buffer.shift_reg_1[93] ;
 wire \u_top_module.u_buffer.shift_reg_1[94] ;
 wire \u_top_module.u_buffer.shift_reg_1[95] ;
 wire \u_top_module.u_buffer.shift_reg_1[96] ;
 wire \u_top_module.u_buffer.shift_reg_1[97] ;
 wire \u_top_module.u_buffer.shift_reg_1[98] ;
 wire \u_top_module.u_buffer.shift_reg_1[99] ;
 wire \u_top_module.u_buffer.shift_reg_1[9] ;
 wire \u_top_module.u_buffer.shift_reg_2[0] ;
 wire \u_top_module.u_buffer.shift_reg_2[100] ;
 wire \u_top_module.u_buffer.shift_reg_2[101] ;
 wire \u_top_module.u_buffer.shift_reg_2[102] ;
 wire \u_top_module.u_buffer.shift_reg_2[103] ;
 wire \u_top_module.u_buffer.shift_reg_2[104] ;
 wire \u_top_module.u_buffer.shift_reg_2[105] ;
 wire \u_top_module.u_buffer.shift_reg_2[106] ;
 wire \u_top_module.u_buffer.shift_reg_2[107] ;
 wire \u_top_module.u_buffer.shift_reg_2[108] ;
 wire \u_top_module.u_buffer.shift_reg_2[109] ;
 wire \u_top_module.u_buffer.shift_reg_2[10] ;
 wire \u_top_module.u_buffer.shift_reg_2[110] ;
 wire \u_top_module.u_buffer.shift_reg_2[111] ;
 wire \u_top_module.u_buffer.shift_reg_2[112] ;
 wire \u_top_module.u_buffer.shift_reg_2[113] ;
 wire \u_top_module.u_buffer.shift_reg_2[114] ;
 wire \u_top_module.u_buffer.shift_reg_2[115] ;
 wire \u_top_module.u_buffer.shift_reg_2[116] ;
 wire \u_top_module.u_buffer.shift_reg_2[117] ;
 wire \u_top_module.u_buffer.shift_reg_2[118] ;
 wire \u_top_module.u_buffer.shift_reg_2[119] ;
 wire \u_top_module.u_buffer.shift_reg_2[11] ;
 wire \u_top_module.u_buffer.shift_reg_2[120] ;
 wire \u_top_module.u_buffer.shift_reg_2[121] ;
 wire \u_top_module.u_buffer.shift_reg_2[122] ;
 wire \u_top_module.u_buffer.shift_reg_2[123] ;
 wire \u_top_module.u_buffer.shift_reg_2[124] ;
 wire \u_top_module.u_buffer.shift_reg_2[125] ;
 wire \u_top_module.u_buffer.shift_reg_2[126] ;
 wire \u_top_module.u_buffer.shift_reg_2[127] ;
 wire \u_top_module.u_buffer.shift_reg_2[128] ;
 wire \u_top_module.u_buffer.shift_reg_2[129] ;
 wire \u_top_module.u_buffer.shift_reg_2[12] ;
 wire \u_top_module.u_buffer.shift_reg_2[130] ;
 wire \u_top_module.u_buffer.shift_reg_2[131] ;
 wire \u_top_module.u_buffer.shift_reg_2[132] ;
 wire \u_top_module.u_buffer.shift_reg_2[133] ;
 wire \u_top_module.u_buffer.shift_reg_2[134] ;
 wire \u_top_module.u_buffer.shift_reg_2[135] ;
 wire \u_top_module.u_buffer.shift_reg_2[136] ;
 wire \u_top_module.u_buffer.shift_reg_2[137] ;
 wire \u_top_module.u_buffer.shift_reg_2[138] ;
 wire \u_top_module.u_buffer.shift_reg_2[139] ;
 wire \u_top_module.u_buffer.shift_reg_2[13] ;
 wire \u_top_module.u_buffer.shift_reg_2[140] ;
 wire \u_top_module.u_buffer.shift_reg_2[141] ;
 wire \u_top_module.u_buffer.shift_reg_2[142] ;
 wire \u_top_module.u_buffer.shift_reg_2[143] ;
 wire \u_top_module.u_buffer.shift_reg_2[144] ;
 wire \u_top_module.u_buffer.shift_reg_2[145] ;
 wire \u_top_module.u_buffer.shift_reg_2[146] ;
 wire \u_top_module.u_buffer.shift_reg_2[147] ;
 wire \u_top_module.u_buffer.shift_reg_2[148] ;
 wire \u_top_module.u_buffer.shift_reg_2[149] ;
 wire \u_top_module.u_buffer.shift_reg_2[14] ;
 wire \u_top_module.u_buffer.shift_reg_2[150] ;
 wire \u_top_module.u_buffer.shift_reg_2[151] ;
 wire \u_top_module.u_buffer.shift_reg_2[152] ;
 wire \u_top_module.u_buffer.shift_reg_2[153] ;
 wire \u_top_module.u_buffer.shift_reg_2[154] ;
 wire \u_top_module.u_buffer.shift_reg_2[155] ;
 wire \u_top_module.u_buffer.shift_reg_2[156] ;
 wire \u_top_module.u_buffer.shift_reg_2[157] ;
 wire \u_top_module.u_buffer.shift_reg_2[158] ;
 wire \u_top_module.u_buffer.shift_reg_2[159] ;
 wire \u_top_module.u_buffer.shift_reg_2[15] ;
 wire \u_top_module.u_buffer.shift_reg_2[160] ;
 wire \u_top_module.u_buffer.shift_reg_2[161] ;
 wire \u_top_module.u_buffer.shift_reg_2[162] ;
 wire \u_top_module.u_buffer.shift_reg_2[163] ;
 wire \u_top_module.u_buffer.shift_reg_2[164] ;
 wire \u_top_module.u_buffer.shift_reg_2[165] ;
 wire \u_top_module.u_buffer.shift_reg_2[166] ;
 wire \u_top_module.u_buffer.shift_reg_2[167] ;
 wire \u_top_module.u_buffer.shift_reg_2[168] ;
 wire \u_top_module.u_buffer.shift_reg_2[169] ;
 wire \u_top_module.u_buffer.shift_reg_2[16] ;
 wire \u_top_module.u_buffer.shift_reg_2[170] ;
 wire \u_top_module.u_buffer.shift_reg_2[171] ;
 wire \u_top_module.u_buffer.shift_reg_2[172] ;
 wire \u_top_module.u_buffer.shift_reg_2[173] ;
 wire \u_top_module.u_buffer.shift_reg_2[174] ;
 wire \u_top_module.u_buffer.shift_reg_2[175] ;
 wire \u_top_module.u_buffer.shift_reg_2[176] ;
 wire \u_top_module.u_buffer.shift_reg_2[177] ;
 wire \u_top_module.u_buffer.shift_reg_2[178] ;
 wire \u_top_module.u_buffer.shift_reg_2[179] ;
 wire \u_top_module.u_buffer.shift_reg_2[17] ;
 wire \u_top_module.u_buffer.shift_reg_2[180] ;
 wire \u_top_module.u_buffer.shift_reg_2[181] ;
 wire \u_top_module.u_buffer.shift_reg_2[182] ;
 wire \u_top_module.u_buffer.shift_reg_2[183] ;
 wire \u_top_module.u_buffer.shift_reg_2[184] ;
 wire \u_top_module.u_buffer.shift_reg_2[185] ;
 wire \u_top_module.u_buffer.shift_reg_2[186] ;
 wire \u_top_module.u_buffer.shift_reg_2[187] ;
 wire \u_top_module.u_buffer.shift_reg_2[188] ;
 wire \u_top_module.u_buffer.shift_reg_2[189] ;
 wire \u_top_module.u_buffer.shift_reg_2[18] ;
 wire \u_top_module.u_buffer.shift_reg_2[190] ;
 wire \u_top_module.u_buffer.shift_reg_2[191] ;
 wire \u_top_module.u_buffer.shift_reg_2[192] ;
 wire \u_top_module.u_buffer.shift_reg_2[193] ;
 wire \u_top_module.u_buffer.shift_reg_2[194] ;
 wire \u_top_module.u_buffer.shift_reg_2[195] ;
 wire \u_top_module.u_buffer.shift_reg_2[196] ;
 wire \u_top_module.u_buffer.shift_reg_2[197] ;
 wire \u_top_module.u_buffer.shift_reg_2[198] ;
 wire \u_top_module.u_buffer.shift_reg_2[199] ;
 wire \u_top_module.u_buffer.shift_reg_2[19] ;
 wire \u_top_module.u_buffer.shift_reg_2[1] ;
 wire \u_top_module.u_buffer.shift_reg_2[200] ;
 wire \u_top_module.u_buffer.shift_reg_2[201] ;
 wire \u_top_module.u_buffer.shift_reg_2[202] ;
 wire \u_top_module.u_buffer.shift_reg_2[203] ;
 wire \u_top_module.u_buffer.shift_reg_2[204] ;
 wire \u_top_module.u_buffer.shift_reg_2[205] ;
 wire \u_top_module.u_buffer.shift_reg_2[206] ;
 wire \u_top_module.u_buffer.shift_reg_2[207] ;
 wire \u_top_module.u_buffer.shift_reg_2[208] ;
 wire \u_top_module.u_buffer.shift_reg_2[209] ;
 wire \u_top_module.u_buffer.shift_reg_2[20] ;
 wire \u_top_module.u_buffer.shift_reg_2[210] ;
 wire \u_top_module.u_buffer.shift_reg_2[211] ;
 wire \u_top_module.u_buffer.shift_reg_2[212] ;
 wire \u_top_module.u_buffer.shift_reg_2[213] ;
 wire \u_top_module.u_buffer.shift_reg_2[214] ;
 wire \u_top_module.u_buffer.shift_reg_2[215] ;
 wire \u_top_module.u_buffer.shift_reg_2[216] ;
 wire \u_top_module.u_buffer.shift_reg_2[217] ;
 wire \u_top_module.u_buffer.shift_reg_2[218] ;
 wire \u_top_module.u_buffer.shift_reg_2[219] ;
 wire \u_top_module.u_buffer.shift_reg_2[21] ;
 wire \u_top_module.u_buffer.shift_reg_2[220] ;
 wire \u_top_module.u_buffer.shift_reg_2[221] ;
 wire \u_top_module.u_buffer.shift_reg_2[222] ;
 wire \u_top_module.u_buffer.shift_reg_2[223] ;
 wire \u_top_module.u_buffer.shift_reg_2[224] ;
 wire \u_top_module.u_buffer.shift_reg_2[225] ;
 wire \u_top_module.u_buffer.shift_reg_2[226] ;
 wire \u_top_module.u_buffer.shift_reg_2[227] ;
 wire \u_top_module.u_buffer.shift_reg_2[228] ;
 wire \u_top_module.u_buffer.shift_reg_2[229] ;
 wire \u_top_module.u_buffer.shift_reg_2[22] ;
 wire \u_top_module.u_buffer.shift_reg_2[230] ;
 wire \u_top_module.u_buffer.shift_reg_2[231] ;
 wire \u_top_module.u_buffer.shift_reg_2[232] ;
 wire \u_top_module.u_buffer.shift_reg_2[233] ;
 wire \u_top_module.u_buffer.shift_reg_2[234] ;
 wire \u_top_module.u_buffer.shift_reg_2[235] ;
 wire \u_top_module.u_buffer.shift_reg_2[236] ;
 wire \u_top_module.u_buffer.shift_reg_2[237] ;
 wire \u_top_module.u_buffer.shift_reg_2[238] ;
 wire \u_top_module.u_buffer.shift_reg_2[239] ;
 wire \u_top_module.u_buffer.shift_reg_2[23] ;
 wire \u_top_module.u_buffer.shift_reg_2[240] ;
 wire \u_top_module.u_buffer.shift_reg_2[241] ;
 wire \u_top_module.u_buffer.shift_reg_2[242] ;
 wire \u_top_module.u_buffer.shift_reg_2[243] ;
 wire \u_top_module.u_buffer.shift_reg_2[244] ;
 wire \u_top_module.u_buffer.shift_reg_2[245] ;
 wire \u_top_module.u_buffer.shift_reg_2[246] ;
 wire \u_top_module.u_buffer.shift_reg_2[247] ;
 wire \u_top_module.u_buffer.shift_reg_2[248] ;
 wire \u_top_module.u_buffer.shift_reg_2[249] ;
 wire \u_top_module.u_buffer.shift_reg_2[24] ;
 wire \u_top_module.u_buffer.shift_reg_2[250] ;
 wire \u_top_module.u_buffer.shift_reg_2[251] ;
 wire \u_top_module.u_buffer.shift_reg_2[252] ;
 wire \u_top_module.u_buffer.shift_reg_2[253] ;
 wire \u_top_module.u_buffer.shift_reg_2[254] ;
 wire \u_top_module.u_buffer.shift_reg_2[255] ;
 wire \u_top_module.u_buffer.shift_reg_2[25] ;
 wire \u_top_module.u_buffer.shift_reg_2[26] ;
 wire \u_top_module.u_buffer.shift_reg_2[27] ;
 wire \u_top_module.u_buffer.shift_reg_2[28] ;
 wire \u_top_module.u_buffer.shift_reg_2[29] ;
 wire \u_top_module.u_buffer.shift_reg_2[2] ;
 wire \u_top_module.u_buffer.shift_reg_2[30] ;
 wire \u_top_module.u_buffer.shift_reg_2[31] ;
 wire \u_top_module.u_buffer.shift_reg_2[32] ;
 wire \u_top_module.u_buffer.shift_reg_2[33] ;
 wire \u_top_module.u_buffer.shift_reg_2[34] ;
 wire \u_top_module.u_buffer.shift_reg_2[35] ;
 wire \u_top_module.u_buffer.shift_reg_2[36] ;
 wire \u_top_module.u_buffer.shift_reg_2[37] ;
 wire \u_top_module.u_buffer.shift_reg_2[38] ;
 wire \u_top_module.u_buffer.shift_reg_2[39] ;
 wire \u_top_module.u_buffer.shift_reg_2[3] ;
 wire \u_top_module.u_buffer.shift_reg_2[40] ;
 wire \u_top_module.u_buffer.shift_reg_2[41] ;
 wire \u_top_module.u_buffer.shift_reg_2[42] ;
 wire \u_top_module.u_buffer.shift_reg_2[43] ;
 wire \u_top_module.u_buffer.shift_reg_2[44] ;
 wire \u_top_module.u_buffer.shift_reg_2[45] ;
 wire \u_top_module.u_buffer.shift_reg_2[46] ;
 wire \u_top_module.u_buffer.shift_reg_2[47] ;
 wire \u_top_module.u_buffer.shift_reg_2[48] ;
 wire \u_top_module.u_buffer.shift_reg_2[49] ;
 wire \u_top_module.u_buffer.shift_reg_2[4] ;
 wire \u_top_module.u_buffer.shift_reg_2[50] ;
 wire \u_top_module.u_buffer.shift_reg_2[51] ;
 wire \u_top_module.u_buffer.shift_reg_2[52] ;
 wire \u_top_module.u_buffer.shift_reg_2[53] ;
 wire \u_top_module.u_buffer.shift_reg_2[54] ;
 wire \u_top_module.u_buffer.shift_reg_2[55] ;
 wire \u_top_module.u_buffer.shift_reg_2[56] ;
 wire \u_top_module.u_buffer.shift_reg_2[57] ;
 wire \u_top_module.u_buffer.shift_reg_2[58] ;
 wire \u_top_module.u_buffer.shift_reg_2[59] ;
 wire \u_top_module.u_buffer.shift_reg_2[5] ;
 wire \u_top_module.u_buffer.shift_reg_2[60] ;
 wire \u_top_module.u_buffer.shift_reg_2[61] ;
 wire \u_top_module.u_buffer.shift_reg_2[62] ;
 wire \u_top_module.u_buffer.shift_reg_2[63] ;
 wire \u_top_module.u_buffer.shift_reg_2[64] ;
 wire \u_top_module.u_buffer.shift_reg_2[65] ;
 wire \u_top_module.u_buffer.shift_reg_2[66] ;
 wire \u_top_module.u_buffer.shift_reg_2[67] ;
 wire \u_top_module.u_buffer.shift_reg_2[68] ;
 wire \u_top_module.u_buffer.shift_reg_2[69] ;
 wire \u_top_module.u_buffer.shift_reg_2[6] ;
 wire \u_top_module.u_buffer.shift_reg_2[70] ;
 wire \u_top_module.u_buffer.shift_reg_2[71] ;
 wire \u_top_module.u_buffer.shift_reg_2[72] ;
 wire \u_top_module.u_buffer.shift_reg_2[73] ;
 wire \u_top_module.u_buffer.shift_reg_2[74] ;
 wire \u_top_module.u_buffer.shift_reg_2[75] ;
 wire \u_top_module.u_buffer.shift_reg_2[76] ;
 wire \u_top_module.u_buffer.shift_reg_2[77] ;
 wire \u_top_module.u_buffer.shift_reg_2[78] ;
 wire \u_top_module.u_buffer.shift_reg_2[79] ;
 wire \u_top_module.u_buffer.shift_reg_2[7] ;
 wire \u_top_module.u_buffer.shift_reg_2[80] ;
 wire \u_top_module.u_buffer.shift_reg_2[81] ;
 wire \u_top_module.u_buffer.shift_reg_2[82] ;
 wire \u_top_module.u_buffer.shift_reg_2[83] ;
 wire \u_top_module.u_buffer.shift_reg_2[84] ;
 wire \u_top_module.u_buffer.shift_reg_2[85] ;
 wire \u_top_module.u_buffer.shift_reg_2[86] ;
 wire \u_top_module.u_buffer.shift_reg_2[87] ;
 wire \u_top_module.u_buffer.shift_reg_2[88] ;
 wire \u_top_module.u_buffer.shift_reg_2[89] ;
 wire \u_top_module.u_buffer.shift_reg_2[8] ;
 wire \u_top_module.u_buffer.shift_reg_2[90] ;
 wire \u_top_module.u_buffer.shift_reg_2[91] ;
 wire \u_top_module.u_buffer.shift_reg_2[92] ;
 wire \u_top_module.u_buffer.shift_reg_2[93] ;
 wire \u_top_module.u_buffer.shift_reg_2[94] ;
 wire \u_top_module.u_buffer.shift_reg_2[95] ;
 wire \u_top_module.u_buffer.shift_reg_2[96] ;
 wire \u_top_module.u_buffer.shift_reg_2[97] ;
 wire \u_top_module.u_buffer.shift_reg_2[98] ;
 wire \u_top_module.u_buffer.shift_reg_2[99] ;
 wire \u_top_module.u_buffer.shift_reg_2[9] ;
 wire \u_top_module.u_decimator_1.counter[0] ;
 wire \u_top_module.u_decimator_1.counter[1] ;
 wire \u_top_module.u_decimator_1.counter[2] ;
 wire \u_top_module.u_decimator_1.counter[3] ;
 wire \u_top_module.u_decimator_1.counter[4] ;
 wire \u_top_module.u_decimator_1.counter[5] ;
 wire \u_top_module.u_decimator_1.counter[6] ;
 wire \u_top_module.u_decimator_1.counter[7] ;
 wire \u_top_module.u_decimator_2.counter[0] ;
 wire \u_top_module.u_decimator_2.counter[1] ;
 wire \u_top_module.u_decimator_2.counter[2] ;
 wire \u_top_module.u_decimator_2.counter[3] ;
 wire \u_top_module.u_decimator_2.counter[4] ;
 wire \u_top_module.u_decimator_2.counter[5] ;
 wire \u_top_module.u_decimator_2.counter[6] ;
 wire \u_top_module.u_decimator_2.counter[7] ;
 wire \u_top_module.u_memory.memory[0][0] ;
 wire \u_top_module.u_memory.memory[0][1] ;
 wire \u_top_module.u_memory.memory[0][2] ;
 wire \u_top_module.u_memory.memory[0][3] ;
 wire \u_top_module.u_memory.memory[0][4] ;
 wire \u_top_module.u_memory.memory[0][5] ;
 wire \u_top_module.u_memory.memory[0][6] ;
 wire \u_top_module.u_memory.memory[0][7] ;
 wire \u_top_module.u_memory.memory[1][0] ;
 wire \u_top_module.u_memory.memory[1][1] ;
 wire \u_top_module.u_memory.memory[1][2] ;
 wire \u_top_module.u_memory.memory[1][3] ;
 wire \u_top_module.u_memory.memory[1][4] ;
 wire \u_top_module.u_memory.memory[1][5] ;
 wire \u_top_module.u_memory.memory[1][6] ;
 wire \u_top_module.u_memory.memory[1][7] ;
 wire \u_top_module.u_memory.memory[2][0] ;
 wire \u_top_module.u_memory.memory[2][1] ;
 wire \u_top_module.u_memory.memory[2][2] ;
 wire \u_top_module.u_memory.memory[2][3] ;
 wire \u_top_module.u_memory.memory[2][4] ;
 wire \u_top_module.u_memory.memory[2][5] ;
 wire \u_top_module.u_memory.memory[2][6] ;
 wire \u_top_module.u_memory.memory[2][7] ;
 wire \u_top_module.u_memory.memory[3][0] ;
 wire \u_top_module.u_memory.memory[3][1] ;
 wire \u_top_module.u_memory.memory[3][2] ;
 wire \u_top_module.u_memory.memory[3][3] ;
 wire \u_top_module.u_memory.memory[3][4] ;
 wire \u_top_module.u_memory.memory[3][5] ;
 wire \u_top_module.u_memory.memory[3][6] ;
 wire \u_top_module.u_memory.memory[3][7] ;
 wire \u_top_module.u_memory.memory[4][0] ;
 wire \u_top_module.u_memory.memory[4][1] ;
 wire \u_top_module.u_memory.memory[4][2] ;
 wire \u_top_module.u_memory.memory[4][3] ;
 wire \u_top_module.u_memory.memory[4][4] ;
 wire \u_top_module.u_memory.memory[4][5] ;
 wire \u_top_module.u_memory.memory[4][6] ;
 wire \u_top_module.u_memory.memory[4][7] ;
 wire \u_top_module.u_memory.memory[5][0] ;
 wire \u_top_module.u_memory.memory[5][1] ;
 wire \u_top_module.u_memory.memory[5][2] ;
 wire \u_top_module.u_memory.memory[5][3] ;
 wire \u_top_module.u_memory.memory[5][4] ;
 wire \u_top_module.u_memory.memory[5][5] ;
 wire \u_top_module.u_memory.memory[5][6] ;
 wire \u_top_module.u_memory.memory[5][7] ;
 wire \u_top_module.u_memory.memory[6][0] ;
 wire \u_top_module.u_memory.memory[6][1] ;
 wire \u_top_module.u_memory.memory[6][2] ;
 wire \u_top_module.u_memory.memory[6][3] ;
 wire \u_top_module.u_memory.memory[6][4] ;
 wire \u_top_module.u_memory.memory[6][5] ;
 wire \u_top_module.u_memory.memory[6][6] ;
 wire \u_top_module.u_memory.memory[6][7] ;
 wire \u_top_module.u_memory.memory[7][0] ;
 wire \u_top_module.u_memory.memory[7][1] ;
 wire \u_top_module.u_memory.memory[7][2] ;
 wire \u_top_module.u_memory.memory[7][3] ;
 wire \u_top_module.u_memory.memory[7][4] ;
 wire \u_top_module.u_memory.memory[7][5] ;
 wire \u_top_module.u_memory.memory[7][6] ;
 wire \u_top_module.u_memory.memory[7][7] ;
 wire \u_top_module.u_spi_port.cs_n_prev ;
 wire \u_top_module.u_spi_port.shift_reg[0] ;
 wire \u_top_module.u_spi_port.shift_reg[10] ;
 wire \u_top_module.u_spi_port.shift_reg[11] ;
 wire \u_top_module.u_spi_port.shift_reg[12] ;
 wire \u_top_module.u_spi_port.shift_reg[13] ;
 wire \u_top_module.u_spi_port.shift_reg[14] ;
 wire \u_top_module.u_spi_port.shift_reg[15] ;
 wire \u_top_module.u_spi_port.shift_reg[1] ;
 wire \u_top_module.u_spi_port.shift_reg[2] ;
 wire \u_top_module.u_spi_port.shift_reg[3] ;
 wire \u_top_module.u_spi_port.shift_reg[4] ;
 wire \u_top_module.u_spi_port.shift_reg[5] ;
 wire \u_top_module.u_spi_port.shift_reg[6] ;
 wire \u_top_module.u_spi_port.shift_reg[7] ;
 wire \u_top_module.u_spi_port.shift_reg[8] ;
 wire \u_top_module.u_spi_port.shift_reg[9] ;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;

 sg13g2_inv_1 _1164_ (.Y(_0026_),
    .A(net2));
 sg13g2_inv_1 _1165_ (.Y(_0166_),
    .A(\u_top_module.addr[1] ));
 sg13g2_inv_1 _1166_ (.Y(_0167_),
    .A(\u_top_module.u_decimator_2.counter[3] ));
 sg13g2_inv_1 _1167_ (.Y(_0168_),
    .A(\u_top_module.u_decimator_2.counter[4] ));
 sg13g2_inv_1 _1168_ (.Y(_0169_),
    .A(_0008_));
 sg13g2_inv_1 _1169_ (.Y(_0170_),
    .A(\u_top_module.u_decimator_1.counter[4] ));
 sg13g2_inv_1 _1170_ (.Y(_0171_),
    .A(\u_top_module.u_decimator_1.counter[3] ));
 sg13g2_inv_1 _1171_ (.Y(_0172_),
    .A(\u_top_module.u_decimator_1.counter[2] ));
 sg13g2_inv_1 _1172_ (.Y(_0173_),
    .A(_0011_));
 sg13g2_inv_1 _1173_ (.Y(_0174_),
    .A(\u_top_module.u_memory.memory[0][0] ));
 sg13g2_inv_1 _1174_ (.Y(_0175_),
    .A(\u_top_module.u_buffer.corr_pos[7] ));
 sg13g2_inv_1 _1175_ (.Y(_0176_),
    .A(\u_top_module.u_buffer.corr_pos[6] ));
 sg13g2_inv_1 _1176_ (.Y(_0177_),
    .A(\u_top_module.u_buffer.corr_neg[6] ));
 sg13g2_inv_1 _1177_ (.Y(_0178_),
    .A(\u_top_module.u_buffer.corr_pos[5] ));
 sg13g2_inv_1 _1178_ (.Y(_0179_),
    .A(net821));
 sg13g2_inv_1 _1179_ (.Y(_0180_),
    .A(\u_top_module.u_buffer.corr_neg[4] ));
 sg13g2_inv_1 _1180_ (.Y(_0181_),
    .A(\u_top_module.u_buffer.corr_pos[4] ));
 sg13g2_inv_1 _1181_ (.Y(_0182_),
    .A(\u_top_module.u_buffer.corr_pos[3] ));
 sg13g2_inv_1 _1182_ (.Y(_0183_),
    .A(\u_top_module.u_buffer.corr_neg[3] ));
 sg13g2_inv_1 _1183_ (.Y(_0184_),
    .A(\u_top_module.u_buffer.corr_pos[2] ));
 sg13g2_inv_1 _1184_ (.Y(_0185_),
    .A(\u_top_module.u_buffer.corr_neg[2] ));
 sg13g2_inv_1 _1185_ (.Y(_0186_),
    .A(\u_top_module.u_buffer.corr_pos[1] ));
 sg13g2_inv_1 _1186_ (.Y(_0187_),
    .A(\u_top_module.u_buffer.corr_neg[1] ));
 sg13g2_inv_1 _1187_ (.Y(_0188_),
    .A(\u_top_module.u_buffer.corr_neg[0] ));
 sg13g2_inv_1 _1188_ (.Y(_0189_),
    .A(uo_out[3]));
 sg13g2_inv_1 _1189_ (.Y(_0190_),
    .A(uo_out[5]));
 sg13g2_nor2_1 _1190_ (.A(\u_top_module.addr[3] ),
    .B(\u_top_module.addr[2] ),
    .Y(_0191_));
 sg13g2_nor4_2 _1191_ (.A(\u_top_module.addr[5] ),
    .B(\u_top_module.addr[4] ),
    .C(\u_top_module.addr[7] ),
    .Y(_0192_),
    .D(\u_top_module.addr[6] ));
 sg13g2_nand2_1 _1192_ (.Y(_0193_),
    .A(_0166_),
    .B(\u_top_module.addr[0] ));
 sg13g2_nand4_1 _1193_ (.B(\u_top_module.addr[0] ),
    .C(_0191_),
    .A(_0166_),
    .Y(_0002_),
    .D(_0192_));
 sg13g2_nor2_2 _1194_ (.A(\u_top_module.addr[1] ),
    .B(\u_top_module.addr[0] ),
    .Y(_0194_));
 sg13g2_nand3_1 _1195_ (.B(_0192_),
    .C(_0194_),
    .A(_0191_),
    .Y(_0001_));
 sg13g2_nor3_1 _1196_ (.A(\u_top_module.decimation_ratio[1] ),
    .B(\u_top_module.decimation_ratio[3] ),
    .C(\u_top_module.decimation_ratio[2] ),
    .Y(_0195_));
 sg13g2_nand2b_1 _1197_ (.Y(_0196_),
    .B(\u_top_module.decimation_ratio[0] ),
    .A_N(\u_top_module.decimation_ratio[7] ));
 sg13g2_nor4_2 _1198_ (.A(\u_top_module.decimation_ratio[5] ),
    .B(\u_top_module.decimation_ratio[4] ),
    .C(\u_top_module.decimation_ratio[6] ),
    .Y(_0197_),
    .D(_0196_));
 sg13g2_and2_1 _1199_ (.A(_0195_),
    .B(_0197_),
    .X(_0198_));
 sg13g2_nand2_2 _1200_ (.Y(_0199_),
    .A(_0195_),
    .B(_0197_));
 sg13g2_mux2_2 _1201_ (.A0(net969),
    .A1(\u_top_module.dec_clk ),
    .S(_0199_),
    .X(\u_top_module.corr_dec_clk ));
 sg13g2_nor2_1 _1202_ (.A(\u_top_module.addr[2] ),
    .B(_0194_),
    .Y(_0200_));
 sg13g2_nor2b_2 _1203_ (.A(_0200_),
    .B_N(_0005_),
    .Y(_0201_));
 sg13g2_o21ai_1 _1204_ (.B1(_0005_),
    .Y(_0202_),
    .A1(\u_top_module.addr[2] ),
    .A2(_0194_));
 sg13g2_nor2_1 _1205_ (.A(\u_top_module.addr[2] ),
    .B(_0193_),
    .Y(_0203_));
 sg13g2_nand2_1 _1206_ (.Y(_0204_),
    .A(\u_top_module.addr[1] ),
    .B(\u_top_module.addr[0] ));
 sg13g2_nor2_1 _1207_ (.A(_0005_),
    .B(_0204_),
    .Y(_0205_));
 sg13g2_a22oi_1 _1208_ (.Y(_0206_),
    .B1(net937),
    .B2(\u_top_module.u_memory.memory[7][0] ),
    .A2(net929),
    .A1(\u_top_module.u_memory.memory[1][0] ));
 sg13g2_nand2b_1 _1209_ (.Y(_0207_),
    .B(\u_top_module.addr[1] ),
    .A_N(\u_top_module.addr[0] ));
 sg13g2_nor2_1 _1210_ (.A(\u_top_module.addr[2] ),
    .B(_0207_),
    .Y(_0208_));
 sg13g2_nand2_1 _1211_ (.Y(_0209_),
    .A(\u_top_module.u_memory.memory[2][0] ),
    .B(net935));
 sg13g2_nor2_1 _1212_ (.A(\u_top_module.addr[2] ),
    .B(_0204_),
    .Y(_0210_));
 sg13g2_nor2_1 _1213_ (.A(_0005_),
    .B(_0207_),
    .Y(_0211_));
 sg13g2_nor2_1 _1214_ (.A(_0005_),
    .B(_0193_),
    .Y(_0212_));
 sg13g2_a22oi_1 _1215_ (.Y(_0213_),
    .B1(net931),
    .B2(\u_top_module.u_memory.memory[6][0] ),
    .A2(_0194_),
    .A1(\u_top_module.u_memory.memory[4][0] ));
 sg13g2_nand3_1 _1216_ (.B(_0209_),
    .C(_0213_),
    .A(_0202_),
    .Y(_0214_));
 sg13g2_a221oi_1 _1217_ (.B2(\u_top_module.u_memory.memory[5][0] ),
    .C1(_0214_),
    .B1(net927),
    .A1(\u_top_module.u_memory.memory[3][0] ),
    .Y(_0215_),
    .A2(net933));
 sg13g2_nor3_1 _1218_ (.A(\u_top_module.addr[1] ),
    .B(\u_top_module.addr[0] ),
    .C(_0005_),
    .Y(_0216_));
 sg13g2_a22oi_1 _1219_ (.Y(_0158_),
    .B1(_0206_),
    .B2(_0215_),
    .A2(_0201_),
    .A1(_0174_));
 sg13g2_a22oi_1 _1220_ (.Y(_0217_),
    .B1(net930),
    .B2(\u_top_module.u_memory.memory[6][1] ),
    .A2(_0201_),
    .A1(\u_top_module.u_memory.memory[0][1] ));
 sg13g2_a22oi_1 _1221_ (.Y(_0218_),
    .B1(net936),
    .B2(\u_top_module.u_memory.memory[7][1] ),
    .A2(net928),
    .A1(\u_top_module.u_memory.memory[1][1] ));
 sg13g2_a22oi_1 _1222_ (.Y(_0219_),
    .B1(net926),
    .B2(\u_top_module.u_memory.memory[5][1] ),
    .A2(net932),
    .A1(\u_top_module.u_memory.memory[3][1] ));
 sg13g2_a22oi_1 _1223_ (.Y(_0220_),
    .B1(net943),
    .B2(\u_top_module.u_memory.memory[4][1] ),
    .A2(net934),
    .A1(\u_top_module.u_memory.memory[2][1] ));
 sg13g2_and2_1 _1224_ (.A(_0219_),
    .B(_0220_),
    .X(_0221_));
 sg13g2_nand3_1 _1225_ (.B(_0218_),
    .C(_0221_),
    .A(_0217_),
    .Y(_0159_));
 sg13g2_a22oi_1 _1226_ (.Y(_0222_),
    .B1(net944),
    .B2(\u_top_module.u_memory.memory[4][2] ),
    .A2(net933),
    .A1(\u_top_module.u_memory.memory[3][2] ));
 sg13g2_a22oi_1 _1227_ (.Y(_0223_),
    .B1(net931),
    .B2(\u_top_module.u_memory.memory[6][2] ),
    .A2(net937),
    .A1(\u_top_module.u_memory.memory[7][2] ));
 sg13g2_a22oi_1 _1228_ (.Y(_0224_),
    .B1(net935),
    .B2(\u_top_module.u_memory.memory[2][2] ),
    .A2(net929),
    .A1(\u_top_module.u_memory.memory[1][2] ));
 sg13g2_a22oi_1 _1229_ (.Y(_0225_),
    .B1(net927),
    .B2(\u_top_module.u_memory.memory[5][2] ),
    .A2(_0201_),
    .A1(\u_top_module.u_memory.memory[0][2] ));
 sg13g2_nand4_1 _1230_ (.B(_0223_),
    .C(_0224_),
    .A(_0222_),
    .Y(_0160_),
    .D(_0225_));
 sg13g2_a22oi_1 _1231_ (.Y(_0226_),
    .B1(net937),
    .B2(\u_top_module.u_memory.memory[7][3] ),
    .A2(_0201_),
    .A1(\u_top_module.u_memory.memory[0][3] ));
 sg13g2_a22oi_1 _1232_ (.Y(_0227_),
    .B1(net927),
    .B2(\u_top_module.u_memory.memory[5][3] ),
    .A2(net935),
    .A1(\u_top_module.u_memory.memory[2][3] ));
 sg13g2_a22oi_1 _1233_ (.Y(_0228_),
    .B1(net944),
    .B2(\u_top_module.u_memory.memory[4][3] ),
    .A2(_0211_),
    .A1(\u_top_module.u_memory.memory[6][3] ));
 sg13g2_a22oi_1 _1234_ (.Y(_0229_),
    .B1(net933),
    .B2(\u_top_module.u_memory.memory[3][3] ),
    .A2(net929),
    .A1(\u_top_module.u_memory.memory[1][3] ));
 sg13g2_and2_1 _1235_ (.A(_0228_),
    .B(_0229_),
    .X(_0230_));
 sg13g2_nand3_1 _1236_ (.B(_0227_),
    .C(_0230_),
    .A(_0226_),
    .Y(_0161_));
 sg13g2_a22oi_1 _1237_ (.Y(_0231_),
    .B1(net934),
    .B2(\u_top_module.u_memory.memory[2][4] ),
    .A2(net936),
    .A1(\u_top_module.u_memory.memory[7][4] ));
 sg13g2_a22oi_1 _1238_ (.Y(_0232_),
    .B1(net930),
    .B2(\u_top_module.u_memory.memory[6][4] ),
    .A2(net928),
    .A1(\u_top_module.u_memory.memory[1][4] ));
 sg13g2_a22oi_1 _1239_ (.Y(_0233_),
    .B1(net943),
    .B2(\u_top_module.u_memory.memory[4][4] ),
    .A2(net932),
    .A1(\u_top_module.u_memory.memory[3][4] ));
 sg13g2_a22oi_1 _1240_ (.Y(_0234_),
    .B1(net926),
    .B2(\u_top_module.u_memory.memory[5][4] ),
    .A2(_0201_),
    .A1(\u_top_module.u_memory.memory[0][4] ));
 sg13g2_nand4_1 _1241_ (.B(_0232_),
    .C(_0233_),
    .A(_0231_),
    .Y(_0162_),
    .D(_0234_));
 sg13g2_a22oi_1 _1242_ (.Y(_0235_),
    .B1(net943),
    .B2(\u_top_module.u_memory.memory[4][5] ),
    .A2(net930),
    .A1(\u_top_module.u_memory.memory[6][5] ));
 sg13g2_a22oi_1 _1243_ (.Y(_0236_),
    .B1(net926),
    .B2(\u_top_module.u_memory.memory[5][5] ),
    .A2(net928),
    .A1(\u_top_module.u_memory.memory[1][5] ));
 sg13g2_a22oi_1 _1244_ (.Y(_0237_),
    .B1(net934),
    .B2(\u_top_module.u_memory.memory[2][5] ),
    .A2(net936),
    .A1(\u_top_module.u_memory.memory[7][5] ));
 sg13g2_a21oi_1 _1245_ (.A1(\u_top_module.u_memory.memory[3][5] ),
    .A2(net932),
    .Y(_0238_),
    .B1(_0201_));
 sg13g2_nand4_1 _1246_ (.B(_0236_),
    .C(_0237_),
    .A(_0235_),
    .Y(_0239_),
    .D(_0238_));
 sg13g2_o21ai_1 _1247_ (.B1(_0239_),
    .Y(_0240_),
    .A1(\u_top_module.u_memory.memory[0][5] ),
    .A2(_0202_));
 sg13g2_inv_1 _1248_ (.Y(_0163_),
    .A(_0240_));
 sg13g2_a22oi_1 _1249_ (.Y(_0241_),
    .B1(net943),
    .B2(\u_top_module.u_memory.memory[4][6] ),
    .A2(net926),
    .A1(\u_top_module.u_memory.memory[5][6] ));
 sg13g2_a22oi_1 _1250_ (.Y(_0242_),
    .B1(net930),
    .B2(\u_top_module.u_memory.memory[6][6] ),
    .A2(net936),
    .A1(\u_top_module.u_memory.memory[7][6] ));
 sg13g2_a22oi_1 _1251_ (.Y(_0243_),
    .B1(net932),
    .B2(\u_top_module.u_memory.memory[3][6] ),
    .A2(net934),
    .A1(\u_top_module.u_memory.memory[2][6] ));
 sg13g2_a21oi_1 _1252_ (.A1(\u_top_module.u_memory.memory[1][6] ),
    .A2(net928),
    .Y(_0244_),
    .B1(_0201_));
 sg13g2_nand4_1 _1253_ (.B(_0242_),
    .C(_0243_),
    .A(_0241_),
    .Y(_0245_),
    .D(_0244_));
 sg13g2_o21ai_1 _1254_ (.B1(_0245_),
    .Y(_0246_),
    .A1(\u_top_module.u_memory.memory[0][6] ),
    .A2(_0202_));
 sg13g2_inv_1 _1255_ (.Y(_0164_),
    .A(_0246_));
 sg13g2_a22oi_1 _1256_ (.Y(_0247_),
    .B1(net937),
    .B2(\u_top_module.u_memory.memory[7][7] ),
    .A2(_0201_),
    .A1(\u_top_module.u_memory.memory[0][7] ));
 sg13g2_a22oi_1 _1257_ (.Y(_0248_),
    .B1(net931),
    .B2(\u_top_module.u_memory.memory[6][7] ),
    .A2(net935),
    .A1(\u_top_module.u_memory.memory[2][7] ));
 sg13g2_a22oi_1 _1258_ (.Y(_0249_),
    .B1(net933),
    .B2(\u_top_module.u_memory.memory[3][7] ),
    .A2(net929),
    .A1(\u_top_module.u_memory.memory[1][7] ));
 sg13g2_a22oi_1 _1259_ (.Y(_0250_),
    .B1(net944),
    .B2(\u_top_module.u_memory.memory[4][7] ),
    .A2(net927),
    .A1(\u_top_module.u_memory.memory[5][7] ));
 sg13g2_and2_1 _1260_ (.A(_0249_),
    .B(_0250_),
    .X(_0251_));
 sg13g2_nand3_1 _1261_ (.B(_0248_),
    .C(_0251_),
    .A(_0247_),
    .Y(_0165_));
 sg13g2_nor2_1 _1262_ (.A(\u_top_module.u_buffer.corr_neg[7] ),
    .B(_0175_),
    .Y(_0252_));
 sg13g2_nand2b_1 _1263_ (.Y(_0253_),
    .B(\u_top_module.u_buffer.corr_pos[7] ),
    .A_N(\u_top_module.u_buffer.corr_neg[7] ));
 sg13g2_a22oi_1 _1264_ (.Y(_0254_),
    .B1(_0176_),
    .B2(\u_top_module.u_buffer.corr_neg[6] ),
    .A2(_0175_),
    .A1(\u_top_module.u_buffer.corr_neg[7] ));
 sg13g2_a22oi_1 _1265_ (.Y(_0255_),
    .B1(\u_top_module.u_buffer.corr_pos[5] ),
    .B2(_0179_),
    .A2(_0177_),
    .A1(\u_top_module.u_buffer.corr_pos[6] ));
 sg13g2_nor2_1 _1266_ (.A(_0180_),
    .B(\u_top_module.u_buffer.corr_pos[4] ),
    .Y(_0256_));
 sg13g2_a21oi_1 _1267_ (.A1(_0178_),
    .A2(net821),
    .Y(_0257_),
    .B1(_0256_));
 sg13g2_nand2_1 _1268_ (.Y(_0258_),
    .A(_0180_),
    .B(\u_top_module.u_buffer.corr_pos[4] ));
 sg13g2_nor2_1 _1269_ (.A(_0182_),
    .B(\u_top_module.u_buffer.corr_neg[3] ),
    .Y(_0259_));
 sg13g2_a21oi_1 _1270_ (.A1(\u_top_module.u_buffer.corr_pos[2] ),
    .A2(_0185_),
    .Y(_0260_),
    .B1(_0259_));
 sg13g2_a22oi_1 _1271_ (.Y(_0261_),
    .B1(_0188_),
    .B2(\u_top_module.u_buffer.corr_pos[0] ),
    .A2(_0187_),
    .A1(\u_top_module.u_buffer.corr_pos[1] ));
 sg13g2_nor2_1 _1272_ (.A(\u_top_module.u_buffer.corr_pos[1] ),
    .B(_0187_),
    .Y(_0262_));
 sg13g2_o21ai_1 _1273_ (.B1(_0260_),
    .Y(_0263_),
    .A1(_0261_),
    .A2(_0262_));
 sg13g2_a22oi_1 _1274_ (.Y(_0264_),
    .B1(_0184_),
    .B2(\u_top_module.u_buffer.corr_neg[2] ),
    .A2(\u_top_module.u_buffer.corr_neg[3] ),
    .A1(_0182_));
 sg13g2_o21ai_1 _1275_ (.B1(_0263_),
    .Y(_0265_),
    .A1(_0259_),
    .A2(_0264_));
 sg13g2_a221oi_1 _1276_ (.B2(_0265_),
    .C1(_0256_),
    .B1(_0258_),
    .A1(_0178_),
    .Y(_0266_),
    .A2(net821));
 sg13g2_nand2b_1 _1277_ (.Y(_0267_),
    .B(_0255_),
    .A_N(_0266_));
 sg13g2_a21o_1 _1278_ (.A2(_0267_),
    .A1(_0254_),
    .B1(_0252_),
    .X(_0000_));
 sg13g2_xor2_1 _1279_ (.B(\u_top_module.u_buffer.shift_reg_1[255] ),
    .A(\u_top_module.u_buffer.shift_reg_2[255] ),
    .X(_0268_));
 sg13g2_xnor2_1 _1280_ (.Y(_0269_),
    .A(\u_top_module.dec_data_2 ),
    .B(\u_top_module.dec_data_1 ));
 sg13g2_xor2_1 _1281_ (.B(_0269_),
    .A(_0268_),
    .X(_0270_));
 sg13g2_xor2_1 _1282_ (.B(_0270_),
    .A(_0014_),
    .X(_0018_));
 sg13g2_a21oi_2 _1283_ (.B1(uo_out[1]),
    .Y(_0271_),
    .A2(_0269_),
    .A1(_0268_));
 sg13g2_and3_1 _1284_ (.X(_0272_),
    .A(uo_out[1]),
    .B(_0268_),
    .C(_0269_));
 sg13g2_or2_1 _1285_ (.X(_0273_),
    .B(_0272_),
    .A(_0271_));
 sg13g2_nor4_2 _1286_ (.A(_0014_),
    .B(_0270_),
    .C(_0271_),
    .Y(_0274_),
    .D(_0272_));
 sg13g2_o21ai_1 _1287_ (.B1(_0273_),
    .Y(_0275_),
    .A1(_0014_),
    .A2(_0270_));
 sg13g2_nor2b_1 _1288_ (.A(_0274_),
    .B_N(_0275_),
    .Y(_0019_));
 sg13g2_nand2b_1 _1289_ (.Y(_0276_),
    .B(uo_out[1]),
    .A_N(uo_out[2]));
 sg13g2_xnor2_1 _1290_ (.Y(_0277_),
    .A(uo_out[1]),
    .B(uo_out[2]));
 sg13g2_o21ai_1 _1291_ (.B1(_0277_),
    .Y(_0278_),
    .A1(_0271_),
    .A2(_0274_));
 sg13g2_or3_1 _1292_ (.A(_0271_),
    .B(_0274_),
    .C(_0277_),
    .X(_0279_));
 sg13g2_and2_1 _1293_ (.A(_0278_),
    .B(_0279_),
    .X(_0020_));
 sg13g2_xor2_1 _1294_ (.B(uo_out[3]),
    .A(uo_out[2]),
    .X(_0280_));
 sg13g2_a21oi_1 _1295_ (.A1(_0276_),
    .A2(_0278_),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_nand3_1 _1296_ (.B(_0278_),
    .C(_0280_),
    .A(_0276_),
    .Y(_0282_));
 sg13g2_nor2b_1 _1297_ (.A(_0281_),
    .B_N(_0282_),
    .Y(_0021_));
 sg13g2_a21oi_2 _1298_ (.B1(_0281_),
    .Y(_0283_),
    .A2(_0189_),
    .A1(uo_out[2]));
 sg13g2_nand2_1 _1299_ (.Y(_0284_),
    .A(_0189_),
    .B(uo_out[4]));
 sg13g2_nand2b_1 _1300_ (.Y(_0285_),
    .B(uo_out[3]),
    .A_N(uo_out[4]));
 sg13g2_and2_1 _1301_ (.A(_0284_),
    .B(_0285_),
    .X(_0286_));
 sg13g2_nand2b_1 _1302_ (.Y(_0287_),
    .B(_0286_),
    .A_N(_0283_));
 sg13g2_xnor2_1 _1303_ (.Y(_0022_),
    .A(_0283_),
    .B(_0286_));
 sg13g2_xor2_1 _1304_ (.B(uo_out[5]),
    .A(uo_out[4]),
    .X(_0288_));
 sg13g2_nand2_1 _1305_ (.Y(_0289_),
    .A(_0285_),
    .B(_0287_));
 sg13g2_xnor2_1 _1306_ (.Y(_0023_),
    .A(_0288_),
    .B(_0289_));
 sg13g2_nor2_1 _1307_ (.A(_0190_),
    .B(uo_out[6]),
    .Y(_0290_));
 sg13g2_nand2_1 _1308_ (.Y(_0291_),
    .A(_0190_),
    .B(uo_out[6]));
 sg13g2_nand2b_1 _1309_ (.Y(_0292_),
    .B(_0291_),
    .A_N(_0290_));
 sg13g2_nand3b_1 _1310_ (.B(_0285_),
    .C(_0284_),
    .Y(_0293_),
    .A_N(_0288_));
 sg13g2_o21ai_1 _1311_ (.B1(_0190_),
    .Y(_0294_),
    .A1(uo_out[3]),
    .A2(uo_out[4]));
 sg13g2_o21ai_1 _1312_ (.B1(_0294_),
    .Y(_0295_),
    .A1(_0283_),
    .A2(_0293_));
 sg13g2_xnor2_1 _1313_ (.Y(_0024_),
    .A(_0292_),
    .B(_0295_));
 sg13g2_a21oi_1 _1314_ (.A1(_0291_),
    .A2(_0295_),
    .Y(_0296_),
    .B1(_0290_));
 sg13g2_xnor2_1 _1315_ (.Y(_0297_),
    .A(uo_out[6]),
    .B(uo_out[7]));
 sg13g2_xnor2_1 _1316_ (.Y(_0025_),
    .A(_0296_),
    .B(_0297_));
 sg13g2_nand4_1 _1317_ (.B(_0260_),
    .C(_0261_),
    .A(_0257_),
    .Y(_0298_),
    .D(_0264_));
 sg13g2_nor2_1 _1318_ (.A(_0188_),
    .B(\u_top_module.u_buffer.corr_pos[0] ),
    .Y(_0299_));
 sg13g2_nand4_1 _1319_ (.B(_0254_),
    .C(_0255_),
    .A(_0253_),
    .Y(_0300_),
    .D(_0258_));
 sg13g2_nor4_2 _1320_ (.A(_0262_),
    .B(_0298_),
    .C(_0299_),
    .Y(_0301_),
    .D(_0300_));
 sg13g2_nor2_1 _1321_ (.A(_0000_),
    .B(_0301_),
    .Y(_0003_));
 sg13g2_or2_1 _1322_ (.X(_0302_),
    .B(\u_top_module.decimation_ratio[1] ),
    .A(\u_top_module.decimation_ratio[0] ));
 sg13g2_or3_2 _1323_ (.A(\u_top_module.decimation_ratio[0] ),
    .B(\u_top_module.decimation_ratio[1] ),
    .C(\u_top_module.decimation_ratio[2] ),
    .X(_0303_));
 sg13g2_nor4_2 _1324_ (.A(\u_top_module.decimation_ratio[0] ),
    .B(\u_top_module.decimation_ratio[1] ),
    .C(\u_top_module.decimation_ratio[3] ),
    .Y(_0304_),
    .D(\u_top_module.decimation_ratio[2] ));
 sg13g2_nor2b_1 _1325_ (.A(\u_top_module.decimation_ratio[4] ),
    .B_N(_0304_),
    .Y(_0305_));
 sg13g2_nor4_1 _1326_ (.A(\u_top_module.decimation_ratio[3] ),
    .B(\u_top_module.decimation_ratio[5] ),
    .C(\u_top_module.decimation_ratio[4] ),
    .D(_0303_),
    .Y(_0306_));
 sg13g2_nor2b_1 _1327_ (.A(\u_top_module.decimation_ratio[6] ),
    .B_N(_0306_),
    .Y(_0307_));
 sg13g2_nor2b_2 _1328_ (.A(\u_top_module.decimation_ratio[7] ),
    .B_N(_0307_),
    .Y(_0308_));
 sg13g2_xnor2_1 _1329_ (.Y(_0309_),
    .A(\u_top_module.decimation_ratio[6] ),
    .B(_0306_));
 sg13g2_inv_1 _1330_ (.Y(_0310_),
    .A(_0309_));
 sg13g2_nor2_1 _1331_ (.A(_0007_),
    .B(_0310_),
    .Y(_0311_));
 sg13g2_nand2_1 _1332_ (.Y(_0312_),
    .A(\u_top_module.u_decimator_2.counter[0] ),
    .B(\u_top_module.u_decimator_2.counter[1] ));
 sg13g2_nor2b_1 _1333_ (.A(\u_top_module.decimation_ratio[0] ),
    .B_N(\u_top_module.u_decimator_2.counter[0] ),
    .Y(_0313_));
 sg13g2_nand2b_1 _1334_ (.Y(_0314_),
    .B(\u_top_module.decimation_ratio[1] ),
    .A_N(\u_top_module.u_decimator_2.counter[1] ));
 sg13g2_o21ai_1 _1335_ (.B1(_0302_),
    .Y(_0315_),
    .A1(_0313_),
    .A2(_0314_));
 sg13g2_o21ai_1 _1336_ (.B1(\u_top_module.decimation_ratio[2] ),
    .Y(_0316_),
    .A1(\u_top_module.decimation_ratio[0] ),
    .A2(\u_top_module.decimation_ratio[1] ));
 sg13g2_nand3_1 _1337_ (.B(_0303_),
    .C(_0316_),
    .A(_0006_),
    .Y(_0317_));
 sg13g2_a21o_1 _1338_ (.A2(_0316_),
    .A1(_0303_),
    .B1(_0006_),
    .X(_0318_));
 sg13g2_a22oi_1 _1339_ (.Y(_0319_),
    .B1(_0317_),
    .B2(_0318_),
    .A2(_0315_),
    .A1(_0312_));
 sg13g2_xnor2_1 _1340_ (.Y(_0320_),
    .A(\u_top_module.decimation_ratio[3] ),
    .B(_0303_));
 sg13g2_nand3_1 _1341_ (.B(_0303_),
    .C(_0316_),
    .A(\u_top_module.u_decimator_2.counter[2] ),
    .Y(_0321_));
 sg13g2_o21ai_1 _1342_ (.B1(_0321_),
    .Y(_0322_),
    .A1(_0167_),
    .A2(_0320_));
 sg13g2_xnor2_1 _1343_ (.Y(_0323_),
    .A(\u_top_module.decimation_ratio[4] ),
    .B(_0304_));
 sg13g2_xor2_1 _1344_ (.B(_0304_),
    .A(\u_top_module.decimation_ratio[4] ),
    .X(_0324_));
 sg13g2_a22oi_1 _1345_ (.Y(_0325_),
    .B1(_0324_),
    .B2(_0168_),
    .A2(_0320_),
    .A1(_0167_));
 sg13g2_o21ai_1 _1346_ (.B1(_0325_),
    .Y(_0326_),
    .A1(_0319_),
    .A2(_0322_));
 sg13g2_xnor2_1 _1347_ (.Y(_0327_),
    .A(\u_top_module.decimation_ratio[5] ),
    .B(_0305_));
 sg13g2_a22oi_1 _1348_ (.Y(_0328_),
    .B1(_0327_),
    .B2(\u_top_module.u_decimator_2.counter[5] ),
    .A2(_0323_),
    .A1(\u_top_module.u_decimator_2.counter[4] ));
 sg13g2_nor2_1 _1349_ (.A(\u_top_module.u_decimator_2.counter[5] ),
    .B(_0327_),
    .Y(_0329_));
 sg13g2_a221oi_1 _1350_ (.B2(_0328_),
    .C1(_0329_),
    .B1(_0326_),
    .A1(_0007_),
    .Y(_0330_),
    .A2(_0310_));
 sg13g2_or2_1 _1351_ (.X(_0331_),
    .B(_0330_),
    .A(_0311_));
 sg13g2_xnor2_1 _1352_ (.Y(_0332_),
    .A(\u_top_module.decimation_ratio[7] ),
    .B(_0307_));
 sg13g2_xor2_1 _1353_ (.B(_0332_),
    .A(\u_top_module.u_decimator_2.counter[7] ),
    .X(_0333_));
 sg13g2_a221oi_1 _1354_ (.B2(_0331_),
    .C1(net919),
    .B1(_0333_),
    .A1(_0169_),
    .Y(_0334_),
    .A2(_0332_));
 sg13g2_nor2_2 _1355_ (.A(_0308_),
    .B(_0334_),
    .Y(_0335_));
 sg13g2_mux2_1 _1356_ (.A0(\u_top_module.dec_data_2 ),
    .A1(net4),
    .S(_0335_),
    .X(_0027_));
 sg13g2_nor2_1 _1357_ (.A(\u_top_module.u_decimator_1.counter[5] ),
    .B(_0327_),
    .Y(_0336_));
 sg13g2_nand2_2 _1358_ (.Y(_0337_),
    .A(\u_top_module.u_decimator_1.counter[1] ),
    .B(\u_top_module.u_decimator_1.counter[0] ));
 sg13g2_nor2b_1 _1359_ (.A(\u_top_module.decimation_ratio[0] ),
    .B_N(\u_top_module.u_decimator_1.counter[0] ),
    .Y(_0338_));
 sg13g2_nand2b_1 _1360_ (.Y(_0339_),
    .B(\u_top_module.decimation_ratio[1] ),
    .A_N(\u_top_module.u_decimator_1.counter[1] ));
 sg13g2_o21ai_1 _1361_ (.B1(_0302_),
    .Y(_0340_),
    .A1(_0338_),
    .A2(_0339_));
 sg13g2_nand3_1 _1362_ (.B(_0303_),
    .C(_0316_),
    .A(_0010_),
    .Y(_0341_));
 sg13g2_a21o_1 _1363_ (.A2(_0316_),
    .A1(_0303_),
    .B1(_0010_),
    .X(_0342_));
 sg13g2_a22oi_1 _1364_ (.Y(_0343_),
    .B1(_0341_),
    .B2(_0342_),
    .A2(_0340_),
    .A1(_0337_));
 sg13g2_nand3_1 _1365_ (.B(_0303_),
    .C(_0316_),
    .A(\u_top_module.u_decimator_1.counter[2] ),
    .Y(_0344_));
 sg13g2_o21ai_1 _1366_ (.B1(_0344_),
    .Y(_0345_),
    .A1(_0171_),
    .A2(_0320_));
 sg13g2_a22oi_1 _1367_ (.Y(_0346_),
    .B1(_0324_),
    .B2(_0170_),
    .A2(_0320_),
    .A1(_0171_));
 sg13g2_o21ai_1 _1368_ (.B1(_0346_),
    .Y(_0347_),
    .A1(_0343_),
    .A2(_0345_));
 sg13g2_a22oi_1 _1369_ (.Y(_0348_),
    .B1(_0327_),
    .B2(\u_top_module.u_decimator_1.counter[5] ),
    .A2(_0323_),
    .A1(\u_top_module.u_decimator_1.counter[4] ));
 sg13g2_xnor2_1 _1370_ (.Y(_0349_),
    .A(\u_top_module.u_decimator_1.counter[7] ),
    .B(_0332_));
 sg13g2_a21oi_1 _1371_ (.A1(_0347_),
    .A2(_0348_),
    .Y(_0350_),
    .B1(_0336_));
 sg13g2_xor2_1 _1372_ (.B(_0309_),
    .A(_0009_),
    .X(_0351_));
 sg13g2_nor2_1 _1373_ (.A(_0349_),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_nor3_1 _1374_ (.A(_0009_),
    .B(_0310_),
    .C(_0349_),
    .Y(_0353_));
 sg13g2_a221oi_1 _1375_ (.B2(_0352_),
    .C1(_0353_),
    .B1(_0350_),
    .A1(_0173_),
    .Y(_0354_),
    .A2(_0332_));
 sg13g2_a21oi_1 _1376_ (.A1(_0199_),
    .A2(_0354_),
    .Y(_0355_),
    .B1(\u_top_module.u_decimator_1.counter[0] ));
 sg13g2_a21oi_1 _1377_ (.A1(\u_top_module.u_decimator_1.counter[0] ),
    .A2(_0199_),
    .Y(_0028_),
    .B1(_0355_));
 sg13g2_nor3_2 _1378_ (.A(net919),
    .B(_0308_),
    .C(_0354_),
    .Y(_0356_));
 sg13g2_nor2_1 _1379_ (.A(net919),
    .B(_0337_),
    .Y(_0357_));
 sg13g2_a21oi_1 _1380_ (.A1(\u_top_module.u_decimator_1.counter[0] ),
    .A2(_0199_),
    .Y(_0358_),
    .B1(\u_top_module.u_decimator_1.counter[1] ));
 sg13g2_nor3_1 _1381_ (.A(_0356_),
    .B(_0357_),
    .C(_0358_),
    .Y(_0029_));
 sg13g2_nand2_1 _1382_ (.Y(_0359_),
    .A(\u_top_module.u_decimator_1.counter[2] ),
    .B(net919));
 sg13g2_a21oi_2 _1383_ (.B1(_0308_),
    .Y(_0360_),
    .A2(_0354_),
    .A1(_0199_));
 sg13g2_xnor2_1 _1384_ (.Y(_0361_),
    .A(_0010_),
    .B(_0337_));
 sg13g2_o21ai_1 _1385_ (.B1(_0359_),
    .Y(_0030_),
    .A1(_0360_),
    .A2(_0361_));
 sg13g2_nor4_1 _1386_ (.A(_0171_),
    .B(_0172_),
    .C(net919),
    .D(_0337_),
    .Y(_0362_));
 sg13g2_a21oi_1 _1387_ (.A1(\u_top_module.u_decimator_1.counter[2] ),
    .A2(_0357_),
    .Y(_0363_),
    .B1(\u_top_module.u_decimator_1.counter[3] ));
 sg13g2_nor3_1 _1388_ (.A(_0356_),
    .B(_0362_),
    .C(_0363_),
    .Y(_0031_));
 sg13g2_nand2_1 _1389_ (.Y(_0364_),
    .A(\u_top_module.u_decimator_1.counter[4] ),
    .B(net918));
 sg13g2_nor3_2 _1390_ (.A(_0171_),
    .B(_0172_),
    .C(_0337_),
    .Y(_0365_));
 sg13g2_xor2_1 _1391_ (.B(_0365_),
    .A(_0013_),
    .X(_0366_));
 sg13g2_o21ai_1 _1392_ (.B1(_0364_),
    .Y(_0032_),
    .A1(_0360_),
    .A2(_0366_));
 sg13g2_nand3_1 _1393_ (.B(_0199_),
    .C(_0365_),
    .A(\u_top_module.u_decimator_1.counter[4] ),
    .Y(_0367_));
 sg13g2_xor2_1 _1394_ (.B(_0367_),
    .A(\u_top_module.u_decimator_1.counter[5] ),
    .X(_0368_));
 sg13g2_nor2_1 _1395_ (.A(_0356_),
    .B(_0368_),
    .Y(_0033_));
 sg13g2_nand2_1 _1396_ (.Y(_0369_),
    .A(\u_top_module.u_decimator_1.counter[6] ),
    .B(net918));
 sg13g2_nand3_1 _1397_ (.B(\u_top_module.u_decimator_1.counter[4] ),
    .C(_0365_),
    .A(\u_top_module.u_decimator_1.counter[5] ),
    .Y(_0370_));
 sg13g2_nor2_1 _1398_ (.A(_0009_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_xnor2_1 _1399_ (.Y(_0372_),
    .A(_0009_),
    .B(_0370_));
 sg13g2_o21ai_1 _1400_ (.B1(_0369_),
    .Y(_0034_),
    .A1(_0360_),
    .A2(_0372_));
 sg13g2_nand2_1 _1401_ (.Y(_0373_),
    .A(\u_top_module.u_decimator_1.counter[7] ),
    .B(net918));
 sg13g2_xnor2_1 _1402_ (.Y(_0374_),
    .A(_0173_),
    .B(_0371_));
 sg13g2_o21ai_1 _1403_ (.B1(_0373_),
    .Y(_0035_),
    .A1(_0360_),
    .A2(_0374_));
 sg13g2_mux2_1 _1404_ (.A0(\u_top_module.dec_clk ),
    .A1(_0004_),
    .S(_0356_),
    .X(_0036_));
 sg13g2_or4_1 _1405_ (.A(\u_top_module.filter_length[6] ),
    .B(\u_top_module.filter_length[5] ),
    .C(\u_top_module.filter_length[4] ),
    .D(\u_top_module.filter_length[3] ),
    .X(_0375_));
 sg13g2_nor4_2 _1406_ (.A(\u_top_module.filter_length[2] ),
    .B(\u_top_module.filter_length[1] ),
    .C(\u_top_module.filter_length[7] ),
    .Y(_0376_),
    .D(_0375_));
 sg13g2_xnor2_1 _1407_ (.Y(_0377_),
    .A(\u_top_module.u_buffer.shift_reg_2[255] ),
    .B(\u_top_module.u_buffer.shift_reg_1[254] ));
 sg13g2_xor2_1 _1408_ (.B(\u_top_module.u_buffer.shift_reg_2[0] ),
    .A(\u_top_module.dec_data_1 ),
    .X(_0378_));
 sg13g2_nor2_1 _1409_ (.A(_0377_),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_xnor2_1 _1410_ (.Y(_0380_),
    .A(_0377_),
    .B(_0378_));
 sg13g2_nor2b_1 _1411_ (.A(_0015_),
    .B_N(_0380_),
    .Y(_0381_));
 sg13g2_xor2_1 _1412_ (.B(_0380_),
    .A(_0015_),
    .X(_0382_));
 sg13g2_nand2_1 _1413_ (.Y(_0383_),
    .A(\u_top_module.u_buffer.corr_pos[0] ),
    .B(net923));
 sg13g2_o21ai_1 _1414_ (.B1(_0383_),
    .Y(_0037_),
    .A1(net923),
    .A2(_0382_));
 sg13g2_nor2_1 _1415_ (.A(\u_top_module.u_buffer.corr_pos[1] ),
    .B(_0379_),
    .Y(_0384_));
 sg13g2_nand2_1 _1416_ (.Y(_0385_),
    .A(\u_top_module.u_buffer.corr_pos[1] ),
    .B(_0379_));
 sg13g2_nand2b_1 _1417_ (.Y(_0386_),
    .B(_0385_),
    .A_N(_0384_));
 sg13g2_xnor2_1 _1418_ (.Y(_0387_),
    .A(_0381_),
    .B(_0386_));
 sg13g2_nor2_1 _1419_ (.A(net923),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_a21oi_1 _1420_ (.A1(_0186_),
    .A2(net923),
    .Y(_0038_),
    .B1(_0388_));
 sg13g2_nand2_1 _1421_ (.Y(_0389_),
    .A(\u_top_module.u_buffer.corr_pos[2] ),
    .B(net923));
 sg13g2_a21o_1 _1422_ (.A2(_0385_),
    .A1(_0381_),
    .B1(_0384_),
    .X(_0390_));
 sg13g2_xor2_1 _1423_ (.B(\u_top_module.u_buffer.corr_pos[1] ),
    .A(\u_top_module.u_buffer.corr_pos[2] ),
    .X(_0391_));
 sg13g2_xnor2_1 _1424_ (.Y(_0392_),
    .A(\u_top_module.u_buffer.corr_pos[2] ),
    .B(\u_top_module.u_buffer.corr_pos[1] ));
 sg13g2_xnor2_1 _1425_ (.Y(_0393_),
    .A(_0390_),
    .B(_0392_));
 sg13g2_o21ai_1 _1426_ (.B1(_0389_),
    .Y(_0039_),
    .A1(net921),
    .A2(_0393_));
 sg13g2_nor2_1 _1427_ (.A(\u_top_module.u_buffer.corr_pos[2] ),
    .B(_0186_),
    .Y(_0394_));
 sg13g2_a21oi_1 _1428_ (.A1(_0390_),
    .A2(_0392_),
    .Y(_0395_),
    .B1(_0394_));
 sg13g2_xor2_1 _1429_ (.B(\u_top_module.u_buffer.corr_pos[2] ),
    .A(\u_top_module.u_buffer.corr_pos[3] ),
    .X(_0396_));
 sg13g2_xor2_1 _1430_ (.B(_0396_),
    .A(_0395_),
    .X(_0397_));
 sg13g2_nor2_1 _1431_ (.A(net921),
    .B(_0397_),
    .Y(_0398_));
 sg13g2_a21oi_1 _1432_ (.A1(_0182_),
    .A2(net921),
    .Y(_0040_),
    .B1(_0398_));
 sg13g2_nand2_1 _1433_ (.Y(_0399_),
    .A(\u_top_module.u_buffer.corr_pos[4] ),
    .B(net921));
 sg13g2_nor2_1 _1434_ (.A(_0391_),
    .B(_0396_),
    .Y(_0400_));
 sg13g2_a21oi_1 _1435_ (.A1(_0184_),
    .A2(_0186_),
    .Y(_0401_),
    .B1(\u_top_module.u_buffer.corr_pos[3] ));
 sg13g2_a21o_1 _1436_ (.A2(_0400_),
    .A1(_0390_),
    .B1(_0401_),
    .X(_0402_));
 sg13g2_nor2_1 _1437_ (.A(\u_top_module.u_buffer.corr_pos[4] ),
    .B(_0182_),
    .Y(_0403_));
 sg13g2_xnor2_1 _1438_ (.Y(_0404_),
    .A(\u_top_module.u_buffer.corr_pos[4] ),
    .B(\u_top_module.u_buffer.corr_pos[3] ));
 sg13g2_inv_1 _1439_ (.Y(_0405_),
    .A(_0404_));
 sg13g2_xnor2_1 _1440_ (.Y(_0406_),
    .A(_0402_),
    .B(_0404_));
 sg13g2_o21ai_1 _1441_ (.B1(_0399_),
    .Y(_0041_),
    .A1(net921),
    .A2(_0406_));
 sg13g2_xor2_1 _1442_ (.B(\u_top_module.u_buffer.corr_pos[4] ),
    .A(\u_top_module.u_buffer.corr_pos[5] ),
    .X(_0407_));
 sg13g2_a21oi_1 _1443_ (.A1(_0402_),
    .A2(_0404_),
    .Y(_0408_),
    .B1(_0403_));
 sg13g2_xnor2_1 _1444_ (.Y(_0409_),
    .A(_0407_),
    .B(_0408_));
 sg13g2_nand2_1 _1445_ (.Y(_0410_),
    .A(\u_top_module.u_buffer.corr_pos[5] ),
    .B(net921));
 sg13g2_o21ai_1 _1446_ (.B1(_0410_),
    .Y(_0042_),
    .A1(net921),
    .A2(_0409_));
 sg13g2_nand2_1 _1447_ (.Y(_0411_),
    .A(_0176_),
    .B(\u_top_module.u_buffer.corr_pos[5] ));
 sg13g2_xor2_1 _1448_ (.B(\u_top_module.u_buffer.corr_pos[5] ),
    .A(\u_top_module.u_buffer.corr_pos[6] ),
    .X(_0412_));
 sg13g2_nor2_1 _1449_ (.A(_0405_),
    .B(_0407_),
    .Y(_0413_));
 sg13g2_a21oi_1 _1450_ (.A1(_0181_),
    .A2(_0182_),
    .Y(_0414_),
    .B1(\u_top_module.u_buffer.corr_pos[5] ));
 sg13g2_a21oi_1 _1451_ (.A1(_0402_),
    .A2(_0413_),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_xor2_1 _1452_ (.B(_0415_),
    .A(_0412_),
    .X(_0416_));
 sg13g2_nor2_1 _1453_ (.A(net921),
    .B(_0416_),
    .Y(_0417_));
 sg13g2_a21oi_1 _1454_ (.A1(_0176_),
    .A2(net920),
    .Y(_0043_),
    .B1(_0417_));
 sg13g2_o21ai_1 _1455_ (.B1(_0411_),
    .Y(_0418_),
    .A1(_0412_),
    .A2(_0415_));
 sg13g2_xnor2_1 _1456_ (.Y(_0419_),
    .A(\u_top_module.u_buffer.corr_pos[7] ),
    .B(\u_top_module.u_buffer.corr_pos[6] ));
 sg13g2_xnor2_1 _1457_ (.Y(_0420_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_nand2_1 _1458_ (.Y(_0421_),
    .A(\u_top_module.u_buffer.corr_pos[7] ),
    .B(net920));
 sg13g2_o21ai_1 _1459_ (.B1(_0421_),
    .Y(_0044_),
    .A1(net920),
    .A2(_0420_));
 sg13g2_mux2_1 _1460_ (.A0(\u_top_module.dec_data_1 ),
    .A1(net3),
    .S(_0360_),
    .X(_0045_));
 sg13g2_nor2_1 _1461_ (.A(\u_top_module.u_decimator_2.counter[0] ),
    .B(_0334_),
    .Y(_0422_));
 sg13g2_a21oi_1 _1462_ (.A1(\u_top_module.u_decimator_2.counter[0] ),
    .A2(_0199_),
    .Y(_0046_),
    .B1(_0422_));
 sg13g2_nand2_1 _1463_ (.Y(_0423_),
    .A(\u_top_module.u_decimator_2.counter[1] ),
    .B(net919));
 sg13g2_xnor2_1 _1464_ (.Y(_0424_),
    .A(\u_top_module.u_decimator_2.counter[0] ),
    .B(\u_top_module.u_decimator_2.counter[1] ));
 sg13g2_o21ai_1 _1465_ (.B1(_0423_),
    .Y(_0047_),
    .A1(_0335_),
    .A2(_0424_));
 sg13g2_nand2_1 _1466_ (.Y(_0425_),
    .A(\u_top_module.u_decimator_2.counter[2] ),
    .B(net919));
 sg13g2_xnor2_1 _1467_ (.Y(_0426_),
    .A(_0006_),
    .B(_0312_));
 sg13g2_o21ai_1 _1468_ (.B1(_0425_),
    .Y(_0048_),
    .A1(_0335_),
    .A2(_0426_));
 sg13g2_nand2_1 _1469_ (.Y(_0427_),
    .A(\u_top_module.u_decimator_2.counter[3] ),
    .B(net918));
 sg13g2_nand3_1 _1470_ (.B(\u_top_module.u_decimator_2.counter[1] ),
    .C(\u_top_module.u_decimator_2.counter[2] ),
    .A(\u_top_module.u_decimator_2.counter[0] ),
    .Y(_0428_));
 sg13g2_nor2_1 _1471_ (.A(_0167_),
    .B(_0428_),
    .Y(_0429_));
 sg13g2_xnor2_1 _1472_ (.Y(_0430_),
    .A(_0167_),
    .B(_0428_));
 sg13g2_o21ai_1 _1473_ (.B1(_0427_),
    .Y(_0049_),
    .A1(_0335_),
    .A2(_0430_));
 sg13g2_nand2_1 _1474_ (.Y(_0431_),
    .A(\u_top_module.u_decimator_2.counter[4] ),
    .B(net918));
 sg13g2_xor2_1 _1475_ (.B(_0429_),
    .A(_0012_),
    .X(_0432_));
 sg13g2_o21ai_1 _1476_ (.B1(_0431_),
    .Y(_0050_),
    .A1(_0335_),
    .A2(_0432_));
 sg13g2_nand2_1 _1477_ (.Y(_0433_),
    .A(\u_top_module.u_decimator_2.counter[5] ),
    .B(net918));
 sg13g2_a21oi_1 _1478_ (.A1(\u_top_module.u_decimator_2.counter[4] ),
    .A2(_0429_),
    .Y(_0434_),
    .B1(\u_top_module.u_decimator_2.counter[5] ));
 sg13g2_nand3_1 _1479_ (.B(\u_top_module.u_decimator_2.counter[4] ),
    .C(_0429_),
    .A(\u_top_module.u_decimator_2.counter[5] ),
    .Y(_0435_));
 sg13g2_nand2b_1 _1480_ (.Y(_0436_),
    .B(_0435_),
    .A_N(_0434_));
 sg13g2_o21ai_1 _1481_ (.B1(_0433_),
    .Y(_0051_),
    .A1(_0335_),
    .A2(_0436_));
 sg13g2_nand2_1 _1482_ (.Y(_0437_),
    .A(\u_top_module.u_decimator_2.counter[6] ),
    .B(net918));
 sg13g2_nor2_1 _1483_ (.A(_0007_),
    .B(_0435_),
    .Y(_0438_));
 sg13g2_xnor2_1 _1484_ (.Y(_0439_),
    .A(_0007_),
    .B(_0435_));
 sg13g2_o21ai_1 _1485_ (.B1(_0437_),
    .Y(_0052_),
    .A1(_0335_),
    .A2(_0439_));
 sg13g2_nand2_1 _1486_ (.Y(_0440_),
    .A(\u_top_module.u_decimator_2.counter[7] ),
    .B(net918));
 sg13g2_xnor2_1 _1487_ (.Y(_0441_),
    .A(_0169_),
    .B(_0438_));
 sg13g2_o21ai_1 _1488_ (.B1(_0440_),
    .Y(_0053_),
    .A1(_0335_),
    .A2(_0441_));
 sg13g2_nor3_1 _1489_ (.A(\u_top_module.addr[2] ),
    .B(\u_top_module.addr[1] ),
    .C(\u_top_module.addr[0] ),
    .Y(_0442_));
 sg13g2_nand2_1 _1490_ (.Y(_0443_),
    .A(net952),
    .B(net942));
 sg13g2_o21ai_1 _1491_ (.B1(_0443_),
    .Y(_0054_),
    .A1(_0174_),
    .A2(net942));
 sg13g2_mux2_1 _1492_ (.A0(\u_top_module.u_memory.memory[0][1] ),
    .A1(\u_top_module.capture_reg[1] ),
    .S(net942),
    .X(_0055_));
 sg13g2_mux2_1 _1493_ (.A0(\u_top_module.u_memory.memory[0][2] ),
    .A1(net950),
    .S(net942),
    .X(_0056_));
 sg13g2_mux2_1 _1494_ (.A0(\u_top_module.u_memory.memory[0][3] ),
    .A1(\u_top_module.capture_reg[3] ),
    .S(net942),
    .X(_0057_));
 sg13g2_mux2_1 _1495_ (.A0(\u_top_module.u_memory.memory[0][4] ),
    .A1(\u_top_module.capture_reg[4] ),
    .S(net942),
    .X(_0058_));
 sg13g2_mux2_1 _1496_ (.A0(\u_top_module.u_memory.memory[0][5] ),
    .A1(\u_top_module.capture_reg[5] ),
    .S(net942),
    .X(_0059_));
 sg13g2_mux2_1 _1497_ (.A0(\u_top_module.u_memory.memory[0][6] ),
    .A1(\u_top_module.capture_reg[6] ),
    .S(net942),
    .X(_0060_));
 sg13g2_mux2_1 _1498_ (.A0(\u_top_module.u_memory.memory[0][7] ),
    .A1(\u_top_module.capture_reg[7] ),
    .S(_0442_),
    .X(_0061_));
 sg13g2_mux2_1 _1499_ (.A0(\u_top_module.u_memory.memory[1][0] ),
    .A1(net952),
    .S(net929),
    .X(_0062_));
 sg13g2_mux2_1 _1500_ (.A0(\u_top_module.u_memory.memory[1][1] ),
    .A1(net951),
    .S(net928),
    .X(_0063_));
 sg13g2_mux2_1 _1501_ (.A0(\u_top_module.u_memory.memory[1][2] ),
    .A1(\u_top_module.capture_reg[2] ),
    .S(net929),
    .X(_0064_));
 sg13g2_mux2_1 _1502_ (.A0(\u_top_module.u_memory.memory[1][3] ),
    .A1(net949),
    .S(net929),
    .X(_0065_));
 sg13g2_mux2_1 _1503_ (.A0(\u_top_module.u_memory.memory[1][4] ),
    .A1(net948),
    .S(net928),
    .X(_0066_));
 sg13g2_mux2_1 _1504_ (.A0(\u_top_module.u_memory.memory[1][5] ),
    .A1(net947),
    .S(net928),
    .X(_0067_));
 sg13g2_mux2_1 _1505_ (.A0(\u_top_module.u_memory.memory[1][6] ),
    .A1(net946),
    .S(net928),
    .X(_0068_));
 sg13g2_mux2_1 _1506_ (.A0(\u_top_module.u_memory.memory[1][7] ),
    .A1(net945),
    .S(net929),
    .X(_0069_));
 sg13g2_mux2_1 _1507_ (.A0(\u_top_module.u_memory.memory[5][0] ),
    .A1(net952),
    .S(net927),
    .X(_0070_));
 sg13g2_mux2_1 _1508_ (.A0(\u_top_module.u_memory.memory[5][1] ),
    .A1(net951),
    .S(net926),
    .X(_0071_));
 sg13g2_mux2_1 _1509_ (.A0(\u_top_module.u_memory.memory[5][2] ),
    .A1(net950),
    .S(net927),
    .X(_0072_));
 sg13g2_mux2_1 _1510_ (.A0(\u_top_module.u_memory.memory[5][3] ),
    .A1(net949),
    .S(net927),
    .X(_0073_));
 sg13g2_mux2_1 _1511_ (.A0(\u_top_module.u_memory.memory[5][4] ),
    .A1(net948),
    .S(net926),
    .X(_0074_));
 sg13g2_mux2_1 _1512_ (.A0(\u_top_module.u_memory.memory[5][5] ),
    .A1(net947),
    .S(net926),
    .X(_0075_));
 sg13g2_mux2_1 _1513_ (.A0(\u_top_module.u_memory.memory[5][6] ),
    .A1(net946),
    .S(net926),
    .X(_0076_));
 sg13g2_mux2_1 _1514_ (.A0(\u_top_module.u_memory.memory[5][7] ),
    .A1(net945),
    .S(net927),
    .X(_0077_));
 sg13g2_mux2_1 _1515_ (.A0(\u_top_module.u_memory.memory[2][0] ),
    .A1(net952),
    .S(net935),
    .X(_0078_));
 sg13g2_mux2_1 _1516_ (.A0(\u_top_module.u_memory.memory[2][1] ),
    .A1(net951),
    .S(net934),
    .X(_0079_));
 sg13g2_mux2_1 _1517_ (.A0(\u_top_module.u_memory.memory[2][2] ),
    .A1(net950),
    .S(net935),
    .X(_0080_));
 sg13g2_mux2_1 _1518_ (.A0(\u_top_module.u_memory.memory[2][3] ),
    .A1(net949),
    .S(net935),
    .X(_0081_));
 sg13g2_mux2_1 _1519_ (.A0(\u_top_module.u_memory.memory[2][4] ),
    .A1(net948),
    .S(net934),
    .X(_0082_));
 sg13g2_mux2_1 _1520_ (.A0(\u_top_module.u_memory.memory[2][5] ),
    .A1(net947),
    .S(net934),
    .X(_0083_));
 sg13g2_mux2_1 _1521_ (.A0(\u_top_module.u_memory.memory[2][6] ),
    .A1(net946),
    .S(net934),
    .X(_0084_));
 sg13g2_mux2_1 _1522_ (.A0(\u_top_module.u_memory.memory[2][7] ),
    .A1(net945),
    .S(net935),
    .X(_0085_));
 sg13g2_mux2_1 _1523_ (.A0(\u_top_module.u_memory.memory[3][0] ),
    .A1(net952),
    .S(net933),
    .X(_0086_));
 sg13g2_mux2_1 _1524_ (.A0(\u_top_module.u_memory.memory[3][1] ),
    .A1(net951),
    .S(net932),
    .X(_0087_));
 sg13g2_mux2_1 _1525_ (.A0(\u_top_module.u_memory.memory[3][2] ),
    .A1(net950),
    .S(net933),
    .X(_0088_));
 sg13g2_mux2_1 _1526_ (.A0(\u_top_module.u_memory.memory[3][3] ),
    .A1(net949),
    .S(net933),
    .X(_0089_));
 sg13g2_mux2_1 _1527_ (.A0(\u_top_module.u_memory.memory[3][4] ),
    .A1(net948),
    .S(net932),
    .X(_0090_));
 sg13g2_mux2_1 _1528_ (.A0(\u_top_module.u_memory.memory[3][5] ),
    .A1(net947),
    .S(net932),
    .X(_0091_));
 sg13g2_mux2_1 _1529_ (.A0(\u_top_module.u_memory.memory[3][6] ),
    .A1(net946),
    .S(net932),
    .X(_0092_));
 sg13g2_mux2_1 _1530_ (.A0(\u_top_module.u_memory.memory[3][7] ),
    .A1(net945),
    .S(net933),
    .X(_0093_));
 sg13g2_mux2_1 _1531_ (.A0(\u_top_module.u_memory.memory[6][0] ),
    .A1(net952),
    .S(net931),
    .X(_0094_));
 sg13g2_mux2_1 _1532_ (.A0(\u_top_module.u_memory.memory[6][1] ),
    .A1(net951),
    .S(net930),
    .X(_0095_));
 sg13g2_mux2_1 _1533_ (.A0(\u_top_module.u_memory.memory[6][2] ),
    .A1(net950),
    .S(net931),
    .X(_0096_));
 sg13g2_mux2_1 _1534_ (.A0(\u_top_module.u_memory.memory[6][3] ),
    .A1(net949),
    .S(net931),
    .X(_0097_));
 sg13g2_mux2_1 _1535_ (.A0(\u_top_module.u_memory.memory[6][4] ),
    .A1(net948),
    .S(net930),
    .X(_0098_));
 sg13g2_mux2_1 _1536_ (.A0(\u_top_module.u_memory.memory[6][5] ),
    .A1(net947),
    .S(net930),
    .X(_0099_));
 sg13g2_mux2_1 _1537_ (.A0(\u_top_module.u_memory.memory[6][6] ),
    .A1(net946),
    .S(net930),
    .X(_0100_));
 sg13g2_mux2_1 _1538_ (.A0(\u_top_module.u_memory.memory[6][7] ),
    .A1(net945),
    .S(net931),
    .X(_0101_));
 sg13g2_mux2_1 _1539_ (.A0(\u_top_module.u_memory.memory[4][0] ),
    .A1(net952),
    .S(net944),
    .X(_0102_));
 sg13g2_mux2_1 _1540_ (.A0(\u_top_module.u_memory.memory[4][1] ),
    .A1(net951),
    .S(net943),
    .X(_0103_));
 sg13g2_mux2_1 _1541_ (.A0(\u_top_module.u_memory.memory[4][2] ),
    .A1(net950),
    .S(net944),
    .X(_0104_));
 sg13g2_mux2_1 _1542_ (.A0(\u_top_module.u_memory.memory[4][3] ),
    .A1(net949),
    .S(net944),
    .X(_0105_));
 sg13g2_mux2_1 _1543_ (.A0(\u_top_module.u_memory.memory[4][4] ),
    .A1(net948),
    .S(net943),
    .X(_0106_));
 sg13g2_mux2_1 _1544_ (.A0(\u_top_module.u_memory.memory[4][5] ),
    .A1(net947),
    .S(net943),
    .X(_0107_));
 sg13g2_mux2_1 _1545_ (.A0(\u_top_module.u_memory.memory[4][6] ),
    .A1(net946),
    .S(net943),
    .X(_0108_));
 sg13g2_mux2_1 _1546_ (.A0(\u_top_module.u_memory.memory[4][7] ),
    .A1(net945),
    .S(net944),
    .X(_0109_));
 sg13g2_nor2_2 _1547_ (.A(_0026_),
    .B(\u_top_module.u_spi_port.cs_n_prev ),
    .Y(_0444_));
 sg13g2_mux2_1 _1548_ (.A0(\u_top_module.capture_reg[0] ),
    .A1(\u_top_module.u_spi_port.shift_reg[0] ),
    .S(net940),
    .X(_0110_));
 sg13g2_mux2_1 _1549_ (.A0(net951),
    .A1(\u_top_module.u_spi_port.shift_reg[1] ),
    .S(net941),
    .X(_0111_));
 sg13g2_mux2_1 _1550_ (.A0(net950),
    .A1(\u_top_module.u_spi_port.shift_reg[2] ),
    .S(net941),
    .X(_0112_));
 sg13g2_mux2_1 _1551_ (.A0(net949),
    .A1(\u_top_module.u_spi_port.shift_reg[3] ),
    .S(net941),
    .X(_0113_));
 sg13g2_mux2_1 _1552_ (.A0(net948),
    .A1(\u_top_module.u_spi_port.shift_reg[4] ),
    .S(net941),
    .X(_0114_));
 sg13g2_mux2_1 _1553_ (.A0(net947),
    .A1(\u_top_module.u_spi_port.shift_reg[5] ),
    .S(net941),
    .X(_0115_));
 sg13g2_mux2_1 _1554_ (.A0(net946),
    .A1(\u_top_module.u_spi_port.shift_reg[6] ),
    .S(net941),
    .X(_0116_));
 sg13g2_mux2_1 _1555_ (.A0(net945),
    .A1(\u_top_module.u_spi_port.shift_reg[7] ),
    .S(net941),
    .X(_0117_));
 sg13g2_mux2_1 _1556_ (.A0(\u_top_module.addr[0] ),
    .A1(\u_top_module.u_spi_port.shift_reg[8] ),
    .S(net940),
    .X(_0118_));
 sg13g2_nand2_1 _1557_ (.Y(_0445_),
    .A(\u_top_module.u_spi_port.shift_reg[9] ),
    .B(net940));
 sg13g2_o21ai_1 _1558_ (.B1(_0445_),
    .Y(_0119_),
    .A1(_0166_),
    .A2(net940));
 sg13g2_mux2_1 _1559_ (.A0(\u_top_module.addr[2] ),
    .A1(\u_top_module.u_spi_port.shift_reg[10] ),
    .S(net940),
    .X(_0120_));
 sg13g2_mux2_1 _1560_ (.A0(\u_top_module.addr[3] ),
    .A1(\u_top_module.u_spi_port.shift_reg[11] ),
    .S(net940),
    .X(_0121_));
 sg13g2_mux2_1 _1561_ (.A0(\u_top_module.addr[4] ),
    .A1(\u_top_module.u_spi_port.shift_reg[12] ),
    .S(_0444_),
    .X(_0122_));
 sg13g2_mux2_1 _1562_ (.A0(\u_top_module.addr[5] ),
    .A1(\u_top_module.u_spi_port.shift_reg[13] ),
    .S(_0444_),
    .X(_0123_));
 sg13g2_mux2_1 _1563_ (.A0(\u_top_module.addr[6] ),
    .A1(\u_top_module.u_spi_port.shift_reg[14] ),
    .S(net940),
    .X(_0124_));
 sg13g2_mux2_1 _1564_ (.A0(\u_top_module.addr[7] ),
    .A1(\u_top_module.u_spi_port.shift_reg[15] ),
    .S(net940),
    .X(_0125_));
 sg13g2_mux2_1 _1565_ (.A0(\u_top_module.u_memory.memory[7][0] ),
    .A1(net952),
    .S(net937),
    .X(_0126_));
 sg13g2_mux2_1 _1566_ (.A0(\u_top_module.u_memory.memory[7][1] ),
    .A1(net951),
    .S(net936),
    .X(_0127_));
 sg13g2_mux2_1 _1567_ (.A0(\u_top_module.u_memory.memory[7][2] ),
    .A1(net950),
    .S(net937),
    .X(_0128_));
 sg13g2_mux2_1 _1568_ (.A0(\u_top_module.u_memory.memory[7][3] ),
    .A1(net949),
    .S(net937),
    .X(_0129_));
 sg13g2_mux2_1 _1569_ (.A0(\u_top_module.u_memory.memory[7][4] ),
    .A1(net948),
    .S(net936),
    .X(_0130_));
 sg13g2_mux2_1 _1570_ (.A0(\u_top_module.u_memory.memory[7][5] ),
    .A1(net947),
    .S(net936),
    .X(_0131_));
 sg13g2_mux2_1 _1571_ (.A0(\u_top_module.u_memory.memory[7][6] ),
    .A1(net946),
    .S(net936),
    .X(_0132_));
 sg13g2_mux2_1 _1572_ (.A0(\u_top_module.u_memory.memory[7][7] ),
    .A1(net945),
    .S(net937),
    .X(_0133_));
 sg13g2_nand2_1 _1573_ (.Y(_0446_),
    .A(_0026_),
    .B(net972));
 sg13g2_mux2_1 _1574_ (.A0(net1),
    .A1(\u_top_module.u_spi_port.shift_reg[0] ),
    .S(net938),
    .X(_0134_));
 sg13g2_mux2_1 _1575_ (.A0(\u_top_module.u_spi_port.shift_reg[0] ),
    .A1(\u_top_module.u_spi_port.shift_reg[1] ),
    .S(net938),
    .X(_0135_));
 sg13g2_mux2_1 _1576_ (.A0(\u_top_module.u_spi_port.shift_reg[1] ),
    .A1(\u_top_module.u_spi_port.shift_reg[2] ),
    .S(net939),
    .X(_0136_));
 sg13g2_mux2_1 _1577_ (.A0(\u_top_module.u_spi_port.shift_reg[2] ),
    .A1(\u_top_module.u_spi_port.shift_reg[3] ),
    .S(net939),
    .X(_0137_));
 sg13g2_mux2_1 _1578_ (.A0(\u_top_module.u_spi_port.shift_reg[3] ),
    .A1(\u_top_module.u_spi_port.shift_reg[4] ),
    .S(net939),
    .X(_0138_));
 sg13g2_mux2_1 _1579_ (.A0(\u_top_module.u_spi_port.shift_reg[4] ),
    .A1(\u_top_module.u_spi_port.shift_reg[5] ),
    .S(net939),
    .X(_0139_));
 sg13g2_mux2_1 _1580_ (.A0(\u_top_module.u_spi_port.shift_reg[5] ),
    .A1(\u_top_module.u_spi_port.shift_reg[6] ),
    .S(net939),
    .X(_0140_));
 sg13g2_mux2_1 _1581_ (.A0(\u_top_module.u_spi_port.shift_reg[6] ),
    .A1(\u_top_module.u_spi_port.shift_reg[7] ),
    .S(net939),
    .X(_0141_));
 sg13g2_mux2_1 _1582_ (.A0(\u_top_module.u_spi_port.shift_reg[7] ),
    .A1(\u_top_module.u_spi_port.shift_reg[8] ),
    .S(net939),
    .X(_0142_));
 sg13g2_mux2_1 _1583_ (.A0(\u_top_module.u_spi_port.shift_reg[8] ),
    .A1(\u_top_module.u_spi_port.shift_reg[9] ),
    .S(net938),
    .X(_0143_));
 sg13g2_mux2_1 _1584_ (.A0(\u_top_module.u_spi_port.shift_reg[9] ),
    .A1(\u_top_module.u_spi_port.shift_reg[10] ),
    .S(net938),
    .X(_0144_));
 sg13g2_mux2_1 _1585_ (.A0(\u_top_module.u_spi_port.shift_reg[10] ),
    .A1(\u_top_module.u_spi_port.shift_reg[11] ),
    .S(net938),
    .X(_0145_));
 sg13g2_mux2_1 _1586_ (.A0(\u_top_module.u_spi_port.shift_reg[11] ),
    .A1(\u_top_module.u_spi_port.shift_reg[12] ),
    .S(_0446_),
    .X(_0146_));
 sg13g2_mux2_1 _1587_ (.A0(\u_top_module.u_spi_port.shift_reg[12] ),
    .A1(\u_top_module.u_spi_port.shift_reg[13] ),
    .S(net938),
    .X(_0147_));
 sg13g2_mux2_1 _1588_ (.A0(\u_top_module.u_spi_port.shift_reg[13] ),
    .A1(\u_top_module.u_spi_port.shift_reg[14] ),
    .S(net938),
    .X(_0148_));
 sg13g2_mux2_1 _1589_ (.A0(\u_top_module.u_spi_port.shift_reg[14] ),
    .A1(\u_top_module.u_spi_port.shift_reg[15] ),
    .S(net938),
    .X(_0149_));
 sg13g2_xnor2_1 _1590_ (.Y(_0447_),
    .A(\u_top_module.u_buffer.shift_reg_1[255] ),
    .B(\u_top_module.u_buffer.shift_reg_2[254] ));
 sg13g2_xor2_1 _1591_ (.B(\u_top_module.u_buffer.shift_reg_1[0] ),
    .A(\u_top_module.dec_data_2 ),
    .X(_0448_));
 sg13g2_nor2_1 _1592_ (.A(_0447_),
    .B(_0448_),
    .Y(_0449_));
 sg13g2_xor2_1 _1593_ (.B(_0448_),
    .A(_0447_),
    .X(_0450_));
 sg13g2_nor2_1 _1594_ (.A(_0016_),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_xnor2_1 _1595_ (.Y(_0452_),
    .A(_0016_),
    .B(_0450_));
 sg13g2_nand2_1 _1596_ (.Y(_0453_),
    .A(\u_top_module.u_buffer.corr_neg[0] ),
    .B(net924));
 sg13g2_o21ai_1 _1597_ (.B1(_0453_),
    .Y(_0150_),
    .A1(net923),
    .A2(_0452_));
 sg13g2_nor2_1 _1598_ (.A(\u_top_module.u_buffer.corr_neg[1] ),
    .B(_0449_),
    .Y(_0454_));
 sg13g2_nand2_1 _1599_ (.Y(_0455_),
    .A(\u_top_module.u_buffer.corr_neg[1] ),
    .B(_0449_));
 sg13g2_nand2b_1 _1600_ (.Y(_0456_),
    .B(_0455_),
    .A_N(_0454_));
 sg13g2_xnor2_1 _1601_ (.Y(_0457_),
    .A(_0451_),
    .B(_0456_));
 sg13g2_nor2_1 _1602_ (.A(net923),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_a21oi_1 _1603_ (.A1(_0187_),
    .A2(net923),
    .Y(_0151_),
    .B1(_0458_));
 sg13g2_a21oi_1 _1604_ (.A1(_0451_),
    .A2(_0455_),
    .Y(_0459_),
    .B1(_0454_));
 sg13g2_a21o_1 _1605_ (.A2(_0455_),
    .A1(_0451_),
    .B1(_0454_),
    .X(_0460_));
 sg13g2_nor2_1 _1606_ (.A(\u_top_module.u_buffer.corr_neg[2] ),
    .B(_0187_),
    .Y(_0461_));
 sg13g2_nor2_1 _1607_ (.A(_0185_),
    .B(\u_top_module.u_buffer.corr_neg[1] ),
    .Y(_0462_));
 sg13g2_nor2_1 _1608_ (.A(_0461_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_xnor2_1 _1609_ (.Y(_0464_),
    .A(_0459_),
    .B(_0463_));
 sg13g2_nor2_1 _1610_ (.A(net924),
    .B(_0464_),
    .Y(_0465_));
 sg13g2_a21oi_1 _1611_ (.A1(_0185_),
    .A2(net924),
    .Y(_0152_),
    .B1(_0465_));
 sg13g2_xor2_1 _1612_ (.B(\u_top_module.u_buffer.corr_neg[2] ),
    .A(\u_top_module.u_buffer.corr_neg[3] ),
    .X(_0466_));
 sg13g2_a21oi_1 _1613_ (.A1(_0460_),
    .A2(_0463_),
    .Y(_0467_),
    .B1(_0461_));
 sg13g2_xor2_1 _1614_ (.B(_0467_),
    .A(_0466_),
    .X(_0468_));
 sg13g2_nor2_1 _1615_ (.A(net924),
    .B(_0468_),
    .Y(_0469_));
 sg13g2_a21oi_1 _1616_ (.A1(_0183_),
    .A2(net924),
    .Y(_0153_),
    .B1(_0469_));
 sg13g2_nand2_1 _1617_ (.Y(_0470_),
    .A(\u_top_module.u_buffer.corr_neg[4] ),
    .B(net922));
 sg13g2_or3_1 _1618_ (.A(_0461_),
    .B(_0462_),
    .C(_0466_),
    .X(_0471_));
 sg13g2_o21ai_1 _1619_ (.B1(_0183_),
    .Y(_0472_),
    .A1(\u_top_module.u_buffer.corr_neg[2] ),
    .A2(\u_top_module.u_buffer.corr_neg[1] ));
 sg13g2_o21ai_1 _1620_ (.B1(_0472_),
    .Y(_0473_),
    .A1(_0459_),
    .A2(_0471_));
 sg13g2_nor2_1 _1621_ (.A(\u_top_module.u_buffer.corr_neg[4] ),
    .B(_0183_),
    .Y(_0474_));
 sg13g2_xnor2_1 _1622_ (.Y(_0475_),
    .A(\u_top_module.u_buffer.corr_neg[4] ),
    .B(\u_top_module.u_buffer.corr_neg[3] ));
 sg13g2_xnor2_1 _1623_ (.Y(_0476_),
    .A(_0473_),
    .B(_0475_));
 sg13g2_o21ai_1 _1624_ (.B1(_0470_),
    .Y(_0154_),
    .A1(net922),
    .A2(_0476_));
 sg13g2_xnor2_1 _1625_ (.Y(_0477_),
    .A(\u_top_module.u_buffer.corr_neg[5] ),
    .B(\u_top_module.u_buffer.corr_neg[4] ));
 sg13g2_a21oi_1 _1626_ (.A1(_0473_),
    .A2(_0475_),
    .Y(_0478_),
    .B1(_0474_));
 sg13g2_xor2_1 _1627_ (.B(_0478_),
    .A(_0477_),
    .X(_0479_));
 sg13g2_nand2_1 _1628_ (.Y(_0480_),
    .A(net821),
    .B(net920));
 sg13g2_o21ai_1 _1629_ (.B1(_0480_),
    .Y(_0155_),
    .A1(net922),
    .A2(_0479_));
 sg13g2_nand2_1 _1630_ (.Y(_0481_),
    .A(_0177_),
    .B(net821));
 sg13g2_nor2_1 _1631_ (.A(_0177_),
    .B(net821),
    .Y(_0482_));
 sg13g2_xnor2_1 _1632_ (.Y(_0483_),
    .A(\u_top_module.u_buffer.corr_neg[6] ),
    .B(net821));
 sg13g2_and2_1 _1633_ (.A(_0475_),
    .B(_0477_),
    .X(_0484_));
 sg13g2_a21oi_1 _1634_ (.A1(_0180_),
    .A2(_0183_),
    .Y(_0485_),
    .B1(net821));
 sg13g2_a21oi_1 _1635_ (.A1(_0473_),
    .A2(_0484_),
    .Y(_0486_),
    .B1(_0485_));
 sg13g2_xnor2_1 _1636_ (.Y(_0487_),
    .A(_0483_),
    .B(_0486_));
 sg13g2_nor2_1 _1637_ (.A(net920),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_a21oi_1 _1638_ (.A1(_0177_),
    .A2(net920),
    .Y(_0156_),
    .B1(_0488_));
 sg13g2_o21ai_1 _1639_ (.B1(_0481_),
    .Y(_0489_),
    .A1(_0482_),
    .A2(_0486_));
 sg13g2_xnor2_1 _1640_ (.Y(_0490_),
    .A(\u_top_module.u_buffer.corr_neg[7] ),
    .B(\u_top_module.u_buffer.corr_neg[6] ));
 sg13g2_xnor2_1 _1641_ (.Y(_0491_),
    .A(_0489_),
    .B(_0490_));
 sg13g2_nand2_1 _1642_ (.Y(_0492_),
    .A(\u_top_module.u_buffer.corr_neg[7] ),
    .B(net920));
 sg13g2_o21ai_1 _1643_ (.B1(_0492_),
    .Y(_0157_),
    .A1(net920),
    .A2(_0491_));
 sg13g2_dfrbp_1 _1644_ (.CLK(net840),
    .RESET_B(net994),
    .D(\u_top_module.u_buffer.shift_reg_2[98] ),
    .Q_N(_0613_),
    .Q(\u_top_module.u_buffer.shift_reg_2[99] ));
 sg13g2_dfrbp_1 _1645_ (.CLK(net840),
    .RESET_B(net994),
    .D(\u_top_module.u_buffer.shift_reg_2[99] ),
    .Q_N(_0614_),
    .Q(\u_top_module.u_buffer.shift_reg_2[100] ));
 sg13g2_dfrbp_1 _1646_ (.CLK(net840),
    .RESET_B(net994),
    .D(\u_top_module.u_buffer.shift_reg_2[100] ),
    .Q_N(_0615_),
    .Q(\u_top_module.u_buffer.shift_reg_2[101] ));
 sg13g2_dfrbp_1 _1647_ (.CLK(net842),
    .RESET_B(net996),
    .D(\u_top_module.u_buffer.shift_reg_2[101] ),
    .Q_N(_0616_),
    .Q(\u_top_module.u_buffer.shift_reg_2[102] ));
 sg13g2_dfrbp_1 _1648_ (.CLK(net842),
    .RESET_B(net996),
    .D(\u_top_module.u_buffer.shift_reg_2[102] ),
    .Q_N(_0617_),
    .Q(\u_top_module.u_buffer.shift_reg_2[103] ));
 sg13g2_dfrbp_1 _1649_ (.CLK(net842),
    .RESET_B(net996),
    .D(\u_top_module.u_buffer.shift_reg_2[103] ),
    .Q_N(_0618_),
    .Q(\u_top_module.u_buffer.shift_reg_2[104] ));
 sg13g2_dfrbp_1 _1650_ (.CLK(net842),
    .RESET_B(net996),
    .D(\u_top_module.u_buffer.shift_reg_2[104] ),
    .Q_N(_0619_),
    .Q(\u_top_module.u_buffer.shift_reg_2[105] ));
 sg13g2_dfrbp_1 _1651_ (.CLK(net842),
    .RESET_B(net996),
    .D(\u_top_module.u_buffer.shift_reg_2[105] ),
    .Q_N(_0620_),
    .Q(\u_top_module.u_buffer.shift_reg_2[106] ));
 sg13g2_dfrbp_1 _1652_ (.CLK(net842),
    .RESET_B(net996),
    .D(\u_top_module.u_buffer.shift_reg_2[106] ),
    .Q_N(_0621_),
    .Q(\u_top_module.u_buffer.shift_reg_2[107] ));
 sg13g2_dfrbp_1 _1653_ (.CLK(net845),
    .RESET_B(net999),
    .D(\u_top_module.u_buffer.shift_reg_2[107] ),
    .Q_N(_0622_),
    .Q(\u_top_module.u_buffer.shift_reg_2[108] ));
 sg13g2_dfrbp_1 _1654_ (.CLK(net845),
    .RESET_B(net999),
    .D(\u_top_module.u_buffer.shift_reg_2[108] ),
    .Q_N(_0623_),
    .Q(\u_top_module.u_buffer.shift_reg_2[109] ));
 sg13g2_dfrbp_1 _1655_ (.CLK(net845),
    .RESET_B(net999),
    .D(\u_top_module.u_buffer.shift_reg_2[109] ),
    .Q_N(_0624_),
    .Q(\u_top_module.u_buffer.shift_reg_2[110] ));
 sg13g2_dfrbp_1 _1656_ (.CLK(net842),
    .RESET_B(net996),
    .D(\u_top_module.u_buffer.shift_reg_2[110] ),
    .Q_N(_0625_),
    .Q(\u_top_module.u_buffer.shift_reg_2[111] ));
 sg13g2_dfrbp_1 _1657_ (.CLK(net842),
    .RESET_B(net996),
    .D(\u_top_module.u_buffer.shift_reg_2[111] ),
    .Q_N(_0626_),
    .Q(\u_top_module.u_buffer.shift_reg_2[112] ));
 sg13g2_dfrbp_1 _1658_ (.CLK(net885),
    .RESET_B(net1040),
    .D(\u_top_module.u_buffer.shift_reg_2[112] ),
    .Q_N(_0627_),
    .Q(\u_top_module.u_buffer.shift_reg_2[113] ));
 sg13g2_dfrbp_1 _1659_ (.CLK(net885),
    .RESET_B(net1040),
    .D(\u_top_module.u_buffer.shift_reg_2[113] ),
    .Q_N(_0628_),
    .Q(\u_top_module.u_buffer.shift_reg_2[114] ));
 sg13g2_dfrbp_1 _1660_ (.CLK(net885),
    .RESET_B(net1040),
    .D(\u_top_module.u_buffer.shift_reg_2[114] ),
    .Q_N(_0629_),
    .Q(\u_top_module.u_buffer.shift_reg_2[115] ));
 sg13g2_dfrbp_1 _1661_ (.CLK(net885),
    .RESET_B(net1040),
    .D(\u_top_module.u_buffer.shift_reg_2[115] ),
    .Q_N(_0630_),
    .Q(\u_top_module.u_buffer.shift_reg_2[116] ));
 sg13g2_dfrbp_1 _1662_ (.CLK(net886),
    .RESET_B(net1043),
    .D(\u_top_module.u_buffer.shift_reg_2[116] ),
    .Q_N(_0631_),
    .Q(\u_top_module.u_buffer.shift_reg_2[117] ));
 sg13g2_dfrbp_1 _1663_ (.CLK(net886),
    .RESET_B(net1043),
    .D(\u_top_module.u_buffer.shift_reg_2[117] ),
    .Q_N(_0632_),
    .Q(\u_top_module.u_buffer.shift_reg_2[118] ));
 sg13g2_dfrbp_1 _1664_ (.CLK(net886),
    .RESET_B(net1041),
    .D(\u_top_module.u_buffer.shift_reg_2[118] ),
    .Q_N(_0633_),
    .Q(\u_top_module.u_buffer.shift_reg_2[119] ));
 sg13g2_dfrbp_1 _1665_ (.CLK(net886),
    .RESET_B(net1041),
    .D(\u_top_module.u_buffer.shift_reg_2[119] ),
    .Q_N(_0634_),
    .Q(\u_top_module.u_buffer.shift_reg_2[120] ));
 sg13g2_dfrbp_1 _1666_ (.CLK(net889),
    .RESET_B(net1044),
    .D(\u_top_module.u_buffer.shift_reg_2[120] ),
    .Q_N(_0635_),
    .Q(\u_top_module.u_buffer.shift_reg_2[121] ));
 sg13g2_dfrbp_1 _1667_ (.CLK(net889),
    .RESET_B(net1044),
    .D(\u_top_module.u_buffer.shift_reg_2[121] ),
    .Q_N(_0636_),
    .Q(\u_top_module.u_buffer.shift_reg_2[122] ));
 sg13g2_dfrbp_1 _1668_ (.CLK(net889),
    .RESET_B(net1044),
    .D(\u_top_module.u_buffer.shift_reg_2[122] ),
    .Q_N(_0637_),
    .Q(\u_top_module.u_buffer.shift_reg_2[123] ));
 sg13g2_dfrbp_1 _1669_ (.CLK(net890),
    .RESET_B(net1045),
    .D(\u_top_module.u_buffer.shift_reg_2[123] ),
    .Q_N(_0638_),
    .Q(\u_top_module.u_buffer.shift_reg_2[124] ));
 sg13g2_dfrbp_1 _1670_ (.CLK(net890),
    .RESET_B(net1045),
    .D(\u_top_module.u_buffer.shift_reg_2[124] ),
    .Q_N(_0639_),
    .Q(\u_top_module.u_buffer.shift_reg_2[125] ));
 sg13g2_dfrbp_1 _1671_ (.CLK(net890),
    .RESET_B(net1045),
    .D(\u_top_module.u_buffer.shift_reg_2[125] ),
    .Q_N(_0640_),
    .Q(\u_top_module.u_buffer.shift_reg_2[126] ));
 sg13g2_dfrbp_1 _1672_ (.CLK(net890),
    .RESET_B(net1045),
    .D(\u_top_module.u_buffer.shift_reg_2[126] ),
    .Q_N(_0641_),
    .Q(\u_top_module.u_buffer.shift_reg_2[127] ));
 sg13g2_dfrbp_1 _1673_ (.CLK(net900),
    .RESET_B(net1054),
    .D(\u_top_module.u_buffer.shift_reg_2[127] ),
    .Q_N(_0642_),
    .Q(\u_top_module.u_buffer.shift_reg_2[128] ));
 sg13g2_dfrbp_1 _1674_ (.CLK(net900),
    .RESET_B(net1054),
    .D(\u_top_module.u_buffer.shift_reg_2[128] ),
    .Q_N(_0643_),
    .Q(\u_top_module.u_buffer.shift_reg_2[129] ));
 sg13g2_dfrbp_1 _1675_ (.CLK(net900),
    .RESET_B(net1054),
    .D(\u_top_module.u_buffer.shift_reg_2[129] ),
    .Q_N(_0644_),
    .Q(\u_top_module.u_buffer.shift_reg_2[130] ));
 sg13g2_dfrbp_1 _1676_ (.CLK(net900),
    .RESET_B(net1054),
    .D(\u_top_module.u_buffer.shift_reg_2[130] ),
    .Q_N(_0645_),
    .Q(\u_top_module.u_buffer.shift_reg_2[131] ));
 sg13g2_dfrbp_1 _1677_ (.CLK(net901),
    .RESET_B(net1055),
    .D(\u_top_module.u_buffer.shift_reg_2[131] ),
    .Q_N(_0646_),
    .Q(\u_top_module.u_buffer.shift_reg_2[132] ));
 sg13g2_dfrbp_1 _1678_ (.CLK(net901),
    .RESET_B(net1055),
    .D(\u_top_module.u_buffer.shift_reg_2[132] ),
    .Q_N(_0647_),
    .Q(\u_top_module.u_buffer.shift_reg_2[133] ));
 sg13g2_dfrbp_1 _1679_ (.CLK(net901),
    .RESET_B(net1055),
    .D(\u_top_module.u_buffer.shift_reg_2[133] ),
    .Q_N(_0648_),
    .Q(\u_top_module.u_buffer.shift_reg_2[134] ));
 sg13g2_dfrbp_1 _1680_ (.CLK(net902),
    .RESET_B(net1056),
    .D(\u_top_module.u_buffer.shift_reg_2[134] ),
    .Q_N(_0649_),
    .Q(\u_top_module.u_buffer.shift_reg_2[135] ));
 sg13g2_dfrbp_1 _1681_ (.CLK(net902),
    .RESET_B(net1056),
    .D(\u_top_module.u_buffer.shift_reg_2[135] ),
    .Q_N(_0650_),
    .Q(\u_top_module.u_buffer.shift_reg_2[136] ));
 sg13g2_dfrbp_1 _1682_ (.CLK(net902),
    .RESET_B(net1056),
    .D(\u_top_module.u_buffer.shift_reg_2[136] ),
    .Q_N(_0651_),
    .Q(\u_top_module.u_buffer.shift_reg_2[137] ));
 sg13g2_dfrbp_1 _1683_ (.CLK(net902),
    .RESET_B(net1056),
    .D(\u_top_module.u_buffer.shift_reg_2[137] ),
    .Q_N(_0652_),
    .Q(\u_top_module.u_buffer.shift_reg_2[138] ));
 sg13g2_dfrbp_1 _1684_ (.CLK(net902),
    .RESET_B(net1056),
    .D(\u_top_module.u_buffer.shift_reg_2[138] ),
    .Q_N(_0653_),
    .Q(\u_top_module.u_buffer.shift_reg_2[139] ));
 sg13g2_dfrbp_1 _1685_ (.CLK(net902),
    .RESET_B(net1056),
    .D(\u_top_module.u_buffer.shift_reg_2[139] ),
    .Q_N(_0654_),
    .Q(\u_top_module.u_buffer.shift_reg_2[140] ));
 sg13g2_dfrbp_1 _1686_ (.CLK(net905),
    .RESET_B(net1059),
    .D(\u_top_module.u_buffer.shift_reg_2[140] ),
    .Q_N(_0655_),
    .Q(\u_top_module.u_buffer.shift_reg_2[141] ));
 sg13g2_dfrbp_1 _1687_ (.CLK(net905),
    .RESET_B(net1059),
    .D(\u_top_module.u_buffer.shift_reg_2[141] ),
    .Q_N(_0656_),
    .Q(\u_top_module.u_buffer.shift_reg_2[142] ));
 sg13g2_dfrbp_1 _1688_ (.CLK(net905),
    .RESET_B(net1059),
    .D(\u_top_module.u_buffer.shift_reg_2[142] ),
    .Q_N(_0657_),
    .Q(\u_top_module.u_buffer.shift_reg_2[143] ));
 sg13g2_dfrbp_1 _1689_ (.CLK(net905),
    .RESET_B(net1059),
    .D(\u_top_module.u_buffer.shift_reg_2[143] ),
    .Q_N(_0658_),
    .Q(\u_top_module.u_buffer.shift_reg_2[144] ));
 sg13g2_dfrbp_1 _1690_ (.CLK(net905),
    .RESET_B(net1059),
    .D(\u_top_module.u_buffer.shift_reg_2[144] ),
    .Q_N(_0659_),
    .Q(\u_top_module.u_buffer.shift_reg_2[145] ));
 sg13g2_dfrbp_1 _1691_ (.CLK(net905),
    .RESET_B(net1059),
    .D(\u_top_module.u_buffer.shift_reg_2[145] ),
    .Q_N(_0660_),
    .Q(\u_top_module.u_buffer.shift_reg_2[146] ));
 sg13g2_dfrbp_1 _1692_ (.CLK(net906),
    .RESET_B(net1060),
    .D(\u_top_module.u_buffer.shift_reg_2[146] ),
    .Q_N(_0661_),
    .Q(\u_top_module.u_buffer.shift_reg_2[147] ));
 sg13g2_dfrbp_1 _1693_ (.CLK(net910),
    .RESET_B(net1060),
    .D(\u_top_module.u_buffer.shift_reg_2[147] ),
    .Q_N(_0662_),
    .Q(\u_top_module.u_buffer.shift_reg_2[148] ));
 sg13g2_dfrbp_1 _1694_ (.CLK(net910),
    .RESET_B(net1066),
    .D(\u_top_module.u_buffer.shift_reg_2[148] ),
    .Q_N(_0663_),
    .Q(\u_top_module.u_buffer.shift_reg_2[149] ));
 sg13g2_dfrbp_1 _1695_ (.CLK(net910),
    .RESET_B(net1066),
    .D(\u_top_module.u_buffer.shift_reg_2[149] ),
    .Q_N(_0664_),
    .Q(\u_top_module.u_buffer.shift_reg_2[150] ));
 sg13g2_dfrbp_1 _1696_ (.CLK(net910),
    .RESET_B(net1060),
    .D(\u_top_module.u_buffer.shift_reg_2[150] ),
    .Q_N(_0665_),
    .Q(\u_top_module.u_buffer.shift_reg_2[151] ));
 sg13g2_dfrbp_1 _1697_ (.CLK(net906),
    .RESET_B(net1060),
    .D(\u_top_module.u_buffer.shift_reg_2[151] ),
    .Q_N(_0666_),
    .Q(\u_top_module.u_buffer.shift_reg_2[152] ));
 sg13g2_dfrbp_1 _1698_ (.CLK(net905),
    .RESET_B(net1059),
    .D(\u_top_module.u_buffer.shift_reg_2[152] ),
    .Q_N(_0667_),
    .Q(\u_top_module.u_buffer.shift_reg_2[153] ));
 sg13g2_dfrbp_1 _1699_ (.CLK(net905),
    .RESET_B(net1059),
    .D(\u_top_module.u_buffer.shift_reg_2[153] ),
    .Q_N(_0668_),
    .Q(\u_top_module.u_buffer.shift_reg_2[154] ));
 sg13g2_dfrbp_1 _1700_ (.CLK(net904),
    .RESET_B(net1057),
    .D(\u_top_module.u_buffer.shift_reg_2[154] ),
    .Q_N(_0669_),
    .Q(\u_top_module.u_buffer.shift_reg_2[155] ));
 sg13g2_dfrbp_1 _1701_ (.CLK(net904),
    .RESET_B(net1057),
    .D(\u_top_module.u_buffer.shift_reg_2[155] ),
    .Q_N(_0670_),
    .Q(\u_top_module.u_buffer.shift_reg_2[156] ));
 sg13g2_dfrbp_1 _1702_ (.CLK(net904),
    .RESET_B(net1058),
    .D(\u_top_module.u_buffer.shift_reg_2[156] ),
    .Q_N(_0671_),
    .Q(\u_top_module.u_buffer.shift_reg_2[157] ));
 sg13g2_dfrbp_1 _1703_ (.CLK(net904),
    .RESET_B(net1058),
    .D(\u_top_module.u_buffer.shift_reg_2[157] ),
    .Q_N(_0672_),
    .Q(\u_top_module.u_buffer.shift_reg_2[158] ));
 sg13g2_dfrbp_1 _1704_ (.CLK(net903),
    .RESET_B(net1058),
    .D(\u_top_module.u_buffer.shift_reg_2[158] ),
    .Q_N(_0673_),
    .Q(\u_top_module.u_buffer.shift_reg_2[159] ));
 sg13g2_dfrbp_1 _1705_ (.CLK(net903),
    .RESET_B(net1058),
    .D(\u_top_module.u_buffer.shift_reg_2[159] ),
    .Q_N(_0674_),
    .Q(\u_top_module.u_buffer.shift_reg_2[160] ));
 sg13g2_dfrbp_1 _1706_ (.CLK(net903),
    .RESET_B(net1057),
    .D(\u_top_module.u_buffer.shift_reg_2[160] ),
    .Q_N(_0675_),
    .Q(\u_top_module.u_buffer.shift_reg_2[161] ));
 sg13g2_dfrbp_1 _1707_ (.CLK(net903),
    .RESET_B(net1057),
    .D(\u_top_module.u_buffer.shift_reg_2[161] ),
    .Q_N(_0676_),
    .Q(\u_top_module.u_buffer.shift_reg_2[162] ));
 sg13g2_dfrbp_1 _1708_ (.CLK(net903),
    .RESET_B(net1057),
    .D(\u_top_module.u_buffer.shift_reg_2[162] ),
    .Q_N(_0677_),
    .Q(\u_top_module.u_buffer.shift_reg_2[163] ));
 sg13g2_dfrbp_1 _1709_ (.CLK(net903),
    .RESET_B(net1057),
    .D(\u_top_module.u_buffer.shift_reg_2[163] ),
    .Q_N(_0678_),
    .Q(\u_top_module.u_buffer.shift_reg_2[164] ));
 sg13g2_dfrbp_1 _1710_ (.CLK(net903),
    .RESET_B(net1057),
    .D(\u_top_module.u_buffer.shift_reg_2[164] ),
    .Q_N(_0679_),
    .Q(\u_top_module.u_buffer.shift_reg_2[165] ));
 sg13g2_dfrbp_1 _1711_ (.CLK(net903),
    .RESET_B(net1057),
    .D(\u_top_module.u_buffer.shift_reg_2[165] ),
    .Q_N(_0680_),
    .Q(\u_top_module.u_buffer.shift_reg_2[166] ));
 sg13g2_dfrbp_1 _1712_ (.CLK(net901),
    .RESET_B(net1055),
    .D(\u_top_module.u_buffer.shift_reg_2[166] ),
    .Q_N(_0681_),
    .Q(\u_top_module.u_buffer.shift_reg_2[167] ));
 sg13g2_dfrbp_1 _1713_ (.CLK(net901),
    .RESET_B(net1055),
    .D(\u_top_module.u_buffer.shift_reg_2[167] ),
    .Q_N(_0682_),
    .Q(\u_top_module.u_buffer.shift_reg_2[168] ));
 sg13g2_dfrbp_1 _1714_ (.CLK(net901),
    .RESET_B(net1055),
    .D(\u_top_module.u_buffer.shift_reg_2[168] ),
    .Q_N(_0683_),
    .Q(\u_top_module.u_buffer.shift_reg_2[169] ));
 sg13g2_dfrbp_1 _1715_ (.CLK(net901),
    .RESET_B(net1055),
    .D(\u_top_module.u_buffer.shift_reg_2[169] ),
    .Q_N(_0684_),
    .Q(\u_top_module.u_buffer.shift_reg_2[170] ));
 sg13g2_dfrbp_1 _1716_ (.CLK(net900),
    .RESET_B(net1054),
    .D(\u_top_module.u_buffer.shift_reg_2[170] ),
    .Q_N(_0685_),
    .Q(\u_top_module.u_buffer.shift_reg_2[171] ));
 sg13g2_dfrbp_1 _1717_ (.CLK(net900),
    .RESET_B(net1054),
    .D(\u_top_module.u_buffer.shift_reg_2[171] ),
    .Q_N(_0686_),
    .Q(\u_top_module.u_buffer.shift_reg_2[172] ));
 sg13g2_dfrbp_1 _1718_ (.CLK(net900),
    .RESET_B(net1054),
    .D(\u_top_module.u_buffer.shift_reg_2[172] ),
    .Q_N(_0687_),
    .Q(\u_top_module.u_buffer.shift_reg_2[173] ));
 sg13g2_dfrbp_1 _1719_ (.CLK(net900),
    .RESET_B(net1054),
    .D(\u_top_module.u_buffer.shift_reg_2[173] ),
    .Q_N(_0688_),
    .Q(\u_top_module.u_buffer.shift_reg_2[174] ));
 sg13g2_dfrbp_1 _1720_ (.CLK(net889),
    .RESET_B(net1044),
    .D(\u_top_module.u_buffer.shift_reg_2[174] ),
    .Q_N(_0689_),
    .Q(\u_top_module.u_buffer.shift_reg_2[175] ));
 sg13g2_dfrbp_1 _1721_ (.CLK(net890),
    .RESET_B(net1044),
    .D(\u_top_module.u_buffer.shift_reg_2[175] ),
    .Q_N(_0690_),
    .Q(\u_top_module.u_buffer.shift_reg_2[176] ));
 sg13g2_dfrbp_1 _1722_ (.CLK(net889),
    .RESET_B(net1045),
    .D(\u_top_module.u_buffer.shift_reg_2[176] ),
    .Q_N(_0691_),
    .Q(\u_top_module.u_buffer.shift_reg_2[177] ));
 sg13g2_dfrbp_1 _1723_ (.CLK(net889),
    .RESET_B(net1044),
    .D(\u_top_module.u_buffer.shift_reg_2[177] ),
    .Q_N(_0692_),
    .Q(\u_top_module.u_buffer.shift_reg_2[178] ));
 sg13g2_dfrbp_1 _1724_ (.CLK(net889),
    .RESET_B(net1044),
    .D(\u_top_module.u_buffer.shift_reg_2[178] ),
    .Q_N(_0693_),
    .Q(\u_top_module.u_buffer.shift_reg_2[179] ));
 sg13g2_dfrbp_1 _1725_ (.CLK(net892),
    .RESET_B(net1047),
    .D(\u_top_module.u_buffer.shift_reg_2[179] ),
    .Q_N(_0694_),
    .Q(\u_top_module.u_buffer.shift_reg_2[180] ));
 sg13g2_dfrbp_1 _1726_ (.CLK(net887),
    .RESET_B(net1042),
    .D(\u_top_module.u_buffer.shift_reg_2[180] ),
    .Q_N(_0695_),
    .Q(\u_top_module.u_buffer.shift_reg_2[181] ));
 sg13g2_dfrbp_1 _1727_ (.CLK(net887),
    .RESET_B(net1042),
    .D(\u_top_module.u_buffer.shift_reg_2[181] ),
    .Q_N(_0696_),
    .Q(\u_top_module.u_buffer.shift_reg_2[182] ));
 sg13g2_dfrbp_1 _1728_ (.CLK(net887),
    .RESET_B(net1043),
    .D(\u_top_module.u_buffer.shift_reg_2[182] ),
    .Q_N(_0697_),
    .Q(\u_top_module.u_buffer.shift_reg_2[183] ));
 sg13g2_dfrbp_1 _1729_ (.CLK(net888),
    .RESET_B(net1043),
    .D(\u_top_module.u_buffer.shift_reg_2[183] ),
    .Q_N(_0698_),
    .Q(\u_top_module.u_buffer.shift_reg_2[184] ));
 sg13g2_dfrbp_1 _1730_ (.CLK(net887),
    .RESET_B(net1042),
    .D(\u_top_module.u_buffer.shift_reg_2[184] ),
    .Q_N(_0699_),
    .Q(\u_top_module.u_buffer.shift_reg_2[185] ));
 sg13g2_dfrbp_1 _1731_ (.CLK(net894),
    .RESET_B(net1049),
    .D(\u_top_module.u_buffer.shift_reg_2[185] ),
    .Q_N(_0700_),
    .Q(\u_top_module.u_buffer.shift_reg_2[186] ));
 sg13g2_dfrbp_1 _1732_ (.CLK(net894),
    .RESET_B(net1049),
    .D(\u_top_module.u_buffer.shift_reg_2[186] ),
    .Q_N(_0701_),
    .Q(\u_top_module.u_buffer.shift_reg_2[187] ));
 sg13g2_dfrbp_1 _1733_ (.CLK(net894),
    .RESET_B(net1049),
    .D(\u_top_module.u_buffer.shift_reg_2[187] ),
    .Q_N(_0702_),
    .Q(\u_top_module.u_buffer.shift_reg_2[188] ));
 sg13g2_dfrbp_1 _1734_ (.CLK(net894),
    .RESET_B(net1049),
    .D(\u_top_module.u_buffer.shift_reg_2[188] ),
    .Q_N(_0703_),
    .Q(\u_top_module.u_buffer.shift_reg_2[189] ));
 sg13g2_dfrbp_1 _1735_ (.CLK(net894),
    .RESET_B(net1049),
    .D(\u_top_module.u_buffer.shift_reg_2[189] ),
    .Q_N(_0704_),
    .Q(\u_top_module.u_buffer.shift_reg_2[190] ));
 sg13g2_dfrbp_1 _1736_ (.CLK(net850),
    .RESET_B(net1004),
    .D(\u_top_module.u_buffer.shift_reg_2[190] ),
    .Q_N(_0705_),
    .Q(\u_top_module.u_buffer.shift_reg_2[191] ));
 sg13g2_dfrbp_1 _1737_ (.CLK(net850),
    .RESET_B(net1004),
    .D(\u_top_module.u_buffer.shift_reg_2[191] ),
    .Q_N(_0706_),
    .Q(\u_top_module.u_buffer.shift_reg_2[192] ));
 sg13g2_dfrbp_1 _1738_ (.CLK(net850),
    .RESET_B(net1004),
    .D(\u_top_module.u_buffer.shift_reg_2[192] ),
    .Q_N(_0707_),
    .Q(\u_top_module.u_buffer.shift_reg_2[193] ));
 sg13g2_dfrbp_1 _1739_ (.CLK(net851),
    .RESET_B(net1006),
    .D(\u_top_module.u_buffer.shift_reg_2[193] ),
    .Q_N(_0708_),
    .Q(\u_top_module.u_buffer.shift_reg_2[194] ));
 sg13g2_dfrbp_1 _1740_ (.CLK(net852),
    .RESET_B(net1006),
    .D(\u_top_module.u_buffer.shift_reg_2[194] ),
    .Q_N(_0709_),
    .Q(\u_top_module.u_buffer.shift_reg_2[195] ));
 sg13g2_dfrbp_1 _1741_ (.CLK(net851),
    .RESET_B(net1005),
    .D(\u_top_module.u_buffer.shift_reg_2[195] ),
    .Q_N(_0710_),
    .Q(\u_top_module.u_buffer.shift_reg_2[196] ));
 sg13g2_dfrbp_1 _1742_ (.CLK(net851),
    .RESET_B(net1005),
    .D(\u_top_module.u_buffer.shift_reg_2[196] ),
    .Q_N(_0711_),
    .Q(\u_top_module.u_buffer.shift_reg_2[197] ));
 sg13g2_dfrbp_1 _1743_ (.CLK(net851),
    .RESET_B(net1005),
    .D(\u_top_module.u_buffer.shift_reg_2[197] ),
    .Q_N(_0712_),
    .Q(\u_top_module.u_buffer.shift_reg_2[198] ));
 sg13g2_dfrbp_1 _1744_ (.CLK(net851),
    .RESET_B(net1005),
    .D(\u_top_module.u_buffer.shift_reg_2[198] ),
    .Q_N(_0713_),
    .Q(\u_top_module.u_buffer.shift_reg_2[199] ));
 sg13g2_dfrbp_1 _1745_ (.CLK(net851),
    .RESET_B(net1005),
    .D(\u_top_module.u_buffer.shift_reg_2[199] ),
    .Q_N(_0714_),
    .Q(\u_top_module.u_buffer.shift_reg_2[200] ));
 sg13g2_dfrbp_1 _1746_ (.CLK(net847),
    .RESET_B(net1002),
    .D(\u_top_module.u_buffer.shift_reg_2[200] ),
    .Q_N(_0715_),
    .Q(\u_top_module.u_buffer.shift_reg_2[201] ));
 sg13g2_dfrbp_1 _1747_ (.CLK(net875),
    .RESET_B(net1002),
    .D(\u_top_module.u_buffer.shift_reg_2[201] ),
    .Q_N(_0716_),
    .Q(\u_top_module.u_buffer.shift_reg_2[202] ));
 sg13g2_dfrbp_1 _1748_ (.CLK(net875),
    .RESET_B(net1027),
    .D(\u_top_module.u_buffer.shift_reg_2[202] ),
    .Q_N(_0717_),
    .Q(\u_top_module.u_buffer.shift_reg_2[203] ));
 sg13g2_dfrbp_1 _1749_ (.CLK(net875),
    .RESET_B(net1027),
    .D(\u_top_module.u_buffer.shift_reg_2[203] ),
    .Q_N(_0718_),
    .Q(\u_top_module.u_buffer.shift_reg_2[204] ));
 sg13g2_dfrbp_1 _1750_ (.CLK(net875),
    .RESET_B(net1027),
    .D(\u_top_module.u_buffer.shift_reg_2[204] ),
    .Q_N(_0719_),
    .Q(\u_top_module.u_buffer.shift_reg_2[205] ));
 sg13g2_dfrbp_1 _1751_ (.CLK(net875),
    .RESET_B(net1027),
    .D(\u_top_module.u_buffer.shift_reg_2[205] ),
    .Q_N(_0720_),
    .Q(\u_top_module.u_buffer.shift_reg_2[206] ));
 sg13g2_dfrbp_1 _1752_ (.CLK(net876),
    .RESET_B(net1027),
    .D(\u_top_module.u_buffer.shift_reg_2[206] ),
    .Q_N(_0721_),
    .Q(\u_top_module.u_buffer.shift_reg_2[207] ));
 sg13g2_dfrbp_1 _1753_ (.CLK(net878),
    .RESET_B(net1028),
    .D(\u_top_module.u_buffer.shift_reg_2[207] ),
    .Q_N(_0722_),
    .Q(\u_top_module.u_buffer.shift_reg_2[208] ));
 sg13g2_dfrbp_1 _1754_ (.CLK(net877),
    .RESET_B(net1028),
    .D(\u_top_module.u_buffer.shift_reg_2[208] ),
    .Q_N(_0723_),
    .Q(\u_top_module.u_buffer.shift_reg_2[209] ));
 sg13g2_dfrbp_1 _1755_ (.CLK(net877),
    .RESET_B(net1029),
    .D(\u_top_module.u_buffer.shift_reg_2[209] ),
    .Q_N(_0724_),
    .Q(\u_top_module.u_buffer.shift_reg_2[210] ));
 sg13g2_dfrbp_1 _1756_ (.CLK(net877),
    .RESET_B(net1029),
    .D(\u_top_module.u_buffer.shift_reg_2[210] ),
    .Q_N(_0725_),
    .Q(\u_top_module.u_buffer.shift_reg_2[211] ));
 sg13g2_dfrbp_1 _1757_ (.CLK(net877),
    .RESET_B(net1029),
    .D(\u_top_module.u_buffer.shift_reg_2[211] ),
    .Q_N(_0726_),
    .Q(\u_top_module.u_buffer.shift_reg_2[212] ));
 sg13g2_dfrbp_1 _1758_ (.CLK(net877),
    .RESET_B(net1029),
    .D(\u_top_module.u_buffer.shift_reg_2[212] ),
    .Q_N(_0727_),
    .Q(\u_top_module.u_buffer.shift_reg_2[213] ));
 sg13g2_dfrbp_1 _1759_ (.CLK(net877),
    .RESET_B(net1029),
    .D(\u_top_module.u_buffer.shift_reg_2[213] ),
    .Q_N(_0728_),
    .Q(\u_top_module.u_buffer.shift_reg_2[214] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(net877),
    .RESET_B(net1029),
    .D(\u_top_module.u_buffer.shift_reg_2[214] ),
    .Q_N(_0729_),
    .Q(\u_top_module.u_buffer.shift_reg_2[215] ));
 sg13g2_dfrbp_1 _1761_ (.CLK(net877),
    .RESET_B(net1029),
    .D(\u_top_module.u_buffer.shift_reg_2[215] ),
    .Q_N(_0730_),
    .Q(\u_top_module.u_buffer.shift_reg_2[216] ));
 sg13g2_dfrbp_1 _1762_ (.CLK(net882),
    .RESET_B(net1029),
    .D(\u_top_module.u_buffer.shift_reg_2[216] ),
    .Q_N(_0731_),
    .Q(\u_top_module.u_buffer.shift_reg_2[217] ));
 sg13g2_dfrbp_1 _1763_ (.CLK(net871),
    .RESET_B(net1016),
    .D(\u_top_module.u_buffer.shift_reg_2[217] ),
    .Q_N(_0732_),
    .Q(\u_top_module.u_buffer.shift_reg_2[218] ));
 sg13g2_dfrbp_1 _1764_ (.CLK(net871),
    .RESET_B(net1022),
    .D(\u_top_module.u_buffer.shift_reg_2[218] ),
    .Q_N(_0733_),
    .Q(\u_top_module.u_buffer.shift_reg_2[219] ));
 sg13g2_dfrbp_1 _1765_ (.CLK(net871),
    .RESET_B(net1022),
    .D(\u_top_module.u_buffer.shift_reg_2[219] ),
    .Q_N(_0734_),
    .Q(\u_top_module.u_buffer.shift_reg_2[220] ));
 sg13g2_dfrbp_1 _1766_ (.CLK(net871),
    .RESET_B(net1022),
    .D(\u_top_module.u_buffer.shift_reg_2[220] ),
    .Q_N(_0735_),
    .Q(\u_top_module.u_buffer.shift_reg_2[221] ));
 sg13g2_dfrbp_1 _1767_ (.CLK(net870),
    .RESET_B(net1022),
    .D(\u_top_module.u_buffer.shift_reg_2[221] ),
    .Q_N(_0736_),
    .Q(\u_top_module.u_buffer.shift_reg_2[222] ));
 sg13g2_dfrbp_1 _1768_ (.CLK(net871),
    .RESET_B(net1022),
    .D(\u_top_module.u_buffer.shift_reg_2[222] ),
    .Q_N(_0737_),
    .Q(\u_top_module.u_buffer.shift_reg_2[223] ));
 sg13g2_dfrbp_1 _1769_ (.CLK(net871),
    .RESET_B(net1023),
    .D(\u_top_module.u_buffer.shift_reg_2[223] ),
    .Q_N(_0738_),
    .Q(\u_top_module.u_buffer.shift_reg_2[224] ));
 sg13g2_dfrbp_1 _1770_ (.CLK(net872),
    .RESET_B(net1022),
    .D(\u_top_module.u_buffer.shift_reg_2[224] ),
    .Q_N(_0739_),
    .Q(\u_top_module.u_buffer.shift_reg_2[225] ));
 sg13g2_dfrbp_1 _1771_ (.CLK(net872),
    .RESET_B(net1022),
    .D(\u_top_module.u_buffer.shift_reg_2[225] ),
    .Q_N(_0740_),
    .Q(\u_top_module.u_buffer.shift_reg_2[226] ));
 sg13g2_dfrbp_1 _1772_ (.CLK(net872),
    .RESET_B(net1022),
    .D(\u_top_module.u_buffer.shift_reg_2[226] ),
    .Q_N(_0741_),
    .Q(\u_top_module.u_buffer.shift_reg_2[227] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(net872),
    .RESET_B(net1025),
    .D(\u_top_module.u_buffer.shift_reg_2[227] ),
    .Q_N(_0742_),
    .Q(\u_top_module.u_buffer.shift_reg_2[228] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(net872),
    .RESET_B(net1025),
    .D(\u_top_module.u_buffer.shift_reg_2[228] ),
    .Q_N(_0743_),
    .Q(\u_top_module.u_buffer.shift_reg_2[229] ));
 sg13g2_dfrbp_1 _1775_ (.CLK(net880),
    .RESET_B(net1034),
    .D(\u_top_module.u_buffer.shift_reg_2[229] ),
    .Q_N(_0744_),
    .Q(\u_top_module.u_buffer.shift_reg_2[230] ));
 sg13g2_dfrbp_1 _1776_ (.CLK(net880),
    .RESET_B(net1034),
    .D(\u_top_module.u_buffer.shift_reg_2[230] ),
    .Q_N(_0745_),
    .Q(\u_top_module.u_buffer.shift_reg_2[231] ));
 sg13g2_dfrbp_1 _1777_ (.CLK(net880),
    .RESET_B(net1034),
    .D(\u_top_module.u_buffer.shift_reg_2[231] ),
    .Q_N(_0746_),
    .Q(\u_top_module.u_buffer.shift_reg_2[232] ));
 sg13g2_dfrbp_1 _1778_ (.CLK(net880),
    .RESET_B(net1036),
    .D(\u_top_module.u_buffer.shift_reg_2[232] ),
    .Q_N(_0747_),
    .Q(\u_top_module.u_buffer.shift_reg_2[233] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(net880),
    .RESET_B(net1036),
    .D(\u_top_module.u_buffer.shift_reg_2[233] ),
    .Q_N(_0748_),
    .Q(\u_top_module.u_buffer.shift_reg_2[234] ));
 sg13g2_dfrbp_1 _1780_ (.CLK(net882),
    .RESET_B(net1036),
    .D(\u_top_module.u_buffer.shift_reg_2[234] ),
    .Q_N(_0749_),
    .Q(\u_top_module.u_buffer.shift_reg_2[235] ));
 sg13g2_dfrbp_1 _1781_ (.CLK(net882),
    .RESET_B(net1036),
    .D(\u_top_module.u_buffer.shift_reg_2[235] ),
    .Q_N(_0750_),
    .Q(\u_top_module.u_buffer.shift_reg_2[236] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(net882),
    .RESET_B(net1036),
    .D(\u_top_module.u_buffer.shift_reg_2[236] ),
    .Q_N(_0751_),
    .Q(\u_top_module.u_buffer.shift_reg_2[237] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(net882),
    .RESET_B(net1036),
    .D(\u_top_module.u_buffer.shift_reg_2[237] ),
    .Q_N(_0752_),
    .Q(\u_top_module.u_buffer.shift_reg_2[238] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(net882),
    .RESET_B(net1036),
    .D(\u_top_module.u_buffer.shift_reg_2[238] ),
    .Q_N(_0753_),
    .Q(\u_top_module.u_buffer.shift_reg_2[239] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(net882),
    .RESET_B(net1030),
    .D(\u_top_module.u_buffer.shift_reg_2[239] ),
    .Q_N(_0754_),
    .Q(\u_top_module.u_buffer.shift_reg_2[240] ));
 sg13g2_dfrbp_1 _1786_ (.CLK(net878),
    .RESET_B(net1030),
    .D(\u_top_module.u_buffer.shift_reg_2[240] ),
    .Q_N(_0755_),
    .Q(\u_top_module.u_buffer.shift_reg_2[241] ));
 sg13g2_dfrbp_1 _1787_ (.CLK(net878),
    .RESET_B(net1030),
    .D(\u_top_module.u_buffer.shift_reg_2[241] ),
    .Q_N(_0756_),
    .Q(\u_top_module.u_buffer.shift_reg_2[242] ));
 sg13g2_dfrbp_1 _1788_ (.CLK(net879),
    .RESET_B(net1033),
    .D(\u_top_module.u_buffer.shift_reg_2[242] ),
    .Q_N(_0757_),
    .Q(\u_top_module.u_buffer.shift_reg_2[243] ));
 sg13g2_dfrbp_1 _1789_ (.CLK(net879),
    .RESET_B(net1033),
    .D(\u_top_module.u_buffer.shift_reg_2[243] ),
    .Q_N(_0758_),
    .Q(\u_top_module.u_buffer.shift_reg_2[244] ));
 sg13g2_dfrbp_1 _1790_ (.CLK(net884),
    .RESET_B(net1033),
    .D(\u_top_module.u_buffer.shift_reg_2[244] ),
    .Q_N(_0759_),
    .Q(\u_top_module.u_buffer.shift_reg_2[245] ));
 sg13g2_dfrbp_1 _1791_ (.CLK(net879),
    .RESET_B(net1033),
    .D(\u_top_module.u_buffer.shift_reg_2[245] ),
    .Q_N(_0760_),
    .Q(\u_top_module.u_buffer.shift_reg_2[246] ));
 sg13g2_dfrbp_1 _1792_ (.CLK(net913),
    .RESET_B(net1069),
    .D(\u_top_module.u_buffer.shift_reg_2[246] ),
    .Q_N(_0761_),
    .Q(\u_top_module.u_buffer.shift_reg_2[247] ));
 sg13g2_dfrbp_1 _1793_ (.CLK(net913),
    .RESET_B(net1069),
    .D(\u_top_module.u_buffer.shift_reg_2[247] ),
    .Q_N(_0762_),
    .Q(\u_top_module.u_buffer.shift_reg_2[248] ));
 sg13g2_dfrbp_1 _1794_ (.CLK(net913),
    .RESET_B(net1069),
    .D(\u_top_module.u_buffer.shift_reg_2[248] ),
    .Q_N(_0763_),
    .Q(\u_top_module.u_buffer.shift_reg_2[249] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(net914),
    .RESET_B(net1073),
    .D(\u_top_module.u_buffer.shift_reg_2[249] ),
    .Q_N(_0764_),
    .Q(\u_top_module.u_buffer.shift_reg_2[250] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(net914),
    .RESET_B(net1073),
    .D(\u_top_module.u_buffer.shift_reg_2[250] ),
    .Q_N(_0765_),
    .Q(\u_top_module.u_buffer.shift_reg_2[251] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(net913),
    .RESET_B(net1073),
    .D(\u_top_module.u_buffer.shift_reg_2[251] ),
    .Q_N(_0766_),
    .Q(\u_top_module.u_buffer.shift_reg_2[252] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(net915),
    .RESET_B(net1078),
    .D(\u_top_module.u_buffer.shift_reg_2[252] ),
    .Q_N(_0767_),
    .Q(\u_top_module.u_buffer.shift_reg_2[253] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(net915),
    .RESET_B(net1078),
    .D(\u_top_module.u_buffer.shift_reg_2[253] ),
    .Q_N(_0768_),
    .Q(\u_top_module.u_buffer.shift_reg_2[254] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(net915),
    .RESET_B(net1078),
    .D(\u_top_module.u_buffer.shift_reg_2[254] ),
    .Q_N(_0612_),
    .Q(\u_top_module.u_buffer.shift_reg_2[255] ));
 sg13g2_dfrbp_1 _1801_ (.CLK(net972),
    .RESET_B(net1085),
    .D(_0027_),
    .Q_N(_0611_),
    .Q(\u_top_module.dec_data_2 ));
 sg13g2_dfrbp_1 _1802_ (.CLK(net969),
    .RESET_B(net1086),
    .D(_0028_),
    .Q_N(_0610_),
    .Q(\u_top_module.u_decimator_1.counter[0] ));
 sg13g2_dfrbp_1 _1803_ (.CLK(net969),
    .RESET_B(net1083),
    .D(_0029_),
    .Q_N(_0609_),
    .Q(\u_top_module.u_decimator_1.counter[1] ));
 sg13g2_dfrbp_1 _1804_ (.CLK(net969),
    .RESET_B(net1083),
    .D(_0030_),
    .Q_N(_0010_),
    .Q(\u_top_module.u_decimator_1.counter[2] ));
 sg13g2_dfrbp_1 _1805_ (.CLK(net969),
    .RESET_B(net1083),
    .D(_0031_),
    .Q_N(_0608_),
    .Q(\u_top_module.u_decimator_1.counter[3] ));
 sg13g2_dfrbp_1 _1806_ (.CLK(net969),
    .RESET_B(net1083),
    .D(_0032_),
    .Q_N(_0013_),
    .Q(\u_top_module.u_decimator_1.counter[4] ));
 sg13g2_dfrbp_1 _1807_ (.CLK(net969),
    .RESET_B(net1083),
    .D(_0033_),
    .Q_N(_0607_),
    .Q(\u_top_module.u_decimator_1.counter[5] ));
 sg13g2_dfrbp_1 _1808_ (.CLK(net971),
    .RESET_B(net1083),
    .D(_0034_),
    .Q_N(_0009_),
    .Q(\u_top_module.u_decimator_1.counter[6] ));
 sg13g2_dfrbp_1 _1809_ (.CLK(net971),
    .RESET_B(net1083),
    .D(_0035_),
    .Q_N(_0011_),
    .Q(\u_top_module.u_decimator_1.counter[7] ));
 sg13g2_dfrbp_1 _1810_ (.CLK(net972),
    .RESET_B(net1085),
    .D(_0036_),
    .Q_N(_0004_),
    .Q(\u_top_module.dec_clk ));
 sg13g2_dfrbp_1 _1811_ (.CLK(net908),
    .RESET_B(net1064),
    .D(_0037_),
    .Q_N(_0015_),
    .Q(\u_top_module.u_buffer.corr_pos[0] ));
 sg13g2_dfrbp_1 _1812_ (.CLK(net907),
    .RESET_B(net1063),
    .D(_0038_),
    .Q_N(_0606_),
    .Q(\u_top_module.u_buffer.corr_pos[1] ));
 sg13g2_dfrbp_1 _1813_ (.CLK(net907),
    .RESET_B(net1062),
    .D(_0039_),
    .Q_N(_0605_),
    .Q(\u_top_module.u_buffer.corr_pos[2] ));
 sg13g2_dfrbp_1 _1814_ (.CLK(net909),
    .RESET_B(net1062),
    .D(_0040_),
    .Q_N(_0604_),
    .Q(\u_top_module.u_buffer.corr_pos[3] ));
 sg13g2_dfrbp_1 _1815_ (.CLK(net909),
    .RESET_B(net1062),
    .D(_0041_),
    .Q_N(_0603_),
    .Q(\u_top_module.u_buffer.corr_pos[4] ));
 sg13g2_dfrbp_1 _1816_ (.CLK(net909),
    .RESET_B(net1062),
    .D(_0042_),
    .Q_N(_0602_),
    .Q(\u_top_module.u_buffer.corr_pos[5] ));
 sg13g2_dfrbp_1 _1817_ (.CLK(net909),
    .RESET_B(net1065),
    .D(_0043_),
    .Q_N(_0601_),
    .Q(\u_top_module.u_buffer.corr_pos[6] ));
 sg13g2_dfrbp_1 _1818_ (.CLK(net909),
    .RESET_B(net1062),
    .D(_0044_),
    .Q_N(_0600_),
    .Q(\u_top_module.u_buffer.corr_pos[7] ));
 sg13g2_dfrbp_1 _1819_ (.CLK(net972),
    .RESET_B(net1085),
    .D(_0045_),
    .Q_N(_0769_),
    .Q(\u_top_module.dec_data_1 ));
 sg13g2_dllrq_1 _1820_ (.D(\u_top_module.mem_out[1] ),
    .GATE_N(_0002_),
    .RESET_B(net17),
    .Q(\u_top_module.filter_length[1] ));
 sg13g2_dllrq_1 _1821_ (.D(\u_top_module.mem_out[2] ),
    .GATE_N(_0002_),
    .RESET_B(net18),
    .Q(\u_top_module.filter_length[2] ));
 sg13g2_dllrq_1 _1822_ (.D(\u_top_module.mem_out[3] ),
    .GATE_N(_0002_),
    .RESET_B(net19),
    .Q(\u_top_module.filter_length[3] ));
 sg13g2_dllrq_1 _1823_ (.D(\u_top_module.mem_out[4] ),
    .GATE_N(_0002_),
    .RESET_B(net20),
    .Q(\u_top_module.filter_length[4] ));
 sg13g2_dllrq_1 _1824_ (.D(\u_top_module.mem_out[5] ),
    .GATE_N(_0002_),
    .RESET_B(net21),
    .Q(\u_top_module.filter_length[5] ));
 sg13g2_dllrq_1 _1825_ (.D(\u_top_module.mem_out[6] ),
    .GATE_N(_0002_),
    .RESET_B(net22),
    .Q(\u_top_module.filter_length[6] ));
 sg13g2_dllrq_1 _1826_ (.D(\u_top_module.mem_out[7] ),
    .GATE_N(_0002_),
    .RESET_B(net23),
    .Q(\u_top_module.filter_length[7] ));
 sg13g2_dllrq_1 _1827_ (.D(\u_top_module.mem_out[0] ),
    .GATE_N(_0001_),
    .RESET_B(net24),
    .Q(\u_top_module.decimation_ratio[0] ));
 sg13g2_dllrq_1 _1828_ (.D(\u_top_module.mem_out[1] ),
    .GATE_N(_0001_),
    .RESET_B(net25),
    .Q(\u_top_module.decimation_ratio[1] ));
 sg13g2_dllrq_1 _1829_ (.D(\u_top_module.mem_out[2] ),
    .GATE_N(_0001_),
    .RESET_B(net26),
    .Q(\u_top_module.decimation_ratio[2] ));
 sg13g2_dllrq_1 _1830_ (.D(\u_top_module.mem_out[3] ),
    .GATE_N(_0001_),
    .RESET_B(net27),
    .Q(\u_top_module.decimation_ratio[3] ));
 sg13g2_dllrq_1 _1831_ (.D(\u_top_module.mem_out[4] ),
    .GATE_N(_0001_),
    .RESET_B(net28),
    .Q(\u_top_module.decimation_ratio[4] ));
 sg13g2_dllrq_1 _1832_ (.D(\u_top_module.mem_out[5] ),
    .GATE_N(_0001_),
    .RESET_B(net29),
    .Q(\u_top_module.decimation_ratio[5] ));
 sg13g2_dllrq_1 _1833_ (.D(\u_top_module.mem_out[6] ),
    .GATE_N(_0001_),
    .RESET_B(net30),
    .Q(\u_top_module.decimation_ratio[6] ));
 sg13g2_dllrq_1 _1834_ (.D(\u_top_module.mem_out[7] ),
    .GATE_N(_0001_),
    .RESET_B(net31),
    .Q(\u_top_module.decimation_ratio[7] ));
 sg13g2_dfrbp_1 _1835_ (.CLK(net973),
    .RESET_B(net32),
    .D(_0158_),
    .Q_N(_0770_),
    .Q(\u_top_module.mem_out[0] ));
 sg13g2_dfrbp_1 _1836_ (.CLK(net961),
    .RESET_B(net33),
    .D(_0159_),
    .Q_N(_0771_),
    .Q(\u_top_module.mem_out[1] ));
 sg13g2_dfrbp_1 _1837_ (.CLK(net963),
    .RESET_B(net34),
    .D(_0160_),
    .Q_N(_0772_),
    .Q(\u_top_module.mem_out[2] ));
 sg13g2_dfrbp_1 _1838_ (.CLK(net963),
    .RESET_B(net35),
    .D(_0161_),
    .Q_N(_0773_),
    .Q(\u_top_module.mem_out[3] ));
 sg13g2_dfrbp_1 _1839_ (.CLK(net961),
    .RESET_B(net36),
    .D(_0162_),
    .Q_N(_0774_),
    .Q(\u_top_module.mem_out[4] ));
 sg13g2_dfrbp_1 _1840_ (.CLK(net963),
    .RESET_B(net37),
    .D(_0163_),
    .Q_N(_0775_),
    .Q(\u_top_module.mem_out[5] ));
 sg13g2_dfrbp_1 _1841_ (.CLK(net962),
    .RESET_B(net39),
    .D(_0164_),
    .Q_N(_0776_),
    .Q(\u_top_module.mem_out[6] ));
 sg13g2_dfrbp_1 _1842_ (.CLK(net973),
    .RESET_B(net38),
    .D(_0165_),
    .Q_N(_0599_),
    .Q(\u_top_module.mem_out[7] ));
 sg13g2_dfrbp_1 _1843_ (.CLK(net970),
    .RESET_B(net1086),
    .D(_0046_),
    .Q_N(_0598_),
    .Q(\u_top_module.u_decimator_2.counter[0] ));
 sg13g2_dfrbp_1 _1844_ (.CLK(net970),
    .RESET_B(net1082),
    .D(_0047_),
    .Q_N(_0597_),
    .Q(\u_top_module.u_decimator_2.counter[1] ));
 sg13g2_dfrbp_1 _1845_ (.CLK(net969),
    .RESET_B(net1082),
    .D(_0048_),
    .Q_N(_0006_),
    .Q(\u_top_module.u_decimator_2.counter[2] ));
 sg13g2_dfrbp_1 _1846_ (.CLK(net970),
    .RESET_B(net1084),
    .D(_0049_),
    .Q_N(_0596_),
    .Q(\u_top_module.u_decimator_2.counter[3] ));
 sg13g2_dfrbp_1 _1847_ (.CLK(net970),
    .RESET_B(net1084),
    .D(_0050_),
    .Q_N(_0012_),
    .Q(\u_top_module.u_decimator_2.counter[4] ));
 sg13g2_dfrbp_1 _1848_ (.CLK(net970),
    .RESET_B(net1083),
    .D(_0051_),
    .Q_N(_0595_),
    .Q(\u_top_module.u_decimator_2.counter[5] ));
 sg13g2_dfrbp_1 _1849_ (.CLK(net971),
    .RESET_B(net1084),
    .D(_0052_),
    .Q_N(_0007_),
    .Q(\u_top_module.u_decimator_2.counter[6] ));
 sg13g2_dfrbp_1 _1850_ (.CLK(net971),
    .RESET_B(net1084),
    .D(_0053_),
    .Q_N(_0008_),
    .Q(\u_top_module.u_decimator_2.counter[7] ));
 sg13g2_dfrbp_1 _1851_ (.CLK(net973),
    .RESET_B(net1082),
    .D(_0054_),
    .Q_N(_0594_),
    .Q(\u_top_module.u_memory.memory[0][0] ));
 sg13g2_dfrbp_1 _1852_ (.CLK(net960),
    .RESET_B(net1075),
    .D(_0055_),
    .Q_N(_0593_),
    .Q(\u_top_module.u_memory.memory[0][1] ));
 sg13g2_dfrbp_1 _1853_ (.CLK(net962),
    .RESET_B(net1076),
    .D(_0056_),
    .Q_N(_0592_),
    .Q(\u_top_module.u_memory.memory[0][2] ));
 sg13g2_dfrbp_1 _1854_ (.CLK(net957),
    .RESET_B(net1071),
    .D(_0057_),
    .Q_N(_0591_),
    .Q(\u_top_module.u_memory.memory[0][3] ));
 sg13g2_dfrbp_1 _1855_ (.CLK(net959),
    .RESET_B(net1075),
    .D(_0058_),
    .Q_N(_0590_),
    .Q(\u_top_module.u_memory.memory[0][4] ));
 sg13g2_dfrbp_1 _1856_ (.CLK(net955),
    .RESET_B(net1070),
    .D(_0059_),
    .Q_N(_0589_),
    .Q(\u_top_module.u_memory.memory[0][5] ));
 sg13g2_dfrbp_1 _1857_ (.CLK(net955),
    .RESET_B(net1070),
    .D(_0060_),
    .Q_N(_0588_),
    .Q(\u_top_module.u_memory.memory[0][6] ));
 sg13g2_dfrbp_1 _1858_ (.CLK(net965),
    .RESET_B(net1072),
    .D(_0061_),
    .Q_N(_0587_),
    .Q(\u_top_module.u_memory.memory[0][7] ));
 sg13g2_dfrbp_1 _1859_ (.CLK(net973),
    .RESET_B(net1082),
    .D(_0062_),
    .Q_N(_0586_),
    .Q(\u_top_module.u_memory.memory[1][0] ));
 sg13g2_dfrbp_1 _1860_ (.CLK(net961),
    .RESET_B(net1077),
    .D(_0063_),
    .Q_N(_0585_),
    .Q(\u_top_module.u_memory.memory[1][1] ));
 sg13g2_dfrbp_1 _1861_ (.CLK(net962),
    .RESET_B(net1076),
    .D(_0064_),
    .Q_N(_0584_),
    .Q(\u_top_module.u_memory.memory[1][2] ));
 sg13g2_dfrbp_1 _1862_ (.CLK(net956),
    .RESET_B(net1071),
    .D(_0065_),
    .Q_N(_0583_),
    .Q(\u_top_module.u_memory.memory[1][3] ));
 sg13g2_dfrbp_1 _1863_ (.CLK(net959),
    .RESET_B(net1037),
    .D(_0066_),
    .Q_N(_0582_),
    .Q(\u_top_module.u_memory.memory[1][4] ));
 sg13g2_dfrbp_1 _1864_ (.CLK(net953),
    .RESET_B(net1032),
    .D(_0067_),
    .Q_N(_0581_),
    .Q(\u_top_module.u_memory.memory[1][5] ));
 sg13g2_dfrbp_1 _1865_ (.CLK(net953),
    .RESET_B(net1031),
    .D(_0068_),
    .Q_N(_0580_),
    .Q(\u_top_module.u_memory.memory[1][6] ));
 sg13g2_dfrbp_1 _1866_ (.CLK(net964),
    .RESET_B(net1072),
    .D(_0069_),
    .Q_N(_0579_),
    .Q(\u_top_module.u_memory.memory[1][7] ));
 sg13g2_dfrbp_1 _1867_ (.CLK(net973),
    .RESET_B(net1082),
    .D(_0070_),
    .Q_N(_0578_),
    .Q(\u_top_module.u_memory.memory[5][0] ));
 sg13g2_dfrbp_1 _1868_ (.CLK(net959),
    .RESET_B(net1075),
    .D(_0071_),
    .Q_N(_0577_),
    .Q(\u_top_module.u_memory.memory[5][1] ));
 sg13g2_dfrbp_1 _1869_ (.CLK(net962),
    .RESET_B(net1076),
    .D(_0072_),
    .Q_N(_0576_),
    .Q(\u_top_module.u_memory.memory[5][2] ));
 sg13g2_dfrbp_1 _1870_ (.CLK(net957),
    .RESET_B(net1071),
    .D(_0073_),
    .Q_N(_0575_),
    .Q(\u_top_module.u_memory.memory[5][3] ));
 sg13g2_dfrbp_1 _1871_ (.CLK(net959),
    .RESET_B(net1037),
    .D(_0074_),
    .Q_N(_0574_),
    .Q(\u_top_module.u_memory.memory[5][4] ));
 sg13g2_dfrbp_1 _1872_ (.CLK(net954),
    .RESET_B(net1032),
    .D(_0075_),
    .Q_N(_0573_),
    .Q(\u_top_module.u_memory.memory[5][5] ));
 sg13g2_dfrbp_1 _1873_ (.CLK(net953),
    .RESET_B(net1031),
    .D(_0076_),
    .Q_N(_0572_),
    .Q(\u_top_module.u_memory.memory[5][6] ));
 sg13g2_dfrbp_1 _1874_ (.CLK(net964),
    .RESET_B(net1072),
    .D(_0077_),
    .Q_N(_0571_),
    .Q(\u_top_module.u_memory.memory[5][7] ));
 sg13g2_dfrbp_1 _1875_ (.CLK(net973),
    .RESET_B(net1082),
    .D(_0078_),
    .Q_N(_0570_),
    .Q(\u_top_module.u_memory.memory[2][0] ));
 sg13g2_dfrbp_1 _1876_ (.CLK(net961),
    .RESET_B(net1077),
    .D(_0079_),
    .Q_N(_0569_),
    .Q(\u_top_module.u_memory.memory[2][1] ));
 sg13g2_dfrbp_1 _1877_ (.CLK(net962),
    .RESET_B(net1076),
    .D(_0080_),
    .Q_N(_0568_),
    .Q(\u_top_module.u_memory.memory[2][2] ));
 sg13g2_dfrbp_1 _1878_ (.CLK(net956),
    .RESET_B(net1071),
    .D(_0081_),
    .Q_N(_0567_),
    .Q(\u_top_module.u_memory.memory[2][3] ));
 sg13g2_dfrbp_1 _1879_ (.CLK(net959),
    .RESET_B(net1037),
    .D(_0082_),
    .Q_N(_0566_),
    .Q(\u_top_module.u_memory.memory[2][4] ));
 sg13g2_dfrbp_1 _1880_ (.CLK(net954),
    .RESET_B(net1032),
    .D(_0083_),
    .Q_N(_0565_),
    .Q(\u_top_module.u_memory.memory[2][5] ));
 sg13g2_dfrbp_1 _1881_ (.CLK(net953),
    .RESET_B(net1031),
    .D(_0084_),
    .Q_N(_0564_),
    .Q(\u_top_module.u_memory.memory[2][6] ));
 sg13g2_dfrbp_1 _1882_ (.CLK(net964),
    .RESET_B(net1072),
    .D(_0085_),
    .Q_N(_0563_),
    .Q(\u_top_module.u_memory.memory[2][7] ));
 sg13g2_dfrbp_1 _1883_ (.CLK(net973),
    .RESET_B(net1082),
    .D(_0086_),
    .Q_N(_0562_),
    .Q(\u_top_module.u_memory.memory[3][0] ));
 sg13g2_dfrbp_1 _1884_ (.CLK(net961),
    .RESET_B(net1075),
    .D(_0087_),
    .Q_N(_0561_),
    .Q(\u_top_module.u_memory.memory[3][1] ));
 sg13g2_dfrbp_1 _1885_ (.CLK(net963),
    .RESET_B(net1076),
    .D(_0088_),
    .Q_N(_0560_),
    .Q(\u_top_module.u_memory.memory[3][2] ));
 sg13g2_dfrbp_1 _1886_ (.CLK(net956),
    .RESET_B(net1071),
    .D(_0089_),
    .Q_N(_0559_),
    .Q(\u_top_module.u_memory.memory[3][3] ));
 sg13g2_dfrbp_1 _1887_ (.CLK(net959),
    .RESET_B(net1037),
    .D(_0090_),
    .Q_N(_0558_),
    .Q(\u_top_module.u_memory.memory[3][4] ));
 sg13g2_dfrbp_1 _1888_ (.CLK(net954),
    .RESET_B(net1031),
    .D(_0091_),
    .Q_N(_0557_),
    .Q(\u_top_module.u_memory.memory[3][5] ));
 sg13g2_dfrbp_1 _1889_ (.CLK(net953),
    .RESET_B(net1031),
    .D(_0092_),
    .Q_N(_0556_),
    .Q(\u_top_module.u_memory.memory[3][6] ));
 sg13g2_dfrbp_1 _1890_ (.CLK(net964),
    .RESET_B(net1072),
    .D(_0093_),
    .Q_N(_0555_),
    .Q(\u_top_module.u_memory.memory[3][7] ));
 sg13g2_dfrbp_1 _1891_ (.CLK(net965),
    .RESET_B(net1079),
    .D(_0094_),
    .Q_N(_0554_),
    .Q(\u_top_module.u_memory.memory[6][0] ));
 sg13g2_dfrbp_1 _1892_ (.CLK(net960),
    .RESET_B(net1075),
    .D(_0095_),
    .Q_N(_0553_),
    .Q(\u_top_module.u_memory.memory[6][1] ));
 sg13g2_dfrbp_1 _1893_ (.CLK(net962),
    .RESET_B(net1076),
    .D(_0096_),
    .Q_N(_0552_),
    .Q(\u_top_module.u_memory.memory[6][2] ));
 sg13g2_dfrbp_1 _1894_ (.CLK(net956),
    .RESET_B(net1071),
    .D(_0097_),
    .Q_N(_0551_),
    .Q(\u_top_module.u_memory.memory[6][3] ));
 sg13g2_dfrbp_1 _1895_ (.CLK(net959),
    .RESET_B(net1037),
    .D(_0098_),
    .Q_N(_0550_),
    .Q(\u_top_module.u_memory.memory[6][4] ));
 sg13g2_dfrbp_1 _1896_ (.CLK(net954),
    .RESET_B(net1032),
    .D(_0099_),
    .Q_N(_0549_),
    .Q(\u_top_module.u_memory.memory[6][5] ));
 sg13g2_dfrbp_1 _1897_ (.CLK(net953),
    .RESET_B(net1031),
    .D(_0100_),
    .Q_N(_0548_),
    .Q(\u_top_module.u_memory.memory[6][6] ));
 sg13g2_dfrbp_1 _1898_ (.CLK(net964),
    .RESET_B(net1079),
    .D(_0101_),
    .Q_N(_0547_),
    .Q(\u_top_module.u_memory.memory[6][7] ));
 sg13g2_dfrbp_1 _1899_ (.CLK(net964),
    .RESET_B(net1079),
    .D(_0102_),
    .Q_N(_0546_),
    .Q(\u_top_module.u_memory.memory[4][0] ));
 sg13g2_dfrbp_1 _1900_ (.CLK(net961),
    .RESET_B(net1075),
    .D(_0103_),
    .Q_N(_0545_),
    .Q(\u_top_module.u_memory.memory[4][1] ));
 sg13g2_dfrbp_1 _1901_ (.CLK(net963),
    .RESET_B(net1077),
    .D(_0104_),
    .Q_N(_0544_),
    .Q(\u_top_module.u_memory.memory[4][2] ));
 sg13g2_dfrbp_1 _1902_ (.CLK(net956),
    .RESET_B(net1071),
    .D(_0105_),
    .Q_N(_0543_),
    .Q(\u_top_module.u_memory.memory[4][3] ));
 sg13g2_dfrbp_1 _1903_ (.CLK(net960),
    .RESET_B(net1037),
    .D(_0106_),
    .Q_N(_0542_),
    .Q(\u_top_module.u_memory.memory[4][4] ));
 sg13g2_dfrbp_1 _1904_ (.CLK(net954),
    .RESET_B(net1032),
    .D(_0107_),
    .Q_N(_0541_),
    .Q(\u_top_module.u_memory.memory[4][5] ));
 sg13g2_dfrbp_1 _1905_ (.CLK(net953),
    .RESET_B(net1031),
    .D(_0108_),
    .Q_N(_0540_),
    .Q(\u_top_module.u_memory.memory[4][6] ));
 sg13g2_dfrbp_1 _1906_ (.CLK(net964),
    .RESET_B(net1072),
    .D(_0109_),
    .Q_N(_0539_),
    .Q(\u_top_module.u_memory.memory[4][7] ));
 sg13g2_dfrbp_1 _1907_ (.CLK(net972),
    .RESET_B(net1085),
    .D(_0026_),
    .Q_N(\u_top_module.u_spi_port.cs_n_prev ),
    .Q(_0017_));
 sg13g2_dfrbp_1 _1908_ (.CLK(net972),
    .RESET_B(net1085),
    .D(_0110_),
    .Q_N(_0538_),
    .Q(\u_top_module.capture_reg[0] ));
 sg13g2_dfrbp_1 _1909_ (.CLK(net960),
    .RESET_B(net1075),
    .D(_0111_),
    .Q_N(_0537_),
    .Q(\u_top_module.capture_reg[1] ));
 sg13g2_dfrbp_1 _1910_ (.CLK(net962),
    .RESET_B(net1076),
    .D(_0112_),
    .Q_N(_0536_),
    .Q(\u_top_module.capture_reg[2] ));
 sg13g2_dfrbp_1 _1911_ (.CLK(net956),
    .RESET_B(net1070),
    .D(_0113_),
    .Q_N(_0535_),
    .Q(\u_top_module.capture_reg[3] ));
 sg13g2_dfrbp_1 _1912_ (.CLK(net960),
    .RESET_B(net1075),
    .D(_0114_),
    .Q_N(_0534_),
    .Q(\u_top_module.capture_reg[4] ));
 sg13g2_dfrbp_1 _1913_ (.CLK(net955),
    .RESET_B(net1070),
    .D(_0115_),
    .Q_N(_0533_),
    .Q(\u_top_module.capture_reg[5] ));
 sg13g2_dfrbp_1 _1914_ (.CLK(net955),
    .RESET_B(net1070),
    .D(_0116_),
    .Q_N(_0532_),
    .Q(\u_top_module.capture_reg[6] ));
 sg13g2_dfrbp_1 _1915_ (.CLK(net958),
    .RESET_B(net1073),
    .D(_0117_),
    .Q_N(_0531_),
    .Q(\u_top_module.capture_reg[7] ));
 sg13g2_dfrbp_1 _1916_ (.CLK(net965),
    .RESET_B(net1079),
    .D(_0118_),
    .Q_N(_0530_),
    .Q(\u_top_module.addr[0] ));
 sg13g2_dfrbp_1 _1917_ (.CLK(net965),
    .RESET_B(net1078),
    .D(_0119_),
    .Q_N(_0529_),
    .Q(\u_top_module.addr[1] ));
 sg13g2_dfrbp_1 _1918_ (.CLK(net965),
    .RESET_B(net1079),
    .D(_0120_),
    .Q_N(_0005_),
    .Q(\u_top_module.addr[2] ));
 sg13g2_dfrbp_1 _1919_ (.CLK(net965),
    .RESET_B(net1079),
    .D(_0121_),
    .Q_N(_0528_),
    .Q(\u_top_module.addr[3] ));
 sg13g2_dfrbp_1 _1920_ (.CLK(net966),
    .RESET_B(net1080),
    .D(_0122_),
    .Q_N(_0527_),
    .Q(\u_top_module.addr[4] ));
 sg13g2_dfrbp_1 _1921_ (.CLK(net966),
    .RESET_B(net1080),
    .D(_0123_),
    .Q_N(_0526_),
    .Q(\u_top_module.addr[5] ));
 sg13g2_dfrbp_1 _1922_ (.CLK(net966),
    .RESET_B(net1080),
    .D(_0124_),
    .Q_N(_0525_),
    .Q(\u_top_module.addr[6] ));
 sg13g2_dfrbp_1 _1923_ (.CLK(net966),
    .RESET_B(net1080),
    .D(_0125_),
    .Q_N(_0524_),
    .Q(\u_top_module.addr[7] ));
 sg13g2_dfrbp_1 _1924_ (.CLK(net973),
    .RESET_B(net1082),
    .D(_0126_),
    .Q_N(_0523_),
    .Q(\u_top_module.u_memory.memory[7][0] ));
 sg13g2_dfrbp_1 _1925_ (.CLK(net961),
    .RESET_B(net1077),
    .D(_0127_),
    .Q_N(_0522_),
    .Q(\u_top_module.u_memory.memory[7][1] ));
 sg13g2_dfrbp_1 _1926_ (.CLK(net962),
    .RESET_B(net1076),
    .D(_0128_),
    .Q_N(_0521_),
    .Q(\u_top_module.u_memory.memory[7][2] ));
 sg13g2_dfrbp_1 _1927_ (.CLK(net957),
    .RESET_B(net1071),
    .D(_0129_),
    .Q_N(_0520_),
    .Q(\u_top_module.u_memory.memory[7][3] ));
 sg13g2_dfrbp_1 _1928_ (.CLK(net959),
    .RESET_B(net1037),
    .D(_0130_),
    .Q_N(_0519_),
    .Q(\u_top_module.u_memory.memory[7][4] ));
 sg13g2_dfrbp_1 _1929_ (.CLK(net954),
    .RESET_B(net1032),
    .D(_0131_),
    .Q_N(_0518_),
    .Q(\u_top_module.u_memory.memory[7][5] ));
 sg13g2_dfrbp_1 _1930_ (.CLK(net953),
    .RESET_B(net1031),
    .D(_0132_),
    .Q_N(_0517_),
    .Q(\u_top_module.u_memory.memory[7][6] ));
 sg13g2_dfrbp_1 _1931_ (.CLK(net964),
    .RESET_B(net1072),
    .D(_0133_),
    .Q_N(_0516_),
    .Q(\u_top_module.u_memory.memory[7][7] ));
 sg13g2_dfrbp_1 _1932_ (.CLK(net972),
    .RESET_B(net1085),
    .D(_0134_),
    .Q_N(_0515_),
    .Q(\u_top_module.u_spi_port.shift_reg[0] ));
 sg13g2_dfrbp_1 _1933_ (.CLK(net966),
    .RESET_B(net1085),
    .D(_0135_),
    .Q_N(_0514_),
    .Q(\u_top_module.u_spi_port.shift_reg[1] ));
 sg13g2_dfrbp_1 _1934_ (.CLK(net956),
    .RESET_B(net1069),
    .D(_0136_),
    .Q_N(_0513_),
    .Q(\u_top_module.u_spi_port.shift_reg[2] ));
 sg13g2_dfrbp_1 _1935_ (.CLK(net956),
    .RESET_B(net1070),
    .D(_0137_),
    .Q_N(_0512_),
    .Q(\u_top_module.u_spi_port.shift_reg[3] ));
 sg13g2_dfrbp_1 _1936_ (.CLK(net955),
    .RESET_B(net1070),
    .D(_0138_),
    .Q_N(_0511_),
    .Q(\u_top_module.u_spi_port.shift_reg[4] ));
 sg13g2_dfrbp_1 _1937_ (.CLK(net958),
    .RESET_B(net1069),
    .D(_0139_),
    .Q_N(_0510_),
    .Q(\u_top_module.u_spi_port.shift_reg[5] ));
 sg13g2_dfrbp_1 _1938_ (.CLK(net958),
    .RESET_B(net1069),
    .D(_0140_),
    .Q_N(_0509_),
    .Q(\u_top_module.u_spi_port.shift_reg[6] ));
 sg13g2_dfrbp_1 _1939_ (.CLK(net958),
    .RESET_B(net1073),
    .D(_0141_),
    .Q_N(_0508_),
    .Q(\u_top_module.u_spi_port.shift_reg[7] ));
 sg13g2_dfrbp_1 _1940_ (.CLK(net968),
    .RESET_B(net1078),
    .D(_0142_),
    .Q_N(_0507_),
    .Q(\u_top_module.u_spi_port.shift_reg[8] ));
 sg13g2_dfrbp_1 _1941_ (.CLK(net968),
    .RESET_B(net1078),
    .D(_0143_),
    .Q_N(_0506_),
    .Q(\u_top_module.u_spi_port.shift_reg[9] ));
 sg13g2_dfrbp_1 _1942_ (.CLK(net965),
    .RESET_B(net1079),
    .D(_0144_),
    .Q_N(_0505_),
    .Q(\u_top_module.u_spi_port.shift_reg[10] ));
 sg13g2_dfrbp_1 _1943_ (.CLK(net966),
    .RESET_B(net1080),
    .D(_0145_),
    .Q_N(_0504_),
    .Q(\u_top_module.u_spi_port.shift_reg[11] ));
 sg13g2_dfrbp_1 _1944_ (.CLK(net966),
    .RESET_B(net1080),
    .D(_0146_),
    .Q_N(_0503_),
    .Q(\u_top_module.u_spi_port.shift_reg[12] ));
 sg13g2_dfrbp_1 _1945_ (.CLK(net967),
    .RESET_B(net1081),
    .D(_0147_),
    .Q_N(_0502_),
    .Q(\u_top_module.u_spi_port.shift_reg[13] ));
 sg13g2_dfrbp_1 _1946_ (.CLK(net967),
    .RESET_B(net1080),
    .D(_0148_),
    .Q_N(_0501_),
    .Q(\u_top_module.u_spi_port.shift_reg[14] ));
 sg13g2_dfrbp_1 _1947_ (.CLK(net966),
    .RESET_B(net1080),
    .D(_0149_),
    .Q_N(_0500_),
    .Q(\u_top_module.u_spi_port.shift_reg[15] ));
 sg13g2_dfrbp_1 _1948_ (.CLK(net907),
    .RESET_B(net1064),
    .D(_0150_),
    .Q_N(_0016_),
    .Q(\u_top_module.u_buffer.corr_neg[0] ));
 sg13g2_dfrbp_1 _1949_ (.CLK(net908),
    .RESET_B(net1064),
    .D(_0151_),
    .Q_N(_0499_),
    .Q(\u_top_module.u_buffer.corr_neg[1] ));
 sg13g2_dfrbp_1 _1950_ (.CLK(net908),
    .RESET_B(net1064),
    .D(_0152_),
    .Q_N(_0498_),
    .Q(\u_top_module.u_buffer.corr_neg[2] ));
 sg13g2_dfrbp_1 _1951_ (.CLK(net908),
    .RESET_B(net1062),
    .D(_0153_),
    .Q_N(_0497_),
    .Q(\u_top_module.u_buffer.corr_neg[3] ));
 sg13g2_dfrbp_1 _1952_ (.CLK(net910),
    .RESET_B(net1066),
    .D(_0154_),
    .Q_N(_0496_),
    .Q(\u_top_module.u_buffer.corr_neg[4] ));
 sg13g2_dfrbp_1 _1953_ (.CLK(net910),
    .RESET_B(net1066),
    .D(_0155_),
    .Q_N(_0495_),
    .Q(\u_top_module.u_buffer.corr_neg[5] ));
 sg13g2_dfrbp_1 _1954_ (.CLK(net909),
    .RESET_B(net1062),
    .D(_0156_),
    .Q_N(_0494_),
    .Q(\u_top_module.u_buffer.corr_neg[6] ));
 sg13g2_dfrbp_1 _1955_ (.CLK(net909),
    .RESET_B(net1062),
    .D(_0157_),
    .Q_N(_0777_),
    .Q(\u_top_module.u_buffer.corr_neg[7] ));
 sg13g2_dfrbp_1 _1956_ (.CLK(net911),
    .RESET_B(net1066),
    .D(_0003_),
    .Q_N(_0778_),
    .Q(\u_top_module.pos ));
 sg13g2_dfrbp_1 _1957_ (.CLK(net915),
    .RESET_B(net1063),
    .D(\u_top_module.dec_data_1 ),
    .Q_N(_0779_),
    .Q(\u_top_module.u_buffer.shift_reg_1[0] ));
 sg13g2_dfrbp_1 _1958_ (.CLK(net907),
    .RESET_B(net1063),
    .D(\u_top_module.u_buffer.shift_reg_1[0] ),
    .Q_N(_0780_),
    .Q(\u_top_module.u_buffer.shift_reg_1[1] ));
 sg13g2_dfrbp_1 _1959_ (.CLK(net907),
    .RESET_B(net1063),
    .D(\u_top_module.u_buffer.shift_reg_1[1] ),
    .Q_N(_0781_),
    .Q(\u_top_module.u_buffer.shift_reg_1[2] ));
 sg13g2_dfrbp_1 _1960_ (.CLK(net907),
    .RESET_B(net1063),
    .D(\u_top_module.u_buffer.shift_reg_1[2] ),
    .Q_N(_0782_),
    .Q(\u_top_module.u_buffer.shift_reg_1[3] ));
 sg13g2_dfrbp_1 _1961_ (.CLK(net898),
    .RESET_B(net1052),
    .D(\u_top_module.u_buffer.shift_reg_1[3] ),
    .Q_N(_0783_),
    .Q(\u_top_module.u_buffer.shift_reg_1[4] ));
 sg13g2_dfrbp_1 _1962_ (.CLK(net898),
    .RESET_B(net1052),
    .D(\u_top_module.u_buffer.shift_reg_1[4] ),
    .Q_N(_0784_),
    .Q(\u_top_module.u_buffer.shift_reg_1[5] ));
 sg13g2_dfrbp_1 _1963_ (.CLK(net898),
    .RESET_B(net1052),
    .D(\u_top_module.u_buffer.shift_reg_1[5] ),
    .Q_N(_0785_),
    .Q(\u_top_module.u_buffer.shift_reg_1[6] ));
 sg13g2_dfrbp_1 _1964_ (.CLK(net898),
    .RESET_B(net1052),
    .D(\u_top_module.u_buffer.shift_reg_1[6] ),
    .Q_N(_0786_),
    .Q(\u_top_module.u_buffer.shift_reg_1[7] ));
 sg13g2_dfrbp_1 _1965_ (.CLK(net898),
    .RESET_B(net1052),
    .D(\u_top_module.u_buffer.shift_reg_1[7] ),
    .Q_N(_0787_),
    .Q(\u_top_module.u_buffer.shift_reg_1[8] ));
 sg13g2_dfrbp_1 _1966_ (.CLK(net896),
    .RESET_B(net1050),
    .D(\u_top_module.u_buffer.shift_reg_1[8] ),
    .Q_N(_0788_),
    .Q(\u_top_module.u_buffer.shift_reg_1[9] ));
 sg13g2_dfrbp_1 _1967_ (.CLK(net896),
    .RESET_B(net1051),
    .D(\u_top_module.u_buffer.shift_reg_1[9] ),
    .Q_N(_0789_),
    .Q(\u_top_module.u_buffer.shift_reg_1[10] ));
 sg13g2_dfrbp_1 _1968_ (.CLK(net896),
    .RESET_B(net1050),
    .D(\u_top_module.u_buffer.shift_reg_1[10] ),
    .Q_N(_0790_),
    .Q(\u_top_module.u_buffer.shift_reg_1[11] ));
 sg13g2_dfrbp_1 _1969_ (.CLK(net896),
    .RESET_B(net1050),
    .D(\u_top_module.u_buffer.shift_reg_1[11] ),
    .Q_N(_0791_),
    .Q(\u_top_module.u_buffer.shift_reg_1[12] ));
 sg13g2_dfrbp_1 _1970_ (.CLK(net879),
    .RESET_B(net1005),
    .D(\u_top_module.u_buffer.shift_reg_1[12] ),
    .Q_N(_0792_),
    .Q(\u_top_module.u_buffer.shift_reg_1[13] ));
 sg13g2_dfrbp_1 _1971_ (.CLK(net879),
    .RESET_B(net1005),
    .D(\u_top_module.u_buffer.shift_reg_1[13] ),
    .Q_N(_0793_),
    .Q(\u_top_module.u_buffer.shift_reg_1[14] ));
 sg13g2_dfrbp_1 _1972_ (.CLK(net879),
    .RESET_B(net1033),
    .D(\u_top_module.u_buffer.shift_reg_1[14] ),
    .Q_N(_0794_),
    .Q(\u_top_module.u_buffer.shift_reg_1[15] ));
 sg13g2_dfrbp_1 _1973_ (.CLK(net879),
    .RESET_B(net1033),
    .D(\u_top_module.u_buffer.shift_reg_1[15] ),
    .Q_N(_0795_),
    .Q(\u_top_module.u_buffer.shift_reg_1[16] ));
 sg13g2_dfrbp_1 _1974_ (.CLK(net875),
    .RESET_B(net1027),
    .D(\u_top_module.u_buffer.shift_reg_1[16] ),
    .Q_N(_0796_),
    .Q(\u_top_module.u_buffer.shift_reg_1[17] ));
 sg13g2_dfrbp_1 _1975_ (.CLK(net875),
    .RESET_B(net1027),
    .D(\u_top_module.u_buffer.shift_reg_1[17] ),
    .Q_N(_0797_),
    .Q(\u_top_module.u_buffer.shift_reg_1[18] ));
 sg13g2_dfrbp_1 _1976_ (.CLK(net875),
    .RESET_B(net1027),
    .D(\u_top_module.u_buffer.shift_reg_1[18] ),
    .Q_N(_0798_),
    .Q(\u_top_module.u_buffer.shift_reg_1[19] ));
 sg13g2_dfrbp_1 _1977_ (.CLK(net876),
    .RESET_B(net1028),
    .D(\u_top_module.u_buffer.shift_reg_1[19] ),
    .Q_N(_0799_),
    .Q(\u_top_module.u_buffer.shift_reg_1[20] ));
 sg13g2_dfrbp_1 _1978_ (.CLK(net876),
    .RESET_B(net1028),
    .D(\u_top_module.u_buffer.shift_reg_1[20] ),
    .Q_N(_0800_),
    .Q(\u_top_module.u_buffer.shift_reg_1[21] ));
 sg13g2_dfrbp_1 _1979_ (.CLK(net876),
    .RESET_B(net1028),
    .D(\u_top_module.u_buffer.shift_reg_1[21] ),
    .Q_N(_0801_),
    .Q(\u_top_module.u_buffer.shift_reg_1[22] ));
 sg13g2_dfrbp_1 _1980_ (.CLK(net860),
    .RESET_B(net1014),
    .D(\u_top_module.u_buffer.shift_reg_1[22] ),
    .Q_N(_0802_),
    .Q(\u_top_module.u_buffer.shift_reg_1[23] ));
 sg13g2_dfrbp_1 _1981_ (.CLK(net860),
    .RESET_B(net1014),
    .D(\u_top_module.u_buffer.shift_reg_1[23] ),
    .Q_N(_0803_),
    .Q(\u_top_module.u_buffer.shift_reg_1[24] ));
 sg13g2_dfrbp_1 _1982_ (.CLK(net863),
    .RESET_B(net1014),
    .D(\u_top_module.u_buffer.shift_reg_1[24] ),
    .Q_N(_0804_),
    .Q(\u_top_module.u_buffer.shift_reg_1[25] ));
 sg13g2_dfrbp_1 _1983_ (.CLK(net863),
    .RESET_B(net1016),
    .D(\u_top_module.u_buffer.shift_reg_1[25] ),
    .Q_N(_0805_),
    .Q(\u_top_module.u_buffer.shift_reg_1[26] ));
 sg13g2_dfrbp_1 _1984_ (.CLK(net863),
    .RESET_B(net1016),
    .D(\u_top_module.u_buffer.shift_reg_1[26] ),
    .Q_N(_0806_),
    .Q(\u_top_module.u_buffer.shift_reg_1[27] ));
 sg13g2_dfrbp_1 _1985_ (.CLK(net863),
    .RESET_B(net1016),
    .D(\u_top_module.u_buffer.shift_reg_1[27] ),
    .Q_N(_0807_),
    .Q(\u_top_module.u_buffer.shift_reg_1[28] ));
 sg13g2_dfrbp_1 _1986_ (.CLK(net862),
    .RESET_B(net1015),
    .D(\u_top_module.u_buffer.shift_reg_1[28] ),
    .Q_N(_0808_),
    .Q(\u_top_module.u_buffer.shift_reg_1[29] ));
 sg13g2_dfrbp_1 _1987_ (.CLK(net862),
    .RESET_B(net1015),
    .D(\u_top_module.u_buffer.shift_reg_1[29] ),
    .Q_N(_0809_),
    .Q(\u_top_module.u_buffer.shift_reg_1[30] ));
 sg13g2_dfrbp_1 _1988_ (.CLK(net862),
    .RESET_B(net1015),
    .D(\u_top_module.u_buffer.shift_reg_1[30] ),
    .Q_N(_0810_),
    .Q(\u_top_module.u_buffer.shift_reg_1[31] ));
 sg13g2_dfrbp_1 _1989_ (.CLK(net858),
    .RESET_B(net1011),
    .D(\u_top_module.u_buffer.shift_reg_1[31] ),
    .Q_N(_0811_),
    .Q(\u_top_module.u_buffer.shift_reg_1[32] ));
 sg13g2_dfrbp_1 _1990_ (.CLK(net857),
    .RESET_B(net1011),
    .D(\u_top_module.u_buffer.shift_reg_1[32] ),
    .Q_N(_0812_),
    .Q(\u_top_module.u_buffer.shift_reg_1[33] ));
 sg13g2_dfrbp_1 _1991_ (.CLK(net857),
    .RESET_B(net1011),
    .D(\u_top_module.u_buffer.shift_reg_1[33] ),
    .Q_N(_0813_),
    .Q(\u_top_module.u_buffer.shift_reg_1[34] ));
 sg13g2_dfrbp_1 _1992_ (.CLK(net857),
    .RESET_B(net1011),
    .D(\u_top_module.u_buffer.shift_reg_1[34] ),
    .Q_N(_0814_),
    .Q(\u_top_module.u_buffer.shift_reg_1[35] ));
 sg13g2_dfrbp_1 _1993_ (.CLK(net857),
    .RESET_B(net1011),
    .D(\u_top_module.u_buffer.shift_reg_1[35] ),
    .Q_N(_0815_),
    .Q(\u_top_module.u_buffer.shift_reg_1[36] ));
 sg13g2_dfrbp_1 _1994_ (.CLK(net859),
    .RESET_B(net1011),
    .D(\u_top_module.u_buffer.shift_reg_1[36] ),
    .Q_N(_0816_),
    .Q(\u_top_module.u_buffer.shift_reg_1[37] ));
 sg13g2_dfrbp_1 _1995_ (.CLK(net859),
    .RESET_B(net1013),
    .D(\u_top_module.u_buffer.shift_reg_1[37] ),
    .Q_N(_0817_),
    .Q(\u_top_module.u_buffer.shift_reg_1[38] ));
 sg13g2_dfrbp_1 _1996_ (.CLK(net858),
    .RESET_B(net1012),
    .D(\u_top_module.u_buffer.shift_reg_1[38] ),
    .Q_N(_0818_),
    .Q(\u_top_module.u_buffer.shift_reg_1[39] ));
 sg13g2_dfrbp_1 _1997_ (.CLK(net859),
    .RESET_B(net1012),
    .D(\u_top_module.u_buffer.shift_reg_1[39] ),
    .Q_N(_0819_),
    .Q(\u_top_module.u_buffer.shift_reg_1[40] ));
 sg13g2_dfrbp_1 _1998_ (.CLK(net859),
    .RESET_B(net1013),
    .D(\u_top_module.u_buffer.shift_reg_1[40] ),
    .Q_N(_0820_),
    .Q(\u_top_module.u_buffer.shift_reg_1[41] ));
 sg13g2_dfrbp_1 _1999_ (.CLK(net859),
    .RESET_B(net1013),
    .D(\u_top_module.u_buffer.shift_reg_1[41] ),
    .Q_N(_0821_),
    .Q(\u_top_module.u_buffer.shift_reg_1[42] ));
 sg13g2_dfrbp_1 _2000_ (.CLK(net867),
    .RESET_B(net1013),
    .D(\u_top_module.u_buffer.shift_reg_1[42] ),
    .Q_N(_0822_),
    .Q(\u_top_module.u_buffer.shift_reg_1[43] ));
 sg13g2_dfrbp_1 _2001_ (.CLK(net867),
    .RESET_B(net1013),
    .D(\u_top_module.u_buffer.shift_reg_1[43] ),
    .Q_N(_0823_),
    .Q(\u_top_module.u_buffer.shift_reg_1[44] ));
 sg13g2_dfrbp_1 _2002_ (.CLK(net866),
    .RESET_B(net1019),
    .D(\u_top_module.u_buffer.shift_reg_1[44] ),
    .Q_N(_0824_),
    .Q(\u_top_module.u_buffer.shift_reg_1[45] ));
 sg13g2_dfrbp_1 _2003_ (.CLK(net866),
    .RESET_B(net1019),
    .D(\u_top_module.u_buffer.shift_reg_1[45] ),
    .Q_N(_0825_),
    .Q(\u_top_module.u_buffer.shift_reg_1[46] ));
 sg13g2_dfrbp_1 _2004_ (.CLK(net867),
    .RESET_B(net1019),
    .D(\u_top_module.u_buffer.shift_reg_1[46] ),
    .Q_N(_0826_),
    .Q(\u_top_module.u_buffer.shift_reg_1[47] ));
 sg13g2_dfrbp_1 _2005_ (.CLK(net867),
    .RESET_B(net1019),
    .D(\u_top_module.u_buffer.shift_reg_1[47] ),
    .Q_N(_0827_),
    .Q(\u_top_module.u_buffer.shift_reg_1[48] ));
 sg13g2_dfrbp_1 _2006_ (.CLK(net866),
    .RESET_B(net1019),
    .D(\u_top_module.u_buffer.shift_reg_1[48] ),
    .Q_N(_0828_),
    .Q(\u_top_module.u_buffer.shift_reg_1[49] ));
 sg13g2_dfrbp_1 _2007_ (.CLK(net867),
    .RESET_B(net1020),
    .D(\u_top_module.u_buffer.shift_reg_1[49] ),
    .Q_N(_0829_),
    .Q(\u_top_module.u_buffer.shift_reg_1[50] ));
 sg13g2_dfrbp_1 _2008_ (.CLK(net866),
    .RESET_B(net1020),
    .D(\u_top_module.u_buffer.shift_reg_1[50] ),
    .Q_N(_0830_),
    .Q(\u_top_module.u_buffer.shift_reg_1[51] ));
 sg13g2_dfrbp_1 _2009_ (.CLK(net866),
    .RESET_B(net1019),
    .D(\u_top_module.u_buffer.shift_reg_1[51] ),
    .Q_N(_0831_),
    .Q(\u_top_module.u_buffer.shift_reg_1[52] ));
 sg13g2_dfrbp_1 _2010_ (.CLK(net866),
    .RESET_B(net1019),
    .D(\u_top_module.u_buffer.shift_reg_1[52] ),
    .Q_N(_0832_),
    .Q(\u_top_module.u_buffer.shift_reg_1[53] ));
 sg13g2_dfrbp_1 _2011_ (.CLK(net866),
    .RESET_B(net1019),
    .D(\u_top_module.u_buffer.shift_reg_1[53] ),
    .Q_N(_0833_),
    .Q(\u_top_module.u_buffer.shift_reg_1[54] ));
 sg13g2_dfrbp_1 _2012_ (.CLK(net866),
    .RESET_B(net1012),
    .D(\u_top_module.u_buffer.shift_reg_1[54] ),
    .Q_N(_0834_),
    .Q(\u_top_module.u_buffer.shift_reg_1[55] ));
 sg13g2_dfrbp_1 _2013_ (.CLK(net858),
    .RESET_B(net1012),
    .D(\u_top_module.u_buffer.shift_reg_1[55] ),
    .Q_N(_0835_),
    .Q(\u_top_module.u_buffer.shift_reg_1[56] ));
 sg13g2_dfrbp_1 _2014_ (.CLK(net858),
    .RESET_B(net1012),
    .D(\u_top_module.u_buffer.shift_reg_1[56] ),
    .Q_N(_0836_),
    .Q(\u_top_module.u_buffer.shift_reg_1[57] ));
 sg13g2_dfrbp_1 _2015_ (.CLK(net858),
    .RESET_B(net1012),
    .D(\u_top_module.u_buffer.shift_reg_1[57] ),
    .Q_N(_0837_),
    .Q(\u_top_module.u_buffer.shift_reg_1[58] ));
 sg13g2_dfrbp_1 _2016_ (.CLK(net858),
    .RESET_B(net1012),
    .D(\u_top_module.u_buffer.shift_reg_1[58] ),
    .Q_N(_0838_),
    .Q(\u_top_module.u_buffer.shift_reg_1[59] ));
 sg13g2_dfrbp_1 _2017_ (.CLK(net858),
    .RESET_B(net1012),
    .D(\u_top_module.u_buffer.shift_reg_1[59] ),
    .Q_N(_0839_),
    .Q(\u_top_module.u_buffer.shift_reg_1[60] ));
 sg13g2_dfrbp_1 _2018_ (.CLK(net858),
    .RESET_B(net1010),
    .D(\u_top_module.u_buffer.shift_reg_1[60] ),
    .Q_N(_0840_),
    .Q(\u_top_module.u_buffer.shift_reg_1[61] ));
 sg13g2_dfrbp_1 _2019_ (.CLK(net856),
    .RESET_B(net1010),
    .D(\u_top_module.u_buffer.shift_reg_1[61] ),
    .Q_N(_0841_),
    .Q(\u_top_module.u_buffer.shift_reg_1[62] ));
 sg13g2_dfrbp_1 _2020_ (.CLK(net856),
    .RESET_B(net1010),
    .D(\u_top_module.u_buffer.shift_reg_1[62] ),
    .Q_N(_0842_),
    .Q(\u_top_module.u_buffer.shift_reg_1[63] ));
 sg13g2_dfrbp_1 _2021_ (.CLK(net856),
    .RESET_B(net1011),
    .D(\u_top_module.u_buffer.shift_reg_1[63] ),
    .Q_N(_0843_),
    .Q(\u_top_module.u_buffer.shift_reg_1[64] ));
 sg13g2_dfrbp_1 _2022_ (.CLK(net857),
    .RESET_B(net1010),
    .D(\u_top_module.u_buffer.shift_reg_1[64] ),
    .Q_N(_0844_),
    .Q(\u_top_module.u_buffer.shift_reg_1[65] ));
 sg13g2_dfrbp_1 _2023_ (.CLK(net857),
    .RESET_B(net1010),
    .D(\u_top_module.u_buffer.shift_reg_1[65] ),
    .Q_N(_0845_),
    .Q(\u_top_module.u_buffer.shift_reg_1[66] ));
 sg13g2_dfrbp_1 _2024_ (.CLK(net856),
    .RESET_B(net1010),
    .D(\u_top_module.u_buffer.shift_reg_1[66] ),
    .Q_N(_0846_),
    .Q(\u_top_module.u_buffer.shift_reg_1[67] ));
 sg13g2_dfrbp_1 _2025_ (.CLK(net856),
    .RESET_B(net1010),
    .D(\u_top_module.u_buffer.shift_reg_1[67] ),
    .Q_N(_0847_),
    .Q(\u_top_module.u_buffer.shift_reg_1[68] ));
 sg13g2_dfrbp_1 _2026_ (.CLK(net856),
    .RESET_B(net1010),
    .D(\u_top_module.u_buffer.shift_reg_1[68] ),
    .Q_N(_0848_),
    .Q(\u_top_module.u_buffer.shift_reg_1[69] ));
 sg13g2_dfrbp_1 _2027_ (.CLK(net856),
    .RESET_B(net985),
    .D(\u_top_module.u_buffer.shift_reg_1[69] ),
    .Q_N(_0849_),
    .Q(\u_top_module.u_buffer.shift_reg_1[70] ));
 sg13g2_dfrbp_1 _2028_ (.CLK(net856),
    .RESET_B(net985),
    .D(\u_top_module.u_buffer.shift_reg_1[70] ),
    .Q_N(_0850_),
    .Q(\u_top_module.u_buffer.shift_reg_1[71] ));
 sg13g2_dfrbp_1 _2029_ (.CLK(net832),
    .RESET_B(net986),
    .D(\u_top_module.u_buffer.shift_reg_1[71] ),
    .Q_N(_0851_),
    .Q(\u_top_module.u_buffer.shift_reg_1[72] ));
 sg13g2_dfrbp_1 _2030_ (.CLK(net832),
    .RESET_B(net985),
    .D(\u_top_module.u_buffer.shift_reg_1[72] ),
    .Q_N(_0852_),
    .Q(\u_top_module.u_buffer.shift_reg_1[73] ));
 sg13g2_dfrbp_1 _2031_ (.CLK(net832),
    .RESET_B(net985),
    .D(\u_top_module.u_buffer.shift_reg_1[73] ),
    .Q_N(_0853_),
    .Q(\u_top_module.u_buffer.shift_reg_1[74] ));
 sg13g2_dfrbp_1 _2032_ (.CLK(net832),
    .RESET_B(net985),
    .D(\u_top_module.u_buffer.shift_reg_1[74] ),
    .Q_N(_0854_),
    .Q(\u_top_module.u_buffer.shift_reg_1[75] ));
 sg13g2_dfrbp_1 _2033_ (.CLK(net832),
    .RESET_B(net985),
    .D(\u_top_module.u_buffer.shift_reg_1[75] ),
    .Q_N(_0855_),
    .Q(\u_top_module.u_buffer.shift_reg_1[76] ));
 sg13g2_dfrbp_1 _2034_ (.CLK(net832),
    .RESET_B(net985),
    .D(\u_top_module.u_buffer.shift_reg_1[76] ),
    .Q_N(_0856_),
    .Q(\u_top_module.u_buffer.shift_reg_1[77] ));
 sg13g2_dfrbp_1 _2035_ (.CLK(net832),
    .RESET_B(net985),
    .D(\u_top_module.u_buffer.shift_reg_1[77] ),
    .Q_N(_0857_),
    .Q(\u_top_module.u_buffer.shift_reg_1[78] ));
 sg13g2_dfrbp_1 _2036_ (.CLK(net832),
    .RESET_B(net983),
    .D(\u_top_module.u_buffer.shift_reg_1[78] ),
    .Q_N(_0858_),
    .Q(\u_top_module.u_buffer.shift_reg_1[79] ));
 sg13g2_dfrbp_1 _2037_ (.CLK(net831),
    .RESET_B(net984),
    .D(\u_top_module.u_buffer.shift_reg_1[79] ),
    .Q_N(_0859_),
    .Q(\u_top_module.u_buffer.shift_reg_1[80] ));
 sg13g2_dfrbp_1 _2038_ (.CLK(net830),
    .RESET_B(net984),
    .D(\u_top_module.u_buffer.shift_reg_1[80] ),
    .Q_N(_0860_),
    .Q(\u_top_module.u_buffer.shift_reg_1[81] ));
 sg13g2_dfrbp_1 _2039_ (.CLK(net831),
    .RESET_B(net983),
    .D(\u_top_module.u_buffer.shift_reg_1[81] ),
    .Q_N(_0861_),
    .Q(\u_top_module.u_buffer.shift_reg_1[82] ));
 sg13g2_dfrbp_1 _2040_ (.CLK(net830),
    .RESET_B(net983),
    .D(\u_top_module.u_buffer.shift_reg_1[82] ),
    .Q_N(_0862_),
    .Q(\u_top_module.u_buffer.shift_reg_1[83] ));
 sg13g2_dfrbp_1 _2041_ (.CLK(net830),
    .RESET_B(net983),
    .D(\u_top_module.u_buffer.shift_reg_1[83] ),
    .Q_N(_0863_),
    .Q(\u_top_module.u_buffer.shift_reg_1[84] ));
 sg13g2_dfrbp_1 _2042_ (.CLK(net830),
    .RESET_B(net983),
    .D(\u_top_module.u_buffer.shift_reg_1[84] ),
    .Q_N(_0864_),
    .Q(\u_top_module.u_buffer.shift_reg_1[85] ));
 sg13g2_dfrbp_1 _2043_ (.CLK(net830),
    .RESET_B(net983),
    .D(\u_top_module.u_buffer.shift_reg_1[85] ),
    .Q_N(_0865_),
    .Q(\u_top_module.u_buffer.shift_reg_1[86] ));
 sg13g2_dfrbp_1 _2044_ (.CLK(net830),
    .RESET_B(net983),
    .D(\u_top_module.u_buffer.shift_reg_1[86] ),
    .Q_N(_0866_),
    .Q(\u_top_module.u_buffer.shift_reg_1[87] ));
 sg13g2_dfrbp_1 _2045_ (.CLK(net830),
    .RESET_B(net983),
    .D(\u_top_module.u_buffer.shift_reg_1[87] ),
    .Q_N(_0867_),
    .Q(\u_top_module.u_buffer.shift_reg_1[88] ));
 sg13g2_dfrbp_1 _2046_ (.CLK(net830),
    .RESET_B(net977),
    .D(\u_top_module.u_buffer.shift_reg_1[88] ),
    .Q_N(_0868_),
    .Q(\u_top_module.u_buffer.shift_reg_1[89] ));
 sg13g2_dfrbp_1 _2047_ (.CLK(net824),
    .RESET_B(net977),
    .D(\u_top_module.u_buffer.shift_reg_1[89] ),
    .Q_N(_0869_),
    .Q(\u_top_module.u_buffer.shift_reg_1[90] ));
 sg13g2_dfrbp_1 _2048_ (.CLK(net824),
    .RESET_B(net977),
    .D(\u_top_module.u_buffer.shift_reg_1[90] ),
    .Q_N(_0870_),
    .Q(\u_top_module.u_buffer.shift_reg_1[91] ));
 sg13g2_dfrbp_1 _2049_ (.CLK(net825),
    .RESET_B(net978),
    .D(\u_top_module.u_buffer.shift_reg_1[91] ),
    .Q_N(_0871_),
    .Q(\u_top_module.u_buffer.shift_reg_1[92] ));
 sg13g2_dfrbp_1 _2050_ (.CLK(net825),
    .RESET_B(net978),
    .D(\u_top_module.u_buffer.shift_reg_1[92] ),
    .Q_N(_0872_),
    .Q(\u_top_module.u_buffer.shift_reg_1[93] ));
 sg13g2_dfrbp_1 _2051_ (.CLK(net825),
    .RESET_B(net978),
    .D(\u_top_module.u_buffer.shift_reg_1[93] ),
    .Q_N(_0873_),
    .Q(\u_top_module.u_buffer.shift_reg_1[94] ));
 sg13g2_dfrbp_1 _2052_ (.CLK(net825),
    .RESET_B(net978),
    .D(\u_top_module.u_buffer.shift_reg_1[94] ),
    .Q_N(_0874_),
    .Q(\u_top_module.u_buffer.shift_reg_1[95] ));
 sg13g2_dfrbp_1 _2053_ (.CLK(net824),
    .RESET_B(net978),
    .D(\u_top_module.u_buffer.shift_reg_1[95] ),
    .Q_N(_0875_),
    .Q(\u_top_module.u_buffer.shift_reg_1[96] ));
 sg13g2_dfrbp_1 _2054_ (.CLK(net824),
    .RESET_B(net977),
    .D(\u_top_module.u_buffer.shift_reg_1[96] ),
    .Q_N(_0876_),
    .Q(\u_top_module.u_buffer.shift_reg_1[97] ));
 sg13g2_dfrbp_1 _2055_ (.CLK(net824),
    .RESET_B(net977),
    .D(\u_top_module.u_buffer.shift_reg_1[97] ),
    .Q_N(_0877_),
    .Q(\u_top_module.u_buffer.shift_reg_1[98] ));
 sg13g2_dfrbp_1 _2056_ (.CLK(net824),
    .RESET_B(net977),
    .D(\u_top_module.u_buffer.shift_reg_1[98] ),
    .Q_N(_0878_),
    .Q(\u_top_module.u_buffer.shift_reg_1[99] ));
 sg13g2_dfrbp_1 _2057_ (.CLK(net824),
    .RESET_B(net977),
    .D(\u_top_module.u_buffer.shift_reg_1[99] ),
    .Q_N(_0879_),
    .Q(\u_top_module.u_buffer.shift_reg_1[100] ));
 sg13g2_dfrbp_1 _2058_ (.CLK(net822),
    .RESET_B(net975),
    .D(\u_top_module.u_buffer.shift_reg_1[100] ),
    .Q_N(_0880_),
    .Q(\u_top_module.u_buffer.shift_reg_1[101] ));
 sg13g2_dfrbp_1 _2059_ (.CLK(net822),
    .RESET_B(net975),
    .D(\u_top_module.u_buffer.shift_reg_1[101] ),
    .Q_N(_0881_),
    .Q(\u_top_module.u_buffer.shift_reg_1[102] ));
 sg13g2_dfrbp_1 _2060_ (.CLK(net822),
    .RESET_B(net975),
    .D(\u_top_module.u_buffer.shift_reg_1[102] ),
    .Q_N(_0882_),
    .Q(\u_top_module.u_buffer.shift_reg_1[103] ));
 sg13g2_dfrbp_1 _2061_ (.CLK(net822),
    .RESET_B(net975),
    .D(\u_top_module.u_buffer.shift_reg_1[103] ),
    .Q_N(_0883_),
    .Q(\u_top_module.u_buffer.shift_reg_1[104] ));
 sg13g2_dfrbp_1 _2062_ (.CLK(net822),
    .RESET_B(net975),
    .D(\u_top_module.u_buffer.shift_reg_1[104] ),
    .Q_N(_0884_),
    .Q(\u_top_module.u_buffer.shift_reg_1[105] ));
 sg13g2_dfrbp_1 _2063_ (.CLK(net822),
    .RESET_B(net975),
    .D(\u_top_module.u_buffer.shift_reg_1[105] ),
    .Q_N(_0885_),
    .Q(\u_top_module.u_buffer.shift_reg_1[106] ));
 sg13g2_dfrbp_1 _2064_ (.CLK(net822),
    .RESET_B(net975),
    .D(\u_top_module.u_buffer.shift_reg_1[106] ),
    .Q_N(_0886_),
    .Q(\u_top_module.u_buffer.shift_reg_1[107] ));
 sg13g2_dfrbp_1 _2065_ (.CLK(net823),
    .RESET_B(net975),
    .D(\u_top_module.u_buffer.shift_reg_1[107] ),
    .Q_N(_0887_),
    .Q(\u_top_module.u_buffer.shift_reg_1[108] ));
 sg13g2_dfrbp_1 _2066_ (.CLK(net823),
    .RESET_B(net976),
    .D(\u_top_module.u_buffer.shift_reg_1[108] ),
    .Q_N(_0888_),
    .Q(\u_top_module.u_buffer.shift_reg_1[109] ));
 sg13g2_dfrbp_1 _2067_ (.CLK(net822),
    .RESET_B(net976),
    .D(\u_top_module.u_buffer.shift_reg_1[109] ),
    .Q_N(_0889_),
    .Q(\u_top_module.u_buffer.shift_reg_1[110] ));
 sg13g2_dfrbp_1 _2068_ (.CLK(net823),
    .RESET_B(net976),
    .D(\u_top_module.u_buffer.shift_reg_1[110] ),
    .Q_N(_0890_),
    .Q(\u_top_module.u_buffer.shift_reg_1[111] ));
 sg13g2_dfrbp_1 _2069_ (.CLK(net823),
    .RESET_B(net976),
    .D(\u_top_module.u_buffer.shift_reg_1[111] ),
    .Q_N(_0891_),
    .Q(\u_top_module.u_buffer.shift_reg_1[112] ));
 sg13g2_dfrbp_1 _2070_ (.CLK(net827),
    .RESET_B(net980),
    .D(\u_top_module.u_buffer.shift_reg_1[112] ),
    .Q_N(_0892_),
    .Q(\u_top_module.u_buffer.shift_reg_1[113] ));
 sg13g2_dfrbp_1 _2071_ (.CLK(net827),
    .RESET_B(net980),
    .D(\u_top_module.u_buffer.shift_reg_1[113] ),
    .Q_N(_0893_),
    .Q(\u_top_module.u_buffer.shift_reg_1[114] ));
 sg13g2_dfrbp_1 _2072_ (.CLK(net827),
    .RESET_B(net980),
    .D(\u_top_module.u_buffer.shift_reg_1[114] ),
    .Q_N(_0894_),
    .Q(\u_top_module.u_buffer.shift_reg_1[115] ));
 sg13g2_dfrbp_1 _2073_ (.CLK(net827),
    .RESET_B(net980),
    .D(\u_top_module.u_buffer.shift_reg_1[115] ),
    .Q_N(_0895_),
    .Q(\u_top_module.u_buffer.shift_reg_1[116] ));
 sg13g2_dfrbp_1 _2074_ (.CLK(net827),
    .RESET_B(net980),
    .D(\u_top_module.u_buffer.shift_reg_1[116] ),
    .Q_N(_0896_),
    .Q(\u_top_module.u_buffer.shift_reg_1[117] ));
 sg13g2_dfrbp_1 _2075_ (.CLK(net827),
    .RESET_B(net980),
    .D(\u_top_module.u_buffer.shift_reg_1[117] ),
    .Q_N(_0897_),
    .Q(\u_top_module.u_buffer.shift_reg_1[118] ));
 sg13g2_dfrbp_1 _2076_ (.CLK(net827),
    .RESET_B(net981),
    .D(\u_top_module.u_buffer.shift_reg_1[118] ),
    .Q_N(_0898_),
    .Q(\u_top_module.u_buffer.shift_reg_1[119] ));
 sg13g2_dfrbp_1 _2077_ (.CLK(net828),
    .RESET_B(net981),
    .D(\u_top_module.u_buffer.shift_reg_1[119] ),
    .Q_N(_0899_),
    .Q(\u_top_module.u_buffer.shift_reg_1[120] ));
 sg13g2_dfrbp_1 _2078_ (.CLK(net828),
    .RESET_B(net981),
    .D(\u_top_module.u_buffer.shift_reg_1[120] ),
    .Q_N(_0900_),
    .Q(\u_top_module.u_buffer.shift_reg_1[121] ));
 sg13g2_dfrbp_1 _2079_ (.CLK(net828),
    .RESET_B(net980),
    .D(\u_top_module.u_buffer.shift_reg_1[121] ),
    .Q_N(_0901_),
    .Q(\u_top_module.u_buffer.shift_reg_1[122] ));
 sg13g2_dfrbp_1 _2080_ (.CLK(net827),
    .RESET_B(net980),
    .D(\u_top_module.u_buffer.shift_reg_1[122] ),
    .Q_N(_0902_),
    .Q(\u_top_module.u_buffer.shift_reg_1[123] ));
 sg13g2_dfrbp_1 _2081_ (.CLK(net839),
    .RESET_B(net993),
    .D(\u_top_module.u_buffer.shift_reg_1[123] ),
    .Q_N(_0903_),
    .Q(\u_top_module.u_buffer.shift_reg_1[124] ));
 sg13g2_dfrbp_1 _2082_ (.CLK(net839),
    .RESET_B(net993),
    .D(\u_top_module.u_buffer.shift_reg_1[124] ),
    .Q_N(_0904_),
    .Q(\u_top_module.u_buffer.shift_reg_1[125] ));
 sg13g2_dfrbp_1 _2083_ (.CLK(net839),
    .RESET_B(net993),
    .D(\u_top_module.u_buffer.shift_reg_1[125] ),
    .Q_N(_0905_),
    .Q(\u_top_module.u_buffer.shift_reg_1[126] ));
 sg13g2_dfrbp_1 _2084_ (.CLK(net839),
    .RESET_B(net993),
    .D(\u_top_module.u_buffer.shift_reg_1[126] ),
    .Q_N(_0906_),
    .Q(\u_top_module.u_buffer.shift_reg_1[127] ));
 sg13g2_dfrbp_1 _2085_ (.CLK(net839),
    .RESET_B(net993),
    .D(\u_top_module.u_buffer.shift_reg_1[127] ),
    .Q_N(_0907_),
    .Q(\u_top_module.u_buffer.shift_reg_1[128] ));
 sg13g2_dfrbp_1 _2086_ (.CLK(net841),
    .RESET_B(net994),
    .D(\u_top_module.u_buffer.shift_reg_1[128] ),
    .Q_N(_0908_),
    .Q(\u_top_module.u_buffer.shift_reg_1[129] ));
 sg13g2_dfrbp_1 _2087_ (.CLK(net840),
    .RESET_B(net994),
    .D(\u_top_module.u_buffer.shift_reg_1[129] ),
    .Q_N(_0909_),
    .Q(\u_top_module.u_buffer.shift_reg_1[130] ));
 sg13g2_dfrbp_1 _2088_ (.CLK(net840),
    .RESET_B(net994),
    .D(\u_top_module.u_buffer.shift_reg_1[130] ),
    .Q_N(_0910_),
    .Q(\u_top_module.u_buffer.shift_reg_1[131] ));
 sg13g2_dfrbp_1 _2089_ (.CLK(net840),
    .RESET_B(net995),
    .D(\u_top_module.u_buffer.shift_reg_1[131] ),
    .Q_N(_0911_),
    .Q(\u_top_module.u_buffer.shift_reg_1[132] ));
 sg13g2_dfrbp_1 _2090_ (.CLK(net854),
    .RESET_B(net1008),
    .D(\u_top_module.u_buffer.shift_reg_1[132] ),
    .Q_N(_0912_),
    .Q(\u_top_module.u_buffer.shift_reg_1[133] ));
 sg13g2_dfrbp_1 _2091_ (.CLK(net843),
    .RESET_B(net997),
    .D(\u_top_module.u_buffer.shift_reg_1[133] ),
    .Q_N(_0913_),
    .Q(\u_top_module.u_buffer.shift_reg_1[134] ));
 sg13g2_dfrbp_1 _2092_ (.CLK(net843),
    .RESET_B(net997),
    .D(\u_top_module.u_buffer.shift_reg_1[134] ),
    .Q_N(_0914_),
    .Q(\u_top_module.u_buffer.shift_reg_1[135] ));
 sg13g2_dfrbp_1 _2093_ (.CLK(net843),
    .RESET_B(net997),
    .D(\u_top_module.u_buffer.shift_reg_1[135] ),
    .Q_N(_0915_),
    .Q(\u_top_module.u_buffer.shift_reg_1[136] ));
 sg13g2_dfrbp_1 _2094_ (.CLK(net843),
    .RESET_B(net997),
    .D(\u_top_module.u_buffer.shift_reg_1[136] ),
    .Q_N(_0916_),
    .Q(\u_top_module.u_buffer.shift_reg_1[137] ));
 sg13g2_dfrbp_1 _2095_ (.CLK(net843),
    .RESET_B(net997),
    .D(\u_top_module.u_buffer.shift_reg_1[137] ),
    .Q_N(_0917_),
    .Q(\u_top_module.u_buffer.shift_reg_1[138] ));
 sg13g2_dfrbp_1 _2096_ (.CLK(net844),
    .RESET_B(net998),
    .D(\u_top_module.u_buffer.shift_reg_1[138] ),
    .Q_N(_0918_),
    .Q(\u_top_module.u_buffer.shift_reg_1[139] ));
 sg13g2_dfrbp_1 _2097_ (.CLK(net844),
    .RESET_B(net998),
    .D(\u_top_module.u_buffer.shift_reg_1[139] ),
    .Q_N(_0919_),
    .Q(\u_top_module.u_buffer.shift_reg_1[140] ));
 sg13g2_dfrbp_1 _2098_ (.CLK(net844),
    .RESET_B(net998),
    .D(\u_top_module.u_buffer.shift_reg_1[140] ),
    .Q_N(_0920_),
    .Q(\u_top_module.u_buffer.shift_reg_1[141] ));
 sg13g2_dfrbp_1 _2099_ (.CLK(net844),
    .RESET_B(net998),
    .D(\u_top_module.u_buffer.shift_reg_1[141] ),
    .Q_N(_0921_),
    .Q(\u_top_module.u_buffer.shift_reg_1[142] ));
 sg13g2_dfrbp_1 _2100_ (.CLK(net887),
    .RESET_B(net1041),
    .D(\u_top_module.u_buffer.shift_reg_1[142] ),
    .Q_N(_0922_),
    .Q(\u_top_module.u_buffer.shift_reg_1[143] ));
 sg13g2_dfrbp_1 _2101_ (.CLK(net885),
    .RESET_B(net1040),
    .D(\u_top_module.u_buffer.shift_reg_1[143] ),
    .Q_N(_0923_),
    .Q(\u_top_module.u_buffer.shift_reg_1[144] ));
 sg13g2_dfrbp_1 _2102_ (.CLK(net885),
    .RESET_B(net1040),
    .D(\u_top_module.u_buffer.shift_reg_1[144] ),
    .Q_N(_0924_),
    .Q(\u_top_module.u_buffer.shift_reg_1[145] ));
 sg13g2_dfrbp_1 _2103_ (.CLK(net885),
    .RESET_B(net1040),
    .D(\u_top_module.u_buffer.shift_reg_1[145] ),
    .Q_N(_0925_),
    .Q(\u_top_module.u_buffer.shift_reg_1[146] ));
 sg13g2_dfrbp_1 _2104_ (.CLK(net885),
    .RESET_B(net1040),
    .D(\u_top_module.u_buffer.shift_reg_1[146] ),
    .Q_N(_0926_),
    .Q(\u_top_module.u_buffer.shift_reg_1[147] ));
 sg13g2_dfrbp_1 _2105_ (.CLK(net886),
    .RESET_B(net1041),
    .D(\u_top_module.u_buffer.shift_reg_1[147] ),
    .Q_N(_0927_),
    .Q(\u_top_module.u_buffer.shift_reg_1[148] ));
 sg13g2_dfrbp_1 _2106_ (.CLK(net886),
    .RESET_B(net1041),
    .D(\u_top_module.u_buffer.shift_reg_1[148] ),
    .Q_N(_0928_),
    .Q(\u_top_module.u_buffer.shift_reg_1[149] ));
 sg13g2_dfrbp_1 _2107_ (.CLK(net886),
    .RESET_B(net1041),
    .D(\u_top_module.u_buffer.shift_reg_1[149] ),
    .Q_N(_0929_),
    .Q(\u_top_module.u_buffer.shift_reg_1[150] ));
 sg13g2_dfrbp_1 _2108_ (.CLK(net886),
    .RESET_B(net1041),
    .D(\u_top_module.u_buffer.shift_reg_1[150] ),
    .Q_N(_0930_),
    .Q(\u_top_module.u_buffer.shift_reg_1[151] ));
 sg13g2_dfrbp_1 _2109_ (.CLK(net889),
    .RESET_B(net1044),
    .D(\u_top_module.u_buffer.shift_reg_1[151] ),
    .Q_N(_0931_),
    .Q(\u_top_module.u_buffer.shift_reg_1[152] ));
 sg13g2_dfrbp_1 _2110_ (.CLK(net892),
    .RESET_B(net1047),
    .D(\u_top_module.u_buffer.shift_reg_1[152] ),
    .Q_N(_0932_),
    .Q(\u_top_module.u_buffer.shift_reg_1[153] ));
 sg13g2_dfrbp_1 _2111_ (.CLK(net892),
    .RESET_B(net1047),
    .D(\u_top_module.u_buffer.shift_reg_1[153] ),
    .Q_N(_0933_),
    .Q(\u_top_module.u_buffer.shift_reg_1[154] ));
 sg13g2_dfrbp_1 _2112_ (.CLK(net892),
    .RESET_B(net1047),
    .D(\u_top_module.u_buffer.shift_reg_1[154] ),
    .Q_N(_0934_),
    .Q(\u_top_module.u_buffer.shift_reg_1[155] ));
 sg13g2_dfrbp_1 _2113_ (.CLK(net891),
    .RESET_B(net1046),
    .D(\u_top_module.u_buffer.shift_reg_1[155] ),
    .Q_N(_0935_),
    .Q(\u_top_module.u_buffer.shift_reg_1[156] ));
 sg13g2_dfrbp_1 _2114_ (.CLK(net891),
    .RESET_B(net1046),
    .D(\u_top_module.u_buffer.shift_reg_1[156] ),
    .Q_N(_0936_),
    .Q(\u_top_module.u_buffer.shift_reg_1[157] ));
 sg13g2_dfrbp_1 _2115_ (.CLK(net891),
    .RESET_B(net1046),
    .D(\u_top_module.u_buffer.shift_reg_1[157] ),
    .Q_N(_0937_),
    .Q(\u_top_module.u_buffer.shift_reg_1[158] ));
 sg13g2_dfrbp_1 _2116_ (.CLK(net891),
    .RESET_B(net1046),
    .D(\u_top_module.u_buffer.shift_reg_1[158] ),
    .Q_N(_0938_),
    .Q(\u_top_module.u_buffer.shift_reg_1[159] ));
 sg13g2_dfrbp_1 _2117_ (.CLK(net891),
    .RESET_B(net1046),
    .D(\u_top_module.u_buffer.shift_reg_1[159] ),
    .Q_N(_0939_),
    .Q(\u_top_module.u_buffer.shift_reg_1[160] ));
 sg13g2_dfrbp_1 _2118_ (.CLK(net892),
    .RESET_B(net1047),
    .D(\u_top_module.u_buffer.shift_reg_1[160] ),
    .Q_N(_0940_),
    .Q(\u_top_module.u_buffer.shift_reg_1[161] ));
 sg13g2_dfrbp_1 _2119_ (.CLK(net891),
    .RESET_B(net1046),
    .D(\u_top_module.u_buffer.shift_reg_1[161] ),
    .Q_N(_0941_),
    .Q(\u_top_module.u_buffer.shift_reg_1[162] ));
 sg13g2_dfrbp_1 _2120_ (.CLK(net891),
    .RESET_B(net1046),
    .D(\u_top_module.u_buffer.shift_reg_1[162] ),
    .Q_N(_0942_),
    .Q(\u_top_module.u_buffer.shift_reg_1[163] ));
 sg13g2_dfrbp_1 _2121_ (.CLK(net891),
    .RESET_B(net1046),
    .D(\u_top_module.u_buffer.shift_reg_1[163] ),
    .Q_N(_0943_),
    .Q(\u_top_module.u_buffer.shift_reg_1[164] ));
 sg13g2_dfrbp_1 _2122_ (.CLK(net892),
    .RESET_B(net1047),
    .D(\u_top_module.u_buffer.shift_reg_1[164] ),
    .Q_N(_0944_),
    .Q(\u_top_module.u_buffer.shift_reg_1[165] ));
 sg13g2_dfrbp_1 _2123_ (.CLK(net899),
    .RESET_B(net1047),
    .D(\u_top_module.u_buffer.shift_reg_1[165] ),
    .Q_N(_0945_),
    .Q(\u_top_module.u_buffer.shift_reg_1[166] ));
 sg13g2_dfrbp_1 _2124_ (.CLK(net899),
    .RESET_B(net1053),
    .D(\u_top_module.u_buffer.shift_reg_1[166] ),
    .Q_N(_0946_),
    .Q(\u_top_module.u_buffer.shift_reg_1[167] ));
 sg13g2_dfrbp_1 _2125_ (.CLK(net899),
    .RESET_B(net1053),
    .D(\u_top_module.u_buffer.shift_reg_1[167] ),
    .Q_N(_0947_),
    .Q(\u_top_module.u_buffer.shift_reg_1[168] ));
 sg13g2_dfrbp_1 _2126_ (.CLK(net894),
    .RESET_B(net1049),
    .D(\u_top_module.u_buffer.shift_reg_1[168] ),
    .Q_N(_0948_),
    .Q(\u_top_module.u_buffer.shift_reg_1[169] ));
 sg13g2_dfrbp_1 _2127_ (.CLK(net894),
    .RESET_B(net1042),
    .D(\u_top_module.u_buffer.shift_reg_1[169] ),
    .Q_N(_0949_),
    .Q(\u_top_module.u_buffer.shift_reg_1[170] ));
 sg13g2_dfrbp_1 _2128_ (.CLK(net894),
    .RESET_B(net1042),
    .D(\u_top_module.u_buffer.shift_reg_1[170] ),
    .Q_N(_0950_),
    .Q(\u_top_module.u_buffer.shift_reg_1[171] ));
 sg13g2_dfrbp_1 _2129_ (.CLK(net887),
    .RESET_B(net1042),
    .D(\u_top_module.u_buffer.shift_reg_1[171] ),
    .Q_N(_0951_),
    .Q(\u_top_module.u_buffer.shift_reg_1[172] ));
 sg13g2_dfrbp_1 _2130_ (.CLK(net887),
    .RESET_B(net1042),
    .D(\u_top_module.u_buffer.shift_reg_1[172] ),
    .Q_N(_0952_),
    .Q(\u_top_module.u_buffer.shift_reg_1[173] ));
 sg13g2_dfrbp_1 _2131_ (.CLK(net887),
    .RESET_B(net1042),
    .D(\u_top_module.u_buffer.shift_reg_1[173] ),
    .Q_N(_0953_),
    .Q(\u_top_module.u_buffer.shift_reg_1[174] ));
 sg13g2_dfrbp_1 _2132_ (.CLK(net843),
    .RESET_B(net997),
    .D(\u_top_module.u_buffer.shift_reg_1[174] ),
    .Q_N(_0954_),
    .Q(\u_top_module.u_buffer.shift_reg_1[175] ));
 sg13g2_dfrbp_1 _2133_ (.CLK(net843),
    .RESET_B(net997),
    .D(\u_top_module.u_buffer.shift_reg_1[175] ),
    .Q_N(_0955_),
    .Q(\u_top_module.u_buffer.shift_reg_1[176] ));
 sg13g2_dfrbp_1 _2134_ (.CLK(net843),
    .RESET_B(net998),
    .D(\u_top_module.u_buffer.shift_reg_1[176] ),
    .Q_N(_0956_),
    .Q(\u_top_module.u_buffer.shift_reg_1[177] ));
 sg13g2_dfrbp_1 _2135_ (.CLK(net850),
    .RESET_B(net998),
    .D(\u_top_module.u_buffer.shift_reg_1[177] ),
    .Q_N(_0957_),
    .Q(\u_top_module.u_buffer.shift_reg_1[178] ));
 sg13g2_dfrbp_1 _2136_ (.CLK(net849),
    .RESET_B(net997),
    .D(\u_top_module.u_buffer.shift_reg_1[178] ),
    .Q_N(_0958_),
    .Q(\u_top_module.u_buffer.shift_reg_1[179] ));
 sg13g2_dfrbp_1 _2137_ (.CLK(net849),
    .RESET_B(net1003),
    .D(\u_top_module.u_buffer.shift_reg_1[179] ),
    .Q_N(_0959_),
    .Q(\u_top_module.u_buffer.shift_reg_1[180] ));
 sg13g2_dfrbp_1 _2138_ (.CLK(net849),
    .RESET_B(net1003),
    .D(\u_top_module.u_buffer.shift_reg_1[180] ),
    .Q_N(_0960_),
    .Q(\u_top_module.u_buffer.shift_reg_1[181] ));
 sg13g2_dfrbp_1 _2139_ (.CLK(net849),
    .RESET_B(net1003),
    .D(\u_top_module.u_buffer.shift_reg_1[181] ),
    .Q_N(_0961_),
    .Q(\u_top_module.u_buffer.shift_reg_1[182] ));
 sg13g2_dfrbp_1 _2140_ (.CLK(net849),
    .RESET_B(net1003),
    .D(\u_top_module.u_buffer.shift_reg_1[182] ),
    .Q_N(_0962_),
    .Q(\u_top_module.u_buffer.shift_reg_1[183] ));
 sg13g2_dfrbp_1 _2141_ (.CLK(net848),
    .RESET_B(net1000),
    .D(\u_top_module.u_buffer.shift_reg_1[183] ),
    .Q_N(_0963_),
    .Q(\u_top_module.u_buffer.shift_reg_1[184] ));
 sg13g2_dfrbp_1 _2142_ (.CLK(net848),
    .RESET_B(net1000),
    .D(\u_top_module.u_buffer.shift_reg_1[184] ),
    .Q_N(_0964_),
    .Q(\u_top_module.u_buffer.shift_reg_1[185] ));
 sg13g2_dfrbp_1 _2143_ (.CLK(net848),
    .RESET_B(net1000),
    .D(\u_top_module.u_buffer.shift_reg_1[185] ),
    .Q_N(_0965_),
    .Q(\u_top_module.u_buffer.shift_reg_1[186] ));
 sg13g2_dfrbp_1 _2144_ (.CLK(net848),
    .RESET_B(net1000),
    .D(\u_top_module.u_buffer.shift_reg_1[186] ),
    .Q_N(_0966_),
    .Q(\u_top_module.u_buffer.shift_reg_1[187] ));
 sg13g2_dfrbp_1 _2145_ (.CLK(net848),
    .RESET_B(net1000),
    .D(\u_top_module.u_buffer.shift_reg_1[187] ),
    .Q_N(_0967_),
    .Q(\u_top_module.u_buffer.shift_reg_1[188] ));
 sg13g2_dfrbp_1 _2146_ (.CLK(net847),
    .RESET_B(net1000),
    .D(\u_top_module.u_buffer.shift_reg_1[188] ),
    .Q_N(_0968_),
    .Q(\u_top_module.u_buffer.shift_reg_1[189] ));
 sg13g2_dfrbp_1 _2147_ (.CLK(net846),
    .RESET_B(net1002),
    .D(\u_top_module.u_buffer.shift_reg_1[189] ),
    .Q_N(_0969_),
    .Q(\u_top_module.u_buffer.shift_reg_1[190] ));
 sg13g2_dfrbp_1 _2148_ (.CLK(net846),
    .RESET_B(net1002),
    .D(\u_top_module.u_buffer.shift_reg_1[190] ),
    .Q_N(_0970_),
    .Q(\u_top_module.u_buffer.shift_reg_1[191] ));
 sg13g2_dfrbp_1 _2149_ (.CLK(net846),
    .RESET_B(net1002),
    .D(\u_top_module.u_buffer.shift_reg_1[191] ),
    .Q_N(_0971_),
    .Q(\u_top_module.u_buffer.shift_reg_1[192] ));
 sg13g2_dfrbp_1 _2150_ (.CLK(net846),
    .RESET_B(net1002),
    .D(\u_top_module.u_buffer.shift_reg_1[192] ),
    .Q_N(_0972_),
    .Q(\u_top_module.u_buffer.shift_reg_1[193] ));
 sg13g2_dfrbp_1 _2151_ (.CLK(net846),
    .RESET_B(net1002),
    .D(\u_top_module.u_buffer.shift_reg_1[193] ),
    .Q_N(_0973_),
    .Q(\u_top_module.u_buffer.shift_reg_1[194] ));
 sg13g2_dfrbp_1 _2152_ (.CLK(net861),
    .RESET_B(net991),
    .D(\u_top_module.u_buffer.shift_reg_1[194] ),
    .Q_N(_0974_),
    .Q(\u_top_module.u_buffer.shift_reg_1[195] ));
 sg13g2_dfrbp_1 _2153_ (.CLK(net861),
    .RESET_B(net1017),
    .D(\u_top_module.u_buffer.shift_reg_1[195] ),
    .Q_N(_0975_),
    .Q(\u_top_module.u_buffer.shift_reg_1[196] ));
 sg13g2_dfrbp_1 _2154_ (.CLK(net861),
    .RESET_B(net1017),
    .D(\u_top_module.u_buffer.shift_reg_1[196] ),
    .Q_N(_0976_),
    .Q(\u_top_module.u_buffer.shift_reg_1[197] ));
 sg13g2_dfrbp_1 _2155_ (.CLK(net861),
    .RESET_B(net1014),
    .D(\u_top_module.u_buffer.shift_reg_1[197] ),
    .Q_N(_0977_),
    .Q(\u_top_module.u_buffer.shift_reg_1[198] ));
 sg13g2_dfrbp_1 _2156_ (.CLK(net860),
    .RESET_B(net1014),
    .D(\u_top_module.u_buffer.shift_reg_1[198] ),
    .Q_N(_0978_),
    .Q(\u_top_module.u_buffer.shift_reg_1[199] ));
 sg13g2_dfrbp_1 _2157_ (.CLK(net860),
    .RESET_B(net1014),
    .D(\u_top_module.u_buffer.shift_reg_1[199] ),
    .Q_N(_0979_),
    .Q(\u_top_module.u_buffer.shift_reg_1[200] ));
 sg13g2_dfrbp_1 _2158_ (.CLK(net862),
    .RESET_B(net1014),
    .D(\u_top_module.u_buffer.shift_reg_1[200] ),
    .Q_N(_0980_),
    .Q(\u_top_module.u_buffer.shift_reg_1[201] ));
 sg13g2_dfrbp_1 _2159_ (.CLK(net862),
    .RESET_B(net1015),
    .D(\u_top_module.u_buffer.shift_reg_1[201] ),
    .Q_N(_0981_),
    .Q(\u_top_module.u_buffer.shift_reg_1[202] ));
 sg13g2_dfrbp_1 _2160_ (.CLK(net862),
    .RESET_B(net1015),
    .D(\u_top_module.u_buffer.shift_reg_1[202] ),
    .Q_N(_0982_),
    .Q(\u_top_module.u_buffer.shift_reg_1[203] ));
 sg13g2_dfrbp_1 _2161_ (.CLK(net862),
    .RESET_B(net1016),
    .D(\u_top_module.u_buffer.shift_reg_1[203] ),
    .Q_N(_0983_),
    .Q(\u_top_module.u_buffer.shift_reg_1[204] ));
 sg13g2_dfrbp_1 _2162_ (.CLK(net862),
    .RESET_B(net1015),
    .D(\u_top_module.u_buffer.shift_reg_1[204] ),
    .Q_N(_0984_),
    .Q(\u_top_module.u_buffer.shift_reg_1[205] ));
 sg13g2_dfrbp_1 _2163_ (.CLK(net870),
    .RESET_B(net1015),
    .D(\u_top_module.u_buffer.shift_reg_1[205] ),
    .Q_N(_0985_),
    .Q(\u_top_module.u_buffer.shift_reg_1[206] ));
 sg13g2_dfrbp_1 _2164_ (.CLK(net870),
    .RESET_B(net1015),
    .D(\u_top_module.u_buffer.shift_reg_1[206] ),
    .Q_N(_0986_),
    .Q(\u_top_module.u_buffer.shift_reg_1[207] ));
 sg13g2_dfrbp_1 _2165_ (.CLK(net870),
    .RESET_B(net1023),
    .D(\u_top_module.u_buffer.shift_reg_1[207] ),
    .Q_N(_0987_),
    .Q(\u_top_module.u_buffer.shift_reg_1[208] ));
 sg13g2_dfrbp_1 _2166_ (.CLK(net870),
    .RESET_B(net1023),
    .D(\u_top_module.u_buffer.shift_reg_1[208] ),
    .Q_N(_0988_),
    .Q(\u_top_module.u_buffer.shift_reg_1[209] ));
 sg13g2_dfrbp_1 _2167_ (.CLK(net870),
    .RESET_B(net1023),
    .D(\u_top_module.u_buffer.shift_reg_1[209] ),
    .Q_N(_0989_),
    .Q(\u_top_module.u_buffer.shift_reg_1[210] ));
 sg13g2_dfrbp_1 _2168_ (.CLK(net870),
    .RESET_B(net1023),
    .D(\u_top_module.u_buffer.shift_reg_1[210] ),
    .Q_N(_0990_),
    .Q(\u_top_module.u_buffer.shift_reg_1[211] ));
 sg13g2_dfrbp_1 _2169_ (.CLK(net870),
    .RESET_B(net1023),
    .D(\u_top_module.u_buffer.shift_reg_1[211] ),
    .Q_N(_0991_),
    .Q(\u_top_module.u_buffer.shift_reg_1[212] ));
 sg13g2_dfrbp_1 _2170_ (.CLK(net868),
    .RESET_B(net1020),
    .D(\u_top_module.u_buffer.shift_reg_1[212] ),
    .Q_N(_0992_),
    .Q(\u_top_module.u_buffer.shift_reg_1[213] ));
 sg13g2_dfrbp_1 _2171_ (.CLK(net868),
    .RESET_B(net1020),
    .D(\u_top_module.u_buffer.shift_reg_1[213] ),
    .Q_N(_0993_),
    .Q(\u_top_module.u_buffer.shift_reg_1[214] ));
 sg13g2_dfrbp_1 _2172_ (.CLK(net868),
    .RESET_B(net1020),
    .D(\u_top_module.u_buffer.shift_reg_1[214] ),
    .Q_N(_0994_),
    .Q(\u_top_module.u_buffer.shift_reg_1[215] ));
 sg13g2_dfrbp_1 _2173_ (.CLK(net868),
    .RESET_B(net1021),
    .D(\u_top_module.u_buffer.shift_reg_1[215] ),
    .Q_N(_0995_),
    .Q(\u_top_module.u_buffer.shift_reg_1[216] ));
 sg13g2_dfrbp_1 _2174_ (.CLK(net868),
    .RESET_B(net1021),
    .D(\u_top_module.u_buffer.shift_reg_1[216] ),
    .Q_N(_0996_),
    .Q(\u_top_module.u_buffer.shift_reg_1[217] ));
 sg13g2_dfrbp_1 _2175_ (.CLK(net869),
    .RESET_B(net1021),
    .D(\u_top_module.u_buffer.shift_reg_1[217] ),
    .Q_N(_0997_),
    .Q(\u_top_module.u_buffer.shift_reg_1[218] ));
 sg13g2_dfrbp_1 _2176_ (.CLK(net869),
    .RESET_B(net1021),
    .D(\u_top_module.u_buffer.shift_reg_1[218] ),
    .Q_N(_0998_),
    .Q(\u_top_module.u_buffer.shift_reg_1[219] ));
 sg13g2_dfrbp_1 _2177_ (.CLK(net869),
    .RESET_B(net1021),
    .D(\u_top_module.u_buffer.shift_reg_1[219] ),
    .Q_N(_0999_),
    .Q(\u_top_module.u_buffer.shift_reg_1[220] ));
 sg13g2_dfrbp_1 _2178_ (.CLK(net868),
    .RESET_B(net1021),
    .D(\u_top_module.u_buffer.shift_reg_1[220] ),
    .Q_N(_1000_),
    .Q(\u_top_module.u_buffer.shift_reg_1[221] ));
 sg13g2_dfrbp_1 _2179_ (.CLK(net868),
    .RESET_B(net1021),
    .D(\u_top_module.u_buffer.shift_reg_1[221] ),
    .Q_N(_1001_),
    .Q(\u_top_module.u_buffer.shift_reg_1[222] ));
 sg13g2_dfrbp_1 _2180_ (.CLK(net869),
    .RESET_B(net1026),
    .D(\u_top_module.u_buffer.shift_reg_1[222] ),
    .Q_N(_1002_),
    .Q(\u_top_module.u_buffer.shift_reg_1[223] ));
 sg13g2_dfrbp_1 _2181_ (.CLK(net868),
    .RESET_B(net1021),
    .D(\u_top_module.u_buffer.shift_reg_1[223] ),
    .Q_N(_1003_),
    .Q(\u_top_module.u_buffer.shift_reg_1[224] ));
 sg13g2_dfrbp_1 _2182_ (.CLK(net873),
    .RESET_B(net1024),
    .D(\u_top_module.u_buffer.shift_reg_1[224] ),
    .Q_N(_1004_),
    .Q(\u_top_module.u_buffer.shift_reg_1[225] ));
 sg13g2_dfrbp_1 _2183_ (.CLK(net873),
    .RESET_B(net1024),
    .D(\u_top_module.u_buffer.shift_reg_1[225] ),
    .Q_N(_1005_),
    .Q(\u_top_module.u_buffer.shift_reg_1[226] ));
 sg13g2_dfrbp_1 _2184_ (.CLK(net873),
    .RESET_B(net1024),
    .D(\u_top_module.u_buffer.shift_reg_1[226] ),
    .Q_N(_1006_),
    .Q(\u_top_module.u_buffer.shift_reg_1[227] ));
 sg13g2_dfrbp_1 _2185_ (.CLK(net873),
    .RESET_B(net1024),
    .D(\u_top_module.u_buffer.shift_reg_1[227] ),
    .Q_N(_1007_),
    .Q(\u_top_module.u_buffer.shift_reg_1[228] ));
 sg13g2_dfrbp_1 _2186_ (.CLK(net873),
    .RESET_B(net1024),
    .D(\u_top_module.u_buffer.shift_reg_1[228] ),
    .Q_N(_1008_),
    .Q(\u_top_module.u_buffer.shift_reg_1[229] ));
 sg13g2_dfrbp_1 _2187_ (.CLK(net872),
    .RESET_B(net1024),
    .D(\u_top_module.u_buffer.shift_reg_1[229] ),
    .Q_N(_1009_),
    .Q(\u_top_module.u_buffer.shift_reg_1[230] ));
 sg13g2_dfrbp_1 _2188_ (.CLK(net872),
    .RESET_B(net1024),
    .D(\u_top_module.u_buffer.shift_reg_1[230] ),
    .Q_N(_1010_),
    .Q(\u_top_module.u_buffer.shift_reg_1[231] ));
 sg13g2_dfrbp_1 _2189_ (.CLK(net873),
    .RESET_B(net1025),
    .D(\u_top_module.u_buffer.shift_reg_1[231] ),
    .Q_N(_1011_),
    .Q(\u_top_module.u_buffer.shift_reg_1[232] ));
 sg13g2_dfrbp_1 _2190_ (.CLK(net872),
    .RESET_B(net1024),
    .D(\u_top_module.u_buffer.shift_reg_1[232] ),
    .Q_N(_1012_),
    .Q(\u_top_module.u_buffer.shift_reg_1[233] ));
 sg13g2_dfrbp_1 _2191_ (.CLK(net881),
    .RESET_B(net1034),
    .D(\u_top_module.u_buffer.shift_reg_1[233] ),
    .Q_N(_1013_),
    .Q(\u_top_module.u_buffer.shift_reg_1[234] ));
 sg13g2_dfrbp_1 _2192_ (.CLK(net881),
    .RESET_B(net1034),
    .D(\u_top_module.u_buffer.shift_reg_1[234] ),
    .Q_N(_1014_),
    .Q(\u_top_module.u_buffer.shift_reg_1[235] ));
 sg13g2_dfrbp_1 _2193_ (.CLK(net880),
    .RESET_B(net1034),
    .D(\u_top_module.u_buffer.shift_reg_1[235] ),
    .Q_N(_1015_),
    .Q(\u_top_module.u_buffer.shift_reg_1[236] ));
 sg13g2_dfrbp_1 _2194_ (.CLK(net880),
    .RESET_B(net1034),
    .D(\u_top_module.u_buffer.shift_reg_1[236] ),
    .Q_N(_1016_),
    .Q(\u_top_module.u_buffer.shift_reg_1[237] ));
 sg13g2_dfrbp_1 _2195_ (.CLK(net880),
    .RESET_B(net1034),
    .D(\u_top_module.u_buffer.shift_reg_1[237] ),
    .Q_N(_1017_),
    .Q(\u_top_module.u_buffer.shift_reg_1[238] ));
 sg13g2_dfrbp_1 _2196_ (.CLK(net881),
    .RESET_B(net1035),
    .D(\u_top_module.u_buffer.shift_reg_1[238] ),
    .Q_N(_1018_),
    .Q(\u_top_module.u_buffer.shift_reg_1[239] ));
 sg13g2_dfrbp_1 _2197_ (.CLK(net881),
    .RESET_B(net1035),
    .D(\u_top_module.u_buffer.shift_reg_1[239] ),
    .Q_N(_1019_),
    .Q(\u_top_module.u_buffer.shift_reg_1[240] ));
 sg13g2_dfrbp_1 _2198_ (.CLK(net881),
    .RESET_B(net1035),
    .D(\u_top_module.u_buffer.shift_reg_1[240] ),
    .Q_N(_1020_),
    .Q(\u_top_module.u_buffer.shift_reg_1[241] ));
 sg13g2_dfrbp_1 _2199_ (.CLK(net881),
    .RESET_B(net1035),
    .D(\u_top_module.u_buffer.shift_reg_1[241] ),
    .Q_N(_1021_),
    .Q(\u_top_module.u_buffer.shift_reg_1[242] ));
 sg13g2_dfrbp_1 _2200_ (.CLK(net881),
    .RESET_B(net1035),
    .D(\u_top_module.u_buffer.shift_reg_1[242] ),
    .Q_N(_1022_),
    .Q(\u_top_module.u_buffer.shift_reg_1[243] ));
 sg13g2_dfrbp_1 _2201_ (.CLK(net883),
    .RESET_B(net1038),
    .D(\u_top_module.u_buffer.shift_reg_1[243] ),
    .Q_N(_1023_),
    .Q(\u_top_module.u_buffer.shift_reg_1[244] ));
 sg13g2_dfrbp_1 _2202_ (.CLK(net883),
    .RESET_B(net1038),
    .D(\u_top_module.u_buffer.shift_reg_1[244] ),
    .Q_N(_1024_),
    .Q(\u_top_module.u_buffer.shift_reg_1[245] ));
 sg13g2_dfrbp_1 _2203_ (.CLK(net883),
    .RESET_B(net1037),
    .D(\u_top_module.u_buffer.shift_reg_1[245] ),
    .Q_N(_1025_),
    .Q(\u_top_module.u_buffer.shift_reg_1[246] ));
 sg13g2_dfrbp_1 _2204_ (.CLK(net883),
    .RESET_B(net1038),
    .D(\u_top_module.u_buffer.shift_reg_1[246] ),
    .Q_N(_1026_),
    .Q(\u_top_module.u_buffer.shift_reg_1[247] ));
 sg13g2_dfrbp_1 _2205_ (.CLK(net851),
    .RESET_B(net1005),
    .D(\u_top_module.u_buffer.shift_reg_1[247] ),
    .Q_N(_1027_),
    .Q(\u_top_module.u_buffer.shift_reg_1[248] ));
 sg13g2_dfrbp_1 _2206_ (.CLK(net913),
    .RESET_B(net1050),
    .D(\u_top_module.u_buffer.shift_reg_1[248] ),
    .Q_N(_1028_),
    .Q(\u_top_module.u_buffer.shift_reg_1[249] ));
 sg13g2_dfrbp_1 _2207_ (.CLK(net913),
    .RESET_B(net1069),
    .D(\u_top_module.u_buffer.shift_reg_1[249] ),
    .Q_N(_1029_),
    .Q(\u_top_module.u_buffer.shift_reg_1[250] ));
 sg13g2_dfrbp_1 _2208_ (.CLK(net913),
    .RESET_B(net1069),
    .D(\u_top_module.u_buffer.shift_reg_1[250] ),
    .Q_N(_1030_),
    .Q(\u_top_module.u_buffer.shift_reg_1[251] ));
 sg13g2_dfrbp_1 _2209_ (.CLK(net913),
    .RESET_B(net1073),
    .D(\u_top_module.u_buffer.shift_reg_1[251] ),
    .Q_N(_1031_),
    .Q(\u_top_module.u_buffer.shift_reg_1[252] ));
 sg13g2_dfrbp_1 _2210_ (.CLK(net914),
    .RESET_B(net1073),
    .D(\u_top_module.u_buffer.shift_reg_1[252] ),
    .Q_N(_1032_),
    .Q(\u_top_module.u_buffer.shift_reg_1[253] ));
 sg13g2_dfrbp_1 _2211_ (.CLK(net915),
    .RESET_B(net1078),
    .D(\u_top_module.u_buffer.shift_reg_1[253] ),
    .Q_N(_1033_),
    .Q(\u_top_module.u_buffer.shift_reg_1[254] ));
 sg13g2_dfrbp_1 _2212_ (.CLK(net915),
    .RESET_B(net1078),
    .D(\u_top_module.u_buffer.shift_reg_1[254] ),
    .Q_N(_1034_),
    .Q(\u_top_module.u_buffer.shift_reg_1[255] ));
 sg13g2_dfrbp_1 _2213_ (.CLK(net910),
    .RESET_B(net1066),
    .D(_0000_),
    .Q_N(_1035_),
    .Q(\u_top_module.neg ));
 sg13g2_dfrbp_1 _2214_ (.CLK(net916),
    .RESET_B(net1081),
    .D(_0018_),
    .Q_N(_0014_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _2215_ (.CLK(net916),
    .RESET_B(net1081),
    .D(_0019_),
    .Q_N(_1036_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _2216_ (.CLK(net916),
    .RESET_B(net1081),
    .D(_0020_),
    .Q_N(_1037_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _2217_ (.CLK(net916),
    .RESET_B(net1081),
    .D(_0021_),
    .Q_N(_1038_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _2218_ (.CLK(net916),
    .RESET_B(net1067),
    .D(_0022_),
    .Q_N(_1039_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2219_ (.CLK(net915),
    .RESET_B(net1067),
    .D(_0023_),
    .Q_N(_1040_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2220_ (.CLK(net910),
    .RESET_B(net1066),
    .D(_0024_),
    .Q_N(_1041_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _2221_ (.CLK(net911),
    .RESET_B(net1066),
    .D(_0025_),
    .Q_N(_1042_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _2222_ (.CLK(net915),
    .RESET_B(net1063),
    .D(\u_top_module.dec_data_2 ),
    .Q_N(_1043_),
    .Q(\u_top_module.u_buffer.shift_reg_2[0] ));
 sg13g2_dfrbp_1 _2223_ (.CLK(net907),
    .RESET_B(net1063),
    .D(\u_top_module.u_buffer.shift_reg_2[0] ),
    .Q_N(_1044_),
    .Q(\u_top_module.u_buffer.shift_reg_2[1] ));
 sg13g2_dfrbp_1 _2224_ (.CLK(net907),
    .RESET_B(net1063),
    .D(\u_top_module.u_buffer.shift_reg_2[1] ),
    .Q_N(_1045_),
    .Q(\u_top_module.u_buffer.shift_reg_2[2] ));
 sg13g2_dfrbp_1 _2225_ (.CLK(net898),
    .RESET_B(net1053),
    .D(\u_top_module.u_buffer.shift_reg_2[2] ),
    .Q_N(_1046_),
    .Q(\u_top_module.u_buffer.shift_reg_2[3] ));
 sg13g2_dfrbp_1 _2226_ (.CLK(net899),
    .RESET_B(net1052),
    .D(\u_top_module.u_buffer.shift_reg_2[3] ),
    .Q_N(_1047_),
    .Q(\u_top_module.u_buffer.shift_reg_2[4] ));
 sg13g2_dfrbp_1 _2227_ (.CLK(net898),
    .RESET_B(net1052),
    .D(\u_top_module.u_buffer.shift_reg_2[4] ),
    .Q_N(_1048_),
    .Q(\u_top_module.u_buffer.shift_reg_2[5] ));
 sg13g2_dfrbp_1 _2228_ (.CLK(net898),
    .RESET_B(net1052),
    .D(\u_top_module.u_buffer.shift_reg_2[5] ),
    .Q_N(_1049_),
    .Q(\u_top_module.u_buffer.shift_reg_2[6] ));
 sg13g2_dfrbp_1 _2229_ (.CLK(net899),
    .RESET_B(net1053),
    .D(\u_top_module.u_buffer.shift_reg_2[6] ),
    .Q_N(_1050_),
    .Q(\u_top_module.u_buffer.shift_reg_2[7] ));
 sg13g2_dfrbp_1 _2230_ (.CLK(net899),
    .RESET_B(net1053),
    .D(\u_top_module.u_buffer.shift_reg_2[7] ),
    .Q_N(_1051_),
    .Q(\u_top_module.u_buffer.shift_reg_2[8] ));
 sg13g2_dfrbp_1 _2231_ (.CLK(net899),
    .RESET_B(net1053),
    .D(\u_top_module.u_buffer.shift_reg_2[8] ),
    .Q_N(_1052_),
    .Q(\u_top_module.u_buffer.shift_reg_2[9] ));
 sg13g2_dfrbp_1 _2232_ (.CLK(net895),
    .RESET_B(net1049),
    .D(\u_top_module.u_buffer.shift_reg_2[9] ),
    .Q_N(_1053_),
    .Q(\u_top_module.u_buffer.shift_reg_2[10] ));
 sg13g2_dfrbp_1 _2233_ (.CLK(net895),
    .RESET_B(net1051),
    .D(\u_top_module.u_buffer.shift_reg_2[10] ),
    .Q_N(_1054_),
    .Q(\u_top_module.u_buffer.shift_reg_2[11] ));
 sg13g2_dfrbp_1 _2234_ (.CLK(net895),
    .RESET_B(net1051),
    .D(\u_top_module.u_buffer.shift_reg_2[11] ),
    .Q_N(_1055_),
    .Q(\u_top_module.u_buffer.shift_reg_2[12] ));
 sg13g2_dfrbp_1 _2235_ (.CLK(net895),
    .RESET_B(net1049),
    .D(\u_top_module.u_buffer.shift_reg_2[12] ),
    .Q_N(_1056_),
    .Q(\u_top_module.u_buffer.shift_reg_2[13] ));
 sg13g2_dfrbp_1 _2236_ (.CLK(net895),
    .RESET_B(net1051),
    .D(\u_top_module.u_buffer.shift_reg_2[13] ),
    .Q_N(_1057_),
    .Q(\u_top_module.u_buffer.shift_reg_2[14] ));
 sg13g2_dfrbp_1 _2237_ (.CLK(net897),
    .RESET_B(net1051),
    .D(\u_top_module.u_buffer.shift_reg_2[14] ),
    .Q_N(_1058_),
    .Q(\u_top_module.u_buffer.shift_reg_2[15] ));
 sg13g2_dfrbp_1 _2238_ (.CLK(net897),
    .RESET_B(net1051),
    .D(\u_top_module.u_buffer.shift_reg_2[15] ),
    .Q_N(_1059_),
    .Q(\u_top_module.u_buffer.shift_reg_2[16] ));
 sg13g2_dfrbp_1 _2239_ (.CLK(net896),
    .RESET_B(net1050),
    .D(\u_top_module.u_buffer.shift_reg_2[16] ),
    .Q_N(_1060_),
    .Q(\u_top_module.u_buffer.shift_reg_2[17] ));
 sg13g2_dfrbp_1 _2240_ (.CLK(net896),
    .RESET_B(net1050),
    .D(\u_top_module.u_buffer.shift_reg_2[17] ),
    .Q_N(_1061_),
    .Q(\u_top_module.u_buffer.shift_reg_2[18] ));
 sg13g2_dfrbp_1 _2241_ (.CLK(net896),
    .RESET_B(net1050),
    .D(\u_top_module.u_buffer.shift_reg_2[18] ),
    .Q_N(_1062_),
    .Q(\u_top_module.u_buffer.shift_reg_2[19] ));
 sg13g2_dfrbp_1 _2242_ (.CLK(net896),
    .RESET_B(net1050),
    .D(\u_top_module.u_buffer.shift_reg_2[19] ),
    .Q_N(_1063_),
    .Q(\u_top_module.u_buffer.shift_reg_2[20] ));
 sg13g2_dfrbp_1 _2243_ (.CLK(net852),
    .RESET_B(net1006),
    .D(\u_top_module.u_buffer.shift_reg_2[20] ),
    .Q_N(_1064_),
    .Q(\u_top_module.u_buffer.shift_reg_2[21] ));
 sg13g2_dfrbp_1 _2244_ (.CLK(net851),
    .RESET_B(net1006),
    .D(\u_top_module.u_buffer.shift_reg_2[21] ),
    .Q_N(_1065_),
    .Q(\u_top_module.u_buffer.shift_reg_2[22] ));
 sg13g2_dfrbp_1 _2245_ (.CLK(net850),
    .RESET_B(net1004),
    .D(\u_top_module.u_buffer.shift_reg_2[22] ),
    .Q_N(_1066_),
    .Q(\u_top_module.u_buffer.shift_reg_2[23] ));
 sg13g2_dfrbp_1 _2246_ (.CLK(net850),
    .RESET_B(net1003),
    .D(\u_top_module.u_buffer.shift_reg_2[23] ),
    .Q_N(_1067_),
    .Q(\u_top_module.u_buffer.shift_reg_2[24] ));
 sg13g2_dfrbp_1 _2247_ (.CLK(net849),
    .RESET_B(net1003),
    .D(\u_top_module.u_buffer.shift_reg_2[24] ),
    .Q_N(_1068_),
    .Q(\u_top_module.u_buffer.shift_reg_2[25] ));
 sg13g2_dfrbp_1 _2248_ (.CLK(net849),
    .RESET_B(net1003),
    .D(\u_top_module.u_buffer.shift_reg_2[25] ),
    .Q_N(_1069_),
    .Q(\u_top_module.u_buffer.shift_reg_2[26] ));
 sg13g2_dfrbp_1 _2249_ (.CLK(net849),
    .RESET_B(net1003),
    .D(\u_top_module.u_buffer.shift_reg_2[26] ),
    .Q_N(_1070_),
    .Q(\u_top_module.u_buffer.shift_reg_2[27] ));
 sg13g2_dfrbp_1 _2250_ (.CLK(net847),
    .RESET_B(net1001),
    .D(\u_top_module.u_buffer.shift_reg_2[27] ),
    .Q_N(_1071_),
    .Q(\u_top_module.u_buffer.shift_reg_2[28] ));
 sg13g2_dfrbp_1 _2251_ (.CLK(net847),
    .RESET_B(net1000),
    .D(\u_top_module.u_buffer.shift_reg_2[28] ),
    .Q_N(_1072_),
    .Q(\u_top_module.u_buffer.shift_reg_2[29] ));
 sg13g2_dfrbp_1 _2252_ (.CLK(net847),
    .RESET_B(net1000),
    .D(\u_top_module.u_buffer.shift_reg_2[29] ),
    .Q_N(_1073_),
    .Q(\u_top_module.u_buffer.shift_reg_2[30] ));
 sg13g2_dfrbp_1 _2253_ (.CLK(net846),
    .RESET_B(net1001),
    .D(\u_top_module.u_buffer.shift_reg_2[30] ),
    .Q_N(_1074_),
    .Q(\u_top_module.u_buffer.shift_reg_2[31] ));
 sg13g2_dfrbp_1 _2254_ (.CLK(net846),
    .RESET_B(net1001),
    .D(\u_top_module.u_buffer.shift_reg_2[31] ),
    .Q_N(_1075_),
    .Q(\u_top_module.u_buffer.shift_reg_2[32] ));
 sg13g2_dfrbp_1 _2255_ (.CLK(net846),
    .RESET_B(net1001),
    .D(\u_top_module.u_buffer.shift_reg_2[32] ),
    .Q_N(_1076_),
    .Q(\u_top_module.u_buffer.shift_reg_2[33] ));
 sg13g2_dfrbp_1 _2256_ (.CLK(net837),
    .RESET_B(net990),
    .D(\u_top_module.u_buffer.shift_reg_2[33] ),
    .Q_N(_1077_),
    .Q(\u_top_module.u_buffer.shift_reg_2[34] ));
 sg13g2_dfrbp_1 _2257_ (.CLK(net837),
    .RESET_B(net990),
    .D(\u_top_module.u_buffer.shift_reg_2[34] ),
    .Q_N(_1078_),
    .Q(\u_top_module.u_buffer.shift_reg_2[35] ));
 sg13g2_dfrbp_1 _2258_ (.CLK(net838),
    .RESET_B(net991),
    .D(\u_top_module.u_buffer.shift_reg_2[35] ),
    .Q_N(_1079_),
    .Q(\u_top_module.u_buffer.shift_reg_2[36] ));
 sg13g2_dfrbp_1 _2259_ (.CLK(net838),
    .RESET_B(net991),
    .D(\u_top_module.u_buffer.shift_reg_2[36] ),
    .Q_N(_1080_),
    .Q(\u_top_module.u_buffer.shift_reg_2[37] ));
 sg13g2_dfrbp_1 _2260_ (.CLK(net837),
    .RESET_B(net991),
    .D(\u_top_module.u_buffer.shift_reg_2[37] ),
    .Q_N(_1081_),
    .Q(\u_top_module.u_buffer.shift_reg_2[38] ));
 sg13g2_dfrbp_1 _2261_ (.CLK(net838),
    .RESET_B(net990),
    .D(\u_top_module.u_buffer.shift_reg_2[38] ),
    .Q_N(_1082_),
    .Q(\u_top_module.u_buffer.shift_reg_2[39] ));
 sg13g2_dfrbp_1 _2262_ (.CLK(net837),
    .RESET_B(net990),
    .D(\u_top_module.u_buffer.shift_reg_2[39] ),
    .Q_N(_1083_),
    .Q(\u_top_module.u_buffer.shift_reg_2[40] ));
 sg13g2_dfrbp_1 _2263_ (.CLK(net837),
    .RESET_B(net990),
    .D(\u_top_module.u_buffer.shift_reg_2[40] ),
    .Q_N(_1084_),
    .Q(\u_top_module.u_buffer.shift_reg_2[41] ));
 sg13g2_dfrbp_1 _2264_ (.CLK(net860),
    .RESET_B(net990),
    .D(\u_top_module.u_buffer.shift_reg_2[41] ),
    .Q_N(_1085_),
    .Q(\u_top_module.u_buffer.shift_reg_2[42] ));
 sg13g2_dfrbp_1 _2265_ (.CLK(net860),
    .RESET_B(net990),
    .D(\u_top_module.u_buffer.shift_reg_2[42] ),
    .Q_N(_1086_),
    .Q(\u_top_module.u_buffer.shift_reg_2[43] ));
 sg13g2_dfrbp_1 _2266_ (.CLK(net860),
    .RESET_B(net1014),
    .D(\u_top_module.u_buffer.shift_reg_2[43] ),
    .Q_N(_1087_),
    .Q(\u_top_module.u_buffer.shift_reg_2[44] ));
 sg13g2_dfrbp_1 _2267_ (.CLK(net860),
    .RESET_B(net990),
    .D(\u_top_module.u_buffer.shift_reg_2[44] ),
    .Q_N(_1088_),
    .Q(\u_top_module.u_buffer.shift_reg_2[45] ));
 sg13g2_dfrbp_1 _2268_ (.CLK(net857),
    .RESET_B(net986),
    .D(\u_top_module.u_buffer.shift_reg_2[45] ),
    .Q_N(_1089_),
    .Q(\u_top_module.u_buffer.shift_reg_2[46] ));
 sg13g2_dfrbp_1 _2269_ (.CLK(net833),
    .RESET_B(net986),
    .D(\u_top_module.u_buffer.shift_reg_2[46] ),
    .Q_N(_1090_),
    .Q(\u_top_module.u_buffer.shift_reg_2[47] ));
 sg13g2_dfrbp_1 _2270_ (.CLK(net833),
    .RESET_B(net987),
    .D(\u_top_module.u_buffer.shift_reg_2[47] ),
    .Q_N(_1091_),
    .Q(\u_top_module.u_buffer.shift_reg_2[48] ));
 sg13g2_dfrbp_1 _2271_ (.CLK(net833),
    .RESET_B(net987),
    .D(\u_top_module.u_buffer.shift_reg_2[48] ),
    .Q_N(_1092_),
    .Q(\u_top_module.u_buffer.shift_reg_2[49] ));
 sg13g2_dfrbp_1 _2272_ (.CLK(net833),
    .RESET_B(net986),
    .D(\u_top_module.u_buffer.shift_reg_2[49] ),
    .Q_N(_1093_),
    .Q(\u_top_module.u_buffer.shift_reg_2[50] ));
 sg13g2_dfrbp_1 _2273_ (.CLK(net833),
    .RESET_B(net986),
    .D(\u_top_module.u_buffer.shift_reg_2[50] ),
    .Q_N(_1094_),
    .Q(\u_top_module.u_buffer.shift_reg_2[51] ));
 sg13g2_dfrbp_1 _2274_ (.CLK(net833),
    .RESET_B(net986),
    .D(\u_top_module.u_buffer.shift_reg_2[51] ),
    .Q_N(_1095_),
    .Q(\u_top_module.u_buffer.shift_reg_2[52] ));
 sg13g2_dfrbp_1 _2275_ (.CLK(net833),
    .RESET_B(net986),
    .D(\u_top_module.u_buffer.shift_reg_2[52] ),
    .Q_N(_1096_),
    .Q(\u_top_module.u_buffer.shift_reg_2[53] ));
 sg13g2_dfrbp_1 _2276_ (.CLK(net833),
    .RESET_B(net984),
    .D(\u_top_module.u_buffer.shift_reg_2[53] ),
    .Q_N(_1097_),
    .Q(\u_top_module.u_buffer.shift_reg_2[54] ));
 sg13g2_dfrbp_1 _2277_ (.CLK(net831),
    .RESET_B(net984),
    .D(\u_top_module.u_buffer.shift_reg_2[54] ),
    .Q_N(_1098_),
    .Q(\u_top_module.u_buffer.shift_reg_2[55] ));
 sg13g2_dfrbp_1 _2278_ (.CLK(net831),
    .RESET_B(net984),
    .D(\u_top_module.u_buffer.shift_reg_2[55] ),
    .Q_N(_1099_),
    .Q(\u_top_module.u_buffer.shift_reg_2[56] ));
 sg13g2_dfrbp_1 _2279_ (.CLK(net831),
    .RESET_B(net984),
    .D(\u_top_module.u_buffer.shift_reg_2[56] ),
    .Q_N(_1100_),
    .Q(\u_top_module.u_buffer.shift_reg_2[57] ));
 sg13g2_dfrbp_1 _2280_ (.CLK(net831),
    .RESET_B(net984),
    .D(\u_top_module.u_buffer.shift_reg_2[57] ),
    .Q_N(_1101_),
    .Q(\u_top_module.u_buffer.shift_reg_2[58] ));
 sg13g2_dfrbp_1 _2281_ (.CLK(net834),
    .RESET_B(net978),
    .D(\u_top_module.u_buffer.shift_reg_2[58] ),
    .Q_N(_1102_),
    .Q(\u_top_module.u_buffer.shift_reg_2[59] ));
 sg13g2_dfrbp_1 _2282_ (.CLK(net824),
    .RESET_B(net978),
    .D(\u_top_module.u_buffer.shift_reg_2[59] ),
    .Q_N(_1103_),
    .Q(\u_top_module.u_buffer.shift_reg_2[60] ));
 sg13g2_dfrbp_1 _2283_ (.CLK(net831),
    .RESET_B(net977),
    .D(\u_top_module.u_buffer.shift_reg_2[60] ),
    .Q_N(_1104_),
    .Q(\u_top_module.u_buffer.shift_reg_2[61] ));
 sg13g2_dfrbp_1 _2284_ (.CLK(net835),
    .RESET_B(net988),
    .D(\u_top_module.u_buffer.shift_reg_2[61] ),
    .Q_N(_1105_),
    .Q(\u_top_module.u_buffer.shift_reg_2[62] ));
 sg13g2_dfrbp_1 _2285_ (.CLK(net835),
    .RESET_B(net988),
    .D(\u_top_module.u_buffer.shift_reg_2[62] ),
    .Q_N(_1106_),
    .Q(\u_top_module.u_buffer.shift_reg_2[63] ));
 sg13g2_dfrbp_1 _2286_ (.CLK(net835),
    .RESET_B(net989),
    .D(\u_top_module.u_buffer.shift_reg_2[63] ),
    .Q_N(_1107_),
    .Q(\u_top_module.u_buffer.shift_reg_2[64] ));
 sg13g2_dfrbp_1 _2287_ (.CLK(net835),
    .RESET_B(net989),
    .D(\u_top_module.u_buffer.shift_reg_2[64] ),
    .Q_N(_1108_),
    .Q(\u_top_module.u_buffer.shift_reg_2[65] ));
 sg13g2_dfrbp_1 _2288_ (.CLK(net835),
    .RESET_B(net988),
    .D(\u_top_module.u_buffer.shift_reg_2[65] ),
    .Q_N(_1109_),
    .Q(\u_top_module.u_buffer.shift_reg_2[66] ));
 sg13g2_dfrbp_1 _2289_ (.CLK(net837),
    .RESET_B(net988),
    .D(\u_top_module.u_buffer.shift_reg_2[66] ),
    .Q_N(_1110_),
    .Q(\u_top_module.u_buffer.shift_reg_2[67] ));
 sg13g2_dfrbp_1 _2290_ (.CLK(net837),
    .RESET_B(net988),
    .D(\u_top_module.u_buffer.shift_reg_2[67] ),
    .Q_N(_1111_),
    .Q(\u_top_module.u_buffer.shift_reg_2[68] ));
 sg13g2_dfrbp_1 _2291_ (.CLK(net837),
    .RESET_B(net988),
    .D(\u_top_module.u_buffer.shift_reg_2[68] ),
    .Q_N(_1112_),
    .Q(\u_top_module.u_buffer.shift_reg_2[69] ));
 sg13g2_dfrbp_1 _2292_ (.CLK(net835),
    .RESET_B(net988),
    .D(\u_top_module.u_buffer.shift_reg_2[69] ),
    .Q_N(_1113_),
    .Q(\u_top_module.u_buffer.shift_reg_2[70] ));
 sg13g2_dfrbp_1 _2293_ (.CLK(net835),
    .RESET_B(net988),
    .D(\u_top_module.u_buffer.shift_reg_2[70] ),
    .Q_N(_1114_),
    .Q(\u_top_module.u_buffer.shift_reg_2[71] ));
 sg13g2_dfrbp_1 _2294_ (.CLK(net836),
    .RESET_B(net992),
    .D(\u_top_module.u_buffer.shift_reg_2[71] ),
    .Q_N(_1115_),
    .Q(\u_top_module.u_buffer.shift_reg_2[72] ));
 sg13g2_dfrbp_1 _2295_ (.CLK(net836),
    .RESET_B(net989),
    .D(\u_top_module.u_buffer.shift_reg_2[72] ),
    .Q_N(_1116_),
    .Q(\u_top_module.u_buffer.shift_reg_2[73] ));
 sg13g2_dfrbp_1 _2296_ (.CLK(net836),
    .RESET_B(net992),
    .D(\u_top_module.u_buffer.shift_reg_2[73] ),
    .Q_N(_1117_),
    .Q(\u_top_module.u_buffer.shift_reg_2[74] ));
 sg13g2_dfrbp_1 _2297_ (.CLK(net836),
    .RESET_B(net989),
    .D(\u_top_module.u_buffer.shift_reg_2[74] ),
    .Q_N(_1118_),
    .Q(\u_top_module.u_buffer.shift_reg_2[75] ));
 sg13g2_dfrbp_1 _2298_ (.CLK(net835),
    .RESET_B(net989),
    .D(\u_top_module.u_buffer.shift_reg_2[75] ),
    .Q_N(_1119_),
    .Q(\u_top_module.u_buffer.shift_reg_2[76] ));
 sg13g2_dfrbp_1 _2299_ (.CLK(net836),
    .RESET_B(net989),
    .D(\u_top_module.u_buffer.shift_reg_2[76] ),
    .Q_N(_1120_),
    .Q(\u_top_module.u_buffer.shift_reg_2[77] ));
 sg13g2_dfrbp_1 _2300_ (.CLK(net836),
    .RESET_B(net989),
    .D(\u_top_module.u_buffer.shift_reg_2[77] ),
    .Q_N(_1121_),
    .Q(\u_top_module.u_buffer.shift_reg_2[78] ));
 sg13g2_dfrbp_1 _2301_ (.CLK(net848),
    .RESET_B(net1001),
    .D(\u_top_module.u_buffer.shift_reg_2[78] ),
    .Q_N(_1122_),
    .Q(\u_top_module.u_buffer.shift_reg_2[79] ));
 sg13g2_dfrbp_1 _2302_ (.CLK(net848),
    .RESET_B(net1001),
    .D(\u_top_module.u_buffer.shift_reg_2[79] ),
    .Q_N(_1123_),
    .Q(\u_top_module.u_buffer.shift_reg_2[80] ));
 sg13g2_dfrbp_1 _2303_ (.CLK(net848),
    .RESET_B(net1001),
    .D(\u_top_module.u_buffer.shift_reg_2[80] ),
    .Q_N(_1124_),
    .Q(\u_top_module.u_buffer.shift_reg_2[81] ));
 sg13g2_dfrbp_1 _2304_ (.CLK(net841),
    .RESET_B(net995),
    .D(\u_top_module.u_buffer.shift_reg_2[81] ),
    .Q_N(_1125_),
    .Q(\u_top_module.u_buffer.shift_reg_2[82] ));
 sg13g2_dfrbp_1 _2305_ (.CLK(net841),
    .RESET_B(net995),
    .D(\u_top_module.u_buffer.shift_reg_2[82] ),
    .Q_N(_1126_),
    .Q(\u_top_module.u_buffer.shift_reg_2[83] ));
 sg13g2_dfrbp_1 _2306_ (.CLK(net841),
    .RESET_B(net995),
    .D(\u_top_module.u_buffer.shift_reg_2[83] ),
    .Q_N(_1127_),
    .Q(\u_top_module.u_buffer.shift_reg_2[84] ));
 sg13g2_dfrbp_1 _2307_ (.CLK(net841),
    .RESET_B(net995),
    .D(\u_top_module.u_buffer.shift_reg_2[84] ),
    .Q_N(_1128_),
    .Q(\u_top_module.u_buffer.shift_reg_2[85] ));
 sg13g2_dfrbp_1 _2308_ (.CLK(net841),
    .RESET_B(net995),
    .D(\u_top_module.u_buffer.shift_reg_2[85] ),
    .Q_N(_1129_),
    .Q(\u_top_module.u_buffer.shift_reg_2[86] ));
 sg13g2_dfrbp_1 _2309_ (.CLK(net841),
    .RESET_B(net995),
    .D(\u_top_module.u_buffer.shift_reg_2[86] ),
    .Q_N(_1130_),
    .Q(\u_top_module.u_buffer.shift_reg_2[87] ));
 sg13g2_dfrbp_1 _2310_ (.CLK(net828),
    .RESET_B(net981),
    .D(\u_top_module.u_buffer.shift_reg_2[87] ),
    .Q_N(_1131_),
    .Q(\u_top_module.u_buffer.shift_reg_2[88] ));
 sg13g2_dfrbp_1 _2311_ (.CLK(net829),
    .RESET_B(net982),
    .D(\u_top_module.u_buffer.shift_reg_2[88] ),
    .Q_N(_1132_),
    .Q(\u_top_module.u_buffer.shift_reg_2[89] ));
 sg13g2_dfrbp_1 _2312_ (.CLK(net828),
    .RESET_B(net981),
    .D(\u_top_module.u_buffer.shift_reg_2[89] ),
    .Q_N(_1133_),
    .Q(\u_top_module.u_buffer.shift_reg_2[90] ));
 sg13g2_dfrbp_1 _2313_ (.CLK(net828),
    .RESET_B(net981),
    .D(\u_top_module.u_buffer.shift_reg_2[90] ),
    .Q_N(_1134_),
    .Q(\u_top_module.u_buffer.shift_reg_2[91] ));
 sg13g2_dfrbp_1 _2314_ (.CLK(net828),
    .RESET_B(net981),
    .D(\u_top_module.u_buffer.shift_reg_2[91] ),
    .Q_N(_1135_),
    .Q(\u_top_module.u_buffer.shift_reg_2[92] ));
 sg13g2_dfrbp_1 _2315_ (.CLK(net829),
    .RESET_B(net982),
    .D(\u_top_module.u_buffer.shift_reg_2[92] ),
    .Q_N(_1136_),
    .Q(\u_top_module.u_buffer.shift_reg_2[93] ));
 sg13g2_dfrbp_1 _2316_ (.CLK(net829),
    .RESET_B(net982),
    .D(\u_top_module.u_buffer.shift_reg_2[93] ),
    .Q_N(_1137_),
    .Q(\u_top_module.u_buffer.shift_reg_2[94] ));
 sg13g2_dfrbp_1 _2317_ (.CLK(net840),
    .RESET_B(net994),
    .D(\u_top_module.u_buffer.shift_reg_2[94] ),
    .Q_N(_1138_),
    .Q(\u_top_module.u_buffer.shift_reg_2[95] ));
 sg13g2_dfrbp_1 _2318_ (.CLK(net839),
    .RESET_B(net993),
    .D(\u_top_module.u_buffer.shift_reg_2[95] ),
    .Q_N(_1139_),
    .Q(\u_top_module.u_buffer.shift_reg_2[96] ));
 sg13g2_dfrbp_1 _2319_ (.CLK(net839),
    .RESET_B(net993),
    .D(\u_top_module.u_buffer.shift_reg_2[96] ),
    .Q_N(_1140_),
    .Q(\u_top_module.u_buffer.shift_reg_2[97] ));
 sg13g2_dfrbp_1 _2320_ (.CLK(net839),
    .RESET_B(net993),
    .D(\u_top_module.u_buffer.shift_reg_2[97] ),
    .Q_N(_0493_),
    .Q(\u_top_module.u_buffer.shift_reg_2[98] ));
 sg13g2_tiehi _1821__18 (.L_HI(net18));
 sg13g2_tiehi _1822__19 (.L_HI(net19));
 sg13g2_tiehi _1823__20 (.L_HI(net20));
 sg13g2_tiehi _1824__21 (.L_HI(net21));
 sg13g2_tiehi _1825__22 (.L_HI(net22));
 sg13g2_tiehi _1826__23 (.L_HI(net23));
 sg13g2_tiehi _1827__24 (.L_HI(net24));
 sg13g2_tiehi _1828__25 (.L_HI(net25));
 sg13g2_tiehi _1829__26 (.L_HI(net26));
 sg13g2_tiehi _1830__27 (.L_HI(net27));
 sg13g2_tiehi _1831__28 (.L_HI(net28));
 sg13g2_tiehi _1832__29 (.L_HI(net29));
 sg13g2_tiehi _1833__30 (.L_HI(net30));
 sg13g2_tiehi _1834__31 (.L_HI(net31));
 sg13g2_tiehi _1835__32 (.L_HI(net32));
 sg13g2_tiehi _1836__33 (.L_HI(net33));
 sg13g2_tiehi _1837__34 (.L_HI(net34));
 sg13g2_tiehi _1838__35 (.L_HI(net35));
 sg13g2_tiehi _1839__36 (.L_HI(net36));
 sg13g2_tiehi _1840__37 (.L_HI(net37));
 sg13g2_tiehi _1842__38 (.L_HI(net38));
 sg13g2_tiehi _1841__39 (.L_HI(net39));
 sg13g2_tiehi tt_um_pdm_correlator_arghunter_40 (.L_HI(net40));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tielo tt_um_pdm_correlator_arghunter_6 (.L_LO(net6));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_7 (.L_LO(net7));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_8 (.L_LO(net8));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_9 (.L_LO(net9));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_10 (.L_LO(net10));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_11 (.L_LO(net11));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_12 (.L_LO(net12));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_13 (.L_LO(net13));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_14 (.L_LO(net14));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_15 (.L_LO(net15));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_16 (.L_LO(net16));
 sg13g2_tiehi _1820__17 (.L_HI(net17));
 sg13g2_buf_1 _2357_ (.A(net967),
    .X(uio_out[0]));
 sg13g2_buf_1 _2358_ (.A(\u_top_module.pos ),
    .X(uio_out[1]));
 sg13g2_buf_1 _2359_ (.A(\u_top_module.neg ),
    .X(uio_out[2]));
 sg13g2_buf_2 fanout821 (.A(\u_top_module.u_buffer.corr_neg[5] ),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(net826),
    .X(net822));
 sg13g2_buf_1 fanout823 (.A(net826),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(net826),
    .X(net824));
 sg13g2_buf_1 fanout825 (.A(net826),
    .X(net825));
 sg13g2_buf_1 fanout826 (.A(net829),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(net828),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(net829),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(net855),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(net831),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(net834),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(net834),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(net834),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(net855),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(net838),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(net838),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(net838),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(net855),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(net840),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(net854),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(net845),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(net845),
    .X(net843));
 sg13g2_buf_1 fanout844 (.A(net845),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(net854),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(net853),
    .X(net846));
 sg13g2_buf_1 fanout847 (.A(net853),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(net853),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net852),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net852),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(net852),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net854),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(net855),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(\u_top_module.corr_dec_clk ),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(net857),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(net865),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(net865),
    .X(net858));
 sg13g2_buf_1 fanout859 (.A(net865),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net864),
    .X(net860));
 sg13g2_buf_1 fanout861 (.A(net864),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(net864),
    .X(net862));
 sg13g2_buf_1 fanout863 (.A(net864),
    .X(net863));
 sg13g2_buf_1 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_1 fanout865 (.A(net884),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(net867),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net874),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(net874),
    .X(net868));
 sg13g2_buf_1 fanout869 (.A(net874),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(net874),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(net874),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(net874),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net884),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(net876),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(net878),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(net879),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(net884),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(net881),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(net882),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(net883),
    .X(net882));
 sg13g2_buf_1 fanout883 (.A(net884),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(\u_top_module.corr_dec_clk ),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(net888),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(net888),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_1 fanout888 (.A(net893),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net893),
    .X(net889));
 sg13g2_buf_1 fanout890 (.A(net893),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(net892),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(net893),
    .X(net892));
 sg13g2_buf_1 fanout893 (.A(net912),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(net897),
    .X(net894));
 sg13g2_buf_1 fanout895 (.A(net897),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(net912),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(net899),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(net912),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(net902),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(net902),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(net912),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(net906),
    .X(net903));
 sg13g2_buf_1 fanout904 (.A(net906),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(net906),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(net912),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(net911),
    .X(net907));
 sg13g2_buf_1 fanout908 (.A(net909),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(net911),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(net911),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_4 fanout912 (.X(net912),
    .A(net917));
 sg13g2_buf_2 fanout913 (.A(net914),
    .X(net913));
 sg13g2_buf_1 fanout914 (.A(net917),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(net917),
    .X(net915));
 sg13g2_buf_1 fanout916 (.A(net917),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(\u_top_module.corr_dec_clk ),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(net919),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_0198_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(net922),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(net925),
    .X(net921));
 sg13g2_buf_1 fanout922 (.A(net925),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(net925),
    .X(net923));
 sg13g2_buf_1 fanout924 (.A(net925),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_0376_),
    .X(net925));
 sg13g2_buf_4 fanout926 (.X(net926),
    .A(_0212_));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(_0212_));
 sg13g2_buf_4 fanout928 (.X(net928),
    .A(_0203_));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(_0203_));
 sg13g2_buf_4 fanout930 (.X(net930),
    .A(net931));
 sg13g2_buf_4 fanout931 (.X(net931),
    .A(_0211_));
 sg13g2_buf_4 fanout932 (.X(net932),
    .A(_0210_));
 sg13g2_buf_4 fanout933 (.X(net933),
    .A(_0210_));
 sg13g2_buf_4 fanout934 (.X(net934),
    .A(_0208_));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(_0208_));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(_0205_));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(_0205_));
 sg13g2_buf_4 fanout938 (.X(net938),
    .A(net939));
 sg13g2_buf_4 fanout939 (.X(net939),
    .A(_0446_));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(net941));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(_0444_));
 sg13g2_buf_4 fanout942 (.X(net942),
    .A(_0442_));
 sg13g2_buf_4 fanout943 (.X(net943),
    .A(_0216_));
 sg13g2_buf_4 fanout944 (.X(net944),
    .A(_0216_));
 sg13g2_buf_2 fanout945 (.A(\u_top_module.capture_reg[7] ),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(\u_top_module.capture_reg[6] ),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(\u_top_module.capture_reg[5] ),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(\u_top_module.capture_reg[4] ),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(\u_top_module.capture_reg[3] ),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(\u_top_module.capture_reg[2] ),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(\u_top_module.capture_reg[1] ),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(\u_top_module.capture_reg[0] ),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(net955),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(net955),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(net958),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(net957),
    .X(net956));
 sg13g2_buf_1 fanout957 (.A(net958),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(net974),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(net960),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(net961),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(net974),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(net963),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(net974),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(net965),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(net968),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(net967),
    .X(net966));
 sg13g2_buf_1 fanout967 (.A(net968),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(net974),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(net971),
    .X(net969));
 sg13g2_buf_1 fanout970 (.A(net971),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(net972),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(net974),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(net974),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(ui_in[0]),
    .X(net974));
 sg13g2_buf_4 fanout975 (.X(net975),
    .A(net979));
 sg13g2_buf_2 fanout976 (.A(net979),
    .X(net976));
 sg13g2_buf_4 fanout977 (.X(net977),
    .A(net979));
 sg13g2_buf_4 fanout978 (.X(net978),
    .A(net979));
 sg13g2_buf_2 fanout979 (.A(net982),
    .X(net979));
 sg13g2_buf_4 fanout980 (.X(net980),
    .A(net981));
 sg13g2_buf_4 fanout981 (.X(net981),
    .A(net982));
 sg13g2_buf_2 fanout982 (.A(net1009),
    .X(net982));
 sg13g2_buf_4 fanout983 (.X(net983),
    .A(net984));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(net987));
 sg13g2_buf_4 fanout985 (.X(net985),
    .A(net986));
 sg13g2_buf_4 fanout986 (.X(net986),
    .A(net987));
 sg13g2_buf_2 fanout987 (.A(net1009),
    .X(net987));
 sg13g2_buf_4 fanout988 (.X(net988),
    .A(net989));
 sg13g2_buf_4 fanout989 (.X(net989),
    .A(net992));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(net992));
 sg13g2_buf_2 fanout991 (.A(net992),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(net1009),
    .X(net992));
 sg13g2_buf_4 fanout993 (.X(net993),
    .A(net994));
 sg13g2_buf_4 fanout994 (.X(net994),
    .A(net995));
 sg13g2_buf_4 fanout995 (.X(net995),
    .A(net1008));
 sg13g2_buf_4 fanout996 (.X(net996),
    .A(net999));
 sg13g2_buf_4 fanout997 (.X(net997),
    .A(net999));
 sg13g2_buf_4 fanout998 (.X(net998),
    .A(net999));
 sg13g2_buf_2 fanout999 (.A(net1008),
    .X(net999));
 sg13g2_buf_4 fanout1000 (.X(net1000),
    .A(net1001));
 sg13g2_buf_4 fanout1001 (.X(net1001),
    .A(net1002));
 sg13g2_buf_4 fanout1002 (.X(net1002),
    .A(net1008));
 sg13g2_buf_4 fanout1003 (.X(net1003),
    .A(net1007));
 sg13g2_buf_2 fanout1004 (.A(net1007),
    .X(net1004));
 sg13g2_buf_4 fanout1005 (.X(net1005),
    .A(net1007));
 sg13g2_buf_2 fanout1006 (.A(net1007),
    .X(net1006));
 sg13g2_buf_1 fanout1007 (.A(net1008),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(net1009),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(rst_n),
    .X(net1009));
 sg13g2_buf_4 fanout1010 (.X(net1010),
    .A(net1011));
 sg13g2_buf_4 fanout1011 (.X(net1011),
    .A(net1018));
 sg13g2_buf_4 fanout1012 (.X(net1012),
    .A(net1018));
 sg13g2_buf_2 fanout1013 (.A(net1018),
    .X(net1013));
 sg13g2_buf_4 fanout1014 (.X(net1014),
    .A(net1017));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(net1016));
 sg13g2_buf_4 fanout1016 (.X(net1016),
    .A(net1017));
 sg13g2_buf_2 fanout1017 (.A(net1018),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(net1039),
    .X(net1018));
 sg13g2_buf_4 fanout1019 (.X(net1019),
    .A(net1020));
 sg13g2_buf_4 fanout1020 (.X(net1020),
    .A(net1026));
 sg13g2_buf_4 fanout1021 (.X(net1021),
    .A(net1026));
 sg13g2_buf_4 fanout1022 (.X(net1022),
    .A(net1023));
 sg13g2_buf_4 fanout1023 (.X(net1023),
    .A(net1025));
 sg13g2_buf_4 fanout1024 (.X(net1024),
    .A(net1025));
 sg13g2_buf_2 fanout1025 (.A(net1026),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(net1039),
    .X(net1026));
 sg13g2_buf_4 fanout1027 (.X(net1027),
    .A(net1028));
 sg13g2_buf_2 fanout1028 (.A(net1030),
    .X(net1028));
 sg13g2_buf_4 fanout1029 (.X(net1029),
    .A(net1030));
 sg13g2_buf_2 fanout1030 (.A(net1039),
    .X(net1030));
 sg13g2_buf_4 fanout1031 (.X(net1031),
    .A(net1033));
 sg13g2_buf_4 fanout1032 (.X(net1032),
    .A(net1033));
 sg13g2_buf_4 fanout1033 (.X(net1033),
    .A(net1039));
 sg13g2_buf_4 fanout1034 (.X(net1034),
    .A(net1038));
 sg13g2_buf_2 fanout1035 (.A(net1036),
    .X(net1035));
 sg13g2_buf_4 fanout1036 (.X(net1036),
    .A(net1038));
 sg13g2_buf_4 fanout1037 (.X(net1037),
    .A(net1038));
 sg13g2_buf_2 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(rst_n),
    .X(net1039));
 sg13g2_buf_4 fanout1040 (.X(net1040),
    .A(net1041));
 sg13g2_buf_4 fanout1041 (.X(net1041),
    .A(net1043));
 sg13g2_buf_4 fanout1042 (.X(net1042),
    .A(net1043));
 sg13g2_buf_2 fanout1043 (.A(net1048),
    .X(net1043));
 sg13g2_buf_4 fanout1044 (.X(net1044),
    .A(net1048));
 sg13g2_buf_2 fanout1045 (.A(net1048),
    .X(net1045));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(net1047));
 sg13g2_buf_4 fanout1047 (.X(net1047),
    .A(net1048));
 sg13g2_buf_2 fanout1048 (.A(net1068),
    .X(net1048));
 sg13g2_buf_4 fanout1049 (.X(net1049),
    .A(net1051));
 sg13g2_buf_4 fanout1050 (.X(net1050),
    .A(net1051));
 sg13g2_buf_4 fanout1051 (.X(net1051),
    .A(net1068));
 sg13g2_buf_4 fanout1052 (.X(net1052),
    .A(net1053));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(net1068));
 sg13g2_buf_4 fanout1054 (.X(net1054),
    .A(net1056));
 sg13g2_buf_4 fanout1055 (.X(net1055),
    .A(net1056));
 sg13g2_buf_4 fanout1056 (.X(net1056),
    .A(net1068));
 sg13g2_buf_4 fanout1057 (.X(net1057),
    .A(net1061));
 sg13g2_buf_2 fanout1058 (.A(net1061),
    .X(net1058));
 sg13g2_buf_4 fanout1059 (.X(net1059),
    .A(net1061));
 sg13g2_buf_2 fanout1060 (.A(net1061),
    .X(net1060));
 sg13g2_buf_1 fanout1061 (.A(net1068),
    .X(net1061));
 sg13g2_buf_4 fanout1062 (.X(net1062),
    .A(net1065));
 sg13g2_buf_4 fanout1063 (.X(net1063),
    .A(net1065));
 sg13g2_buf_2 fanout1064 (.A(net1065),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(net1067),
    .X(net1065));
 sg13g2_buf_4 fanout1066 (.X(net1066),
    .A(net1067));
 sg13g2_buf_2 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(net1088));
 sg13g2_buf_4 fanout1069 (.X(net1069),
    .A(net1074));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(net1074));
 sg13g2_buf_4 fanout1071 (.X(net1071),
    .A(net1074));
 sg13g2_buf_4 fanout1072 (.X(net1072),
    .A(net1073));
 sg13g2_buf_4 fanout1073 (.X(net1073),
    .A(net1074));
 sg13g2_buf_2 fanout1074 (.A(net1088),
    .X(net1074));
 sg13g2_buf_4 fanout1075 (.X(net1075),
    .A(net1077));
 sg13g2_buf_4 fanout1076 (.X(net1076),
    .A(net1077));
 sg13g2_buf_2 fanout1077 (.A(net1088),
    .X(net1077));
 sg13g2_buf_4 fanout1078 (.X(net1078),
    .A(net1087));
 sg13g2_buf_4 fanout1079 (.X(net1079),
    .A(net1087));
 sg13g2_buf_4 fanout1080 (.X(net1080),
    .A(net1081));
 sg13g2_buf_4 fanout1081 (.X(net1081),
    .A(net1087));
 sg13g2_buf_4 fanout1082 (.X(net1082),
    .A(net1086));
 sg13g2_buf_4 fanout1083 (.X(net1083),
    .A(net1084));
 sg13g2_buf_2 fanout1084 (.A(net1085),
    .X(net1084));
 sg13g2_buf_4 fanout1085 (.X(net1085),
    .A(net1086));
 sg13g2_buf_2 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(net1088),
    .X(net1087));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_tielo tt_um_pdm_correlator_arghunter_5 (.L_LO(net5));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_fill_2 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_fill_2 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_4 FILLER_0_182 ();
 sg13g2_fill_1 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_fill_1 FILLER_0_246 ();
 sg13g2_fill_2 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_4 FILLER_0_308 ();
 sg13g2_fill_2 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_fill_2 FILLER_1_35 ();
 sg13g2_fill_1 FILLER_1_37 ();
 sg13g2_decap_8 FILLER_1_64 ();
 sg13g2_decap_4 FILLER_1_71 ();
 sg13g2_decap_4 FILLER_1_101 ();
 sg13g2_fill_2 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_237 ();
 sg13g2_fill_2 FILLER_1_244 ();
 sg13g2_decap_4 FILLER_1_298 ();
 sg13g2_decap_8 FILLER_1_328 ();
 sg13g2_decap_8 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_342 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_61 ();
 sg13g2_decap_4 FILLER_2_68 ();
 sg13g2_fill_1 FILLER_2_72 ();
 sg13g2_decap_8 FILLER_2_125 ();
 sg13g2_decap_4 FILLER_2_132 ();
 sg13g2_decap_8 FILLER_2_162 ();
 sg13g2_fill_1 FILLER_2_169 ();
 sg13g2_fill_2 FILLER_2_196 ();
 sg13g2_fill_1 FILLER_2_198 ();
 sg13g2_decap_8 FILLER_2_225 ();
 sg13g2_decap_8 FILLER_2_232 ();
 sg13g2_decap_8 FILLER_2_239 ();
 sg13g2_decap_4 FILLER_2_246 ();
 sg13g2_fill_1 FILLER_2_250 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_fill_1 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_337 ();
 sg13g2_decap_8 FILLER_2_344 ();
 sg13g2_decap_8 FILLER_2_351 ();
 sg13g2_decap_8 FILLER_2_358 ();
 sg13g2_decap_8 FILLER_2_365 ();
 sg13g2_decap_8 FILLER_2_372 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_fill_2 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_110 ();
 sg13g2_decap_8 FILLER_3_117 ();
 sg13g2_decap_4 FILLER_3_124 ();
 sg13g2_fill_1 FILLER_3_128 ();
 sg13g2_decap_8 FILLER_3_155 ();
 sg13g2_decap_4 FILLER_3_162 ();
 sg13g2_decap_4 FILLER_3_192 ();
 sg13g2_fill_1 FILLER_3_196 ();
 sg13g2_fill_2 FILLER_3_223 ();
 sg13g2_fill_1 FILLER_3_225 ();
 sg13g2_decap_4 FILLER_3_278 ();
 sg13g2_fill_1 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_335 ();
 sg13g2_decap_8 FILLER_3_342 ();
 sg13g2_decap_8 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_356 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_61 ();
 sg13g2_fill_1 FILLER_4_68 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_fill_2 FILLER_4_109 ();
 sg13g2_fill_1 FILLER_4_111 ();
 sg13g2_decap_4 FILLER_4_138 ();
 sg13g2_fill_1 FILLER_4_142 ();
 sg13g2_fill_2 FILLER_4_195 ();
 sg13g2_fill_1 FILLER_4_197 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_4 FILLER_5_28 ();
 sg13g2_fill_2 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_fill_2 FILLER_5_67 ();
 sg13g2_fill_1 FILLER_5_69 ();
 sg13g2_decap_8 FILLER_5_96 ();
 sg13g2_decap_4 FILLER_5_103 ();
 sg13g2_decap_4 FILLER_5_159 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_4 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_264 ();
 sg13g2_decap_8 FILLER_5_271 ();
 sg13g2_fill_2 FILLER_5_278 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_4 FILLER_5_403 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_fill_1 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_76 ();
 sg13g2_fill_2 FILLER_6_83 ();
 sg13g2_fill_1 FILLER_6_85 ();
 sg13g2_fill_1 FILLER_6_117 ();
 sg13g2_decap_8 FILLER_6_204 ();
 sg13g2_decap_8 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_218 ();
 sg13g2_decap_8 FILLER_6_225 ();
 sg13g2_decap_8 FILLER_6_240 ();
 sg13g2_decap_8 FILLER_6_247 ();
 sg13g2_decap_8 FILLER_6_254 ();
 sg13g2_decap_8 FILLER_6_261 ();
 sg13g2_decap_8 FILLER_6_268 ();
 sg13g2_decap_8 FILLER_6_275 ();
 sg13g2_decap_8 FILLER_6_282 ();
 sg13g2_decap_8 FILLER_6_289 ();
 sg13g2_decap_8 FILLER_6_296 ();
 sg13g2_decap_8 FILLER_6_303 ();
 sg13g2_decap_8 FILLER_6_310 ();
 sg13g2_decap_8 FILLER_6_317 ();
 sg13g2_fill_1 FILLER_6_324 ();
 sg13g2_fill_1 FILLER_6_351 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_4 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_32 ();
 sg13g2_decap_8 FILLER_7_60 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_4 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_152 ();
 sg13g2_decap_8 FILLER_7_159 ();
 sg13g2_decap_8 FILLER_7_166 ();
 sg13g2_decap_8 FILLER_7_173 ();
 sg13g2_decap_8 FILLER_7_180 ();
 sg13g2_decap_8 FILLER_7_187 ();
 sg13g2_decap_8 FILLER_7_194 ();
 sg13g2_decap_8 FILLER_7_201 ();
 sg13g2_decap_8 FILLER_7_208 ();
 sg13g2_decap_8 FILLER_7_215 ();
 sg13g2_decap_8 FILLER_7_222 ();
 sg13g2_decap_8 FILLER_7_229 ();
 sg13g2_decap_8 FILLER_7_236 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_decap_8 FILLER_7_250 ();
 sg13g2_fill_2 FILLER_7_257 ();
 sg13g2_fill_1 FILLER_7_259 ();
 sg13g2_decap_4 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_272 ();
 sg13g2_decap_8 FILLER_7_299 ();
 sg13g2_fill_1 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_338 ();
 sg13g2_decap_8 FILLER_7_345 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_359 ();
 sg13g2_decap_8 FILLER_7_366 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_8 FILLER_7_380 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_76 ();
 sg13g2_decap_8 FILLER_8_83 ();
 sg13g2_decap_4 FILLER_8_90 ();
 sg13g2_fill_1 FILLER_8_94 ();
 sg13g2_decap_8 FILLER_8_152 ();
 sg13g2_decap_8 FILLER_8_159 ();
 sg13g2_decap_8 FILLER_8_166 ();
 sg13g2_decap_8 FILLER_8_173 ();
 sg13g2_decap_8 FILLER_8_180 ();
 sg13g2_decap_4 FILLER_8_239 ();
 sg13g2_fill_1 FILLER_8_243 ();
 sg13g2_fill_1 FILLER_8_322 ();
 sg13g2_fill_2 FILLER_8_331 ();
 sg13g2_fill_1 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_367 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_fill_2 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_78 ();
 sg13g2_fill_1 FILLER_9_89 ();
 sg13g2_fill_1 FILLER_9_116 ();
 sg13g2_decap_8 FILLER_9_169 ();
 sg13g2_decap_8 FILLER_9_176 ();
 sg13g2_fill_2 FILLER_9_183 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_37 ();
 sg13g2_decap_8 FILLER_10_44 ();
 sg13g2_decap_8 FILLER_10_107 ();
 sg13g2_fill_1 FILLER_10_114 ();
 sg13g2_fill_2 FILLER_10_120 ();
 sg13g2_fill_1 FILLER_10_153 ();
 sg13g2_decap_8 FILLER_10_206 ();
 sg13g2_fill_1 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_4 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_14 ();
 sg13g2_decap_4 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_46 ();
 sg13g2_fill_2 FILLER_11_83 ();
 sg13g2_decap_4 FILLER_11_93 ();
 sg13g2_decap_4 FILLER_11_227 ();
 sg13g2_fill_2 FILLER_11_231 ();
 sg13g2_fill_2 FILLER_11_238 ();
 sg13g2_fill_1 FILLER_11_245 ();
 sg13g2_fill_2 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_260 ();
 sg13g2_decap_8 FILLER_11_272 ();
 sg13g2_decap_8 FILLER_11_279 ();
 sg13g2_decap_8 FILLER_11_286 ();
 sg13g2_decap_8 FILLER_11_293 ();
 sg13g2_fill_2 FILLER_11_300 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_fill_1 FILLER_11_354 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_4 FILLER_12_21 ();
 sg13g2_decap_4 FILLER_12_51 ();
 sg13g2_fill_2 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_124 ();
 sg13g2_decap_8 FILLER_12_131 ();
 sg13g2_decap_8 FILLER_12_138 ();
 sg13g2_decap_4 FILLER_12_145 ();
 sg13g2_fill_2 FILLER_12_149 ();
 sg13g2_decap_8 FILLER_12_177 ();
 sg13g2_decap_8 FILLER_12_184 ();
 sg13g2_decap_8 FILLER_12_191 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_decap_8 FILLER_12_205 ();
 sg13g2_decap_8 FILLER_12_212 ();
 sg13g2_decap_8 FILLER_12_219 ();
 sg13g2_decap_8 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_233 ();
 sg13g2_decap_8 FILLER_12_240 ();
 sg13g2_decap_8 FILLER_12_247 ();
 sg13g2_decap_8 FILLER_12_254 ();
 sg13g2_decap_8 FILLER_12_261 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_decap_4 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_4 FILLER_12_333 ();
 sg13g2_fill_1 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_4 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_25 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_fill_2 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_fill_1 FILLER_13_85 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_105 ();
 sg13g2_fill_1 FILLER_13_107 ();
 sg13g2_decap_8 FILLER_13_113 ();
 sg13g2_decap_8 FILLER_13_120 ();
 sg13g2_fill_2 FILLER_13_127 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_decap_8 FILLER_13_138 ();
 sg13g2_decap_8 FILLER_13_145 ();
 sg13g2_fill_1 FILLER_13_152 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_fill_2 FILLER_13_170 ();
 sg13g2_fill_2 FILLER_13_224 ();
 sg13g2_fill_2 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_34 ();
 sg13g2_decap_8 FILLER_14_41 ();
 sg13g2_decap_8 FILLER_14_48 ();
 sg13g2_decap_8 FILLER_14_55 ();
 sg13g2_decap_8 FILLER_14_62 ();
 sg13g2_decap_8 FILLER_14_69 ();
 sg13g2_decap_8 FILLER_14_76 ();
 sg13g2_decap_8 FILLER_14_83 ();
 sg13g2_fill_2 FILLER_14_90 ();
 sg13g2_fill_1 FILLER_14_92 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_4 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_187 ();
 sg13g2_fill_1 FILLER_15_194 ();
 sg13g2_fill_2 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_fill_1 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_7 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_fill_1 FILLER_16_142 ();
 sg13g2_decap_4 FILLER_16_156 ();
 sg13g2_fill_1 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_178 ();
 sg13g2_decap_8 FILLER_16_185 ();
 sg13g2_decap_8 FILLER_16_192 ();
 sg13g2_decap_8 FILLER_16_199 ();
 sg13g2_decap_8 FILLER_16_206 ();
 sg13g2_decap_8 FILLER_16_213 ();
 sg13g2_fill_2 FILLER_16_220 ();
 sg13g2_fill_1 FILLER_16_222 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_4 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_decap_4 FILLER_16_255 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_fill_1 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_fill_1 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_4 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_25 ();
 sg13g2_fill_1 FILLER_17_83 ();
 sg13g2_decap_8 FILLER_17_110 ();
 sg13g2_decap_8 FILLER_17_117 ();
 sg13g2_decap_8 FILLER_17_124 ();
 sg13g2_decap_4 FILLER_17_131 ();
 sg13g2_fill_2 FILLER_17_135 ();
 sg13g2_fill_1 FILLER_17_163 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_fill_2 FILLER_17_178 ();
 sg13g2_fill_1 FILLER_17_180 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_225 ();
 sg13g2_decap_8 FILLER_17_232 ();
 sg13g2_decap_4 FILLER_17_239 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_4 FILLER_17_319 ();
 sg13g2_fill_2 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_fill_1 FILLER_17_345 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_93 ();
 sg13g2_fill_2 FILLER_18_100 ();
 sg13g2_fill_1 FILLER_18_102 ();
 sg13g2_decap_4 FILLER_18_129 ();
 sg13g2_fill_2 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_213 ();
 sg13g2_fill_1 FILLER_18_215 ();
 sg13g2_fill_1 FILLER_18_242 ();
 sg13g2_fill_2 FILLER_18_251 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_fill_2 FILLER_18_286 ();
 sg13g2_fill_1 FILLER_18_288 ();
 sg13g2_fill_2 FILLER_18_367 ();
 sg13g2_fill_1 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_4 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_47 ();
 sg13g2_decap_4 FILLER_19_54 ();
 sg13g2_fill_1 FILLER_19_58 ();
 sg13g2_decap_4 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_89 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_14 ();
 sg13g2_fill_2 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_fill_2 FILLER_20_67 ();
 sg13g2_fill_1 FILLER_20_69 ();
 sg13g2_fill_2 FILLER_20_148 ();
 sg13g2_decap_8 FILLER_20_155 ();
 sg13g2_fill_2 FILLER_20_162 ();
 sg13g2_fill_1 FILLER_20_164 ();
 sg13g2_decap_8 FILLER_20_191 ();
 sg13g2_fill_1 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_20_251 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_293 ();
 sg13g2_decap_4 FILLER_20_346 ();
 sg13g2_fill_2 FILLER_20_350 ();
 sg13g2_decap_4 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_4 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_32 ();
 sg13g2_decap_8 FILLER_21_59 ();
 sg13g2_decap_8 FILLER_21_66 ();
 sg13g2_decap_8 FILLER_21_73 ();
 sg13g2_fill_1 FILLER_21_80 ();
 sg13g2_decap_4 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_fill_2 FILLER_21_138 ();
 sg13g2_decap_8 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_180 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_215 ();
 sg13g2_decap_8 FILLER_21_222 ();
 sg13g2_decap_8 FILLER_21_229 ();
 sg13g2_decap_8 FILLER_21_236 ();
 sg13g2_decap_8 FILLER_21_243 ();
 sg13g2_decap_8 FILLER_21_250 ();
 sg13g2_decap_8 FILLER_21_257 ();
 sg13g2_decap_8 FILLER_21_264 ();
 sg13g2_decap_8 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_278 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_decap_4 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_65 ();
 sg13g2_decap_8 FILLER_22_72 ();
 sg13g2_fill_1 FILLER_22_79 ();
 sg13g2_decap_8 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_113 ();
 sg13g2_decap_8 FILLER_22_120 ();
 sg13g2_decap_8 FILLER_22_127 ();
 sg13g2_fill_2 FILLER_22_134 ();
 sg13g2_decap_8 FILLER_22_162 ();
 sg13g2_decap_8 FILLER_22_169 ();
 sg13g2_decap_8 FILLER_22_176 ();
 sg13g2_decap_8 FILLER_22_183 ();
 sg13g2_decap_8 FILLER_22_190 ();
 sg13g2_decap_4 FILLER_22_197 ();
 sg13g2_decap_4 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_fill_2 FILLER_22_219 ();
 sg13g2_fill_1 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_227 ();
 sg13g2_decap_8 FILLER_22_234 ();
 sg13g2_decap_8 FILLER_22_241 ();
 sg13g2_decap_4 FILLER_22_248 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_fill_1 FILLER_22_355 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_41 ();
 sg13g2_decap_8 FILLER_23_48 ();
 sg13g2_decap_8 FILLER_23_107 ();
 sg13g2_decap_8 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_121 ();
 sg13g2_decap_8 FILLER_23_128 ();
 sg13g2_decap_4 FILLER_23_135 ();
 sg13g2_fill_2 FILLER_23_139 ();
 sg13g2_decap_8 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_174 ();
 sg13g2_decap_4 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_fill_2 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_266 ();
 sg13g2_fill_2 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_354 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_47 ();
 sg13g2_fill_1 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_107 ();
 sg13g2_decap_8 FILLER_24_134 ();
 sg13g2_decap_8 FILLER_24_141 ();
 sg13g2_decap_8 FILLER_24_148 ();
 sg13g2_decap_8 FILLER_24_155 ();
 sg13g2_fill_2 FILLER_24_162 ();
 sg13g2_fill_1 FILLER_24_164 ();
 sg13g2_fill_2 FILLER_24_295 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_fill_2 FILLER_24_363 ();
 sg13g2_fill_1 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_4 FILLER_24_378 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_77 ();
 sg13g2_fill_1 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_fill_1 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_decap_4 FILLER_25_284 ();
 sg13g2_fill_2 FILLER_25_288 ();
 sg13g2_decap_8 FILLER_25_298 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_4 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_fill_2 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_fill_1 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_69 ();
 sg13g2_decap_8 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_83 ();
 sg13g2_decap_8 FILLER_26_89 ();
 sg13g2_decap_8 FILLER_26_96 ();
 sg13g2_decap_4 FILLER_26_103 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_173 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_262 ();
 sg13g2_decap_8 FILLER_26_269 ();
 sg13g2_decap_8 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_290 ();
 sg13g2_decap_4 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_25 ();
 sg13g2_decap_4 FILLER_27_52 ();
 sg13g2_decap_4 FILLER_27_90 ();
 sg13g2_decap_8 FILLER_27_125 ();
 sg13g2_decap_4 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_fill_2 FILLER_27_163 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_342 ();
 sg13g2_decap_4 FILLER_27_377 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_fill_1 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_88 ();
 sg13g2_decap_4 FILLER_28_97 ();
 sg13g2_decap_4 FILLER_28_106 ();
 sg13g2_decap_8 FILLER_28_149 ();
 sg13g2_decap_4 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_213 ();
 sg13g2_fill_2 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_234 ();
 sg13g2_decap_8 FILLER_28_240 ();
 sg13g2_decap_4 FILLER_28_247 ();
 sg13g2_fill_1 FILLER_28_251 ();
 sg13g2_decap_8 FILLER_28_257 ();
 sg13g2_fill_1 FILLER_28_315 ();
 sg13g2_decap_4 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_44 ();
 sg13g2_decap_8 FILLER_29_51 ();
 sg13g2_decap_8 FILLER_29_58 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_fill_1 FILLER_29_67 ();
 sg13g2_fill_2 FILLER_29_94 ();
 sg13g2_fill_1 FILLER_29_187 ();
 sg13g2_decap_4 FILLER_29_240 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_4 FILLER_29_259 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_decap_4 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_4 FILLER_30_70 ();
 sg13g2_fill_2 FILLER_30_74 ();
 sg13g2_decap_4 FILLER_30_162 ();
 sg13g2_fill_2 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_298 ();
 sg13g2_decap_8 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_355 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_82 ();
 sg13g2_decap_4 FILLER_31_89 ();
 sg13g2_fill_2 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_215 ();
 sg13g2_decap_4 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_253 ();
 sg13g2_decap_4 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_decap_4 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_324 ();
 sg13g2_fill_2 FILLER_31_331 ();
 sg13g2_fill_1 FILLER_31_333 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_31_400 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_89 ();
 sg13g2_decap_8 FILLER_32_96 ();
 sg13g2_decap_8 FILLER_32_108 ();
 sg13g2_decap_8 FILLER_32_115 ();
 sg13g2_decap_8 FILLER_32_122 ();
 sg13g2_decap_8 FILLER_32_129 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_174 ();
 sg13g2_decap_8 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_188 ();
 sg13g2_decap_8 FILLER_32_195 ();
 sg13g2_decap_8 FILLER_32_202 ();
 sg13g2_decap_8 FILLER_32_209 ();
 sg13g2_decap_4 FILLER_32_216 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_decap_4 FILLER_32_248 ();
 sg13g2_decap_4 FILLER_32_278 ();
 sg13g2_decap_8 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_299 ();
 sg13g2_fill_2 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_360 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_102 ();
 sg13g2_decap_8 FILLER_33_109 ();
 sg13g2_decap_8 FILLER_33_116 ();
 sg13g2_decap_8 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_130 ();
 sg13g2_fill_2 FILLER_33_137 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_decap_4 FILLER_33_150 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_decap_4 FILLER_33_159 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_decap_8 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_198 ();
 sg13g2_decap_8 FILLER_33_205 ();
 sg13g2_fill_2 FILLER_33_212 ();
 sg13g2_decap_8 FILLER_33_240 ();
 sg13g2_decap_4 FILLER_33_247 ();
 sg13g2_decap_4 FILLER_33_293 ();
 sg13g2_decap_8 FILLER_33_313 ();
 sg13g2_decap_8 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_decap_8 FILLER_33_356 ();
 sg13g2_decap_4 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_367 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_78 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_fill_1 FILLER_34_135 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_230 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_244 ();
 sg13g2_decap_8 FILLER_34_251 ();
 sg13g2_decap_8 FILLER_34_258 ();
 sg13g2_fill_2 FILLER_34_265 ();
 sg13g2_decap_8 FILLER_34_289 ();
 sg13g2_fill_2 FILLER_34_296 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_fill_2 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_57 ();
 sg13g2_decap_4 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_76 ();
 sg13g2_fill_1 FILLER_35_85 ();
 sg13g2_fill_2 FILLER_35_190 ();
 sg13g2_fill_1 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_219 ();
 sg13g2_decap_8 FILLER_35_226 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_decap_8 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_247 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_288 ();
 sg13g2_decap_8 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_26 ();
 sg13g2_decap_4 FILLER_36_33 ();
 sg13g2_fill_1 FILLER_36_37 ();
 sg13g2_fill_1 FILLER_36_68 ();
 sg13g2_decap_8 FILLER_36_95 ();
 sg13g2_decap_4 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_208 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_fill_2 FILLER_36_286 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_fill_2 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_40 ();
 sg13g2_fill_1 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_69 ();
 sg13g2_decap_4 FILLER_37_76 ();
 sg13g2_fill_1 FILLER_37_80 ();
 sg13g2_fill_2 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_109 ();
 sg13g2_decap_8 FILLER_37_136 ();
 sg13g2_decap_8 FILLER_37_143 ();
 sg13g2_decap_8 FILLER_37_150 ();
 sg13g2_decap_8 FILLER_37_157 ();
 sg13g2_fill_2 FILLER_37_164 ();
 sg13g2_decap_8 FILLER_37_171 ();
 sg13g2_fill_2 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_180 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_fill_1 FILLER_37_317 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_44 ();
 sg13g2_decap_8 FILLER_38_71 ();
 sg13g2_decap_8 FILLER_38_78 ();
 sg13g2_decap_8 FILLER_38_85 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_8 FILLER_38_122 ();
 sg13g2_decap_8 FILLER_38_129 ();
 sg13g2_decap_4 FILLER_38_136 ();
 sg13g2_decap_4 FILLER_38_145 ();
 sg13g2_fill_1 FILLER_38_149 ();
 sg13g2_fill_2 FILLER_38_233 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_fill_1 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_26 ();
 sg13g2_decap_8 FILLER_39_33 ();
 sg13g2_decap_4 FILLER_39_40 ();
 sg13g2_decap_4 FILLER_39_70 ();
 sg13g2_fill_1 FILLER_39_74 ();
 sg13g2_fill_2 FILLER_39_101 ();
 sg13g2_fill_1 FILLER_39_103 ();
 sg13g2_decap_4 FILLER_39_130 ();
 sg13g2_fill_2 FILLER_39_134 ();
 sg13g2_decap_8 FILLER_39_188 ();
 sg13g2_decap_8 FILLER_39_195 ();
 sg13g2_decap_8 FILLER_39_202 ();
 sg13g2_decap_8 FILLER_39_209 ();
 sg13g2_fill_1 FILLER_39_216 ();
 sg13g2_decap_8 FILLER_39_247 ();
 sg13g2_fill_2 FILLER_39_254 ();
 sg13g2_fill_1 FILLER_39_302 ();
 sg13g2_decap_8 FILLER_39_313 ();
 sg13g2_decap_4 FILLER_39_320 ();
 sg13g2_fill_1 FILLER_39_324 ();
 sg13g2_decap_8 FILLER_39_355 ();
 sg13g2_decap_8 FILLER_39_362 ();
 sg13g2_decap_8 FILLER_39_369 ();
 sg13g2_decap_8 FILLER_39_376 ();
 sg13g2_decap_8 FILLER_39_383 ();
 sg13g2_decap_8 FILLER_39_390 ();
 sg13g2_decap_8 FILLER_39_397 ();
 sg13g2_decap_4 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_26 ();
 sg13g2_decap_8 FILLER_40_33 ();
 sg13g2_decap_8 FILLER_40_40 ();
 sg13g2_decap_8 FILLER_40_47 ();
 sg13g2_decap_8 FILLER_40_54 ();
 sg13g2_decap_8 FILLER_40_61 ();
 sg13g2_decap_8 FILLER_40_68 ();
 sg13g2_decap_8 FILLER_40_75 ();
 sg13g2_decap_4 FILLER_40_82 ();
 sg13g2_decap_8 FILLER_40_216 ();
 sg13g2_decap_4 FILLER_40_223 ();
 sg13g2_fill_2 FILLER_40_227 ();
 sg13g2_decap_8 FILLER_40_244 ();
 sg13g2_decap_4 FILLER_40_251 ();
 sg13g2_fill_2 FILLER_40_255 ();
 sg13g2_fill_2 FILLER_40_283 ();
 sg13g2_fill_1 FILLER_40_285 ();
 sg13g2_fill_1 FILLER_40_291 ();
 sg13g2_decap_8 FILLER_40_297 ();
 sg13g2_decap_8 FILLER_40_304 ();
 sg13g2_fill_2 FILLER_40_337 ();
 sg13g2_decap_8 FILLER_40_365 ();
 sg13g2_decap_8 FILLER_40_372 ();
 sg13g2_decap_8 FILLER_40_379 ();
 sg13g2_decap_8 FILLER_40_386 ();
 sg13g2_decap_8 FILLER_40_393 ();
 sg13g2_decap_8 FILLER_40_400 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_4 FILLER_41_26 ();
 sg13g2_fill_2 FILLER_41_30 ();
 sg13g2_decap_8 FILLER_41_58 ();
 sg13g2_decap_8 FILLER_41_65 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_fill_1 FILLER_41_133 ();
 sg13g2_fill_1 FILLER_41_160 ();
 sg13g2_decap_4 FILLER_41_187 ();
 sg13g2_decap_4 FILLER_41_217 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_decap_8 FILLER_41_232 ();
 sg13g2_decap_8 FILLER_41_239 ();
 sg13g2_decap_8 FILLER_41_246 ();
 sg13g2_fill_2 FILLER_41_253 ();
 sg13g2_decap_8 FILLER_41_265 ();
 sg13g2_decap_8 FILLER_41_272 ();
 sg13g2_decap_8 FILLER_41_279 ();
 sg13g2_decap_8 FILLER_41_286 ();
 sg13g2_decap_4 FILLER_41_293 ();
 sg13g2_fill_2 FILLER_41_303 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_fill_1 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_347 ();
 sg13g2_decap_8 FILLER_41_354 ();
 sg13g2_decap_8 FILLER_41_361 ();
 sg13g2_decap_8 FILLER_41_368 ();
 sg13g2_decap_8 FILLER_41_375 ();
 sg13g2_decap_8 FILLER_41_382 ();
 sg13g2_decap_8 FILLER_41_389 ();
 sg13g2_decap_8 FILLER_41_396 ();
 sg13g2_decap_4 FILLER_41_403 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_9 ();
 sg13g2_decap_8 FILLER_42_44 ();
 sg13g2_fill_2 FILLER_42_51 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_fill_2 FILLER_42_133 ();
 sg13g2_fill_1 FILLER_42_135 ();
 sg13g2_decap_8 FILLER_42_162 ();
 sg13g2_decap_8 FILLER_42_169 ();
 sg13g2_decap_8 FILLER_42_176 ();
 sg13g2_decap_8 FILLER_42_183 ();
 sg13g2_fill_1 FILLER_42_190 ();
 sg13g2_fill_1 FILLER_42_217 ();
 sg13g2_decap_4 FILLER_42_244 ();
 sg13g2_fill_2 FILLER_42_248 ();
 sg13g2_fill_2 FILLER_42_265 ();
 sg13g2_decap_8 FILLER_42_277 ();
 sg13g2_fill_2 FILLER_42_284 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_fill_2 FILLER_42_327 ();
 sg13g2_fill_1 FILLER_42_329 ();
 sg13g2_fill_2 FILLER_42_340 ();
 sg13g2_decap_8 FILLER_42_368 ();
 sg13g2_decap_8 FILLER_42_375 ();
 sg13g2_decap_8 FILLER_42_382 ();
 sg13g2_decap_8 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_4 FILLER_42_403 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_fill_2 FILLER_43_26 ();
 sg13g2_fill_2 FILLER_43_54 ();
 sg13g2_decap_8 FILLER_43_82 ();
 sg13g2_decap_4 FILLER_43_89 ();
 sg13g2_decap_8 FILLER_43_145 ();
 sg13g2_decap_8 FILLER_43_152 ();
 sg13g2_fill_1 FILLER_43_159 ();
 sg13g2_decap_8 FILLER_43_186 ();
 sg13g2_decap_8 FILLER_43_193 ();
 sg13g2_decap_8 FILLER_43_200 ();
 sg13g2_decap_8 FILLER_43_207 ();
 sg13g2_fill_1 FILLER_43_214 ();
 sg13g2_decap_4 FILLER_43_303 ();
 sg13g2_fill_1 FILLER_43_307 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_fill_1 FILLER_44_57 ();
 sg13g2_decap_8 FILLER_44_144 ();
 sg13g2_decap_8 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_158 ();
 sg13g2_decap_8 FILLER_44_165 ();
 sg13g2_decap_4 FILLER_44_172 ();
 sg13g2_fill_2 FILLER_44_176 ();
 sg13g2_decap_8 FILLER_44_204 ();
 sg13g2_decap_8 FILLER_44_211 ();
 sg13g2_decap_4 FILLER_44_218 ();
 sg13g2_decap_8 FILLER_44_242 ();
 sg13g2_fill_2 FILLER_44_249 ();
 sg13g2_fill_1 FILLER_44_251 ();
 sg13g2_decap_8 FILLER_44_262 ();
 sg13g2_fill_2 FILLER_44_321 ();
 sg13g2_fill_1 FILLER_44_323 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_27 ();
 sg13g2_fill_1 FILLER_45_81 ();
 sg13g2_decap_4 FILLER_45_186 ();
 sg13g2_decap_8 FILLER_45_216 ();
 sg13g2_fill_2 FILLER_45_235 ();
 sg13g2_decap_8 FILLER_45_263 ();
 sg13g2_fill_2 FILLER_45_270 ();
 sg13g2_decap_8 FILLER_45_298 ();
 sg13g2_decap_8 FILLER_45_310 ();
 sg13g2_fill_2 FILLER_45_332 ();
 sg13g2_fill_1 FILLER_45_334 ();
 sg13g2_decap_8 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_347 ();
 sg13g2_decap_8 FILLER_45_354 ();
 sg13g2_decap_8 FILLER_45_361 ();
 sg13g2_decap_8 FILLER_45_368 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_382 ();
 sg13g2_decap_8 FILLER_45_389 ();
 sg13g2_decap_8 FILLER_45_396 ();
 sg13g2_decap_4 FILLER_45_403 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_4 FILLER_46_26 ();
 sg13g2_decap_8 FILLER_46_90 ();
 sg13g2_decap_8 FILLER_46_97 ();
 sg13g2_decap_8 FILLER_46_104 ();
 sg13g2_decap_8 FILLER_46_111 ();
 sg13g2_decap_8 FILLER_46_118 ();
 sg13g2_fill_1 FILLER_46_229 ();
 sg13g2_fill_2 FILLER_46_235 ();
 sg13g2_fill_2 FILLER_46_283 ();
 sg13g2_fill_1 FILLER_46_285 ();
 sg13g2_decap_8 FILLER_46_354 ();
 sg13g2_decap_8 FILLER_46_361 ();
 sg13g2_decap_8 FILLER_46_368 ();
 sg13g2_decap_8 FILLER_46_375 ();
 sg13g2_decap_8 FILLER_46_382 ();
 sg13g2_decap_8 FILLER_46_389 ();
 sg13g2_decap_8 FILLER_46_396 ();
 sg13g2_decap_4 FILLER_46_403 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_9 ();
 sg13g2_fill_1 FILLER_47_88 ();
 sg13g2_decap_8 FILLER_47_115 ();
 sg13g2_decap_8 FILLER_47_122 ();
 sg13g2_decap_4 FILLER_47_129 ();
 sg13g2_fill_1 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_138 ();
 sg13g2_decap_8 FILLER_47_145 ();
 sg13g2_fill_2 FILLER_47_157 ();
 sg13g2_fill_1 FILLER_47_159 ();
 sg13g2_decap_8 FILLER_47_186 ();
 sg13g2_decap_8 FILLER_47_193 ();
 sg13g2_decap_8 FILLER_47_200 ();
 sg13g2_fill_2 FILLER_47_207 ();
 sg13g2_fill_1 FILLER_47_209 ();
 sg13g2_fill_2 FILLER_47_228 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_fill_1 FILLER_47_264 ();
 sg13g2_fill_2 FILLER_47_286 ();
 sg13g2_fill_1 FILLER_47_288 ();
 sg13g2_fill_1 FILLER_47_305 ();
 sg13g2_decap_8 FILLER_47_314 ();
 sg13g2_fill_2 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_367 ();
 sg13g2_decap_8 FILLER_47_374 ();
 sg13g2_decap_8 FILLER_47_381 ();
 sg13g2_decap_8 FILLER_47_388 ();
 sg13g2_decap_8 FILLER_47_395 ();
 sg13g2_decap_8 FILLER_47_402 ();
 sg13g2_decap_4 FILLER_48_26 ();
 sg13g2_fill_2 FILLER_48_30 ();
 sg13g2_fill_2 FILLER_48_37 ();
 sg13g2_decap_8 FILLER_48_48 ();
 sg13g2_fill_2 FILLER_48_60 ();
 sg13g2_decap_8 FILLER_48_88 ();
 sg13g2_fill_2 FILLER_48_95 ();
 sg13g2_fill_1 FILLER_48_97 ();
 sg13g2_decap_4 FILLER_48_124 ();
 sg13g2_fill_2 FILLER_48_128 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_4 FILLER_48_175 ();
 sg13g2_fill_2 FILLER_48_179 ();
 sg13g2_decap_4 FILLER_48_243 ();
 sg13g2_fill_1 FILLER_48_247 ();
 sg13g2_decap_4 FILLER_48_258 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_decap_8 FILLER_48_304 ();
 sg13g2_decap_8 FILLER_48_311 ();
 sg13g2_decap_8 FILLER_48_318 ();
 sg13g2_decap_4 FILLER_48_325 ();
 sg13g2_fill_2 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_369 ();
 sg13g2_decap_8 FILLER_48_376 ();
 sg13g2_decap_8 FILLER_48_383 ();
 sg13g2_decap_8 FILLER_48_390 ();
 sg13g2_decap_8 FILLER_48_397 ();
 sg13g2_decap_4 FILLER_48_404 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_4 FILLER_49_56 ();
 sg13g2_fill_1 FILLER_49_60 ();
 sg13g2_decap_8 FILLER_49_65 ();
 sg13g2_decap_4 FILLER_49_72 ();
 sg13g2_fill_2 FILLER_49_76 ();
 sg13g2_fill_2 FILLER_49_161 ();
 sg13g2_fill_1 FILLER_49_163 ();
 sg13g2_decap_8 FILLER_49_198 ();
 sg13g2_decap_8 FILLER_49_205 ();
 sg13g2_fill_2 FILLER_49_212 ();
 sg13g2_fill_1 FILLER_49_214 ();
 sg13g2_decap_8 FILLER_49_223 ();
 sg13g2_decap_4 FILLER_49_230 ();
 sg13g2_decap_4 FILLER_49_260 ();
 sg13g2_fill_1 FILLER_49_264 ();
 sg13g2_fill_1 FILLER_49_297 ();
 sg13g2_decap_4 FILLER_49_345 ();
 sg13g2_fill_2 FILLER_49_349 ();
 sg13g2_decap_8 FILLER_49_355 ();
 sg13g2_decap_8 FILLER_49_362 ();
 sg13g2_decap_8 FILLER_49_369 ();
 sg13g2_decap_8 FILLER_49_376 ();
 sg13g2_decap_8 FILLER_49_383 ();
 sg13g2_decap_8 FILLER_49_390 ();
 sg13g2_decap_8 FILLER_49_397 ();
 sg13g2_decap_4 FILLER_49_404 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_14 ();
 sg13g2_fill_1 FILLER_50_46 ();
 sg13g2_decap_8 FILLER_50_55 ();
 sg13g2_decap_8 FILLER_50_62 ();
 sg13g2_decap_8 FILLER_50_69 ();
 sg13g2_decap_8 FILLER_50_76 ();
 sg13g2_fill_2 FILLER_50_83 ();
 sg13g2_fill_2 FILLER_50_111 ();
 sg13g2_fill_1 FILLER_50_113 ();
 sg13g2_fill_2 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_194 ();
 sg13g2_decap_8 FILLER_50_201 ();
 sg13g2_decap_8 FILLER_50_208 ();
 sg13g2_decap_8 FILLER_50_215 ();
 sg13g2_decap_4 FILLER_50_222 ();
 sg13g2_decap_8 FILLER_50_236 ();
 sg13g2_decap_8 FILLER_50_243 ();
 sg13g2_fill_2 FILLER_50_250 ();
 sg13g2_fill_1 FILLER_50_252 ();
 sg13g2_decap_4 FILLER_50_259 ();
 sg13g2_fill_1 FILLER_50_263 ();
 sg13g2_fill_2 FILLER_50_284 ();
 sg13g2_decap_8 FILLER_50_374 ();
 sg13g2_decap_8 FILLER_50_381 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_4 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_4 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_103 ();
 sg13g2_decap_8 FILLER_51_110 ();
 sg13g2_decap_8 FILLER_51_117 ();
 sg13g2_decap_4 FILLER_51_124 ();
 sg13g2_fill_2 FILLER_51_128 ();
 sg13g2_decap_4 FILLER_51_156 ();
 sg13g2_fill_1 FILLER_51_160 ();
 sg13g2_decap_8 FILLER_51_264 ();
 sg13g2_decap_8 FILLER_51_271 ();
 sg13g2_decap_8 FILLER_51_278 ();
 sg13g2_decap_4 FILLER_51_285 ();
 sg13g2_fill_2 FILLER_51_289 ();
 sg13g2_decap_4 FILLER_51_312 ();
 sg13g2_fill_1 FILLER_51_316 ();
 sg13g2_decap_8 FILLER_51_369 ();
 sg13g2_decap_8 FILLER_51_376 ();
 sg13g2_decap_8 FILLER_51_383 ();
 sg13g2_decap_8 FILLER_51_390 ();
 sg13g2_decap_8 FILLER_51_397 ();
 sg13g2_decap_4 FILLER_51_404 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_44 ();
 sg13g2_decap_8 FILLER_52_51 ();
 sg13g2_fill_1 FILLER_52_118 ();
 sg13g2_decap_8 FILLER_52_145 ();
 sg13g2_decap_8 FILLER_52_152 ();
 sg13g2_fill_2 FILLER_52_159 ();
 sg13g2_fill_1 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_170 ();
 sg13g2_decap_4 FILLER_52_177 ();
 sg13g2_fill_1 FILLER_52_181 ();
 sg13g2_fill_2 FILLER_52_270 ();
 sg13g2_decap_8 FILLER_52_280 ();
 sg13g2_decap_8 FILLER_52_291 ();
 sg13g2_decap_8 FILLER_52_298 ();
 sg13g2_decap_8 FILLER_52_305 ();
 sg13g2_decap_8 FILLER_52_312 ();
 sg13g2_fill_2 FILLER_52_319 ();
 sg13g2_decap_8 FILLER_52_331 ();
 sg13g2_decap_8 FILLER_52_338 ();
 sg13g2_decap_4 FILLER_52_345 ();
 sg13g2_fill_1 FILLER_52_349 ();
 sg13g2_decap_8 FILLER_52_354 ();
 sg13g2_decap_8 FILLER_52_361 ();
 sg13g2_decap_8 FILLER_52_368 ();
 sg13g2_decap_8 FILLER_52_375 ();
 sg13g2_decap_8 FILLER_52_382 ();
 sg13g2_decap_8 FILLER_52_389 ();
 sg13g2_decap_8 FILLER_52_396 ();
 sg13g2_decap_4 FILLER_52_403 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_21 ();
 sg13g2_fill_1 FILLER_53_23 ();
 sg13g2_decap_8 FILLER_53_128 ();
 sg13g2_fill_1 FILLER_53_135 ();
 sg13g2_decap_8 FILLER_53_162 ();
 sg13g2_decap_8 FILLER_53_169 ();
 sg13g2_decap_8 FILLER_53_176 ();
 sg13g2_fill_2 FILLER_53_183 ();
 sg13g2_decap_8 FILLER_53_211 ();
 sg13g2_decap_8 FILLER_53_218 ();
 sg13g2_fill_1 FILLER_53_225 ();
 sg13g2_fill_1 FILLER_53_270 ();
 sg13g2_decap_8 FILLER_53_299 ();
 sg13g2_decap_4 FILLER_53_306 ();
 sg13g2_fill_1 FILLER_53_310 ();
 sg13g2_decap_8 FILLER_53_316 ();
 sg13g2_decap_8 FILLER_53_323 ();
 sg13g2_decap_4 FILLER_53_330 ();
 sg13g2_fill_1 FILLER_53_334 ();
 sg13g2_fill_1 FILLER_53_351 ();
 sg13g2_decap_8 FILLER_53_368 ();
 sg13g2_decap_8 FILLER_53_375 ();
 sg13g2_decap_8 FILLER_53_382 ();
 sg13g2_decap_8 FILLER_53_389 ();
 sg13g2_decap_8 FILLER_53_396 ();
 sg13g2_decap_4 FILLER_53_403 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_4 FILLER_54_14 ();
 sg13g2_fill_1 FILLER_54_18 ();
 sg13g2_decap_4 FILLER_54_45 ();
 sg13g2_fill_1 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_55 ();
 sg13g2_fill_2 FILLER_54_62 ();
 sg13g2_decap_4 FILLER_54_168 ();
 sg13g2_fill_2 FILLER_54_172 ();
 sg13g2_decap_4 FILLER_54_182 ();
 sg13g2_fill_2 FILLER_54_186 ();
 sg13g2_decap_8 FILLER_54_218 ();
 sg13g2_decap_8 FILLER_54_225 ();
 sg13g2_fill_2 FILLER_54_232 ();
 sg13g2_fill_1 FILLER_54_234 ();
 sg13g2_decap_8 FILLER_54_241 ();
 sg13g2_decap_8 FILLER_54_248 ();
 sg13g2_decap_4 FILLER_54_261 ();
 sg13g2_fill_2 FILLER_54_328 ();
 sg13g2_fill_1 FILLER_54_330 ();
 sg13g2_decap_8 FILLER_54_371 ();
 sg13g2_decap_8 FILLER_54_378 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_399 ();
 sg13g2_fill_2 FILLER_54_406 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_4 ();
 sg13g2_decap_8 FILLER_55_75 ();
 sg13g2_decap_8 FILLER_55_82 ();
 sg13g2_decap_8 FILLER_55_89 ();
 sg13g2_decap_4 FILLER_55_96 ();
 sg13g2_fill_1 FILLER_55_100 ();
 sg13g2_decap_8 FILLER_55_106 ();
 sg13g2_decap_8 FILLER_55_191 ();
 sg13g2_decap_8 FILLER_55_198 ();
 sg13g2_decap_8 FILLER_55_205 ();
 sg13g2_decap_8 FILLER_55_212 ();
 sg13g2_fill_1 FILLER_55_219 ();
 sg13g2_decap_8 FILLER_55_230 ();
 sg13g2_fill_1 FILLER_55_237 ();
 sg13g2_decap_8 FILLER_55_243 ();
 sg13g2_decap_8 FILLER_55_250 ();
 sg13g2_decap_8 FILLER_55_257 ();
 sg13g2_decap_8 FILLER_55_264 ();
 sg13g2_fill_1 FILLER_55_271 ();
 sg13g2_fill_2 FILLER_55_297 ();
 sg13g2_decap_8 FILLER_55_333 ();
 sg13g2_fill_2 FILLER_55_348 ();
 sg13g2_decap_8 FILLER_55_374 ();
 sg13g2_decap_8 FILLER_55_381 ();
 sg13g2_decap_8 FILLER_55_388 ();
 sg13g2_decap_8 FILLER_55_395 ();
 sg13g2_decap_8 FILLER_55_402 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_4 FILLER_56_28 ();
 sg13g2_fill_2 FILLER_56_32 ();
 sg13g2_decap_8 FILLER_56_60 ();
 sg13g2_decap_8 FILLER_56_67 ();
 sg13g2_decap_8 FILLER_56_74 ();
 sg13g2_decap_8 FILLER_56_81 ();
 sg13g2_decap_8 FILLER_56_88 ();
 sg13g2_decap_8 FILLER_56_95 ();
 sg13g2_fill_1 FILLER_56_102 ();
 sg13g2_decap_8 FILLER_56_129 ();
 sg13g2_decap_8 FILLER_56_136 ();
 sg13g2_decap_8 FILLER_56_143 ();
 sg13g2_decap_4 FILLER_56_150 ();
 sg13g2_fill_2 FILLER_56_154 ();
 sg13g2_decap_4 FILLER_56_208 ();
 sg13g2_fill_2 FILLER_56_212 ();
 sg13g2_fill_1 FILLER_56_240 ();
 sg13g2_fill_2 FILLER_56_246 ();
 sg13g2_decap_8 FILLER_56_258 ();
 sg13g2_decap_8 FILLER_56_265 ();
 sg13g2_decap_4 FILLER_56_272 ();
 sg13g2_fill_2 FILLER_56_280 ();
 sg13g2_fill_1 FILLER_56_282 ();
 sg13g2_decap_8 FILLER_56_292 ();
 sg13g2_decap_4 FILLER_56_299 ();
 sg13g2_decap_8 FILLER_56_333 ();
 sg13g2_fill_2 FILLER_56_340 ();
 sg13g2_decap_8 FILLER_56_370 ();
 sg13g2_decap_8 FILLER_56_377 ();
 sg13g2_decap_8 FILLER_56_384 ();
 sg13g2_decap_8 FILLER_56_391 ();
 sg13g2_decap_8 FILLER_56_398 ();
 sg13g2_decap_4 FILLER_56_405 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_fill_2 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_16 ();
 sg13g2_decap_8 FILLER_57_47 ();
 sg13g2_fill_2 FILLER_57_54 ();
 sg13g2_fill_1 FILLER_57_56 ();
 sg13g2_fill_1 FILLER_57_83 ();
 sg13g2_decap_8 FILLER_57_110 ();
 sg13g2_decap_8 FILLER_57_117 ();
 sg13g2_decap_8 FILLER_57_124 ();
 sg13g2_decap_8 FILLER_57_131 ();
 sg13g2_decap_8 FILLER_57_138 ();
 sg13g2_decap_8 FILLER_57_145 ();
 sg13g2_decap_8 FILLER_57_152 ();
 sg13g2_decap_8 FILLER_57_163 ();
 sg13g2_decap_8 FILLER_57_170 ();
 sg13g2_decap_4 FILLER_57_177 ();
 sg13g2_fill_2 FILLER_57_181 ();
 sg13g2_fill_2 FILLER_57_209 ();
 sg13g2_fill_1 FILLER_57_211 ();
 sg13g2_fill_2 FILLER_57_238 ();
 sg13g2_fill_1 FILLER_57_240 ();
 sg13g2_fill_2 FILLER_57_280 ();
 sg13g2_fill_1 FILLER_57_293 ();
 sg13g2_decap_8 FILLER_57_302 ();
 sg13g2_decap_8 FILLER_57_309 ();
 sg13g2_decap_8 FILLER_57_316 ();
 sg13g2_decap_4 FILLER_57_323 ();
 sg13g2_fill_2 FILLER_57_347 ();
 sg13g2_fill_1 FILLER_57_349 ();
 sg13g2_decap_8 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_385 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_fill_2 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_4 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_110 ();
 sg13g2_fill_1 FILLER_58_117 ();
 sg13g2_fill_2 FILLER_58_144 ();
 sg13g2_fill_2 FILLER_58_172 ();
 sg13g2_fill_1 FILLER_58_174 ();
 sg13g2_fill_2 FILLER_58_180 ();
 sg13g2_fill_1 FILLER_58_182 ();
 sg13g2_fill_2 FILLER_58_209 ();
 sg13g2_fill_2 FILLER_58_237 ();
 sg13g2_fill_1 FILLER_58_239 ();
 sg13g2_decap_4 FILLER_58_272 ();
 sg13g2_fill_1 FILLER_58_286 ();
 sg13g2_fill_2 FILLER_58_297 ();
 sg13g2_decap_8 FILLER_58_325 ();
 sg13g2_fill_2 FILLER_58_352 ();
 sg13g2_decap_8 FILLER_58_374 ();
 sg13g2_decap_8 FILLER_58_381 ();
 sg13g2_decap_8 FILLER_58_388 ();
 sg13g2_decap_8 FILLER_58_395 ();
 sg13g2_decap_8 FILLER_58_402 ();
 sg13g2_decap_8 FILLER_59_26 ();
 sg13g2_decap_4 FILLER_59_33 ();
 sg13g2_fill_1 FILLER_59_37 ();
 sg13g2_decap_4 FILLER_59_64 ();
 sg13g2_fill_2 FILLER_59_102 ();
 sg13g2_fill_2 FILLER_59_139 ();
 sg13g2_fill_1 FILLER_59_141 ();
 sg13g2_fill_2 FILLER_59_147 ();
 sg13g2_fill_1 FILLER_59_167 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_decap_4 FILLER_59_210 ();
 sg13g2_fill_2 FILLER_59_214 ();
 sg13g2_fill_2 FILLER_59_224 ();
 sg13g2_fill_2 FILLER_59_246 ();
 sg13g2_fill_1 FILLER_59_248 ();
 sg13g2_fill_1 FILLER_59_259 ();
 sg13g2_decap_4 FILLER_59_348 ();
 sg13g2_decap_8 FILLER_59_356 ();
 sg13g2_decap_8 FILLER_59_363 ();
 sg13g2_decap_8 FILLER_59_370 ();
 sg13g2_decap_8 FILLER_59_377 ();
 sg13g2_decap_8 FILLER_59_384 ();
 sg13g2_decap_8 FILLER_59_391 ();
 sg13g2_decap_8 FILLER_59_398 ();
 sg13g2_decap_4 FILLER_59_405 ();
 sg13g2_decap_8 FILLER_60_26 ();
 sg13g2_fill_2 FILLER_60_33 ();
 sg13g2_decap_8 FILLER_60_61 ();
 sg13g2_decap_8 FILLER_60_68 ();
 sg13g2_decap_8 FILLER_60_75 ();
 sg13g2_fill_1 FILLER_60_82 ();
 sg13g2_decap_4 FILLER_60_109 ();
 sg13g2_fill_2 FILLER_60_113 ();
 sg13g2_fill_2 FILLER_60_163 ();
 sg13g2_decap_8 FILLER_60_191 ();
 sg13g2_decap_8 FILLER_60_198 ();
 sg13g2_fill_1 FILLER_60_205 ();
 sg13g2_decap_8 FILLER_60_214 ();
 sg13g2_decap_8 FILLER_60_221 ();
 sg13g2_fill_2 FILLER_60_249 ();
 sg13g2_fill_1 FILLER_60_251 ();
 sg13g2_fill_2 FILLER_60_263 ();
 sg13g2_decap_8 FILLER_60_331 ();
 sg13g2_decap_4 FILLER_60_338 ();
 sg13g2_fill_1 FILLER_60_367 ();
 sg13g2_decap_8 FILLER_60_381 ();
 sg13g2_decap_8 FILLER_60_388 ();
 sg13g2_decap_8 FILLER_60_395 ();
 sg13g2_decap_8 FILLER_60_402 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_decap_8 FILLER_61_107 ();
 sg13g2_fill_2 FILLER_61_114 ();
 sg13g2_fill_1 FILLER_61_185 ();
 sg13g2_decap_8 FILLER_61_212 ();
 sg13g2_fill_2 FILLER_61_245 ();
 sg13g2_decap_4 FILLER_61_278 ();
 sg13g2_fill_2 FILLER_61_282 ();
 sg13g2_fill_1 FILLER_61_293 ();
 sg13g2_decap_8 FILLER_61_304 ();
 sg13g2_decap_8 FILLER_61_311 ();
 sg13g2_decap_8 FILLER_61_318 ();
 sg13g2_decap_8 FILLER_61_325 ();
 sg13g2_decap_8 FILLER_61_391 ();
 sg13g2_decap_8 FILLER_61_398 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_11 ();
 sg13g2_decap_8 FILLER_62_65 ();
 sg13g2_decap_8 FILLER_62_72 ();
 sg13g2_decap_4 FILLER_62_79 ();
 sg13g2_decap_8 FILLER_62_109 ();
 sg13g2_fill_2 FILLER_62_147 ();
 sg13g2_fill_2 FILLER_62_168 ();
 sg13g2_fill_1 FILLER_62_183 ();
 sg13g2_decap_4 FILLER_62_214 ();
 sg13g2_decap_8 FILLER_62_270 ();
 sg13g2_decap_8 FILLER_62_277 ();
 sg13g2_decap_4 FILLER_62_284 ();
 sg13g2_decap_4 FILLER_62_294 ();
 sg13g2_fill_1 FILLER_62_298 ();
 sg13g2_fill_2 FILLER_62_305 ();
 sg13g2_fill_1 FILLER_62_349 ();
 sg13g2_decap_8 FILLER_62_384 ();
 sg13g2_decap_8 FILLER_62_391 ();
 sg13g2_decap_8 FILLER_62_398 ();
 sg13g2_decap_4 FILLER_62_405 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_41 ();
 sg13g2_decap_8 FILLER_63_48 ();
 sg13g2_decap_8 FILLER_63_55 ();
 sg13g2_fill_2 FILLER_63_62 ();
 sg13g2_fill_1 FILLER_63_64 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_4 FILLER_63_105 ();
 sg13g2_fill_2 FILLER_63_109 ();
 sg13g2_decap_4 FILLER_63_123 ();
 sg13g2_fill_2 FILLER_63_127 ();
 sg13g2_decap_8 FILLER_63_137 ();
 sg13g2_decap_8 FILLER_63_144 ();
 sg13g2_fill_1 FILLER_63_151 ();
 sg13g2_decap_4 FILLER_63_157 ();
 sg13g2_fill_1 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_165 ();
 sg13g2_fill_2 FILLER_63_196 ();
 sg13g2_decap_4 FILLER_63_224 ();
 sg13g2_fill_1 FILLER_63_228 ();
 sg13g2_fill_2 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_267 ();
 sg13g2_fill_1 FILLER_63_274 ();
 sg13g2_decap_4 FILLER_63_326 ();
 sg13g2_fill_1 FILLER_63_330 ();
 sg13g2_fill_1 FILLER_63_351 ();
 sg13g2_decap_4 FILLER_63_360 ();
 sg13g2_decap_8 FILLER_63_377 ();
 sg13g2_decap_8 FILLER_63_384 ();
 sg13g2_decap_8 FILLER_63_391 ();
 sg13g2_decap_8 FILLER_63_398 ();
 sg13g2_decap_4 FILLER_63_405 ();
 sg13g2_decap_8 FILLER_64_86 ();
 sg13g2_decap_8 FILLER_64_93 ();
 sg13g2_fill_2 FILLER_64_100 ();
 sg13g2_fill_1 FILLER_64_102 ();
 sg13g2_decap_4 FILLER_64_129 ();
 sg13g2_fill_2 FILLER_64_141 ();
 sg13g2_fill_1 FILLER_64_143 ();
 sg13g2_decap_4 FILLER_64_148 ();
 sg13g2_fill_1 FILLER_64_152 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_fill_2 FILLER_64_168 ();
 sg13g2_fill_1 FILLER_64_170 ();
 sg13g2_fill_1 FILLER_64_176 ();
 sg13g2_decap_8 FILLER_64_185 ();
 sg13g2_decap_4 FILLER_64_192 ();
 sg13g2_fill_1 FILLER_64_196 ();
 sg13g2_decap_8 FILLER_64_223 ();
 sg13g2_decap_8 FILLER_64_230 ();
 sg13g2_decap_8 FILLER_64_237 ();
 sg13g2_decap_8 FILLER_64_244 ();
 sg13g2_decap_4 FILLER_64_251 ();
 sg13g2_fill_1 FILLER_64_255 ();
 sg13g2_fill_2 FILLER_64_282 ();
 sg13g2_fill_1 FILLER_64_284 ();
 sg13g2_decap_8 FILLER_64_289 ();
 sg13g2_decap_4 FILLER_64_296 ();
 sg13g2_decap_4 FILLER_64_309 ();
 sg13g2_fill_1 FILLER_64_313 ();
 sg13g2_decap_8 FILLER_64_321 ();
 sg13g2_decap_8 FILLER_64_328 ();
 sg13g2_decap_8 FILLER_64_335 ();
 sg13g2_decap_8 FILLER_64_350 ();
 sg13g2_decap_4 FILLER_64_357 ();
 sg13g2_decap_8 FILLER_64_372 ();
 sg13g2_decap_4 FILLER_64_379 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_14 ();
 sg13g2_fill_1 FILLER_65_16 ();
 sg13g2_fill_1 FILLER_65_74 ();
 sg13g2_decap_4 FILLER_65_101 ();
 sg13g2_fill_2 FILLER_65_127 ();
 sg13g2_fill_1 FILLER_65_129 ();
 sg13g2_fill_1 FILLER_65_139 ();
 sg13g2_fill_2 FILLER_65_155 ();
 sg13g2_fill_1 FILLER_65_157 ();
 sg13g2_decap_4 FILLER_65_202 ();
 sg13g2_fill_2 FILLER_65_206 ();
 sg13g2_fill_2 FILLER_65_216 ();
 sg13g2_decap_8 FILLER_65_226 ();
 sg13g2_decap_8 FILLER_65_233 ();
 sg13g2_decap_8 FILLER_65_240 ();
 sg13g2_decap_8 FILLER_65_247 ();
 sg13g2_decap_4 FILLER_65_254 ();
 sg13g2_fill_1 FILLER_65_258 ();
 sg13g2_fill_1 FILLER_65_290 ();
 sg13g2_decap_8 FILLER_65_323 ();
 sg13g2_decap_8 FILLER_65_330 ();
 sg13g2_decap_8 FILLER_65_337 ();
 sg13g2_fill_2 FILLER_65_344 ();
 sg13g2_fill_2 FILLER_65_364 ();
 sg13g2_fill_1 FILLER_65_366 ();
 sg13g2_fill_1 FILLER_65_393 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_fill_2 FILLER_66_26 ();
 sg13g2_fill_1 FILLER_66_28 ();
 sg13g2_fill_2 FILLER_66_63 ();
 sg13g2_decap_4 FILLER_66_99 ();
 sg13g2_fill_2 FILLER_66_122 ();
 sg13g2_fill_2 FILLER_66_197 ();
 sg13g2_fill_2 FILLER_66_225 ();
 sg13g2_decap_4 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_241 ();
 sg13g2_fill_2 FILLER_66_252 ();
 sg13g2_decap_4 FILLER_66_268 ();
 sg13g2_decap_8 FILLER_66_280 ();
 sg13g2_decap_8 FILLER_66_323 ();
 sg13g2_fill_2 FILLER_66_330 ();
 sg13g2_fill_1 FILLER_66_332 ();
 sg13g2_fill_2 FILLER_66_359 ();
 sg13g2_decap_4 FILLER_67_26 ();
 sg13g2_fill_2 FILLER_67_30 ();
 sg13g2_decap_8 FILLER_67_37 ();
 sg13g2_decap_8 FILLER_67_44 ();
 sg13g2_decap_8 FILLER_67_51 ();
 sg13g2_decap_4 FILLER_67_58 ();
 sg13g2_fill_1 FILLER_67_62 ();
 sg13g2_decap_4 FILLER_67_94 ();
 sg13g2_fill_1 FILLER_67_98 ();
 sg13g2_fill_2 FILLER_67_143 ();
 sg13g2_fill_1 FILLER_67_150 ();
 sg13g2_fill_2 FILLER_67_156 ();
 sg13g2_fill_2 FILLER_67_172 ();
 sg13g2_decap_4 FILLER_67_183 ();
 sg13g2_fill_2 FILLER_67_229 ();
 sg13g2_fill_1 FILLER_67_257 ();
 sg13g2_fill_2 FILLER_67_302 ();
 sg13g2_decap_4 FILLER_67_314 ();
 sg13g2_fill_2 FILLER_67_318 ();
 sg13g2_fill_2 FILLER_67_351 ();
 sg13g2_fill_1 FILLER_67_353 ();
 sg13g2_fill_1 FILLER_67_365 ();
 sg13g2_fill_2 FILLER_67_382 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_4 FILLER_68_28 ();
 sg13g2_fill_2 FILLER_68_32 ();
 sg13g2_decap_8 FILLER_68_86 ();
 sg13g2_decap_8 FILLER_68_93 ();
 sg13g2_decap_4 FILLER_68_100 ();
 sg13g2_fill_2 FILLER_68_104 ();
 sg13g2_fill_1 FILLER_68_115 ();
 sg13g2_fill_2 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_139 ();
 sg13g2_decap_8 FILLER_68_146 ();
 sg13g2_decap_8 FILLER_68_153 ();
 sg13g2_decap_4 FILLER_68_160 ();
 sg13g2_decap_8 FILLER_68_171 ();
 sg13g2_decap_4 FILLER_68_178 ();
 sg13g2_fill_1 FILLER_68_182 ();
 sg13g2_fill_1 FILLER_68_195 ();
 sg13g2_fill_1 FILLER_68_200 ();
 sg13g2_decap_4 FILLER_68_227 ();
 sg13g2_fill_2 FILLER_68_231 ();
 sg13g2_fill_2 FILLER_68_264 ();
 sg13g2_decap_8 FILLER_68_296 ();
 sg13g2_decap_8 FILLER_68_303 ();
 sg13g2_decap_4 FILLER_68_310 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_fill_1 FILLER_68_324 ();
 sg13g2_fill_2 FILLER_68_371 ();
 sg13g2_fill_1 FILLER_68_373 ();
 sg13g2_decap_8 FILLER_68_384 ();
 sg13g2_fill_2 FILLER_68_391 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_4 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_65 ();
 sg13g2_decap_8 FILLER_69_72 ();
 sg13g2_decap_8 FILLER_69_79 ();
 sg13g2_decap_8 FILLER_69_86 ();
 sg13g2_decap_8 FILLER_69_93 ();
 sg13g2_decap_8 FILLER_69_100 ();
 sg13g2_decap_4 FILLER_69_107 ();
 sg13g2_fill_2 FILLER_69_111 ();
 sg13g2_fill_2 FILLER_69_118 ();
 sg13g2_fill_1 FILLER_69_120 ();
 sg13g2_fill_2 FILLER_69_125 ();
 sg13g2_decap_8 FILLER_69_131 ();
 sg13g2_decap_4 FILLER_69_138 ();
 sg13g2_fill_1 FILLER_69_142 ();
 sg13g2_decap_4 FILLER_69_147 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_fill_1 FILLER_69_160 ();
 sg13g2_fill_1 FILLER_69_170 ();
 sg13g2_fill_1 FILLER_69_176 ();
 sg13g2_decap_4 FILLER_69_181 ();
 sg13g2_decap_8 FILLER_69_202 ();
 sg13g2_decap_8 FILLER_69_209 ();
 sg13g2_decap_8 FILLER_69_216 ();
 sg13g2_decap_8 FILLER_69_223 ();
 sg13g2_fill_1 FILLER_69_230 ();
 sg13g2_fill_1 FILLER_69_246 ();
 sg13g2_decap_8 FILLER_69_283 ();
 sg13g2_fill_2 FILLER_69_290 ();
 sg13g2_fill_1 FILLER_69_292 ();
 sg13g2_decap_8 FILLER_69_298 ();
 sg13g2_decap_8 FILLER_69_310 ();
 sg13g2_decap_8 FILLER_69_317 ();
 sg13g2_decap_4 FILLER_69_328 ();
 sg13g2_fill_2 FILLER_69_332 ();
 sg13g2_fill_2 FILLER_69_339 ();
 sg13g2_fill_1 FILLER_69_341 ();
 sg13g2_decap_4 FILLER_69_361 ();
 sg13g2_decap_4 FILLER_69_370 ();
 sg13g2_fill_2 FILLER_69_374 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_47 ();
 sg13g2_decap_8 FILLER_70_54 ();
 sg13g2_decap_8 FILLER_70_61 ();
 sg13g2_decap_8 FILLER_70_68 ();
 sg13g2_fill_1 FILLER_70_135 ();
 sg13g2_decap_8 FILLER_70_208 ();
 sg13g2_decap_8 FILLER_70_215 ();
 sg13g2_fill_1 FILLER_70_222 ();
 sg13g2_decap_8 FILLER_70_231 ();
 sg13g2_decap_8 FILLER_70_246 ();
 sg13g2_decap_8 FILLER_70_253 ();
 sg13g2_fill_2 FILLER_70_260 ();
 sg13g2_decap_8 FILLER_70_272 ();
 sg13g2_fill_1 FILLER_70_279 ();
 sg13g2_decap_8 FILLER_70_290 ();
 sg13g2_decap_4 FILLER_70_297 ();
 sg13g2_fill_1 FILLER_70_301 ();
 sg13g2_fill_2 FILLER_70_307 ();
 sg13g2_fill_1 FILLER_70_309 ();
 sg13g2_fill_2 FILLER_70_315 ();
 sg13g2_fill_1 FILLER_70_317 ();
 sg13g2_fill_2 FILLER_70_348 ();
 sg13g2_decap_8 FILLER_70_360 ();
 sg13g2_fill_1 FILLER_70_367 ();
 sg13g2_fill_1 FILLER_70_382 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_fill_1 FILLER_71_21 ();
 sg13g2_fill_1 FILLER_71_131 ();
 sg13g2_fill_1 FILLER_71_202 ();
 sg13g2_decap_8 FILLER_71_237 ();
 sg13g2_fill_2 FILLER_71_254 ();
 sg13g2_fill_1 FILLER_71_256 ();
 sg13g2_decap_8 FILLER_71_265 ();
 sg13g2_fill_2 FILLER_71_272 ();
 sg13g2_fill_2 FILLER_71_284 ();
 sg13g2_fill_1 FILLER_71_286 ();
 sg13g2_decap_8 FILLER_71_339 ();
 sg13g2_fill_1 FILLER_71_356 ();
 sg13g2_fill_2 FILLER_71_372 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_4 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_fill_2 FILLER_72_77 ();
 sg13g2_fill_2 FILLER_72_153 ();
 sg13g2_fill_1 FILLER_72_155 ();
 sg13g2_fill_1 FILLER_72_176 ();
 sg13g2_decap_8 FILLER_72_182 ();
 sg13g2_decap_4 FILLER_72_189 ();
 sg13g2_fill_1 FILLER_72_193 ();
 sg13g2_decap_4 FILLER_72_242 ();
 sg13g2_decap_4 FILLER_72_308 ();
 sg13g2_fill_1 FILLER_72_312 ();
 sg13g2_decap_8 FILLER_72_328 ();
 sg13g2_decap_8 FILLER_72_335 ();
 sg13g2_decap_4 FILLER_72_342 ();
 sg13g2_fill_2 FILLER_72_346 ();
 sg13g2_fill_1 FILLER_72_360 ();
 sg13g2_decap_4 FILLER_72_381 ();
 sg13g2_fill_2 FILLER_72_385 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_fill_1 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_48 ();
 sg13g2_decap_8 FILLER_73_55 ();
 sg13g2_fill_1 FILLER_73_62 ();
 sg13g2_decap_4 FILLER_73_71 ();
 sg13g2_fill_1 FILLER_73_75 ();
 sg13g2_decap_8 FILLER_73_102 ();
 sg13g2_fill_1 FILLER_73_109 ();
 sg13g2_fill_2 FILLER_73_122 ();
 sg13g2_fill_1 FILLER_73_124 ();
 sg13g2_decap_4 FILLER_73_153 ();
 sg13g2_fill_2 FILLER_73_157 ();
 sg13g2_decap_4 FILLER_73_176 ();
 sg13g2_fill_1 FILLER_73_180 ();
 sg13g2_decap_8 FILLER_73_186 ();
 sg13g2_decap_8 FILLER_73_198 ();
 sg13g2_decap_4 FILLER_73_205 ();
 sg13g2_fill_2 FILLER_73_209 ();
 sg13g2_fill_2 FILLER_73_219 ();
 sg13g2_fill_1 FILLER_73_284 ();
 sg13g2_decap_4 FILLER_73_311 ();
 sg13g2_fill_2 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_363 ();
 sg13g2_fill_2 FILLER_73_382 ();
 sg13g2_fill_2 FILLER_73_388 ();
 sg13g2_decap_8 FILLER_73_395 ();
 sg13g2_decap_8 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_fill_1 FILLER_74_21 ();
 sg13g2_decap_4 FILLER_74_48 ();
 sg13g2_fill_1 FILLER_74_78 ();
 sg13g2_fill_1 FILLER_74_83 ();
 sg13g2_decap_8 FILLER_74_92 ();
 sg13g2_decap_8 FILLER_74_99 ();
 sg13g2_decap_8 FILLER_74_106 ();
 sg13g2_decap_8 FILLER_74_113 ();
 sg13g2_fill_1 FILLER_74_120 ();
 sg13g2_fill_1 FILLER_74_126 ();
 sg13g2_decap_4 FILLER_74_131 ();
 sg13g2_fill_2 FILLER_74_135 ();
 sg13g2_decap_8 FILLER_74_146 ();
 sg13g2_decap_8 FILLER_74_153 ();
 sg13g2_decap_8 FILLER_74_160 ();
 sg13g2_decap_8 FILLER_74_167 ();
 sg13g2_decap_8 FILLER_74_174 ();
 sg13g2_decap_4 FILLER_74_181 ();
 sg13g2_fill_1 FILLER_74_185 ();
 sg13g2_decap_8 FILLER_74_212 ();
 sg13g2_decap_8 FILLER_74_229 ();
 sg13g2_decap_4 FILLER_74_236 ();
 sg13g2_fill_1 FILLER_74_240 ();
 sg13g2_decap_8 FILLER_74_253 ();
 sg13g2_decap_8 FILLER_74_260 ();
 sg13g2_decap_4 FILLER_74_267 ();
 sg13g2_fill_1 FILLER_74_271 ();
 sg13g2_decap_8 FILLER_74_282 ();
 sg13g2_fill_2 FILLER_74_289 ();
 sg13g2_fill_1 FILLER_74_291 ();
 sg13g2_fill_2 FILLER_74_296 ();
 sg13g2_decap_8 FILLER_74_306 ();
 sg13g2_fill_2 FILLER_74_313 ();
 sg13g2_fill_1 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_324 ();
 sg13g2_fill_1 FILLER_74_331 ();
 sg13g2_decap_4 FILLER_74_362 ();
 sg13g2_fill_2 FILLER_74_366 ();
 sg13g2_fill_1 FILLER_74_373 ();
 sg13g2_decap_8 FILLER_74_395 ();
 sg13g2_decap_8 FILLER_74_402 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_fill_1 FILLER_75_78 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_fill_2 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_163 ();
 sg13g2_decap_4 FILLER_75_170 ();
 sg13g2_fill_2 FILLER_75_174 ();
 sg13g2_decap_8 FILLER_75_184 ();
 sg13g2_decap_4 FILLER_75_191 ();
 sg13g2_fill_2 FILLER_75_195 ();
 sg13g2_decap_8 FILLER_75_204 ();
 sg13g2_decap_8 FILLER_75_211 ();
 sg13g2_decap_4 FILLER_75_218 ();
 sg13g2_fill_1 FILLER_75_222 ();
 sg13g2_decap_4 FILLER_75_233 ();
 sg13g2_fill_2 FILLER_75_237 ();
 sg13g2_decap_8 FILLER_75_261 ();
 sg13g2_decap_4 FILLER_75_268 ();
 sg13g2_fill_2 FILLER_75_272 ();
 sg13g2_decap_4 FILLER_75_309 ();
 sg13g2_fill_2 FILLER_75_313 ();
 sg13g2_decap_4 FILLER_75_320 ();
 sg13g2_decap_4 FILLER_75_329 ();
 sg13g2_fill_2 FILLER_75_333 ();
 sg13g2_fill_1 FILLER_75_340 ();
 sg13g2_decap_4 FILLER_75_357 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_decap_4 FILLER_75_404 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_fill_2 FILLER_76_63 ();
 sg13g2_fill_1 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_76 ();
 sg13g2_decap_8 FILLER_76_83 ();
 sg13g2_decap_4 FILLER_76_121 ();
 sg13g2_fill_1 FILLER_76_125 ();
 sg13g2_fill_1 FILLER_76_187 ();
 sg13g2_fill_2 FILLER_76_214 ();
 sg13g2_fill_1 FILLER_76_216 ();
 sg13g2_fill_1 FILLER_76_237 ();
 sg13g2_fill_2 FILLER_76_269 ();
 sg13g2_decap_4 FILLER_76_281 ();
 sg13g2_decap_8 FILLER_76_334 ();
 sg13g2_fill_1 FILLER_76_341 ();
 sg13g2_fill_2 FILLER_76_352 ();
 sg13g2_fill_2 FILLER_76_363 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_4 FILLER_77_42 ();
 sg13g2_fill_2 FILLER_77_46 ();
 sg13g2_fill_2 FILLER_77_105 ();
 sg13g2_fill_1 FILLER_77_107 ();
 sg13g2_decap_8 FILLER_77_134 ();
 sg13g2_decap_8 FILLER_77_141 ();
 sg13g2_decap_4 FILLER_77_148 ();
 sg13g2_fill_2 FILLER_77_157 ();
 sg13g2_fill_2 FILLER_77_206 ();
 sg13g2_fill_2 FILLER_77_239 ();
 sg13g2_fill_1 FILLER_77_241 ();
 sg13g2_fill_2 FILLER_77_304 ();
 sg13g2_fill_1 FILLER_77_332 ();
 sg13g2_fill_1 FILLER_77_347 ();
 sg13g2_fill_1 FILLER_77_380 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_fill_1 FILLER_78_73 ();
 sg13g2_decap_4 FILLER_78_152 ();
 sg13g2_fill_2 FILLER_78_156 ();
 sg13g2_decap_8 FILLER_78_236 ();
 sg13g2_fill_1 FILLER_78_243 ();
 sg13g2_decap_4 FILLER_78_270 ();
 sg13g2_fill_2 FILLER_78_300 ();
 sg13g2_fill_1 FILLER_78_302 ();
 sg13g2_fill_1 FILLER_78_381 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_4 FILLER_79_65 ();
 sg13g2_fill_1 FILLER_79_69 ();
 sg13g2_decap_8 FILLER_79_122 ();
 sg13g2_decap_8 FILLER_79_129 ();
 sg13g2_decap_4 FILLER_79_136 ();
 sg13g2_fill_2 FILLER_79_174 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_4 FILLER_79_252 ();
 sg13g2_fill_1 FILLER_79_266 ();
 sg13g2_fill_2 FILLER_79_277 ();
 sg13g2_decap_4 FILLER_79_305 ();
 sg13g2_fill_1 FILLER_79_309 ();
 sg13g2_decap_8 FILLER_79_320 ();
 sg13g2_fill_1 FILLER_79_327 ();
 sg13g2_decap_4 FILLER_79_354 ();
 sg13g2_fill_2 FILLER_79_358 ();
 sg13g2_fill_1 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_389 ();
 sg13g2_decap_8 FILLER_79_396 ();
 sg13g2_decap_4 FILLER_79_403 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_8 FILLER_80_166 ();
 sg13g2_decap_8 FILLER_80_173 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_188 ();
 sg13g2_fill_1 FILLER_80_192 ();
 sg13g2_decap_4 FILLER_80_208 ();
 sg13g2_fill_2 FILLER_80_212 ();
 sg13g2_decap_8 FILLER_80_219 ();
 sg13g2_decap_8 FILLER_80_226 ();
 sg13g2_decap_8 FILLER_80_233 ();
 sg13g2_decap_8 FILLER_80_240 ();
 sg13g2_decap_8 FILLER_80_247 ();
 sg13g2_decap_8 FILLER_80_254 ();
 sg13g2_decap_8 FILLER_80_261 ();
 sg13g2_decap_4 FILLER_80_268 ();
 sg13g2_fill_1 FILLER_80_272 ();
 sg13g2_decap_8 FILLER_80_283 ();
 sg13g2_decap_8 FILLER_80_290 ();
 sg13g2_decap_8 FILLER_80_297 ();
 sg13g2_decap_8 FILLER_80_304 ();
 sg13g2_decap_8 FILLER_80_311 ();
 sg13g2_decap_4 FILLER_80_318 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_decap_4 FILLER_80_348 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_decap_8 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_371 ();
 sg13g2_decap_8 FILLER_80_378 ();
 sg13g2_decap_8 FILLER_80_385 ();
 sg13g2_decap_8 FILLER_80_392 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net40;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule

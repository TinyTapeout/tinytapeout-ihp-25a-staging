module tt_um_tiny_ternary_tapeout_csa (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire \bit_select[0] ;
 wire \bit_select[1] ;
 wire \bit_select[2] ;
 wire \bit_select[3] ;
 wire \bit_select[4] ;
 wire \bit_select[5] ;
 wire \bit_select[6] ;
 wire \bit_select[7] ;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \count[4] ;
 wire \count[5] ;
 wire \count[6] ;
 wire \count[7] ;
 wire load_ena;
 wire \load_weights[0] ;
 wire \load_weights[100] ;
 wire \load_weights[101] ;
 wire \load_weights[102] ;
 wire \load_weights[103] ;
 wire \load_weights[104] ;
 wire \load_weights[105] ;
 wire \load_weights[106] ;
 wire \load_weights[107] ;
 wire \load_weights[108] ;
 wire \load_weights[109] ;
 wire \load_weights[10] ;
 wire \load_weights[110] ;
 wire \load_weights[111] ;
 wire \load_weights[112] ;
 wire \load_weights[113] ;
 wire \load_weights[114] ;
 wire \load_weights[115] ;
 wire \load_weights[116] ;
 wire \load_weights[117] ;
 wire \load_weights[118] ;
 wire \load_weights[119] ;
 wire \load_weights[11] ;
 wire \load_weights[120] ;
 wire \load_weights[121] ;
 wire \load_weights[122] ;
 wire \load_weights[123] ;
 wire \load_weights[124] ;
 wire \load_weights[125] ;
 wire \load_weights[126] ;
 wire \load_weights[127] ;
 wire \load_weights[128] ;
 wire \load_weights[129] ;
 wire \load_weights[12] ;
 wire \load_weights[130] ;
 wire \load_weights[131] ;
 wire \load_weights[132] ;
 wire \load_weights[133] ;
 wire \load_weights[134] ;
 wire \load_weights[135] ;
 wire \load_weights[136] ;
 wire \load_weights[137] ;
 wire \load_weights[138] ;
 wire \load_weights[139] ;
 wire \load_weights[13] ;
 wire \load_weights[140] ;
 wire \load_weights[141] ;
 wire \load_weights[142] ;
 wire \load_weights[143] ;
 wire \load_weights[144] ;
 wire \load_weights[145] ;
 wire \load_weights[146] ;
 wire \load_weights[147] ;
 wire \load_weights[148] ;
 wire \load_weights[149] ;
 wire \load_weights[14] ;
 wire \load_weights[150] ;
 wire \load_weights[151] ;
 wire \load_weights[152] ;
 wire \load_weights[153] ;
 wire \load_weights[154] ;
 wire \load_weights[155] ;
 wire \load_weights[156] ;
 wire \load_weights[157] ;
 wire \load_weights[158] ;
 wire \load_weights[159] ;
 wire \load_weights[15] ;
 wire \load_weights[160] ;
 wire \load_weights[161] ;
 wire \load_weights[162] ;
 wire \load_weights[163] ;
 wire \load_weights[164] ;
 wire \load_weights[165] ;
 wire \load_weights[166] ;
 wire \load_weights[167] ;
 wire \load_weights[168] ;
 wire \load_weights[169] ;
 wire \load_weights[16] ;
 wire \load_weights[170] ;
 wire \load_weights[171] ;
 wire \load_weights[172] ;
 wire \load_weights[173] ;
 wire \load_weights[174] ;
 wire \load_weights[175] ;
 wire \load_weights[176] ;
 wire \load_weights[177] ;
 wire \load_weights[178] ;
 wire \load_weights[179] ;
 wire \load_weights[17] ;
 wire \load_weights[180] ;
 wire \load_weights[181] ;
 wire \load_weights[182] ;
 wire \load_weights[183] ;
 wire \load_weights[184] ;
 wire \load_weights[185] ;
 wire \load_weights[186] ;
 wire \load_weights[187] ;
 wire \load_weights[188] ;
 wire \load_weights[189] ;
 wire \load_weights[18] ;
 wire \load_weights[190] ;
 wire \load_weights[191] ;
 wire \load_weights[192] ;
 wire \load_weights[193] ;
 wire \load_weights[194] ;
 wire \load_weights[195] ;
 wire \load_weights[196] ;
 wire \load_weights[197] ;
 wire \load_weights[198] ;
 wire \load_weights[199] ;
 wire \load_weights[19] ;
 wire \load_weights[1] ;
 wire \load_weights[200] ;
 wire \load_weights[201] ;
 wire \load_weights[202] ;
 wire \load_weights[203] ;
 wire \load_weights[204] ;
 wire \load_weights[205] ;
 wire \load_weights[206] ;
 wire \load_weights[207] ;
 wire \load_weights[208] ;
 wire \load_weights[209] ;
 wire \load_weights[20] ;
 wire \load_weights[210] ;
 wire \load_weights[211] ;
 wire \load_weights[212] ;
 wire \load_weights[213] ;
 wire \load_weights[214] ;
 wire \load_weights[215] ;
 wire \load_weights[216] ;
 wire \load_weights[217] ;
 wire \load_weights[218] ;
 wire \load_weights[219] ;
 wire \load_weights[21] ;
 wire \load_weights[220] ;
 wire \load_weights[221] ;
 wire \load_weights[222] ;
 wire \load_weights[223] ;
 wire \load_weights[224] ;
 wire \load_weights[225] ;
 wire \load_weights[226] ;
 wire \load_weights[227] ;
 wire \load_weights[228] ;
 wire \load_weights[229] ;
 wire \load_weights[22] ;
 wire \load_weights[230] ;
 wire \load_weights[231] ;
 wire \load_weights[232] ;
 wire \load_weights[233] ;
 wire \load_weights[234] ;
 wire \load_weights[235] ;
 wire \load_weights[236] ;
 wire \load_weights[237] ;
 wire \load_weights[238] ;
 wire \load_weights[239] ;
 wire \load_weights[23] ;
 wire \load_weights[240] ;
 wire \load_weights[241] ;
 wire \load_weights[242] ;
 wire \load_weights[243] ;
 wire \load_weights[244] ;
 wire \load_weights[245] ;
 wire \load_weights[246] ;
 wire \load_weights[247] ;
 wire \load_weights[248] ;
 wire \load_weights[249] ;
 wire \load_weights[24] ;
 wire \load_weights[250] ;
 wire \load_weights[251] ;
 wire \load_weights[252] ;
 wire \load_weights[253] ;
 wire \load_weights[254] ;
 wire \load_weights[255] ;
 wire \load_weights[256] ;
 wire \load_weights[257] ;
 wire \load_weights[258] ;
 wire \load_weights[259] ;
 wire \load_weights[25] ;
 wire \load_weights[260] ;
 wire \load_weights[261] ;
 wire \load_weights[262] ;
 wire \load_weights[263] ;
 wire \load_weights[264] ;
 wire \load_weights[265] ;
 wire \load_weights[266] ;
 wire \load_weights[267] ;
 wire \load_weights[268] ;
 wire \load_weights[269] ;
 wire \load_weights[26] ;
 wire \load_weights[270] ;
 wire \load_weights[271] ;
 wire \load_weights[272] ;
 wire \load_weights[273] ;
 wire \load_weights[274] ;
 wire \load_weights[275] ;
 wire \load_weights[276] ;
 wire \load_weights[277] ;
 wire \load_weights[278] ;
 wire \load_weights[279] ;
 wire \load_weights[27] ;
 wire \load_weights[280] ;
 wire \load_weights[281] ;
 wire \load_weights[282] ;
 wire \load_weights[283] ;
 wire \load_weights[284] ;
 wire \load_weights[285] ;
 wire \load_weights[286] ;
 wire \load_weights[287] ;
 wire \load_weights[28] ;
 wire \load_weights[29] ;
 wire \load_weights[2] ;
 wire \load_weights[30] ;
 wire \load_weights[31] ;
 wire \load_weights[32] ;
 wire \load_weights[33] ;
 wire \load_weights[34] ;
 wire \load_weights[35] ;
 wire \load_weights[36] ;
 wire \load_weights[37] ;
 wire \load_weights[38] ;
 wire \load_weights[39] ;
 wire \load_weights[3] ;
 wire \load_weights[40] ;
 wire \load_weights[41] ;
 wire \load_weights[42] ;
 wire \load_weights[43] ;
 wire \load_weights[44] ;
 wire \load_weights[45] ;
 wire \load_weights[46] ;
 wire \load_weights[47] ;
 wire \load_weights[48] ;
 wire \load_weights[49] ;
 wire \load_weights[4] ;
 wire \load_weights[50] ;
 wire \load_weights[51] ;
 wire \load_weights[52] ;
 wire \load_weights[53] ;
 wire \load_weights[54] ;
 wire \load_weights[55] ;
 wire \load_weights[56] ;
 wire \load_weights[57] ;
 wire \load_weights[58] ;
 wire \load_weights[59] ;
 wire \load_weights[5] ;
 wire \load_weights[60] ;
 wire \load_weights[61] ;
 wire \load_weights[62] ;
 wire \load_weights[63] ;
 wire \load_weights[64] ;
 wire \load_weights[65] ;
 wire \load_weights[66] ;
 wire \load_weights[67] ;
 wire \load_weights[68] ;
 wire \load_weights[69] ;
 wire \load_weights[6] ;
 wire \load_weights[70] ;
 wire \load_weights[71] ;
 wire \load_weights[72] ;
 wire \load_weights[73] ;
 wire \load_weights[74] ;
 wire \load_weights[75] ;
 wire \load_weights[76] ;
 wire \load_weights[77] ;
 wire \load_weights[78] ;
 wire \load_weights[79] ;
 wire \load_weights[7] ;
 wire \load_weights[80] ;
 wire \load_weights[81] ;
 wire \load_weights[82] ;
 wire \load_weights[83] ;
 wire \load_weights[84] ;
 wire \load_weights[85] ;
 wire \load_weights[86] ;
 wire \load_weights[87] ;
 wire \load_weights[88] ;
 wire \load_weights[89] ;
 wire \load_weights[8] ;
 wire \load_weights[90] ;
 wire \load_weights[91] ;
 wire \load_weights[92] ;
 wire \load_weights[93] ;
 wire \load_weights[94] ;
 wire \load_weights[95] ;
 wire \load_weights[96] ;
 wire \load_weights[97] ;
 wire \load_weights[98] ;
 wire \load_weights[99] ;
 wire \load_weights[9] ;
 wire mult_ena;
 wire \tt_um_mult_inst.genblk1[0].carry[0] ;
 wire \tt_um_mult_inst.genblk1[0].carry[1] ;
 wire \tt_um_mult_inst.genblk1[0].carry[2] ;
 wire \tt_um_mult_inst.genblk1[0].carry[3] ;
 wire \tt_um_mult_inst.genblk1[0].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[0].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[0].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[0].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[0].out ;
 wire \tt_um_mult_inst.genblk1[0].out_q ;
 wire \tt_um_mult_inst.genblk1[10].carry[0] ;
 wire \tt_um_mult_inst.genblk1[10].carry[1] ;
 wire \tt_um_mult_inst.genblk1[10].carry[2] ;
 wire \tt_um_mult_inst.genblk1[10].carry[3] ;
 wire \tt_um_mult_inst.genblk1[10].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[10].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[10].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[10].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[10].out ;
 wire \tt_um_mult_inst.genblk1[10].out_q ;
 wire \tt_um_mult_inst.genblk1[11].carry[0] ;
 wire \tt_um_mult_inst.genblk1[11].carry[1] ;
 wire \tt_um_mult_inst.genblk1[11].carry[2] ;
 wire \tt_um_mult_inst.genblk1[11].carry[3] ;
 wire \tt_um_mult_inst.genblk1[11].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[11].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[11].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[11].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[11].out ;
 wire \tt_um_mult_inst.genblk1[11].out_q ;
 wire \tt_um_mult_inst.genblk1[1].carry[0] ;
 wire \tt_um_mult_inst.genblk1[1].carry[1] ;
 wire \tt_um_mult_inst.genblk1[1].carry[2] ;
 wire \tt_um_mult_inst.genblk1[1].carry[3] ;
 wire \tt_um_mult_inst.genblk1[1].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[1].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[1].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[1].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[1].out ;
 wire \tt_um_mult_inst.genblk1[1].out_q ;
 wire \tt_um_mult_inst.genblk1[2].carry[0] ;
 wire \tt_um_mult_inst.genblk1[2].carry[1] ;
 wire \tt_um_mult_inst.genblk1[2].carry[2] ;
 wire \tt_um_mult_inst.genblk1[2].carry[3] ;
 wire \tt_um_mult_inst.genblk1[2].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[2].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[2].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[2].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[2].out ;
 wire \tt_um_mult_inst.genblk1[2].out_q ;
 wire \tt_um_mult_inst.genblk1[3].carry[0] ;
 wire \tt_um_mult_inst.genblk1[3].carry[1] ;
 wire \tt_um_mult_inst.genblk1[3].carry[2] ;
 wire \tt_um_mult_inst.genblk1[3].carry[3] ;
 wire \tt_um_mult_inst.genblk1[3].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[3].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[3].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[3].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[3].out ;
 wire \tt_um_mult_inst.genblk1[3].out_q ;
 wire \tt_um_mult_inst.genblk1[4].carry[0] ;
 wire \tt_um_mult_inst.genblk1[4].carry[1] ;
 wire \tt_um_mult_inst.genblk1[4].carry[2] ;
 wire \tt_um_mult_inst.genblk1[4].carry[3] ;
 wire \tt_um_mult_inst.genblk1[4].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[4].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[4].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[4].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[4].out ;
 wire \tt_um_mult_inst.genblk1[4].out_q ;
 wire \tt_um_mult_inst.genblk1[5].carry[0] ;
 wire \tt_um_mult_inst.genblk1[5].carry[1] ;
 wire \tt_um_mult_inst.genblk1[5].carry[2] ;
 wire \tt_um_mult_inst.genblk1[5].carry[3] ;
 wire \tt_um_mult_inst.genblk1[5].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[5].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[5].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[5].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[5].out ;
 wire \tt_um_mult_inst.genblk1[5].out_q ;
 wire \tt_um_mult_inst.genblk1[6].carry[0] ;
 wire \tt_um_mult_inst.genblk1[6].carry[1] ;
 wire \tt_um_mult_inst.genblk1[6].carry[2] ;
 wire \tt_um_mult_inst.genblk1[6].carry[3] ;
 wire \tt_um_mult_inst.genblk1[6].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[6].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[6].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[6].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[6].out ;
 wire \tt_um_mult_inst.genblk1[6].out_q ;
 wire \tt_um_mult_inst.genblk1[7].carry[0] ;
 wire \tt_um_mult_inst.genblk1[7].carry[1] ;
 wire \tt_um_mult_inst.genblk1[7].carry[2] ;
 wire \tt_um_mult_inst.genblk1[7].carry[3] ;
 wire \tt_um_mult_inst.genblk1[7].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[7].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[7].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[7].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[7].out ;
 wire \tt_um_mult_inst.genblk1[7].out_q ;
 wire \tt_um_mult_inst.genblk1[8].carry[0] ;
 wire \tt_um_mult_inst.genblk1[8].carry[1] ;
 wire \tt_um_mult_inst.genblk1[8].carry[2] ;
 wire \tt_um_mult_inst.genblk1[8].carry[3] ;
 wire \tt_um_mult_inst.genblk1[8].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[8].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[8].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[8].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[8].out ;
 wire \tt_um_mult_inst.genblk1[8].out_q ;
 wire \tt_um_mult_inst.genblk1[9].carry[0] ;
 wire \tt_um_mult_inst.genblk1[9].carry[1] ;
 wire \tt_um_mult_inst.genblk1[9].carry[2] ;
 wire \tt_um_mult_inst.genblk1[9].carry[3] ;
 wire \tt_um_mult_inst.genblk1[9].carry_q[0] ;
 wire \tt_um_mult_inst.genblk1[9].carry_q[1] ;
 wire \tt_um_mult_inst.genblk1[9].carry_q[2] ;
 wire \tt_um_mult_inst.genblk1[9].carry_q[3] ;
 wire \tt_um_mult_inst.genblk1[9].out ;
 wire \tt_um_mult_inst.genblk1[9].out_q ;
 wire net377;
 wire net378;
 wire net379;
 wire clknet_leaf_0_clk;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net1;
 wire net2;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;

 sg13g2_o21ai_1 _2857_ (.B1(_1785_),
    .Y(_1805_),
    .A1(_1780_),
    .A2(_1786_));
 sg13g2_nand2_1 _2858_ (.Y(_1806_),
    .A(_1781_),
    .B(_1805_));
 sg13g2_xor2_1 _2859_ (.B(_1805_),
    .A(_1781_),
    .X(_1807_));
 sg13g2_or2_1 _2860_ (.X(_1808_),
    .B(_1807_),
    .A(_1804_));
 sg13g2_a21oi_1 _2861_ (.A1(_1804_),
    .A2(_1807_),
    .Y(_1809_),
    .B1(net428));
 sg13g2_a22oi_1 _2862_ (.Y(_1810_),
    .B1(_1808_),
    .B2(_1809_),
    .A2(net428),
    .A1(\tt_um_mult_inst.genblk1[2].carry[2] ));
 sg13g2_nor2_1 _2863_ (.A(_1793_),
    .B(_1810_),
    .Y(_1811_));
 sg13g2_xnor2_1 _2864_ (.Y(_1812_),
    .A(_1793_),
    .B(_1810_));
 sg13g2_a21oi_2 _2865_ (.B1(_1812_),
    .Y(_1813_),
    .A2(_1797_),
    .A1(_1795_));
 sg13g2_nand3_1 _2866_ (.B(_1797_),
    .C(_1812_),
    .A(_1795_),
    .Y(_1814_));
 sg13g2_nand2b_1 _2867_ (.Y(_1815_),
    .B(_1814_),
    .A_N(_1813_));
 sg13g2_nor2_1 _2868_ (.A(_1800_),
    .B(_1815_),
    .Y(_1816_));
 sg13g2_xor2_1 _2869_ (.B(_1815_),
    .A(_1800_),
    .X(_1817_));
 sg13g2_o21ai_1 _2870_ (.B1(_1802_),
    .Y(_1818_),
    .A1(_1773_),
    .A2(_1803_));
 sg13g2_xor2_1 _2871_ (.B(_1818_),
    .A(_1817_),
    .X(\tt_um_mult_inst.genblk1[2].carry_q[1] ));
 sg13g2_a21oi_1 _2872_ (.A1(_1817_),
    .A2(_1818_),
    .Y(_1819_),
    .B1(_1816_));
 sg13g2_a22oi_1 _2873_ (.Y(_1820_),
    .B1(_1806_),
    .B2(_1809_),
    .A2(net428),
    .A1(net918));
 sg13g2_nand2_1 _2874_ (.Y(_1821_),
    .A(_1811_),
    .B(_1820_));
 sg13g2_xor2_1 _2875_ (.B(_1820_),
    .A(_1811_),
    .X(_1822_));
 sg13g2_xor2_1 _2876_ (.B(_1822_),
    .A(_1813_),
    .X(_1823_));
 sg13g2_xnor2_1 _2877_ (.Y(\tt_um_mult_inst.genblk1[2].carry_q[2] ),
    .A(_1819_),
    .B(_1823_));
 sg13g2_nand3_1 _2878_ (.B(_1818_),
    .C(_1823_),
    .A(_1817_),
    .Y(_1824_));
 sg13g2_o21ai_1 _2879_ (.B1(_1822_),
    .Y(_1825_),
    .A1(_1813_),
    .A2(_1816_));
 sg13g2_nand3_1 _2880_ (.B(_1824_),
    .C(_1825_),
    .A(net919),
    .Y(\tt_um_mult_inst.genblk1[2].carry_q[3] ));
 sg13g2_mux2_1 _2881_ (.A0(net662),
    .A1(net523),
    .S(net487),
    .X(_0029_));
 sg13g2_mux2_1 _2882_ (.A0(net666),
    .A1(net519),
    .S(net487),
    .X(_0030_));
 sg13g2_mux2_1 _2883_ (.A0(net659),
    .A1(net513),
    .S(net488),
    .X(_0031_));
 sg13g2_mux2_1 _2884_ (.A0(net653),
    .A1(net509),
    .S(net488),
    .X(_0032_));
 sg13g2_mux2_1 _2885_ (.A0(net380),
    .A1(net560),
    .S(net479),
    .X(_0033_));
 sg13g2_mux2_1 _2886_ (.A0(net656),
    .A1(net555),
    .S(net488),
    .X(_0034_));
 sg13g2_mux2_1 _2887_ (.A0(net646),
    .A1(net550),
    .S(net481),
    .X(_0035_));
 sg13g2_mux2_1 _2888_ (.A0(net572),
    .A1(net546),
    .S(net484),
    .X(_0036_));
 sg13g2_mux2_1 _2889_ (.A0(net615),
    .A1(net541),
    .S(net478),
    .X(_0037_));
 sg13g2_mux2_1 _2890_ (.A0(net780),
    .A1(net537),
    .S(net485),
    .X(_0038_));
 sg13g2_mux2_1 _2891_ (.A0(net405),
    .A1(net532),
    .S(net481),
    .X(_0039_));
 sg13g2_mux2_1 _2892_ (.A0(net638),
    .A1(net528),
    .S(net486),
    .X(_0040_));
 sg13g2_mux2_1 _2893_ (.A0(\load_weights[12] ),
    .A1(net662),
    .S(net487),
    .X(_0041_));
 sg13g2_mux2_1 _2894_ (.A0(net756),
    .A1(net666),
    .S(net487),
    .X(_0042_));
 sg13g2_mux2_1 _2895_ (.A0(net773),
    .A1(net659),
    .S(net488),
    .X(_0043_));
 sg13g2_mux2_1 _2896_ (.A0(net698),
    .A1(net653),
    .S(net487),
    .X(_0044_));
 sg13g2_nand2_1 _2897_ (.Y(_1826_),
    .A(net479),
    .B(net380));
 sg13g2_o21ai_1 _2898_ (.B1(_1826_),
    .Y(_0045_),
    .A1(net479),
    .A2(_1956_));
 sg13g2_mux2_1 _2899_ (.A0(net604),
    .A1(net656),
    .S(net488),
    .X(_0046_));
 sg13g2_mux2_1 _2900_ (.A0(net651),
    .A1(net646),
    .S(net480),
    .X(_0047_));
 sg13g2_mux2_1 _2901_ (.A0(\load_weights[19] ),
    .A1(net572),
    .S(net484),
    .X(_0048_));
 sg13g2_mux2_1 _2902_ (.A0(\load_weights[20] ),
    .A1(net615),
    .S(net479),
    .X(_0049_));
 sg13g2_mux2_1 _2903_ (.A0(net761),
    .A1(net780),
    .S(net485),
    .X(_0050_));
 sg13g2_nand2_1 _2904_ (.Y(_1827_),
    .A(net479),
    .B(net405));
 sg13g2_o21ai_1 _2905_ (.B1(_1827_),
    .Y(_0051_),
    .A1(net478),
    .A2(_1957_));
 sg13g2_mux2_1 _2906_ (.A0(net676),
    .A1(net638),
    .S(net484),
    .X(_0052_));
 sg13g2_mux2_1 _2907_ (.A0(net747),
    .A1(net798),
    .S(net487),
    .X(_0053_));
 sg13g2_mux2_1 _2908_ (.A0(net682),
    .A1(\load_weights[13] ),
    .S(net487),
    .X(_0054_));
 sg13g2_mux2_1 _2909_ (.A0(net886),
    .A1(net773),
    .S(net484),
    .X(_0055_));
 sg13g2_mux2_1 _2910_ (.A0(net386),
    .A1(net698),
    .S(net488),
    .X(_0056_));
 sg13g2_nor2_1 _2911_ (.A(net487),
    .B(net647),
    .Y(_1828_));
 sg13g2_a21oi_1 _2912_ (.A1(net478),
    .A2(_1956_),
    .Y(_0057_),
    .B1(_1828_));
 sg13g2_mux2_1 _2913_ (.A0(net384),
    .A1(net604),
    .S(net484),
    .X(_0058_));
 sg13g2_mux2_1 _2914_ (.A0(net707),
    .A1(net651),
    .S(net479),
    .X(_0059_));
 sg13g2_mux2_1 _2915_ (.A0(net416),
    .A1(net608),
    .S(net485),
    .X(_0060_));
 sg13g2_mux2_1 _2916_ (.A0(net619),
    .A1(\load_weights[20] ),
    .S(net478),
    .X(_0061_));
 sg13g2_mux2_1 _2917_ (.A0(net711),
    .A1(net761),
    .S(net485),
    .X(_0062_));
 sg13g2_nor2_1 _2918_ (.A(net478),
    .B(net579),
    .Y(_1829_));
 sg13g2_a21oi_1 _2919_ (.A1(net478),
    .A2(_1957_),
    .Y(_0063_),
    .B1(_1829_));
 sg13g2_mux2_1 _2920_ (.A0(net791),
    .A1(net676),
    .S(net483),
    .X(_0064_));
 sg13g2_mux2_1 _2921_ (.A0(net700),
    .A1(net747),
    .S(net483),
    .X(_0065_));
 sg13g2_mux2_1 _2922_ (.A0(net702),
    .A1(net682),
    .S(net483),
    .X(_0066_));
 sg13g2_mux2_1 _2923_ (.A0(net887),
    .A1(net886),
    .S(net482),
    .X(_0067_));
 sg13g2_nand2_1 _2924_ (.Y(_1830_),
    .A(net484),
    .B(net386));
 sg13g2_o21ai_1 _2925_ (.B1(_1830_),
    .Y(_0068_),
    .A1(net484),
    .A2(_1951_));
 sg13g2_mux2_1 _2926_ (.A0(net868),
    .A1(net647),
    .S(net483),
    .X(_0069_));
 sg13g2_nand2_1 _2927_ (.Y(_1831_),
    .A(net484),
    .B(net384));
 sg13g2_o21ai_1 _2928_ (.B1(_1831_),
    .Y(_0070_),
    .A1(net485),
    .A2(_1950_));
 sg13g2_mux2_1 _2929_ (.A0(net804),
    .A1(net707),
    .S(net478),
    .X(_0071_));
 sg13g2_nand2_1 _2930_ (.Y(_1832_),
    .A(net485),
    .B(net416));
 sg13g2_o21ai_1 _2931_ (.B1(_1832_),
    .Y(_0072_),
    .A1(net485),
    .A2(_1949_));
 sg13g2_mux2_1 _2932_ (.A0(net640),
    .A1(net619),
    .S(net478),
    .X(_0073_));
 sg13g2_mux2_1 _2933_ (.A0(\load_weights[45] ),
    .A1(net711),
    .S(net485),
    .X(_0074_));
 sg13g2_mux2_1 _2934_ (.A0(net834),
    .A1(net579),
    .S(net479),
    .X(_0075_));
 sg13g2_mux2_1 _2935_ (.A0(net818),
    .A1(net791),
    .S(net482),
    .X(_0076_));
 sg13g2_mux2_1 _2936_ (.A0(net566),
    .A1(net700),
    .S(net476),
    .X(_0077_));
 sg13g2_mux2_1 _2937_ (.A0(net771),
    .A1(net702),
    .S(net476),
    .X(_0078_));
 sg13g2_mux2_1 _2938_ (.A0(net792),
    .A1(\load_weights[38] ),
    .S(net482),
    .X(_0079_));
 sg13g2_nor2_1 _2939_ (.A(net483),
    .B(net750),
    .Y(_1833_));
 sg13g2_a21oi_1 _2940_ (.A1(net483),
    .A2(_1951_),
    .Y(_0080_),
    .B1(_1833_));
 sg13g2_mux2_1 _2941_ (.A0(net799),
    .A1(\load_weights[40] ),
    .S(net476),
    .X(_0081_));
 sg13g2_nor2_1 _2942_ (.A(net482),
    .B(net408),
    .Y(_1834_));
 sg13g2_a21oi_1 _2943_ (.A1(net482),
    .A2(_1950_),
    .Y(_0082_),
    .B1(_1834_));
 sg13g2_mux2_1 _2944_ (.A0(net742),
    .A1(\load_weights[42] ),
    .S(net480),
    .X(_0083_));
 sg13g2_nor2_1 _2945_ (.A(net476),
    .B(net420),
    .Y(_1835_));
 sg13g2_a21oi_1 _2946_ (.A1(net482),
    .A2(_1949_),
    .Y(_0084_),
    .B1(_1835_));
 sg13g2_mux2_1 _2947_ (.A0(net631),
    .A1(net640),
    .S(net480),
    .X(_0085_));
 sg13g2_mux2_1 _2948_ (.A0(net719),
    .A1(net885),
    .S(net482),
    .X(_0086_));
 sg13g2_mux2_1 _2949_ (.A0(net654),
    .A1(\load_weights[46] ),
    .S(net480),
    .X(_0087_));
 sg13g2_mux2_1 _2950_ (.A0(\load_weights[59] ),
    .A1(net818),
    .S(net482),
    .X(_0088_));
 sg13g2_mux2_1 _2951_ (.A0(\load_weights[60] ),
    .A1(net566),
    .S(net481),
    .X(_0089_));
 sg13g2_mux2_1 _2952_ (.A0(\load_weights[61] ),
    .A1(net771),
    .S(net477),
    .X(_0090_));
 sg13g2_mux2_1 _2953_ (.A0(net827),
    .A1(net792),
    .S(net476),
    .X(_0091_));
 sg13g2_nand2_1 _2954_ (.Y(_1836_),
    .A(net477),
    .B(net750));
 sg13g2_o21ai_1 _2955_ (.B1(_1836_),
    .Y(_0092_),
    .A1(net477),
    .A2(_1963_));
 sg13g2_mux2_1 _2956_ (.A0(net806),
    .A1(net799),
    .S(net476),
    .X(_0093_));
 sg13g2_mux2_1 _2957_ (.A0(net796),
    .A1(net408),
    .S(net476),
    .X(_0094_));
 sg13g2_mux2_1 _2958_ (.A0(net745),
    .A1(net742),
    .S(net480),
    .X(_0095_));
 sg13g2_mux2_1 _2959_ (.A0(net828),
    .A1(net420),
    .S(net476),
    .X(_0096_));
 sg13g2_mux2_1 _2960_ (.A0(\load_weights[68] ),
    .A1(net631),
    .S(net480),
    .X(_0097_));
 sg13g2_nand2_1 _2961_ (.Y(_1837_),
    .A(net477),
    .B(net719));
 sg13g2_o21ai_1 _2962_ (.B1(_1837_),
    .Y(_0098_),
    .A1(net477),
    .A2(_1962_));
 sg13g2_mux2_1 _2963_ (.A0(net783),
    .A1(net654),
    .S(net480),
    .X(_0099_));
 sg13g2_mux2_1 _2964_ (.A0(net850),
    .A1(net867),
    .S(net477),
    .X(_0100_));
 sg13g2_mux2_1 _2965_ (.A0(net786),
    .A1(\load_weights[60] ),
    .S(net477),
    .X(_0101_));
 sg13g2_mux2_1 _2966_ (.A0(net733),
    .A1(\load_weights[61] ),
    .S(net453),
    .X(_0102_));
 sg13g2_mux2_1 _2967_ (.A0(net902),
    .A1(net827),
    .S(net452),
    .X(_0103_));
 sg13g2_nor2_1 _2968_ (.A(net453),
    .B(net592),
    .Y(_1838_));
 sg13g2_a21oi_1 _2969_ (.A1(net453),
    .A2(_1963_),
    .Y(_0104_),
    .B1(_1838_));
 sg13g2_mux2_1 _2970_ (.A0(net911),
    .A1(net806),
    .S(net452),
    .X(_0105_));
 sg13g2_mux2_1 _2971_ (.A0(net753),
    .A1(net796),
    .S(net453),
    .X(_0106_));
 sg13g2_mux2_1 _2972_ (.A0(net810),
    .A1(net745),
    .S(net458),
    .X(_0107_));
 sg13g2_mux2_1 _2973_ (.A0(net674),
    .A1(\load_weights[67] ),
    .S(net452),
    .X(_0108_));
 sg13g2_mux2_1 _2974_ (.A0(net808),
    .A1(\load_weights[68] ),
    .S(net458),
    .X(_0109_));
 sg13g2_nor2_1 _2975_ (.A(net452),
    .B(net415),
    .Y(_1839_));
 sg13g2_a21oi_1 _2976_ (.A1(net452),
    .A2(_1962_),
    .Y(_0110_),
    .B1(_1839_));
 sg13g2_mux2_1 _2977_ (.A0(net837),
    .A1(net783),
    .S(net458),
    .X(_0111_));
 sg13g2_mux2_1 _2978_ (.A0(net841),
    .A1(net850),
    .S(net452),
    .X(_0112_));
 sg13g2_mux2_1 _2979_ (.A0(net824),
    .A1(net786),
    .S(net453),
    .X(_0113_));
 sg13g2_mux2_1 _2980_ (.A0(net716),
    .A1(net733),
    .S(net453),
    .X(_0114_));
 sg13g2_mux2_1 _2981_ (.A0(\load_weights[86] ),
    .A1(net902),
    .S(net451),
    .X(_0115_));
 sg13g2_nand2_1 _2982_ (.Y(_1840_),
    .A(net452),
    .B(net592));
 sg13g2_o21ai_1 _2983_ (.B1(_1840_),
    .Y(_0116_),
    .A1(net451),
    .A2(_1943_));
 sg13g2_mux2_1 _2984_ (.A0(net913),
    .A1(net911),
    .S(net443),
    .X(_0117_));
 sg13g2_mux2_1 _2985_ (.A0(net630),
    .A1(net753),
    .S(net453),
    .X(_0118_));
 sg13g2_mux2_1 _2986_ (.A0(net869),
    .A1(net810),
    .S(net458),
    .X(_0119_));
 sg13g2_mux2_1 _2987_ (.A0(net639),
    .A1(net674),
    .S(net452),
    .X(_0120_));
 sg13g2_mux2_1 _2988_ (.A0(net860),
    .A1(net808),
    .S(net457),
    .X(_0121_));
 sg13g2_nand2_1 _2989_ (.Y(_1841_),
    .A(net451),
    .B(net415));
 sg13g2_o21ai_1 _2990_ (.B1(_1841_),
    .Y(_0122_),
    .A1(net451),
    .A2(_1942_));
 sg13g2_mux2_1 _2991_ (.A0(net844),
    .A1(net837),
    .S(net457),
    .X(_0123_));
 sg13g2_mux2_1 _2992_ (.A0(net778),
    .A1(net841),
    .S(net451),
    .X(_0124_));
 sg13g2_mux2_1 _2993_ (.A0(net704),
    .A1(\load_weights[84] ),
    .S(net445),
    .X(_0125_));
 sg13g2_mux2_1 _2994_ (.A0(net677),
    .A1(net716),
    .S(net443),
    .X(_0126_));
 sg13g2_mux2_1 _2995_ (.A0(net684),
    .A1(\load_weights[86] ),
    .S(net443),
    .X(_0127_));
 sg13g2_nor2_1 _2996_ (.A(net451),
    .B(net606),
    .Y(_1842_));
 sg13g2_a21oi_1 _2997_ (.A1(net451),
    .A2(_1943_),
    .Y(_0128_),
    .B1(_1842_));
 sg13g2_mux2_1 _2998_ (.A0(net660),
    .A1(\load_weights[88] ),
    .S(net443),
    .X(_0129_));
 sg13g2_mux2_1 _2999_ (.A0(net388),
    .A1(net630),
    .S(net454),
    .X(_0130_));
 sg13g2_mux2_1 _3000_ (.A0(net896),
    .A1(net869),
    .S(net444),
    .X(_0131_));
 sg13g2_mux2_1 _3001_ (.A0(net382),
    .A1(net639),
    .S(net451),
    .X(_0132_));
 sg13g2_mux2_1 _3002_ (.A0(net851),
    .A1(\load_weights[92] ),
    .S(net444),
    .X(_0133_));
 sg13g2_nor2_1 _3003_ (.A(net443),
    .B(net413),
    .Y(_1843_));
 sg13g2_a21oi_1 _3004_ (.A1(net443),
    .A2(_1942_),
    .Y(_0134_),
    .B1(_1843_));
 sg13g2_mux2_1 _3005_ (.A0(net854),
    .A1(net844),
    .S(net455),
    .X(_0135_));
 sg13g2_mux2_1 _3006_ (.A0(net754),
    .A1(net778),
    .S(net443),
    .X(_0136_));
 sg13g2_mux2_1 _3007_ (.A0(net708),
    .A1(net704),
    .S(net445),
    .X(_0137_));
 sg13g2_mux2_1 _3008_ (.A0(\load_weights[109] ),
    .A1(net677),
    .S(net444),
    .X(_0138_));
 sg13g2_mux2_1 _3009_ (.A0(net727),
    .A1(net684),
    .S(net445),
    .X(_0139_));
 sg13g2_nand2_1 _3010_ (.Y(_1844_),
    .A(net449),
    .B(net606));
 sg13g2_o21ai_1 _3011_ (.B1(_1844_),
    .Y(_0140_),
    .A1(net449),
    .A2(_1948_));
 sg13g2_mux2_1 _3012_ (.A0(net717),
    .A1(net660),
    .S(net445),
    .X(_0141_));
 sg13g2_nand2_1 _3013_ (.Y(_1845_),
    .A(net455),
    .B(net388));
 sg13g2_o21ai_1 _3014_ (.B1(_1845_),
    .Y(_0142_),
    .A1(net455),
    .A2(_1945_));
 sg13g2_mux2_1 _3015_ (.A0(net898),
    .A1(net896),
    .S(net445),
    .X(_0143_));
 sg13g2_nand2_1 _3016_ (.Y(_1846_),
    .A(net444),
    .B(net382));
 sg13g2_o21ai_1 _3017_ (.B1(_1846_),
    .Y(_0144_),
    .A1(net444),
    .A2(_1946_));
 sg13g2_mux2_1 _3018_ (.A0(net876),
    .A1(net851),
    .S(net447),
    .X(_0145_));
 sg13g2_nand2_1 _3019_ (.Y(_1847_),
    .A(net444),
    .B(net413));
 sg13g2_o21ai_1 _3020_ (.B1(_1847_),
    .Y(_0146_),
    .A1(net443),
    .A2(_1947_));
 sg13g2_mux2_1 _3021_ (.A0(net587),
    .A1(net854),
    .S(net449),
    .X(_0147_));
 sg13g2_mux2_1 _3022_ (.A0(\load_weights[119] ),
    .A1(net754),
    .S(net444),
    .X(_0148_));
 sg13g2_mux2_1 _3023_ (.A0(net746),
    .A1(net708),
    .S(net446),
    .X(_0149_));
 sg13g2_mux2_1 _3024_ (.A0(net590),
    .A1(\load_weights[109] ),
    .S(net447),
    .X(_0150_));
 sg13g2_mux2_1 _3025_ (.A0(net644),
    .A1(\load_weights[110] ),
    .S(net446),
    .X(_0151_));
 sg13g2_nor2_1 _3026_ (.A(net449),
    .B(net394),
    .Y(_1848_));
 sg13g2_a21oi_1 _3027_ (.A1(net449),
    .A2(_1948_),
    .Y(_0152_),
    .B1(_1848_));
 sg13g2_mux2_1 _3028_ (.A0(net718),
    .A1(net717),
    .S(net446),
    .X(_0153_));
 sg13g2_nor2_1 _3029_ (.A(net455),
    .B(net392),
    .Y(_1849_));
 sg13g2_a21oi_1 _3030_ (.A1(net455),
    .A2(_1945_),
    .Y(_0154_),
    .B1(_1849_));
 sg13g2_mux2_1 _3031_ (.A0(net822),
    .A1(\load_weights[114] ),
    .S(net446),
    .X(_0155_));
 sg13g2_nor2_1 _3032_ (.A(net455),
    .B(net418),
    .Y(_1850_));
 sg13g2_a21oi_1 _3033_ (.A1(net455),
    .A2(_1946_),
    .Y(_0156_),
    .B1(_1850_));
 sg13g2_mux2_1 _3034_ (.A0(net585),
    .A1(\load_weights[116] ),
    .S(net446),
    .X(_0157_));
 sg13g2_nor2_1 _3035_ (.A(net455),
    .B(net398),
    .Y(_1851_));
 sg13g2_a21oi_1 _3036_ (.A1(net449),
    .A2(_1947_),
    .Y(_0158_),
    .B1(_1851_));
 sg13g2_mux2_1 _3037_ (.A0(net583),
    .A1(net587),
    .S(net447),
    .X(_0159_));
 sg13g2_mux2_1 _3038_ (.A0(\load_weights[131] ),
    .A1(net757),
    .S(net449),
    .X(_0160_));
 sg13g2_mux2_1 _3039_ (.A0(net703),
    .A1(net746),
    .S(net446),
    .X(_0161_));
 sg13g2_mux2_1 _3040_ (.A0(net614),
    .A1(net590),
    .S(net447),
    .X(_0162_));
 sg13g2_mux2_1 _3041_ (.A0(net736),
    .A1(net644),
    .S(net446),
    .X(_0163_));
 sg13g2_nand2_1 _3042_ (.Y(_1852_),
    .A(net449),
    .B(net394));
 sg13g2_o21ai_1 _3043_ (.B1(_1852_),
    .Y(_0164_),
    .A1(net456),
    .A2(_1955_));
 sg13g2_mux2_1 _3044_ (.A0(net664),
    .A1(net718),
    .S(net448),
    .X(_0165_));
 sg13g2_nand2_1 _3045_ (.Y(_1853_),
    .A(net457),
    .B(net392));
 sg13g2_o21ai_1 _3046_ (.B1(_1853_),
    .Y(_0166_),
    .A1(net456),
    .A2(_1953_));
 sg13g2_mux2_1 _3047_ (.A0(net849),
    .A1(net822),
    .S(net446),
    .X(_0167_));
 sg13g2_nand2_1 _3048_ (.Y(_1854_),
    .A(net456),
    .B(net418));
 sg13g2_o21ai_1 _3049_ (.B1(_1854_),
    .Y(_0168_),
    .A1(net456),
    .A2(_1952_));
 sg13g2_mux2_1 _3050_ (.A0(net617),
    .A1(net585),
    .S(net448),
    .X(_0169_));
 sg13g2_nand2_1 _3051_ (.Y(_1855_),
    .A(net456),
    .B(net398));
 sg13g2_o21ai_1 _3052_ (.B1(_1855_),
    .Y(_0170_),
    .A1(net456),
    .A2(_1954_));
 sg13g2_mux2_1 _3053_ (.A0(\load_weights[142] ),
    .A1(net583),
    .S(net448),
    .X(_0171_));
 sg13g2_mux2_1 _3054_ (.A0(\load_weights[143] ),
    .A1(net825),
    .S(net450),
    .X(_0172_));
 sg13g2_mux2_1 _3055_ (.A0(net588),
    .A1(net703),
    .S(net448),
    .X(_0173_));
 sg13g2_mux2_1 _3056_ (.A0(net618),
    .A1(net614),
    .S(net460),
    .X(_0174_));
 sg13g2_mux2_1 _3057_ (.A0(net600),
    .A1(\load_weights[134] ),
    .S(net459),
    .X(_0175_));
 sg13g2_nor2_1 _3058_ (.A(net461),
    .B(net605),
    .Y(_1856_));
 sg13g2_a21oi_1 _3059_ (.A1(net461),
    .A2(_1955_),
    .Y(_0176_),
    .B1(_1856_));
 sg13g2_mux2_1 _3060_ (.A0(net401),
    .A1(net664),
    .S(net459),
    .X(_0177_));
 sg13g2_nor2_1 _3061_ (.A(net467),
    .B(net720),
    .Y(_1857_));
 sg13g2_a21oi_1 _3062_ (.A1(net456),
    .A2(_1953_),
    .Y(_0178_),
    .B1(_1857_));
 sg13g2_mux2_1 _3063_ (.A0(net687),
    .A1(\load_weights[138] ),
    .S(net459),
    .X(_0179_));
 sg13g2_nor2_1 _3064_ (.A(net467),
    .B(net633),
    .Y(_1858_));
 sg13g2_a21oi_1 _3065_ (.A1(net467),
    .A2(_1952_),
    .Y(_0180_),
    .B1(_1858_));
 sg13g2_mux2_1 _3066_ (.A0(net779),
    .A1(net617),
    .S(net459),
    .X(_0181_));
 sg13g2_nor2_1 _3067_ (.A(net467),
    .B(net691),
    .Y(_1859_));
 sg13g2_a21oi_1 _3068_ (.A1(net456),
    .A2(_1954_),
    .Y(_0182_),
    .B1(_1859_));
 sg13g2_mux2_1 _3069_ (.A0(net390),
    .A1(net713),
    .S(net459),
    .X(_0183_));
 sg13g2_mux2_1 _3070_ (.A0(net612),
    .A1(\load_weights[143] ),
    .S(net461),
    .X(_0184_));
 sg13g2_mux2_1 _3071_ (.A0(\load_weights[156] ),
    .A1(net588),
    .S(net459),
    .X(_0185_));
 sg13g2_mux2_1 _3072_ (.A0(net672),
    .A1(net618),
    .S(net459),
    .X(_0186_));
 sg13g2_mux2_1 _3073_ (.A0(net611),
    .A1(net600),
    .S(net459),
    .X(_0187_));
 sg13g2_mux2_1 _3074_ (.A0(net853),
    .A1(net605),
    .S(net461),
    .X(_0188_));
 sg13g2_nand2_1 _3075_ (.Y(_1860_),
    .A(net460),
    .B(net401));
 sg13g2_o21ai_1 _3076_ (.B1(_1860_),
    .Y(_0189_),
    .A1(net460),
    .A2(_1940_));
 sg13g2_mux2_1 _3077_ (.A0(\load_weights[161] ),
    .A1(net720),
    .S(net467),
    .X(_0190_));
 sg13g2_mux2_1 _3078_ (.A0(net729),
    .A1(net687),
    .S(net462),
    .X(_0191_));
 sg13g2_mux2_1 _3079_ (.A0(net710),
    .A1(net633),
    .S(net461),
    .X(_0192_));
 sg13g2_mux2_1 _3080_ (.A0(net785),
    .A1(net779),
    .S(net460),
    .X(_0193_));
 sg13g2_mux2_1 _3081_ (.A0(\load_weights[165] ),
    .A1(net691),
    .S(net467),
    .X(_0194_));
 sg13g2_nand2_1 _3082_ (.Y(_1861_),
    .A(net460),
    .B(net390));
 sg13g2_o21ai_1 _3083_ (.B1(_1861_),
    .Y(_0195_),
    .A1(net460),
    .A2(_1939_));
 sg13g2_mux2_1 _3084_ (.A0(net723),
    .A1(net612),
    .S(net461),
    .X(_0196_));
 sg13g2_mux2_1 _3085_ (.A0(net621),
    .A1(\load_weights[156] ),
    .S(net460),
    .X(_0197_));
 sg13g2_mux2_1 _3086_ (.A0(net628),
    .A1(\load_weights[157] ),
    .S(net462),
    .X(_0198_));
 sg13g2_mux2_1 _3087_ (.A0(net701),
    .A1(net611),
    .S(net463),
    .X(_0199_));
 sg13g2_mux2_1 _3088_ (.A0(net668),
    .A1(\load_weights[159] ),
    .S(net466),
    .X(_0200_));
 sg13g2_nor2_1 _3089_ (.A(net463),
    .B(net570),
    .Y(_1862_));
 sg13g2_a21oi_1 _3090_ (.A1(net463),
    .A2(_1940_),
    .Y(_0201_),
    .B1(_1862_));
 sg13g2_mux2_1 _3091_ (.A0(net649),
    .A1(\load_weights[161] ),
    .S(net461),
    .X(_0202_));
 sg13g2_mux2_1 _3092_ (.A0(net680),
    .A1(net729),
    .S(net463),
    .X(_0203_));
 sg13g2_mux2_1 _3093_ (.A0(net594),
    .A1(\load_weights[163] ),
    .S(net468),
    .X(_0204_));
 sg13g2_mux2_1 _3094_ (.A0(net626),
    .A1(\load_weights[164] ),
    .S(net463),
    .X(_0205_));
 sg13g2_mux2_1 _3095_ (.A0(net576),
    .A1(\load_weights[165] ),
    .S(net468),
    .X(_0206_));
 sg13g2_nor2_1 _3096_ (.A(net464),
    .B(net396),
    .Y(_1863_));
 sg13g2_a21oi_1 _3097_ (.A1(net464),
    .A2(_1939_),
    .Y(_0207_),
    .B1(_1863_));
 sg13g2_mux2_1 _3098_ (.A0(net695),
    .A1(\load_weights[167] ),
    .S(net461),
    .X(_0208_));
 sg13g2_mux2_1 _3099_ (.A0(net643),
    .A1(net621),
    .S(net463),
    .X(_0209_));
 sg13g2_mux2_1 _3100_ (.A0(net739),
    .A1(net628),
    .S(net474),
    .X(_0210_));
 sg13g2_mux2_1 _3101_ (.A0(net767),
    .A1(net701),
    .S(net463),
    .X(_0211_));
 sg13g2_mux2_1 _3102_ (.A0(net759),
    .A1(net668),
    .S(net466),
    .X(_0212_));
 sg13g2_nand2_1 _3103_ (.Y(_1864_),
    .A(net464),
    .B(net570));
 sg13g2_o21ai_1 _3104_ (.B1(_1864_),
    .Y(_0213_),
    .A1(net464),
    .A2(_1960_));
 sg13g2_mux2_1 _3105_ (.A0(net803),
    .A1(net649),
    .S(net474),
    .X(_0214_));
 sg13g2_mux2_1 _3106_ (.A0(\load_weights[186] ),
    .A1(net680),
    .S(net464),
    .X(_0215_));
 sg13g2_mux2_1 _3107_ (.A0(net610),
    .A1(net594),
    .S(net468),
    .X(_0216_));
 sg13g2_mux2_1 _3108_ (.A0(net732),
    .A1(net626),
    .S(net463),
    .X(_0217_));
 sg13g2_mux2_1 _3109_ (.A0(net697),
    .A1(net576),
    .S(net468),
    .X(_0218_));
 sg13g2_nand2_1 _3110_ (.Y(_1865_),
    .A(net465),
    .B(net396));
 sg13g2_o21ai_1 _3111_ (.B1(_1865_),
    .Y(_0219_),
    .A1(net465),
    .A2(_1959_));
 sg13g2_mux2_1 _3112_ (.A0(net744),
    .A1(net695),
    .S(net468),
    .X(_0220_));
 sg13g2_mux2_1 _3113_ (.A0(net789),
    .A1(net643),
    .S(net468),
    .X(_0221_));
 sg13g2_mux2_1 _3114_ (.A0(net714),
    .A1(net739),
    .S(net470),
    .X(_0222_));
 sg13g2_mux2_1 _3115_ (.A0(net689),
    .A1(\load_weights[182] ),
    .S(net469),
    .X(_0223_));
 sg13g2_mux2_1 _3116_ (.A0(net805),
    .A1(net759),
    .S(net468),
    .X(_0224_));
 sg13g2_nor2_1 _3117_ (.A(net470),
    .B(net830),
    .Y(_1866_));
 sg13g2_a21oi_1 _3118_ (.A1(net472),
    .A2(_1960_),
    .Y(_0225_),
    .B1(_1866_));
 sg13g2_mux2_1 _3119_ (.A0(net748),
    .A1(\load_weights[185] ),
    .S(net470),
    .X(_0226_));
 sg13g2_mux2_1 _3120_ (.A0(net861),
    .A1(\load_weights[186] ),
    .S(net474),
    .X(_0227_));
 sg13g2_mux2_1 _3121_ (.A0(net835),
    .A1(net610),
    .S(net467),
    .X(_0228_));
 sg13g2_mux2_1 _3122_ (.A0(net811),
    .A1(net732),
    .S(net472),
    .X(_0229_));
 sg13g2_mux2_1 _3123_ (.A0(net797),
    .A1(net697),
    .S(net467),
    .X(_0230_));
 sg13g2_nor2_1 _3124_ (.A(net472),
    .B(net846),
    .Y(_1867_));
 sg13g2_a21oi_1 _3125_ (.A1(net472),
    .A2(_1959_),
    .Y(_0231_),
    .B1(_1867_));
 sg13g2_mux2_1 _3126_ (.A0(net848),
    .A1(net744),
    .S(net468),
    .X(_0232_));
 sg13g2_mux2_1 _3127_ (.A0(\load_weights[204] ),
    .A1(net789),
    .S(net490),
    .X(_0233_));
 sg13g2_mux2_1 _3128_ (.A0(\load_weights[205] ),
    .A1(net714),
    .S(net490),
    .X(_0234_));
 sg13g2_mux2_1 _3129_ (.A0(net784),
    .A1(net689),
    .S(net469),
    .X(_0235_));
 sg13g2_mux2_1 _3130_ (.A0(net842),
    .A1(net805),
    .S(net470),
    .X(_0236_));
 sg13g2_nand2_1 _3131_ (.Y(_1868_),
    .A(net469),
    .B(net830));
 sg13g2_o21ai_1 _3132_ (.B1(_1868_),
    .Y(_0237_),
    .A1(net469),
    .A2(_1937_));
 sg13g2_mux2_1 _3133_ (.A0(net815),
    .A1(net748),
    .S(net490),
    .X(_0238_));
 sg13g2_mux2_1 _3134_ (.A0(net863),
    .A1(net861),
    .S(net469),
    .X(_0239_));
 sg13g2_mux2_1 _3135_ (.A0(\load_weights[211] ),
    .A1(net835),
    .S(net469),
    .X(_0240_));
 sg13g2_mux2_1 _3136_ (.A0(net829),
    .A1(net811),
    .S(net470),
    .X(_0241_));
 sg13g2_mux2_1 _3137_ (.A0(net820),
    .A1(net797),
    .S(net469),
    .X(_0242_));
 sg13g2_nand2_1 _3138_ (.Y(_1869_),
    .A(net470),
    .B(net846));
 sg13g2_o21ai_1 _3139_ (.B1(_1869_),
    .Y(_0243_),
    .A1(net490),
    .A2(_1936_));
 sg13g2_mux2_1 _3140_ (.A0(net855),
    .A1(net848),
    .S(net469),
    .X(_0244_));
 sg13g2_mux2_1 _3141_ (.A0(net914),
    .A1(\load_weights[204] ),
    .S(net490),
    .X(_0245_));
 sg13g2_mux2_1 _3142_ (.A0(net858),
    .A1(\load_weights[205] ),
    .S(net490),
    .X(_0246_));
 sg13g2_mux2_1 _3143_ (.A0(net890),
    .A1(net784),
    .S(net493),
    .X(_0247_));
 sg13g2_mux2_1 _3144_ (.A0(net774),
    .A1(\load_weights[207] ),
    .S(net490),
    .X(_0248_));
 sg13g2_nor2_1 _3145_ (.A(net499),
    .B(net410),
    .Y(_1870_));
 sg13g2_a21oi_1 _3146_ (.A1(net499),
    .A2(_1937_),
    .Y(_0249_),
    .B1(_1870_));
 sg13g2_mux2_1 _3147_ (.A0(net882),
    .A1(net815),
    .S(net491),
    .X(_0250_));
 sg13g2_mux2_1 _3148_ (.A0(net838),
    .A1(\load_weights[210] ),
    .S(net491),
    .X(_0251_));
 sg13g2_mux2_1 _3149_ (.A0(net724),
    .A1(\load_weights[211] ),
    .S(net491),
    .X(_0252_));
 sg13g2_mux2_1 _3150_ (.A0(net888),
    .A1(net829),
    .S(net490),
    .X(_0253_));
 sg13g2_mux2_1 _3151_ (.A0(net769),
    .A1(net820),
    .S(net491),
    .X(_0254_));
 sg13g2_nor2_1 _3152_ (.A(net491),
    .B(net564),
    .Y(_1871_));
 sg13g2_a21oi_1 _3153_ (.A1(net491),
    .A2(_1936_),
    .Y(_0255_),
    .B1(_1871_));
 sg13g2_mux2_1 _3154_ (.A0(net763),
    .A1(\load_weights[215] ),
    .S(net491),
    .X(_0256_));
 sg13g2_mux2_1 _3155_ (.A0(net909),
    .A1(\load_weights[216] ),
    .S(net503),
    .X(_0257_));
 sg13g2_mux2_1 _3156_ (.A0(net899),
    .A1(net858),
    .S(net492),
    .X(_0258_));
 sg13g2_mux2_1 _3157_ (.A0(\load_weights[230] ),
    .A1(net890),
    .S(net500),
    .X(_0259_));
 sg13g2_mux2_1 _3158_ (.A0(net625),
    .A1(net774),
    .S(net492),
    .X(_0260_));
 sg13g2_nand2_1 _3159_ (.Y(_1872_),
    .A(net499),
    .B(net410));
 sg13g2_o21ai_1 _3160_ (.B1(_1872_),
    .Y(_0261_),
    .A1(net499),
    .A2(_1931_));
 sg13g2_mux2_1 _3161_ (.A0(net906),
    .A1(net882),
    .S(net500),
    .X(_0262_));
 sg13g2_mux2_1 _3162_ (.A0(net879),
    .A1(net838),
    .S(net499),
    .X(_0263_));
 sg13g2_mux2_1 _3163_ (.A0(net762),
    .A1(net724),
    .S(net491),
    .X(_0264_));
 sg13g2_mux2_1 _3164_ (.A0(net905),
    .A1(net888),
    .S(net500),
    .X(_0265_));
 sg13g2_mux2_1 _3165_ (.A0(\load_weights[237] ),
    .A1(net769),
    .S(net499),
    .X(_0266_));
 sg13g2_nand2_1 _3166_ (.Y(_1873_),
    .A(net500),
    .B(net564));
 sg13g2_o21ai_1 _3167_ (.B1(_1873_),
    .Y(_0267_),
    .A1(net499),
    .A2(_1930_));
 sg13g2_mux2_1 _3168_ (.A0(net788),
    .A1(net763),
    .S(net492),
    .X(_0268_));
 sg13g2_mux2_1 _3169_ (.A0(net812),
    .A1(\load_weights[228] ),
    .S(net503),
    .X(_0269_));
 sg13g2_mux2_1 _3170_ (.A0(net602),
    .A1(\load_weights[229] ),
    .S(net492),
    .X(_0270_));
 sg13g2_mux2_1 _3171_ (.A0(net635),
    .A1(\load_weights[230] ),
    .S(net501),
    .X(_0271_));
 sg13g2_mux2_1 _3172_ (.A0(net598),
    .A1(net625),
    .S(net496),
    .X(_0272_));
 sg13g2_nor2_1 _3173_ (.A(net501),
    .B(net581),
    .Y(_1874_));
 sg13g2_a21oi_1 _3174_ (.A1(net501),
    .A2(_1931_),
    .Y(_0273_),
    .B1(_1874_));
 sg13g2_mux2_1 _3175_ (.A0(net730),
    .A1(\load_weights[233] ),
    .S(net501),
    .X(_0274_));
 sg13g2_mux2_1 _3176_ (.A0(net781),
    .A1(\load_weights[234] ),
    .S(net501),
    .X(_0275_));
 sg13g2_mux2_1 _3177_ (.A0(net670),
    .A1(\load_weights[235] ),
    .S(net492),
    .X(_0276_));
 sg13g2_mux2_1 _3178_ (.A0(net641),
    .A1(\load_weights[236] ),
    .S(net496),
    .X(_0277_));
 sg13g2_mux2_1 _3179_ (.A0(net596),
    .A1(\load_weights[237] ),
    .S(net499),
    .X(_0278_));
 sg13g2_nor2_1 _3180_ (.A(net496),
    .B(net568),
    .Y(_1875_));
 sg13g2_a21oi_1 _3181_ (.A1(net496),
    .A2(_1930_),
    .Y(_0279_),
    .B1(_1875_));
 sg13g2_mux2_1 _3182_ (.A0(net737),
    .A1(net788),
    .S(net492),
    .X(_0280_));
 sg13g2_mux2_1 _3183_ (.A0(net814),
    .A1(net812),
    .S(net501),
    .X(_0281_));
 sg13g2_mux2_1 _3184_ (.A0(net673),
    .A1(net602),
    .S(net497),
    .X(_0282_));
 sg13g2_mux2_1 _3185_ (.A0(net741),
    .A1(net635),
    .S(net501),
    .X(_0283_));
 sg13g2_mux2_1 _3186_ (.A0(\load_weights[255] ),
    .A1(net598),
    .S(net496),
    .X(_0284_));
 sg13g2_nand2_1 _3187_ (.Y(_1876_),
    .A(net502),
    .B(net581));
 sg13g2_o21ai_1 _3188_ (.B1(_1876_),
    .Y(_0285_),
    .A1(net502),
    .A2(_1928_));
 sg13g2_mux2_1 _3189_ (.A0(net752),
    .A1(net730),
    .S(net501),
    .X(_0286_));
 sg13g2_mux2_1 _3190_ (.A0(net794),
    .A1(net781),
    .S(net496),
    .X(_0287_));
 sg13g2_mux2_1 _3191_ (.A0(net726),
    .A1(net670),
    .S(net496),
    .X(_0288_));
 sg13g2_mux2_1 _3192_ (.A0(net699),
    .A1(net641),
    .S(net497),
    .X(_0289_));
 sg13g2_mux2_1 _3193_ (.A0(net694),
    .A1(net596),
    .S(net502),
    .X(_0290_));
 sg13g2_nand2_1 _3194_ (.Y(_1877_),
    .A(net497),
    .B(net568));
 sg13g2_o21ai_1 _3195_ (.B1(_1877_),
    .Y(_0291_),
    .A1(net497),
    .A2(_1927_));
 sg13g2_mux2_1 _3196_ (.A0(\load_weights[263] ),
    .A1(net737),
    .S(net496),
    .X(_0292_));
 sg13g2_mux2_1 _3197_ (.A0(net801),
    .A1(\load_weights[252] ),
    .S(net495),
    .X(_0293_));
 sg13g2_mux2_1 _3198_ (.A0(net821),
    .A1(net673),
    .S(net495),
    .X(_0294_));
 sg13g2_mux2_1 _3199_ (.A0(net900),
    .A1(net741),
    .S(net494),
    .X(_0295_));
 sg13g2_mux2_1 _3200_ (.A0(net880),
    .A1(\load_weights[255] ),
    .S(net498),
    .X(_0296_));
 sg13g2_nor2_1 _3201_ (.A(net497),
    .B(net816),
    .Y(_1878_));
 sg13g2_a21oi_1 _3202_ (.A1(net497),
    .A2(_1928_),
    .Y(_0297_),
    .B1(_1878_));
 sg13g2_mux2_1 _3203_ (.A0(net623),
    .A1(\load_weights[257] ),
    .S(net495),
    .X(_0298_));
 sg13g2_mux2_1 _3204_ (.A0(net894),
    .A1(net794),
    .S(net498),
    .X(_0299_));
 sg13g2_mux2_1 _3205_ (.A0(net657),
    .A1(\load_weights[259] ),
    .S(net495),
    .X(_0300_));
 sg13g2_mux2_1 _3206_ (.A0(net874),
    .A1(net699),
    .S(net494),
    .X(_0301_));
 sg13g2_mux2_1 _3207_ (.A0(net740),
    .A1(net694),
    .S(net495),
    .X(_0302_));
 sg13g2_nor2_1 _3208_ (.A(net494),
    .B(net765),
    .Y(_1879_));
 sg13g2_a21oi_1 _3209_ (.A1(net494),
    .A2(_1927_),
    .Y(_0303_),
    .B1(_1879_));
 sg13g2_mux2_1 _3210_ (.A0(net776),
    .A1(\load_weights[263] ),
    .S(net495),
    .X(_0304_));
 sg13g2_mux2_1 _3211_ (.A0(net840),
    .A1(net801),
    .S(net472),
    .X(_0305_));
 sg13g2_mux2_1 _3212_ (.A0(net845),
    .A1(net821),
    .S(net472),
    .X(_0306_));
 sg13g2_mux2_1 _3213_ (.A0(net901),
    .A1(net900),
    .S(net473),
    .X(_0307_));
 sg13g2_mux2_1 _3214_ (.A0(net897),
    .A1(net880),
    .S(net473),
    .X(_0308_));
 sg13g2_nand2_1 _3215_ (.Y(_1880_),
    .A(net472),
    .B(net816));
 sg13g2_o21ai_1 _3216_ (.B1(_1880_),
    .Y(_0309_),
    .A1(net473),
    .A2(_1934_));
 sg13g2_mux2_1 _3217_ (.A0(net679),
    .A1(net623),
    .S(net494),
    .X(_0310_));
 sg13g2_mux2_1 _3218_ (.A0(\load_weights[282] ),
    .A1(net894),
    .S(net473),
    .X(_0311_));
 sg13g2_mux2_1 _3219_ (.A0(net693),
    .A1(net657),
    .S(net495),
    .X(_0312_));
 sg13g2_mux2_1 _3220_ (.A0(net889),
    .A1(net874),
    .S(net494),
    .X(_0313_));
 sg13g2_mux2_1 _3221_ (.A0(net751),
    .A1(net740),
    .S(net495),
    .X(_0314_));
 sg13g2_nand2_1 _3222_ (.Y(_1881_),
    .A(net494),
    .B(net765));
 sg13g2_o21ai_1 _3223_ (.B1(_1881_),
    .Y(_0315_),
    .A1(net494),
    .A2(_1933_));
 sg13g2_mux2_1 _3224_ (.A0(net795),
    .A1(net776),
    .S(net472),
    .X(_0316_));
 sg13g2_nor4_1 _3225_ (.A(net519),
    .B(net524),
    .C(net509),
    .D(net514),
    .Y(_1882_));
 sg13g2_nor4_2 _3226_ (.A(net538),
    .B(net542),
    .C(net529),
    .Y(_1883_),
    .D(net533));
 sg13g2_nor4_1 _3227_ (.A(net556),
    .B(net561),
    .C(net547),
    .D(net551),
    .Y(_1884_));
 sg13g2_nand3_1 _3228_ (.B(_1883_),
    .C(_1884_),
    .A(_1882_),
    .Y(_1885_));
 sg13g2_nor2b_1 _3229_ (.A(net892),
    .B_N(_1885_),
    .Y(_1886_));
 sg13g2_nand3b_1 _3230_ (.B(_1886_),
    .C(net1),
    .Y(_1887_),
    .A_N(net502));
 sg13g2_nor2_1 _3231_ (.A(net561),
    .B(_1887_),
    .Y(_1888_));
 sg13g2_a21oi_1 _3232_ (.A1(_1924_),
    .A2(net421),
    .Y(_0317_),
    .B1(_1888_));
 sg13g2_nor2_1 _3233_ (.A(net556),
    .B(_1887_),
    .Y(_1889_));
 sg13g2_a21oi_1 _3234_ (.A1(_1925_),
    .A2(net421),
    .Y(_0318_),
    .B1(_1889_));
 sg13g2_nor2_1 _3235_ (.A(net551),
    .B(_1887_),
    .Y(_1890_));
 sg13g2_a21oi_1 _3236_ (.A1(_1926_),
    .A2(net421),
    .Y(_0319_),
    .B1(_1890_));
 sg13g2_mux2_1 _3237_ (.A0(net547),
    .A1(net807),
    .S(net421),
    .X(_0320_));
 sg13g2_mux2_1 _3238_ (.A0(net542),
    .A1(net843),
    .S(net421),
    .X(_0321_));
 sg13g2_mux2_1 _3239_ (.A0(net537),
    .A1(net856),
    .S(net421),
    .X(_0322_));
 sg13g2_mux2_1 _3240_ (.A0(net533),
    .A1(net760),
    .S(net421),
    .X(_0323_));
 sg13g2_mux2_1 _3241_ (.A0(net528),
    .A1(net667),
    .S(net421),
    .X(_0324_));
 sg13g2_and3_1 _3242_ (.X(_1891_),
    .A(\count[1] ),
    .B(\count[0] ),
    .C(net831));
 sg13g2_and4_1 _3243_ (.A(net502),
    .B(net917),
    .C(_1989_),
    .D(_1891_),
    .X(_1892_));
 sg13g2_o21ai_1 _3244_ (.B1(net1),
    .Y(_1893_),
    .A1(net892),
    .A2(_1892_));
 sg13g2_inv_1 _3245_ (.Y(_0325_),
    .A(net893));
 sg13g2_nor2_1 _3246_ (.A(net502),
    .B(_1886_),
    .Y(_1894_));
 sg13g2_nor3_1 _3247_ (.A(_1922_),
    .B(_1892_),
    .C(_1894_),
    .Y(_0326_));
 sg13g2_nand2b_1 _3248_ (.Y(_1895_),
    .B(\bit_select[0] ),
    .A_N(\count[0] ));
 sg13g2_xnor2_1 _3249_ (.Y(_1896_),
    .A(\count[3] ),
    .B(\bit_select[3] ));
 sg13g2_nor2_1 _3250_ (.A(_1923_),
    .B(\bit_select[4] ),
    .Y(_1897_));
 sg13g2_nor2_1 _3251_ (.A(\count[1] ),
    .B(_1925_),
    .Y(_1898_));
 sg13g2_xnor2_1 _3252_ (.Y(_1899_),
    .A(\count[7] ),
    .B(\bit_select[7] ));
 sg13g2_nor2_1 _3253_ (.A(\count[2] ),
    .B(_1926_),
    .Y(_1900_));
 sg13g2_a22oi_1 _3254_ (.Y(_1901_),
    .B1(_1926_),
    .B2(\count[2] ),
    .A2(_1924_),
    .A1(\count[0] ));
 sg13g2_a22oi_1 _3255_ (.Y(_1902_),
    .B1(\bit_select[4] ),
    .B2(_1923_),
    .A2(_1925_),
    .A1(\count[1] ));
 sg13g2_xnor2_1 _3256_ (.Y(_1903_),
    .A(\count[5] ),
    .B(\bit_select[5] ));
 sg13g2_xnor2_1 _3257_ (.Y(_1904_),
    .A(\count[6] ),
    .B(\bit_select[6] ));
 sg13g2_nand4_1 _3258_ (.B(_1902_),
    .C(_1903_),
    .A(_1896_),
    .Y(_1905_),
    .D(_1904_));
 sg13g2_nor4_1 _3259_ (.A(_1897_),
    .B(_1898_),
    .C(_1900_),
    .D(_1905_),
    .Y(_1906_));
 sg13g2_nand4_1 _3260_ (.B(_1899_),
    .C(_1901_),
    .A(_1895_),
    .Y(_1907_),
    .D(_1906_));
 sg13g2_a21oi_1 _3261_ (.A1(net892),
    .A2(_1907_),
    .Y(_1908_),
    .B1(net502));
 sg13g2_nand2b_2 _3262_ (.Y(_1909_),
    .B(net1),
    .A_N(_1908_));
 sg13g2_nor2_1 _3263_ (.A(net864),
    .B(_1909_),
    .Y(_0327_));
 sg13g2_xnor2_1 _3264_ (.Y(_1910_),
    .A(net908),
    .B(net864));
 sg13g2_nor2_1 _3265_ (.A(_1909_),
    .B(_1910_),
    .Y(_0328_));
 sg13g2_a21oi_1 _3266_ (.A1(\count[1] ),
    .A2(\count[0] ),
    .Y(_1911_),
    .B1(net831));
 sg13g2_nor3_1 _3267_ (.A(_1891_),
    .B(_1909_),
    .C(net832),
    .Y(_0329_));
 sg13g2_or2_1 _3268_ (.X(_1912_),
    .B(_1909_),
    .A(_1892_));
 sg13g2_and2_1 _3269_ (.A(net883),
    .B(_1891_),
    .X(_1913_));
 sg13g2_nor2_1 _3270_ (.A(net883),
    .B(_1891_),
    .Y(_1914_));
 sg13g2_nor3_1 _3271_ (.A(_1912_),
    .B(_1913_),
    .C(net884),
    .Y(_0330_));
 sg13g2_and2_1 _3272_ (.A(net877),
    .B(_1913_),
    .X(_1915_));
 sg13g2_nor2_1 _3273_ (.A(net877),
    .B(_1913_),
    .Y(_1916_));
 sg13g2_nor3_1 _3274_ (.A(_1912_),
    .B(_1915_),
    .C(net878),
    .Y(_0331_));
 sg13g2_and2_1 _3275_ (.A(net871),
    .B(_1915_),
    .X(_1917_));
 sg13g2_nor2_1 _3276_ (.A(net871),
    .B(_1915_),
    .Y(_1918_));
 sg13g2_nor3_1 _3277_ (.A(_1909_),
    .B(_1917_),
    .C(net872),
    .Y(_0332_));
 sg13g2_nand2_1 _3278_ (.Y(_1919_),
    .A(net904),
    .B(_1917_));
 sg13g2_xnor2_1 _3279_ (.Y(_1920_),
    .A(net904),
    .B(_1917_));
 sg13g2_nor2_1 _3280_ (.A(_1909_),
    .B(_1920_),
    .Y(_0333_));
 sg13g2_xor2_1 _3281_ (.B(_1919_),
    .A(net912),
    .X(_1921_));
 sg13g2_nor2_1 _3282_ (.A(_1909_),
    .B(_1921_),
    .Y(_0334_));
 sg13g2_inv_1 _3283_ (.Y(_1922_),
    .A(net1));
 sg13g2_inv_1 _3284_ (.Y(_1923_),
    .A(\count[4] ));
 sg13g2_inv_1 _3285_ (.Y(_1924_),
    .A(net403));
 sg13g2_inv_1 _3286_ (.Y(_1925_),
    .A(net575));
 sg13g2_inv_1 _3287_ (.Y(_1926_),
    .A(net706));
 sg13g2_inv_1 _3288_ (.Y(_1927_),
    .A(net875));
 sg13g2_inv_2 _3289_ (.Y(_1928_),
    .A(\load_weights[256] ));
 sg13g2_inv_1 _3290_ (.Y(_1929_),
    .A(_0022_));
 sg13g2_inv_1 _3291_ (.Y(_1930_),
    .A(net686));
 sg13g2_inv_1 _3292_ (.Y(_1931_),
    .A(net609));
 sg13g2_inv_1 _3293_ (.Y(_1932_),
    .A(_0024_));
 sg13g2_inv_1 _3294_ (.Y(_1933_),
    .A(\load_weights[286] ));
 sg13g2_inv_1 _3295_ (.Y(_1934_),
    .A(net866));
 sg13g2_inv_1 _3296_ (.Y(_1935_),
    .A(_0026_));
 sg13g2_inv_1 _3297_ (.Y(_1936_),
    .A(net637));
 sg13g2_inv_2 _3298_ (.Y(_1937_),
    .A(net722));
 sg13g2_inv_1 _3299_ (.Y(_1938_),
    .A(_0028_));
 sg13g2_inv_1 _3300_ (.Y(_1939_),
    .A(net412));
 sg13g2_inv_1 _3301_ (.Y(_1940_),
    .A(net768));
 sg13g2_inv_1 _3302_ (.Y(_1941_),
    .A(_0001_));
 sg13g2_inv_1 _3303_ (.Y(_1942_),
    .A(net414));
 sg13g2_inv_1 _3304_ (.Y(_1943_),
    .A(\load_weights[87] ));
 sg13g2_inv_1 _3305_ (.Y(_1944_),
    .A(_0003_));
 sg13g2_inv_1 _3306_ (.Y(_1945_),
    .A(net578));
 sg13g2_inv_2 _3307_ (.Y(_1946_),
    .A(net574));
 sg13g2_inv_2 _3308_ (.Y(_1947_),
    .A(net400));
 sg13g2_inv_1 _3309_ (.Y(_1948_),
    .A(net665));
 sg13g2_inv_2 _3310_ (.Y(_1949_),
    .A(\load_weights[43] ));
 sg13g2_inv_2 _3311_ (.Y(_1950_),
    .A(\load_weights[41] ));
 sg13g2_inv_1 _3312_ (.Y(_1951_),
    .A(net870));
 sg13g2_inv_1 _3313_ (.Y(_1952_),
    .A(\load_weights[139] ));
 sg13g2_inv_1 _3314_ (.Y(_1953_),
    .A(net728));
 sg13g2_inv_1 _3315_ (.Y(_1954_),
    .A(net735));
 sg13g2_inv_1 _3316_ (.Y(_1955_),
    .A(net407));
 sg13g2_inv_1 _3317_ (.Y(_1956_),
    .A(\load_weights[16] ));
 sg13g2_inv_1 _3318_ (.Y(_1957_),
    .A(\load_weights[22] ));
 sg13g2_inv_1 _3319_ (.Y(_1958_),
    .A(_0015_));
 sg13g2_inv_2 _3320_ (.Y(_1959_),
    .A(\load_weights[190] ));
 sg13g2_inv_2 _3321_ (.Y(_1960_),
    .A(net857));
 sg13g2_inv_1 _3322_ (.Y(_1961_),
    .A(_0017_));
 sg13g2_inv_1 _3323_ (.Y(_1962_),
    .A(net709));
 sg13g2_inv_1 _3324_ (.Y(_1963_),
    .A(net652));
 sg13g2_inv_1 _3325_ (.Y(_1964_),
    .A(_0019_));
 sg13g2_a21oi_1 _3326_ (.A1(net551),
    .A2(\load_weights[246] ),
    .Y(_1965_),
    .B1(\load_weights[258] ));
 sg13g2_a21o_1 _3327_ (.A2(\load_weights[258] ),
    .A1(net550),
    .B1(_1965_),
    .X(_1966_));
 sg13g2_a21oi_1 _3328_ (.A1(net510),
    .A2(\load_weights[243] ),
    .Y(_1967_),
    .B1(\load_weights[255] ));
 sg13g2_a21o_1 _3329_ (.A2(\load_weights[255] ),
    .A1(net510),
    .B1(_1967_),
    .X(_1968_));
 sg13g2_xor2_1 _3330_ (.B(_1968_),
    .A(_1966_),
    .X(_1969_));
 sg13g2_a21oi_1 _3331_ (.A1(net518),
    .A2(\load_weights[241] ),
    .Y(_1970_),
    .B1(\load_weights[253] ));
 sg13g2_a21oi_1 _3332_ (.A1(net518),
    .A2(\load_weights[253] ),
    .Y(_1971_),
    .B1(_1970_));
 sg13g2_nand2_1 _3333_ (.Y(_1972_),
    .A(_1969_),
    .B(_1971_));
 sg13g2_xnor2_1 _3334_ (.Y(_1973_),
    .A(_1969_),
    .B(_1971_));
 sg13g2_inv_1 _3335_ (.Y(_1974_),
    .A(_1973_));
 sg13g2_a21oi_1 _3336_ (.A1(net528),
    .A2(\load_weights[251] ),
    .Y(_1975_),
    .B1(\load_weights[263] ));
 sg13g2_a21o_1 _3337_ (.A2(\load_weights[263] ),
    .A1(net528),
    .B1(_1975_),
    .X(_1976_));
 sg13g2_a21oi_1 _3338_ (.A1(net533),
    .A2(\load_weights[250] ),
    .Y(_1977_),
    .B1(\load_weights[262] ));
 sg13g2_a21o_1 _3339_ (.A2(\load_weights[262] ),
    .A1(net533),
    .B1(_1977_),
    .X(_1978_));
 sg13g2_xor2_1 _3340_ (.B(_1978_),
    .A(_1976_),
    .X(_1979_));
 sg13g2_a21oi_1 _3341_ (.A1(net542),
    .A2(\load_weights[248] ),
    .Y(_1980_),
    .B1(\load_weights[260] ));
 sg13g2_a21o_1 _3342_ (.A2(\load_weights[260] ),
    .A1(net541),
    .B1(_1980_),
    .X(_1981_));
 sg13g2_inv_1 _3343_ (.Y(_1982_),
    .A(_1981_));
 sg13g2_nand2_1 _3344_ (.Y(_1983_),
    .A(_1979_),
    .B(_1982_));
 sg13g2_nand2b_1 _3345_ (.Y(_1984_),
    .B(_1981_),
    .A_N(_1979_));
 sg13g2_nand2_1 _3346_ (.Y(_1985_),
    .A(_1979_),
    .B(_1981_));
 sg13g2_nand2b_1 _3347_ (.Y(_1986_),
    .B(_1982_),
    .A_N(_1979_));
 sg13g2_nand2_1 _3348_ (.Y(_1987_),
    .A(_1983_),
    .B(_1984_));
 sg13g2_inv_1 _3349_ (.Y(_1988_),
    .A(_1987_));
 sg13g2_nor4_2 _3350_ (.A(\count[3] ),
    .B(\count[5] ),
    .C(\count[7] ),
    .Y(_1989_),
    .D(\count[6] ));
 sg13g2_nor4_2 _3351_ (.A(\count[1] ),
    .B(\count[0] ),
    .C(\count[2] ),
    .Y(_1990_),
    .D(\count[4] ));
 sg13g2_and2_2 _3352_ (.A(_1989_),
    .B(_1990_),
    .X(_1991_));
 sg13g2_nand2_2 _3353_ (.Y(_1992_),
    .A(_1989_),
    .B(_1990_));
 sg13g2_nand2_1 _3354_ (.Y(_1993_),
    .A(\load_weights[252] ),
    .B(\load_weights[253] ));
 sg13g2_xnor2_1 _3355_ (.Y(_1994_),
    .A(\load_weights[252] ),
    .B(\load_weights[253] ));
 sg13g2_and2_1 _3356_ (.A(\load_weights[254] ),
    .B(\load_weights[255] ),
    .X(_1995_));
 sg13g2_xor2_1 _3357_ (.B(\load_weights[255] ),
    .A(\load_weights[254] ),
    .X(_1996_));
 sg13g2_xnor2_1 _3358_ (.Y(_1997_),
    .A(\load_weights[257] ),
    .B(_1996_));
 sg13g2_nor2_1 _3359_ (.A(_1994_),
    .B(_1997_),
    .Y(_1998_));
 sg13g2_xnor2_1 _3360_ (.Y(_1999_),
    .A(_1994_),
    .B(_1997_));
 sg13g2_and2_1 _3361_ (.A(\load_weights[259] ),
    .B(\load_weights[261] ),
    .X(_2000_));
 sg13g2_xor2_1 _3362_ (.B(\load_weights[261] ),
    .A(\load_weights[259] ),
    .X(_2001_));
 sg13g2_xnor2_1 _3363_ (.Y(_2002_),
    .A(\load_weights[263] ),
    .B(_2001_));
 sg13g2_nor2_1 _3364_ (.A(_1999_),
    .B(_2002_),
    .Y(_2003_));
 sg13g2_xor2_1 _3365_ (.B(_2002_),
    .A(_1999_),
    .X(_2004_));
 sg13g2_nand2_1 _3366_ (.Y(_2005_),
    .A(\load_weights[260] ),
    .B(_2004_));
 sg13g2_xnor2_1 _3367_ (.Y(_2006_),
    .A(\load_weights[260] ),
    .B(_2004_));
 sg13g2_xnor2_1 _3368_ (.Y(_2007_),
    .A(\load_weights[262] ),
    .B(_2006_));
 sg13g2_nand2_1 _3369_ (.Y(_2008_),
    .A(\load_weights[258] ),
    .B(_2007_));
 sg13g2_xor2_1 _3370_ (.B(_2007_),
    .A(\load_weights[258] ),
    .X(_2009_));
 sg13g2_xnor2_1 _3371_ (.Y(_2010_),
    .A(\load_weights[258] ),
    .B(_2007_));
 sg13g2_nand2_1 _3372_ (.Y(_2011_),
    .A(\load_weights[256] ),
    .B(_2009_));
 sg13g2_a21oi_1 _3373_ (.A1(_1928_),
    .A2(_2010_),
    .Y(_2012_),
    .B1(net433));
 sg13g2_xnor2_1 _3374_ (.Y(_2013_),
    .A(\load_weights[256] ),
    .B(_2009_));
 sg13g2_nor2_1 _3375_ (.A(_1929_),
    .B(net442),
    .Y(_2014_));
 sg13g2_a221oi_1 _3376_ (.B2(_2013_),
    .C1(_2014_),
    .B1(net442),
    .A1(_1985_),
    .Y(_2015_),
    .A2(_1986_));
 sg13g2_a221oi_1 _3377_ (.B2(_2012_),
    .C1(_1988_),
    .B1(_2011_),
    .A1(_1929_),
    .Y(_2016_),
    .A2(net433));
 sg13g2_a221oi_1 _3378_ (.B2(_2012_),
    .C1(_1987_),
    .B1(_2011_),
    .A1(_1929_),
    .Y(_2017_),
    .A2(net432));
 sg13g2_a221oi_1 _3379_ (.B2(_2013_),
    .C1(_2014_),
    .B1(net441),
    .A1(_1983_),
    .Y(_2018_),
    .A2(_1984_));
 sg13g2_nor3_1 _3380_ (.A(_1973_),
    .B(_2015_),
    .C(_2016_),
    .Y(_2019_));
 sg13g2_o21ai_1 _3381_ (.B1(_1974_),
    .Y(_2020_),
    .A1(_2017_),
    .A2(_2018_));
 sg13g2_nor3_1 _3382_ (.A(_1974_),
    .B(_2017_),
    .C(_2018_),
    .Y(_2021_));
 sg13g2_o21ai_1 _3383_ (.B1(_1973_),
    .Y(_2022_),
    .A1(_2015_),
    .A2(_2016_));
 sg13g2_a21oi_1 _3384_ (.A1(net514),
    .A2(\load_weights[242] ),
    .Y(_2023_),
    .B1(\load_weights[254] ));
 sg13g2_a21oi_1 _3385_ (.A1(net514),
    .A2(\load_weights[254] ),
    .Y(_2024_),
    .B1(_2023_));
 sg13g2_a21o_1 _3386_ (.A2(\load_weights[254] ),
    .A1(net514),
    .B1(_2023_),
    .X(_2025_));
 sg13g2_nor3_1 _3387_ (.A(_2019_),
    .B(_2021_),
    .C(_2025_),
    .Y(_2026_));
 sg13g2_nand3_1 _3388_ (.B(_2022_),
    .C(_2024_),
    .A(_2020_),
    .Y(_2027_));
 sg13g2_a21oi_1 _3389_ (.A1(_2020_),
    .A2(_2022_),
    .Y(_2028_),
    .B1(_2024_));
 sg13g2_o21ai_1 _3390_ (.B1(_2025_),
    .Y(_2029_),
    .A1(_2019_),
    .A2(_2021_));
 sg13g2_a21oi_1 _3391_ (.A1(net523),
    .A2(\load_weights[240] ),
    .Y(_2030_),
    .B1(\load_weights[252] ));
 sg13g2_a21oi_1 _3392_ (.A1(net524),
    .A2(\load_weights[252] ),
    .Y(_2031_),
    .B1(_2030_));
 sg13g2_a21o_1 _3393_ (.A2(\load_weights[252] ),
    .A1(net523),
    .B1(_2030_),
    .X(_2032_));
 sg13g2_nor3_1 _3394_ (.A(_2026_),
    .B(_2028_),
    .C(_2032_),
    .Y(_2033_));
 sg13g2_nand3_1 _3395_ (.B(_2029_),
    .C(_2031_),
    .A(_2027_),
    .Y(_2034_));
 sg13g2_a21oi_1 _3396_ (.A1(_2027_),
    .A2(_2029_),
    .Y(_2035_),
    .B1(_2031_));
 sg13g2_o21ai_1 _3397_ (.B1(_2032_),
    .Y(_2036_),
    .A1(_2026_),
    .A2(_2028_));
 sg13g2_a21oi_1 _3398_ (.A1(net556),
    .A2(\load_weights[245] ),
    .Y(_2037_),
    .B1(\load_weights[257] ));
 sg13g2_a21oi_1 _3399_ (.A1(net555),
    .A2(\load_weights[257] ),
    .Y(_2038_),
    .B1(_2037_));
 sg13g2_a21o_1 _3400_ (.A2(\load_weights[257] ),
    .A1(net555),
    .B1(_2037_),
    .X(_2039_));
 sg13g2_nor3_1 _3401_ (.A(_2033_),
    .B(_2035_),
    .C(_2039_),
    .Y(_2040_));
 sg13g2_nand3_1 _3402_ (.B(_2036_),
    .C(_2038_),
    .A(_2034_),
    .Y(_2041_));
 sg13g2_a21oi_1 _3403_ (.A1(_2034_),
    .A2(_2036_),
    .Y(_2042_),
    .B1(_2038_));
 sg13g2_o21ai_1 _3404_ (.B1(_2039_),
    .Y(_2043_),
    .A1(_2033_),
    .A2(_2035_));
 sg13g2_a21oi_1 _3405_ (.A1(net561),
    .A2(\load_weights[244] ),
    .Y(_2044_),
    .B1(\load_weights[256] ));
 sg13g2_a21o_1 _3406_ (.A2(\load_weights[256] ),
    .A1(net561),
    .B1(_2044_),
    .X(_2045_));
 sg13g2_inv_1 _3407_ (.Y(_2046_),
    .A(_2045_));
 sg13g2_nor3_1 _3408_ (.A(_2040_),
    .B(_2042_),
    .C(_2045_),
    .Y(_2047_));
 sg13g2_a21oi_1 _3409_ (.A1(_2041_),
    .A2(_2043_),
    .Y(_2048_),
    .B1(_2046_));
 sg13g2_nand3_1 _3410_ (.B(_2043_),
    .C(_2045_),
    .A(_2041_),
    .Y(_2049_));
 sg13g2_o21ai_1 _3411_ (.B1(_2046_),
    .Y(_2050_),
    .A1(_2040_),
    .A2(_2042_));
 sg13g2_a21oi_1 _3412_ (.A1(net546),
    .A2(\load_weights[247] ),
    .Y(_2051_),
    .B1(\load_weights[259] ));
 sg13g2_a21o_1 _3413_ (.A2(\load_weights[259] ),
    .A1(net547),
    .B1(_2051_),
    .X(_2052_));
 sg13g2_nor3_1 _3414_ (.A(_2047_),
    .B(_2048_),
    .C(_2052_),
    .Y(_2053_));
 sg13g2_and3_1 _3415_ (.X(_2054_),
    .A(_2049_),
    .B(_2050_),
    .C(_2052_));
 sg13g2_o21ai_1 _3416_ (.B1(_2052_),
    .Y(_2055_),
    .A1(_2047_),
    .A2(_2048_));
 sg13g2_a21oi_1 _3417_ (.A1(net537),
    .A2(net596),
    .Y(_2056_),
    .B1(\load_weights[261] ));
 sg13g2_a21oi_1 _3418_ (.A1(net537),
    .A2(\load_weights[261] ),
    .Y(_2057_),
    .B1(_2056_));
 sg13g2_nor3_1 _3419_ (.A(_2053_),
    .B(_2054_),
    .C(_2057_),
    .Y(_2058_));
 sg13g2_o21ai_1 _3420_ (.B1(_2057_),
    .Y(_2059_),
    .A1(_2053_),
    .A2(_2054_));
 sg13g2_nand2b_1 _3421_ (.Y(\tt_um_mult_inst.genblk1[10].out_q ),
    .B(_2059_),
    .A_N(_2058_));
 sg13g2_a21oi_1 _3422_ (.A1(_2055_),
    .A2(_2057_),
    .Y(_2060_),
    .B1(_2053_));
 sg13g2_o21ai_1 _3423_ (.B1(_1972_),
    .Y(_2061_),
    .A1(_1966_),
    .A2(_1968_));
 sg13g2_nand2b_1 _3424_ (.Y(_2062_),
    .B(_2020_),
    .A_N(_2015_));
 sg13g2_o21ai_1 _3425_ (.B1(_1983_),
    .Y(_2063_),
    .A1(_1976_),
    .A2(_1978_));
 sg13g2_nor2_1 _3426_ (.A(\tt_um_mult_inst.genblk1[10].carry[1] ),
    .B(net441),
    .Y(_2064_));
 sg13g2_nand2_1 _3427_ (.Y(_2065_),
    .A(_2008_),
    .B(_2011_));
 sg13g2_a21oi_1 _3428_ (.A1(\load_weights[263] ),
    .A2(_2001_),
    .Y(_2066_),
    .B1(_2000_));
 sg13g2_a21oi_1 _3429_ (.A1(\load_weights[257] ),
    .A2(_1996_),
    .Y(_2067_),
    .B1(_1995_));
 sg13g2_nor2_1 _3430_ (.A(_1993_),
    .B(_2067_),
    .Y(_2068_));
 sg13g2_xnor2_1 _3431_ (.Y(_2069_),
    .A(_1993_),
    .B(_2067_));
 sg13g2_nor2_1 _3432_ (.A(_1998_),
    .B(_2003_),
    .Y(_2070_));
 sg13g2_nor2_1 _3433_ (.A(_2069_),
    .B(_2070_),
    .Y(_2071_));
 sg13g2_xnor2_1 _3434_ (.Y(_2072_),
    .A(_2069_),
    .B(_2070_));
 sg13g2_nor2_1 _3435_ (.A(_2066_),
    .B(_2072_),
    .Y(_2073_));
 sg13g2_xor2_1 _3436_ (.B(_2072_),
    .A(_2066_),
    .X(_2074_));
 sg13g2_o21ai_1 _3437_ (.B1(_2005_),
    .Y(_2075_),
    .A1(_1927_),
    .A2(_2006_));
 sg13g2_and2_1 _3438_ (.A(_2074_),
    .B(_2075_),
    .X(_2076_));
 sg13g2_xor2_1 _3439_ (.B(_2075_),
    .A(_2074_),
    .X(_2077_));
 sg13g2_xnor2_1 _3440_ (.Y(_2078_),
    .A(_2065_),
    .B(_2077_));
 sg13g2_a21oi_1 _3441_ (.A1(net441),
    .A2(_2078_),
    .Y(_2079_),
    .B1(_2064_));
 sg13g2_nand2_1 _3442_ (.Y(_2080_),
    .A(_2063_),
    .B(_2079_));
 sg13g2_xor2_1 _3443_ (.B(_2079_),
    .A(_2063_),
    .X(_2081_));
 sg13g2_nand2_1 _3444_ (.Y(_2082_),
    .A(_2062_),
    .B(_2081_));
 sg13g2_xnor2_1 _3445_ (.Y(_2083_),
    .A(_2062_),
    .B(_2081_));
 sg13g2_nand2b_1 _3446_ (.Y(_2084_),
    .B(_2061_),
    .A_N(_2083_));
 sg13g2_xor2_1 _3447_ (.B(_2083_),
    .A(_2061_),
    .X(_2085_));
 sg13g2_nand2_1 _3448_ (.Y(_2086_),
    .A(_2027_),
    .B(_2034_));
 sg13g2_nand2b_1 _3449_ (.Y(_2087_),
    .B(_2086_),
    .A_N(_2085_));
 sg13g2_xnor2_1 _3450_ (.Y(_2088_),
    .A(_2085_),
    .B(_2086_));
 sg13g2_o21ai_1 _3451_ (.B1(_2041_),
    .Y(_2089_),
    .A1(_2042_),
    .A2(_2045_));
 sg13g2_nand2_1 _3452_ (.Y(_2090_),
    .A(_2088_),
    .B(_2089_));
 sg13g2_xnor2_1 _3453_ (.Y(_2091_),
    .A(_2088_),
    .B(_2089_));
 sg13g2_xor2_1 _3454_ (.B(_2091_),
    .A(_2060_),
    .X(\tt_um_mult_inst.genblk1[10].carry_q[0] ));
 sg13g2_o21ai_1 _3455_ (.B1(_2090_),
    .Y(_2092_),
    .A1(_2060_),
    .A2(_2091_));
 sg13g2_nand2_1 _3456_ (.Y(_2093_),
    .A(_2068_),
    .B(_2073_));
 sg13g2_nor3_1 _3457_ (.A(_2068_),
    .B(_2071_),
    .C(_2073_),
    .Y(_2094_));
 sg13g2_a21oi_1 _3458_ (.A1(_2068_),
    .A2(_2073_),
    .Y(_2095_),
    .B1(_2094_));
 sg13g2_a21o_1 _3459_ (.A2(_2077_),
    .A1(_2065_),
    .B1(_2076_),
    .X(_2096_));
 sg13g2_or2_1 _3460_ (.X(_2097_),
    .B(_2096_),
    .A(_2095_));
 sg13g2_a21oi_1 _3461_ (.A1(_2095_),
    .A2(_2096_),
    .Y(_2098_),
    .B1(net433));
 sg13g2_a22oi_1 _3462_ (.Y(_2099_),
    .B1(_2097_),
    .B2(_2098_),
    .A2(net432),
    .A1(\tt_um_mult_inst.genblk1[10].carry[2] ));
 sg13g2_nor2_1 _3463_ (.A(_2080_),
    .B(_2099_),
    .Y(_2100_));
 sg13g2_xnor2_1 _3464_ (.Y(_2101_),
    .A(_2080_),
    .B(_2099_));
 sg13g2_a21o_1 _3465_ (.A2(_2084_),
    .A1(_2082_),
    .B1(_2101_),
    .X(_2102_));
 sg13g2_nand3_1 _3466_ (.B(_2084_),
    .C(_2101_),
    .A(_2082_),
    .Y(_2103_));
 sg13g2_nand2_1 _3467_ (.Y(_2104_),
    .A(_2102_),
    .B(_2103_));
 sg13g2_nor2_1 _3468_ (.A(_2087_),
    .B(_2104_),
    .Y(_2105_));
 sg13g2_xor2_1 _3469_ (.B(_2104_),
    .A(_2087_),
    .X(_2106_));
 sg13g2_xor2_1 _3470_ (.B(_2106_),
    .A(_2092_),
    .X(\tt_um_mult_inst.genblk1[10].carry_q[1] ));
 sg13g2_a22oi_1 _3471_ (.Y(_2107_),
    .B1(_2093_),
    .B2(_2098_),
    .A2(net433),
    .A1(net927));
 sg13g2_xnor2_1 _3472_ (.Y(_2108_),
    .A(_2100_),
    .B(_2107_));
 sg13g2_nor2_1 _3473_ (.A(_2102_),
    .B(_2108_),
    .Y(_2109_));
 sg13g2_xor2_1 _3474_ (.B(_2108_),
    .A(_2102_),
    .X(_2110_));
 sg13g2_a21oi_1 _3475_ (.A1(_2092_),
    .A2(_2106_),
    .Y(_2111_),
    .B1(_2105_));
 sg13g2_nand2b_1 _3476_ (.Y(_2112_),
    .B(_2110_),
    .A_N(_2111_));
 sg13g2_xnor2_1 _3477_ (.Y(\tt_um_mult_inst.genblk1[10].carry_q[2] ),
    .A(_2110_),
    .B(_2111_));
 sg13g2_a21oi_1 _3478_ (.A1(_2100_),
    .A2(_2107_),
    .Y(_2113_),
    .B1(_2109_));
 sg13g2_nand2_1 _3479_ (.Y(\tt_um_mult_inst.genblk1[10].carry_q[3] ),
    .A(_2112_),
    .B(_2113_));
 sg13g2_a21oi_1 _3480_ (.A1(net538),
    .A2(\load_weights[225] ),
    .Y(_2114_),
    .B1(\load_weights[237] ));
 sg13g2_a21o_1 _3481_ (.A2(\load_weights[237] ),
    .A1(net538),
    .B1(_2114_),
    .X(_2115_));
 sg13g2_a21oi_1 _3482_ (.A1(net547),
    .A2(\load_weights[223] ),
    .Y(_2116_),
    .B1(\load_weights[235] ));
 sg13g2_a21o_1 _3483_ (.A2(\load_weights[235] ),
    .A1(net547),
    .B1(_2116_),
    .X(_2117_));
 sg13g2_xor2_1 _3484_ (.B(_2117_),
    .A(_2115_),
    .X(_2118_));
 sg13g2_a21oi_1 _3485_ (.A1(net509),
    .A2(\load_weights[219] ),
    .Y(_2119_),
    .B1(\load_weights[231] ));
 sg13g2_a21oi_2 _3486_ (.B1(_2119_),
    .Y(_2120_),
    .A2(\load_weights[231] ),
    .A1(net509));
 sg13g2_nand2_1 _3487_ (.Y(_2121_),
    .A(_2118_),
    .B(_2120_));
 sg13g2_xnor2_1 _3488_ (.Y(_2122_),
    .A(_2118_),
    .B(_2120_));
 sg13g2_inv_1 _3489_ (.Y(_2123_),
    .A(_2122_));
 sg13g2_a21oi_1 _3490_ (.A1(net551),
    .A2(\load_weights[222] ),
    .Y(_2124_),
    .B1(\load_weights[234] ));
 sg13g2_a21o_1 _3491_ (.A2(\load_weights[234] ),
    .A1(net551),
    .B1(_2124_),
    .X(_2125_));
 sg13g2_a21oi_1 _3492_ (.A1(net513),
    .A2(\load_weights[218] ),
    .Y(_2126_),
    .B1(\load_weights[230] ));
 sg13g2_a21o_1 _3493_ (.A2(\load_weights[230] ),
    .A1(net514),
    .B1(_2126_),
    .X(_2127_));
 sg13g2_xor2_1 _3494_ (.B(_2127_),
    .A(_2125_),
    .X(_2128_));
 sg13g2_a21oi_1 _3495_ (.A1(net529),
    .A2(\load_weights[227] ),
    .Y(_2129_),
    .B1(\load_weights[239] ));
 sg13g2_a21o_1 _3496_ (.A2(\load_weights[239] ),
    .A1(net529),
    .B1(_2129_),
    .X(_2130_));
 sg13g2_inv_1 _3497_ (.Y(_2131_),
    .A(_2130_));
 sg13g2_nand2_1 _3498_ (.Y(_2132_),
    .A(_2128_),
    .B(_2131_));
 sg13g2_nand2b_1 _3499_ (.Y(_2133_),
    .B(_2130_),
    .A_N(_2128_));
 sg13g2_nand2_1 _3500_ (.Y(_2134_),
    .A(_2128_),
    .B(_2130_));
 sg13g2_nand2b_1 _3501_ (.Y(_2135_),
    .B(_2131_),
    .A_N(_2128_));
 sg13g2_nand2_1 _3502_ (.Y(_2136_),
    .A(_2132_),
    .B(_2133_));
 sg13g2_inv_1 _3503_ (.Y(_2137_),
    .A(_2136_));
 sg13g2_nand2_1 _3504_ (.Y(_2138_),
    .A(\load_weights[228] ),
    .B(\load_weights[229] ));
 sg13g2_xnor2_1 _3505_ (.Y(_2139_),
    .A(\load_weights[228] ),
    .B(\load_weights[229] ));
 sg13g2_and2_1 _3506_ (.A(\load_weights[230] ),
    .B(\load_weights[231] ),
    .X(_2140_));
 sg13g2_xor2_1 _3507_ (.B(\load_weights[231] ),
    .A(\load_weights[230] ),
    .X(_2141_));
 sg13g2_xnor2_1 _3508_ (.Y(_2142_),
    .A(\load_weights[233] ),
    .B(_2141_));
 sg13g2_nor2_1 _3509_ (.A(_2139_),
    .B(_2142_),
    .Y(_2143_));
 sg13g2_xnor2_1 _3510_ (.Y(_2144_),
    .A(_2139_),
    .B(_2142_));
 sg13g2_and2_1 _3511_ (.A(\load_weights[235] ),
    .B(\load_weights[237] ),
    .X(_2145_));
 sg13g2_xor2_1 _3512_ (.B(\load_weights[237] ),
    .A(\load_weights[235] ),
    .X(_2146_));
 sg13g2_xnor2_1 _3513_ (.Y(_2147_),
    .A(\load_weights[239] ),
    .B(_2146_));
 sg13g2_nor2_1 _3514_ (.A(_2144_),
    .B(_2147_),
    .Y(_2148_));
 sg13g2_xor2_1 _3515_ (.B(_2147_),
    .A(_2144_),
    .X(_2149_));
 sg13g2_nand2_1 _3516_ (.Y(_2150_),
    .A(\load_weights[236] ),
    .B(_2149_));
 sg13g2_xnor2_1 _3517_ (.Y(_2151_),
    .A(\load_weights[236] ),
    .B(_2149_));
 sg13g2_xnor2_1 _3518_ (.Y(_2152_),
    .A(\load_weights[238] ),
    .B(_2151_));
 sg13g2_nand2_1 _3519_ (.Y(_2153_),
    .A(\load_weights[234] ),
    .B(_2152_));
 sg13g2_xor2_1 _3520_ (.B(_2152_),
    .A(\load_weights[234] ),
    .X(_0335_));
 sg13g2_xnor2_1 _3521_ (.Y(_0336_),
    .A(\load_weights[234] ),
    .B(_2152_));
 sg13g2_nand2_1 _3522_ (.Y(_0337_),
    .A(\load_weights[232] ),
    .B(_0335_));
 sg13g2_a21oi_1 _3523_ (.A1(_1931_),
    .A2(_0336_),
    .Y(_0338_),
    .B1(net432));
 sg13g2_xnor2_1 _3524_ (.Y(_0339_),
    .A(\load_weights[232] ),
    .B(_0335_));
 sg13g2_nor2_1 _3525_ (.A(_1932_),
    .B(net441),
    .Y(_0340_));
 sg13g2_a221oi_1 _3526_ (.B2(net441),
    .C1(_0340_),
    .B1(_0339_),
    .A1(_2134_),
    .Y(_0341_),
    .A2(_2135_));
 sg13g2_a221oi_1 _3527_ (.B2(_0338_),
    .C1(_2137_),
    .B1(_0337_),
    .A1(_1932_),
    .Y(_0342_),
    .A2(net432));
 sg13g2_a221oi_1 _3528_ (.B2(_0338_),
    .C1(_2136_),
    .B1(_0337_),
    .A1(_1932_),
    .Y(_0343_),
    .A2(net432));
 sg13g2_a221oi_1 _3529_ (.B2(net441),
    .C1(_0340_),
    .B1(_0339_),
    .A1(_2132_),
    .Y(_0344_),
    .A2(_2133_));
 sg13g2_nor3_1 _3530_ (.A(_2122_),
    .B(_0341_),
    .C(_0342_),
    .Y(_0345_));
 sg13g2_o21ai_1 _3531_ (.B1(_2123_),
    .Y(_0346_),
    .A1(_0343_),
    .A2(_0344_));
 sg13g2_nor3_1 _3532_ (.A(_2123_),
    .B(_0343_),
    .C(_0344_),
    .Y(_0347_));
 sg13g2_o21ai_1 _3533_ (.B1(_2122_),
    .Y(_0348_),
    .A1(_0341_),
    .A2(_0342_));
 sg13g2_a21oi_1 _3534_ (.A1(net556),
    .A2(\load_weights[221] ),
    .Y(_0349_),
    .B1(\load_weights[233] ));
 sg13g2_a21oi_1 _3535_ (.A1(net556),
    .A2(\load_weights[233] ),
    .Y(_0350_),
    .B1(_0349_));
 sg13g2_a21o_1 _3536_ (.A2(\load_weights[233] ),
    .A1(net556),
    .B1(_0349_),
    .X(_0351_));
 sg13g2_nor3_1 _3537_ (.A(_0345_),
    .B(_0347_),
    .C(_0351_),
    .Y(_0352_));
 sg13g2_nand3_1 _3538_ (.B(_0348_),
    .C(_0350_),
    .A(_0346_),
    .Y(_0353_));
 sg13g2_a21oi_1 _3539_ (.A1(_0346_),
    .A2(_0348_),
    .Y(_0354_),
    .B1(_0350_));
 sg13g2_o21ai_1 _3540_ (.B1(_0351_),
    .Y(_0355_),
    .A1(_0345_),
    .A2(_0347_));
 sg13g2_a21oi_1 _3541_ (.A1(net518),
    .A2(\load_weights[217] ),
    .Y(_0356_),
    .B1(\load_weights[229] ));
 sg13g2_a21oi_2 _3542_ (.B1(_0356_),
    .Y(_0357_),
    .A2(\load_weights[229] ),
    .A1(net518));
 sg13g2_a21o_1 _3543_ (.A2(\load_weights[229] ),
    .A1(net518),
    .B1(_0356_),
    .X(_0358_));
 sg13g2_nor3_1 _3544_ (.A(_0352_),
    .B(_0354_),
    .C(_0358_),
    .Y(_0359_));
 sg13g2_nand3_1 _3545_ (.B(_0355_),
    .C(_0357_),
    .A(_0353_),
    .Y(_0360_));
 sg13g2_a21oi_1 _3546_ (.A1(_0353_),
    .A2(_0355_),
    .Y(_0361_),
    .B1(_0357_));
 sg13g2_o21ai_1 _3547_ (.B1(_0358_),
    .Y(_0362_),
    .A1(_0352_),
    .A2(_0354_));
 sg13g2_a21oi_1 _3548_ (.A1(net542),
    .A2(\load_weights[224] ),
    .Y(_0363_),
    .B1(\load_weights[236] ));
 sg13g2_a21oi_1 _3549_ (.A1(net542),
    .A2(\load_weights[236] ),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_a21o_1 _3550_ (.A2(\load_weights[236] ),
    .A1(net542),
    .B1(_0363_),
    .X(_0365_));
 sg13g2_nor3_1 _3551_ (.A(_0359_),
    .B(_0361_),
    .C(_0365_),
    .Y(_0366_));
 sg13g2_nand3_1 _3552_ (.B(_0362_),
    .C(_0364_),
    .A(_0360_),
    .Y(_0367_));
 sg13g2_a21oi_1 _3553_ (.A1(_0360_),
    .A2(_0362_),
    .Y(_0368_),
    .B1(_0364_));
 sg13g2_o21ai_1 _3554_ (.B1(_0365_),
    .Y(_0369_),
    .A1(_0359_),
    .A2(_0361_));
 sg13g2_a21oi_1 _3555_ (.A1(net524),
    .A2(\load_weights[216] ),
    .Y(_0370_),
    .B1(\load_weights[228] ));
 sg13g2_a21o_1 _3556_ (.A2(\load_weights[228] ),
    .A1(net524),
    .B1(_0370_),
    .X(_0371_));
 sg13g2_inv_1 _3557_ (.Y(_0372_),
    .A(_0371_));
 sg13g2_nor3_1 _3558_ (.A(_0366_),
    .B(_0368_),
    .C(_0371_),
    .Y(_0373_));
 sg13g2_a21oi_1 _3559_ (.A1(_0367_),
    .A2(_0369_),
    .Y(_0374_),
    .B1(_0372_));
 sg13g2_nand3_1 _3560_ (.B(_0369_),
    .C(_0371_),
    .A(_0367_),
    .Y(_0375_));
 sg13g2_o21ai_1 _3561_ (.B1(_0372_),
    .Y(_0376_),
    .A1(_0366_),
    .A2(_0368_));
 sg13g2_a21oi_1 _3562_ (.A1(net533),
    .A2(\load_weights[226] ),
    .Y(_0377_),
    .B1(\load_weights[238] ));
 sg13g2_a21o_1 _3563_ (.A2(\load_weights[238] ),
    .A1(net533),
    .B1(_0377_),
    .X(_0378_));
 sg13g2_nor3_2 _3564_ (.A(_0373_),
    .B(_0374_),
    .C(_0378_),
    .Y(_0379_));
 sg13g2_and3_1 _3565_ (.X(_0380_),
    .A(_0375_),
    .B(_0376_),
    .C(_0378_));
 sg13g2_o21ai_1 _3566_ (.B1(_0378_),
    .Y(_0381_),
    .A1(_0373_),
    .A2(_0374_));
 sg13g2_a21oi_1 _3567_ (.A1(net561),
    .A2(net410),
    .Y(_0382_),
    .B1(net609));
 sg13g2_a21oi_2 _3568_ (.B1(_0382_),
    .Y(_0383_),
    .A2(net609),
    .A1(net560));
 sg13g2_nor3_1 _3569_ (.A(_0379_),
    .B(_0380_),
    .C(_0383_),
    .Y(_0384_));
 sg13g2_o21ai_1 _3570_ (.B1(_0383_),
    .Y(_0385_),
    .A1(_0379_),
    .A2(_0380_));
 sg13g2_nand2b_1 _3571_ (.Y(\tt_um_mult_inst.genblk1[9].out_q ),
    .B(_0385_),
    .A_N(_0384_));
 sg13g2_a21oi_2 _3572_ (.B1(_0379_),
    .Y(_0386_),
    .A2(_0383_),
    .A1(_0381_));
 sg13g2_o21ai_1 _3573_ (.B1(_2121_),
    .Y(_0387_),
    .A1(_2115_),
    .A2(_2117_));
 sg13g2_nand2b_1 _3574_ (.Y(_0388_),
    .B(_0346_),
    .A_N(_0341_));
 sg13g2_o21ai_1 _3575_ (.B1(_2132_),
    .Y(_0389_),
    .A1(_2125_),
    .A2(_2127_));
 sg13g2_nor2_1 _3576_ (.A(\tt_um_mult_inst.genblk1[9].carry[1] ),
    .B(net441),
    .Y(_0390_));
 sg13g2_nand2_1 _3577_ (.Y(_0391_),
    .A(_2153_),
    .B(_0337_));
 sg13g2_a21oi_2 _3578_ (.B1(_2145_),
    .Y(_0392_),
    .A2(_2146_),
    .A1(\load_weights[239] ));
 sg13g2_a21oi_1 _3579_ (.A1(\load_weights[233] ),
    .A2(_2141_),
    .Y(_0393_),
    .B1(_2140_));
 sg13g2_nor2_1 _3580_ (.A(_2138_),
    .B(_0393_),
    .Y(_0394_));
 sg13g2_xnor2_1 _3581_ (.Y(_0395_),
    .A(_2138_),
    .B(_0393_));
 sg13g2_nor2_1 _3582_ (.A(_2143_),
    .B(_2148_),
    .Y(_0396_));
 sg13g2_nor2_1 _3583_ (.A(_0395_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_xnor2_1 _3584_ (.Y(_0398_),
    .A(_0395_),
    .B(_0396_));
 sg13g2_nor2_1 _3585_ (.A(_0392_),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_xor2_1 _3586_ (.B(_0398_),
    .A(_0392_),
    .X(_0400_));
 sg13g2_o21ai_1 _3587_ (.B1(_2150_),
    .Y(_0401_),
    .A1(_1930_),
    .A2(_2151_));
 sg13g2_and2_1 _3588_ (.A(_0400_),
    .B(_0401_),
    .X(_0402_));
 sg13g2_xor2_1 _3589_ (.B(_0401_),
    .A(_0400_),
    .X(_0403_));
 sg13g2_xnor2_1 _3590_ (.Y(_0404_),
    .A(_0391_),
    .B(_0403_));
 sg13g2_a21oi_1 _3591_ (.A1(net441),
    .A2(_0404_),
    .Y(_0405_),
    .B1(_0390_));
 sg13g2_nand2_1 _3592_ (.Y(_0406_),
    .A(_0389_),
    .B(_0405_));
 sg13g2_xor2_1 _3593_ (.B(_0405_),
    .A(_0389_),
    .X(_0407_));
 sg13g2_nand2_1 _3594_ (.Y(_0408_),
    .A(_0388_),
    .B(_0407_));
 sg13g2_xnor2_1 _3595_ (.Y(_0409_),
    .A(_0388_),
    .B(_0407_));
 sg13g2_nand2b_1 _3596_ (.Y(_0410_),
    .B(_0387_),
    .A_N(_0409_));
 sg13g2_xor2_1 _3597_ (.B(_0409_),
    .A(_0387_),
    .X(_0411_));
 sg13g2_nand2_1 _3598_ (.Y(_0412_),
    .A(_0353_),
    .B(_0360_));
 sg13g2_nand2b_1 _3599_ (.Y(_0413_),
    .B(_0412_),
    .A_N(_0411_));
 sg13g2_xnor2_1 _3600_ (.Y(_0414_),
    .A(_0411_),
    .B(_0412_));
 sg13g2_o21ai_1 _3601_ (.B1(_0367_),
    .Y(_0415_),
    .A1(_0368_),
    .A2(_0371_));
 sg13g2_nand2_1 _3602_ (.Y(_0416_),
    .A(_0414_),
    .B(_0415_));
 sg13g2_xnor2_1 _3603_ (.Y(_0417_),
    .A(_0414_),
    .B(_0415_));
 sg13g2_xor2_1 _3604_ (.B(_0417_),
    .A(_0386_),
    .X(\tt_um_mult_inst.genblk1[9].carry_q[0] ));
 sg13g2_o21ai_1 _3605_ (.B1(_0416_),
    .Y(_0418_),
    .A1(_0386_),
    .A2(_0417_));
 sg13g2_nand2_1 _3606_ (.Y(_0419_),
    .A(_0394_),
    .B(_0399_));
 sg13g2_nor3_1 _3607_ (.A(_0394_),
    .B(_0397_),
    .C(_0399_),
    .Y(_0420_));
 sg13g2_a21oi_1 _3608_ (.A1(_0394_),
    .A2(_0399_),
    .Y(_0421_),
    .B1(_0420_));
 sg13g2_a21o_1 _3609_ (.A2(_0403_),
    .A1(_0391_),
    .B1(_0402_),
    .X(_0422_));
 sg13g2_or2_1 _3610_ (.X(_0423_),
    .B(_0422_),
    .A(_0421_));
 sg13g2_a21oi_1 _3611_ (.A1(_0421_),
    .A2(_0422_),
    .Y(_0424_),
    .B1(net432));
 sg13g2_a22oi_1 _3612_ (.Y(_0425_),
    .B1(_0423_),
    .B2(_0424_),
    .A2(net432),
    .A1(\tt_um_mult_inst.genblk1[9].carry[2] ));
 sg13g2_xnor2_1 _3613_ (.Y(_0426_),
    .A(_0406_),
    .B(_0425_));
 sg13g2_a21o_1 _3614_ (.A2(_0410_),
    .A1(_0408_),
    .B1(_0426_),
    .X(_0427_));
 sg13g2_nand3_1 _3615_ (.B(_0410_),
    .C(_0426_),
    .A(_0408_),
    .Y(_0428_));
 sg13g2_nand2_1 _3616_ (.Y(_0429_),
    .A(_0427_),
    .B(_0428_));
 sg13g2_nor2_1 _3617_ (.A(_0413_),
    .B(_0429_),
    .Y(_0430_));
 sg13g2_xor2_1 _3618_ (.B(_0429_),
    .A(_0413_),
    .X(_0431_));
 sg13g2_xor2_1 _3619_ (.B(_0431_),
    .A(_0418_),
    .X(\tt_um_mult_inst.genblk1[9].carry_q[1] ));
 sg13g2_a21oi_1 _3620_ (.A1(_0418_),
    .A2(_0431_),
    .Y(_0432_),
    .B1(_0430_));
 sg13g2_a22oi_1 _3621_ (.Y(_0433_),
    .B1(_0419_),
    .B2(_0424_),
    .A2(net432),
    .A1(net920));
 sg13g2_o21ai_1 _3622_ (.B1(_0427_),
    .Y(_0434_),
    .A1(_0406_),
    .A2(_0425_));
 sg13g2_xor2_1 _3623_ (.B(_0434_),
    .A(_0433_),
    .X(_0435_));
 sg13g2_nor2b_1 _3624_ (.A(_0432_),
    .B_N(_0435_),
    .Y(_0436_));
 sg13g2_xnor2_1 _3625_ (.Y(\tt_um_mult_inst.genblk1[9].carry_q[2] ),
    .A(_0432_),
    .B(_0435_));
 sg13g2_a21o_1 _3626_ (.A2(_0434_),
    .A1(_0433_),
    .B1(_0436_),
    .X(\tt_um_mult_inst.genblk1[9].carry_q[3] ));
 sg13g2_a21oi_1 _3627_ (.A1(net548),
    .A2(\load_weights[270] ),
    .Y(_0437_),
    .B1(\load_weights[282] ));
 sg13g2_a21o_1 _3628_ (.A2(\load_weights[282] ),
    .A1(net548),
    .B1(_0437_),
    .X(_0438_));
 sg13g2_a21oi_1 _3629_ (.A1(net559),
    .A2(\load_weights[268] ),
    .Y(_0439_),
    .B1(\load_weights[280] ));
 sg13g2_a21o_1 _3630_ (.A2(\load_weights[280] ),
    .A1(net558),
    .B1(_0439_),
    .X(_0440_));
 sg13g2_xor2_1 _3631_ (.B(_0440_),
    .A(_0438_),
    .X(_0441_));
 sg13g2_a21oi_1 _3632_ (.A1(net512),
    .A2(\load_weights[266] ),
    .Y(_0442_),
    .B1(\load_weights[278] ));
 sg13g2_a21oi_1 _3633_ (.A1(net512),
    .A2(\load_weights[278] ),
    .Y(_0443_),
    .B1(_0442_));
 sg13g2_nand2_1 _3634_ (.Y(_0444_),
    .A(_0441_),
    .B(_0443_));
 sg13g2_xnor2_1 _3635_ (.Y(_0445_),
    .A(_0441_),
    .B(_0443_));
 sg13g2_inv_1 _3636_ (.Y(_0446_),
    .A(_0445_));
 sg13g2_a21oi_1 _3637_ (.A1(net527),
    .A2(\load_weights[275] ),
    .Y(_0447_),
    .B1(\load_weights[287] ));
 sg13g2_a21o_1 _3638_ (.A2(\load_weights[287] ),
    .A1(net527),
    .B1(_0447_),
    .X(_0448_));
 sg13g2_a21oi_1 _3639_ (.A1(net531),
    .A2(\load_weights[274] ),
    .Y(_0449_),
    .B1(\load_weights[286] ));
 sg13g2_a21o_1 _3640_ (.A2(\load_weights[286] ),
    .A1(net531),
    .B1(_0449_),
    .X(_0450_));
 sg13g2_xor2_1 _3641_ (.B(_0450_),
    .A(_0448_),
    .X(_0451_));
 sg13g2_a21oi_1 _3642_ (.A1(net540),
    .A2(\load_weights[272] ),
    .Y(_0452_),
    .B1(\load_weights[284] ));
 sg13g2_a21o_1 _3643_ (.A2(\load_weights[284] ),
    .A1(net540),
    .B1(_0452_),
    .X(_0453_));
 sg13g2_inv_1 _3644_ (.Y(_0454_),
    .A(_0453_));
 sg13g2_nand2_1 _3645_ (.Y(_0455_),
    .A(_0451_),
    .B(_0454_));
 sg13g2_nand2b_1 _3646_ (.Y(_0456_),
    .B(_0453_),
    .A_N(_0451_));
 sg13g2_nand2_1 _3647_ (.Y(_0457_),
    .A(_0451_),
    .B(_0453_));
 sg13g2_nand2b_1 _3648_ (.Y(_0458_),
    .B(_0454_),
    .A_N(_0451_));
 sg13g2_nand2_1 _3649_ (.Y(_0459_),
    .A(_0455_),
    .B(_0456_));
 sg13g2_inv_1 _3650_ (.Y(_0460_),
    .A(_0459_));
 sg13g2_nand2_1 _3651_ (.Y(_0461_),
    .A(\load_weights[276] ),
    .B(\load_weights[277] ));
 sg13g2_xnor2_1 _3652_ (.Y(_0462_),
    .A(\load_weights[276] ),
    .B(\load_weights[277] ));
 sg13g2_and2_1 _3653_ (.A(\load_weights[278] ),
    .B(\load_weights[279] ),
    .X(_0463_));
 sg13g2_xor2_1 _3654_ (.B(\load_weights[279] ),
    .A(\load_weights[278] ),
    .X(_0464_));
 sg13g2_xnor2_1 _3655_ (.Y(_0465_),
    .A(\load_weights[281] ),
    .B(_0464_));
 sg13g2_nor2_1 _3656_ (.A(_0462_),
    .B(_0465_),
    .Y(_0466_));
 sg13g2_xnor2_1 _3657_ (.Y(_0467_),
    .A(_0462_),
    .B(_0465_));
 sg13g2_and2_1 _3658_ (.A(\load_weights[283] ),
    .B(\load_weights[285] ),
    .X(_0468_));
 sg13g2_xor2_1 _3659_ (.B(\load_weights[285] ),
    .A(\load_weights[283] ),
    .X(_0469_));
 sg13g2_xnor2_1 _3660_ (.Y(_0470_),
    .A(\load_weights[287] ),
    .B(_0469_));
 sg13g2_nor2_1 _3661_ (.A(_0467_),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_xor2_1 _3662_ (.B(_0470_),
    .A(_0467_),
    .X(_0472_));
 sg13g2_nand2_1 _3663_ (.Y(_0473_),
    .A(\load_weights[284] ),
    .B(_0472_));
 sg13g2_xnor2_1 _3664_ (.Y(_0474_),
    .A(\load_weights[284] ),
    .B(_0472_));
 sg13g2_xnor2_1 _3665_ (.Y(_0475_),
    .A(\load_weights[286] ),
    .B(_0474_));
 sg13g2_nand2_1 _3666_ (.Y(_0476_),
    .A(\load_weights[282] ),
    .B(_0475_));
 sg13g2_xor2_1 _3667_ (.B(_0475_),
    .A(\load_weights[282] ),
    .X(_0477_));
 sg13g2_xnor2_1 _3668_ (.Y(_0478_),
    .A(\load_weights[282] ),
    .B(_0475_));
 sg13g2_nand2_1 _3669_ (.Y(_0479_),
    .A(\load_weights[280] ),
    .B(_0477_));
 sg13g2_a21oi_1 _3670_ (.A1(_1934_),
    .A2(_0478_),
    .Y(_0480_),
    .B1(net427));
 sg13g2_xnor2_1 _3671_ (.Y(_0481_),
    .A(\load_weights[280] ),
    .B(_0477_));
 sg13g2_nor2_1 _3672_ (.A(_1935_),
    .B(net438),
    .Y(_0482_));
 sg13g2_a221oi_1 _3673_ (.B2(net438),
    .C1(_0482_),
    .B1(_0481_),
    .A1(_0457_),
    .Y(_0483_),
    .A2(_0458_));
 sg13g2_a221oi_1 _3674_ (.B2(_0480_),
    .C1(_0460_),
    .B1(_0479_),
    .A1(_1935_),
    .Y(_0484_),
    .A2(net427));
 sg13g2_a221oi_1 _3675_ (.B2(_0480_),
    .C1(_0459_),
    .B1(_0479_),
    .A1(_1935_),
    .Y(_0485_),
    .A2(net426));
 sg13g2_a221oi_1 _3676_ (.B2(net438),
    .C1(_0482_),
    .B1(_0481_),
    .A1(_0455_),
    .Y(_0486_),
    .A2(_0456_));
 sg13g2_nor3_1 _3677_ (.A(_0445_),
    .B(_0483_),
    .C(_0484_),
    .Y(_0487_));
 sg13g2_o21ai_1 _3678_ (.B1(_0446_),
    .Y(_0488_),
    .A1(_0485_),
    .A2(_0486_));
 sg13g2_nor3_1 _3679_ (.A(_0446_),
    .B(_0485_),
    .C(_0486_),
    .Y(_0489_));
 sg13g2_o21ai_1 _3680_ (.B1(_0445_),
    .Y(_0490_),
    .A1(_0483_),
    .A2(_0484_));
 sg13g2_a21oi_1 _3681_ (.A1(net507),
    .A2(\load_weights[267] ),
    .Y(_0491_),
    .B1(\load_weights[279] ));
 sg13g2_a21oi_1 _3682_ (.A1(net507),
    .A2(\load_weights[279] ),
    .Y(_0492_),
    .B1(_0491_));
 sg13g2_a21o_1 _3683_ (.A2(\load_weights[279] ),
    .A1(net507),
    .B1(_0491_),
    .X(_0493_));
 sg13g2_nor3_1 _3684_ (.A(_0487_),
    .B(_0489_),
    .C(_0493_),
    .Y(_0494_));
 sg13g2_nand3_1 _3685_ (.B(_0490_),
    .C(_0492_),
    .A(_0488_),
    .Y(_0495_));
 sg13g2_a21oi_1 _3686_ (.A1(_0488_),
    .A2(_0490_),
    .Y(_0496_),
    .B1(_0492_));
 sg13g2_o21ai_1 _3687_ (.B1(_0493_),
    .Y(_0497_),
    .A1(_0487_),
    .A2(_0489_));
 sg13g2_a21oi_1 _3688_ (.A1(net517),
    .A2(\load_weights[265] ),
    .Y(_0498_),
    .B1(\load_weights[277] ));
 sg13g2_a21oi_1 _3689_ (.A1(net517),
    .A2(\load_weights[277] ),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_a21o_1 _3690_ (.A2(\load_weights[277] ),
    .A1(net517),
    .B1(_0498_),
    .X(_0500_));
 sg13g2_nor3_1 _3691_ (.A(_0494_),
    .B(_0496_),
    .C(_0500_),
    .Y(_0501_));
 sg13g2_nand3_1 _3692_ (.B(_0497_),
    .C(_0499_),
    .A(_0495_),
    .Y(_0502_));
 sg13g2_a21oi_1 _3693_ (.A1(_0495_),
    .A2(_0497_),
    .Y(_0503_),
    .B1(_0499_));
 sg13g2_o21ai_1 _3694_ (.B1(_0500_),
    .Y(_0504_),
    .A1(_0494_),
    .A2(_0496_));
 sg13g2_a21oi_1 _3695_ (.A1(net557),
    .A2(\load_weights[269] ),
    .Y(_0505_),
    .B1(\load_weights[281] ));
 sg13g2_a21oi_1 _3696_ (.A1(net557),
    .A2(\load_weights[281] ),
    .Y(_0506_),
    .B1(_0505_));
 sg13g2_a21o_1 _3697_ (.A2(\load_weights[281] ),
    .A1(net557),
    .B1(_0505_),
    .X(_0507_));
 sg13g2_nor3_1 _3698_ (.A(_0501_),
    .B(_0503_),
    .C(_0507_),
    .Y(_0508_));
 sg13g2_nand3_1 _3699_ (.B(_0504_),
    .C(_0506_),
    .A(_0502_),
    .Y(_0509_));
 sg13g2_a21oi_1 _3700_ (.A1(_0502_),
    .A2(_0504_),
    .Y(_0510_),
    .B1(_0506_));
 sg13g2_o21ai_1 _3701_ (.B1(_0507_),
    .Y(_0511_),
    .A1(_0501_),
    .A2(_0503_));
 sg13g2_a21oi_1 _3702_ (.A1(net522),
    .A2(\load_weights[264] ),
    .Y(_0512_),
    .B1(\load_weights[276] ));
 sg13g2_a21o_1 _3703_ (.A2(\load_weights[276] ),
    .A1(net522),
    .B1(_0512_),
    .X(_0513_));
 sg13g2_inv_1 _3704_ (.Y(_0514_),
    .A(_0513_));
 sg13g2_nor3_1 _3705_ (.A(_0508_),
    .B(_0510_),
    .C(_0513_),
    .Y(_0515_));
 sg13g2_a21oi_1 _3706_ (.A1(_0509_),
    .A2(_0511_),
    .Y(_0516_),
    .B1(_0514_));
 sg13g2_nand3_1 _3707_ (.B(_0511_),
    .C(_0513_),
    .A(_0509_),
    .Y(_0517_));
 sg13g2_o21ai_1 _3708_ (.B1(_0514_),
    .Y(_0518_),
    .A1(_0508_),
    .A2(_0510_));
 sg13g2_a21oi_1 _3709_ (.A1(net544),
    .A2(\load_weights[271] ),
    .Y(_0519_),
    .B1(\load_weights[283] ));
 sg13g2_a21o_1 _3710_ (.A2(\load_weights[283] ),
    .A1(net545),
    .B1(_0519_),
    .X(_0520_));
 sg13g2_nor3_2 _3711_ (.A(_0515_),
    .B(_0516_),
    .C(_0520_),
    .Y(_0521_));
 sg13g2_and3_1 _3712_ (.X(_0522_),
    .A(_0517_),
    .B(_0518_),
    .C(_0520_));
 sg13g2_o21ai_1 _3713_ (.B1(_0520_),
    .Y(_0523_),
    .A1(_0515_),
    .A2(_0516_));
 sg13g2_a21oi_1 _3714_ (.A1(net538),
    .A2(\load_weights[273] ),
    .Y(_0524_),
    .B1(\load_weights[285] ));
 sg13g2_a21oi_2 _3715_ (.B1(_0524_),
    .Y(_0525_),
    .A2(\load_weights[285] ),
    .A1(net536));
 sg13g2_nor3_1 _3716_ (.A(_0521_),
    .B(_0522_),
    .C(_0525_),
    .Y(_0526_));
 sg13g2_o21ai_1 _3717_ (.B1(_0525_),
    .Y(_0527_),
    .A1(_0521_),
    .A2(_0522_));
 sg13g2_nand2b_2 _3718_ (.Y(\tt_um_mult_inst.genblk1[11].out_q ),
    .B(_0527_),
    .A_N(_0526_));
 sg13g2_a21oi_2 _3719_ (.B1(_0521_),
    .Y(_0528_),
    .A2(_0525_),
    .A1(_0523_));
 sg13g2_o21ai_1 _3720_ (.B1(_0444_),
    .Y(_0529_),
    .A1(_0438_),
    .A2(_0440_));
 sg13g2_nand2b_1 _3721_ (.Y(_0530_),
    .B(_0488_),
    .A_N(_0483_));
 sg13g2_o21ai_1 _3722_ (.B1(_0455_),
    .Y(_0531_),
    .A1(_0448_),
    .A2(_0450_));
 sg13g2_nand2_1 _3723_ (.Y(_0532_),
    .A(\tt_um_mult_inst.genblk1[11].carry[1] ),
    .B(net426));
 sg13g2_nand2_1 _3724_ (.Y(_0533_),
    .A(_0476_),
    .B(_0479_));
 sg13g2_a21oi_2 _3725_ (.B1(_0468_),
    .Y(_0534_),
    .A2(_0469_),
    .A1(\load_weights[287] ));
 sg13g2_a21oi_1 _3726_ (.A1(\load_weights[281] ),
    .A2(_0464_),
    .Y(_0535_),
    .B1(_0463_));
 sg13g2_nor2_1 _3727_ (.A(_0461_),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_xnor2_1 _3728_ (.Y(_0537_),
    .A(_0461_),
    .B(_0535_));
 sg13g2_nor2_1 _3729_ (.A(_0466_),
    .B(_0471_),
    .Y(_0538_));
 sg13g2_nor2_1 _3730_ (.A(_0537_),
    .B(_0538_),
    .Y(_0539_));
 sg13g2_xnor2_1 _3731_ (.Y(_0540_),
    .A(_0537_),
    .B(_0538_));
 sg13g2_nor2_1 _3732_ (.A(_0534_),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_xor2_1 _3733_ (.B(_0540_),
    .A(_0534_),
    .X(_0542_));
 sg13g2_o21ai_1 _3734_ (.B1(_0473_),
    .Y(_0543_),
    .A1(_1933_),
    .A2(_0474_));
 sg13g2_and2_1 _3735_ (.A(_0542_),
    .B(_0543_),
    .X(_0544_));
 sg13g2_xor2_1 _3736_ (.B(_0543_),
    .A(_0542_),
    .X(_0545_));
 sg13g2_xnor2_1 _3737_ (.Y(_0546_),
    .A(_0533_),
    .B(_0545_));
 sg13g2_o21ai_1 _3738_ (.B1(_0532_),
    .Y(_0547_),
    .A1(net426),
    .A2(_0546_));
 sg13g2_nand2_1 _3739_ (.Y(_0548_),
    .A(_0531_),
    .B(_0547_));
 sg13g2_xor2_1 _3740_ (.B(_0547_),
    .A(_0531_),
    .X(_0549_));
 sg13g2_nand2_1 _3741_ (.Y(_0550_),
    .A(_0530_),
    .B(_0549_));
 sg13g2_xnor2_1 _3742_ (.Y(_0551_),
    .A(_0530_),
    .B(_0549_));
 sg13g2_nand2b_1 _3743_ (.Y(_0552_),
    .B(_0529_),
    .A_N(_0551_));
 sg13g2_xor2_1 _3744_ (.B(_0551_),
    .A(_0529_),
    .X(_0553_));
 sg13g2_nand2_2 _3745_ (.Y(_0554_),
    .A(_0495_),
    .B(_0502_));
 sg13g2_nand2b_1 _3746_ (.Y(_0555_),
    .B(_0554_),
    .A_N(_0553_));
 sg13g2_xnor2_1 _3747_ (.Y(_0556_),
    .A(_0553_),
    .B(_0554_));
 sg13g2_o21ai_1 _3748_ (.B1(_0509_),
    .Y(_0557_),
    .A1(_0510_),
    .A2(_0513_));
 sg13g2_nand2_1 _3749_ (.Y(_0558_),
    .A(_0556_),
    .B(_0557_));
 sg13g2_xnor2_1 _3750_ (.Y(_0559_),
    .A(_0556_),
    .B(_0557_));
 sg13g2_xor2_1 _3751_ (.B(_0559_),
    .A(_0528_),
    .X(\tt_um_mult_inst.genblk1[11].carry_q[0] ));
 sg13g2_o21ai_1 _3752_ (.B1(_0558_),
    .Y(_0560_),
    .A1(_0528_),
    .A2(_0559_));
 sg13g2_nand2_1 _3753_ (.Y(_0561_),
    .A(_0536_),
    .B(_0541_));
 sg13g2_nor3_1 _3754_ (.A(_0536_),
    .B(_0539_),
    .C(_0541_),
    .Y(_0562_));
 sg13g2_a21oi_1 _3755_ (.A1(_0536_),
    .A2(_0541_),
    .Y(_0563_),
    .B1(_0562_));
 sg13g2_a21o_1 _3756_ (.A2(_0545_),
    .A1(_0533_),
    .B1(_0544_),
    .X(_0564_));
 sg13g2_or2_1 _3757_ (.X(_0565_),
    .B(_0564_),
    .A(_0563_));
 sg13g2_a21oi_1 _3758_ (.A1(_0563_),
    .A2(_0564_),
    .Y(_0566_),
    .B1(net426));
 sg13g2_a22oi_1 _3759_ (.Y(_0567_),
    .B1(_0565_),
    .B2(_0566_),
    .A2(net426),
    .A1(\tt_um_mult_inst.genblk1[11].carry[2] ));
 sg13g2_nor2_1 _3760_ (.A(_0548_),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_xnor2_1 _3761_ (.Y(_0569_),
    .A(_0548_),
    .B(_0567_));
 sg13g2_a21o_1 _3762_ (.A2(_0552_),
    .A1(_0550_),
    .B1(_0569_),
    .X(_0570_));
 sg13g2_nand3_1 _3763_ (.B(_0552_),
    .C(_0569_),
    .A(_0550_),
    .Y(_0571_));
 sg13g2_nand2_1 _3764_ (.Y(_0572_),
    .A(_0570_),
    .B(_0571_));
 sg13g2_nor2_1 _3765_ (.A(_0555_),
    .B(_0572_),
    .Y(_0573_));
 sg13g2_xor2_1 _3766_ (.B(_0572_),
    .A(_0555_),
    .X(_0574_));
 sg13g2_xor2_1 _3767_ (.B(_0574_),
    .A(_0560_),
    .X(\tt_um_mult_inst.genblk1[11].carry_q[1] ));
 sg13g2_a22oi_1 _3768_ (.Y(_0575_),
    .B1(_0561_),
    .B2(_0566_),
    .A2(net426),
    .A1(net922));
 sg13g2_xnor2_1 _3769_ (.Y(_0576_),
    .A(_0568_),
    .B(_0575_));
 sg13g2_nor2_1 _3770_ (.A(_0570_),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_xor2_1 _3771_ (.B(_0576_),
    .A(_0570_),
    .X(_0578_));
 sg13g2_a21oi_1 _3772_ (.A1(_0560_),
    .A2(_0574_),
    .Y(_0579_),
    .B1(_0573_));
 sg13g2_nand2b_1 _3773_ (.Y(_0580_),
    .B(_0578_),
    .A_N(_0579_));
 sg13g2_xnor2_1 _3774_ (.Y(\tt_um_mult_inst.genblk1[11].carry_q[2] ),
    .A(_0578_),
    .B(_0579_));
 sg13g2_a21oi_1 _3775_ (.A1(_0568_),
    .A2(_0575_),
    .Y(_0581_),
    .B1(_0577_));
 sg13g2_nand2_1 _3776_ (.Y(\tt_um_mult_inst.genblk1[11].carry_q[3] ),
    .A(_0580_),
    .B(net923));
 sg13g2_a21oi_1 _3777_ (.A1(net548),
    .A2(\load_weights[198] ),
    .Y(_0582_),
    .B1(\load_weights[210] ));
 sg13g2_a21o_1 _3778_ (.A2(\load_weights[210] ),
    .A1(net552),
    .B1(_0582_),
    .X(_0583_));
 sg13g2_a21oi_1 _3779_ (.A1(net559),
    .A2(\load_weights[196] ),
    .Y(_0584_),
    .B1(\load_weights[208] ));
 sg13g2_a21o_1 _3780_ (.A2(\load_weights[208] ),
    .A1(net559),
    .B1(_0584_),
    .X(_0585_));
 sg13g2_xor2_1 _3781_ (.B(_0585_),
    .A(_0583_),
    .X(_0586_));
 sg13g2_a21oi_1 _3782_ (.A1(net512),
    .A2(\load_weights[194] ),
    .Y(_0587_),
    .B1(\load_weights[206] ));
 sg13g2_a21oi_1 _3783_ (.A1(net512),
    .A2(\load_weights[206] ),
    .Y(_0588_),
    .B1(_0587_));
 sg13g2_nand2_1 _3784_ (.Y(_0589_),
    .A(_0586_),
    .B(_0588_));
 sg13g2_xnor2_1 _3785_ (.Y(_0590_),
    .A(_0586_),
    .B(_0588_));
 sg13g2_inv_1 _3786_ (.Y(_0591_),
    .A(_0590_));
 sg13g2_a21oi_1 _3787_ (.A1(net527),
    .A2(\load_weights[203] ),
    .Y(_0592_),
    .B1(\load_weights[215] ));
 sg13g2_a21o_1 _3788_ (.A2(\load_weights[215] ),
    .A1(net527),
    .B1(_0592_),
    .X(_0593_));
 sg13g2_a21oi_1 _3789_ (.A1(net531),
    .A2(\load_weights[202] ),
    .Y(_0594_),
    .B1(\load_weights[214] ));
 sg13g2_a21o_1 _3790_ (.A2(\load_weights[214] ),
    .A1(net530),
    .B1(_0594_),
    .X(_0595_));
 sg13g2_xor2_1 _3791_ (.B(_0595_),
    .A(_0593_),
    .X(_0596_));
 sg13g2_a21oi_1 _3792_ (.A1(net540),
    .A2(\load_weights[200] ),
    .Y(_0597_),
    .B1(\load_weights[212] ));
 sg13g2_a21o_1 _3793_ (.A2(\load_weights[212] ),
    .A1(net540),
    .B1(_0597_),
    .X(_0598_));
 sg13g2_inv_1 _3794_ (.Y(_0599_),
    .A(_0598_));
 sg13g2_nand2_1 _3795_ (.Y(_0600_),
    .A(_0596_),
    .B(_0599_));
 sg13g2_nand2b_1 _3796_ (.Y(_0601_),
    .B(_0598_),
    .A_N(_0596_));
 sg13g2_nand2_1 _3797_ (.Y(_0602_),
    .A(_0596_),
    .B(_0598_));
 sg13g2_nand2b_1 _3798_ (.Y(_0603_),
    .B(_0599_),
    .A_N(_0596_));
 sg13g2_nand2_1 _3799_ (.Y(_0604_),
    .A(_0600_),
    .B(_0601_));
 sg13g2_inv_1 _3800_ (.Y(_0605_),
    .A(_0604_));
 sg13g2_nand2_1 _3801_ (.Y(_0606_),
    .A(\load_weights[204] ),
    .B(\load_weights[205] ));
 sg13g2_xnor2_1 _3802_ (.Y(_0607_),
    .A(\load_weights[204] ),
    .B(\load_weights[205] ));
 sg13g2_and2_1 _3803_ (.A(\load_weights[206] ),
    .B(\load_weights[207] ),
    .X(_0608_));
 sg13g2_xor2_1 _3804_ (.B(\load_weights[207] ),
    .A(\load_weights[206] ),
    .X(_0609_));
 sg13g2_xnor2_1 _3805_ (.Y(_0610_),
    .A(\load_weights[209] ),
    .B(_0609_));
 sg13g2_nor2_1 _3806_ (.A(_0607_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_xnor2_1 _3807_ (.Y(_0612_),
    .A(_0607_),
    .B(_0610_));
 sg13g2_and2_1 _3808_ (.A(\load_weights[211] ),
    .B(\load_weights[213] ),
    .X(_0613_));
 sg13g2_xor2_1 _3809_ (.B(\load_weights[213] ),
    .A(\load_weights[211] ),
    .X(_0614_));
 sg13g2_xnor2_1 _3810_ (.Y(_0615_),
    .A(\load_weights[215] ),
    .B(_0614_));
 sg13g2_nor2_1 _3811_ (.A(_0612_),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_xor2_1 _3812_ (.B(_0615_),
    .A(_0612_),
    .X(_0617_));
 sg13g2_nand2_1 _3813_ (.Y(_0618_),
    .A(\load_weights[212] ),
    .B(_0617_));
 sg13g2_xnor2_1 _3814_ (.Y(_0619_),
    .A(\load_weights[212] ),
    .B(_0617_));
 sg13g2_xnor2_1 _3815_ (.Y(_0620_),
    .A(\load_weights[214] ),
    .B(_0619_));
 sg13g2_nand2_1 _3816_ (.Y(_0621_),
    .A(\load_weights[210] ),
    .B(_0620_));
 sg13g2_xor2_1 _3817_ (.B(_0620_),
    .A(\load_weights[210] ),
    .X(_0622_));
 sg13g2_xnor2_1 _3818_ (.Y(_0623_),
    .A(\load_weights[210] ),
    .B(_0620_));
 sg13g2_nand2_1 _3819_ (.Y(_0624_),
    .A(\load_weights[208] ),
    .B(_0622_));
 sg13g2_a21oi_1 _3820_ (.A1(_1937_),
    .A2(_0623_),
    .Y(_0625_),
    .B1(net433));
 sg13g2_xnor2_1 _3821_ (.Y(_0626_),
    .A(\load_weights[208] ),
    .B(_0622_));
 sg13g2_nor2_1 _3822_ (.A(_1938_),
    .B(net439),
    .Y(_0627_));
 sg13g2_a221oi_1 _3823_ (.B2(net435),
    .C1(_0627_),
    .B1(_0626_),
    .A1(_0602_),
    .Y(_0628_),
    .A2(_0603_));
 sg13g2_a221oi_1 _3824_ (.B2(_0625_),
    .C1(_0605_),
    .B1(_0624_),
    .A1(_1938_),
    .Y(_0629_),
    .A2(net433));
 sg13g2_a221oi_1 _3825_ (.B2(_0625_),
    .C1(_0604_),
    .B1(_0624_),
    .A1(_1938_),
    .Y(_0630_),
    .A2(net433));
 sg13g2_a221oi_1 _3826_ (.B2(net435),
    .C1(_0627_),
    .B1(_0626_),
    .A1(_0600_),
    .Y(_0631_),
    .A2(_0601_));
 sg13g2_nor3_1 _3827_ (.A(_0590_),
    .B(_0628_),
    .C(_0629_),
    .Y(_0632_));
 sg13g2_o21ai_1 _3828_ (.B1(_0591_),
    .Y(_0633_),
    .A1(_0630_),
    .A2(_0631_));
 sg13g2_nor3_1 _3829_ (.A(_0591_),
    .B(_0630_),
    .C(_0631_),
    .Y(_0634_));
 sg13g2_o21ai_1 _3830_ (.B1(_0590_),
    .Y(_0635_),
    .A1(_0628_),
    .A2(_0629_));
 sg13g2_a21oi_1 _3831_ (.A1(net507),
    .A2(\load_weights[195] ),
    .Y(_0636_),
    .B1(\load_weights[207] ));
 sg13g2_a21oi_1 _3832_ (.A1(net506),
    .A2(\load_weights[207] ),
    .Y(_0637_),
    .B1(_0636_));
 sg13g2_a21o_1 _3833_ (.A2(\load_weights[207] ),
    .A1(net506),
    .B1(_0636_),
    .X(_0638_));
 sg13g2_nor3_1 _3834_ (.A(_0632_),
    .B(_0634_),
    .C(_0638_),
    .Y(_0639_));
 sg13g2_nand3_1 _3835_ (.B(_0635_),
    .C(_0637_),
    .A(_0633_),
    .Y(_0640_));
 sg13g2_a21oi_1 _3836_ (.A1(_0633_),
    .A2(_0635_),
    .Y(_0641_),
    .B1(_0637_));
 sg13g2_o21ai_1 _3837_ (.B1(_0638_),
    .Y(_0642_),
    .A1(_0632_),
    .A2(_0634_));
 sg13g2_a21oi_1 _3838_ (.A1(net517),
    .A2(\load_weights[193] ),
    .Y(_0643_),
    .B1(\load_weights[205] ));
 sg13g2_a21oi_1 _3839_ (.A1(net517),
    .A2(\load_weights[205] ),
    .Y(_0644_),
    .B1(_0643_));
 sg13g2_a21o_1 _3840_ (.A2(\load_weights[205] ),
    .A1(net517),
    .B1(_0643_),
    .X(_0645_));
 sg13g2_nor3_1 _3841_ (.A(_0639_),
    .B(_0641_),
    .C(_0645_),
    .Y(_0646_));
 sg13g2_nand3_1 _3842_ (.B(_0642_),
    .C(_0644_),
    .A(_0640_),
    .Y(_0647_));
 sg13g2_a21oi_1 _3843_ (.A1(_0640_),
    .A2(_0642_),
    .Y(_0648_),
    .B1(_0644_));
 sg13g2_o21ai_1 _3844_ (.B1(_0645_),
    .Y(_0649_),
    .A1(_0639_),
    .A2(_0641_));
 sg13g2_a21oi_1 _3845_ (.A1(net553),
    .A2(\load_weights[197] ),
    .Y(_0650_),
    .B1(\load_weights[209] ));
 sg13g2_a21oi_1 _3846_ (.A1(net553),
    .A2(\load_weights[209] ),
    .Y(_0651_),
    .B1(_0650_));
 sg13g2_a21o_1 _3847_ (.A2(\load_weights[209] ),
    .A1(net553),
    .B1(_0650_),
    .X(_0652_));
 sg13g2_nor3_1 _3848_ (.A(_0646_),
    .B(_0648_),
    .C(_0652_),
    .Y(_0653_));
 sg13g2_nand3_1 _3849_ (.B(_0649_),
    .C(_0651_),
    .A(_0647_),
    .Y(_0654_));
 sg13g2_a21oi_1 _3850_ (.A1(_0647_),
    .A2(_0649_),
    .Y(_0655_),
    .B1(_0651_));
 sg13g2_o21ai_1 _3851_ (.B1(_0652_),
    .Y(_0656_),
    .A1(_0646_),
    .A2(_0648_));
 sg13g2_a21oi_1 _3852_ (.A1(net522),
    .A2(\load_weights[192] ),
    .Y(_0657_),
    .B1(\load_weights[204] ));
 sg13g2_a21o_1 _3853_ (.A2(\load_weights[204] ),
    .A1(net522),
    .B1(_0657_),
    .X(_0658_));
 sg13g2_inv_1 _3854_ (.Y(_0659_),
    .A(_0658_));
 sg13g2_nor3_1 _3855_ (.A(_0653_),
    .B(_0655_),
    .C(_0658_),
    .Y(_0660_));
 sg13g2_a21oi_1 _3856_ (.A1(_0654_),
    .A2(_0656_),
    .Y(_0661_),
    .B1(_0659_));
 sg13g2_nand3_1 _3857_ (.B(_0656_),
    .C(_0658_),
    .A(_0654_),
    .Y(_0662_));
 sg13g2_o21ai_1 _3858_ (.B1(_0659_),
    .Y(_0663_),
    .A1(_0653_),
    .A2(_0655_));
 sg13g2_a21oi_1 _3859_ (.A1(net544),
    .A2(\load_weights[199] ),
    .Y(_0664_),
    .B1(\load_weights[211] ));
 sg13g2_a21o_1 _3860_ (.A2(\load_weights[211] ),
    .A1(net544),
    .B1(_0664_),
    .X(_0665_));
 sg13g2_nor3_1 _3861_ (.A(_0660_),
    .B(_0661_),
    .C(_0665_),
    .Y(_0666_));
 sg13g2_and3_1 _3862_ (.X(_0667_),
    .A(_0662_),
    .B(_0663_),
    .C(_0665_));
 sg13g2_o21ai_1 _3863_ (.B1(_0665_),
    .Y(_0668_),
    .A1(_0660_),
    .A2(_0661_));
 sg13g2_a21oi_1 _3864_ (.A1(net538),
    .A2(net797),
    .Y(_0669_),
    .B1(net820));
 sg13g2_a21oi_1 _3865_ (.A1(net536),
    .A2(net932),
    .Y(_0670_),
    .B1(_0669_));
 sg13g2_nor3_1 _3866_ (.A(_0666_),
    .B(_0667_),
    .C(_0670_),
    .Y(_0671_));
 sg13g2_o21ai_1 _3867_ (.B1(_0670_),
    .Y(_0672_),
    .A1(_0666_),
    .A2(_0667_));
 sg13g2_nand2b_1 _3868_ (.Y(\tt_um_mult_inst.genblk1[8].out_q ),
    .B(_0672_),
    .A_N(_0671_));
 sg13g2_a21oi_1 _3869_ (.A1(_0668_),
    .A2(_0670_),
    .Y(_0673_),
    .B1(_0666_));
 sg13g2_o21ai_1 _3870_ (.B1(_0589_),
    .Y(_0674_),
    .A1(_0583_),
    .A2(_0585_));
 sg13g2_nand2b_1 _3871_ (.Y(_0675_),
    .B(_0633_),
    .A_N(_0628_));
 sg13g2_o21ai_1 _3872_ (.B1(_0600_),
    .Y(_0676_),
    .A1(_0593_),
    .A2(_0595_));
 sg13g2_nor2_1 _3873_ (.A(\tt_um_mult_inst.genblk1[8].carry[1] ),
    .B(net436),
    .Y(_0677_));
 sg13g2_nand2_1 _3874_ (.Y(_0678_),
    .A(_0621_),
    .B(_0624_));
 sg13g2_a21oi_1 _3875_ (.A1(\load_weights[215] ),
    .A2(_0614_),
    .Y(_0679_),
    .B1(_0613_));
 sg13g2_a21oi_1 _3876_ (.A1(\load_weights[209] ),
    .A2(_0609_),
    .Y(_0680_),
    .B1(_0608_));
 sg13g2_nor2_1 _3877_ (.A(_0606_),
    .B(_0680_),
    .Y(_0681_));
 sg13g2_xnor2_1 _3878_ (.Y(_0682_),
    .A(_0606_),
    .B(_0680_));
 sg13g2_nor2_1 _3879_ (.A(_0611_),
    .B(_0616_),
    .Y(_0683_));
 sg13g2_nor2_1 _3880_ (.A(_0682_),
    .B(_0683_),
    .Y(_0684_));
 sg13g2_xnor2_1 _3881_ (.Y(_0685_),
    .A(_0682_),
    .B(_0683_));
 sg13g2_nor2_1 _3882_ (.A(_0679_),
    .B(_0685_),
    .Y(_0686_));
 sg13g2_xor2_1 _3883_ (.B(_0685_),
    .A(_0679_),
    .X(_0687_));
 sg13g2_o21ai_1 _3884_ (.B1(_0618_),
    .Y(_0688_),
    .A1(_1936_),
    .A2(_0619_));
 sg13g2_and2_1 _3885_ (.A(_0687_),
    .B(_0688_),
    .X(_0689_));
 sg13g2_xor2_1 _3886_ (.B(_0688_),
    .A(_0687_),
    .X(_0690_));
 sg13g2_xnor2_1 _3887_ (.Y(_0691_),
    .A(_0678_),
    .B(_0690_));
 sg13g2_a21oi_1 _3888_ (.A1(net435),
    .A2(_0691_),
    .Y(_0692_),
    .B1(_0677_));
 sg13g2_nand2_1 _3889_ (.Y(_0693_),
    .A(_0676_),
    .B(_0692_));
 sg13g2_xor2_1 _3890_ (.B(_0692_),
    .A(_0676_),
    .X(_0694_));
 sg13g2_nand2_1 _3891_ (.Y(_0695_),
    .A(_0675_),
    .B(_0694_));
 sg13g2_xnor2_1 _3892_ (.Y(_0696_),
    .A(_0675_),
    .B(_0694_));
 sg13g2_nand2b_1 _3893_ (.Y(_0697_),
    .B(_0674_),
    .A_N(_0696_));
 sg13g2_xor2_1 _3894_ (.B(_0696_),
    .A(_0674_),
    .X(_0698_));
 sg13g2_nand2_1 _3895_ (.Y(_0699_),
    .A(_0640_),
    .B(_0647_));
 sg13g2_nand2b_1 _3896_ (.Y(_0700_),
    .B(_0699_),
    .A_N(_0698_));
 sg13g2_xnor2_1 _3897_ (.Y(_0701_),
    .A(_0698_),
    .B(_0699_));
 sg13g2_o21ai_1 _3898_ (.B1(_0654_),
    .Y(_0702_),
    .A1(_0655_),
    .A2(_0658_));
 sg13g2_nand2_1 _3899_ (.Y(_0703_),
    .A(_0701_),
    .B(_0702_));
 sg13g2_xnor2_1 _3900_ (.Y(_0704_),
    .A(_0701_),
    .B(_0702_));
 sg13g2_xor2_1 _3901_ (.B(_0704_),
    .A(_0673_),
    .X(\tt_um_mult_inst.genblk1[8].carry_q[0] ));
 sg13g2_o21ai_1 _3902_ (.B1(_0703_),
    .Y(_0705_),
    .A1(_0673_),
    .A2(_0704_));
 sg13g2_nand2_1 _3903_ (.Y(_0706_),
    .A(_0681_),
    .B(_0686_));
 sg13g2_nor3_1 _3904_ (.A(_0681_),
    .B(_0684_),
    .C(_0686_),
    .Y(_0707_));
 sg13g2_a21oi_1 _3905_ (.A1(_0681_),
    .A2(_0686_),
    .Y(_0708_),
    .B1(_0707_));
 sg13g2_a21o_1 _3906_ (.A2(_0690_),
    .A1(_0678_),
    .B1(_0689_),
    .X(_0709_));
 sg13g2_or2_1 _3907_ (.X(_0710_),
    .B(_0709_),
    .A(_0708_));
 sg13g2_a21oi_1 _3908_ (.A1(_0708_),
    .A2(_0709_),
    .Y(_0711_),
    .B1(net431));
 sg13g2_a22oi_1 _3909_ (.Y(_0712_),
    .B1(_0710_),
    .B2(_0711_),
    .A2(net428),
    .A1(\tt_um_mult_inst.genblk1[8].carry[2] ));
 sg13g2_xnor2_1 _3910_ (.Y(_0713_),
    .A(_0693_),
    .B(_0712_));
 sg13g2_a21o_1 _3911_ (.A2(_0697_),
    .A1(_0695_),
    .B1(_0713_),
    .X(_0714_));
 sg13g2_nand3_1 _3912_ (.B(_0697_),
    .C(_0713_),
    .A(_0695_),
    .Y(_0715_));
 sg13g2_nand2_1 _3913_ (.Y(_0716_),
    .A(_0714_),
    .B(_0715_));
 sg13g2_nor2_1 _3914_ (.A(_0700_),
    .B(_0716_),
    .Y(_0717_));
 sg13g2_xor2_1 _3915_ (.B(_0716_),
    .A(_0700_),
    .X(_0718_));
 sg13g2_xor2_1 _3916_ (.B(_0718_),
    .A(_0705_),
    .X(\tt_um_mult_inst.genblk1[8].carry_q[1] ));
 sg13g2_a21oi_2 _3917_ (.B1(_0717_),
    .Y(_0719_),
    .A2(_0718_),
    .A1(_0705_));
 sg13g2_a22oi_1 _3918_ (.Y(_0720_),
    .B1(_0706_),
    .B2(_0711_),
    .A2(net428),
    .A1(net916));
 sg13g2_o21ai_1 _3919_ (.B1(_0714_),
    .Y(_0721_),
    .A1(_0693_),
    .A2(_0712_));
 sg13g2_xor2_1 _3920_ (.B(_0721_),
    .A(_0720_),
    .X(_0722_));
 sg13g2_nor2b_1 _3921_ (.A(_0719_),
    .B_N(_0722_),
    .Y(_0723_));
 sg13g2_xnor2_1 _3922_ (.Y(\tt_um_mult_inst.genblk1[8].carry_q[2] ),
    .A(_0719_),
    .B(_0722_));
 sg13g2_a21o_1 _3923_ (.A2(_0721_),
    .A1(_0720_),
    .B1(_0723_),
    .X(\tt_um_mult_inst.genblk1[8].carry_q[3] ));
 sg13g2_a21oi_1 _3924_ (.A1(net548),
    .A2(\load_weights[150] ),
    .Y(_0724_),
    .B1(\load_weights[162] ));
 sg13g2_a21o_1 _3925_ (.A2(\load_weights[162] ),
    .A1(net548),
    .B1(_0724_),
    .X(_0725_));
 sg13g2_a21oi_1 _3926_ (.A1(net558),
    .A2(\load_weights[148] ),
    .Y(_0726_),
    .B1(\load_weights[160] ));
 sg13g2_a21o_1 _3927_ (.A2(\load_weights[160] ),
    .A1(net559),
    .B1(_0726_),
    .X(_0727_));
 sg13g2_xor2_1 _3928_ (.B(_0727_),
    .A(_0725_),
    .X(_0728_));
 sg13g2_a21oi_1 _3929_ (.A1(net512),
    .A2(\load_weights[146] ),
    .Y(_0729_),
    .B1(\load_weights[158] ));
 sg13g2_a21oi_1 _3930_ (.A1(net512),
    .A2(\load_weights[158] ),
    .Y(_0730_),
    .B1(_0729_));
 sg13g2_nand2_1 _3931_ (.Y(_0731_),
    .A(_0728_),
    .B(_0730_));
 sg13g2_xnor2_1 _3932_ (.Y(_0732_),
    .A(_0728_),
    .B(_0730_));
 sg13g2_inv_1 _3933_ (.Y(_0733_),
    .A(_0732_));
 sg13g2_a21oi_1 _3934_ (.A1(net527),
    .A2(\load_weights[155] ),
    .Y(_0734_),
    .B1(\load_weights[167] ));
 sg13g2_a21o_2 _3935_ (.A2(\load_weights[167] ),
    .A1(net527),
    .B1(_0734_),
    .X(_0735_));
 sg13g2_a21oi_1 _3936_ (.A1(net531),
    .A2(\load_weights[154] ),
    .Y(_0736_),
    .B1(\load_weights[166] ));
 sg13g2_a21o_1 _3937_ (.A2(\load_weights[166] ),
    .A1(net531),
    .B1(_0736_),
    .X(_0737_));
 sg13g2_xor2_1 _3938_ (.B(_0737_),
    .A(_0735_),
    .X(_0738_));
 sg13g2_a21oi_1 _3939_ (.A1(net539),
    .A2(\load_weights[152] ),
    .Y(_0739_),
    .B1(\load_weights[164] ));
 sg13g2_a21o_1 _3940_ (.A2(\load_weights[164] ),
    .A1(net539),
    .B1(_0739_),
    .X(_0740_));
 sg13g2_inv_1 _3941_ (.Y(_0741_),
    .A(_0740_));
 sg13g2_nand2_1 _3942_ (.Y(_0742_),
    .A(_0738_),
    .B(_0741_));
 sg13g2_nand2b_1 _3943_ (.Y(_0743_),
    .B(_0740_),
    .A_N(_0738_));
 sg13g2_nand2_1 _3944_ (.Y(_0744_),
    .A(_0742_),
    .B(_0743_));
 sg13g2_nand2_1 _3945_ (.Y(_0745_),
    .A(\load_weights[156] ),
    .B(\load_weights[157] ));
 sg13g2_xnor2_1 _3946_ (.Y(_0746_),
    .A(\load_weights[156] ),
    .B(\load_weights[157] ));
 sg13g2_and2_1 _3947_ (.A(\load_weights[158] ),
    .B(\load_weights[159] ),
    .X(_0747_));
 sg13g2_xor2_1 _3948_ (.B(\load_weights[159] ),
    .A(\load_weights[158] ),
    .X(_0748_));
 sg13g2_xnor2_1 _3949_ (.Y(_0749_),
    .A(\load_weights[161] ),
    .B(_0748_));
 sg13g2_nor2_1 _3950_ (.A(_0746_),
    .B(_0749_),
    .Y(_0750_));
 sg13g2_xnor2_1 _3951_ (.Y(_0751_),
    .A(_0746_),
    .B(_0749_));
 sg13g2_and2_1 _3952_ (.A(\load_weights[163] ),
    .B(\load_weights[165] ),
    .X(_0752_));
 sg13g2_xor2_1 _3953_ (.B(\load_weights[165] ),
    .A(\load_weights[163] ),
    .X(_0753_));
 sg13g2_xnor2_1 _3954_ (.Y(_0754_),
    .A(\load_weights[167] ),
    .B(_0753_));
 sg13g2_nor2_1 _3955_ (.A(_0751_),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_xor2_1 _3956_ (.B(_0754_),
    .A(_0751_),
    .X(_0756_));
 sg13g2_nand2_1 _3957_ (.Y(_0757_),
    .A(\load_weights[164] ),
    .B(_0756_));
 sg13g2_xnor2_1 _3958_ (.Y(_0758_),
    .A(\load_weights[164] ),
    .B(_0756_));
 sg13g2_xnor2_1 _3959_ (.Y(_0759_),
    .A(\load_weights[166] ),
    .B(_0758_));
 sg13g2_nand2_1 _3960_ (.Y(_0760_),
    .A(\load_weights[162] ),
    .B(_0759_));
 sg13g2_xor2_1 _3961_ (.B(_0759_),
    .A(\load_weights[162] ),
    .X(_0761_));
 sg13g2_nand2_1 _3962_ (.Y(_0762_),
    .A(\load_weights[160] ),
    .B(_0761_));
 sg13g2_nor2_1 _3963_ (.A(\load_weights[160] ),
    .B(_0761_),
    .Y(_0763_));
 sg13g2_nor2_1 _3964_ (.A(net424),
    .B(_0763_),
    .Y(_0764_));
 sg13g2_xnor2_1 _3965_ (.Y(_0765_),
    .A(\load_weights[160] ),
    .B(_0761_));
 sg13g2_nor2_1 _3966_ (.A(_1941_),
    .B(net437),
    .Y(_0766_));
 sg13g2_a21oi_1 _3967_ (.A1(net437),
    .A2(_0765_),
    .Y(_0767_),
    .B1(_0766_));
 sg13g2_nor2b_1 _3968_ (.A(_0744_),
    .B_N(_0767_),
    .Y(_0768_));
 sg13g2_nor2b_1 _3969_ (.A(_0767_),
    .B_N(_0744_),
    .Y(_0769_));
 sg13g2_a221oi_1 _3970_ (.B2(_0764_),
    .C1(_0744_),
    .B1(_0762_),
    .A1(_1941_),
    .Y(_0770_),
    .A2(net424));
 sg13g2_a221oi_1 _3971_ (.B2(net437),
    .C1(_0766_),
    .B1(_0765_),
    .A1(_0742_),
    .Y(_0771_),
    .A2(_0743_));
 sg13g2_nor3_2 _3972_ (.A(_0732_),
    .B(_0768_),
    .C(_0769_),
    .Y(_0772_));
 sg13g2_o21ai_1 _3973_ (.B1(_0733_),
    .Y(_0773_),
    .A1(_0770_),
    .A2(_0771_));
 sg13g2_nor3_2 _3974_ (.A(_0733_),
    .B(_0770_),
    .C(_0771_),
    .Y(_0774_));
 sg13g2_o21ai_1 _3975_ (.B1(_0732_),
    .Y(_0775_),
    .A1(_0768_),
    .A2(_0769_));
 sg13g2_a21oi_1 _3976_ (.A1(net506),
    .A2(\load_weights[147] ),
    .Y(_0776_),
    .B1(\load_weights[159] ));
 sg13g2_a21oi_1 _3977_ (.A1(net506),
    .A2(\load_weights[159] ),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_a21o_1 _3978_ (.A2(\load_weights[159] ),
    .A1(net506),
    .B1(_0776_),
    .X(_0778_));
 sg13g2_nor3_1 _3979_ (.A(_0772_),
    .B(_0774_),
    .C(_0778_),
    .Y(_0779_));
 sg13g2_nand3_1 _3980_ (.B(_0775_),
    .C(_0777_),
    .A(_0773_),
    .Y(_0780_));
 sg13g2_a21oi_1 _3981_ (.A1(_0773_),
    .A2(_0775_),
    .Y(_0781_),
    .B1(_0777_));
 sg13g2_o21ai_1 _3982_ (.B1(_0778_),
    .Y(_0782_),
    .A1(_0772_),
    .A2(_0774_));
 sg13g2_a21oi_1 _3983_ (.A1(net516),
    .A2(\load_weights[145] ),
    .Y(_0783_),
    .B1(\load_weights[157] ));
 sg13g2_a21oi_1 _3984_ (.A1(net517),
    .A2(\load_weights[157] ),
    .Y(_0784_),
    .B1(_0783_));
 sg13g2_a21o_1 _3985_ (.A2(\load_weights[157] ),
    .A1(net516),
    .B1(_0783_),
    .X(_0785_));
 sg13g2_nor3_1 _3986_ (.A(_0779_),
    .B(_0781_),
    .C(_0785_),
    .Y(_0786_));
 sg13g2_nand3_1 _3987_ (.B(_0782_),
    .C(_0784_),
    .A(_0780_),
    .Y(_0787_));
 sg13g2_a21oi_1 _3988_ (.A1(_0780_),
    .A2(_0782_),
    .Y(_0788_),
    .B1(_0784_));
 sg13g2_o21ai_1 _3989_ (.B1(_0785_),
    .Y(_0789_),
    .A1(_0779_),
    .A2(_0781_));
 sg13g2_a21oi_1 _3990_ (.A1(net553),
    .A2(\load_weights[149] ),
    .Y(_0790_),
    .B1(\load_weights[161] ));
 sg13g2_a21oi_1 _3991_ (.A1(net553),
    .A2(\load_weights[161] ),
    .Y(_0791_),
    .B1(_0790_));
 sg13g2_a21o_1 _3992_ (.A2(\load_weights[161] ),
    .A1(net553),
    .B1(_0790_),
    .X(_0792_));
 sg13g2_nor3_1 _3993_ (.A(_0786_),
    .B(_0788_),
    .C(_0792_),
    .Y(_0793_));
 sg13g2_nand3_1 _3994_ (.B(_0789_),
    .C(_0791_),
    .A(_0787_),
    .Y(_0794_));
 sg13g2_a21oi_1 _3995_ (.A1(_0787_),
    .A2(_0789_),
    .Y(_0795_),
    .B1(_0791_));
 sg13g2_o21ai_1 _3996_ (.B1(_0792_),
    .Y(_0796_),
    .A1(_0786_),
    .A2(_0788_));
 sg13g2_a21oi_1 _3997_ (.A1(net521),
    .A2(\load_weights[144] ),
    .Y(_0797_),
    .B1(\load_weights[156] ));
 sg13g2_a21o_2 _3998_ (.A2(\load_weights[156] ),
    .A1(net521),
    .B1(_0797_),
    .X(_0798_));
 sg13g2_inv_1 _3999_ (.Y(_0799_),
    .A(_0798_));
 sg13g2_nor3_1 _4000_ (.A(_0793_),
    .B(_0795_),
    .C(_0798_),
    .Y(_0800_));
 sg13g2_a21oi_1 _4001_ (.A1(_0794_),
    .A2(_0796_),
    .Y(_0801_),
    .B1(_0799_));
 sg13g2_nand3_1 _4002_ (.B(_0796_),
    .C(_0798_),
    .A(_0794_),
    .Y(_0802_));
 sg13g2_o21ai_1 _4003_ (.B1(_0799_),
    .Y(_0803_),
    .A1(_0793_),
    .A2(_0795_));
 sg13g2_a21oi_1 _4004_ (.A1(net544),
    .A2(\load_weights[151] ),
    .Y(_0804_),
    .B1(\load_weights[163] ));
 sg13g2_a21o_1 _4005_ (.A2(\load_weights[163] ),
    .A1(net544),
    .B1(_0804_),
    .X(_0805_));
 sg13g2_nor3_2 _4006_ (.A(_0800_),
    .B(_0801_),
    .C(_0805_),
    .Y(_0806_));
 sg13g2_and3_1 _4007_ (.X(_0807_),
    .A(_0802_),
    .B(_0803_),
    .C(_0805_));
 sg13g2_o21ai_1 _4008_ (.B1(_0805_),
    .Y(_0808_),
    .A1(_0800_),
    .A2(_0801_));
 sg13g2_a21oi_1 _4009_ (.A1(net536),
    .A2(\load_weights[153] ),
    .Y(_0809_),
    .B1(\load_weights[165] ));
 sg13g2_a21oi_2 _4010_ (.B1(_0809_),
    .Y(_0810_),
    .A2(\load_weights[165] ),
    .A1(net536));
 sg13g2_nor3_1 _4011_ (.A(_0806_),
    .B(_0807_),
    .C(_0810_),
    .Y(_0811_));
 sg13g2_o21ai_1 _4012_ (.B1(_0810_),
    .Y(_0812_),
    .A1(_0806_),
    .A2(_0807_));
 sg13g2_nand2b_2 _4013_ (.Y(\tt_um_mult_inst.genblk1[6].out_q ),
    .B(_0812_),
    .A_N(_0811_));
 sg13g2_a21oi_2 _4014_ (.B1(_0806_),
    .Y(_0813_),
    .A2(_0810_),
    .A1(_0808_));
 sg13g2_o21ai_1 _4015_ (.B1(_0731_),
    .Y(_0814_),
    .A1(_0725_),
    .A2(_0727_));
 sg13g2_nand2b_1 _4016_ (.Y(_0815_),
    .B(_0773_),
    .A_N(_0768_));
 sg13g2_o21ai_1 _4017_ (.B1(_0742_),
    .Y(_0816_),
    .A1(_0735_),
    .A2(_0737_));
 sg13g2_nor2_1 _4018_ (.A(\tt_um_mult_inst.genblk1[6].carry[1] ),
    .B(net437),
    .Y(_0817_));
 sg13g2_nand2_1 _4019_ (.Y(_0818_),
    .A(_0760_),
    .B(_0762_));
 sg13g2_a21oi_2 _4020_ (.B1(_0752_),
    .Y(_0819_),
    .A2(_0753_),
    .A1(\load_weights[167] ));
 sg13g2_a21oi_1 _4021_ (.A1(\load_weights[161] ),
    .A2(_0748_),
    .Y(_0820_),
    .B1(_0747_));
 sg13g2_nor2_1 _4022_ (.A(_0745_),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_xnor2_1 _4023_ (.Y(_0822_),
    .A(_0745_),
    .B(_0820_));
 sg13g2_nor2_1 _4024_ (.A(_0750_),
    .B(_0755_),
    .Y(_0823_));
 sg13g2_nor2_1 _4025_ (.A(_0822_),
    .B(_0823_),
    .Y(_0824_));
 sg13g2_xnor2_1 _4026_ (.Y(_0825_),
    .A(_0822_),
    .B(_0823_));
 sg13g2_nor2_1 _4027_ (.A(_0819_),
    .B(_0825_),
    .Y(_0826_));
 sg13g2_xor2_1 _4028_ (.B(_0825_),
    .A(_0819_),
    .X(_0827_));
 sg13g2_o21ai_1 _4029_ (.B1(_0757_),
    .Y(_0828_),
    .A1(_1939_),
    .A2(_0758_));
 sg13g2_and2_1 _4030_ (.A(_0827_),
    .B(_0828_),
    .X(_0829_));
 sg13g2_xor2_1 _4031_ (.B(_0828_),
    .A(_0827_),
    .X(_0830_));
 sg13g2_xnor2_1 _4032_ (.Y(_0831_),
    .A(_0818_),
    .B(_0830_));
 sg13g2_a21oi_1 _4033_ (.A1(net437),
    .A2(_0831_),
    .Y(_0832_),
    .B1(_0817_));
 sg13g2_nand2_1 _4034_ (.Y(_0833_),
    .A(_0816_),
    .B(_0832_));
 sg13g2_xor2_1 _4035_ (.B(_0832_),
    .A(_0816_),
    .X(_0834_));
 sg13g2_nand2_1 _4036_ (.Y(_0835_),
    .A(_0815_),
    .B(_0834_));
 sg13g2_xnor2_1 _4037_ (.Y(_0836_),
    .A(_0815_),
    .B(_0834_));
 sg13g2_nand2b_1 _4038_ (.Y(_0837_),
    .B(_0814_),
    .A_N(_0836_));
 sg13g2_xor2_1 _4039_ (.B(_0836_),
    .A(_0814_),
    .X(_0838_));
 sg13g2_nand2_1 _4040_ (.Y(_0839_),
    .A(_0780_),
    .B(_0787_));
 sg13g2_nand2b_1 _4041_ (.Y(_0840_),
    .B(_0839_),
    .A_N(_0838_));
 sg13g2_xnor2_1 _4042_ (.Y(_0841_),
    .A(_0838_),
    .B(_0839_));
 sg13g2_o21ai_1 _4043_ (.B1(_0794_),
    .Y(_0842_),
    .A1(_0795_),
    .A2(_0798_));
 sg13g2_nand2_1 _4044_ (.Y(_0843_),
    .A(_0841_),
    .B(_0842_));
 sg13g2_xnor2_1 _4045_ (.Y(_0844_),
    .A(_0841_),
    .B(_0842_));
 sg13g2_xor2_1 _4046_ (.B(_0844_),
    .A(_0813_),
    .X(\tt_um_mult_inst.genblk1[6].carry_q[0] ));
 sg13g2_o21ai_1 _4047_ (.B1(_0843_),
    .Y(_0845_),
    .A1(_0813_),
    .A2(_0844_));
 sg13g2_nand2_1 _4048_ (.Y(_0846_),
    .A(_0821_),
    .B(_0826_));
 sg13g2_nor3_1 _4049_ (.A(_0821_),
    .B(_0824_),
    .C(_0826_),
    .Y(_0847_));
 sg13g2_a21oi_1 _4050_ (.A1(_0821_),
    .A2(_0826_),
    .Y(_0848_),
    .B1(_0847_));
 sg13g2_a21o_1 _4051_ (.A2(_0830_),
    .A1(_0818_),
    .B1(_0829_),
    .X(_0849_));
 sg13g2_or2_1 _4052_ (.X(_0850_),
    .B(_0849_),
    .A(_0848_));
 sg13g2_a21oi_1 _4053_ (.A1(_0848_),
    .A2(_0849_),
    .Y(_0851_),
    .B1(net424));
 sg13g2_a22oi_1 _4054_ (.Y(_0852_),
    .B1(_0850_),
    .B2(_0851_),
    .A2(net424),
    .A1(\tt_um_mult_inst.genblk1[6].carry[2] ));
 sg13g2_xnor2_1 _4055_ (.Y(_0853_),
    .A(_0833_),
    .B(_0852_));
 sg13g2_a21o_1 _4056_ (.A2(_0837_),
    .A1(_0835_),
    .B1(_0853_),
    .X(_0854_));
 sg13g2_nand3_1 _4057_ (.B(_0837_),
    .C(_0853_),
    .A(_0835_),
    .Y(_0855_));
 sg13g2_nand2_1 _4058_ (.Y(_0856_),
    .A(_0854_),
    .B(_0855_));
 sg13g2_nor2_1 _4059_ (.A(_0840_),
    .B(_0856_),
    .Y(_0857_));
 sg13g2_xor2_1 _4060_ (.B(_0856_),
    .A(_0840_),
    .X(_0858_));
 sg13g2_xor2_1 _4061_ (.B(_0858_),
    .A(_0845_),
    .X(\tt_um_mult_inst.genblk1[6].carry_q[1] ));
 sg13g2_a21oi_1 _4062_ (.A1(_0845_),
    .A2(_0858_),
    .Y(_0859_),
    .B1(_0857_));
 sg13g2_a22oi_1 _4063_ (.Y(_0860_),
    .B1(_0846_),
    .B2(_0851_),
    .A2(net424),
    .A1(net907));
 sg13g2_o21ai_1 _4064_ (.B1(_0854_),
    .Y(_0861_),
    .A1(_0833_),
    .A2(_0852_));
 sg13g2_xnor2_1 _4065_ (.Y(_0862_),
    .A(_0860_),
    .B(_0861_));
 sg13g2_xor2_1 _4066_ (.B(_0862_),
    .A(_0859_),
    .X(\tt_um_mult_inst.genblk1[6].carry_q[2] ));
 sg13g2_nand2_1 _4067_ (.Y(_0863_),
    .A(_0860_),
    .B(_0861_));
 sg13g2_o21ai_1 _4068_ (.B1(_0863_),
    .Y(\tt_um_mult_inst.genblk1[6].carry_q[3] ),
    .A1(_0859_),
    .A2(_0862_));
 sg13g2_a21oi_1 _4069_ (.A1(net530),
    .A2(\load_weights[82] ),
    .Y(_0864_),
    .B1(\load_weights[94] ));
 sg13g2_a21o_1 _4070_ (.A2(\load_weights[94] ),
    .A1(net530),
    .B1(_0864_),
    .X(_0865_));
 sg13g2_a21oi_1 _4071_ (.A1(net540),
    .A2(\load_weights[80] ),
    .Y(_0866_),
    .B1(\load_weights[92] ));
 sg13g2_a21o_1 _4072_ (.A2(\load_weights[92] ),
    .A1(net540),
    .B1(_0866_),
    .X(_0867_));
 sg13g2_xor2_1 _4073_ (.B(_0867_),
    .A(_0865_),
    .X(_0868_));
 sg13g2_a21oi_1 _4074_ (.A1(net554),
    .A2(\load_weights[77] ),
    .Y(_0869_),
    .B1(\load_weights[89] ));
 sg13g2_a21oi_1 _4075_ (.A1(net554),
    .A2(\load_weights[89] ),
    .Y(_0870_),
    .B1(_0869_));
 sg13g2_nand2_1 _4076_ (.Y(_0871_),
    .A(_0868_),
    .B(_0870_));
 sg13g2_xnor2_1 _4077_ (.Y(_0872_),
    .A(_0868_),
    .B(_0870_));
 sg13g2_inv_1 _4078_ (.Y(_0873_),
    .A(_0872_));
 sg13g2_a21oi_1 _4079_ (.A1(net511),
    .A2(\load_weights[74] ),
    .Y(_0874_),
    .B1(\load_weights[86] ));
 sg13g2_a21o_1 _4080_ (.A2(\load_weights[86] ),
    .A1(net511),
    .B1(_0874_),
    .X(_0875_));
 sg13g2_a21oi_1 _4081_ (.A1(net558),
    .A2(\load_weights[76] ),
    .Y(_0876_),
    .B1(\load_weights[88] ));
 sg13g2_a21o_1 _4082_ (.A2(\load_weights[88] ),
    .A1(net558),
    .B1(_0876_),
    .X(_0877_));
 sg13g2_xor2_1 _4083_ (.B(_0877_),
    .A(_0875_),
    .X(_0878_));
 sg13g2_a21oi_1 _4084_ (.A1(net520),
    .A2(\load_weights[73] ),
    .Y(_0879_),
    .B1(\load_weights[85] ));
 sg13g2_a21o_1 _4085_ (.A2(\load_weights[85] ),
    .A1(net520),
    .B1(_0879_),
    .X(_0880_));
 sg13g2_inv_1 _4086_ (.Y(_0881_),
    .A(_0880_));
 sg13g2_nand2_1 _4087_ (.Y(_0882_),
    .A(_0878_),
    .B(_0881_));
 sg13g2_nand2b_1 _4088_ (.Y(_0883_),
    .B(_0880_),
    .A_N(_0878_));
 sg13g2_nand2_1 _4089_ (.Y(_0884_),
    .A(_0878_),
    .B(_0880_));
 sg13g2_nand2b_1 _4090_ (.Y(_0885_),
    .B(_0881_),
    .A_N(_0878_));
 sg13g2_nand2_1 _4091_ (.Y(_0886_),
    .A(_0882_),
    .B(_0883_));
 sg13g2_inv_1 _4092_ (.Y(_0887_),
    .A(_0886_));
 sg13g2_and2_1 _4093_ (.A(\load_weights[85] ),
    .B(\load_weights[84] ),
    .X(_0888_));
 sg13g2_xor2_1 _4094_ (.B(\load_weights[84] ),
    .A(\load_weights[85] ),
    .X(_0889_));
 sg13g2_xnor2_1 _4095_ (.Y(_0890_),
    .A(\load_weights[86] ),
    .B(_0889_));
 sg13g2_inv_1 _4096_ (.Y(_0891_),
    .A(_0890_));
 sg13g2_nand2_1 _4097_ (.Y(_0892_),
    .A(\load_weights[88] ),
    .B(_0891_));
 sg13g2_xor2_1 _4098_ (.B(_0890_),
    .A(\load_weights[88] ),
    .X(_0893_));
 sg13g2_xor2_1 _4099_ (.B(_0893_),
    .A(_0004_),
    .X(_0894_));
 sg13g2_and2_1 _4100_ (.A(\load_weights[90] ),
    .B(\load_weights[92] ),
    .X(_0895_));
 sg13g2_xor2_1 _4101_ (.B(\load_weights[92] ),
    .A(\load_weights[90] ),
    .X(_0896_));
 sg13g2_xor2_1 _4102_ (.B(_0896_),
    .A(\load_weights[94] ),
    .X(_0897_));
 sg13g2_nand2_1 _4103_ (.Y(_0898_),
    .A(_0894_),
    .B(_0897_));
 sg13g2_xnor2_1 _4104_ (.Y(_0899_),
    .A(_0894_),
    .B(_0897_));
 sg13g2_inv_1 _4105_ (.Y(_0900_),
    .A(_0899_));
 sg13g2_xor2_1 _4106_ (.B(_0899_),
    .A(\load_weights[91] ),
    .X(_0901_));
 sg13g2_nor2_1 _4107_ (.A(_1942_),
    .B(_0901_),
    .Y(_0902_));
 sg13g2_xnor2_1 _4108_ (.Y(_0903_),
    .A(\load_weights[93] ),
    .B(_0901_));
 sg13g2_nand2_1 _4109_ (.Y(_0904_),
    .A(\load_weights[89] ),
    .B(_0903_));
 sg13g2_xor2_1 _4110_ (.B(_0903_),
    .A(\load_weights[89] ),
    .X(_0905_));
 sg13g2_xnor2_1 _4111_ (.Y(_0906_),
    .A(\load_weights[89] ),
    .B(_0903_));
 sg13g2_nand2_1 _4112_ (.Y(_0907_),
    .A(\load_weights[87] ),
    .B(_0905_));
 sg13g2_a21oi_1 _4113_ (.A1(_1943_),
    .A2(_0906_),
    .Y(_0908_),
    .B1(net423));
 sg13g2_xnor2_1 _4114_ (.Y(_0909_),
    .A(\load_weights[87] ),
    .B(_0905_));
 sg13g2_nor2_1 _4115_ (.A(_1944_),
    .B(net435),
    .Y(_0910_));
 sg13g2_a221oi_1 _4116_ (.B2(net435),
    .C1(_0910_),
    .B1(_0909_),
    .A1(_0884_),
    .Y(_0911_),
    .A2(_0885_));
 sg13g2_a221oi_1 _4117_ (.B2(_0908_),
    .C1(_0887_),
    .B1(_0907_),
    .A1(_1944_),
    .Y(_0912_),
    .A2(net423));
 sg13g2_a221oi_1 _4118_ (.B2(_0908_),
    .C1(_0886_),
    .B1(_0907_),
    .A1(_1944_),
    .Y(_0913_),
    .A2(net423));
 sg13g2_a221oi_1 _4119_ (.B2(net435),
    .C1(_0910_),
    .B1(_0909_),
    .A1(_0882_),
    .Y(_0914_),
    .A2(_0883_));
 sg13g2_nor3_1 _4120_ (.A(_0872_),
    .B(_0911_),
    .C(_0912_),
    .Y(_0915_));
 sg13g2_o21ai_1 _4121_ (.B1(_0873_),
    .Y(_0916_),
    .A1(_0913_),
    .A2(_0914_));
 sg13g2_nor3_1 _4122_ (.A(_0873_),
    .B(_0913_),
    .C(_0914_),
    .Y(_0917_));
 sg13g2_o21ai_1 _4123_ (.B1(_0872_),
    .Y(_0918_),
    .A1(_0911_),
    .A2(_0912_));
 sg13g2_a21oi_1 _4124_ (.A1(net549),
    .A2(\load_weights[78] ),
    .Y(_0919_),
    .B1(\load_weights[90] ));
 sg13g2_a21oi_1 _4125_ (.A1(net549),
    .A2(\load_weights[90] ),
    .Y(_0920_),
    .B1(_0919_));
 sg13g2_a21o_1 _4126_ (.A2(\load_weights[90] ),
    .A1(net549),
    .B1(_0919_),
    .X(_0921_));
 sg13g2_nor3_1 _4127_ (.A(_0915_),
    .B(_0917_),
    .C(_0921_),
    .Y(_0922_));
 sg13g2_nand3_1 _4128_ (.B(_0918_),
    .C(_0920_),
    .A(_0916_),
    .Y(_0923_));
 sg13g2_a21oi_1 _4129_ (.A1(_0916_),
    .A2(_0918_),
    .Y(_0924_),
    .B1(_0920_));
 sg13g2_o21ai_1 _4130_ (.B1(_0921_),
    .Y(_0925_),
    .A1(_0915_),
    .A2(_0917_));
 sg13g2_a21oi_1 _4131_ (.A1(net522),
    .A2(\load_weights[72] ),
    .Y(_0926_),
    .B1(\load_weights[84] ));
 sg13g2_a21oi_1 _4132_ (.A1(net522),
    .A2(\load_weights[84] ),
    .Y(_0927_),
    .B1(_0926_));
 sg13g2_a21o_1 _4133_ (.A2(\load_weights[84] ),
    .A1(net522),
    .B1(_0926_),
    .X(_0928_));
 sg13g2_nor3_1 _4134_ (.A(_0922_),
    .B(_0924_),
    .C(_0928_),
    .Y(_0929_));
 sg13g2_nand3_1 _4135_ (.B(_0925_),
    .C(_0927_),
    .A(_0923_),
    .Y(_0930_));
 sg13g2_a21oi_1 _4136_ (.A1(_0923_),
    .A2(_0925_),
    .Y(_0931_),
    .B1(_0927_));
 sg13g2_o21ai_1 _4137_ (.B1(_0928_),
    .Y(_0932_),
    .A1(_0922_),
    .A2(_0924_));
 sg13g2_a21oi_1 _4138_ (.A1(net535),
    .A2(\load_weights[81] ),
    .Y(_0933_),
    .B1(\load_weights[93] ));
 sg13g2_a21oi_1 _4139_ (.A1(net535),
    .A2(\load_weights[93] ),
    .Y(_0934_),
    .B1(_0933_));
 sg13g2_a21o_1 _4140_ (.A2(\load_weights[93] ),
    .A1(net535),
    .B1(_0933_),
    .X(_0935_));
 sg13g2_nor3_1 _4141_ (.A(_0929_),
    .B(_0931_),
    .C(_0935_),
    .Y(_0936_));
 sg13g2_nand3_1 _4142_ (.B(_0932_),
    .C(_0934_),
    .A(_0930_),
    .Y(_0937_));
 sg13g2_a21oi_1 _4143_ (.A1(_0930_),
    .A2(_0932_),
    .Y(_0938_),
    .B1(_0934_));
 sg13g2_o21ai_1 _4144_ (.B1(_0935_),
    .Y(_0939_),
    .A1(_0929_),
    .A2(_0931_));
 sg13g2_a21oi_1 _4145_ (.A1(net508),
    .A2(\load_weights[75] ),
    .Y(_0940_),
    .B1(\load_weights[87] ));
 sg13g2_a21o_1 _4146_ (.A2(\load_weights[87] ),
    .A1(net505),
    .B1(_0940_),
    .X(_0941_));
 sg13g2_inv_1 _4147_ (.Y(_0942_),
    .A(_0941_));
 sg13g2_nor3_1 _4148_ (.A(_0936_),
    .B(_0938_),
    .C(_0941_),
    .Y(_0943_));
 sg13g2_a21oi_1 _4149_ (.A1(_0937_),
    .A2(_0939_),
    .Y(_0944_),
    .B1(_0942_));
 sg13g2_nand3_1 _4150_ (.B(_0939_),
    .C(_0941_),
    .A(_0937_),
    .Y(_0945_));
 sg13g2_o21ai_1 _4151_ (.B1(_0942_),
    .Y(_0946_),
    .A1(_0936_),
    .A2(_0938_));
 sg13g2_a21oi_1 _4152_ (.A1(net526),
    .A2(\load_weights[83] ),
    .Y(_0947_),
    .B1(\load_weights[95] ));
 sg13g2_a21o_2 _4153_ (.A2(\load_weights[95] ),
    .A1(net526),
    .B1(_0947_),
    .X(_0948_));
 sg13g2_nor3_1 _4154_ (.A(_0943_),
    .B(_0944_),
    .C(_0948_),
    .Y(_0949_));
 sg13g2_and3_1 _4155_ (.X(_0950_),
    .A(_0945_),
    .B(_0946_),
    .C(_0948_));
 sg13g2_o21ai_1 _4156_ (.B1(_0948_),
    .Y(_0951_),
    .A1(_0943_),
    .A2(_0944_));
 sg13g2_a21oi_1 _4157_ (.A1(net545),
    .A2(net935),
    .Y(_0952_),
    .B1(\load_weights[91] ));
 sg13g2_a21oi_1 _4158_ (.A1(net545),
    .A2(\load_weights[91] ),
    .Y(_0953_),
    .B1(_0952_));
 sg13g2_nor3_1 _4159_ (.A(_0949_),
    .B(_0950_),
    .C(_0953_),
    .Y(_0954_));
 sg13g2_o21ai_1 _4160_ (.B1(_0953_),
    .Y(_0955_),
    .A1(_0949_),
    .A2(_0950_));
 sg13g2_nand2b_2 _4161_ (.Y(\tt_um_mult_inst.genblk1[3].out_q ),
    .B(_0955_),
    .A_N(_0954_));
 sg13g2_a21oi_1 _4162_ (.A1(_0951_),
    .A2(_0953_),
    .Y(_0956_),
    .B1(_0949_));
 sg13g2_o21ai_1 _4163_ (.B1(_0937_),
    .Y(_0957_),
    .A1(_0938_),
    .A2(_0941_));
 sg13g2_o21ai_1 _4164_ (.B1(_0871_),
    .Y(_0958_),
    .A1(_0865_),
    .A2(_0867_));
 sg13g2_nand2b_1 _4165_ (.Y(_0959_),
    .B(_0916_),
    .A_N(_0911_));
 sg13g2_o21ai_1 _4166_ (.B1(_0882_),
    .Y(_0960_),
    .A1(_0875_),
    .A2(_0877_));
 sg13g2_nor2_1 _4167_ (.A(\tt_um_mult_inst.genblk1[3].carry[1] ),
    .B(net435),
    .Y(_0961_));
 sg13g2_nand2_1 _4168_ (.Y(_0962_),
    .A(_0904_),
    .B(_0907_));
 sg13g2_a21oi_2 _4169_ (.B1(_0895_),
    .Y(_0963_),
    .A2(_0896_),
    .A1(\load_weights[94] ));
 sg13g2_and3_1 _4170_ (.X(_0964_),
    .A(\load_weights[86] ),
    .B(\load_weights[88] ),
    .C(_0888_));
 sg13g2_a21oi_1 _4171_ (.A1(\load_weights[86] ),
    .A2(_0889_),
    .Y(_0965_),
    .B1(_0888_));
 sg13g2_a21oi_1 _4172_ (.A1(_0892_),
    .A2(_0965_),
    .Y(_0966_),
    .B1(_0964_));
 sg13g2_o21ai_1 _4173_ (.B1(_0898_),
    .Y(_0967_),
    .A1(_0004_),
    .A2(_0893_));
 sg13g2_nand2_1 _4174_ (.Y(_0968_),
    .A(_0966_),
    .B(_0967_));
 sg13g2_xnor2_1 _4175_ (.Y(_0969_),
    .A(_0966_),
    .B(_0967_));
 sg13g2_xor2_1 _4176_ (.B(_0969_),
    .A(_0963_),
    .X(_0970_));
 sg13g2_a21oi_1 _4177_ (.A1(\load_weights[91] ),
    .A2(_0900_),
    .Y(_0971_),
    .B1(_0902_));
 sg13g2_nor2b_1 _4178_ (.A(_0971_),
    .B_N(_0970_),
    .Y(_0972_));
 sg13g2_xnor2_1 _4179_ (.Y(_0973_),
    .A(_0970_),
    .B(_0971_));
 sg13g2_xnor2_1 _4180_ (.Y(_0974_),
    .A(_0962_),
    .B(_0973_));
 sg13g2_a21oi_1 _4181_ (.A1(net435),
    .A2(_0974_),
    .Y(_0975_),
    .B1(_0961_));
 sg13g2_nand2_1 _4182_ (.Y(_0976_),
    .A(_0960_),
    .B(_0975_));
 sg13g2_xor2_1 _4183_ (.B(_0975_),
    .A(_0960_),
    .X(_0977_));
 sg13g2_nand2_1 _4184_ (.Y(_0978_),
    .A(_0959_),
    .B(_0977_));
 sg13g2_xnor2_1 _4185_ (.Y(_0979_),
    .A(_0959_),
    .B(_0977_));
 sg13g2_nand2b_1 _4186_ (.Y(_0980_),
    .B(_0958_),
    .A_N(_0979_));
 sg13g2_xor2_1 _4187_ (.B(_0979_),
    .A(_0958_),
    .X(_0981_));
 sg13g2_nand2_1 _4188_ (.Y(_0982_),
    .A(_0923_),
    .B(_0930_));
 sg13g2_nand2b_1 _4189_ (.Y(_0983_),
    .B(_0982_),
    .A_N(_0981_));
 sg13g2_xnor2_1 _4190_ (.Y(_0984_),
    .A(_0981_),
    .B(_0982_));
 sg13g2_nand2_1 _4191_ (.Y(_0985_),
    .A(_0957_),
    .B(_0984_));
 sg13g2_xnor2_1 _4192_ (.Y(_0986_),
    .A(_0957_),
    .B(_0984_));
 sg13g2_xor2_1 _4193_ (.B(_0986_),
    .A(_0956_),
    .X(\tt_um_mult_inst.genblk1[3].carry_q[0] ));
 sg13g2_a21o_1 _4194_ (.A2(_0973_),
    .A1(_0962_),
    .B1(_0972_),
    .X(_0987_));
 sg13g2_o21ai_1 _4195_ (.B1(_0968_),
    .Y(_0988_),
    .A1(_0963_),
    .A2(_0969_));
 sg13g2_nand2_1 _4196_ (.Y(_0989_),
    .A(_0964_),
    .B(_0988_));
 sg13g2_xor2_1 _4197_ (.B(_0988_),
    .A(_0964_),
    .X(_0990_));
 sg13g2_or2_1 _4198_ (.X(_0991_),
    .B(_0990_),
    .A(_0987_));
 sg13g2_a21oi_1 _4199_ (.A1(_0987_),
    .A2(_0990_),
    .Y(_0992_),
    .B1(net423));
 sg13g2_a22oi_1 _4200_ (.Y(_0993_),
    .B1(_0991_),
    .B2(_0992_),
    .A2(net423),
    .A1(\tt_um_mult_inst.genblk1[3].carry[2] ));
 sg13g2_nor2_1 _4201_ (.A(_0976_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_xnor2_1 _4202_ (.Y(_0995_),
    .A(_0976_),
    .B(_0993_));
 sg13g2_nand3_1 _4203_ (.B(_0980_),
    .C(_0995_),
    .A(_0978_),
    .Y(_0996_));
 sg13g2_a21o_1 _4204_ (.A2(_0980_),
    .A1(_0978_),
    .B1(_0995_),
    .X(_0997_));
 sg13g2_nand2_1 _4205_ (.Y(_0998_),
    .A(_0996_),
    .B(_0997_));
 sg13g2_nor2_1 _4206_ (.A(_0983_),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_xor2_1 _4207_ (.B(_0998_),
    .A(_0983_),
    .X(_1000_));
 sg13g2_o21ai_1 _4208_ (.B1(_0985_),
    .Y(_1001_),
    .A1(_0956_),
    .A2(_0986_));
 sg13g2_xor2_1 _4209_ (.B(_1001_),
    .A(_1000_),
    .X(\tt_um_mult_inst.genblk1[3].carry_q[1] ));
 sg13g2_a22oi_1 _4210_ (.Y(_1002_),
    .B1(_0989_),
    .B2(_0992_),
    .A2(net423),
    .A1(net924));
 sg13g2_xnor2_1 _4211_ (.Y(_1003_),
    .A(_0994_),
    .B(_1002_));
 sg13g2_nand2_1 _4212_ (.Y(_1004_),
    .A(_0997_),
    .B(_1003_));
 sg13g2_nor2_1 _4213_ (.A(_0997_),
    .B(_1003_),
    .Y(_1005_));
 sg13g2_xor2_1 _4214_ (.B(_1003_),
    .A(_0997_),
    .X(_1006_));
 sg13g2_a21oi_1 _4215_ (.A1(_1000_),
    .A2(_1001_),
    .Y(_1007_),
    .B1(_0999_));
 sg13g2_xnor2_1 _4216_ (.Y(\tt_um_mult_inst.genblk1[3].carry_q[2] ),
    .A(_1006_),
    .B(_1007_));
 sg13g2_nand3_1 _4217_ (.B(_1001_),
    .C(_1004_),
    .A(_1000_),
    .Y(_1008_));
 sg13g2_nand2_1 _4218_ (.Y(_1009_),
    .A(_0999_),
    .B(_1004_));
 sg13g2_a21oi_1 _4219_ (.A1(_0994_),
    .A2(_1002_),
    .Y(_1010_),
    .B1(_1005_));
 sg13g2_nand3_1 _4220_ (.B(_1009_),
    .C(_1010_),
    .A(_1008_),
    .Y(\tt_um_mult_inst.genblk1[3].carry_q[3] ));
 sg13g2_a21oi_1 _4221_ (.A1(net535),
    .A2(\load_weights[105] ),
    .Y(_1011_),
    .B1(\load_weights[117] ));
 sg13g2_a21o_1 _4222_ (.A2(\load_weights[117] ),
    .A1(net535),
    .B1(_1011_),
    .X(_1012_));
 sg13g2_a21oi_1 _4223_ (.A1(net549),
    .A2(\load_weights[102] ),
    .Y(_1013_),
    .B1(\load_weights[114] ));
 sg13g2_a21o_1 _4224_ (.A2(\load_weights[114] ),
    .A1(net549),
    .B1(_1013_),
    .X(_1014_));
 sg13g2_xor2_1 _4225_ (.B(_1014_),
    .A(_1012_),
    .X(_1015_));
 sg13g2_a21oi_1 _4226_ (.A1(net521),
    .A2(\load_weights[96] ),
    .Y(_1016_),
    .B1(\load_weights[108] ));
 sg13g2_a21oi_1 _4227_ (.A1(net521),
    .A2(\load_weights[108] ),
    .Y(_1017_),
    .B1(_1016_));
 sg13g2_nand2_1 _4228_ (.Y(_1018_),
    .A(_1015_),
    .B(_1017_));
 sg13g2_xnor2_1 _4229_ (.Y(_1019_),
    .A(_1015_),
    .B(_1017_));
 sg13g2_a21oi_1 _4230_ (.A1(net516),
    .A2(\load_weights[97] ),
    .Y(_1020_),
    .B1(\load_weights[109] ));
 sg13g2_a21o_1 _4231_ (.A2(\load_weights[109] ),
    .A1(net516),
    .B1(_1020_),
    .X(_1021_));
 sg13g2_a21oi_1 _4232_ (.A1(net554),
    .A2(\load_weights[101] ),
    .Y(_1022_),
    .B1(\load_weights[113] ));
 sg13g2_a21o_1 _4233_ (.A2(\load_weights[113] ),
    .A1(net554),
    .B1(_1022_),
    .X(_1023_));
 sg13g2_xor2_1 _4234_ (.B(_1023_),
    .A(_1021_),
    .X(_1024_));
 sg13g2_a21oi_1 _4235_ (.A1(net526),
    .A2(\load_weights[107] ),
    .Y(_1025_),
    .B1(\load_weights[119] ));
 sg13g2_a21o_1 _4236_ (.A2(\load_weights[119] ),
    .A1(net526),
    .B1(_1025_),
    .X(_1026_));
 sg13g2_inv_1 _4237_ (.Y(_1027_),
    .A(_1026_));
 sg13g2_nand2_1 _4238_ (.Y(_1028_),
    .A(_1024_),
    .B(_1027_));
 sg13g2_nand2b_1 _4239_ (.Y(_1029_),
    .B(_1026_),
    .A_N(_1024_));
 sg13g2_nand2_1 _4240_ (.Y(_1030_),
    .A(_1024_),
    .B(_1026_));
 sg13g2_nand2b_1 _4241_ (.Y(_1031_),
    .B(_1027_),
    .A_N(_1024_));
 sg13g2_nor2_1 _4242_ (.A(_0006_),
    .B(net434),
    .Y(_1032_));
 sg13g2_and2_1 _4243_ (.A(\load_weights[109] ),
    .B(\load_weights[108] ),
    .X(_1033_));
 sg13g2_xor2_1 _4244_ (.B(\load_weights[108] ),
    .A(\load_weights[109] ),
    .X(_1034_));
 sg13g2_xnor2_1 _4245_ (.Y(_1035_),
    .A(\load_weights[110] ),
    .B(_1034_));
 sg13g2_inv_1 _4246_ (.Y(_1036_),
    .A(_1035_));
 sg13g2_nand2_1 _4247_ (.Y(_1037_),
    .A(\load_weights[112] ),
    .B(_1036_));
 sg13g2_xor2_1 _4248_ (.B(_1035_),
    .A(\load_weights[112] ),
    .X(_1038_));
 sg13g2_xor2_1 _4249_ (.B(_1038_),
    .A(_0007_),
    .X(_1039_));
 sg13g2_and2_1 _4250_ (.A(\load_weights[114] ),
    .B(\load_weights[116] ),
    .X(_1040_));
 sg13g2_xor2_1 _4251_ (.B(\load_weights[116] ),
    .A(\load_weights[114] ),
    .X(_1041_));
 sg13g2_xor2_1 _4252_ (.B(_1041_),
    .A(\load_weights[118] ),
    .X(_1042_));
 sg13g2_nand2_1 _4253_ (.Y(_1043_),
    .A(_1039_),
    .B(_1042_));
 sg13g2_xnor2_1 _4254_ (.Y(_1044_),
    .A(_1039_),
    .B(_1042_));
 sg13g2_or2_1 _4255_ (.X(_1045_),
    .B(_1044_),
    .A(_1946_));
 sg13g2_xnor2_1 _4256_ (.Y(_1046_),
    .A(_1946_),
    .B(_1044_));
 sg13g2_xnor2_1 _4257_ (.Y(_1047_),
    .A(_1947_),
    .B(_1046_));
 sg13g2_nor2_1 _4258_ (.A(_1945_),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_xnor2_1 _4259_ (.Y(_1049_),
    .A(\load_weights[113] ),
    .B(_1047_));
 sg13g2_xnor2_1 _4260_ (.Y(_1050_),
    .A(_1948_),
    .B(_1049_));
 sg13g2_xnor2_1 _4261_ (.Y(_1051_),
    .A(\load_weights[111] ),
    .B(_1049_));
 sg13g2_and2_1 _4262_ (.A(_0006_),
    .B(net422),
    .X(_1052_));
 sg13g2_a221oi_1 _4263_ (.B2(net434),
    .C1(_1052_),
    .B1(_1051_),
    .A1(_1030_),
    .Y(_1053_),
    .A2(_1031_));
 sg13g2_a221oi_1 _4264_ (.B2(net434),
    .C1(_1032_),
    .B1(_1050_),
    .A1(_1028_),
    .Y(_1054_),
    .A2(_1029_));
 sg13g2_or3_1 _4265_ (.A(_1019_),
    .B(_1053_),
    .C(_1054_),
    .X(_1055_));
 sg13g2_o21ai_1 _4266_ (.B1(_1019_),
    .Y(_1056_),
    .A1(_1053_),
    .A2(_1054_));
 sg13g2_a21oi_1 _4267_ (.A1(net511),
    .A2(\load_weights[98] ),
    .Y(_1057_),
    .B1(\load_weights[110] ));
 sg13g2_a21oi_1 _4268_ (.A1(net511),
    .A2(\load_weights[110] ),
    .Y(_1058_),
    .B1(_1057_));
 sg13g2_nand3_1 _4269_ (.B(_1056_),
    .C(_1058_),
    .A(_1055_),
    .Y(_1059_));
 sg13g2_a21o_1 _4270_ (.A2(_1056_),
    .A1(_1055_),
    .B1(_1058_),
    .X(_1060_));
 sg13g2_a21oi_1 _4271_ (.A1(net558),
    .A2(\load_weights[100] ),
    .Y(_1061_),
    .B1(\load_weights[112] ));
 sg13g2_a21oi_1 _4272_ (.A1(net558),
    .A2(\load_weights[112] ),
    .Y(_1062_),
    .B1(_1061_));
 sg13g2_nand3_1 _4273_ (.B(_1060_),
    .C(_1062_),
    .A(_1059_),
    .Y(_1063_));
 sg13g2_a21o_1 _4274_ (.A2(_1060_),
    .A1(_1059_),
    .B1(_1062_),
    .X(_1064_));
 sg13g2_a21oi_1 _4275_ (.A1(net539),
    .A2(\load_weights[104] ),
    .Y(_1065_),
    .B1(\load_weights[116] ));
 sg13g2_a21oi_2 _4276_ (.B1(_1065_),
    .Y(_1066_),
    .A2(\load_weights[116] ),
    .A1(net539));
 sg13g2_nand3_1 _4277_ (.B(_1064_),
    .C(_1066_),
    .A(_1063_),
    .Y(_1067_));
 sg13g2_a21oi_1 _4278_ (.A1(_1063_),
    .A2(_1064_),
    .Y(_1068_),
    .B1(_1066_));
 sg13g2_a21o_1 _4279_ (.A2(_1064_),
    .A1(_1063_),
    .B1(_1066_),
    .X(_1069_));
 sg13g2_a21oi_1 _4280_ (.A1(net545),
    .A2(\load_weights[103] ),
    .Y(_1070_),
    .B1(\load_weights[115] ));
 sg13g2_a21o_1 _4281_ (.A2(\load_weights[115] ),
    .A1(net545),
    .B1(_1070_),
    .X(_1071_));
 sg13g2_inv_1 _4282_ (.Y(_1072_),
    .A(_1071_));
 sg13g2_and3_1 _4283_ (.X(_1073_),
    .A(_1067_),
    .B(_1069_),
    .C(_1072_));
 sg13g2_a21oi_1 _4284_ (.A1(_1067_),
    .A2(_1069_),
    .Y(_1074_),
    .B1(_1072_));
 sg13g2_a21oi_1 _4285_ (.A1(net530),
    .A2(\load_weights[106] ),
    .Y(_1075_),
    .B1(\load_weights[118] ));
 sg13g2_a21o_1 _4286_ (.A2(\load_weights[118] ),
    .A1(net530),
    .B1(_1075_),
    .X(_1076_));
 sg13g2_nor3_1 _4287_ (.A(_1073_),
    .B(_1074_),
    .C(_1076_),
    .Y(_1077_));
 sg13g2_o21ai_1 _4288_ (.B1(_1076_),
    .Y(_1078_),
    .A1(_1073_),
    .A2(_1074_));
 sg13g2_nand2b_1 _4289_ (.Y(_1079_),
    .B(_1078_),
    .A_N(_1077_));
 sg13g2_a21oi_1 _4290_ (.A1(net505),
    .A2(net933),
    .Y(_1080_),
    .B1(\load_weights[111] ));
 sg13g2_a21oi_2 _4291_ (.B1(net934),
    .Y(_1081_),
    .A2(net665),
    .A1(net505));
 sg13g2_xnor2_1 _4292_ (.Y(\tt_um_mult_inst.genblk1[4].out_q ),
    .A(_1079_),
    .B(_1081_));
 sg13g2_a21oi_1 _4293_ (.A1(_1078_),
    .A2(_1081_),
    .Y(_1082_),
    .B1(_1077_));
 sg13g2_o21ai_1 _4294_ (.B1(_1067_),
    .Y(_1083_),
    .A1(_1068_),
    .A2(_1071_));
 sg13g2_o21ai_1 _4295_ (.B1(_1018_),
    .Y(_1084_),
    .A1(_1012_),
    .A2(_1014_));
 sg13g2_nand2b_1 _4296_ (.Y(_1085_),
    .B(_1055_),
    .A_N(_1053_));
 sg13g2_o21ai_1 _4297_ (.B1(_1028_),
    .Y(_1086_),
    .A1(_1021_),
    .A2(_1023_));
 sg13g2_nor2_1 _4298_ (.A(\tt_um_mult_inst.genblk1[4].carry[1] ),
    .B(net434),
    .Y(_1087_));
 sg13g2_a21oi_2 _4299_ (.B1(_1048_),
    .Y(_1088_),
    .A2(_1049_),
    .A1(\load_weights[111] ));
 sg13g2_a21oi_1 _4300_ (.A1(\load_weights[118] ),
    .A2(_1041_),
    .Y(_1089_),
    .B1(_1040_));
 sg13g2_and3_1 _4301_ (.X(_1090_),
    .A(\load_weights[110] ),
    .B(\load_weights[112] ),
    .C(_1033_));
 sg13g2_a21oi_1 _4302_ (.A1(\load_weights[110] ),
    .A2(_1034_),
    .Y(_1091_),
    .B1(_1033_));
 sg13g2_a21oi_1 _4303_ (.A1(_1037_),
    .A2(_1091_),
    .Y(_1092_),
    .B1(_1090_));
 sg13g2_o21ai_1 _4304_ (.B1(_1043_),
    .Y(_1093_),
    .A1(_0007_),
    .A2(_1038_));
 sg13g2_xnor2_1 _4305_ (.Y(_1094_),
    .A(_1092_),
    .B(_1093_));
 sg13g2_nor2_1 _4306_ (.A(_1089_),
    .B(_1094_),
    .Y(_1095_));
 sg13g2_xor2_1 _4307_ (.B(_1094_),
    .A(_1089_),
    .X(_1096_));
 sg13g2_o21ai_1 _4308_ (.B1(_1045_),
    .Y(_1097_),
    .A1(_1947_),
    .A2(_1046_));
 sg13g2_xor2_1 _4309_ (.B(_1097_),
    .A(_1096_),
    .X(_1098_));
 sg13g2_nor2b_1 _4310_ (.A(_1088_),
    .B_N(_1098_),
    .Y(_1099_));
 sg13g2_xor2_1 _4311_ (.B(_1098_),
    .A(_1088_),
    .X(_1100_));
 sg13g2_a21oi_1 _4312_ (.A1(net434),
    .A2(_1100_),
    .Y(_1101_),
    .B1(_1087_));
 sg13g2_nand2_1 _4313_ (.Y(_1102_),
    .A(_1086_),
    .B(_1101_));
 sg13g2_xor2_1 _4314_ (.B(_1101_),
    .A(_1086_),
    .X(_1103_));
 sg13g2_xnor2_1 _4315_ (.Y(_1104_),
    .A(_1085_),
    .B(_1103_));
 sg13g2_nor2b_1 _4316_ (.A(_1104_),
    .B_N(_1084_),
    .Y(_1105_));
 sg13g2_xor2_1 _4317_ (.B(_1104_),
    .A(_1084_),
    .X(_1106_));
 sg13g2_nand2_1 _4318_ (.Y(_1107_),
    .A(_1059_),
    .B(_1063_));
 sg13g2_nand2b_1 _4319_ (.Y(_1108_),
    .B(_1107_),
    .A_N(_1106_));
 sg13g2_xnor2_1 _4320_ (.Y(_1109_),
    .A(_1106_),
    .B(_1107_));
 sg13g2_nand2_1 _4321_ (.Y(_1110_),
    .A(_1083_),
    .B(_1109_));
 sg13g2_xnor2_1 _4322_ (.Y(_1111_),
    .A(_1083_),
    .B(_1109_));
 sg13g2_xor2_1 _4323_ (.B(_1111_),
    .A(_1082_),
    .X(\tt_um_mult_inst.genblk1[4].carry_q[0] ));
 sg13g2_a21o_1 _4324_ (.A2(_1103_),
    .A1(_1085_),
    .B1(_1105_),
    .X(_1112_));
 sg13g2_a21o_1 _4325_ (.A2(_1097_),
    .A1(_1096_),
    .B1(_1099_),
    .X(_1113_));
 sg13g2_a21o_1 _4326_ (.A2(_1093_),
    .A1(_1092_),
    .B1(_1095_),
    .X(_1114_));
 sg13g2_nand2_1 _4327_ (.Y(_1115_),
    .A(_1090_),
    .B(_1114_));
 sg13g2_xor2_1 _4328_ (.B(_1114_),
    .A(_1090_),
    .X(_1116_));
 sg13g2_a21oi_1 _4329_ (.A1(_1113_),
    .A2(_1116_),
    .Y(_1117_),
    .B1(net422));
 sg13g2_o21ai_1 _4330_ (.B1(_1117_),
    .Y(_1118_),
    .A1(_1113_),
    .A2(_1116_));
 sg13g2_nand2_1 _4331_ (.Y(_1119_),
    .A(\tt_um_mult_inst.genblk1[4].carry[2] ),
    .B(net422));
 sg13g2_a21oi_2 _4332_ (.B1(_1102_),
    .Y(_1120_),
    .A2(_1119_),
    .A1(_1118_));
 sg13g2_nand3_1 _4333_ (.B(_1118_),
    .C(_1119_),
    .A(_1102_),
    .Y(_1121_));
 sg13g2_nand2b_1 _4334_ (.Y(_1122_),
    .B(_1121_),
    .A_N(_1120_));
 sg13g2_nand2b_1 _4335_ (.Y(_1123_),
    .B(_1112_),
    .A_N(_1122_));
 sg13g2_xor2_1 _4336_ (.B(_1122_),
    .A(_1112_),
    .X(_1124_));
 sg13g2_nor2_1 _4337_ (.A(_1108_),
    .B(_1124_),
    .Y(_1125_));
 sg13g2_xor2_1 _4338_ (.B(_1124_),
    .A(_1108_),
    .X(_1126_));
 sg13g2_o21ai_1 _4339_ (.B1(_1110_),
    .Y(_1127_),
    .A1(_1082_),
    .A2(_1111_));
 sg13g2_xor2_1 _4340_ (.B(_1127_),
    .A(_1126_),
    .X(\tt_um_mult_inst.genblk1[4].carry_q[1] ));
 sg13g2_a22oi_1 _4341_ (.Y(_1128_),
    .B1(_1115_),
    .B2(_1117_),
    .A2(net422),
    .A1(net928));
 sg13g2_xnor2_1 _4342_ (.Y(_1129_),
    .A(_1120_),
    .B(_1128_));
 sg13g2_nor2_1 _4343_ (.A(_1123_),
    .B(_1129_),
    .Y(_1130_));
 sg13g2_nand2_1 _4344_ (.Y(_1131_),
    .A(_1123_),
    .B(_1129_));
 sg13g2_nor2b_1 _4345_ (.A(_1130_),
    .B_N(_1131_),
    .Y(_1132_));
 sg13g2_a21oi_1 _4346_ (.A1(_1126_),
    .A2(_1127_),
    .Y(_1133_),
    .B1(_1125_));
 sg13g2_xnor2_1 _4347_ (.Y(\tt_um_mult_inst.genblk1[4].carry_q[2] ),
    .A(_1132_),
    .B(_1133_));
 sg13g2_nand3_1 _4348_ (.B(_1127_),
    .C(_1131_),
    .A(_1126_),
    .Y(_1134_));
 sg13g2_or3_1 _4349_ (.A(_1108_),
    .B(_1124_),
    .C(_1129_),
    .X(_1135_));
 sg13g2_a21oi_1 _4350_ (.A1(_1120_),
    .A2(_1128_),
    .Y(_1136_),
    .B1(_1130_));
 sg13g2_nand3_1 _4351_ (.B(_1135_),
    .C(_1136_),
    .A(_1134_),
    .Y(\tt_um_mult_inst.genblk1[4].carry_q[3] ));
 sg13g2_a21oi_1 _4352_ (.A1(net550),
    .A2(\load_weights[30] ),
    .Y(_1137_),
    .B1(\load_weights[42] ));
 sg13g2_a21o_1 _4353_ (.A2(\load_weights[42] ),
    .A1(net550),
    .B1(_1137_),
    .X(_1138_));
 sg13g2_a21oi_1 _4354_ (.A1(net560),
    .A2(\load_weights[28] ),
    .Y(_1139_),
    .B1(\load_weights[40] ));
 sg13g2_a21o_1 _4355_ (.A2(\load_weights[40] ),
    .A1(net560),
    .B1(_1139_),
    .X(_1140_));
 sg13g2_xor2_1 _4356_ (.B(_1140_),
    .A(_1138_),
    .X(_1141_));
 sg13g2_a21oi_1 _4357_ (.A1(net513),
    .A2(\load_weights[26] ),
    .Y(_1142_),
    .B1(\load_weights[38] ));
 sg13g2_a21oi_1 _4358_ (.A1(net513),
    .A2(\load_weights[38] ),
    .Y(_1143_),
    .B1(_1142_));
 sg13g2_nand2_1 _4359_ (.Y(_1144_),
    .A(_1141_),
    .B(_1143_));
 sg13g2_xnor2_1 _4360_ (.Y(_1145_),
    .A(_1141_),
    .B(_1143_));
 sg13g2_a21oi_1 _4361_ (.A1(net528),
    .A2(\load_weights[35] ),
    .Y(_1146_),
    .B1(\load_weights[47] ));
 sg13g2_a21o_1 _4362_ (.A2(\load_weights[47] ),
    .A1(net528),
    .B1(_1146_),
    .X(_1147_));
 sg13g2_a21oi_1 _4363_ (.A1(net532),
    .A2(\load_weights[34] ),
    .Y(_1148_),
    .B1(\load_weights[46] ));
 sg13g2_a21o_1 _4364_ (.A2(\load_weights[46] ),
    .A1(net532),
    .B1(_1148_),
    .X(_1149_));
 sg13g2_xor2_1 _4365_ (.B(_1149_),
    .A(_1147_),
    .X(_1150_));
 sg13g2_a21oi_1 _4366_ (.A1(net541),
    .A2(\load_weights[32] ),
    .Y(_1151_),
    .B1(\load_weights[44] ));
 sg13g2_a21o_1 _4367_ (.A2(\load_weights[44] ),
    .A1(net541),
    .B1(_1151_),
    .X(_1152_));
 sg13g2_inv_1 _4368_ (.Y(_1153_),
    .A(_1152_));
 sg13g2_nand2_1 _4369_ (.Y(_1154_),
    .A(_1150_),
    .B(_1153_));
 sg13g2_nand2b_1 _4370_ (.Y(_1155_),
    .B(_1152_),
    .A_N(_1150_));
 sg13g2_nand2_1 _4371_ (.Y(_1156_),
    .A(_1150_),
    .B(_1152_));
 sg13g2_nand2b_1 _4372_ (.Y(_1157_),
    .B(_1153_),
    .A_N(_1150_));
 sg13g2_nor2_1 _4373_ (.A(_0009_),
    .B(net440),
    .Y(_1158_));
 sg13g2_and2_1 _4374_ (.A(\load_weights[36] ),
    .B(\load_weights[37] ),
    .X(_1159_));
 sg13g2_xor2_1 _4375_ (.B(\load_weights[37] ),
    .A(\load_weights[36] ),
    .X(_1160_));
 sg13g2_xnor2_1 _4376_ (.Y(_1161_),
    .A(\load_weights[38] ),
    .B(_1160_));
 sg13g2_inv_1 _4377_ (.Y(_1162_),
    .A(_1161_));
 sg13g2_nand2_1 _4378_ (.Y(_1163_),
    .A(\load_weights[40] ),
    .B(_1162_));
 sg13g2_xor2_1 _4379_ (.B(_1161_),
    .A(\load_weights[40] ),
    .X(_1164_));
 sg13g2_xor2_1 _4380_ (.B(_1164_),
    .A(_0010_),
    .X(_1165_));
 sg13g2_and2_1 _4381_ (.A(\load_weights[44] ),
    .B(\load_weights[42] ),
    .X(_1166_));
 sg13g2_xor2_1 _4382_ (.B(\load_weights[42] ),
    .A(\load_weights[44] ),
    .X(_1167_));
 sg13g2_xnor2_1 _4383_ (.Y(_1168_),
    .A(\load_weights[46] ),
    .B(_1167_));
 sg13g2_inv_1 _4384_ (.Y(_1169_),
    .A(_1168_));
 sg13g2_nand2_1 _4385_ (.Y(_1170_),
    .A(_1165_),
    .B(_1169_));
 sg13g2_xnor2_1 _4386_ (.Y(_1171_),
    .A(_1165_),
    .B(_1169_));
 sg13g2_nor2_1 _4387_ (.A(_1949_),
    .B(_1171_),
    .Y(_1172_));
 sg13g2_xnor2_1 _4388_ (.Y(_1173_),
    .A(_1949_),
    .B(_1171_));
 sg13g2_inv_1 _4389_ (.Y(_1174_),
    .A(_1173_));
 sg13g2_xor2_1 _4390_ (.B(_1173_),
    .A(\load_weights[45] ),
    .X(_1175_));
 sg13g2_xnor2_1 _4391_ (.Y(_1176_),
    .A(\load_weights[41] ),
    .B(_1175_));
 sg13g2_nand2_1 _4392_ (.Y(_1177_),
    .A(\load_weights[39] ),
    .B(_1176_));
 sg13g2_xnor2_1 _4393_ (.Y(_1178_),
    .A(_1951_),
    .B(_1176_));
 sg13g2_xnor2_1 _4394_ (.Y(_1179_),
    .A(\load_weights[39] ),
    .B(_1176_));
 sg13g2_and2_1 _4395_ (.A(_0009_),
    .B(net429),
    .X(_1180_));
 sg13g2_a221oi_1 _4396_ (.B2(net439),
    .C1(_1180_),
    .B1(_1179_),
    .A1(_1156_),
    .Y(_1181_),
    .A2(_1157_));
 sg13g2_a221oi_1 _4397_ (.B2(net439),
    .C1(_1158_),
    .B1(_1178_),
    .A1(_1154_),
    .Y(_1182_),
    .A2(_1155_));
 sg13g2_or3_1 _4398_ (.A(_1145_),
    .B(_1181_),
    .C(_1182_),
    .X(_1183_));
 sg13g2_o21ai_1 _4399_ (.B1(_1145_),
    .Y(_1184_),
    .A1(_1181_),
    .A2(_1182_));
 sg13g2_a21oi_1 _4400_ (.A1(net509),
    .A2(\load_weights[27] ),
    .Y(_1185_),
    .B1(\load_weights[39] ));
 sg13g2_a21oi_1 _4401_ (.A1(net509),
    .A2(\load_weights[39] ),
    .Y(_1186_),
    .B1(_1185_));
 sg13g2_nand3_1 _4402_ (.B(_1184_),
    .C(_1186_),
    .A(_1183_),
    .Y(_1187_));
 sg13g2_a21o_1 _4403_ (.A2(_1184_),
    .A1(_1183_),
    .B1(_1186_),
    .X(_1188_));
 sg13g2_a21oi_1 _4404_ (.A1(net519),
    .A2(\load_weights[25] ),
    .Y(_1189_),
    .B1(\load_weights[37] ));
 sg13g2_a21oi_1 _4405_ (.A1(net519),
    .A2(\load_weights[37] ),
    .Y(_1190_),
    .B1(_1189_));
 sg13g2_nand3_1 _4406_ (.B(_1188_),
    .C(_1190_),
    .A(_1187_),
    .Y(_1191_));
 sg13g2_a21o_1 _4407_ (.A2(_1188_),
    .A1(_1187_),
    .B1(_1190_),
    .X(_1192_));
 sg13g2_a21oi_1 _4408_ (.A1(net555),
    .A2(\load_weights[29] ),
    .Y(_1193_),
    .B1(\load_weights[41] ));
 sg13g2_a21oi_1 _4409_ (.A1(net555),
    .A2(\load_weights[41] ),
    .Y(_1194_),
    .B1(_1193_));
 sg13g2_nand3_1 _4410_ (.B(_1192_),
    .C(_1194_),
    .A(_1191_),
    .Y(_1195_));
 sg13g2_a21oi_1 _4411_ (.A1(_1191_),
    .A2(_1192_),
    .Y(_1196_),
    .B1(_1194_));
 sg13g2_a21o_1 _4412_ (.A2(_1192_),
    .A1(_1191_),
    .B1(_1194_),
    .X(_1197_));
 sg13g2_a21oi_1 _4413_ (.A1(net523),
    .A2(\load_weights[24] ),
    .Y(_1198_),
    .B1(\load_weights[36] ));
 sg13g2_a21o_1 _4414_ (.A2(\load_weights[36] ),
    .A1(net523),
    .B1(_1198_),
    .X(_1199_));
 sg13g2_inv_1 _4415_ (.Y(_1200_),
    .A(_1199_));
 sg13g2_and3_1 _4416_ (.X(_1201_),
    .A(_1195_),
    .B(_1197_),
    .C(_1200_));
 sg13g2_a21oi_1 _4417_ (.A1(_1195_),
    .A2(_1197_),
    .Y(_1202_),
    .B1(_1200_));
 sg13g2_a21oi_1 _4418_ (.A1(net546),
    .A2(\load_weights[31] ),
    .Y(_1203_),
    .B1(\load_weights[43] ));
 sg13g2_a21o_1 _4419_ (.A2(\load_weights[43] ),
    .A1(net546),
    .B1(_1203_),
    .X(_1204_));
 sg13g2_nor3_1 _4420_ (.A(_1201_),
    .B(_1202_),
    .C(_1204_),
    .Y(_1205_));
 sg13g2_o21ai_1 _4421_ (.B1(_1204_),
    .Y(_1206_),
    .A1(_1201_),
    .A2(_1202_));
 sg13g2_nand2b_1 _4422_ (.Y(_1207_),
    .B(_1206_),
    .A_N(_1205_));
 sg13g2_a21oi_1 _4423_ (.A1(net537),
    .A2(net711),
    .Y(_1208_),
    .B1(net929));
 sg13g2_a21oi_1 _4424_ (.A1(net537),
    .A2(net929),
    .Y(_1209_),
    .B1(_1208_));
 sg13g2_xnor2_1 _4425_ (.Y(\tt_um_mult_inst.genblk1[1].out_q ),
    .A(_1207_),
    .B(_1209_));
 sg13g2_a21oi_1 _4426_ (.A1(_1206_),
    .A2(_1209_),
    .Y(_1210_),
    .B1(_1205_));
 sg13g2_o21ai_1 _4427_ (.B1(_1195_),
    .Y(_1211_),
    .A1(_1196_),
    .A2(_1199_));
 sg13g2_o21ai_1 _4428_ (.B1(_1144_),
    .Y(_1212_),
    .A1(_1138_),
    .A2(_1140_));
 sg13g2_nand2b_1 _4429_ (.Y(_1213_),
    .B(_1183_),
    .A_N(_1181_));
 sg13g2_o21ai_1 _4430_ (.B1(_1154_),
    .Y(_1214_),
    .A1(_1147_),
    .A2(_1149_));
 sg13g2_nand2_1 _4431_ (.Y(_1215_),
    .A(\tt_um_mult_inst.genblk1[1].carry[1] ),
    .B(net429));
 sg13g2_o21ai_1 _4432_ (.B1(_1177_),
    .Y(_1216_),
    .A1(_1950_),
    .A2(_1175_));
 sg13g2_a21oi_1 _4433_ (.A1(\load_weights[45] ),
    .A2(_1174_),
    .Y(_1217_),
    .B1(_1172_));
 sg13g2_a21oi_2 _4434_ (.B1(_1166_),
    .Y(_1218_),
    .A2(_1167_),
    .A1(\load_weights[46] ));
 sg13g2_and3_1 _4435_ (.X(_1219_),
    .A(\load_weights[38] ),
    .B(\load_weights[40] ),
    .C(_1159_));
 sg13g2_a21oi_1 _4436_ (.A1(\load_weights[38] ),
    .A2(_1160_),
    .Y(_1220_),
    .B1(_1159_));
 sg13g2_a21oi_1 _4437_ (.A1(_1163_),
    .A2(_1220_),
    .Y(_1221_),
    .B1(_1219_));
 sg13g2_o21ai_1 _4438_ (.B1(_1170_),
    .Y(_1222_),
    .A1(_0010_),
    .A2(_1164_));
 sg13g2_nand2_1 _4439_ (.Y(_1223_),
    .A(_1221_),
    .B(_1222_));
 sg13g2_xnor2_1 _4440_ (.Y(_1224_),
    .A(_1221_),
    .B(_1222_));
 sg13g2_xor2_1 _4441_ (.B(_1224_),
    .A(_1218_),
    .X(_1225_));
 sg13g2_nor2b_1 _4442_ (.A(_1217_),
    .B_N(_1225_),
    .Y(_1226_));
 sg13g2_xnor2_1 _4443_ (.Y(_1227_),
    .A(_1217_),
    .B(_1225_));
 sg13g2_xnor2_1 _4444_ (.Y(_1228_),
    .A(_1216_),
    .B(_1227_));
 sg13g2_o21ai_1 _4445_ (.B1(_1215_),
    .Y(_1229_),
    .A1(net429),
    .A2(_1228_));
 sg13g2_nand2_1 _4446_ (.Y(_1230_),
    .A(_1214_),
    .B(_1229_));
 sg13g2_xor2_1 _4447_ (.B(_1229_),
    .A(_1214_),
    .X(_1231_));
 sg13g2_nand2_1 _4448_ (.Y(_1232_),
    .A(_1213_),
    .B(_1231_));
 sg13g2_xnor2_1 _4449_ (.Y(_1233_),
    .A(_1213_),
    .B(_1231_));
 sg13g2_nand2b_1 _4450_ (.Y(_1234_),
    .B(_1212_),
    .A_N(_1233_));
 sg13g2_xor2_1 _4451_ (.B(_1233_),
    .A(_1212_),
    .X(_1235_));
 sg13g2_nand2_1 _4452_ (.Y(_1236_),
    .A(_1187_),
    .B(_1191_));
 sg13g2_nand2b_1 _4453_ (.Y(_1237_),
    .B(_1236_),
    .A_N(_1235_));
 sg13g2_xor2_1 _4454_ (.B(_1236_),
    .A(_1235_),
    .X(_1238_));
 sg13g2_nand2b_1 _4455_ (.Y(_1239_),
    .B(_1211_),
    .A_N(_1238_));
 sg13g2_xor2_1 _4456_ (.B(_1238_),
    .A(_1211_),
    .X(_1240_));
 sg13g2_xor2_1 _4457_ (.B(_1240_),
    .A(_1210_),
    .X(\tt_um_mult_inst.genblk1[1].carry_q[0] ));
 sg13g2_o21ai_1 _4458_ (.B1(_1223_),
    .Y(_1241_),
    .A1(_1218_),
    .A2(_1224_));
 sg13g2_nand2_1 _4459_ (.Y(_1242_),
    .A(_1219_),
    .B(_1241_));
 sg13g2_xor2_1 _4460_ (.B(_1241_),
    .A(_1219_),
    .X(_1243_));
 sg13g2_a21o_1 _4461_ (.A2(_1227_),
    .A1(_1216_),
    .B1(_1226_),
    .X(_1244_));
 sg13g2_or2_1 _4462_ (.X(_1245_),
    .B(_1244_),
    .A(_1243_));
 sg13g2_a21oi_1 _4463_ (.A1(_1243_),
    .A2(_1244_),
    .Y(_1246_),
    .B1(net429));
 sg13g2_a22oi_1 _4464_ (.Y(_1247_),
    .B1(_1245_),
    .B2(_1246_),
    .A2(net429),
    .A1(\tt_um_mult_inst.genblk1[1].carry[2] ));
 sg13g2_nor2_1 _4465_ (.A(_1230_),
    .B(_1247_),
    .Y(_1248_));
 sg13g2_xnor2_1 _4466_ (.Y(_1249_),
    .A(_1230_),
    .B(_1247_));
 sg13g2_nand3_1 _4467_ (.B(_1234_),
    .C(_1249_),
    .A(_1232_),
    .Y(_1250_));
 sg13g2_a21o_1 _4468_ (.A2(_1234_),
    .A1(_1232_),
    .B1(_1249_),
    .X(_1251_));
 sg13g2_nand2_1 _4469_ (.Y(_1252_),
    .A(_1250_),
    .B(_1251_));
 sg13g2_nor2_1 _4470_ (.A(_1237_),
    .B(_1252_),
    .Y(_1253_));
 sg13g2_xor2_1 _4471_ (.B(_1252_),
    .A(_1237_),
    .X(_1254_));
 sg13g2_o21ai_1 _4472_ (.B1(_1239_),
    .Y(_1255_),
    .A1(_1210_),
    .A2(_1240_));
 sg13g2_xor2_1 _4473_ (.B(_1255_),
    .A(_1254_),
    .X(\tt_um_mult_inst.genblk1[1].carry_q[1] ));
 sg13g2_a21oi_1 _4474_ (.A1(_1254_),
    .A2(_1255_),
    .Y(_1256_),
    .B1(_1253_));
 sg13g2_a22oi_1 _4475_ (.Y(_1257_),
    .B1(_1242_),
    .B2(_1246_),
    .A2(net429),
    .A1(net930));
 sg13g2_nand2_1 _4476_ (.Y(_1258_),
    .A(_1248_),
    .B(_1257_));
 sg13g2_nor2_1 _4477_ (.A(_1248_),
    .B(_1257_),
    .Y(_1259_));
 sg13g2_xnor2_1 _4478_ (.Y(_1260_),
    .A(_1248_),
    .B(_1257_));
 sg13g2_xor2_1 _4479_ (.B(_1260_),
    .A(_1251_),
    .X(_1261_));
 sg13g2_xnor2_1 _4480_ (.Y(\tt_um_mult_inst.genblk1[1].carry_q[2] ),
    .A(_1256_),
    .B(_1261_));
 sg13g2_nand3_1 _4481_ (.B(_1255_),
    .C(_1261_),
    .A(_1254_),
    .Y(_1262_));
 sg13g2_nand2_1 _4482_ (.Y(_1263_),
    .A(_1251_),
    .B(_1258_));
 sg13g2_nor2_1 _4483_ (.A(_1253_),
    .B(_1263_),
    .Y(_1264_));
 sg13g2_o21ai_1 _4484_ (.B1(_1262_),
    .Y(\tt_um_mult_inst.genblk1[1].carry_q[3] ),
    .A1(_1259_),
    .A2(_1264_));
 sg13g2_a21oi_1 _4485_ (.A1(net535),
    .A2(\load_weights[129] ),
    .Y(_1265_),
    .B1(\load_weights[141] ));
 sg13g2_a21o_1 _4486_ (.A2(\load_weights[141] ),
    .A1(net535),
    .B1(_1265_),
    .X(_1266_));
 sg13g2_a21oi_1 _4487_ (.A1(net549),
    .A2(\load_weights[126] ),
    .Y(_1267_),
    .B1(\load_weights[138] ));
 sg13g2_a21o_1 _4488_ (.A2(\load_weights[138] ),
    .A1(net549),
    .B1(_1267_),
    .X(_1268_));
 sg13g2_xor2_1 _4489_ (.B(_1268_),
    .A(_1266_),
    .X(_1269_));
 sg13g2_a21oi_1 _4490_ (.A1(net521),
    .A2(\load_weights[120] ),
    .Y(_1270_),
    .B1(\load_weights[132] ));
 sg13g2_a21oi_2 _4491_ (.B1(_1270_),
    .Y(_1271_),
    .A2(\load_weights[132] ),
    .A1(net521));
 sg13g2_nand2_1 _4492_ (.Y(_1272_),
    .A(_1269_),
    .B(_1271_));
 sg13g2_xnor2_1 _4493_ (.Y(_1273_),
    .A(_1269_),
    .B(_1271_));
 sg13g2_a21oi_1 _4494_ (.A1(net545),
    .A2(\load_weights[127] ),
    .Y(_1274_),
    .B1(\load_weights[139] ));
 sg13g2_a21o_1 _4495_ (.A2(\load_weights[139] ),
    .A1(net545),
    .B1(_1274_),
    .X(_1275_));
 sg13g2_a21oi_1 _4496_ (.A1(net554),
    .A2(\load_weights[125] ),
    .Y(_1276_),
    .B1(\load_weights[137] ));
 sg13g2_a21o_1 _4497_ (.A2(\load_weights[137] ),
    .A1(net554),
    .B1(_1276_),
    .X(_1277_));
 sg13g2_xor2_1 _4498_ (.B(_1277_),
    .A(_1275_),
    .X(_1278_));
 sg13g2_a21oi_1 _4499_ (.A1(net526),
    .A2(\load_weights[131] ),
    .Y(_1279_),
    .B1(\load_weights[143] ));
 sg13g2_a21o_1 _4500_ (.A2(\load_weights[143] ),
    .A1(net526),
    .B1(_1279_),
    .X(_1280_));
 sg13g2_inv_1 _4501_ (.Y(_1281_),
    .A(_1280_));
 sg13g2_nand2_1 _4502_ (.Y(_1282_),
    .A(_1278_),
    .B(_1281_));
 sg13g2_nand2b_1 _4503_ (.Y(_1283_),
    .B(_1280_),
    .A_N(_1278_));
 sg13g2_nand2_1 _4504_ (.Y(_1284_),
    .A(_1278_),
    .B(_1280_));
 sg13g2_nand2b_1 _4505_ (.Y(_1285_),
    .B(_1281_),
    .A_N(_1278_));
 sg13g2_nor2_1 _4506_ (.A(_0012_),
    .B(net436),
    .Y(_1286_));
 sg13g2_and2_1 _4507_ (.A(\load_weights[132] ),
    .B(\load_weights[133] ),
    .X(_1287_));
 sg13g2_xor2_1 _4508_ (.B(\load_weights[133] ),
    .A(\load_weights[132] ),
    .X(_1288_));
 sg13g2_xnor2_1 _4509_ (.Y(_1289_),
    .A(\load_weights[134] ),
    .B(_1288_));
 sg13g2_inv_1 _4510_ (.Y(_1290_),
    .A(_1289_));
 sg13g2_nand2_1 _4511_ (.Y(_1291_),
    .A(\load_weights[136] ),
    .B(_1290_));
 sg13g2_xor2_1 _4512_ (.B(_1289_),
    .A(\load_weights[136] ),
    .X(_1292_));
 sg13g2_xor2_1 _4513_ (.B(_1292_),
    .A(_0013_),
    .X(_1293_));
 sg13g2_and2_1 _4514_ (.A(\load_weights[138] ),
    .B(\load_weights[140] ),
    .X(_1294_));
 sg13g2_xor2_1 _4515_ (.B(\load_weights[140] ),
    .A(\load_weights[138] ),
    .X(_1295_));
 sg13g2_xor2_1 _4516_ (.B(_1295_),
    .A(\load_weights[142] ),
    .X(_1296_));
 sg13g2_nand2_1 _4517_ (.Y(_1297_),
    .A(_1293_),
    .B(_1296_));
 sg13g2_xnor2_1 _4518_ (.Y(_1298_),
    .A(_1293_),
    .B(_1296_));
 sg13g2_or2_1 _4519_ (.X(_1299_),
    .B(_1298_),
    .A(_1952_));
 sg13g2_xnor2_1 _4520_ (.Y(_1300_),
    .A(_1952_),
    .B(_1298_));
 sg13g2_xnor2_1 _4521_ (.Y(_1301_),
    .A(_1954_),
    .B(_1300_));
 sg13g2_nor2_1 _4522_ (.A(_1953_),
    .B(_1301_),
    .Y(_1302_));
 sg13g2_xnor2_1 _4523_ (.Y(_1303_),
    .A(\load_weights[137] ),
    .B(_1301_));
 sg13g2_xnor2_1 _4524_ (.Y(_1304_),
    .A(_1955_),
    .B(_1303_));
 sg13g2_xnor2_1 _4525_ (.Y(_1305_),
    .A(\load_weights[135] ),
    .B(_1303_));
 sg13g2_and2_1 _4526_ (.A(_0012_),
    .B(net422),
    .X(_1306_));
 sg13g2_a221oi_1 _4527_ (.B2(net436),
    .C1(_1306_),
    .B1(_1305_),
    .A1(_1284_),
    .Y(_1307_),
    .A2(_1285_));
 sg13g2_a221oi_1 _4528_ (.B2(net434),
    .C1(_1286_),
    .B1(_1304_),
    .A1(_1282_),
    .Y(_1308_),
    .A2(_1283_));
 sg13g2_or3_1 _4529_ (.A(_1273_),
    .B(_1307_),
    .C(_1308_),
    .X(_1309_));
 sg13g2_o21ai_1 _4530_ (.B1(_1273_),
    .Y(_1310_),
    .A1(_1307_),
    .A2(_1308_));
 sg13g2_a21oi_1 _4531_ (.A1(net558),
    .A2(\load_weights[124] ),
    .Y(_1311_),
    .B1(\load_weights[136] ));
 sg13g2_a21oi_1 _4532_ (.A1(net558),
    .A2(\load_weights[136] ),
    .Y(_1312_),
    .B1(_1311_));
 sg13g2_nand3_1 _4533_ (.B(_1310_),
    .C(_1312_),
    .A(_1309_),
    .Y(_1313_));
 sg13g2_a21o_1 _4534_ (.A2(_1310_),
    .A1(_1309_),
    .B1(_1312_),
    .X(_1314_));
 sg13g2_a21oi_1 _4535_ (.A1(net516),
    .A2(\load_weights[121] ),
    .Y(_1315_),
    .B1(\load_weights[133] ));
 sg13g2_a21oi_1 _4536_ (.A1(net516),
    .A2(\load_weights[133] ),
    .Y(_1316_),
    .B1(_1315_));
 sg13g2_nand3_1 _4537_ (.B(_1314_),
    .C(_1316_),
    .A(_1313_),
    .Y(_1317_));
 sg13g2_a21o_1 _4538_ (.A2(_1314_),
    .A1(_1313_),
    .B1(_1316_),
    .X(_1318_));
 sg13g2_a21oi_1 _4539_ (.A1(net539),
    .A2(\load_weights[128] ),
    .Y(_1319_),
    .B1(\load_weights[140] ));
 sg13g2_a21oi_2 _4540_ (.B1(_1319_),
    .Y(_1320_),
    .A2(\load_weights[140] ),
    .A1(net539));
 sg13g2_nand3_1 _4541_ (.B(_1318_),
    .C(_1320_),
    .A(_1317_),
    .Y(_1321_));
 sg13g2_a21oi_1 _4542_ (.A1(_1317_),
    .A2(_1318_),
    .Y(_1322_),
    .B1(_1320_));
 sg13g2_a21o_1 _4543_ (.A2(_1318_),
    .A1(_1317_),
    .B1(_1320_),
    .X(_1323_));
 sg13g2_a21oi_1 _4544_ (.A1(net511),
    .A2(\load_weights[122] ),
    .Y(_1324_),
    .B1(\load_weights[134] ));
 sg13g2_a21o_1 _4545_ (.A2(\load_weights[134] ),
    .A1(net511),
    .B1(_1324_),
    .X(_1325_));
 sg13g2_inv_1 _4546_ (.Y(_1326_),
    .A(_1325_));
 sg13g2_and3_1 _4547_ (.X(_1327_),
    .A(_1321_),
    .B(_1323_),
    .C(_1326_));
 sg13g2_a21oi_1 _4548_ (.A1(_1321_),
    .A2(_1323_),
    .Y(_1328_),
    .B1(_1326_));
 sg13g2_a21oi_1 _4549_ (.A1(net530),
    .A2(\load_weights[130] ),
    .Y(_1329_),
    .B1(\load_weights[142] ));
 sg13g2_a21o_1 _4550_ (.A2(\load_weights[142] ),
    .A1(net530),
    .B1(_1329_),
    .X(_1330_));
 sg13g2_nor3_1 _4551_ (.A(_1327_),
    .B(_1328_),
    .C(_1330_),
    .Y(_1331_));
 sg13g2_o21ai_1 _4552_ (.B1(_1330_),
    .Y(_1332_),
    .A1(_1327_),
    .A2(_1328_));
 sg13g2_nand2b_1 _4553_ (.Y(_1333_),
    .B(_1332_),
    .A_N(_1331_));
 sg13g2_a21oi_1 _4554_ (.A1(net505),
    .A2(net936),
    .Y(_1334_),
    .B1(\load_weights[135] ));
 sg13g2_a21oi_1 _4555_ (.A1(net505),
    .A2(\load_weights[135] ),
    .Y(_1335_),
    .B1(_1334_));
 sg13g2_xnor2_1 _4556_ (.Y(\tt_um_mult_inst.genblk1[5].out_q ),
    .A(_1333_),
    .B(_1335_));
 sg13g2_a21oi_1 _4557_ (.A1(_1332_),
    .A2(_1335_),
    .Y(_1336_),
    .B1(_1331_));
 sg13g2_o21ai_1 _4558_ (.B1(_1321_),
    .Y(_1337_),
    .A1(_1322_),
    .A2(_1325_));
 sg13g2_o21ai_1 _4559_ (.B1(_1272_),
    .Y(_1338_),
    .A1(_1266_),
    .A2(_1268_));
 sg13g2_nand2b_1 _4560_ (.Y(_1339_),
    .B(_1309_),
    .A_N(_1307_));
 sg13g2_o21ai_1 _4561_ (.B1(_1282_),
    .Y(_1340_),
    .A1(_1275_),
    .A2(_1277_));
 sg13g2_a21oi_1 _4562_ (.A1(\load_weights[135] ),
    .A2(_1303_),
    .Y(_1341_),
    .B1(_1302_));
 sg13g2_a21oi_2 _4563_ (.B1(_1294_),
    .Y(_1342_),
    .A2(_1295_),
    .A1(\load_weights[142] ));
 sg13g2_and3_1 _4564_ (.X(_1343_),
    .A(\load_weights[134] ),
    .B(\load_weights[136] ),
    .C(_1287_));
 sg13g2_a21oi_1 _4565_ (.A1(\load_weights[134] ),
    .A2(_1288_),
    .Y(_1344_),
    .B1(_1287_));
 sg13g2_a21oi_1 _4566_ (.A1(_1291_),
    .A2(_1344_),
    .Y(_1345_),
    .B1(_1343_));
 sg13g2_o21ai_1 _4567_ (.B1(_1297_),
    .Y(_1346_),
    .A1(_0013_),
    .A2(_1292_));
 sg13g2_xnor2_1 _4568_ (.Y(_1347_),
    .A(_1345_),
    .B(_1346_));
 sg13g2_nor2_1 _4569_ (.A(_1342_),
    .B(_1347_),
    .Y(_1348_));
 sg13g2_xor2_1 _4570_ (.B(_1347_),
    .A(_1342_),
    .X(_1349_));
 sg13g2_o21ai_1 _4571_ (.B1(_1299_),
    .Y(_1350_),
    .A1(_1954_),
    .A2(_1300_));
 sg13g2_xor2_1 _4572_ (.B(_1350_),
    .A(_1349_),
    .X(_1351_));
 sg13g2_nor2b_1 _4573_ (.A(_1341_),
    .B_N(_1351_),
    .Y(_1352_));
 sg13g2_xor2_1 _4574_ (.B(_1351_),
    .A(_1341_),
    .X(_1353_));
 sg13g2_nor2_1 _4575_ (.A(\tt_um_mult_inst.genblk1[5].carry[1] ),
    .B(net434),
    .Y(_1354_));
 sg13g2_a21oi_1 _4576_ (.A1(net434),
    .A2(_1353_),
    .Y(_1355_),
    .B1(_1354_));
 sg13g2_nand2_1 _4577_ (.Y(_1356_),
    .A(_1340_),
    .B(_1355_));
 sg13g2_xor2_1 _4578_ (.B(_1355_),
    .A(_1340_),
    .X(_1357_));
 sg13g2_xnor2_1 _4579_ (.Y(_1358_),
    .A(_1339_),
    .B(_1357_));
 sg13g2_nor2b_1 _4580_ (.A(_1358_),
    .B_N(_1338_),
    .Y(_1359_));
 sg13g2_xor2_1 _4581_ (.B(_1358_),
    .A(_1338_),
    .X(_1360_));
 sg13g2_nand2_1 _4582_ (.Y(_1361_),
    .A(_1313_),
    .B(_1317_));
 sg13g2_nand2b_1 _4583_ (.Y(_1362_),
    .B(_1361_),
    .A_N(_1360_));
 sg13g2_xnor2_1 _4584_ (.Y(_1363_),
    .A(_1360_),
    .B(_1361_));
 sg13g2_nand2_1 _4585_ (.Y(_1364_),
    .A(_1337_),
    .B(_1363_));
 sg13g2_xnor2_1 _4586_ (.Y(_1365_),
    .A(_1337_),
    .B(_1363_));
 sg13g2_xor2_1 _4587_ (.B(_1365_),
    .A(_1336_),
    .X(\tt_um_mult_inst.genblk1[5].carry_q[0] ));
 sg13g2_a21o_1 _4588_ (.A2(_1357_),
    .A1(_1339_),
    .B1(_1359_),
    .X(_1366_));
 sg13g2_a21o_1 _4589_ (.A2(_1350_),
    .A1(_1349_),
    .B1(_1352_),
    .X(_1367_));
 sg13g2_a21o_1 _4590_ (.A2(_1346_),
    .A1(_1345_),
    .B1(_1348_),
    .X(_1368_));
 sg13g2_nand2_1 _4591_ (.Y(_1369_),
    .A(_1343_),
    .B(_1368_));
 sg13g2_xor2_1 _4592_ (.B(_1368_),
    .A(_1343_),
    .X(_1370_));
 sg13g2_a21oi_1 _4593_ (.A1(_1367_),
    .A2(_1370_),
    .Y(_1371_),
    .B1(net422));
 sg13g2_o21ai_1 _4594_ (.B1(_1371_),
    .Y(_1372_),
    .A1(_1367_),
    .A2(_1370_));
 sg13g2_nand2_1 _4595_ (.Y(_1373_),
    .A(\tt_um_mult_inst.genblk1[5].carry[2] ),
    .B(net422));
 sg13g2_a21oi_1 _4596_ (.A1(_1372_),
    .A2(_1373_),
    .Y(_1374_),
    .B1(_1356_));
 sg13g2_nand3_1 _4597_ (.B(_1372_),
    .C(_1373_),
    .A(_1356_),
    .Y(_1375_));
 sg13g2_nand2b_1 _4598_ (.Y(_1376_),
    .B(_1375_),
    .A_N(_1374_));
 sg13g2_nand2b_1 _4599_ (.Y(_1377_),
    .B(_1366_),
    .A_N(_1376_));
 sg13g2_xor2_1 _4600_ (.B(_1376_),
    .A(_1366_),
    .X(_1378_));
 sg13g2_nor2_1 _4601_ (.A(_1362_),
    .B(_1378_),
    .Y(_1379_));
 sg13g2_xor2_1 _4602_ (.B(_1378_),
    .A(_1362_),
    .X(_1380_));
 sg13g2_o21ai_1 _4603_ (.B1(_1364_),
    .Y(_1381_),
    .A1(_1336_),
    .A2(_1365_));
 sg13g2_xor2_1 _4604_ (.B(_1381_),
    .A(_1380_),
    .X(\tt_um_mult_inst.genblk1[5].carry_q[1] ));
 sg13g2_a22oi_1 _4605_ (.Y(_1382_),
    .B1(_1369_),
    .B2(_1371_),
    .A2(net422),
    .A1(net926));
 sg13g2_xnor2_1 _4606_ (.Y(_1383_),
    .A(_1374_),
    .B(_1382_));
 sg13g2_nor2_1 _4607_ (.A(_1377_),
    .B(_1383_),
    .Y(_1384_));
 sg13g2_and2_1 _4608_ (.A(_1377_),
    .B(_1383_),
    .X(_1385_));
 sg13g2_nor2_1 _4609_ (.A(_1384_),
    .B(_1385_),
    .Y(_1386_));
 sg13g2_a21oi_1 _4610_ (.A1(_1380_),
    .A2(_1381_),
    .Y(_1387_),
    .B1(_1379_));
 sg13g2_xnor2_1 _4611_ (.Y(\tt_um_mult_inst.genblk1[5].carry_q[2] ),
    .A(_1386_),
    .B(_1387_));
 sg13g2_nor3_1 _4612_ (.A(_1362_),
    .B(_1378_),
    .C(_1383_),
    .Y(_1388_));
 sg13g2_a21oi_1 _4613_ (.A1(_1374_),
    .A2(_1382_),
    .Y(_1389_),
    .B1(_1388_));
 sg13g2_a21oi_1 _4614_ (.A1(_1380_),
    .A2(_1381_),
    .Y(_1390_),
    .B1(_1384_));
 sg13g2_o21ai_1 _4615_ (.B1(_1389_),
    .Y(\tt_um_mult_inst.genblk1[5].carry_q[3] ),
    .A1(_1385_),
    .A2(_1390_));
 sg13g2_a21oi_1 _4616_ (.A1(net513),
    .A2(\load_weights[2] ),
    .Y(_1391_),
    .B1(\load_weights[14] ));
 sg13g2_a21o_1 _4617_ (.A2(\load_weights[14] ),
    .A1(net513),
    .B1(_1391_),
    .X(_1392_));
 sg13g2_a21oi_1 _4618_ (.A1(net528),
    .A2(\load_weights[11] ),
    .Y(_1393_),
    .B1(\load_weights[23] ));
 sg13g2_a21o_1 _4619_ (.A2(\load_weights[23] ),
    .A1(net528),
    .B1(_1393_),
    .X(_1394_));
 sg13g2_xor2_1 _4620_ (.B(_1394_),
    .A(_1392_),
    .X(_1395_));
 sg13g2_a21oi_1 _4621_ (.A1(net537),
    .A2(\load_weights[9] ),
    .Y(_1396_),
    .B1(\load_weights[21] ));
 sg13g2_a21oi_1 _4622_ (.A1(net537),
    .A2(\load_weights[21] ),
    .Y(_1397_),
    .B1(_1396_));
 sg13g2_nand2_1 _4623_ (.Y(_1398_),
    .A(_1395_),
    .B(_1397_));
 sg13g2_xnor2_1 _4624_ (.Y(_1399_),
    .A(_1395_),
    .B(_1397_));
 sg13g2_inv_1 _4625_ (.Y(_1400_),
    .A(_1399_));
 sg13g2_a21oi_1 _4626_ (.A1(net509),
    .A2(\load_weights[3] ),
    .Y(_1401_),
    .B1(\load_weights[15] ));
 sg13g2_a21o_1 _4627_ (.A2(\load_weights[15] ),
    .A1(net509),
    .B1(_1401_),
    .X(_1402_));
 sg13g2_a21oi_1 _4628_ (.A1(net519),
    .A2(\load_weights[1] ),
    .Y(_1403_),
    .B1(\load_weights[13] ));
 sg13g2_a21o_1 _4629_ (.A2(\load_weights[13] ),
    .A1(net519),
    .B1(_1403_),
    .X(_1404_));
 sg13g2_xor2_1 _4630_ (.B(_1404_),
    .A(_1402_),
    .X(_1405_));
 sg13g2_a21oi_1 _4631_ (.A1(net560),
    .A2(\load_weights[4] ),
    .Y(_1406_),
    .B1(\load_weights[16] ));
 sg13g2_a21o_1 _4632_ (.A2(\load_weights[16] ),
    .A1(net560),
    .B1(_1406_),
    .X(_1407_));
 sg13g2_inv_1 _4633_ (.Y(_1408_),
    .A(_1407_));
 sg13g2_nand2_1 _4634_ (.Y(_1409_),
    .A(_1405_),
    .B(_1408_));
 sg13g2_nand2b_1 _4635_ (.Y(_1410_),
    .B(_1407_),
    .A_N(_1405_));
 sg13g2_nand2_1 _4636_ (.Y(_1411_),
    .A(_1405_),
    .B(_1407_));
 sg13g2_nand2b_1 _4637_ (.Y(_1412_),
    .B(_1408_),
    .A_N(_1405_));
 sg13g2_nand2_1 _4638_ (.Y(_1413_),
    .A(_1409_),
    .B(_1410_));
 sg13g2_inv_1 _4639_ (.Y(_1414_),
    .A(_1413_));
 sg13g2_nand2_1 _4640_ (.Y(_1415_),
    .A(\load_weights[13] ),
    .B(\load_weights[12] ));
 sg13g2_xnor2_1 _4641_ (.Y(_1416_),
    .A(\load_weights[13] ),
    .B(\load_weights[12] ));
 sg13g2_and2_1 _4642_ (.A(\load_weights[15] ),
    .B(\load_weights[14] ),
    .X(_1417_));
 sg13g2_xor2_1 _4643_ (.B(\load_weights[14] ),
    .A(\load_weights[15] ),
    .X(_1418_));
 sg13g2_xnor2_1 _4644_ (.Y(_1419_),
    .A(\load_weights[17] ),
    .B(_1418_));
 sg13g2_nor2_1 _4645_ (.A(_1416_),
    .B(_1419_),
    .Y(_1420_));
 sg13g2_xnor2_1 _4646_ (.Y(_1421_),
    .A(_1416_),
    .B(_1419_));
 sg13g2_and2_1 _4647_ (.A(\load_weights[19] ),
    .B(\load_weights[21] ),
    .X(_1422_));
 sg13g2_xor2_1 _4648_ (.B(\load_weights[21] ),
    .A(\load_weights[19] ),
    .X(_1423_));
 sg13g2_xnor2_1 _4649_ (.Y(_1424_),
    .A(\load_weights[23] ),
    .B(_1423_));
 sg13g2_nor2_1 _4650_ (.A(_1421_),
    .B(_1424_),
    .Y(_1425_));
 sg13g2_xor2_1 _4651_ (.B(_1424_),
    .A(_1421_),
    .X(_1426_));
 sg13g2_nand2_1 _4652_ (.Y(_1427_),
    .A(\load_weights[20] ),
    .B(_1426_));
 sg13g2_xnor2_1 _4653_ (.Y(_1428_),
    .A(\load_weights[20] ),
    .B(_1426_));
 sg13g2_xnor2_1 _4654_ (.Y(_1429_),
    .A(\load_weights[22] ),
    .B(_1428_));
 sg13g2_nand2_1 _4655_ (.Y(_1430_),
    .A(\load_weights[18] ),
    .B(_1429_));
 sg13g2_xor2_1 _4656_ (.B(_1429_),
    .A(\load_weights[18] ),
    .X(_1431_));
 sg13g2_xnor2_1 _4657_ (.Y(_1432_),
    .A(\load_weights[18] ),
    .B(_1429_));
 sg13g2_nand2_1 _4658_ (.Y(_1433_),
    .A(\load_weights[16] ),
    .B(_1431_));
 sg13g2_a21oi_1 _4659_ (.A1(_1956_),
    .A2(_1432_),
    .Y(_1434_),
    .B1(net430));
 sg13g2_xnor2_1 _4660_ (.Y(_1435_),
    .A(\load_weights[16] ),
    .B(_1431_));
 sg13g2_nor2_1 _4661_ (.A(_1958_),
    .B(net440),
    .Y(_1436_));
 sg13g2_a221oi_1 _4662_ (.B2(net440),
    .C1(_1436_),
    .B1(_1435_),
    .A1(_1411_),
    .Y(_1437_),
    .A2(_1412_));
 sg13g2_a221oi_1 _4663_ (.B2(_1434_),
    .C1(_1414_),
    .B1(_1433_),
    .A1(_1958_),
    .Y(_1438_),
    .A2(net430));
 sg13g2_a221oi_1 _4664_ (.B2(_1434_),
    .C1(_1413_),
    .B1(_1433_),
    .A1(_1958_),
    .Y(_1439_),
    .A2(net430));
 sg13g2_a221oi_1 _4665_ (.B2(net440),
    .C1(_1436_),
    .B1(_1435_),
    .A1(_1409_),
    .Y(_1440_),
    .A2(_1410_));
 sg13g2_nor3_1 _4666_ (.A(_1399_),
    .B(_1437_),
    .C(_1438_),
    .Y(_1441_));
 sg13g2_o21ai_1 _4667_ (.B1(_1400_),
    .Y(_1442_),
    .A1(_1439_),
    .A2(_1440_));
 sg13g2_nor3_1 _4668_ (.A(_1400_),
    .B(_1439_),
    .C(_1440_),
    .Y(_1443_));
 sg13g2_o21ai_1 _4669_ (.B1(_1399_),
    .Y(_1444_),
    .A1(_1437_),
    .A2(_1438_));
 sg13g2_a21oi_1 _4670_ (.A1(net532),
    .A2(\load_weights[10] ),
    .Y(_1445_),
    .B1(\load_weights[22] ));
 sg13g2_a21oi_1 _4671_ (.A1(net532),
    .A2(\load_weights[22] ),
    .Y(_1446_),
    .B1(_1445_));
 sg13g2_a21o_1 _4672_ (.A2(\load_weights[22] ),
    .A1(net532),
    .B1(_1445_),
    .X(_1447_));
 sg13g2_nor3_1 _4673_ (.A(_1441_),
    .B(_1443_),
    .C(_1447_),
    .Y(_1448_));
 sg13g2_nand3_1 _4674_ (.B(_1444_),
    .C(_1446_),
    .A(_1442_),
    .Y(_1449_));
 sg13g2_a21oi_1 _4675_ (.A1(_1442_),
    .A2(_1444_),
    .Y(_1450_),
    .B1(_1446_));
 sg13g2_o21ai_1 _4676_ (.B1(_1447_),
    .Y(_1451_),
    .A1(_1441_),
    .A2(_1443_));
 sg13g2_a21oi_1 _4677_ (.A1(net541),
    .A2(\load_weights[8] ),
    .Y(_1452_),
    .B1(\load_weights[20] ));
 sg13g2_a21oi_2 _4678_ (.B1(_1452_),
    .Y(_1453_),
    .A2(\load_weights[20] ),
    .A1(net543));
 sg13g2_a21o_1 _4679_ (.A2(\load_weights[20] ),
    .A1(net542),
    .B1(_1452_),
    .X(_1454_));
 sg13g2_nor3_1 _4680_ (.A(_1448_),
    .B(_1450_),
    .C(_1454_),
    .Y(_1455_));
 sg13g2_nand3_1 _4681_ (.B(_1451_),
    .C(_1453_),
    .A(_1449_),
    .Y(_1456_));
 sg13g2_a21oi_1 _4682_ (.A1(_1449_),
    .A2(_1451_),
    .Y(_1457_),
    .B1(_1453_));
 sg13g2_o21ai_1 _4683_ (.B1(_1454_),
    .Y(_1458_),
    .A1(_1448_),
    .A2(_1450_));
 sg13g2_a21oi_1 _4684_ (.A1(net523),
    .A2(\load_weights[0] ),
    .Y(_1459_),
    .B1(\load_weights[12] ));
 sg13g2_a21oi_1 _4685_ (.A1(net523),
    .A2(\load_weights[12] ),
    .Y(_1460_),
    .B1(_1459_));
 sg13g2_a21o_1 _4686_ (.A2(\load_weights[12] ),
    .A1(net523),
    .B1(_1459_),
    .X(_1461_));
 sg13g2_nor3_1 _4687_ (.A(_1455_),
    .B(_1457_),
    .C(_1461_),
    .Y(_1462_));
 sg13g2_nand3_1 _4688_ (.B(_1458_),
    .C(_1460_),
    .A(_1456_),
    .Y(_1463_));
 sg13g2_a21oi_1 _4689_ (.A1(_1456_),
    .A2(_1458_),
    .Y(_1464_),
    .B1(_1460_));
 sg13g2_o21ai_1 _4690_ (.B1(_1461_),
    .Y(_1465_),
    .A1(_1455_),
    .A2(_1457_));
 sg13g2_a21oi_1 _4691_ (.A1(net546),
    .A2(\load_weights[7] ),
    .Y(_1466_),
    .B1(\load_weights[19] ));
 sg13g2_a21o_2 _4692_ (.A2(\load_weights[19] ),
    .A1(net546),
    .B1(_1466_),
    .X(_1467_));
 sg13g2_inv_1 _4693_ (.Y(_1468_),
    .A(_1467_));
 sg13g2_nor3_1 _4694_ (.A(_1462_),
    .B(_1464_),
    .C(_1467_),
    .Y(_1469_));
 sg13g2_a21oi_1 _4695_ (.A1(_1463_),
    .A2(_1465_),
    .Y(_1470_),
    .B1(_1468_));
 sg13g2_nand3_1 _4696_ (.B(_1465_),
    .C(_1467_),
    .A(_1463_),
    .Y(_1471_));
 sg13g2_o21ai_1 _4697_ (.B1(_1468_),
    .Y(_1472_),
    .A1(_1462_),
    .A2(_1464_));
 sg13g2_a21oi_1 _4698_ (.A1(net555),
    .A2(\load_weights[5] ),
    .Y(_1473_),
    .B1(\load_weights[17] ));
 sg13g2_a21o_1 _4699_ (.A2(\load_weights[17] ),
    .A1(net555),
    .B1(_1473_),
    .X(_1474_));
 sg13g2_nor3_1 _4700_ (.A(_1469_),
    .B(_1470_),
    .C(_1474_),
    .Y(_1475_));
 sg13g2_and3_1 _4701_ (.X(_1476_),
    .A(_1471_),
    .B(_1472_),
    .C(_1474_));
 sg13g2_o21ai_1 _4702_ (.B1(_1474_),
    .Y(_1477_),
    .A1(_1469_),
    .A2(_1470_));
 sg13g2_a21oi_1 _4703_ (.A1(net550),
    .A2(\load_weights[6] ),
    .Y(_1478_),
    .B1(\load_weights[18] ));
 sg13g2_a21oi_2 _4704_ (.B1(_1478_),
    .Y(_1479_),
    .A2(\load_weights[18] ),
    .A1(net550));
 sg13g2_nor3_1 _4705_ (.A(_1475_),
    .B(_1476_),
    .C(_1479_),
    .Y(_1480_));
 sg13g2_o21ai_1 _4706_ (.B1(_1479_),
    .Y(_1481_),
    .A1(_1475_),
    .A2(_1476_));
 sg13g2_nand2b_1 _4707_ (.Y(\tt_um_mult_inst.genblk1[0].out_q ),
    .B(_1481_),
    .A_N(_1480_));
 sg13g2_a21oi_1 _4708_ (.A1(_1477_),
    .A2(_1479_),
    .Y(_1482_),
    .B1(_1475_));
 sg13g2_o21ai_1 _4709_ (.B1(_1398_),
    .Y(_1483_),
    .A1(_1392_),
    .A2(_1394_));
 sg13g2_nand2b_1 _4710_ (.Y(_1484_),
    .B(_1442_),
    .A_N(_1437_));
 sg13g2_o21ai_1 _4711_ (.B1(_1409_),
    .Y(_1485_),
    .A1(_1402_),
    .A2(_1404_));
 sg13g2_nand2_1 _4712_ (.Y(_1486_),
    .A(\tt_um_mult_inst.genblk1[0].carry[1] ),
    .B(net430));
 sg13g2_nand2_2 _4713_ (.Y(_1487_),
    .A(_1430_),
    .B(_1433_));
 sg13g2_a21oi_1 _4714_ (.A1(\load_weights[23] ),
    .A2(_1423_),
    .Y(_1488_),
    .B1(_1422_));
 sg13g2_a21oi_1 _4715_ (.A1(\load_weights[17] ),
    .A2(_1418_),
    .Y(_1489_),
    .B1(_1417_));
 sg13g2_nor2_1 _4716_ (.A(_1415_),
    .B(_1489_),
    .Y(_1490_));
 sg13g2_xnor2_1 _4717_ (.Y(_1491_),
    .A(_1415_),
    .B(_1489_));
 sg13g2_nor2_1 _4718_ (.A(_1420_),
    .B(_1425_),
    .Y(_1492_));
 sg13g2_nor2_1 _4719_ (.A(_1491_),
    .B(_1492_),
    .Y(_1493_));
 sg13g2_xnor2_1 _4720_ (.Y(_1494_),
    .A(_1491_),
    .B(_1492_));
 sg13g2_nor2_1 _4721_ (.A(_1488_),
    .B(_1494_),
    .Y(_1495_));
 sg13g2_xor2_1 _4722_ (.B(_1494_),
    .A(_1488_),
    .X(_1496_));
 sg13g2_o21ai_1 _4723_ (.B1(_1427_),
    .Y(_1497_),
    .A1(_1957_),
    .A2(_1428_));
 sg13g2_and2_1 _4724_ (.A(_1496_),
    .B(_1497_),
    .X(_1498_));
 sg13g2_xor2_1 _4725_ (.B(_1497_),
    .A(_1496_),
    .X(_1499_));
 sg13g2_xnor2_1 _4726_ (.Y(_1500_),
    .A(_1487_),
    .B(_1499_));
 sg13g2_o21ai_1 _4727_ (.B1(_1486_),
    .Y(_1501_),
    .A1(net430),
    .A2(_1500_));
 sg13g2_nand2_1 _4728_ (.Y(_1502_),
    .A(_1485_),
    .B(_1501_));
 sg13g2_xor2_1 _4729_ (.B(_1501_),
    .A(_1485_),
    .X(_1503_));
 sg13g2_nand2_1 _4730_ (.Y(_1504_),
    .A(_1484_),
    .B(_1503_));
 sg13g2_xnor2_1 _4731_ (.Y(_1505_),
    .A(_1484_),
    .B(_1503_));
 sg13g2_nand2b_1 _4732_ (.Y(_1506_),
    .B(_1483_),
    .A_N(_1505_));
 sg13g2_xor2_1 _4733_ (.B(_1505_),
    .A(_1483_),
    .X(_1507_));
 sg13g2_nand2_1 _4734_ (.Y(_1508_),
    .A(_1449_),
    .B(_1456_));
 sg13g2_nand2b_1 _4735_ (.Y(_1509_),
    .B(_1508_),
    .A_N(_1507_));
 sg13g2_xnor2_1 _4736_ (.Y(_1510_),
    .A(_1507_),
    .B(_1508_));
 sg13g2_o21ai_1 _4737_ (.B1(_1463_),
    .Y(_1511_),
    .A1(_1464_),
    .A2(_1467_));
 sg13g2_nand2_1 _4738_ (.Y(_1512_),
    .A(_1510_),
    .B(_1511_));
 sg13g2_xnor2_1 _4739_ (.Y(_1513_),
    .A(_1510_),
    .B(_1511_));
 sg13g2_xor2_1 _4740_ (.B(_1513_),
    .A(_1482_),
    .X(\tt_um_mult_inst.genblk1[0].carry_q[0] ));
 sg13g2_o21ai_1 _4741_ (.B1(_1512_),
    .Y(_1514_),
    .A1(_1482_),
    .A2(_1513_));
 sg13g2_nand2_1 _4742_ (.Y(_1515_),
    .A(_1490_),
    .B(_1495_));
 sg13g2_nor3_1 _4743_ (.A(_1490_),
    .B(_1493_),
    .C(_1495_),
    .Y(_1516_));
 sg13g2_a21oi_1 _4744_ (.A1(_1490_),
    .A2(_1495_),
    .Y(_1517_),
    .B1(_1516_));
 sg13g2_a21o_1 _4745_ (.A2(_1499_),
    .A1(_1487_),
    .B1(_1498_),
    .X(_1518_));
 sg13g2_or2_1 _4746_ (.X(_1519_),
    .B(_1518_),
    .A(_1517_));
 sg13g2_a21oi_1 _4747_ (.A1(_1517_),
    .A2(_1518_),
    .Y(_1520_),
    .B1(net429));
 sg13g2_a22oi_1 _4748_ (.Y(_1521_),
    .B1(_1519_),
    .B2(_1520_),
    .A2(net429),
    .A1(\tt_um_mult_inst.genblk1[0].carry[2] ));
 sg13g2_nor2_1 _4749_ (.A(_1502_),
    .B(_1521_),
    .Y(_1522_));
 sg13g2_xnor2_1 _4750_ (.Y(_1523_),
    .A(_1502_),
    .B(_1521_));
 sg13g2_a21o_1 _4751_ (.A2(_1506_),
    .A1(_1504_),
    .B1(_1523_),
    .X(_1524_));
 sg13g2_nand3_1 _4752_ (.B(_1506_),
    .C(_1523_),
    .A(_1504_),
    .Y(_1525_));
 sg13g2_nand2_1 _4753_ (.Y(_1526_),
    .A(_1524_),
    .B(_1525_));
 sg13g2_nor2_1 _4754_ (.A(_1509_),
    .B(_1526_),
    .Y(_1527_));
 sg13g2_xor2_1 _4755_ (.B(_1526_),
    .A(_1509_),
    .X(_1528_));
 sg13g2_xor2_1 _4756_ (.B(_1528_),
    .A(_1514_),
    .X(\tt_um_mult_inst.genblk1[0].carry_q[1] ));
 sg13g2_a22oi_1 _4757_ (.Y(_1529_),
    .B1(_1515_),
    .B2(_1520_),
    .A2(net430),
    .A1(net921));
 sg13g2_xnor2_1 _4758_ (.Y(_1530_),
    .A(_1522_),
    .B(_1529_));
 sg13g2_nor2_1 _4759_ (.A(_1524_),
    .B(_1530_),
    .Y(_1531_));
 sg13g2_xor2_1 _4760_ (.B(_1530_),
    .A(_1524_),
    .X(_1532_));
 sg13g2_a21oi_1 _4761_ (.A1(_1514_),
    .A2(_1528_),
    .Y(_1533_),
    .B1(_1527_));
 sg13g2_nand2b_1 _4762_ (.Y(_1534_),
    .B(_1532_),
    .A_N(_1533_));
 sg13g2_xnor2_1 _4763_ (.Y(\tt_um_mult_inst.genblk1[0].carry_q[2] ),
    .A(_1532_),
    .B(_1533_));
 sg13g2_a21oi_1 _4764_ (.A1(_1522_),
    .A2(_1529_),
    .Y(_1535_),
    .B1(_1531_));
 sg13g2_nand2_1 _4765_ (.Y(\tt_um_mult_inst.genblk1[0].carry_q[3] ),
    .A(_1534_),
    .B(_1535_));
 sg13g2_a21oi_1 _4766_ (.A1(net539),
    .A2(\load_weights[176] ),
    .Y(_1536_),
    .B1(\load_weights[188] ));
 sg13g2_a21o_1 _4767_ (.A2(\load_weights[188] ),
    .A1(net539),
    .B1(_1536_),
    .X(_1537_));
 sg13g2_a21oi_1 _4768_ (.A1(net553),
    .A2(\load_weights[173] ),
    .Y(_1538_),
    .B1(\load_weights[185] ));
 sg13g2_a21o_1 _4769_ (.A2(\load_weights[185] ),
    .A1(net553),
    .B1(_1538_),
    .X(_1539_));
 sg13g2_xor2_1 _4770_ (.B(_1539_),
    .A(_1537_),
    .X(_1540_));
 sg13g2_a21oi_1 _4771_ (.A1(net516),
    .A2(\load_weights[169] ),
    .Y(_1541_),
    .B1(\load_weights[181] ));
 sg13g2_a21oi_1 _4772_ (.A1(net516),
    .A2(\load_weights[181] ),
    .Y(_1542_),
    .B1(_1541_));
 sg13g2_nand2_1 _4773_ (.Y(_1543_),
    .A(_1540_),
    .B(_1542_));
 sg13g2_xnor2_1 _4774_ (.Y(_1544_),
    .A(_1540_),
    .B(_1542_));
 sg13g2_inv_1 _4775_ (.Y(_1545_),
    .A(_1544_));
 sg13g2_a21oi_1 _4776_ (.A1(net521),
    .A2(\load_weights[168] ),
    .Y(_1546_),
    .B1(\load_weights[180] ));
 sg13g2_a21o_1 _4777_ (.A2(\load_weights[180] ),
    .A1(net521),
    .B1(_1546_),
    .X(_1547_));
 sg13g2_a21oi_1 _4778_ (.A1(net511),
    .A2(\load_weights[170] ),
    .Y(_1548_),
    .B1(\load_weights[182] ));
 sg13g2_a21o_1 _4779_ (.A2(\load_weights[182] ),
    .A1(net511),
    .B1(_1548_),
    .X(_1549_));
 sg13g2_xor2_1 _4780_ (.B(_1549_),
    .A(_1547_),
    .X(_1550_));
 sg13g2_a21oi_1 _4781_ (.A1(net531),
    .A2(\load_weights[178] ),
    .Y(_1551_),
    .B1(\load_weights[190] ));
 sg13g2_a21o_1 _4782_ (.A2(\load_weights[190] ),
    .A1(net530),
    .B1(_1551_),
    .X(_1552_));
 sg13g2_inv_1 _4783_ (.Y(_1553_),
    .A(_1552_));
 sg13g2_nand2_1 _4784_ (.Y(_1554_),
    .A(_1550_),
    .B(_1553_));
 sg13g2_nand2b_1 _4785_ (.Y(_1555_),
    .B(_1552_),
    .A_N(_1550_));
 sg13g2_nand2_1 _4786_ (.Y(_1556_),
    .A(_1550_),
    .B(_1552_));
 sg13g2_nand2b_1 _4787_ (.Y(_1557_),
    .B(_1553_),
    .A_N(_1550_));
 sg13g2_nand2_1 _4788_ (.Y(_1558_),
    .A(_1554_),
    .B(_1555_));
 sg13g2_inv_1 _4789_ (.Y(_1559_),
    .A(_1558_));
 sg13g2_nand2_1 _4790_ (.Y(_1560_),
    .A(\load_weights[180] ),
    .B(\load_weights[181] ));
 sg13g2_xnor2_1 _4791_ (.Y(_1561_),
    .A(\load_weights[180] ),
    .B(\load_weights[181] ));
 sg13g2_and2_1 _4792_ (.A(\load_weights[182] ),
    .B(\load_weights[183] ),
    .X(_1562_));
 sg13g2_xor2_1 _4793_ (.B(\load_weights[183] ),
    .A(\load_weights[182] ),
    .X(_1563_));
 sg13g2_xnor2_1 _4794_ (.Y(_1564_),
    .A(\load_weights[185] ),
    .B(_1563_));
 sg13g2_nor2_1 _4795_ (.A(_1561_),
    .B(_1564_),
    .Y(_1565_));
 sg13g2_xnor2_1 _4796_ (.Y(_1566_),
    .A(_1561_),
    .B(_1564_));
 sg13g2_and2_1 _4797_ (.A(\load_weights[187] ),
    .B(\load_weights[189] ),
    .X(_1567_));
 sg13g2_xor2_1 _4798_ (.B(\load_weights[189] ),
    .A(\load_weights[187] ),
    .X(_1568_));
 sg13g2_xnor2_1 _4799_ (.Y(_1569_),
    .A(\load_weights[191] ),
    .B(_1568_));
 sg13g2_nor2_1 _4800_ (.A(_1566_),
    .B(_1569_),
    .Y(_1570_));
 sg13g2_xor2_1 _4801_ (.B(_1569_),
    .A(_1566_),
    .X(_1571_));
 sg13g2_nand2_1 _4802_ (.Y(_1572_),
    .A(\load_weights[188] ),
    .B(_1571_));
 sg13g2_xnor2_1 _4803_ (.Y(_1573_),
    .A(\load_weights[188] ),
    .B(_1571_));
 sg13g2_xnor2_1 _4804_ (.Y(_1574_),
    .A(\load_weights[190] ),
    .B(_1573_));
 sg13g2_nand2_1 _4805_ (.Y(_1575_),
    .A(\load_weights[186] ),
    .B(_1574_));
 sg13g2_xor2_1 _4806_ (.B(_1574_),
    .A(\load_weights[186] ),
    .X(_1576_));
 sg13g2_xnor2_1 _4807_ (.Y(_1577_),
    .A(\load_weights[186] ),
    .B(_1574_));
 sg13g2_nand2_1 _4808_ (.Y(_1578_),
    .A(\load_weights[184] ),
    .B(_1576_));
 sg13g2_a21oi_1 _4809_ (.A1(_1960_),
    .A2(_1577_),
    .Y(_1579_),
    .B1(net424));
 sg13g2_xnor2_1 _4810_ (.Y(_1580_),
    .A(\load_weights[184] ),
    .B(_1576_));
 sg13g2_nor2_1 _4811_ (.A(_1961_),
    .B(net437),
    .Y(_1581_));
 sg13g2_a221oi_1 _4812_ (.B2(net437),
    .C1(_1581_),
    .B1(_1580_),
    .A1(_1556_),
    .Y(_1582_),
    .A2(_1557_));
 sg13g2_a221oi_1 _4813_ (.B2(_1579_),
    .C1(_1559_),
    .B1(_1578_),
    .A1(_1961_),
    .Y(_1583_),
    .A2(net424));
 sg13g2_a221oi_1 _4814_ (.B2(_1579_),
    .C1(_1558_),
    .B1(_1578_),
    .A1(_1961_),
    .Y(_1584_),
    .A2(net424));
 sg13g2_a221oi_1 _4815_ (.B2(net437),
    .C1(_1581_),
    .B1(_1580_),
    .A1(_1554_),
    .Y(_1585_),
    .A2(_1555_));
 sg13g2_nor3_1 _4816_ (.A(_1544_),
    .B(_1582_),
    .C(_1583_),
    .Y(_1586_));
 sg13g2_o21ai_1 _4817_ (.B1(_1545_),
    .Y(_1587_),
    .A1(_1584_),
    .A2(_1585_));
 sg13g2_nor3_1 _4818_ (.A(_1545_),
    .B(_1584_),
    .C(_1585_),
    .Y(_1588_));
 sg13g2_o21ai_1 _4819_ (.B1(_1544_),
    .Y(_1589_),
    .A1(_1582_),
    .A2(_1583_));
 sg13g2_a21oi_1 _4820_ (.A1(net506),
    .A2(\load_weights[171] ),
    .Y(_1590_),
    .B1(\load_weights[183] ));
 sg13g2_a21oi_1 _4821_ (.A1(net506),
    .A2(\load_weights[183] ),
    .Y(_1591_),
    .B1(_1590_));
 sg13g2_a21o_1 _4822_ (.A2(\load_weights[183] ),
    .A1(net506),
    .B1(_1590_),
    .X(_1592_));
 sg13g2_nor3_1 _4823_ (.A(_1586_),
    .B(_1588_),
    .C(_1592_),
    .Y(_1593_));
 sg13g2_nand3_1 _4824_ (.B(_1589_),
    .C(_1591_),
    .A(_1587_),
    .Y(_1594_));
 sg13g2_a21oi_1 _4825_ (.A1(_1587_),
    .A2(_1589_),
    .Y(_1595_),
    .B1(_1591_));
 sg13g2_o21ai_1 _4826_ (.B1(_1592_),
    .Y(_1596_),
    .A1(_1586_),
    .A2(_1588_));
 sg13g2_a21oi_1 _4827_ (.A1(net548),
    .A2(\load_weights[174] ),
    .Y(_1597_),
    .B1(\load_weights[186] ));
 sg13g2_a21oi_1 _4828_ (.A1(net548),
    .A2(\load_weights[186] ),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_a21o_1 _4829_ (.A2(\load_weights[186] ),
    .A1(net548),
    .B1(_1597_),
    .X(_1599_));
 sg13g2_nor3_1 _4830_ (.A(_1593_),
    .B(_1595_),
    .C(_1599_),
    .Y(_1600_));
 sg13g2_nand3_1 _4831_ (.B(_1596_),
    .C(_1598_),
    .A(_1594_),
    .Y(_1601_));
 sg13g2_a21oi_1 _4832_ (.A1(_1594_),
    .A2(_1596_),
    .Y(_1602_),
    .B1(_1598_));
 sg13g2_o21ai_1 _4833_ (.B1(_1599_),
    .Y(_1603_),
    .A1(_1593_),
    .A2(_1595_));
 sg13g2_a21oi_1 _4834_ (.A1(net544),
    .A2(\load_weights[175] ),
    .Y(_1604_),
    .B1(\load_weights[187] ));
 sg13g2_a21oi_2 _4835_ (.B1(_1604_),
    .Y(_1605_),
    .A2(\load_weights[187] ),
    .A1(net544));
 sg13g2_a21o_1 _4836_ (.A2(\load_weights[187] ),
    .A1(net544),
    .B1(_1604_),
    .X(_1606_));
 sg13g2_nor3_1 _4837_ (.A(_1600_),
    .B(_1602_),
    .C(_1606_),
    .Y(_1607_));
 sg13g2_nand3_1 _4838_ (.B(_1603_),
    .C(_1605_),
    .A(_1601_),
    .Y(_1608_));
 sg13g2_a21oi_1 _4839_ (.A1(_1601_),
    .A2(_1603_),
    .Y(_1609_),
    .B1(_1605_));
 sg13g2_o21ai_1 _4840_ (.B1(_1606_),
    .Y(_1610_),
    .A1(_1600_),
    .A2(_1602_));
 sg13g2_a21oi_1 _4841_ (.A1(net559),
    .A2(\load_weights[172] ),
    .Y(_1611_),
    .B1(\load_weights[184] ));
 sg13g2_a21o_1 _4842_ (.A2(\load_weights[184] ),
    .A1(net559),
    .B1(_1611_),
    .X(_1612_));
 sg13g2_inv_1 _4843_ (.Y(_1613_),
    .A(_1612_));
 sg13g2_nor3_1 _4844_ (.A(_1607_),
    .B(_1609_),
    .C(_1612_),
    .Y(_1614_));
 sg13g2_a21oi_1 _4845_ (.A1(_1608_),
    .A2(_1610_),
    .Y(_1615_),
    .B1(_1613_));
 sg13g2_nand3_1 _4846_ (.B(_1610_),
    .C(_1612_),
    .A(_1608_),
    .Y(_1616_));
 sg13g2_o21ai_1 _4847_ (.B1(_1613_),
    .Y(_1617_),
    .A1(_1607_),
    .A2(_1609_));
 sg13g2_a21oi_1 _4848_ (.A1(net536),
    .A2(\load_weights[177] ),
    .Y(_1618_),
    .B1(\load_weights[189] ));
 sg13g2_a21o_2 _4849_ (.A2(\load_weights[189] ),
    .A1(net536),
    .B1(_1618_),
    .X(_1619_));
 sg13g2_nor3_2 _4850_ (.A(_1614_),
    .B(_1615_),
    .C(_1619_),
    .Y(_1620_));
 sg13g2_and3_1 _4851_ (.X(_1621_),
    .A(_1616_),
    .B(_1617_),
    .C(_1619_));
 sg13g2_o21ai_1 _4852_ (.B1(_1619_),
    .Y(_1622_),
    .A1(_1614_),
    .A2(_1615_));
 sg13g2_a21oi_1 _4853_ (.A1(net527),
    .A2(\load_weights[179] ),
    .Y(_1623_),
    .B1(\load_weights[191] ));
 sg13g2_a21oi_2 _4854_ (.B1(_1623_),
    .Y(_1624_),
    .A2(\load_weights[191] ),
    .A1(net527));
 sg13g2_nor3_1 _4855_ (.A(_1620_),
    .B(_1621_),
    .C(_1624_),
    .Y(_1625_));
 sg13g2_o21ai_1 _4856_ (.B1(_1624_),
    .Y(_1626_),
    .A1(_1620_),
    .A2(_1621_));
 sg13g2_nand2b_2 _4857_ (.Y(\tt_um_mult_inst.genblk1[7].out_q ),
    .B(_1626_),
    .A_N(_1625_));
 sg13g2_a21oi_2 _4858_ (.B1(_1620_),
    .Y(_1627_),
    .A2(_1624_),
    .A1(_1622_));
 sg13g2_o21ai_1 _4859_ (.B1(_1543_),
    .Y(_1628_),
    .A1(_1537_),
    .A2(_1539_));
 sg13g2_nand2b_1 _4860_ (.Y(_1629_),
    .B(_1587_),
    .A_N(_1582_));
 sg13g2_o21ai_1 _4861_ (.B1(_1554_),
    .Y(_1630_),
    .A1(_1547_),
    .A2(_1549_));
 sg13g2_nand2_1 _4862_ (.Y(_1631_),
    .A(\tt_um_mult_inst.genblk1[7].carry[1] ),
    .B(net425));
 sg13g2_nand2_1 _4863_ (.Y(_1632_),
    .A(_1575_),
    .B(_1578_));
 sg13g2_a21oi_2 _4864_ (.B1(_1567_),
    .Y(_1633_),
    .A2(_1568_),
    .A1(\load_weights[191] ));
 sg13g2_a21oi_1 _4865_ (.A1(\load_weights[185] ),
    .A2(_1563_),
    .Y(_1634_),
    .B1(_1562_));
 sg13g2_nor2_1 _4866_ (.A(_1560_),
    .B(_1634_),
    .Y(_1635_));
 sg13g2_xnor2_1 _4867_ (.Y(_1636_),
    .A(_1560_),
    .B(_1634_));
 sg13g2_nor2_1 _4868_ (.A(_1565_),
    .B(_1570_),
    .Y(_1637_));
 sg13g2_nor2_1 _4869_ (.A(_1636_),
    .B(_1637_),
    .Y(_1638_));
 sg13g2_xnor2_1 _4870_ (.Y(_1639_),
    .A(_1636_),
    .B(_1637_));
 sg13g2_nor2_1 _4871_ (.A(_1633_),
    .B(_1639_),
    .Y(_1640_));
 sg13g2_xor2_1 _4872_ (.B(_1639_),
    .A(_1633_),
    .X(_1641_));
 sg13g2_o21ai_1 _4873_ (.B1(_1572_),
    .Y(_1642_),
    .A1(_1959_),
    .A2(_1573_));
 sg13g2_and2_1 _4874_ (.A(_1641_),
    .B(_1642_),
    .X(_1643_));
 sg13g2_xor2_1 _4875_ (.B(_1642_),
    .A(_1641_),
    .X(_1644_));
 sg13g2_xnor2_1 _4876_ (.Y(_1645_),
    .A(_1632_),
    .B(_1644_));
 sg13g2_o21ai_1 _4877_ (.B1(_1631_),
    .Y(_1646_),
    .A1(net425),
    .A2(_1645_));
 sg13g2_nand2_1 _4878_ (.Y(_1647_),
    .A(_1630_),
    .B(_1646_));
 sg13g2_xor2_1 _4879_ (.B(_1646_),
    .A(_1630_),
    .X(_1648_));
 sg13g2_nand2_1 _4880_ (.Y(_1649_),
    .A(_1629_),
    .B(_1648_));
 sg13g2_xnor2_1 _4881_ (.Y(_1650_),
    .A(_1629_),
    .B(_1648_));
 sg13g2_nand2b_1 _4882_ (.Y(_1651_),
    .B(_1628_),
    .A_N(_1650_));
 sg13g2_xor2_1 _4883_ (.B(_1650_),
    .A(_1628_),
    .X(_1652_));
 sg13g2_nand2_1 _4884_ (.Y(_1653_),
    .A(_1594_),
    .B(_1601_));
 sg13g2_nand2b_1 _4885_ (.Y(_1654_),
    .B(_1653_),
    .A_N(_1652_));
 sg13g2_xnor2_1 _4886_ (.Y(_1655_),
    .A(_1652_),
    .B(_1653_));
 sg13g2_o21ai_1 _4887_ (.B1(_1608_),
    .Y(_1656_),
    .A1(_1609_),
    .A2(_1612_));
 sg13g2_nand2_1 _4888_ (.Y(_1657_),
    .A(_1655_),
    .B(_1656_));
 sg13g2_xnor2_1 _4889_ (.Y(_1658_),
    .A(_1655_),
    .B(_1656_));
 sg13g2_xor2_1 _4890_ (.B(_1658_),
    .A(_1627_),
    .X(\tt_um_mult_inst.genblk1[7].carry_q[0] ));
 sg13g2_o21ai_1 _4891_ (.B1(_1657_),
    .Y(_1659_),
    .A1(_1627_),
    .A2(_1658_));
 sg13g2_nand2_1 _4892_ (.Y(_1660_),
    .A(_1635_),
    .B(_1640_));
 sg13g2_nor3_1 _4893_ (.A(_1635_),
    .B(_1638_),
    .C(_1640_),
    .Y(_1661_));
 sg13g2_a21oi_1 _4894_ (.A1(_1635_),
    .A2(_1640_),
    .Y(_1662_),
    .B1(_1661_));
 sg13g2_a21o_1 _4895_ (.A2(_1644_),
    .A1(_1632_),
    .B1(_1643_),
    .X(_1663_));
 sg13g2_or2_1 _4896_ (.X(_1664_),
    .B(_1663_),
    .A(_1662_));
 sg13g2_a21oi_1 _4897_ (.A1(_1662_),
    .A2(_1663_),
    .Y(_1665_),
    .B1(net425));
 sg13g2_a22oi_1 _4898_ (.Y(_1666_),
    .B1(_1664_),
    .B2(_1665_),
    .A2(net425),
    .A1(\tt_um_mult_inst.genblk1[7].carry[2] ));
 sg13g2_nor2_1 _4899_ (.A(_1647_),
    .B(_1666_),
    .Y(_1667_));
 sg13g2_xnor2_1 _4900_ (.Y(_1668_),
    .A(_1647_),
    .B(_1666_));
 sg13g2_a21o_1 _4901_ (.A2(_1651_),
    .A1(_1649_),
    .B1(_1668_),
    .X(_1669_));
 sg13g2_nand3_1 _4902_ (.B(_1651_),
    .C(_1668_),
    .A(_1649_),
    .Y(_1670_));
 sg13g2_nand2_1 _4903_ (.Y(_1671_),
    .A(_1669_),
    .B(_1670_));
 sg13g2_nor2_1 _4904_ (.A(_1654_),
    .B(_1671_),
    .Y(_1672_));
 sg13g2_xor2_1 _4905_ (.B(_1671_),
    .A(_1654_),
    .X(_1673_));
 sg13g2_xor2_1 _4906_ (.B(_1673_),
    .A(_1659_),
    .X(\tt_um_mult_inst.genblk1[7].carry_q[1] ));
 sg13g2_a22oi_1 _4907_ (.Y(_1674_),
    .B1(_1660_),
    .B2(_1665_),
    .A2(net425),
    .A1(net925));
 sg13g2_xnor2_1 _4908_ (.Y(_1675_),
    .A(_1667_),
    .B(_1674_));
 sg13g2_nor2_1 _4909_ (.A(_1669_),
    .B(_1675_),
    .Y(_1676_));
 sg13g2_xor2_1 _4910_ (.B(_1675_),
    .A(_1669_),
    .X(_1677_));
 sg13g2_a21oi_1 _4911_ (.A1(_1659_),
    .A2(_1673_),
    .Y(_1678_),
    .B1(_1672_));
 sg13g2_nand2b_1 _4912_ (.Y(_1679_),
    .B(_1677_),
    .A_N(_1678_));
 sg13g2_xnor2_1 _4913_ (.Y(\tt_um_mult_inst.genblk1[7].carry_q[2] ),
    .A(_1677_),
    .B(_1678_));
 sg13g2_a21oi_1 _4914_ (.A1(_1667_),
    .A2(_1674_),
    .Y(_1680_),
    .B1(_1676_));
 sg13g2_nand2_1 _4915_ (.Y(\tt_um_mult_inst.genblk1[7].carry_q[3] ),
    .A(_1679_),
    .B(_1680_));
 sg13g2_a21oi_1 _4916_ (.A1(net536),
    .A2(\load_weights[57] ),
    .Y(_1681_),
    .B1(\load_weights[69] ));
 sg13g2_a21o_1 _4917_ (.A2(\load_weights[69] ),
    .A1(net535),
    .B1(_1681_),
    .X(_1682_));
 sg13g2_a21oi_1 _4918_ (.A1(net560),
    .A2(\load_weights[52] ),
    .Y(_1683_),
    .B1(\load_weights[64] ));
 sg13g2_a21o_1 _4919_ (.A2(\load_weights[64] ),
    .A1(net560),
    .B1(_1683_),
    .X(_1684_));
 sg13g2_xor2_1 _4920_ (.B(_1684_),
    .A(_1682_),
    .X(_1685_));
 sg13g2_a21oi_1 _4921_ (.A1(net513),
    .A2(\load_weights[50] ),
    .Y(_1686_),
    .B1(\load_weights[62] ));
 sg13g2_a21oi_1 _4922_ (.A1(net513),
    .A2(\load_weights[62] ),
    .Y(_1687_),
    .B1(_1686_));
 sg13g2_nand2_1 _4923_ (.Y(_1688_),
    .A(_1685_),
    .B(_1687_));
 sg13g2_xnor2_1 _4924_ (.Y(_1689_),
    .A(_1685_),
    .B(_1687_));
 sg13g2_inv_1 _4925_ (.Y(_1690_),
    .A(_1689_));
 sg13g2_a21oi_1 _4926_ (.A1(net550),
    .A2(\load_weights[54] ),
    .Y(_1691_),
    .B1(\load_weights[66] ));
 sg13g2_a21o_1 _4927_ (.A2(\load_weights[66] ),
    .A1(net550),
    .B1(_1691_),
    .X(_1692_));
 sg13g2_a21oi_1 _4928_ (.A1(net555),
    .A2(\load_weights[53] ),
    .Y(_1693_),
    .B1(\load_weights[65] ));
 sg13g2_a21o_1 _4929_ (.A2(\load_weights[65] ),
    .A1(net554),
    .B1(_1693_),
    .X(_1694_));
 sg13g2_xor2_1 _4930_ (.B(_1694_),
    .A(_1692_),
    .X(_1695_));
 sg13g2_a21oi_1 _4931_ (.A1(net526),
    .A2(\load_weights[59] ),
    .Y(_1696_),
    .B1(\load_weights[71] ));
 sg13g2_a21o_1 _4932_ (.A2(\load_weights[71] ),
    .A1(net526),
    .B1(_1696_),
    .X(_1697_));
 sg13g2_inv_1 _4933_ (.Y(_1698_),
    .A(_1697_));
 sg13g2_nand2_1 _4934_ (.Y(_1699_),
    .A(_1695_),
    .B(_1698_));
 sg13g2_nand2b_1 _4935_ (.Y(_1700_),
    .B(_1697_),
    .A_N(_1695_));
 sg13g2_nand2_1 _4936_ (.Y(_1701_),
    .A(_1695_),
    .B(_1697_));
 sg13g2_nand2b_1 _4937_ (.Y(_1702_),
    .B(_1698_),
    .A_N(_1695_));
 sg13g2_nand2_1 _4938_ (.Y(_1703_),
    .A(_1699_),
    .B(_1700_));
 sg13g2_inv_1 _4939_ (.Y(_1704_),
    .A(_1703_));
 sg13g2_and2_1 _4940_ (.A(\load_weights[60] ),
    .B(\load_weights[61] ),
    .X(_1705_));
 sg13g2_xor2_1 _4941_ (.B(\load_weights[61] ),
    .A(\load_weights[60] ),
    .X(_1706_));
 sg13g2_xnor2_1 _4942_ (.Y(_1707_),
    .A(\load_weights[62] ),
    .B(_1706_));
 sg13g2_inv_1 _4943_ (.Y(_1708_),
    .A(_1707_));
 sg13g2_nand2_1 _4944_ (.Y(_1709_),
    .A(\load_weights[64] ),
    .B(_1708_));
 sg13g2_xor2_1 _4945_ (.B(_1707_),
    .A(\load_weights[64] ),
    .X(_1710_));
 sg13g2_xor2_1 _4946_ (.B(_1710_),
    .A(_0020_),
    .X(_1711_));
 sg13g2_and2_1 _4947_ (.A(\load_weights[66] ),
    .B(\load_weights[68] ),
    .X(_1712_));
 sg13g2_xor2_1 _4948_ (.B(\load_weights[68] ),
    .A(\load_weights[66] ),
    .X(_1713_));
 sg13g2_xor2_1 _4949_ (.B(_1713_),
    .A(\load_weights[70] ),
    .X(_1714_));
 sg13g2_nand2_1 _4950_ (.Y(_1715_),
    .A(_1711_),
    .B(_1714_));
 sg13g2_xnor2_1 _4951_ (.Y(_1716_),
    .A(_1711_),
    .B(_1714_));
 sg13g2_inv_1 _4952_ (.Y(_1717_),
    .A(_1716_));
 sg13g2_xor2_1 _4953_ (.B(_1716_),
    .A(\load_weights[67] ),
    .X(_1718_));
 sg13g2_nor2_1 _4954_ (.A(_1962_),
    .B(_1718_),
    .Y(_1719_));
 sg13g2_xnor2_1 _4955_ (.Y(_1720_),
    .A(\load_weights[69] ),
    .B(_1718_));
 sg13g2_nand2_1 _4956_ (.Y(_1721_),
    .A(\load_weights[65] ),
    .B(_1720_));
 sg13g2_xor2_1 _4957_ (.B(_1720_),
    .A(\load_weights[65] ),
    .X(_1722_));
 sg13g2_xnor2_1 _4958_ (.Y(_1723_),
    .A(\load_weights[65] ),
    .B(_1720_));
 sg13g2_nand2_1 _4959_ (.Y(_1724_),
    .A(\load_weights[63] ),
    .B(_1722_));
 sg13g2_a21oi_1 _4960_ (.A1(_1963_),
    .A2(_1723_),
    .Y(_1725_),
    .B1(net428));
 sg13g2_xnor2_1 _4961_ (.Y(_1726_),
    .A(\load_weights[63] ),
    .B(_1722_));
 sg13g2_nor2_1 _4962_ (.A(_1964_),
    .B(net439),
    .Y(_1727_));
 sg13g2_a221oi_1 _4963_ (.B2(net439),
    .C1(_1727_),
    .B1(_1726_),
    .A1(_1701_),
    .Y(_1728_),
    .A2(_1702_));
 sg13g2_a221oi_1 _4964_ (.B2(_1725_),
    .C1(_1704_),
    .B1(_1724_),
    .A1(_1964_),
    .Y(_1729_),
    .A2(net428));
 sg13g2_a221oi_1 _4965_ (.B2(_1725_),
    .C1(_1703_),
    .B1(_1724_),
    .A1(_1964_),
    .Y(_1730_),
    .A2(net428));
 sg13g2_a221oi_1 _4966_ (.B2(net439),
    .C1(_1727_),
    .B1(_1726_),
    .A1(_1699_),
    .Y(_1731_),
    .A2(_1700_));
 sg13g2_nor3_1 _4967_ (.A(_1689_),
    .B(_1728_),
    .C(_1729_),
    .Y(_1732_));
 sg13g2_o21ai_1 _4968_ (.B1(_1690_),
    .Y(_1733_),
    .A1(_1730_),
    .A2(_1731_));
 sg13g2_nor3_1 _4969_ (.A(_1690_),
    .B(_1730_),
    .C(_1731_),
    .Y(_1734_));
 sg13g2_o21ai_1 _4970_ (.B1(_1689_),
    .Y(_1735_),
    .A1(_1728_),
    .A2(_1729_));
 sg13g2_a21oi_1 _4971_ (.A1(net505),
    .A2(\load_weights[51] ),
    .Y(_1736_),
    .B1(\load_weights[63] ));
 sg13g2_a21oi_1 _4972_ (.A1(net505),
    .A2(\load_weights[63] ),
    .Y(_1737_),
    .B1(_1736_));
 sg13g2_a21o_1 _4973_ (.A2(\load_weights[63] ),
    .A1(net505),
    .B1(_1736_),
    .X(_1738_));
 sg13g2_nor3_1 _4974_ (.A(_1732_),
    .B(_1734_),
    .C(_1738_),
    .Y(_1739_));
 sg13g2_nand3_1 _4975_ (.B(_1735_),
    .C(_1737_),
    .A(_1733_),
    .Y(_1740_));
 sg13g2_a21oi_1 _4976_ (.A1(_1733_),
    .A2(_1735_),
    .Y(_1741_),
    .B1(_1737_));
 sg13g2_o21ai_1 _4977_ (.B1(_1738_),
    .Y(_1742_),
    .A1(_1732_),
    .A2(_1734_));
 sg13g2_a21oi_1 _4978_ (.A1(net518),
    .A2(\load_weights[49] ),
    .Y(_1743_),
    .B1(\load_weights[61] ));
 sg13g2_a21oi_1 _4979_ (.A1(net518),
    .A2(\load_weights[61] ),
    .Y(_1744_),
    .B1(_1743_));
 sg13g2_a21o_1 _4980_ (.A2(\load_weights[61] ),
    .A1(net518),
    .B1(_1743_),
    .X(_1745_));
 sg13g2_nor3_1 _4981_ (.A(_1739_),
    .B(_1741_),
    .C(_1745_),
    .Y(_1746_));
 sg13g2_nand3_1 _4982_ (.B(_1742_),
    .C(_1744_),
    .A(_1740_),
    .Y(_1747_));
 sg13g2_a21oi_1 _4983_ (.A1(_1740_),
    .A2(_1742_),
    .Y(_1748_),
    .B1(_1744_));
 sg13g2_o21ai_1 _4984_ (.B1(_1745_),
    .Y(_1749_),
    .A1(_1739_),
    .A2(_1741_));
 sg13g2_a21oi_1 _4985_ (.A1(net541),
    .A2(\load_weights[56] ),
    .Y(_1750_),
    .B1(\load_weights[68] ));
 sg13g2_a21oi_1 _4986_ (.A1(net541),
    .A2(\load_weights[68] ),
    .Y(_1751_),
    .B1(_1750_));
 sg13g2_a21o_1 _4987_ (.A2(\load_weights[68] ),
    .A1(net541),
    .B1(_1750_),
    .X(_1752_));
 sg13g2_nor3_1 _4988_ (.A(_1746_),
    .B(_1748_),
    .C(_1752_),
    .Y(_1753_));
 sg13g2_nand3_1 _4989_ (.B(_1749_),
    .C(_1751_),
    .A(_1747_),
    .Y(_1754_));
 sg13g2_a21oi_1 _4990_ (.A1(_1747_),
    .A2(_1749_),
    .Y(_1755_),
    .B1(_1751_));
 sg13g2_o21ai_1 _4991_ (.B1(_1752_),
    .Y(_1756_),
    .A1(_1746_),
    .A2(_1748_));
 sg13g2_a21oi_1 _4992_ (.A1(net525),
    .A2(\load_weights[48] ),
    .Y(_1757_),
    .B1(\load_weights[60] ));
 sg13g2_a21o_1 _4993_ (.A2(\load_weights[60] ),
    .A1(net525),
    .B1(_1757_),
    .X(_1758_));
 sg13g2_inv_1 _4994_ (.Y(_1759_),
    .A(_1758_));
 sg13g2_nor3_1 _4995_ (.A(_1753_),
    .B(_1755_),
    .C(_1758_),
    .Y(_1760_));
 sg13g2_a21oi_1 _4996_ (.A1(_1754_),
    .A2(_1756_),
    .Y(_1761_),
    .B1(_1759_));
 sg13g2_nand3_1 _4997_ (.B(_1756_),
    .C(_1758_),
    .A(_1754_),
    .Y(_1762_));
 sg13g2_o21ai_1 _4998_ (.B1(_1759_),
    .Y(_1763_),
    .A1(_1753_),
    .A2(_1755_));
 sg13g2_a21oi_1 _4999_ (.A1(net532),
    .A2(\load_weights[58] ),
    .Y(_1764_),
    .B1(\load_weights[70] ));
 sg13g2_a21o_1 _5000_ (.A2(\load_weights[70] ),
    .A1(net532),
    .B1(_1764_),
    .X(_1765_));
 sg13g2_nor3_1 _5001_ (.A(_1760_),
    .B(_1761_),
    .C(_1765_),
    .Y(_1766_));
 sg13g2_and3_1 _5002_ (.X(_1767_),
    .A(_1762_),
    .B(_1763_),
    .C(_1765_));
 sg13g2_o21ai_1 _5003_ (.B1(_1765_),
    .Y(_1768_),
    .A1(_1760_),
    .A2(_1761_));
 sg13g2_a21oi_1 _5004_ (.A1(net546),
    .A2(net420),
    .Y(_1769_),
    .B1(net828));
 sg13g2_a21oi_2 _5005_ (.B1(_1769_),
    .Y(_1770_),
    .A2(net931),
    .A1(net546));
 sg13g2_nor3_1 _5006_ (.A(_1766_),
    .B(_1767_),
    .C(_1770_),
    .Y(_1771_));
 sg13g2_o21ai_1 _5007_ (.B1(_1770_),
    .Y(_1772_),
    .A1(_1766_),
    .A2(_1767_));
 sg13g2_nand2b_1 _5008_ (.Y(\tt_um_mult_inst.genblk1[2].out_q ),
    .B(_1772_),
    .A_N(_1771_));
 sg13g2_a21oi_1 _5009_ (.A1(_1768_),
    .A2(_1770_),
    .Y(_1773_),
    .B1(_1766_));
 sg13g2_o21ai_1 _5010_ (.B1(_1754_),
    .Y(_1774_),
    .A1(_1755_),
    .A2(_1758_));
 sg13g2_o21ai_1 _5011_ (.B1(_1688_),
    .Y(_1775_),
    .A1(_1682_),
    .A2(_1684_));
 sg13g2_nand2b_1 _5012_ (.Y(_1776_),
    .B(_1733_),
    .A_N(_1728_));
 sg13g2_o21ai_1 _5013_ (.B1(_1699_),
    .Y(_1777_),
    .A1(_1692_),
    .A2(_1694_));
 sg13g2_nor2_1 _5014_ (.A(\tt_um_mult_inst.genblk1[2].carry[1] ),
    .B(net439),
    .Y(_1778_));
 sg13g2_nand2_1 _5015_ (.Y(_1779_),
    .A(_1721_),
    .B(_1724_));
 sg13g2_a21oi_2 _5016_ (.B1(_1712_),
    .Y(_1780_),
    .A2(_1713_),
    .A1(\load_weights[70] ));
 sg13g2_and3_1 _5017_ (.X(_1781_),
    .A(\load_weights[62] ),
    .B(\load_weights[64] ),
    .C(_1705_));
 sg13g2_a21oi_1 _5018_ (.A1(\load_weights[62] ),
    .A2(_1706_),
    .Y(_1782_),
    .B1(_1705_));
 sg13g2_a21oi_1 _5019_ (.A1(_1709_),
    .A2(_1782_),
    .Y(_1783_),
    .B1(_1781_));
 sg13g2_o21ai_1 _5020_ (.B1(_1715_),
    .Y(_1784_),
    .A1(_0020_),
    .A2(_1710_));
 sg13g2_nand2_1 _5021_ (.Y(_1785_),
    .A(_1783_),
    .B(_1784_));
 sg13g2_xnor2_1 _5022_ (.Y(_1786_),
    .A(_1783_),
    .B(_1784_));
 sg13g2_xor2_1 _5023_ (.B(_1786_),
    .A(_1780_),
    .X(_1787_));
 sg13g2_a21oi_1 _5024_ (.A1(\load_weights[67] ),
    .A2(_1717_),
    .Y(_1788_),
    .B1(_1719_));
 sg13g2_nor2b_1 _5025_ (.A(_1788_),
    .B_N(_1787_),
    .Y(_1789_));
 sg13g2_xnor2_1 _5026_ (.Y(_1790_),
    .A(_1787_),
    .B(_1788_));
 sg13g2_xnor2_1 _5027_ (.Y(_1791_),
    .A(_1779_),
    .B(_1790_));
 sg13g2_a21oi_1 _5028_ (.A1(net439),
    .A2(_1791_),
    .Y(_1792_),
    .B1(_1778_));
 sg13g2_nand2_1 _5029_ (.Y(_1793_),
    .A(_1777_),
    .B(_1792_));
 sg13g2_xor2_1 _5030_ (.B(_1792_),
    .A(_1777_),
    .X(_1794_));
 sg13g2_nand2_1 _5031_ (.Y(_1795_),
    .A(_1776_),
    .B(_1794_));
 sg13g2_xnor2_1 _5032_ (.Y(_1796_),
    .A(_1776_),
    .B(_1794_));
 sg13g2_nand2b_1 _5033_ (.Y(_1797_),
    .B(_1775_),
    .A_N(_1796_));
 sg13g2_xor2_1 _5034_ (.B(_1796_),
    .A(_1775_),
    .X(_1798_));
 sg13g2_nand2_1 _5035_ (.Y(_1799_),
    .A(_1740_),
    .B(_1747_));
 sg13g2_nand2b_1 _5036_ (.Y(_1800_),
    .B(_1799_),
    .A_N(_1798_));
 sg13g2_xnor2_1 _5037_ (.Y(_1801_),
    .A(_1798_),
    .B(_1799_));
 sg13g2_nand2_1 _5038_ (.Y(_1802_),
    .A(_1774_),
    .B(_1801_));
 sg13g2_xnor2_1 _5039_ (.Y(_1803_),
    .A(_1774_),
    .B(_1801_));
 sg13g2_xor2_1 _5040_ (.B(_1803_),
    .A(_1773_),
    .X(\tt_um_mult_inst.genblk1[2].carry_q[0] ));
 sg13g2_a21o_1 _5041_ (.A2(_1790_),
    .A1(_1779_),
    .B1(_1789_),
    .X(_1804_));
 sg13g2_dfrbp_1 _5042_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net316),
    .D(_0029_),
    .Q_N(_2453_),
    .Q(\load_weights[0] ));
 sg13g2_dfrbp_1 _5043_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net86),
    .D(_0030_),
    .Q_N(_2452_),
    .Q(\load_weights[1] ));
 sg13g2_dfrbp_1 _5044_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net85),
    .D(_0031_),
    .Q_N(_2451_),
    .Q(\load_weights[2] ));
 sg13g2_dfrbp_1 _5045_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net84),
    .D(_0032_),
    .Q_N(_2450_),
    .Q(\load_weights[3] ));
 sg13g2_dfrbp_1 _5046_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net83),
    .D(_0033_),
    .Q_N(_2449_),
    .Q(\load_weights[4] ));
 sg13g2_dfrbp_1 _5047_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net82),
    .D(_0034_),
    .Q_N(_2448_),
    .Q(\load_weights[5] ));
 sg13g2_dfrbp_1 _5048_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net81),
    .D(_0035_),
    .Q_N(_2447_),
    .Q(\load_weights[6] ));
 sg13g2_dfrbp_1 _5049_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net80),
    .D(_0036_),
    .Q_N(_2446_),
    .Q(\load_weights[7] ));
 sg13g2_dfrbp_1 _5050_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net79),
    .D(_0037_),
    .Q_N(_2445_),
    .Q(\load_weights[8] ));
 sg13g2_dfrbp_1 _5051_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net78),
    .D(_0038_),
    .Q_N(_2444_),
    .Q(\load_weights[9] ));
 sg13g2_dfrbp_1 _5052_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net77),
    .D(_0039_),
    .Q_N(_2443_),
    .Q(\load_weights[10] ));
 sg13g2_dfrbp_1 _5053_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net76),
    .D(_0040_),
    .Q_N(_2442_),
    .Q(\load_weights[11] ));
 sg13g2_dfrbp_1 _5054_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net75),
    .D(net663),
    .Q_N(_2441_),
    .Q(\load_weights[12] ));
 sg13g2_dfrbp_1 _5055_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net74),
    .D(_0042_),
    .Q_N(_2440_),
    .Q(\load_weights[13] ));
 sg13g2_dfrbp_1 _5056_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net73),
    .D(_0043_),
    .Q_N(_2439_),
    .Q(\load_weights[14] ));
 sg13g2_dfrbp_1 _5057_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net72),
    .D(_0044_),
    .Q_N(_2438_),
    .Q(\load_weights[15] ));
 sg13g2_dfrbp_1 _5058_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net71),
    .D(net381),
    .Q_N(_2437_),
    .Q(\load_weights[16] ));
 sg13g2_dfrbp_1 _5059_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net70),
    .D(_0046_),
    .Q_N(_2436_),
    .Q(\load_weights[17] ));
 sg13g2_dfrbp_1 _5060_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net69),
    .D(_0047_),
    .Q_N(_2435_),
    .Q(\load_weights[18] ));
 sg13g2_dfrbp_1 _5061_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net68),
    .D(net573),
    .Q_N(_2434_),
    .Q(\load_weights[19] ));
 sg13g2_dfrbp_1 _5062_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net67),
    .D(net616),
    .Q_N(_2433_),
    .Q(\load_weights[20] ));
 sg13g2_dfrbp_1 _5063_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net66),
    .D(_0050_),
    .Q_N(_2432_),
    .Q(\load_weights[21] ));
 sg13g2_dfrbp_1 _5064_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net65),
    .D(net406),
    .Q_N(_2431_),
    .Q(\load_weights[22] ));
 sg13g2_dfrbp_1 _5065_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net64),
    .D(_0052_),
    .Q_N(_2430_),
    .Q(\load_weights[23] ));
 sg13g2_dfrbp_1 _5066_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net63),
    .D(_0053_),
    .Q_N(_2429_),
    .Q(\load_weights[24] ));
 sg13g2_dfrbp_1 _5067_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net62),
    .D(net683),
    .Q_N(_2428_),
    .Q(\load_weights[25] ));
 sg13g2_dfrbp_1 _5068_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net61),
    .D(_0055_),
    .Q_N(_2427_),
    .Q(\load_weights[26] ));
 sg13g2_dfrbp_1 _5069_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net60),
    .D(_0056_),
    .Q_N(_2426_),
    .Q(\load_weights[27] ));
 sg13g2_dfrbp_1 _5070_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net59),
    .D(net648),
    .Q_N(_2425_),
    .Q(\load_weights[28] ));
 sg13g2_dfrbp_1 _5071_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net58),
    .D(_0058_),
    .Q_N(_2424_),
    .Q(\load_weights[29] ));
 sg13g2_dfrbp_1 _5072_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net57),
    .D(_0059_),
    .Q_N(_2423_),
    .Q(\load_weights[30] ));
 sg13g2_dfrbp_1 _5073_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net56),
    .D(_0060_),
    .Q_N(_2422_),
    .Q(\load_weights[31] ));
 sg13g2_dfrbp_1 _5074_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net55),
    .D(net620),
    .Q_N(_2421_),
    .Q(\load_weights[32] ));
 sg13g2_dfrbp_1 _5075_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net54),
    .D(_0062_),
    .Q_N(_2420_),
    .Q(\load_weights[33] ));
 sg13g2_dfrbp_1 _5076_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net53),
    .D(net580),
    .Q_N(_2419_),
    .Q(\load_weights[34] ));
 sg13g2_dfrbp_1 _5077_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net52),
    .D(_0064_),
    .Q_N(_2418_),
    .Q(\load_weights[35] ));
 sg13g2_dfrbp_1 _5078_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net51),
    .D(_0065_),
    .Q_N(_2417_),
    .Q(\load_weights[36] ));
 sg13g2_dfrbp_1 _5079_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net50),
    .D(_0066_),
    .Q_N(_2416_),
    .Q(\load_weights[37] ));
 sg13g2_dfrbp_1 _5080_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net49),
    .D(_0067_),
    .Q_N(_2415_),
    .Q(\load_weights[38] ));
 sg13g2_dfrbp_1 _5081_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net48),
    .D(net387),
    .Q_N(_2414_),
    .Q(\load_weights[39] ));
 sg13g2_dfrbp_1 _5082_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net47),
    .D(_0069_),
    .Q_N(_2413_),
    .Q(\load_weights[40] ));
 sg13g2_dfrbp_1 _5083_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net46),
    .D(net385),
    .Q_N(_2412_),
    .Q(\load_weights[41] ));
 sg13g2_dfrbp_1 _5084_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net45),
    .D(_0071_),
    .Q_N(_2411_),
    .Q(\load_weights[42] ));
 sg13g2_dfrbp_1 _5085_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net44),
    .D(net417),
    .Q_N(_2410_),
    .Q(\load_weights[43] ));
 sg13g2_dfrbp_1 _5086_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net43),
    .D(_0073_),
    .Q_N(_2409_),
    .Q(\load_weights[44] ));
 sg13g2_dfrbp_1 _5087_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net42),
    .D(net712),
    .Q_N(_2408_),
    .Q(\load_weights[45] ));
 sg13g2_dfrbp_1 _5088_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net41),
    .D(_0075_),
    .Q_N(_2407_),
    .Q(\load_weights[46] ));
 sg13g2_dfrbp_1 _5089_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net40),
    .D(_0076_),
    .Q_N(_0010_),
    .Q(\load_weights[47] ));
 sg13g2_dfrbp_1 _5090_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net39),
    .D(_0077_),
    .Q_N(_2406_),
    .Q(\load_weights[48] ));
 sg13g2_dfrbp_1 _5091_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net38),
    .D(_0078_),
    .Q_N(_2405_),
    .Q(\load_weights[49] ));
 sg13g2_dfrbp_1 _5092_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net37),
    .D(net793),
    .Q_N(_2404_),
    .Q(\load_weights[50] ));
 sg13g2_dfrbp_1 _5093_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net36),
    .D(_0080_),
    .Q_N(_2403_),
    .Q(\load_weights[51] ));
 sg13g2_dfrbp_1 _5094_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net35),
    .D(net800),
    .Q_N(_2402_),
    .Q(\load_weights[52] ));
 sg13g2_dfrbp_1 _5095_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net34),
    .D(net409),
    .Q_N(_2401_),
    .Q(\load_weights[53] ));
 sg13g2_dfrbp_1 _5096_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net33),
    .D(net743),
    .Q_N(_2400_),
    .Q(\load_weights[54] ));
 sg13g2_dfrbp_1 _5097_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net32),
    .D(net563),
    .Q_N(_2399_),
    .Q(\load_weights[55] ));
 sg13g2_dfrbp_1 _5098_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net31),
    .D(_0085_),
    .Q_N(_2398_),
    .Q(\load_weights[56] ));
 sg13g2_dfrbp_1 _5099_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net30),
    .D(_0086_),
    .Q_N(_2397_),
    .Q(\load_weights[57] ));
 sg13g2_dfrbp_1 _5100_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net29),
    .D(net655),
    .Q_N(_2396_),
    .Q(\load_weights[58] ));
 sg13g2_dfrbp_1 _5101_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net28),
    .D(net819),
    .Q_N(_2395_),
    .Q(\load_weights[59] ));
 sg13g2_dfrbp_1 _5102_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net27),
    .D(net567),
    .Q_N(_2394_),
    .Q(\load_weights[60] ));
 sg13g2_dfrbp_1 _5103_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net26),
    .D(net772),
    .Q_N(_2393_),
    .Q(\load_weights[61] ));
 sg13g2_dfrbp_1 _5104_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net25),
    .D(_0091_),
    .Q_N(_2392_),
    .Q(\load_weights[62] ));
 sg13g2_dfrbp_1 _5105_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net24),
    .D(_0092_),
    .Q_N(_2391_),
    .Q(\load_weights[63] ));
 sg13g2_dfrbp_1 _5106_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net23),
    .D(_0093_),
    .Q_N(_2390_),
    .Q(\load_weights[64] ));
 sg13g2_dfrbp_1 _5107_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net22),
    .D(_0094_),
    .Q_N(_2389_),
    .Q(\load_weights[65] ));
 sg13g2_dfrbp_1 _5108_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net21),
    .D(_0095_),
    .Q_N(_2388_),
    .Q(\load_weights[66] ));
 sg13g2_dfrbp_1 _5109_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net20),
    .D(_0096_),
    .Q_N(_2387_),
    .Q(\load_weights[67] ));
 sg13g2_dfrbp_1 _5110_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net19),
    .D(net632),
    .Q_N(_2386_),
    .Q(\load_weights[68] ));
 sg13g2_dfrbp_1 _5111_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net18),
    .D(_0098_),
    .Q_N(_2385_),
    .Q(\load_weights[69] ));
 sg13g2_dfrbp_1 _5112_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net17),
    .D(_0099_),
    .Q_N(_2384_),
    .Q(\load_weights[70] ));
 sg13g2_dfrbp_1 _5113_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net16),
    .D(_0100_),
    .Q_N(_0020_),
    .Q(\load_weights[71] ));
 sg13g2_dfrbp_1 _5114_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net15),
    .D(net787),
    .Q_N(_2383_),
    .Q(\load_weights[72] ));
 sg13g2_dfrbp_1 _5115_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net14),
    .D(net734),
    .Q_N(_2382_),
    .Q(\load_weights[73] ));
 sg13g2_dfrbp_1 _5116_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net13),
    .D(_0103_),
    .Q_N(_2381_),
    .Q(\load_weights[74] ));
 sg13g2_dfrbp_1 _5117_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net12),
    .D(_0104_),
    .Q_N(_2380_),
    .Q(\load_weights[75] ));
 sg13g2_dfrbp_1 _5118_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net11),
    .D(_0105_),
    .Q_N(_2379_),
    .Q(\load_weights[76] ));
 sg13g2_dfrbp_1 _5119_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net10),
    .D(_0106_),
    .Q_N(_2378_),
    .Q(\load_weights[77] ));
 sg13g2_dfrbp_1 _5120_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net315),
    .D(_0107_),
    .Q_N(_2377_),
    .Q(\load_weights[78] ));
 sg13g2_dfrbp_1 _5121_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net314),
    .D(net675),
    .Q_N(_2376_),
    .Q(\load_weights[79] ));
 sg13g2_dfrbp_1 _5122_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net313),
    .D(net809),
    .Q_N(_2375_),
    .Q(\load_weights[80] ));
 sg13g2_dfrbp_1 _5123_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net312),
    .D(_0110_),
    .Q_N(_2374_),
    .Q(\load_weights[81] ));
 sg13g2_dfrbp_1 _5124_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net311),
    .D(_0111_),
    .Q_N(_2373_),
    .Q(\load_weights[82] ));
 sg13g2_dfrbp_1 _5125_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net310),
    .D(_0112_),
    .Q_N(_2372_),
    .Q(\load_weights[83] ));
 sg13g2_dfrbp_1 _5126_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net309),
    .D(_0113_),
    .Q_N(_2371_),
    .Q(\load_weights[84] ));
 sg13g2_dfrbp_1 _5127_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net308),
    .D(_0114_),
    .Q_N(_2370_),
    .Q(\load_weights[85] ));
 sg13g2_dfrbp_1 _5128_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net307),
    .D(net903),
    .Q_N(_2369_),
    .Q(\load_weights[86] ));
 sg13g2_dfrbp_1 _5129_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net306),
    .D(net593),
    .Q_N(_2368_),
    .Q(\load_weights[87] ));
 sg13g2_dfrbp_1 _5130_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net305),
    .D(_0117_),
    .Q_N(_2367_),
    .Q(\load_weights[88] ));
 sg13g2_dfrbp_1 _5131_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net304),
    .D(_0118_),
    .Q_N(_2366_),
    .Q(\load_weights[89] ));
 sg13g2_dfrbp_1 _5132_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net303),
    .D(_0119_),
    .Q_N(_2365_),
    .Q(\load_weights[90] ));
 sg13g2_dfrbp_1 _5133_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net302),
    .D(_0120_),
    .Q_N(_2364_),
    .Q(\load_weights[91] ));
 sg13g2_dfrbp_1 _5134_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net301),
    .D(_0121_),
    .Q_N(_2363_),
    .Q(\load_weights[92] ));
 sg13g2_dfrbp_1 _5135_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net300),
    .D(_0122_),
    .Q_N(_2362_),
    .Q(\load_weights[93] ));
 sg13g2_dfrbp_1 _5136_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net299),
    .D(_0123_),
    .Q_N(_2361_),
    .Q(\load_weights[94] ));
 sg13g2_dfrbp_1 _5137_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net298),
    .D(_0124_),
    .Q_N(_0004_),
    .Q(\load_weights[95] ));
 sg13g2_dfrbp_1 _5138_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net297),
    .D(net705),
    .Q_N(_2360_),
    .Q(\load_weights[96] ));
 sg13g2_dfrbp_1 _5139_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net296),
    .D(_0126_),
    .Q_N(_2359_),
    .Q(\load_weights[97] ));
 sg13g2_dfrbp_1 _5140_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net295),
    .D(net685),
    .Q_N(_2358_),
    .Q(\load_weights[98] ));
 sg13g2_dfrbp_1 _5141_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net294),
    .D(net607),
    .Q_N(_2357_),
    .Q(\load_weights[99] ));
 sg13g2_dfrbp_1 _5142_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net293),
    .D(net661),
    .Q_N(_2356_),
    .Q(\load_weights[100] ));
 sg13g2_dfrbp_1 _5143_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net292),
    .D(_0130_),
    .Q_N(_2355_),
    .Q(\load_weights[101] ));
 sg13g2_dfrbp_1 _5144_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net291),
    .D(_0131_),
    .Q_N(_2354_),
    .Q(\load_weights[102] ));
 sg13g2_dfrbp_1 _5145_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net290),
    .D(_0132_),
    .Q_N(_2353_),
    .Q(\load_weights[103] ));
 sg13g2_dfrbp_1 _5146_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net289),
    .D(net852),
    .Q_N(_2352_),
    .Q(\load_weights[104] ));
 sg13g2_dfrbp_1 _5147_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net288),
    .D(_0134_),
    .Q_N(_2351_),
    .Q(\load_weights[105] ));
 sg13g2_dfrbp_1 _5148_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net287),
    .D(_0135_),
    .Q_N(_2350_),
    .Q(\load_weights[106] ));
 sg13g2_dfrbp_1 _5149_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net286),
    .D(_0136_),
    .Q_N(_2349_),
    .Q(\load_weights[107] ));
 sg13g2_dfrbp_1 _5150_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net285),
    .D(_0137_),
    .Q_N(_2348_),
    .Q(\load_weights[108] ));
 sg13g2_dfrbp_1 _5151_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net284),
    .D(net678),
    .Q_N(_2347_),
    .Q(\load_weights[109] ));
 sg13g2_dfrbp_1 _5152_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net283),
    .D(_0139_),
    .Q_N(_2346_),
    .Q(\load_weights[110] ));
 sg13g2_dfrbp_1 _5153_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net282),
    .D(_0140_),
    .Q_N(_2345_),
    .Q(\load_weights[111] ));
 sg13g2_dfrbp_1 _5154_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net281),
    .D(_0141_),
    .Q_N(_2344_),
    .Q(\load_weights[112] ));
 sg13g2_dfrbp_1 _5155_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net280),
    .D(net389),
    .Q_N(_2343_),
    .Q(\load_weights[113] ));
 sg13g2_dfrbp_1 _5156_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net279),
    .D(_0143_),
    .Q_N(_2342_),
    .Q(\load_weights[114] ));
 sg13g2_dfrbp_1 _5157_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net278),
    .D(net383),
    .Q_N(_2341_),
    .Q(\load_weights[115] ));
 sg13g2_dfrbp_1 _5158_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net277),
    .D(_0145_),
    .Q_N(_2340_),
    .Q(\load_weights[116] ));
 sg13g2_dfrbp_1 _5159_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net276),
    .D(_0146_),
    .Q_N(_2339_),
    .Q(\load_weights[117] ));
 sg13g2_dfrbp_1 _5160_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net275),
    .D(_0147_),
    .Q_N(_2338_),
    .Q(\load_weights[118] ));
 sg13g2_dfrbp_1 _5161_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net274),
    .D(net755),
    .Q_N(_0007_),
    .Q(\load_weights[119] ));
 sg13g2_dfrbp_1 _5162_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net273),
    .D(_0149_),
    .Q_N(_2337_),
    .Q(\load_weights[120] ));
 sg13g2_dfrbp_1 _5163_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net272),
    .D(net591),
    .Q_N(_2336_),
    .Q(\load_weights[121] ));
 sg13g2_dfrbp_1 _5164_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net271),
    .D(net645),
    .Q_N(_2335_),
    .Q(\load_weights[122] ));
 sg13g2_dfrbp_1 _5165_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net270),
    .D(net395),
    .Q_N(_2334_),
    .Q(\load_weights[123] ));
 sg13g2_dfrbp_1 _5166_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net269),
    .D(_0153_),
    .Q_N(_2333_),
    .Q(\load_weights[124] ));
 sg13g2_dfrbp_1 _5167_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net268),
    .D(_0154_),
    .Q_N(_2332_),
    .Q(\load_weights[125] ));
 sg13g2_dfrbp_1 _5168_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net267),
    .D(net823),
    .Q_N(_2331_),
    .Q(\load_weights[126] ));
 sg13g2_dfrbp_1 _5169_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net266),
    .D(_0156_),
    .Q_N(_2330_),
    .Q(\load_weights[127] ));
 sg13g2_dfrbp_1 _5170_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net265),
    .D(net586),
    .Q_N(_2329_),
    .Q(\load_weights[128] ));
 sg13g2_dfrbp_1 _5171_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net264),
    .D(_0158_),
    .Q_N(_2328_),
    .Q(\load_weights[129] ));
 sg13g2_dfrbp_1 _5172_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net263),
    .D(_0159_),
    .Q_N(_2327_),
    .Q(\load_weights[130] ));
 sg13g2_dfrbp_1 _5173_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net262),
    .D(net758),
    .Q_N(_2326_),
    .Q(\load_weights[131] ));
 sg13g2_dfrbp_1 _5174_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net261),
    .D(_0161_),
    .Q_N(_2325_),
    .Q(\load_weights[132] ));
 sg13g2_dfrbp_1 _5175_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net260),
    .D(_0162_),
    .Q_N(_2324_),
    .Q(\load_weights[133] ));
 sg13g2_dfrbp_1 _5176_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net259),
    .D(_0163_),
    .Q_N(_2323_),
    .Q(\load_weights[134] ));
 sg13g2_dfrbp_1 _5177_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net258),
    .D(_0164_),
    .Q_N(_2322_),
    .Q(\load_weights[135] ));
 sg13g2_dfrbp_1 _5178_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net257),
    .D(_0165_),
    .Q_N(_2321_),
    .Q(\load_weights[136] ));
 sg13g2_dfrbp_1 _5179_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net256),
    .D(net393),
    .Q_N(_2320_),
    .Q(\load_weights[137] ));
 sg13g2_dfrbp_1 _5180_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net255),
    .D(_0167_),
    .Q_N(_2319_),
    .Q(\load_weights[138] ));
 sg13g2_dfrbp_1 _5181_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net254),
    .D(net419),
    .Q_N(_2318_),
    .Q(\load_weights[139] ));
 sg13g2_dfrbp_1 _5182_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net253),
    .D(_0169_),
    .Q_N(_2317_),
    .Q(\load_weights[140] ));
 sg13g2_dfrbp_1 _5183_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net252),
    .D(net399),
    .Q_N(_2316_),
    .Q(\load_weights[141] ));
 sg13g2_dfrbp_1 _5184_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net251),
    .D(net584),
    .Q_N(_2315_),
    .Q(\load_weights[142] ));
 sg13g2_dfrbp_1 _5185_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net250),
    .D(net826),
    .Q_N(_0013_),
    .Q(\load_weights[143] ));
 sg13g2_dfrbp_1 _5186_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net249),
    .D(_0173_),
    .Q_N(_2314_),
    .Q(\load_weights[144] ));
 sg13g2_dfrbp_1 _5187_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net248),
    .D(_0174_),
    .Q_N(_2313_),
    .Q(\load_weights[145] ));
 sg13g2_dfrbp_1 _5188_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net247),
    .D(net601),
    .Q_N(_2312_),
    .Q(\load_weights[146] ));
 sg13g2_dfrbp_1 _5189_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net246),
    .D(_0176_),
    .Q_N(_2311_),
    .Q(\load_weights[147] ));
 sg13g2_dfrbp_1 _5190_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net245),
    .D(_0177_),
    .Q_N(_2310_),
    .Q(\load_weights[148] ));
 sg13g2_dfrbp_1 _5191_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net244),
    .D(_0178_),
    .Q_N(_2309_),
    .Q(\load_weights[149] ));
 sg13g2_dfrbp_1 _5192_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net243),
    .D(net688),
    .Q_N(_2308_),
    .Q(\load_weights[150] ));
 sg13g2_dfrbp_1 _5193_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net242),
    .D(net634),
    .Q_N(_2307_),
    .Q(\load_weights[151] ));
 sg13g2_dfrbp_1 _5194_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net241),
    .D(_0181_),
    .Q_N(_2306_),
    .Q(\load_weights[152] ));
 sg13g2_dfrbp_1 _5195_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net240),
    .D(_0182_),
    .Q_N(_2305_),
    .Q(\load_weights[153] ));
 sg13g2_dfrbp_1 _5196_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net239),
    .D(_0183_),
    .Q_N(_2304_),
    .Q(\load_weights[154] ));
 sg13g2_dfrbp_1 _5197_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net238),
    .D(net613),
    .Q_N(_2303_),
    .Q(\load_weights[155] ));
 sg13g2_dfrbp_1 _5198_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net237),
    .D(net589),
    .Q_N(_2302_),
    .Q(\load_weights[156] ));
 sg13g2_dfrbp_1 _5199_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net236),
    .D(_0186_),
    .Q_N(_2301_),
    .Q(\load_weights[157] ));
 sg13g2_dfrbp_1 _5200_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net235),
    .D(_0187_),
    .Q_N(_2300_),
    .Q(\load_weights[158] ));
 sg13g2_dfrbp_1 _5201_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net234),
    .D(_0188_),
    .Q_N(_2299_),
    .Q(\load_weights[159] ));
 sg13g2_dfrbp_1 _5202_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net233),
    .D(net402),
    .Q_N(_2298_),
    .Q(\load_weights[160] ));
 sg13g2_dfrbp_1 _5203_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net232),
    .D(net721),
    .Q_N(_2297_),
    .Q(\load_weights[161] ));
 sg13g2_dfrbp_1 _5204_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net231),
    .D(_0191_),
    .Q_N(_2296_),
    .Q(\load_weights[162] ));
 sg13g2_dfrbp_1 _5205_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net230),
    .D(_0192_),
    .Q_N(_2295_),
    .Q(\load_weights[163] ));
 sg13g2_dfrbp_1 _5206_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net229),
    .D(_0193_),
    .Q_N(_2294_),
    .Q(\load_weights[164] ));
 sg13g2_dfrbp_1 _5207_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net228),
    .D(net692),
    .Q_N(_2293_),
    .Q(\load_weights[165] ));
 sg13g2_dfrbp_1 _5208_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net227),
    .D(net391),
    .Q_N(_2292_),
    .Q(\load_weights[166] ));
 sg13g2_dfrbp_1 _5209_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net226),
    .D(_0196_),
    .Q_N(_2291_),
    .Q(\load_weights[167] ));
 sg13g2_dfrbp_1 _5210_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net225),
    .D(net622),
    .Q_N(_2290_),
    .Q(\load_weights[168] ));
 sg13g2_dfrbp_1 _5211_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net224),
    .D(net629),
    .Q_N(_2289_),
    .Q(\load_weights[169] ));
 sg13g2_dfrbp_1 _5212_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net223),
    .D(_0199_),
    .Q_N(_2288_),
    .Q(\load_weights[170] ));
 sg13g2_dfrbp_1 _5213_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net222),
    .D(net669),
    .Q_N(_2287_),
    .Q(\load_weights[171] ));
 sg13g2_dfrbp_1 _5214_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net221),
    .D(_0201_),
    .Q_N(_2286_),
    .Q(\load_weights[172] ));
 sg13g2_dfrbp_1 _5215_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net220),
    .D(net650),
    .Q_N(_2285_),
    .Q(\load_weights[173] ));
 sg13g2_dfrbp_1 _5216_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net219),
    .D(_0203_),
    .Q_N(_2284_),
    .Q(\load_weights[174] ));
 sg13g2_dfrbp_1 _5217_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net218),
    .D(net595),
    .Q_N(_2283_),
    .Q(\load_weights[175] ));
 sg13g2_dfrbp_1 _5218_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net217),
    .D(net627),
    .Q_N(_2282_),
    .Q(\load_weights[176] ));
 sg13g2_dfrbp_1 _5219_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net216),
    .D(net577),
    .Q_N(_2281_),
    .Q(\load_weights[177] ));
 sg13g2_dfrbp_1 _5220_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net215),
    .D(_0207_),
    .Q_N(_2280_),
    .Q(\load_weights[178] ));
 sg13g2_dfrbp_1 _5221_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net214),
    .D(net696),
    .Q_N(_2279_),
    .Q(\load_weights[179] ));
 sg13g2_dfrbp_1 _5222_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net213),
    .D(_0209_),
    .Q_N(_2278_),
    .Q(\load_weights[180] ));
 sg13g2_dfrbp_1 _5223_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net212),
    .D(_0210_),
    .Q_N(_2277_),
    .Q(\load_weights[181] ));
 sg13g2_dfrbp_1 _5224_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net211),
    .D(_0211_),
    .Q_N(_2276_),
    .Q(\load_weights[182] ));
 sg13g2_dfrbp_1 _5225_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net210),
    .D(_0212_),
    .Q_N(_2275_),
    .Q(\load_weights[183] ));
 sg13g2_dfrbp_1 _5226_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net209),
    .D(net571),
    .Q_N(_2274_),
    .Q(\load_weights[184] ));
 sg13g2_dfrbp_1 _5227_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net208),
    .D(_0214_),
    .Q_N(_2273_),
    .Q(\load_weights[185] ));
 sg13g2_dfrbp_1 _5228_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net207),
    .D(net681),
    .Q_N(_2272_),
    .Q(\load_weights[186] ));
 sg13g2_dfrbp_1 _5229_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net206),
    .D(_0216_),
    .Q_N(_2271_),
    .Q(\load_weights[187] ));
 sg13g2_dfrbp_1 _5230_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net205),
    .D(_0217_),
    .Q_N(_2270_),
    .Q(\load_weights[188] ));
 sg13g2_dfrbp_1 _5231_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net204),
    .D(_0218_),
    .Q_N(_2269_),
    .Q(\load_weights[189] ));
 sg13g2_dfrbp_1 _5232_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net203),
    .D(net397),
    .Q_N(_2268_),
    .Q(\load_weights[190] ));
 sg13g2_dfrbp_1 _5233_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net202),
    .D(_0220_),
    .Q_N(_2267_),
    .Q(\load_weights[191] ));
 sg13g2_dfrbp_1 _5234_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net201),
    .D(_0221_),
    .Q_N(_2266_),
    .Q(\load_weights[192] ));
 sg13g2_dfrbp_1 _5235_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net200),
    .D(_0222_),
    .Q_N(_2265_),
    .Q(\load_weights[193] ));
 sg13g2_dfrbp_1 _5236_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net199),
    .D(net690),
    .Q_N(_2264_),
    .Q(\load_weights[194] ));
 sg13g2_dfrbp_1 _5237_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net198),
    .D(_0224_),
    .Q_N(_2263_),
    .Q(\load_weights[195] ));
 sg13g2_dfrbp_1 _5238_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net197),
    .D(_0225_),
    .Q_N(_2262_),
    .Q(\load_weights[196] ));
 sg13g2_dfrbp_1 _5239_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net196),
    .D(net749),
    .Q_N(_2261_),
    .Q(\load_weights[197] ));
 sg13g2_dfrbp_1 _5240_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net195),
    .D(net862),
    .Q_N(_2260_),
    .Q(\load_weights[198] ));
 sg13g2_dfrbp_1 _5241_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net194),
    .D(_0228_),
    .Q_N(_2259_),
    .Q(\load_weights[199] ));
 sg13g2_dfrbp_1 _5242_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net193),
    .D(_0229_),
    .Q_N(_2258_),
    .Q(\load_weights[200] ));
 sg13g2_dfrbp_1 _5243_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net192),
    .D(_0230_),
    .Q_N(_2257_),
    .Q(\load_weights[201] ));
 sg13g2_dfrbp_1 _5244_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net191),
    .D(net847),
    .Q_N(_2256_),
    .Q(\load_weights[202] ));
 sg13g2_dfrbp_1 _5245_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net190),
    .D(_0232_),
    .Q_N(_2255_),
    .Q(\load_weights[203] ));
 sg13g2_dfrbp_1 _5246_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net189),
    .D(net790),
    .Q_N(_2254_),
    .Q(\load_weights[204] ));
 sg13g2_dfrbp_1 _5247_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net188),
    .D(net715),
    .Q_N(_2253_),
    .Q(\load_weights[205] ));
 sg13g2_dfrbp_1 _5248_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net187),
    .D(_0235_),
    .Q_N(_2252_),
    .Q(\load_weights[206] ));
 sg13g2_dfrbp_1 _5249_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net186),
    .D(_0236_),
    .Q_N(_2251_),
    .Q(\load_weights[207] ));
 sg13g2_dfrbp_1 _5250_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net185),
    .D(_0237_),
    .Q_N(_2250_),
    .Q(\load_weights[208] ));
 sg13g2_dfrbp_1 _5251_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net184),
    .D(_0238_),
    .Q_N(_2249_),
    .Q(\load_weights[209] ));
 sg13g2_dfrbp_1 _5252_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net183),
    .D(_0239_),
    .Q_N(_2248_),
    .Q(\load_weights[210] ));
 sg13g2_dfrbp_1 _5253_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net182),
    .D(net836),
    .Q_N(_2247_),
    .Q(\load_weights[211] ));
 sg13g2_dfrbp_1 _5254_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net181),
    .D(_0241_),
    .Q_N(_2246_),
    .Q(\load_weights[212] ));
 sg13g2_dfrbp_1 _5255_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net180),
    .D(_0242_),
    .Q_N(_2245_),
    .Q(\load_weights[213] ));
 sg13g2_dfrbp_1 _5256_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net179),
    .D(_0243_),
    .Q_N(_2244_),
    .Q(\load_weights[214] ));
 sg13g2_dfrbp_1 _5257_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net178),
    .D(_0244_),
    .Q_N(_2243_),
    .Q(\load_weights[215] ));
 sg13g2_dfrbp_1 _5258_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net177),
    .D(net915),
    .Q_N(_2242_),
    .Q(\load_weights[216] ));
 sg13g2_dfrbp_1 _5259_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net176),
    .D(net859),
    .Q_N(_2241_),
    .Q(\load_weights[217] ));
 sg13g2_dfrbp_1 _5260_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net175),
    .D(_0247_),
    .Q_N(_2240_),
    .Q(\load_weights[218] ));
 sg13g2_dfrbp_1 _5261_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net174),
    .D(net775),
    .Q_N(_2239_),
    .Q(\load_weights[219] ));
 sg13g2_dfrbp_1 _5262_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net173),
    .D(_0249_),
    .Q_N(_2238_),
    .Q(\load_weights[220] ));
 sg13g2_dfrbp_1 _5263_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net172),
    .D(_0250_),
    .Q_N(_2237_),
    .Q(\load_weights[221] ));
 sg13g2_dfrbp_1 _5264_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net171),
    .D(net839),
    .Q_N(_2236_),
    .Q(\load_weights[222] ));
 sg13g2_dfrbp_1 _5265_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net170),
    .D(net725),
    .Q_N(_2235_),
    .Q(\load_weights[223] ));
 sg13g2_dfrbp_1 _5266_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net169),
    .D(_0253_),
    .Q_N(_2234_),
    .Q(\load_weights[224] ));
 sg13g2_dfrbp_1 _5267_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net168),
    .D(_0254_),
    .Q_N(_2233_),
    .Q(\load_weights[225] ));
 sg13g2_dfrbp_1 _5268_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net167),
    .D(_0255_),
    .Q_N(_2232_),
    .Q(\load_weights[226] ));
 sg13g2_dfrbp_1 _5269_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net166),
    .D(net764),
    .Q_N(_2231_),
    .Q(\load_weights[227] ));
 sg13g2_dfrbp_1 _5270_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net165),
    .D(net910),
    .Q_N(_2230_),
    .Q(\load_weights[228] ));
 sg13g2_dfrbp_1 _5271_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net164),
    .D(_0258_),
    .Q_N(_2229_),
    .Q(\load_weights[229] ));
 sg13g2_dfrbp_1 _5272_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net163),
    .D(net891),
    .Q_N(_2228_),
    .Q(\load_weights[230] ));
 sg13g2_dfrbp_1 _5273_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net162),
    .D(_0260_),
    .Q_N(_2227_),
    .Q(\load_weights[231] ));
 sg13g2_dfrbp_1 _5274_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net161),
    .D(net411),
    .Q_N(_2226_),
    .Q(\load_weights[232] ));
 sg13g2_dfrbp_1 _5275_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net160),
    .D(_0262_),
    .Q_N(_2225_),
    .Q(\load_weights[233] ));
 sg13g2_dfrbp_1 _5276_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net159),
    .D(_0263_),
    .Q_N(_2224_),
    .Q(\load_weights[234] ));
 sg13g2_dfrbp_1 _5277_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net158),
    .D(_0264_),
    .Q_N(_2223_),
    .Q(\load_weights[235] ));
 sg13g2_dfrbp_1 _5278_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net157),
    .D(_0265_),
    .Q_N(_2222_),
    .Q(\load_weights[236] ));
 sg13g2_dfrbp_1 _5279_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net156),
    .D(net770),
    .Q_N(_2221_),
    .Q(\load_weights[237] ));
 sg13g2_dfrbp_1 _5280_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net155),
    .D(net565),
    .Q_N(_2220_),
    .Q(\load_weights[238] ));
 sg13g2_dfrbp_1 _5281_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net154),
    .D(_0268_),
    .Q_N(_2219_),
    .Q(\load_weights[239] ));
 sg13g2_dfrbp_1 _5282_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net153),
    .D(net813),
    .Q_N(_2218_),
    .Q(\load_weights[240] ));
 sg13g2_dfrbp_1 _5283_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net152),
    .D(net603),
    .Q_N(_2217_),
    .Q(\load_weights[241] ));
 sg13g2_dfrbp_1 _5284_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net151),
    .D(net636),
    .Q_N(_2216_),
    .Q(\load_weights[242] ));
 sg13g2_dfrbp_1 _5285_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net150),
    .D(_0272_),
    .Q_N(_2215_),
    .Q(\load_weights[243] ));
 sg13g2_dfrbp_1 _5286_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net149),
    .D(_0273_),
    .Q_N(_2214_),
    .Q(\load_weights[244] ));
 sg13g2_dfrbp_1 _5287_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net148),
    .D(net731),
    .Q_N(_2213_),
    .Q(\load_weights[245] ));
 sg13g2_dfrbp_1 _5288_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net147),
    .D(net782),
    .Q_N(_2212_),
    .Q(\load_weights[246] ));
 sg13g2_dfrbp_1 _5289_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net146),
    .D(net671),
    .Q_N(_2211_),
    .Q(\load_weights[247] ));
 sg13g2_dfrbp_1 _5290_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net145),
    .D(net642),
    .Q_N(_2210_),
    .Q(\load_weights[248] ));
 sg13g2_dfrbp_1 _5291_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net144),
    .D(net597),
    .Q_N(_2209_),
    .Q(\load_weights[249] ));
 sg13g2_dfrbp_1 _5292_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net143),
    .D(_0279_),
    .Q_N(_2208_),
    .Q(\load_weights[250] ));
 sg13g2_dfrbp_1 _5293_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net142),
    .D(_0280_),
    .Q_N(_2207_),
    .Q(\load_weights[251] ));
 sg13g2_dfrbp_1 _5294_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net141),
    .D(_0281_),
    .Q_N(_2206_),
    .Q(\load_weights[252] ));
 sg13g2_dfrbp_1 _5295_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net140),
    .D(_0282_),
    .Q_N(_2205_),
    .Q(\load_weights[253] ));
 sg13g2_dfrbp_1 _5296_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net139),
    .D(_0283_),
    .Q_N(_2204_),
    .Q(\load_weights[254] ));
 sg13g2_dfrbp_1 _5297_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net138),
    .D(net599),
    .Q_N(_2203_),
    .Q(\load_weights[255] ));
 sg13g2_dfrbp_1 _5298_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net137),
    .D(net582),
    .Q_N(_2202_),
    .Q(\load_weights[256] ));
 sg13g2_dfrbp_1 _5299_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net136),
    .D(_0286_),
    .Q_N(_2201_),
    .Q(\load_weights[257] ));
 sg13g2_dfrbp_1 _5300_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net135),
    .D(_0287_),
    .Q_N(_2200_),
    .Q(\load_weights[258] ));
 sg13g2_dfrbp_1 _5301_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net134),
    .D(_0288_),
    .Q_N(_2199_),
    .Q(\load_weights[259] ));
 sg13g2_dfrbp_1 _5302_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net133),
    .D(_0289_),
    .Q_N(_2198_),
    .Q(\load_weights[260] ));
 sg13g2_dfrbp_1 _5303_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net132),
    .D(_0290_),
    .Q_N(_2197_),
    .Q(\load_weights[261] ));
 sg13g2_dfrbp_1 _5304_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net131),
    .D(net569),
    .Q_N(_2196_),
    .Q(\load_weights[262] ));
 sg13g2_dfrbp_1 _5305_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net130),
    .D(net738),
    .Q_N(_2195_),
    .Q(\load_weights[263] ));
 sg13g2_dfrbp_1 _5306_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net129),
    .D(net802),
    .Q_N(_2194_),
    .Q(\load_weights[264] ));
 sg13g2_dfrbp_1 _5307_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net128),
    .D(_0294_),
    .Q_N(_2193_),
    .Q(\load_weights[265] ));
 sg13g2_dfrbp_1 _5308_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net127),
    .D(_0295_),
    .Q_N(_2192_),
    .Q(\load_weights[266] ));
 sg13g2_dfrbp_1 _5309_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net126),
    .D(net881),
    .Q_N(_2191_),
    .Q(\load_weights[267] ));
 sg13g2_dfrbp_1 _5310_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net125),
    .D(net817),
    .Q_N(_2190_),
    .Q(\load_weights[268] ));
 sg13g2_dfrbp_1 _5311_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net124),
    .D(net624),
    .Q_N(_2189_),
    .Q(\load_weights[269] ));
 sg13g2_dfrbp_1 _5312_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net123),
    .D(_0299_),
    .Q_N(_2188_),
    .Q(\load_weights[270] ));
 sg13g2_dfrbp_1 _5313_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net122),
    .D(net658),
    .Q_N(_2187_),
    .Q(\load_weights[271] ));
 sg13g2_dfrbp_1 _5314_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net121),
    .D(_0301_),
    .Q_N(_2186_),
    .Q(\load_weights[272] ));
 sg13g2_dfrbp_1 _5315_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net120),
    .D(_0302_),
    .Q_N(_2185_),
    .Q(\load_weights[273] ));
 sg13g2_dfrbp_1 _5316_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net119),
    .D(_0303_),
    .Q_N(_2184_),
    .Q(\load_weights[274] ));
 sg13g2_dfrbp_1 _5317_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net118),
    .D(net777),
    .Q_N(_2183_),
    .Q(\load_weights[275] ));
 sg13g2_dfrbp_1 _5318_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net117),
    .D(_0305_),
    .Q_N(_2182_),
    .Q(\load_weights[276] ));
 sg13g2_dfrbp_1 _5319_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net116),
    .D(_0306_),
    .Q_N(_2181_),
    .Q(\load_weights[277] ));
 sg13g2_dfrbp_1 _5320_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net115),
    .D(_0307_),
    .Q_N(_2180_),
    .Q(\load_weights[278] ));
 sg13g2_dfrbp_1 _5321_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net114),
    .D(_0308_),
    .Q_N(_2179_),
    .Q(\load_weights[279] ));
 sg13g2_dfrbp_1 _5322_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net113),
    .D(_0309_),
    .Q_N(_2178_),
    .Q(\load_weights[280] ));
 sg13g2_dfrbp_1 _5323_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net112),
    .D(_0310_),
    .Q_N(_2177_),
    .Q(\load_weights[281] ));
 sg13g2_dfrbp_1 _5324_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net111),
    .D(net895),
    .Q_N(_2176_),
    .Q(\load_weights[282] ));
 sg13g2_dfrbp_1 _5325_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net110),
    .D(_0312_),
    .Q_N(_2175_),
    .Q(\load_weights[283] ));
 sg13g2_dfrbp_1 _5326_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net109),
    .D(_0313_),
    .Q_N(_2174_),
    .Q(\load_weights[284] ));
 sg13g2_dfrbp_1 _5327_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net108),
    .D(_0314_),
    .Q_N(_2173_),
    .Q(\load_weights[285] ));
 sg13g2_dfrbp_1 _5328_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net107),
    .D(net766),
    .Q_N(_2172_),
    .Q(\load_weights[286] ));
 sg13g2_dfrbp_1 _5329_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net106),
    .D(_0316_),
    .Q_N(_2171_),
    .Q(\load_weights[287] ));
 sg13g2_dfrbp_1 _5330_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net105),
    .D(net404),
    .Q_N(_2170_),
    .Q(\bit_select[0] ));
 sg13g2_dfrbp_1 _5331_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net104),
    .D(_0318_),
    .Q_N(_2169_),
    .Q(\bit_select[1] ));
 sg13g2_dfrbp_1 _5332_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net103),
    .D(_0319_),
    .Q_N(_2168_),
    .Q(\bit_select[2] ));
 sg13g2_dfrbp_1 _5333_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net102),
    .D(_0320_),
    .Q_N(_2167_),
    .Q(\bit_select[3] ));
 sg13g2_dfrbp_1 _5334_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net101),
    .D(_0321_),
    .Q_N(_2166_),
    .Q(\bit_select[4] ));
 sg13g2_dfrbp_1 _5335_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net100),
    .D(_0322_),
    .Q_N(_2165_),
    .Q(\bit_select[5] ));
 sg13g2_dfrbp_1 _5336_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net99),
    .D(_0323_),
    .Q_N(_2164_),
    .Q(\bit_select[6] ));
 sg13g2_dfrbp_1 _5337_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net98),
    .D(_0324_),
    .Q_N(_2163_),
    .Q(\bit_select[7] ));
 sg13g2_dfrbp_1 _5338_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net97),
    .D(_0325_),
    .Q_N(_2162_),
    .Q(mult_ena));
 sg13g2_dfrbp_1 _5339_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net95),
    .D(_0326_),
    .Q_N(_2161_),
    .Q(load_ena));
 sg13g2_dfrbp_1 _5340_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net94),
    .D(net865),
    .Q_N(_2160_),
    .Q(\count[0] ));
 sg13g2_dfrbp_1 _5341_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net93),
    .D(_0328_),
    .Q_N(_2159_),
    .Q(\count[1] ));
 sg13g2_dfrbp_1 _5342_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net92),
    .D(net833),
    .Q_N(_2158_),
    .Q(\count[2] ));
 sg13g2_dfrbp_1 _5343_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net91),
    .D(_0330_),
    .Q_N(_2157_),
    .Q(\count[3] ));
 sg13g2_dfrbp_1 _5344_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net90),
    .D(_0331_),
    .Q_N(_2156_),
    .Q(\count[4] ));
 sg13g2_dfrbp_1 _5345_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net89),
    .D(net873),
    .Q_N(_2155_),
    .Q(\count[5] ));
 sg13g2_dfrbp_1 _5346_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net88),
    .D(_0333_),
    .Q_N(_2154_),
    .Q(\count[6] ));
 sg13g2_dfrbp_1 _5347_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net317),
    .D(_0334_),
    .Q_N(_2454_),
    .Q(\count[7] ));
 sg13g2_dfrbp_1 _5348_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net318),
    .D(\tt_um_mult_inst.genblk1[0].out_q ),
    .Q_N(_2455_),
    .Q(\tt_um_mult_inst.genblk1[0].out ));
 sg13g2_dfrbp_1 _5349_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net319),
    .D(\tt_um_mult_inst.genblk1[0].carry_q[0] ),
    .Q_N(_0015_),
    .Q(\tt_um_mult_inst.genblk1[0].carry[0] ));
 sg13g2_dfrbp_1 _5350_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net320),
    .D(\tt_um_mult_inst.genblk1[0].carry_q[1] ),
    .Q_N(_2456_),
    .Q(\tt_um_mult_inst.genblk1[0].carry[1] ));
 sg13g2_dfrbp_1 _5351_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net321),
    .D(\tt_um_mult_inst.genblk1[0].carry_q[2] ),
    .Q_N(_2457_),
    .Q(\tt_um_mult_inst.genblk1[0].carry[2] ));
 sg13g2_dfrbp_1 _5352_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net322),
    .D(\tt_um_mult_inst.genblk1[0].carry_q[3] ),
    .Q_N(_0016_),
    .Q(\tt_um_mult_inst.genblk1[0].carry[3] ));
 sg13g2_dfrbp_1 _5353_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net323),
    .D(\tt_um_mult_inst.genblk1[1].out_q ),
    .Q_N(_2458_),
    .Q(\tt_um_mult_inst.genblk1[1].out ));
 sg13g2_dfrbp_1 _5354_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net324),
    .D(\tt_um_mult_inst.genblk1[1].carry_q[0] ),
    .Q_N(_0009_),
    .Q(\tt_um_mult_inst.genblk1[1].carry[0] ));
 sg13g2_dfrbp_1 _5355_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net325),
    .D(\tt_um_mult_inst.genblk1[1].carry_q[1] ),
    .Q_N(_2459_),
    .Q(\tt_um_mult_inst.genblk1[1].carry[1] ));
 sg13g2_dfrbp_1 _5356_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net326),
    .D(\tt_um_mult_inst.genblk1[1].carry_q[2] ),
    .Q_N(_2460_),
    .Q(\tt_um_mult_inst.genblk1[1].carry[2] ));
 sg13g2_dfrbp_1 _5357_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net327),
    .D(\tt_um_mult_inst.genblk1[1].carry_q[3] ),
    .Q_N(_0011_),
    .Q(\tt_um_mult_inst.genblk1[1].carry[3] ));
 sg13g2_dfrbp_1 _5358_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net328),
    .D(\tt_um_mult_inst.genblk1[2].out_q ),
    .Q_N(_2461_),
    .Q(\tt_um_mult_inst.genblk1[2].out ));
 sg13g2_dfrbp_1 _5359_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net329),
    .D(\tt_um_mult_inst.genblk1[2].carry_q[0] ),
    .Q_N(_0019_),
    .Q(\tt_um_mult_inst.genblk1[2].carry[0] ));
 sg13g2_dfrbp_1 _5360_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net330),
    .D(\tt_um_mult_inst.genblk1[2].carry_q[1] ),
    .Q_N(_2462_),
    .Q(\tt_um_mult_inst.genblk1[2].carry[1] ));
 sg13g2_dfrbp_1 _5361_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net331),
    .D(\tt_um_mult_inst.genblk1[2].carry_q[2] ),
    .Q_N(_2463_),
    .Q(\tt_um_mult_inst.genblk1[2].carry[2] ));
 sg13g2_dfrbp_1 _5362_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net332),
    .D(\tt_um_mult_inst.genblk1[2].carry_q[3] ),
    .Q_N(_0021_),
    .Q(\tt_um_mult_inst.genblk1[2].carry[3] ));
 sg13g2_dfrbp_1 _5363_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net333),
    .D(\tt_um_mult_inst.genblk1[3].out_q ),
    .Q_N(_2464_),
    .Q(\tt_um_mult_inst.genblk1[3].out ));
 sg13g2_dfrbp_1 _5364_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net334),
    .D(\tt_um_mult_inst.genblk1[3].carry_q[0] ),
    .Q_N(_0003_),
    .Q(\tt_um_mult_inst.genblk1[3].carry[0] ));
 sg13g2_dfrbp_1 _5365_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net335),
    .D(\tt_um_mult_inst.genblk1[3].carry_q[1] ),
    .Q_N(_2465_),
    .Q(\tt_um_mult_inst.genblk1[3].carry[1] ));
 sg13g2_dfrbp_1 _5366_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net336),
    .D(\tt_um_mult_inst.genblk1[3].carry_q[2] ),
    .Q_N(_2466_),
    .Q(\tt_um_mult_inst.genblk1[3].carry[2] ));
 sg13g2_dfrbp_1 _5367_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net337),
    .D(\tt_um_mult_inst.genblk1[3].carry_q[3] ),
    .Q_N(_0005_),
    .Q(\tt_um_mult_inst.genblk1[3].carry[3] ));
 sg13g2_dfrbp_1 _5368_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net338),
    .D(\tt_um_mult_inst.genblk1[4].out_q ),
    .Q_N(_2467_),
    .Q(\tt_um_mult_inst.genblk1[4].out ));
 sg13g2_dfrbp_1 _5369_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net339),
    .D(\tt_um_mult_inst.genblk1[4].carry_q[0] ),
    .Q_N(_0006_),
    .Q(\tt_um_mult_inst.genblk1[4].carry[0] ));
 sg13g2_dfrbp_1 _5370_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net340),
    .D(\tt_um_mult_inst.genblk1[4].carry_q[1] ),
    .Q_N(_2468_),
    .Q(\tt_um_mult_inst.genblk1[4].carry[1] ));
 sg13g2_dfrbp_1 _5371_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net341),
    .D(\tt_um_mult_inst.genblk1[4].carry_q[2] ),
    .Q_N(_2469_),
    .Q(\tt_um_mult_inst.genblk1[4].carry[2] ));
 sg13g2_dfrbp_1 _5372_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net342),
    .D(\tt_um_mult_inst.genblk1[4].carry_q[3] ),
    .Q_N(_0008_),
    .Q(\tt_um_mult_inst.genblk1[4].carry[3] ));
 sg13g2_dfrbp_1 _5373_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net343),
    .D(\tt_um_mult_inst.genblk1[5].out_q ),
    .Q_N(_2470_),
    .Q(\tt_um_mult_inst.genblk1[5].out ));
 sg13g2_dfrbp_1 _5374_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net344),
    .D(\tt_um_mult_inst.genblk1[5].carry_q[0] ),
    .Q_N(_0012_),
    .Q(\tt_um_mult_inst.genblk1[5].carry[0] ));
 sg13g2_dfrbp_1 _5375_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net345),
    .D(\tt_um_mult_inst.genblk1[5].carry_q[1] ),
    .Q_N(_2471_),
    .Q(\tt_um_mult_inst.genblk1[5].carry[1] ));
 sg13g2_dfrbp_1 _5376_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net346),
    .D(\tt_um_mult_inst.genblk1[5].carry_q[2] ),
    .Q_N(_2472_),
    .Q(\tt_um_mult_inst.genblk1[5].carry[2] ));
 sg13g2_dfrbp_1 _5377_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net347),
    .D(\tt_um_mult_inst.genblk1[5].carry_q[3] ),
    .Q_N(_0014_),
    .Q(\tt_um_mult_inst.genblk1[5].carry[3] ));
 sg13g2_dfrbp_1 _5378_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net348),
    .D(\tt_um_mult_inst.genblk1[6].out_q ),
    .Q_N(_2473_),
    .Q(\tt_um_mult_inst.genblk1[6].out ));
 sg13g2_dfrbp_1 _5379_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net349),
    .D(\tt_um_mult_inst.genblk1[6].carry_q[0] ),
    .Q_N(_0001_),
    .Q(\tt_um_mult_inst.genblk1[6].carry[0] ));
 sg13g2_dfrbp_1 _5380_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net350),
    .D(\tt_um_mult_inst.genblk1[6].carry_q[1] ),
    .Q_N(_2474_),
    .Q(\tt_um_mult_inst.genblk1[6].carry[1] ));
 sg13g2_dfrbp_1 _5381_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net351),
    .D(\tt_um_mult_inst.genblk1[6].carry_q[2] ),
    .Q_N(_2475_),
    .Q(\tt_um_mult_inst.genblk1[6].carry[2] ));
 sg13g2_dfrbp_1 _5382_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net352),
    .D(\tt_um_mult_inst.genblk1[6].carry_q[3] ),
    .Q_N(_0002_),
    .Q(\tt_um_mult_inst.genblk1[6].carry[3] ));
 sg13g2_dfrbp_1 _5383_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net353),
    .D(\tt_um_mult_inst.genblk1[7].out_q ),
    .Q_N(_2476_),
    .Q(\tt_um_mult_inst.genblk1[7].out ));
 sg13g2_dfrbp_1 _5384_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net354),
    .D(\tt_um_mult_inst.genblk1[7].carry_q[0] ),
    .Q_N(_0017_),
    .Q(\tt_um_mult_inst.genblk1[7].carry[0] ));
 sg13g2_dfrbp_1 _5385_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net355),
    .D(\tt_um_mult_inst.genblk1[7].carry_q[1] ),
    .Q_N(_2477_),
    .Q(\tt_um_mult_inst.genblk1[7].carry[1] ));
 sg13g2_dfrbp_1 _5386_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net356),
    .D(\tt_um_mult_inst.genblk1[7].carry_q[2] ),
    .Q_N(_2478_),
    .Q(\tt_um_mult_inst.genblk1[7].carry[2] ));
 sg13g2_dfrbp_1 _5387_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net357),
    .D(\tt_um_mult_inst.genblk1[7].carry_q[3] ),
    .Q_N(_0018_),
    .Q(\tt_um_mult_inst.genblk1[7].carry[3] ));
 sg13g2_dfrbp_1 _5388_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net358),
    .D(\tt_um_mult_inst.genblk1[8].out_q ),
    .Q_N(_2479_),
    .Q(\tt_um_mult_inst.genblk1[8].out ));
 sg13g2_dfrbp_1 _5389_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net359),
    .D(\tt_um_mult_inst.genblk1[8].carry_q[0] ),
    .Q_N(_0028_),
    .Q(\tt_um_mult_inst.genblk1[8].carry[0] ));
 sg13g2_dfrbp_1 _5390_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net360),
    .D(\tt_um_mult_inst.genblk1[8].carry_q[1] ),
    .Q_N(_2480_),
    .Q(\tt_um_mult_inst.genblk1[8].carry[1] ));
 sg13g2_dfrbp_1 _5391_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net361),
    .D(\tt_um_mult_inst.genblk1[8].carry_q[2] ),
    .Q_N(_2481_),
    .Q(\tt_um_mult_inst.genblk1[8].carry[2] ));
 sg13g2_dfrbp_1 _5392_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net362),
    .D(\tt_um_mult_inst.genblk1[8].carry_q[3] ),
    .Q_N(_0000_),
    .Q(\tt_um_mult_inst.genblk1[8].carry[3] ));
 sg13g2_dfrbp_1 _5393_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net363),
    .D(\tt_um_mult_inst.genblk1[9].out_q ),
    .Q_N(_2482_),
    .Q(\tt_um_mult_inst.genblk1[9].out ));
 sg13g2_dfrbp_1 _5394_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net364),
    .D(\tt_um_mult_inst.genblk1[9].carry_q[0] ),
    .Q_N(_0024_),
    .Q(\tt_um_mult_inst.genblk1[9].carry[0] ));
 sg13g2_dfrbp_1 _5395_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net365),
    .D(\tt_um_mult_inst.genblk1[9].carry_q[1] ),
    .Q_N(_2483_),
    .Q(\tt_um_mult_inst.genblk1[9].carry[1] ));
 sg13g2_dfrbp_1 _5396_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net366),
    .D(\tt_um_mult_inst.genblk1[9].carry_q[2] ),
    .Q_N(_2484_),
    .Q(\tt_um_mult_inst.genblk1[9].carry[2] ));
 sg13g2_dfrbp_1 _5397_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net367),
    .D(\tt_um_mult_inst.genblk1[9].carry_q[3] ),
    .Q_N(_0025_),
    .Q(\tt_um_mult_inst.genblk1[9].carry[3] ));
 sg13g2_dfrbp_1 _5398_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net368),
    .D(\tt_um_mult_inst.genblk1[10].out_q ),
    .Q_N(_2485_),
    .Q(\tt_um_mult_inst.genblk1[10].out ));
 sg13g2_dfrbp_1 _5399_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net369),
    .D(\tt_um_mult_inst.genblk1[10].carry_q[0] ),
    .Q_N(_0022_),
    .Q(\tt_um_mult_inst.genblk1[10].carry[0] ));
 sg13g2_dfrbp_1 _5400_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net370),
    .D(\tt_um_mult_inst.genblk1[10].carry_q[1] ),
    .Q_N(_2486_),
    .Q(\tt_um_mult_inst.genblk1[10].carry[1] ));
 sg13g2_dfrbp_1 _5401_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net371),
    .D(\tt_um_mult_inst.genblk1[10].carry_q[2] ),
    .Q_N(_2487_),
    .Q(\tt_um_mult_inst.genblk1[10].carry[2] ));
 sg13g2_dfrbp_1 _5402_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net372),
    .D(\tt_um_mult_inst.genblk1[10].carry_q[3] ),
    .Q_N(_0023_),
    .Q(\tt_um_mult_inst.genblk1[10].carry[3] ));
 sg13g2_dfrbp_1 _5403_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net373),
    .D(\tt_um_mult_inst.genblk1[11].out_q ),
    .Q_N(_2488_),
    .Q(\tt_um_mult_inst.genblk1[11].out ));
 sg13g2_dfrbp_1 _5404_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net374),
    .D(\tt_um_mult_inst.genblk1[11].carry_q[0] ),
    .Q_N(_0026_),
    .Q(\tt_um_mult_inst.genblk1[11].carry[0] ));
 sg13g2_dfrbp_1 _5405_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net375),
    .D(\tt_um_mult_inst.genblk1[11].carry_q[1] ),
    .Q_N(_2489_),
    .Q(\tt_um_mult_inst.genblk1[11].carry[1] ));
 sg13g2_dfrbp_1 _5406_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net96),
    .D(\tt_um_mult_inst.genblk1[11].carry_q[2] ),
    .Q_N(_2490_),
    .Q(\tt_um_mult_inst.genblk1[11].carry[2] ));
 sg13g2_dfrbp_1 _5407_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net87),
    .D(\tt_um_mult_inst.genblk1[11].carry_q[3] ),
    .Q_N(_0027_),
    .Q(\tt_um_mult_inst.genblk1[11].carry[3] ));
 sg13g2_tiehi _5118__11 (.L_HI(net11));
 sg13g2_tiehi _5117__12 (.L_HI(net12));
 sg13g2_tiehi _5116__13 (.L_HI(net13));
 sg13g2_tiehi _5115__14 (.L_HI(net14));
 sg13g2_tiehi _5114__15 (.L_HI(net15));
 sg13g2_tiehi _5113__16 (.L_HI(net16));
 sg13g2_tiehi _5112__17 (.L_HI(net17));
 sg13g2_tiehi _5111__18 (.L_HI(net18));
 sg13g2_tiehi _5110__19 (.L_HI(net19));
 sg13g2_tiehi _5109__20 (.L_HI(net20));
 sg13g2_tiehi _5108__21 (.L_HI(net21));
 sg13g2_tiehi _5107__22 (.L_HI(net22));
 sg13g2_tiehi _5106__23 (.L_HI(net23));
 sg13g2_tiehi _5105__24 (.L_HI(net24));
 sg13g2_tiehi _5104__25 (.L_HI(net25));
 sg13g2_tiehi _5103__26 (.L_HI(net26));
 sg13g2_tiehi _5102__27 (.L_HI(net27));
 sg13g2_tiehi _5101__28 (.L_HI(net28));
 sg13g2_tiehi _5100__29 (.L_HI(net29));
 sg13g2_tiehi _5099__30 (.L_HI(net30));
 sg13g2_tiehi _5098__31 (.L_HI(net31));
 sg13g2_tiehi _5097__32 (.L_HI(net32));
 sg13g2_tiehi _5096__33 (.L_HI(net33));
 sg13g2_tiehi _5095__34 (.L_HI(net34));
 sg13g2_tiehi _5094__35 (.L_HI(net35));
 sg13g2_tiehi _5093__36 (.L_HI(net36));
 sg13g2_tiehi _5092__37 (.L_HI(net37));
 sg13g2_tiehi _5091__38 (.L_HI(net38));
 sg13g2_tiehi _5090__39 (.L_HI(net39));
 sg13g2_tiehi _5089__40 (.L_HI(net40));
 sg13g2_tiehi _5088__41 (.L_HI(net41));
 sg13g2_tiehi _5087__42 (.L_HI(net42));
 sg13g2_tiehi _5086__43 (.L_HI(net43));
 sg13g2_tiehi _5085__44 (.L_HI(net44));
 sg13g2_tiehi _5084__45 (.L_HI(net45));
 sg13g2_tiehi _5083__46 (.L_HI(net46));
 sg13g2_tiehi _5082__47 (.L_HI(net47));
 sg13g2_tiehi _5081__48 (.L_HI(net48));
 sg13g2_tiehi _5080__49 (.L_HI(net49));
 sg13g2_tiehi _5079__50 (.L_HI(net50));
 sg13g2_tiehi _5078__51 (.L_HI(net51));
 sg13g2_tiehi _5077__52 (.L_HI(net52));
 sg13g2_tiehi _5076__53 (.L_HI(net53));
 sg13g2_tiehi _5075__54 (.L_HI(net54));
 sg13g2_tiehi _5074__55 (.L_HI(net55));
 sg13g2_tiehi _5073__56 (.L_HI(net56));
 sg13g2_tiehi _5072__57 (.L_HI(net57));
 sg13g2_tiehi _5071__58 (.L_HI(net58));
 sg13g2_tiehi _5070__59 (.L_HI(net59));
 sg13g2_tiehi _5069__60 (.L_HI(net60));
 sg13g2_tiehi _5068__61 (.L_HI(net61));
 sg13g2_tiehi _5067__62 (.L_HI(net62));
 sg13g2_tiehi _5066__63 (.L_HI(net63));
 sg13g2_tiehi _5065__64 (.L_HI(net64));
 sg13g2_tiehi _5064__65 (.L_HI(net65));
 sg13g2_tiehi _5063__66 (.L_HI(net66));
 sg13g2_tiehi _5062__67 (.L_HI(net67));
 sg13g2_tiehi _5061__68 (.L_HI(net68));
 sg13g2_tiehi _5060__69 (.L_HI(net69));
 sg13g2_tiehi _5059__70 (.L_HI(net70));
 sg13g2_tiehi _5058__71 (.L_HI(net71));
 sg13g2_tiehi _5057__72 (.L_HI(net72));
 sg13g2_tiehi _5056__73 (.L_HI(net73));
 sg13g2_tiehi _5055__74 (.L_HI(net74));
 sg13g2_tiehi _5054__75 (.L_HI(net75));
 sg13g2_tiehi _5053__76 (.L_HI(net76));
 sg13g2_tiehi _5052__77 (.L_HI(net77));
 sg13g2_tiehi _5051__78 (.L_HI(net78));
 sg13g2_tiehi _5050__79 (.L_HI(net79));
 sg13g2_tiehi _5049__80 (.L_HI(net80));
 sg13g2_tiehi _5048__81 (.L_HI(net81));
 sg13g2_tiehi _5047__82 (.L_HI(net82));
 sg13g2_tiehi _5046__83 (.L_HI(net83));
 sg13g2_tiehi _5045__84 (.L_HI(net84));
 sg13g2_tiehi _5044__85 (.L_HI(net85));
 sg13g2_tiehi _5043__86 (.L_HI(net86));
 sg13g2_tiehi _5407__87 (.L_HI(net87));
 sg13g2_tiehi _5346__88 (.L_HI(net88));
 sg13g2_tiehi _5345__89 (.L_HI(net89));
 sg13g2_tiehi _5344__90 (.L_HI(net90));
 sg13g2_tiehi _5343__91 (.L_HI(net91));
 sg13g2_tiehi _5342__92 (.L_HI(net92));
 sg13g2_tiehi _5341__93 (.L_HI(net93));
 sg13g2_tiehi _5340__94 (.L_HI(net94));
 sg13g2_tiehi _5339__95 (.L_HI(net95));
 sg13g2_tiehi _5406__96 (.L_HI(net96));
 sg13g2_tiehi _5338__97 (.L_HI(net97));
 sg13g2_tiehi _5337__98 (.L_HI(net98));
 sg13g2_tiehi _5336__99 (.L_HI(net99));
 sg13g2_tiehi _5335__100 (.L_HI(net100));
 sg13g2_tiehi _5334__101 (.L_HI(net101));
 sg13g2_tiehi _5333__102 (.L_HI(net102));
 sg13g2_tiehi _5332__103 (.L_HI(net103));
 sg13g2_tiehi _5331__104 (.L_HI(net104));
 sg13g2_tiehi _5330__105 (.L_HI(net105));
 sg13g2_tiehi _5329__106 (.L_HI(net106));
 sg13g2_tiehi _5328__107 (.L_HI(net107));
 sg13g2_tiehi _5327__108 (.L_HI(net108));
 sg13g2_tiehi _5326__109 (.L_HI(net109));
 sg13g2_tiehi _5325__110 (.L_HI(net110));
 sg13g2_tiehi _5324__111 (.L_HI(net111));
 sg13g2_tiehi _5323__112 (.L_HI(net112));
 sg13g2_tiehi _5322__113 (.L_HI(net113));
 sg13g2_tiehi _5321__114 (.L_HI(net114));
 sg13g2_tiehi _5320__115 (.L_HI(net115));
 sg13g2_tiehi _5319__116 (.L_HI(net116));
 sg13g2_tiehi _5318__117 (.L_HI(net117));
 sg13g2_tiehi _5317__118 (.L_HI(net118));
 sg13g2_tiehi _5316__119 (.L_HI(net119));
 sg13g2_tiehi _5315__120 (.L_HI(net120));
 sg13g2_tiehi _5314__121 (.L_HI(net121));
 sg13g2_tiehi _5313__122 (.L_HI(net122));
 sg13g2_tiehi _5312__123 (.L_HI(net123));
 sg13g2_tiehi _5311__124 (.L_HI(net124));
 sg13g2_tiehi _5310__125 (.L_HI(net125));
 sg13g2_tiehi _5309__126 (.L_HI(net126));
 sg13g2_tiehi _5308__127 (.L_HI(net127));
 sg13g2_tiehi _5307__128 (.L_HI(net128));
 sg13g2_tiehi _5306__129 (.L_HI(net129));
 sg13g2_tiehi _5305__130 (.L_HI(net130));
 sg13g2_tiehi _5304__131 (.L_HI(net131));
 sg13g2_tiehi _5303__132 (.L_HI(net132));
 sg13g2_tiehi _5302__133 (.L_HI(net133));
 sg13g2_tiehi _5301__134 (.L_HI(net134));
 sg13g2_tiehi _5300__135 (.L_HI(net135));
 sg13g2_tiehi _5299__136 (.L_HI(net136));
 sg13g2_tiehi _5298__137 (.L_HI(net137));
 sg13g2_tiehi _5297__138 (.L_HI(net138));
 sg13g2_tiehi _5296__139 (.L_HI(net139));
 sg13g2_tiehi _5295__140 (.L_HI(net140));
 sg13g2_tiehi _5294__141 (.L_HI(net141));
 sg13g2_tiehi _5293__142 (.L_HI(net142));
 sg13g2_tiehi _5292__143 (.L_HI(net143));
 sg13g2_tiehi _5291__144 (.L_HI(net144));
 sg13g2_tiehi _5290__145 (.L_HI(net145));
 sg13g2_tiehi _5289__146 (.L_HI(net146));
 sg13g2_tiehi _5288__147 (.L_HI(net147));
 sg13g2_tiehi _5287__148 (.L_HI(net148));
 sg13g2_tiehi _5286__149 (.L_HI(net149));
 sg13g2_tiehi _5285__150 (.L_HI(net150));
 sg13g2_tiehi _5284__151 (.L_HI(net151));
 sg13g2_tiehi _5283__152 (.L_HI(net152));
 sg13g2_tiehi _5282__153 (.L_HI(net153));
 sg13g2_tiehi _5281__154 (.L_HI(net154));
 sg13g2_tiehi _5280__155 (.L_HI(net155));
 sg13g2_tiehi _5279__156 (.L_HI(net156));
 sg13g2_tiehi _5278__157 (.L_HI(net157));
 sg13g2_tiehi _5277__158 (.L_HI(net158));
 sg13g2_tiehi _5276__159 (.L_HI(net159));
 sg13g2_tiehi _5275__160 (.L_HI(net160));
 sg13g2_tiehi _5274__161 (.L_HI(net161));
 sg13g2_tiehi _5273__162 (.L_HI(net162));
 sg13g2_tiehi _5272__163 (.L_HI(net163));
 sg13g2_tiehi _5271__164 (.L_HI(net164));
 sg13g2_tiehi _5270__165 (.L_HI(net165));
 sg13g2_tiehi _5269__166 (.L_HI(net166));
 sg13g2_tiehi _5268__167 (.L_HI(net167));
 sg13g2_tiehi _5267__168 (.L_HI(net168));
 sg13g2_tiehi _5266__169 (.L_HI(net169));
 sg13g2_tiehi _5265__170 (.L_HI(net170));
 sg13g2_tiehi _5264__171 (.L_HI(net171));
 sg13g2_tiehi _5263__172 (.L_HI(net172));
 sg13g2_tiehi _5262__173 (.L_HI(net173));
 sg13g2_tiehi _5261__174 (.L_HI(net174));
 sg13g2_tiehi _5260__175 (.L_HI(net175));
 sg13g2_tiehi _5259__176 (.L_HI(net176));
 sg13g2_tiehi _5258__177 (.L_HI(net177));
 sg13g2_tiehi _5257__178 (.L_HI(net178));
 sg13g2_tiehi _5256__179 (.L_HI(net179));
 sg13g2_tiehi _5255__180 (.L_HI(net180));
 sg13g2_tiehi _5254__181 (.L_HI(net181));
 sg13g2_tiehi _5253__182 (.L_HI(net182));
 sg13g2_tiehi _5252__183 (.L_HI(net183));
 sg13g2_tiehi _5251__184 (.L_HI(net184));
 sg13g2_tiehi _5250__185 (.L_HI(net185));
 sg13g2_tiehi _5249__186 (.L_HI(net186));
 sg13g2_tiehi _5248__187 (.L_HI(net187));
 sg13g2_tiehi _5247__188 (.L_HI(net188));
 sg13g2_tiehi _5246__189 (.L_HI(net189));
 sg13g2_tiehi _5245__190 (.L_HI(net190));
 sg13g2_tiehi _5244__191 (.L_HI(net191));
 sg13g2_tiehi _5243__192 (.L_HI(net192));
 sg13g2_tiehi _5242__193 (.L_HI(net193));
 sg13g2_tiehi _5241__194 (.L_HI(net194));
 sg13g2_tiehi _5240__195 (.L_HI(net195));
 sg13g2_tiehi _5239__196 (.L_HI(net196));
 sg13g2_tiehi _5238__197 (.L_HI(net197));
 sg13g2_tiehi _5237__198 (.L_HI(net198));
 sg13g2_tiehi _5236__199 (.L_HI(net199));
 sg13g2_tiehi _5235__200 (.L_HI(net200));
 sg13g2_tiehi _5234__201 (.L_HI(net201));
 sg13g2_tiehi _5233__202 (.L_HI(net202));
 sg13g2_tiehi _5232__203 (.L_HI(net203));
 sg13g2_tiehi _5231__204 (.L_HI(net204));
 sg13g2_tiehi _5230__205 (.L_HI(net205));
 sg13g2_tiehi _5229__206 (.L_HI(net206));
 sg13g2_tiehi _5228__207 (.L_HI(net207));
 sg13g2_tiehi _5227__208 (.L_HI(net208));
 sg13g2_tiehi _5226__209 (.L_HI(net209));
 sg13g2_tiehi _5225__210 (.L_HI(net210));
 sg13g2_tiehi _5224__211 (.L_HI(net211));
 sg13g2_tiehi _5223__212 (.L_HI(net212));
 sg13g2_tiehi _5222__213 (.L_HI(net213));
 sg13g2_tiehi _5221__214 (.L_HI(net214));
 sg13g2_tiehi _5220__215 (.L_HI(net215));
 sg13g2_tiehi _5219__216 (.L_HI(net216));
 sg13g2_tiehi _5218__217 (.L_HI(net217));
 sg13g2_tiehi _5217__218 (.L_HI(net218));
 sg13g2_tiehi _5216__219 (.L_HI(net219));
 sg13g2_tiehi _5215__220 (.L_HI(net220));
 sg13g2_tiehi _5214__221 (.L_HI(net221));
 sg13g2_tiehi _5213__222 (.L_HI(net222));
 sg13g2_tiehi _5212__223 (.L_HI(net223));
 sg13g2_tiehi _5211__224 (.L_HI(net224));
 sg13g2_tiehi _5210__225 (.L_HI(net225));
 sg13g2_tiehi _5209__226 (.L_HI(net226));
 sg13g2_tiehi _5208__227 (.L_HI(net227));
 sg13g2_tiehi _5207__228 (.L_HI(net228));
 sg13g2_tiehi _5206__229 (.L_HI(net229));
 sg13g2_tiehi _5205__230 (.L_HI(net230));
 sg13g2_tiehi _5204__231 (.L_HI(net231));
 sg13g2_tiehi _5203__232 (.L_HI(net232));
 sg13g2_tiehi _5202__233 (.L_HI(net233));
 sg13g2_tiehi _5201__234 (.L_HI(net234));
 sg13g2_tiehi _5200__235 (.L_HI(net235));
 sg13g2_tiehi _5199__236 (.L_HI(net236));
 sg13g2_tiehi _5198__237 (.L_HI(net237));
 sg13g2_tiehi _5197__238 (.L_HI(net238));
 sg13g2_tiehi _5196__239 (.L_HI(net239));
 sg13g2_tiehi _5195__240 (.L_HI(net240));
 sg13g2_tiehi _5194__241 (.L_HI(net241));
 sg13g2_tiehi _5193__242 (.L_HI(net242));
 sg13g2_tiehi _5192__243 (.L_HI(net243));
 sg13g2_tiehi _5191__244 (.L_HI(net244));
 sg13g2_tiehi _5190__245 (.L_HI(net245));
 sg13g2_tiehi _5189__246 (.L_HI(net246));
 sg13g2_tiehi _5188__247 (.L_HI(net247));
 sg13g2_tiehi _5187__248 (.L_HI(net248));
 sg13g2_tiehi _5186__249 (.L_HI(net249));
 sg13g2_tiehi _5185__250 (.L_HI(net250));
 sg13g2_tiehi _5184__251 (.L_HI(net251));
 sg13g2_tiehi _5183__252 (.L_HI(net252));
 sg13g2_tiehi _5182__253 (.L_HI(net253));
 sg13g2_tiehi _5181__254 (.L_HI(net254));
 sg13g2_tiehi _5180__255 (.L_HI(net255));
 sg13g2_tiehi _5179__256 (.L_HI(net256));
 sg13g2_tiehi _5178__257 (.L_HI(net257));
 sg13g2_tiehi _5177__258 (.L_HI(net258));
 sg13g2_tiehi _5176__259 (.L_HI(net259));
 sg13g2_tiehi _5175__260 (.L_HI(net260));
 sg13g2_tiehi _5174__261 (.L_HI(net261));
 sg13g2_tiehi _5173__262 (.L_HI(net262));
 sg13g2_tiehi _5172__263 (.L_HI(net263));
 sg13g2_tiehi _5171__264 (.L_HI(net264));
 sg13g2_tiehi _5170__265 (.L_HI(net265));
 sg13g2_tiehi _5169__266 (.L_HI(net266));
 sg13g2_tiehi _5168__267 (.L_HI(net267));
 sg13g2_tiehi _5167__268 (.L_HI(net268));
 sg13g2_tiehi _5166__269 (.L_HI(net269));
 sg13g2_tiehi _5165__270 (.L_HI(net270));
 sg13g2_tiehi _5164__271 (.L_HI(net271));
 sg13g2_tiehi _5163__272 (.L_HI(net272));
 sg13g2_tiehi _5162__273 (.L_HI(net273));
 sg13g2_tiehi _5161__274 (.L_HI(net274));
 sg13g2_tiehi _5160__275 (.L_HI(net275));
 sg13g2_tiehi _5159__276 (.L_HI(net276));
 sg13g2_tiehi _5158__277 (.L_HI(net277));
 sg13g2_tiehi _5157__278 (.L_HI(net278));
 sg13g2_tiehi _5156__279 (.L_HI(net279));
 sg13g2_tiehi _5155__280 (.L_HI(net280));
 sg13g2_tiehi _5154__281 (.L_HI(net281));
 sg13g2_tiehi _5153__282 (.L_HI(net282));
 sg13g2_tiehi _5152__283 (.L_HI(net283));
 sg13g2_tiehi _5151__284 (.L_HI(net284));
 sg13g2_tiehi _5150__285 (.L_HI(net285));
 sg13g2_tiehi _5149__286 (.L_HI(net286));
 sg13g2_tiehi _5148__287 (.L_HI(net287));
 sg13g2_tiehi _5147__288 (.L_HI(net288));
 sg13g2_tiehi _5146__289 (.L_HI(net289));
 sg13g2_tiehi _5145__290 (.L_HI(net290));
 sg13g2_tiehi _5144__291 (.L_HI(net291));
 sg13g2_tiehi _5143__292 (.L_HI(net292));
 sg13g2_tiehi _5142__293 (.L_HI(net293));
 sg13g2_tiehi _5141__294 (.L_HI(net294));
 sg13g2_tiehi _5140__295 (.L_HI(net295));
 sg13g2_tiehi _5139__296 (.L_HI(net296));
 sg13g2_tiehi _5138__297 (.L_HI(net297));
 sg13g2_tiehi _5137__298 (.L_HI(net298));
 sg13g2_tiehi _5136__299 (.L_HI(net299));
 sg13g2_tiehi _5135__300 (.L_HI(net300));
 sg13g2_tiehi _5134__301 (.L_HI(net301));
 sg13g2_tiehi _5133__302 (.L_HI(net302));
 sg13g2_tiehi _5132__303 (.L_HI(net303));
 sg13g2_tiehi _5131__304 (.L_HI(net304));
 sg13g2_tiehi _5130__305 (.L_HI(net305));
 sg13g2_tiehi _5129__306 (.L_HI(net306));
 sg13g2_tiehi _5128__307 (.L_HI(net307));
 sg13g2_tiehi _5127__308 (.L_HI(net308));
 sg13g2_tiehi _5126__309 (.L_HI(net309));
 sg13g2_tiehi _5125__310 (.L_HI(net310));
 sg13g2_tiehi _5124__311 (.L_HI(net311));
 sg13g2_tiehi _5123__312 (.L_HI(net312));
 sg13g2_tiehi _5122__313 (.L_HI(net313));
 sg13g2_tiehi _5121__314 (.L_HI(net314));
 sg13g2_tiehi _5120__315 (.L_HI(net315));
 sg13g2_tiehi _5042__316 (.L_HI(net316));
 sg13g2_tiehi _5347__317 (.L_HI(net317));
 sg13g2_tiehi _5348__318 (.L_HI(net318));
 sg13g2_tiehi _5349__319 (.L_HI(net319));
 sg13g2_tiehi _5350__320 (.L_HI(net320));
 sg13g2_tiehi _5351__321 (.L_HI(net321));
 sg13g2_tiehi _5352__322 (.L_HI(net322));
 sg13g2_tiehi _5353__323 (.L_HI(net323));
 sg13g2_tiehi _5354__324 (.L_HI(net324));
 sg13g2_tiehi _5355__325 (.L_HI(net325));
 sg13g2_tiehi _5356__326 (.L_HI(net326));
 sg13g2_tiehi _5357__327 (.L_HI(net327));
 sg13g2_tiehi _5358__328 (.L_HI(net328));
 sg13g2_tiehi _5359__329 (.L_HI(net329));
 sg13g2_tiehi _5360__330 (.L_HI(net330));
 sg13g2_tiehi _5361__331 (.L_HI(net331));
 sg13g2_tiehi _5362__332 (.L_HI(net332));
 sg13g2_tiehi _5363__333 (.L_HI(net333));
 sg13g2_tiehi _5364__334 (.L_HI(net334));
 sg13g2_tiehi _5365__335 (.L_HI(net335));
 sg13g2_tiehi _5366__336 (.L_HI(net336));
 sg13g2_tiehi _5367__337 (.L_HI(net337));
 sg13g2_tiehi _5368__338 (.L_HI(net338));
 sg13g2_tiehi _5369__339 (.L_HI(net339));
 sg13g2_tiehi _5370__340 (.L_HI(net340));
 sg13g2_tiehi _5371__341 (.L_HI(net341));
 sg13g2_tiehi _5372__342 (.L_HI(net342));
 sg13g2_tiehi _5373__343 (.L_HI(net343));
 sg13g2_tiehi _5374__344 (.L_HI(net344));
 sg13g2_tiehi _5375__345 (.L_HI(net345));
 sg13g2_tiehi _5376__346 (.L_HI(net346));
 sg13g2_tiehi _5377__347 (.L_HI(net347));
 sg13g2_tiehi _5378__348 (.L_HI(net348));
 sg13g2_tiehi _5379__349 (.L_HI(net349));
 sg13g2_tiehi _5380__350 (.L_HI(net350));
 sg13g2_tiehi _5381__351 (.L_HI(net351));
 sg13g2_tiehi _5382__352 (.L_HI(net352));
 sg13g2_tiehi _5383__353 (.L_HI(net353));
 sg13g2_tiehi _5384__354 (.L_HI(net354));
 sg13g2_tiehi _5385__355 (.L_HI(net355));
 sg13g2_tiehi _5386__356 (.L_HI(net356));
 sg13g2_tiehi _5387__357 (.L_HI(net357));
 sg13g2_tiehi _5388__358 (.L_HI(net358));
 sg13g2_tiehi _5389__359 (.L_HI(net359));
 sg13g2_tiehi _5390__360 (.L_HI(net360));
 sg13g2_tiehi _5391__361 (.L_HI(net361));
 sg13g2_tiehi _5392__362 (.L_HI(net362));
 sg13g2_tiehi _5393__363 (.L_HI(net363));
 sg13g2_tiehi _5394__364 (.L_HI(net364));
 sg13g2_tiehi _5395__365 (.L_HI(net365));
 sg13g2_tiehi _5396__366 (.L_HI(net366));
 sg13g2_tiehi _5397__367 (.L_HI(net367));
 sg13g2_tiehi _5398__368 (.L_HI(net368));
 sg13g2_tiehi _5399__369 (.L_HI(net369));
 sg13g2_tiehi _5400__370 (.L_HI(net370));
 sg13g2_tiehi _5401__371 (.L_HI(net371));
 sg13g2_tiehi _5402__372 (.L_HI(net372));
 sg13g2_tiehi _5403__373 (.L_HI(net373));
 sg13g2_tiehi _5404__374 (.L_HI(net374));
 sg13g2_tiehi _5405__375 (.L_HI(net375));
 sg13g2_tiehi tt_um_tiny_ternary_tapeout_csa_376 (.L_HI(net376));
 sg13g2_tiehi tt_um_tiny_ternary_tapeout_csa_377 (.L_HI(net377));
 sg13g2_tiehi tt_um_tiny_ternary_tapeout_csa_378 (.L_HI(net378));
 sg13g2_tiehi tt_um_tiny_ternary_tapeout_csa_379 (.L_HI(net379));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_csa_3 (.L_LO(net3));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_csa_4 (.L_LO(net4));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_csa_5 (.L_LO(net5));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_csa_6 (.L_LO(net6));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_csa_7 (.L_LO(net7));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_csa_8 (.L_LO(net8));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_csa_9 (.L_LO(net9));
 sg13g2_tiehi _5119__10 (.L_HI(net10));
 sg13g2_buf_1 _5786_ (.A(\tt_um_mult_inst.genblk1[0].out ),
    .X(uio_out[0]));
 sg13g2_buf_1 _5787_ (.A(\tt_um_mult_inst.genblk1[1].out ),
    .X(uio_out[1]));
 sg13g2_buf_2 _5788_ (.A(\tt_um_mult_inst.genblk1[2].out ),
    .X(uio_out[2]));
 sg13g2_buf_4 _5789_ (.X(uio_out[3]),
    .A(\tt_um_mult_inst.genblk1[3].out ));
 sg13g2_buf_4 _5790_ (.X(uo_out[0]),
    .A(\tt_um_mult_inst.genblk1[4].out ));
 sg13g2_buf_2 _5791_ (.A(\tt_um_mult_inst.genblk1[5].out ),
    .X(uo_out[1]));
 sg13g2_buf_1 _5792_ (.A(\tt_um_mult_inst.genblk1[6].out ),
    .X(uo_out[2]));
 sg13g2_buf_1 _5793_ (.A(\tt_um_mult_inst.genblk1[7].out ),
    .X(uo_out[3]));
 sg13g2_buf_2 _5794_ (.A(\tt_um_mult_inst.genblk1[8].out ),
    .X(uo_out[4]));
 sg13g2_buf_1 _5795_ (.A(\tt_um_mult_inst.genblk1[9].out ),
    .X(uo_out[5]));
 sg13g2_buf_2 _5796_ (.A(\tt_um_mult_inst.genblk1[10].out ),
    .X(uo_out[6]));
 sg13g2_buf_1 _5797_ (.A(\tt_um_mult_inst.genblk1[11].out ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(_1887_));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(net427));
 sg13g2_buf_2 fanout423 (.A(net427),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(net426),
    .X(net424));
 sg13g2_buf_1 fanout425 (.A(net426),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(net427),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_1992_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(net431),
    .X(net428));
 sg13g2_buf_4 fanout429 (.X(net429),
    .A(net431));
 sg13g2_buf_2 fanout430 (.A(net431),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_1992_),
    .X(net431));
 sg13g2_buf_4 fanout432 (.X(net432),
    .A(net433));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(_1992_));
 sg13g2_buf_4 fanout434 (.X(net434),
    .A(net436));
 sg13g2_buf_4 fanout435 (.X(net435),
    .A(net436));
 sg13g2_buf_2 fanout436 (.A(net438),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(net438),
    .X(net437));
 sg13g2_buf_4 fanout438 (.X(net438),
    .A(_1991_));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(net442));
 sg13g2_buf_2 fanout440 (.A(net442),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(net442),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_1991_),
    .X(net442));
 sg13g2_buf_4 fanout443 (.X(net443),
    .A(net445));
 sg13g2_buf_2 fanout444 (.A(net445),
    .X(net444));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(net450));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(net448));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(net450),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(net475),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(net454),
    .X(net451));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(net454));
 sg13g2_buf_2 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(net475),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(net457),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(net457),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(net458),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(net475),
    .X(net458));
 sg13g2_buf_4 fanout459 (.X(net459),
    .A(net460));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(net462));
 sg13g2_buf_4 fanout461 (.X(net461),
    .A(net462));
 sg13g2_buf_2 fanout462 (.A(net466),
    .X(net462));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(net465));
 sg13g2_buf_1 fanout464 (.A(net465),
    .X(net464));
 sg13g2_buf_1 fanout465 (.A(net466),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(net475),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(net471),
    .X(net467));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(net471));
 sg13g2_buf_4 fanout469 (.X(net469),
    .A(net471));
 sg13g2_buf_2 fanout470 (.A(net471),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(net475),
    .X(net471));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(net474));
 sg13g2_buf_2 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_4 fanout475 (.X(net475),
    .A(load_ena));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(net477));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(net481));
 sg13g2_buf_2 fanout478 (.A(net479),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(net481));
 sg13g2_buf_2 fanout481 (.A(net489),
    .X(net481));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(net486));
 sg13g2_buf_2 fanout483 (.A(net486),
    .X(net483));
 sg13g2_buf_4 fanout484 (.X(net484),
    .A(net486));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(net489),
    .X(net486));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(net489));
 sg13g2_buf_2 fanout488 (.A(net489),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(net504),
    .X(net489));
 sg13g2_buf_4 fanout490 (.X(net490),
    .A(net493));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net493));
 sg13g2_buf_2 fanout492 (.A(net493),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(net504),
    .X(net493));
 sg13g2_buf_4 fanout494 (.X(net494),
    .A(net498));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(net498));
 sg13g2_buf_4 fanout496 (.X(net496),
    .A(net497));
 sg13g2_buf_2 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(net504),
    .X(net498));
 sg13g2_buf_4 fanout499 (.X(net499),
    .A(net503));
 sg13g2_buf_2 fanout500 (.A(net503),
    .X(net500));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(net502));
 sg13g2_buf_2 fanout502 (.A(net503),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(net504),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(load_ena),
    .X(net504));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(net508));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(net508));
 sg13g2_buf_1 fanout507 (.A(net508),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net510),
    .X(net508));
 sg13g2_buf_4 fanout509 (.X(net509),
    .A(net510));
 sg13g2_buf_2 fanout510 (.A(uio_in[7]),
    .X(net510));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(net515));
 sg13g2_buf_4 fanout512 (.X(net512),
    .A(net515));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(net515));
 sg13g2_buf_2 fanout514 (.A(net515),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(uio_in[6]),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(net517),
    .X(net516));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(net520));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(net520));
 sg13g2_buf_2 fanout519 (.A(net520),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(uio_in[5]),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(uio_in[4]),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(uio_in[4]),
    .X(net522));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(net525));
 sg13g2_buf_2 fanout524 (.A(net525),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(uio_in[4]),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(net529));
 sg13g2_buf_4 fanout527 (.X(net527),
    .A(net529));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(net529));
 sg13g2_buf_8 fanout529 (.A(ui_in[7]),
    .X(net529));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(net534));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(net534));
 sg13g2_buf_2 fanout532 (.A(net534),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(ui_in[6]),
    .X(net534));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(net536));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net538));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(net538));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(ui_in[5]));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(net543));
 sg13g2_buf_2 fanout540 (.A(net543),
    .X(net540));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(net542));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(net543));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(ui_in[4]));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(net545));
 sg13g2_buf_4 fanout545 (.X(net545),
    .A(ui_in[3]));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(ui_in[3]));
 sg13g2_buf_2 fanout547 (.A(ui_in[3]),
    .X(net547));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(net549));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(net552));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(net552));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(ui_in[2]),
    .X(net552));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(net554));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(net557));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(net557));
 sg13g2_buf_2 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(ui_in[1]),
    .X(net557));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(net562));
 sg13g2_buf_4 fanout559 (.X(net559),
    .A(net562));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(net562));
 sg13g2_buf_2 fanout561 (.A(net562),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(ui_in[0]),
    .X(net562));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_tiny_ternary_tapeout_csa_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_46_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_49_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_50_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_45_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_37_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_38_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_39_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_40_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_42_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_20_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_36_clk));
 sg13g2_inv_8 clkload17 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_11_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_16_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_17_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_28_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_22_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\load_weights[4] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0045_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold3 (.A(\load_weights[103] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0144_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold5 (.A(\load_weights[29] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0070_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold7 (.A(\load_weights[27] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0068_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold9 (.A(\load_weights[101] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0142_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold11 (.A(\load_weights[154] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0195_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold13 (.A(\load_weights[125] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0166_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold15 (.A(\load_weights[123] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0152_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold17 (.A(\load_weights[178] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0219_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold19 (.A(\load_weights[129] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0170_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold21 (.A(\load_weights[117] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold22 (.A(\load_weights[148] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0189_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold24 (.A(\bit_select[0] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0317_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold26 (.A(\load_weights[10] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0051_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold28 (.A(\load_weights[135] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold29 (.A(\load_weights[53] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0082_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold31 (.A(\load_weights[220] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0261_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold33 (.A(\load_weights[166] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold34 (.A(\load_weights[105] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold35 (.A(\load_weights[93] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold36 (.A(\load_weights[81] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold37 (.A(\load_weights[31] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0072_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold39 (.A(\load_weights[127] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0168_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold41 (.A(\load_weights[55] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0084_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold43 (.A(\load_weights[226] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0267_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold45 (.A(\load_weights[48] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0089_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold47 (.A(\load_weights[250] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0291_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold49 (.A(\load_weights[172] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0213_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold51 (.A(\load_weights[7] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0048_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold53 (.A(\load_weights[115] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold54 (.A(\bit_select[1] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold55 (.A(\load_weights[177] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0206_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold57 (.A(\load_weights[113] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold58 (.A(\load_weights[34] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0063_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold60 (.A(\load_weights[244] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0285_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold62 (.A(\load_weights[130] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0171_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold64 (.A(\load_weights[128] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0157_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold66 (.A(\load_weights[118] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold67 (.A(\load_weights[144] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0185_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold69 (.A(\load_weights[121] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0150_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold71 (.A(\load_weights[75] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0116_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold73 (.A(\load_weights[175] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0204_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold75 (.A(\load_weights[249] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0278_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold77 (.A(\load_weights[243] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0284_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold79 (.A(\load_weights[146] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0175_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold81 (.A(\load_weights[241] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0270_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold83 (.A(\load_weights[17] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold84 (.A(\load_weights[147] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold85 (.A(\load_weights[99] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0128_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold87 (.A(\load_weights[19] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold88 (.A(\load_weights[232] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold89 (.A(\load_weights[187] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold90 (.A(\load_weights[158] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold91 (.A(\load_weights[155] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0184_),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold93 (.A(\load_weights[133] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold94 (.A(\load_weights[8] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0049_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold96 (.A(\load_weights[140] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold97 (.A(\load_weights[145] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold98 (.A(\load_weights[32] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0061_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold100 (.A(\load_weights[168] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0197_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold102 (.A(\load_weights[269] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0298_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold104 (.A(\load_weights[231] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold105 (.A(\load_weights[176] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0205_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold107 (.A(\load_weights[169] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0198_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold109 (.A(\load_weights[89] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold110 (.A(\load_weights[56] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0097_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold112 (.A(\load_weights[151] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0180_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold114 (.A(\load_weights[242] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0271_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold116 (.A(\load_weights[214] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold117 (.A(\load_weights[11] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold118 (.A(\load_weights[91] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold119 (.A(\load_weights[44] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold120 (.A(\load_weights[248] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0277_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold122 (.A(\load_weights[180] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold123 (.A(\load_weights[122] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0151_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold125 (.A(\load_weights[6] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold126 (.A(\load_weights[28] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0057_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold128 (.A(\load_weights[173] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0202_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold130 (.A(\load_weights[18] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold131 (.A(\load_weights[63] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold132 (.A(\load_weights[3] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold133 (.A(\load_weights[58] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0087_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold135 (.A(\load_weights[5] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold136 (.A(\load_weights[271] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0300_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold138 (.A(\load_weights[2] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold139 (.A(\load_weights[100] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0129_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold141 (.A(\load_weights[0] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0041_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold143 (.A(\load_weights[136] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold144 (.A(\load_weights[111] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold145 (.A(\load_weights[1] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold146 (.A(\bit_select[7] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold147 (.A(\load_weights[171] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0200_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold149 (.A(\load_weights[247] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0276_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold151 (.A(\load_weights[157] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold152 (.A(\load_weights[253] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold153 (.A(\load_weights[79] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0108_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold155 (.A(\load_weights[23] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold156 (.A(\load_weights[97] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0138_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold158 (.A(\load_weights[281] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold159 (.A(\load_weights[174] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0215_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold161 (.A(\load_weights[25] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0054_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold163 (.A(\load_weights[98] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0127_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold165 (.A(\load_weights[238] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold166 (.A(\load_weights[150] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0179_),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold168 (.A(\load_weights[194] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0223_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold170 (.A(\load_weights[153] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0194_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold172 (.A(\load_weights[283] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold173 (.A(\load_weights[261] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold174 (.A(\load_weights[179] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0208_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold176 (.A(\load_weights[189] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold177 (.A(\load_weights[15] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold178 (.A(\load_weights[260] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold179 (.A(\load_weights[36] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold180 (.A(\load_weights[170] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold181 (.A(\load_weights[37] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold182 (.A(\load_weights[132] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold183 (.A(\load_weights[96] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0125_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold185 (.A(\bit_select[2] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold186 (.A(\load_weights[30] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold187 (.A(\load_weights[108] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold188 (.A(\load_weights[69] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold189 (.A(\load_weights[163] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold190 (.A(\load_weights[33] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0074_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold192 (.A(\load_weights[142] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold193 (.A(\load_weights[193] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0234_),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold195 (.A(\load_weights[85] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold196 (.A(\load_weights[112] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold197 (.A(\load_weights[124] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold198 (.A(\load_weights[57] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold199 (.A(\load_weights[149] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0190_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold201 (.A(\load_weights[208] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold202 (.A(\load_weights[167] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold203 (.A(\load_weights[223] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0252_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold205 (.A(\load_weights[259] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold206 (.A(\load_weights[110] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold207 (.A(\load_weights[137] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold208 (.A(\load_weights[162] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold209 (.A(\load_weights[245] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0274_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold211 (.A(\load_weights[188] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold212 (.A(\load_weights[73] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0102_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold214 (.A(\load_weights[141] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold215 (.A(\load_weights[134] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold216 (.A(\load_weights[251] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0292_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold218 (.A(\load_weights[181] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold219 (.A(\load_weights[273] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold220 (.A(\load_weights[254] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold221 (.A(\load_weights[54] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0083_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold223 (.A(\load_weights[191] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold224 (.A(\load_weights[66] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold225 (.A(\load_weights[120] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold226 (.A(\load_weights[24] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold227 (.A(\load_weights[197] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0226_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold229 (.A(\load_weights[51] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold230 (.A(\load_weights[285] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold231 (.A(\load_weights[257] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold232 (.A(\load_weights[77] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold233 (.A(\load_weights[107] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0148_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold235 (.A(\load_weights[13] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold236 (.A(\load_weights[119] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0160_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold238 (.A(\load_weights[183] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold239 (.A(\bit_select[6] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold240 (.A(\load_weights[21] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold241 (.A(\load_weights[235] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold242 (.A(\load_weights[227] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0256_),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold244 (.A(\load_weights[274] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0315_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold246 (.A(\load_weights[182] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold247 (.A(\load_weights[160] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold248 (.A(\load_weights[225] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0266_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold250 (.A(\load_weights[49] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0090_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold252 (.A(\load_weights[14] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold253 (.A(\load_weights[219] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0248_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold255 (.A(\load_weights[275] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0304_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold257 (.A(\load_weights[95] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold258 (.A(\load_weights[152] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold259 (.A(\load_weights[9] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold260 (.A(\load_weights[246] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0275_),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold262 (.A(\load_weights[70] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold263 (.A(\load_weights[206] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold264 (.A(\load_weights[164] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold265 (.A(\load_weights[72] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0101_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold267 (.A(\load_weights[239] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold268 (.A(\load_weights[192] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0233_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold270 (.A(\load_weights[35] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold271 (.A(\load_weights[50] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0079_),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold273 (.A(\load_weights[258] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold274 (.A(\load_weights[287] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold275 (.A(\load_weights[65] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold276 (.A(\load_weights[201] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold277 (.A(\load_weights[12] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold278 (.A(\load_weights[52] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0081_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold280 (.A(\load_weights[264] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0293_),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold282 (.A(\load_weights[185] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold283 (.A(\load_weights[42] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold284 (.A(\load_weights[195] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold285 (.A(\load_weights[64] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold286 (.A(\bit_select[3] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold287 (.A(\load_weights[80] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0109_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold289 (.A(\load_weights[78] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold290 (.A(\load_weights[200] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold291 (.A(\load_weights[240] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0269_),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold293 (.A(\load_weights[252] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold294 (.A(\load_weights[209] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold295 (.A(\load_weights[268] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0297_),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold297 (.A(\load_weights[47] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0088_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold299 (.A(\load_weights[213] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold300 (.A(\load_weights[265] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold301 (.A(\load_weights[126] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0155_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold303 (.A(\load_weights[84] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold304 (.A(\load_weights[131] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0172_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold306 (.A(\load_weights[62] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold307 (.A(\load_weights[67] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold308 (.A(\load_weights[212] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold309 (.A(\load_weights[196] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold310 (.A(\count[2] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold311 (.A(_1911_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0329_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold313 (.A(\load_weights[46] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold314 (.A(\load_weights[199] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0240_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold316 (.A(\load_weights[82] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold317 (.A(\load_weights[222] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0251_),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold319 (.A(\load_weights[276] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold320 (.A(\load_weights[83] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold321 (.A(\load_weights[207] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold322 (.A(\bit_select[4] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold323 (.A(\load_weights[94] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold324 (.A(\load_weights[277] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold325 (.A(\load_weights[202] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0231_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold327 (.A(\load_weights[203] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold328 (.A(\load_weights[138] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold329 (.A(\load_weights[71] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold330 (.A(\load_weights[104] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0133_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold332 (.A(\load_weights[159] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold333 (.A(\load_weights[106] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold334 (.A(\load_weights[215] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold335 (.A(\bit_select[5] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold336 (.A(\load_weights[184] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold337 (.A(\load_weights[217] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0246_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold339 (.A(\load_weights[92] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold340 (.A(\load_weights[198] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0227_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold342 (.A(\load_weights[210] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold343 (.A(\count[0] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0327_),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold345 (.A(\load_weights[280] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold346 (.A(\load_weights[59] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold347 (.A(\load_weights[40] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold348 (.A(\load_weights[90] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold349 (.A(\load_weights[39] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold350 (.A(\count[5] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold351 (.A(_1918_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0332_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold353 (.A(\load_weights[272] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold354 (.A(\load_weights[262] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold355 (.A(\load_weights[116] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold356 (.A(\count[4] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold357 (.A(_1916_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold358 (.A(\load_weights[234] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold359 (.A(\load_weights[267] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0296_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold361 (.A(\load_weights[221] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold362 (.A(\count[3] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold363 (.A(_1914_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold364 (.A(\load_weights[45] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold365 (.A(\load_weights[26] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold366 (.A(\load_weights[38] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold367 (.A(\load_weights[224] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold368 (.A(\load_weights[284] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold369 (.A(\load_weights[218] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0259_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold371 (.A(mult_ena),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold372 (.A(_1893_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold373 (.A(\load_weights[270] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0311_),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold375 (.A(\load_weights[102] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold376 (.A(\load_weights[279] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold377 (.A(\load_weights[114] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold378 (.A(\load_weights[229] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold379 (.A(\load_weights[266] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold380 (.A(\load_weights[278] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold381 (.A(\load_weights[74] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0115_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold383 (.A(\count[6] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold384 (.A(\load_weights[236] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold385 (.A(\load_weights[233] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0002_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold387 (.A(\count[1] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold388 (.A(\load_weights[228] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0257_),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold390 (.A(\load_weights[76] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold391 (.A(\count[7] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold392 (.A(\load_weights[88] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold393 (.A(\load_weights[216] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0245_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0000_),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold396 (.A(\count[4] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0021_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold398 (.A(_1821_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0025_),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0016_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0027_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0581_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0005_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0018_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0014_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0023_),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0008_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold408 (.A(\load_weights[45] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0011_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold410 (.A(\load_weights[67] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold411 (.A(\load_weights[213] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold412 (.A(\load_weights[99] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold413 (.A(_1080_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold414 (.A(\load_weights[79] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold415 (.A(\load_weights[123] ),
    .X(net936));
 sg13g2_antennanp ANTENNA_1 (.A(\tt_um_mult_inst.genblk1[6].out_q ));
 sg13g2_antennanp ANTENNA_2 (.A(ui_in[0]));
 sg13g2_antennanp ANTENNA_3 (.A(ui_in[4]));
 sg13g2_antennanp ANTENNA_4 (.A(uio_in[6]));
 sg13g2_antennanp ANTENNA_5 (.A(ui_in[4]));
 sg13g2_antennanp ANTENNA_6 (.A(uio_in[6]));
 sg13g2_antennanp ANTENNA_7 (.A(ui_in[4]));
 sg13g2_antennanp ANTENNA_8 (.A(uio_in[6]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_4 FILLER_0_63 ();
 sg13g2_fill_2 FILLER_0_67 ();
 sg13g2_decap_8 FILLER_0_107 ();
 sg13g2_decap_8 FILLER_0_114 ();
 sg13g2_fill_2 FILLER_0_121 ();
 sg13g2_fill_1 FILLER_0_123 ();
 sg13g2_fill_2 FILLER_0_128 ();
 sg13g2_fill_1 FILLER_0_130 ();
 sg13g2_fill_2 FILLER_0_148 ();
 sg13g2_fill_1 FILLER_0_150 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_fill_1 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_177 ();
 sg13g2_fill_1 FILLER_0_184 ();
 sg13g2_decap_4 FILLER_0_194 ();
 sg13g2_fill_2 FILLER_0_226 ();
 sg13g2_fill_1 FILLER_0_228 ();
 sg13g2_fill_1 FILLER_0_233 ();
 sg13g2_decap_4 FILLER_0_238 ();
 sg13g2_fill_1 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_fill_2 FILLER_0_261 ();
 sg13g2_fill_1 FILLER_0_263 ();
 sg13g2_fill_2 FILLER_0_310 ();
 sg13g2_decap_4 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_4 FILLER_1_49 ();
 sg13g2_fill_2 FILLER_1_117 ();
 sg13g2_fill_2 FILLER_1_160 ();
 sg13g2_fill_1 FILLER_1_162 ();
 sg13g2_fill_2 FILLER_1_238 ();
 sg13g2_fill_1 FILLER_1_240 ();
 sg13g2_fill_1 FILLER_1_293 ();
 sg13g2_fill_2 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_fill_2 FILLER_2_75 ();
 sg13g2_fill_1 FILLER_2_77 ();
 sg13g2_fill_2 FILLER_2_82 ();
 sg13g2_fill_2 FILLER_2_88 ();
 sg13g2_fill_2 FILLER_2_186 ();
 sg13g2_fill_2 FILLER_2_214 ();
 sg13g2_fill_1 FILLER_2_242 ();
 sg13g2_fill_1 FILLER_2_257 ();
 sg13g2_fill_2 FILLER_2_273 ();
 sg13g2_fill_1 FILLER_2_337 ();
 sg13g2_fill_2 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_fill_2 FILLER_3_176 ();
 sg13g2_fill_1 FILLER_3_178 ();
 sg13g2_decap_8 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_386 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_fill_1 FILLER_4_28 ();
 sg13g2_fill_2 FILLER_4_115 ();
 sg13g2_fill_1 FILLER_4_164 ();
 sg13g2_fill_2 FILLER_4_199 ();
 sg13g2_fill_1 FILLER_4_233 ();
 sg13g2_fill_1 FILLER_4_260 ();
 sg13g2_fill_1 FILLER_4_274 ();
 sg13g2_fill_2 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_4 FILLER_5_21 ();
 sg13g2_fill_2 FILLER_5_25 ();
 sg13g2_fill_2 FILLER_5_53 ();
 sg13g2_fill_1 FILLER_5_55 ();
 sg13g2_fill_1 FILLER_5_68 ();
 sg13g2_fill_2 FILLER_5_87 ();
 sg13g2_fill_1 FILLER_5_125 ();
 sg13g2_fill_1 FILLER_5_135 ();
 sg13g2_fill_1 FILLER_5_145 ();
 sg13g2_fill_1 FILLER_5_238 ();
 sg13g2_fill_1 FILLER_5_267 ();
 sg13g2_fill_2 FILLER_5_348 ();
 sg13g2_fill_1 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_68 ();
 sg13g2_fill_2 FILLER_6_151 ();
 sg13g2_fill_1 FILLER_6_184 ();
 sg13g2_decap_4 FILLER_6_236 ();
 sg13g2_fill_1 FILLER_6_240 ();
 sg13g2_fill_1 FILLER_6_246 ();
 sg13g2_fill_1 FILLER_6_304 ();
 sg13g2_fill_2 FILLER_6_331 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_4 FILLER_7_14 ();
 sg13g2_fill_2 FILLER_7_18 ();
 sg13g2_fill_2 FILLER_7_42 ();
 sg13g2_fill_1 FILLER_7_44 ();
 sg13g2_fill_2 FILLER_7_54 ();
 sg13g2_fill_2 FILLER_7_66 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_fill_1 FILLER_7_90 ();
 sg13g2_fill_2 FILLER_7_183 ();
 sg13g2_fill_2 FILLER_7_229 ();
 sg13g2_fill_1 FILLER_7_231 ();
 sg13g2_fill_2 FILLER_7_251 ();
 sg13g2_fill_1 FILLER_7_253 ();
 sg13g2_fill_2 FILLER_7_279 ();
 sg13g2_fill_2 FILLER_7_299 ();
 sg13g2_fill_1 FILLER_7_301 ();
 sg13g2_fill_2 FILLER_7_313 ();
 sg13g2_fill_1 FILLER_7_315 ();
 sg13g2_fill_1 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_fill_2 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_30 ();
 sg13g2_fill_2 FILLER_8_90 ();
 sg13g2_fill_1 FILLER_8_92 ();
 sg13g2_fill_2 FILLER_8_115 ();
 sg13g2_fill_1 FILLER_8_132 ();
 sg13g2_fill_2 FILLER_8_164 ();
 sg13g2_fill_1 FILLER_8_166 ();
 sg13g2_fill_1 FILLER_8_176 ();
 sg13g2_fill_2 FILLER_8_202 ();
 sg13g2_fill_1 FILLER_8_204 ();
 sg13g2_fill_1 FILLER_8_244 ();
 sg13g2_fill_2 FILLER_8_255 ();
 sg13g2_fill_1 FILLER_8_270 ();
 sg13g2_fill_2 FILLER_8_283 ();
 sg13g2_fill_1 FILLER_8_285 ();
 sg13g2_fill_2 FILLER_8_305 ();
 sg13g2_fill_2 FILLER_8_320 ();
 sg13g2_fill_1 FILLER_8_341 ();
 sg13g2_fill_2 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_46 ();
 sg13g2_fill_1 FILLER_9_94 ();
 sg13g2_fill_2 FILLER_9_116 ();
 sg13g2_fill_1 FILLER_9_118 ();
 sg13g2_fill_2 FILLER_9_127 ();
 sg13g2_fill_1 FILLER_9_129 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_142 ();
 sg13g2_fill_1 FILLER_9_190 ();
 sg13g2_fill_2 FILLER_9_242 ();
 sg13g2_decap_8 FILLER_9_276 ();
 sg13g2_fill_1 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_292 ();
 sg13g2_fill_1 FILLER_9_355 ();
 sg13g2_fill_1 FILLER_9_368 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_63 ();
 sg13g2_fill_2 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_132 ();
 sg13g2_fill_2 FILLER_10_148 ();
 sg13g2_fill_2 FILLER_10_176 ();
 sg13g2_fill_2 FILLER_10_224 ();
 sg13g2_fill_1 FILLER_10_250 ();
 sg13g2_decap_8 FILLER_10_267 ();
 sg13g2_decap_4 FILLER_10_274 ();
 sg13g2_fill_2 FILLER_10_278 ();
 sg13g2_fill_2 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_327 ();
 sg13g2_fill_1 FILLER_10_329 ();
 sg13g2_decap_4 FILLER_10_356 ();
 sg13g2_fill_2 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_4 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_fill_2 FILLER_11_36 ();
 sg13g2_fill_1 FILLER_11_38 ();
 sg13g2_fill_2 FILLER_11_48 ();
 sg13g2_fill_2 FILLER_11_70 ();
 sg13g2_fill_2 FILLER_11_87 ();
 sg13g2_fill_1 FILLER_11_89 ();
 sg13g2_fill_2 FILLER_11_106 ();
 sg13g2_fill_1 FILLER_11_108 ();
 sg13g2_fill_1 FILLER_11_117 ();
 sg13g2_fill_2 FILLER_11_200 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_fill_2 FILLER_11_207 ();
 sg13g2_fill_1 FILLER_11_218 ();
 sg13g2_fill_1 FILLER_11_231 ();
 sg13g2_fill_2 FILLER_11_281 ();
 sg13g2_decap_4 FILLER_11_295 ();
 sg13g2_fill_1 FILLER_11_299 ();
 sg13g2_fill_2 FILLER_11_329 ();
 sg13g2_fill_1 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_fill_1 FILLER_12_18 ();
 sg13g2_decap_4 FILLER_12_29 ();
 sg13g2_fill_2 FILLER_12_67 ();
 sg13g2_fill_2 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_79 ();
 sg13g2_fill_2 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_113 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_fill_2 FILLER_12_184 ();
 sg13g2_fill_2 FILLER_12_199 ();
 sg13g2_fill_1 FILLER_12_201 ();
 sg13g2_fill_2 FILLER_12_215 ();
 sg13g2_fill_2 FILLER_12_226 ();
 sg13g2_fill_1 FILLER_12_228 ();
 sg13g2_fill_1 FILLER_12_241 ();
 sg13g2_fill_1 FILLER_12_255 ();
 sg13g2_fill_2 FILLER_12_299 ();
 sg13g2_fill_1 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_323 ();
 sg13g2_fill_2 FILLER_12_345 ();
 sg13g2_fill_1 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_fill_2 FILLER_12_359 ();
 sg13g2_fill_1 FILLER_12_361 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_16 ();
 sg13g2_fill_2 FILLER_13_43 ();
 sg13g2_fill_2 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_fill_2 FILLER_13_305 ();
 sg13g2_fill_1 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_fill_2 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_358 ();
 sg13g2_decap_4 FILLER_13_364 ();
 sg13g2_fill_2 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_18 ();
 sg13g2_fill_2 FILLER_14_23 ();
 sg13g2_fill_1 FILLER_14_60 ();
 sg13g2_fill_2 FILLER_14_92 ();
 sg13g2_fill_1 FILLER_14_94 ();
 sg13g2_fill_2 FILLER_14_169 ();
 sg13g2_fill_1 FILLER_14_171 ();
 sg13g2_fill_2 FILLER_14_203 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_276 ();
 sg13g2_fill_2 FILLER_14_301 ();
 sg13g2_fill_2 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_fill_1 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_34 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_164 ();
 sg13g2_decap_4 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_207 ();
 sg13g2_fill_2 FILLER_15_253 ();
 sg13g2_fill_1 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_fill_1 FILLER_15_341 ();
 sg13g2_decap_4 FILLER_15_392 ();
 sg13g2_decap_4 FILLER_16_26 ();
 sg13g2_fill_2 FILLER_16_114 ();
 sg13g2_fill_1 FILLER_16_116 ();
 sg13g2_fill_2 FILLER_16_143 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_fill_2 FILLER_16_192 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_fill_2 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_219 ();
 sg13g2_decap_4 FILLER_16_224 ();
 sg13g2_decap_4 FILLER_16_260 ();
 sg13g2_fill_2 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_fill_1 FILLER_16_277 ();
 sg13g2_fill_2 FILLER_16_335 ();
 sg13g2_decap_4 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_346 ();
 sg13g2_decap_4 FILLER_16_362 ();
 sg13g2_fill_1 FILLER_16_391 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_25 ();
 sg13g2_fill_2 FILLER_17_51 ();
 sg13g2_decap_4 FILLER_17_78 ();
 sg13g2_fill_1 FILLER_17_103 ();
 sg13g2_fill_2 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_172 ();
 sg13g2_fill_2 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_263 ();
 sg13g2_fill_2 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_fill_1 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_decap_4 FILLER_17_348 ();
 sg13g2_fill_1 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_4 FILLER_17_387 ();
 sg13g2_fill_2 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_16 ();
 sg13g2_decap_8 FILLER_18_22 ();
 sg13g2_fill_2 FILLER_18_54 ();
 sg13g2_fill_1 FILLER_18_71 ();
 sg13g2_decap_4 FILLER_18_76 ();
 sg13g2_fill_2 FILLER_18_80 ();
 sg13g2_decap_4 FILLER_18_90 ();
 sg13g2_fill_1 FILLER_18_94 ();
 sg13g2_fill_1 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_138 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_fill_2 FILLER_18_204 ();
 sg13g2_fill_1 FILLER_18_206 ();
 sg13g2_fill_1 FILLER_18_235 ();
 sg13g2_decap_4 FILLER_18_330 ();
 sg13g2_fill_1 FILLER_18_339 ();
 sg13g2_fill_2 FILLER_18_348 ();
 sg13g2_fill_1 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_fill_2 FILLER_18_397 ();
 sg13g2_fill_1 FILLER_18_399 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_20 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_99 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_136 ();
 sg13g2_fill_1 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_193 ();
 sg13g2_fill_2 FILLER_19_295 ();
 sg13g2_fill_1 FILLER_19_297 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_decap_4 FILLER_19_378 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_147 ();
 sg13g2_decap_4 FILLER_20_213 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_241 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_fill_2 FILLER_20_276 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_fill_2 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_370 ();
 sg13g2_fill_2 FILLER_21_36 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_75 ();
 sg13g2_fill_1 FILLER_21_134 ();
 sg13g2_fill_2 FILLER_21_149 ();
 sg13g2_fill_1 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_decap_8 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_fill_2 FILLER_21_221 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_fill_2 FILLER_21_242 ();
 sg13g2_fill_1 FILLER_21_253 ();
 sg13g2_fill_2 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_265 ();
 sg13g2_fill_2 FILLER_21_310 ();
 sg13g2_fill_1 FILLER_21_312 ();
 sg13g2_decap_4 FILLER_21_351 ();
 sg13g2_fill_2 FILLER_21_359 ();
 sg13g2_fill_1 FILLER_21_361 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_fill_1 FILLER_22_19 ();
 sg13g2_fill_2 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_35 ();
 sg13g2_decap_4 FILLER_22_170 ();
 sg13g2_fill_2 FILLER_22_174 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_decap_4 FILLER_22_229 ();
 sg13g2_fill_1 FILLER_22_233 ();
 sg13g2_decap_4 FILLER_22_288 ();
 sg13g2_fill_1 FILLER_22_305 ();
 sg13g2_fill_2 FILLER_22_316 ();
 sg13g2_fill_1 FILLER_22_323 ();
 sg13g2_fill_2 FILLER_22_346 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_fill_1 FILLER_22_394 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_4 ();
 sg13g2_fill_1 FILLER_23_9 ();
 sg13g2_fill_1 FILLER_23_40 ();
 sg13g2_fill_2 FILLER_23_72 ();
 sg13g2_fill_2 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_133 ();
 sg13g2_fill_1 FILLER_23_135 ();
 sg13g2_decap_8 FILLER_23_174 ();
 sg13g2_decap_8 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_fill_1 FILLER_23_335 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_1 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_24_34 ();
 sg13g2_fill_1 FILLER_24_36 ();
 sg13g2_fill_1 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_107 ();
 sg13g2_fill_2 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_128 ();
 sg13g2_fill_2 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_362 ();
 sg13g2_fill_2 FILLER_24_388 ();
 sg13g2_fill_1 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_74 ();
 sg13g2_fill_2 FILLER_25_99 ();
 sg13g2_fill_1 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_191 ();
 sg13g2_fill_1 FILLER_25_228 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_348 ();
 sg13g2_fill_2 FILLER_25_355 ();
 sg13g2_fill_2 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_fill_1 FILLER_25_384 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_fill_2 FILLER_26_201 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_219 ();
 sg13g2_fill_1 FILLER_26_221 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_fill_2 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_fill_1 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_339 ();
 sg13g2_decap_8 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_27_44 ();
 sg13g2_fill_1 FILLER_27_50 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_1 FILLER_27_111 ();
 sg13g2_fill_2 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_fill_2 FILLER_27_227 ();
 sg13g2_fill_1 FILLER_27_229 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_332 ();
 sg13g2_fill_1 FILLER_28_25 ();
 sg13g2_fill_2 FILLER_28_48 ();
 sg13g2_fill_1 FILLER_28_75 ();
 sg13g2_fill_1 FILLER_28_90 ();
 sg13g2_fill_2 FILLER_28_122 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_fill_1 FILLER_28_307 ();
 sg13g2_decap_4 FILLER_28_317 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_fill_2 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_fill_2 FILLER_28_394 ();
 sg13g2_fill_1 FILLER_29_16 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_fill_1 FILLER_29_74 ();
 sg13g2_fill_1 FILLER_29_79 ();
 sg13g2_fill_2 FILLER_29_173 ();
 sg13g2_fill_2 FILLER_29_237 ();
 sg13g2_fill_1 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_263 ();
 sg13g2_fill_2 FILLER_29_383 ();
 sg13g2_fill_2 FILLER_29_398 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_2 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_fill_2 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_45 ();
 sg13g2_fill_2 FILLER_31_76 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_fill_1 FILLER_31_243 ();
 sg13g2_fill_2 FILLER_31_324 ();
 sg13g2_fill_1 FILLER_31_326 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_5 ();
 sg13g2_decap_8 FILLER_32_12 ();
 sg13g2_fill_2 FILLER_32_37 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_fill_2 FILLER_32_69 ();
 sg13g2_fill_2 FILLER_32_102 ();
 sg13g2_fill_1 FILLER_32_104 ();
 sg13g2_fill_1 FILLER_32_112 ();
 sg13g2_decap_4 FILLER_32_177 ();
 sg13g2_fill_2 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_186 ();
 sg13g2_fill_2 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_decap_4 FILLER_32_200 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_fill_2 FILLER_32_245 ();
 sg13g2_fill_1 FILLER_32_273 ();
 sg13g2_fill_2 FILLER_32_348 ();
 sg13g2_fill_1 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_16 ();
 sg13g2_fill_1 FILLER_33_64 ();
 sg13g2_fill_1 FILLER_33_146 ();
 sg13g2_fill_2 FILLER_33_152 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_decap_8 FILLER_33_174 ();
 sg13g2_decap_8 FILLER_33_181 ();
 sg13g2_decap_4 FILLER_33_188 ();
 sg13g2_decap_4 FILLER_33_201 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_fill_2 FILLER_33_219 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_fill_2 FILLER_33_268 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_289 ();
 sg13g2_fill_1 FILLER_33_374 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_1 FILLER_34_39 ();
 sg13g2_fill_1 FILLER_34_66 ();
 sg13g2_fill_1 FILLER_34_110 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_decap_8 FILLER_34_164 ();
 sg13g2_decap_8 FILLER_34_171 ();
 sg13g2_fill_2 FILLER_34_178 ();
 sg13g2_fill_2 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_218 ();
 sg13g2_fill_2 FILLER_34_243 ();
 sg13g2_fill_2 FILLER_34_258 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_fill_2 FILLER_34_312 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_fill_1 FILLER_34_390 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_52 ();
 sg13g2_decap_8 FILLER_35_58 ();
 sg13g2_decap_8 FILLER_35_65 ();
 sg13g2_decap_8 FILLER_35_72 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_decap_4 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_88 ();
 sg13g2_decap_4 FILLER_35_107 ();
 sg13g2_fill_1 FILLER_35_115 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_decap_4 FILLER_35_167 ();
 sg13g2_fill_2 FILLER_35_171 ();
 sg13g2_decap_8 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_211 ();
 sg13g2_decap_4 FILLER_35_218 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_286 ();
 sg13g2_decap_4 FILLER_35_331 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_24 ();
 sg13g2_fill_2 FILLER_36_30 ();
 sg13g2_decap_8 FILLER_36_50 ();
 sg13g2_decap_8 FILLER_36_57 ();
 sg13g2_decap_8 FILLER_36_64 ();
 sg13g2_decap_8 FILLER_36_71 ();
 sg13g2_fill_2 FILLER_36_78 ();
 sg13g2_fill_1 FILLER_36_84 ();
 sg13g2_decap_4 FILLER_36_104 ();
 sg13g2_fill_2 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_140 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_204 ();
 sg13g2_decap_4 FILLER_36_234 ();
 sg13g2_fill_2 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_15 ();
 sg13g2_fill_2 FILLER_37_27 ();
 sg13g2_fill_1 FILLER_37_29 ();
 sg13g2_fill_2 FILLER_37_43 ();
 sg13g2_fill_1 FILLER_37_45 ();
 sg13g2_decap_8 FILLER_37_59 ();
 sg13g2_fill_2 FILLER_37_66 ();
 sg13g2_decap_8 FILLER_37_124 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_decap_8 FILLER_37_138 ();
 sg13g2_decap_4 FILLER_37_145 ();
 sg13g2_fill_2 FILLER_37_149 ();
 sg13g2_fill_2 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_241 ();
 sg13g2_fill_2 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_333 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_376 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_65 ();
 sg13g2_fill_1 FILLER_38_98 ();
 sg13g2_decap_4 FILLER_38_125 ();
 sg13g2_fill_2 FILLER_38_129 ();
 sg13g2_decap_4 FILLER_38_135 ();
 sg13g2_fill_2 FILLER_38_139 ();
 sg13g2_decap_8 FILLER_38_149 ();
 sg13g2_decap_8 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_163 ();
 sg13g2_fill_1 FILLER_38_206 ();
 sg13g2_fill_1 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_246 ();
 sg13g2_fill_2 FILLER_38_260 ();
 sg13g2_fill_2 FILLER_38_322 ();
 sg13g2_decap_4 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_385 ();
 sg13g2_fill_2 FILLER_38_390 ();
 sg13g2_fill_2 FILLER_38_396 ();
 sg13g2_fill_2 FILLER_38_402 ();
 sg13g2_fill_1 FILLER_38_404 ();
 sg13g2_fill_2 FILLER_39_45 ();
 sg13g2_fill_2 FILLER_39_83 ();
 sg13g2_decap_4 FILLER_39_157 ();
 sg13g2_fill_1 FILLER_39_161 ();
 sg13g2_fill_2 FILLER_39_200 ();
 sg13g2_fill_1 FILLER_39_202 ();
 sg13g2_fill_2 FILLER_39_213 ();
 sg13g2_fill_2 FILLER_39_254 ();
 sg13g2_fill_2 FILLER_39_291 ();
 sg13g2_fill_2 FILLER_39_307 ();
 sg13g2_fill_1 FILLER_39_309 ();
 sg13g2_decap_4 FILLER_39_328 ();
 sg13g2_fill_1 FILLER_39_332 ();
 sg13g2_fill_1 FILLER_40_73 ();
 sg13g2_fill_2 FILLER_40_171 ();
 sg13g2_fill_2 FILLER_40_189 ();
 sg13g2_decap_4 FILLER_40_215 ();
 sg13g2_fill_1 FILLER_40_219 ();
 sg13g2_fill_1 FILLER_40_238 ();
 sg13g2_fill_2 FILLER_40_247 ();
 sg13g2_fill_1 FILLER_40_249 ();
 sg13g2_fill_2 FILLER_40_308 ();
 sg13g2_fill_1 FILLER_40_351 ();
 sg13g2_fill_2 FILLER_40_390 ();
 sg13g2_fill_1 FILLER_40_392 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_76 ();
 sg13g2_fill_2 FILLER_41_109 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_fill_2 FILLER_41_131 ();
 sg13g2_fill_2 FILLER_41_169 ();
 sg13g2_fill_1 FILLER_41_171 ();
 sg13g2_decap_8 FILLER_41_205 ();
 sg13g2_decap_8 FILLER_41_212 ();
 sg13g2_decap_4 FILLER_41_219 ();
 sg13g2_fill_1 FILLER_41_228 ();
 sg13g2_fill_2 FILLER_41_242 ();
 sg13g2_fill_2 FILLER_41_252 ();
 sg13g2_fill_1 FILLER_41_254 ();
 sg13g2_fill_2 FILLER_41_262 ();
 sg13g2_fill_2 FILLER_41_356 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_fill_2 FILLER_42_59 ();
 sg13g2_fill_2 FILLER_42_66 ();
 sg13g2_fill_1 FILLER_42_68 ();
 sg13g2_decap_4 FILLER_42_80 ();
 sg13g2_fill_2 FILLER_42_84 ();
 sg13g2_fill_1 FILLER_42_89 ();
 sg13g2_fill_1 FILLER_42_94 ();
 sg13g2_decap_4 FILLER_42_99 ();
 sg13g2_fill_1 FILLER_42_116 ();
 sg13g2_fill_2 FILLER_42_169 ();
 sg13g2_fill_2 FILLER_42_179 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_fill_1 FILLER_42_223 ();
 sg13g2_fill_1 FILLER_42_262 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_4 FILLER_42_287 ();
 sg13g2_fill_1 FILLER_42_291 ();
 sg13g2_decap_8 FILLER_42_305 ();
 sg13g2_decap_8 FILLER_42_325 ();
 sg13g2_decap_4 FILLER_42_332 ();
 sg13g2_fill_1 FILLER_42_336 ();
 sg13g2_fill_1 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_365 ();
 sg13g2_fill_2 FILLER_42_372 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_4 ();
 sg13g2_fill_1 FILLER_43_16 ();
 sg13g2_fill_2 FILLER_43_61 ();
 sg13g2_fill_1 FILLER_43_63 ();
 sg13g2_fill_2 FILLER_43_127 ();
 sg13g2_fill_1 FILLER_43_129 ();
 sg13g2_decap_4 FILLER_43_142 ();
 sg13g2_fill_1 FILLER_43_146 ();
 sg13g2_decap_4 FILLER_43_178 ();
 sg13g2_fill_2 FILLER_43_182 ();
 sg13g2_fill_2 FILLER_43_192 ();
 sg13g2_fill_1 FILLER_43_194 ();
 sg13g2_fill_2 FILLER_43_221 ();
 sg13g2_fill_1 FILLER_43_312 ();
 sg13g2_decap_4 FILLER_43_323 ();
 sg13g2_fill_2 FILLER_43_327 ();
 sg13g2_fill_2 FILLER_43_333 ();
 sg13g2_fill_1 FILLER_43_335 ();
 sg13g2_fill_1 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_4 FILLER_44_7 ();
 sg13g2_fill_2 FILLER_44_15 ();
 sg13g2_decap_8 FILLER_44_22 ();
 sg13g2_fill_2 FILLER_44_41 ();
 sg13g2_fill_2 FILLER_44_63 ();
 sg13g2_fill_2 FILLER_44_109 ();
 sg13g2_fill_1 FILLER_44_119 ();
 sg13g2_fill_1 FILLER_44_139 ();
 sg13g2_fill_2 FILLER_44_150 ();
 sg13g2_decap_8 FILLER_44_174 ();
 sg13g2_fill_1 FILLER_44_181 ();
 sg13g2_decap_4 FILLER_44_211 ();
 sg13g2_fill_2 FILLER_44_238 ();
 sg13g2_fill_1 FILLER_44_248 ();
 sg13g2_fill_2 FILLER_44_252 ();
 sg13g2_decap_4 FILLER_44_299 ();
 sg13g2_fill_2 FILLER_44_329 ();
 sg13g2_fill_1 FILLER_44_351 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_27 ();
 sg13g2_fill_2 FILLER_45_34 ();
 sg13g2_fill_1 FILLER_45_36 ();
 sg13g2_fill_2 FILLER_45_47 ();
 sg13g2_fill_1 FILLER_45_53 ();
 sg13g2_fill_2 FILLER_45_104 ();
 sg13g2_fill_1 FILLER_45_106 ();
 sg13g2_decap_8 FILLER_45_194 ();
 sg13g2_fill_1 FILLER_45_201 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_fill_2 FILLER_45_217 ();
 sg13g2_fill_1 FILLER_45_219 ();
 sg13g2_fill_1 FILLER_45_224 ();
 sg13g2_fill_2 FILLER_45_320 ();
 sg13g2_fill_2 FILLER_45_362 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_54 ();
 sg13g2_fill_1 FILLER_46_56 ();
 sg13g2_fill_1 FILLER_46_103 ();
 sg13g2_fill_1 FILLER_46_113 ();
 sg13g2_fill_2 FILLER_46_159 ();
 sg13g2_fill_2 FILLER_46_223 ();
 sg13g2_fill_1 FILLER_46_225 ();
 sg13g2_fill_2 FILLER_46_230 ();
 sg13g2_fill_1 FILLER_46_232 ();
 sg13g2_fill_1 FILLER_46_241 ();
 sg13g2_decap_4 FILLER_46_251 ();
 sg13g2_fill_1 FILLER_46_304 ();
 sg13g2_fill_1 FILLER_46_353 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_fill_1 FILLER_47_34 ();
 sg13g2_fill_2 FILLER_47_48 ();
 sg13g2_decap_4 FILLER_47_110 ();
 sg13g2_decap_4 FILLER_47_126 ();
 sg13g2_fill_2 FILLER_47_130 ();
 sg13g2_fill_2 FILLER_47_136 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_decap_4 FILLER_47_202 ();
 sg13g2_fill_2 FILLER_47_214 ();
 sg13g2_fill_1 FILLER_47_216 ();
 sg13g2_decap_8 FILLER_47_267 ();
 sg13g2_decap_4 FILLER_47_274 ();
 sg13g2_fill_1 FILLER_47_278 ();
 sg13g2_fill_2 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_322 ();
 sg13g2_fill_1 FILLER_47_342 ();
 sg13g2_fill_2 FILLER_47_398 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_4 ();
 sg13g2_fill_1 FILLER_48_40 ();
 sg13g2_fill_2 FILLER_48_71 ();
 sg13g2_fill_1 FILLER_48_92 ();
 sg13g2_fill_2 FILLER_48_115 ();
 sg13g2_fill_1 FILLER_48_136 ();
 sg13g2_decap_8 FILLER_48_141 ();
 sg13g2_decap_8 FILLER_48_152 ();
 sg13g2_decap_8 FILLER_48_159 ();
 sg13g2_decap_8 FILLER_48_166 ();
 sg13g2_fill_1 FILLER_48_173 ();
 sg13g2_fill_2 FILLER_48_198 ();
 sg13g2_fill_1 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_48_235 ();
 sg13g2_fill_1 FILLER_48_241 ();
 sg13g2_decap_4 FILLER_48_252 ();
 sg13g2_fill_2 FILLER_48_256 ();
 sg13g2_fill_2 FILLER_48_317 ();
 sg13g2_fill_2 FILLER_48_324 ();
 sg13g2_fill_1 FILLER_48_326 ();
 sg13g2_fill_2 FILLER_48_353 ();
 sg13g2_fill_1 FILLER_48_382 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_fill_2 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_81 ();
 sg13g2_fill_1 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_fill_1 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_163 ();
 sg13g2_decap_8 FILLER_49_170 ();
 sg13g2_decap_4 FILLER_49_177 ();
 sg13g2_fill_1 FILLER_49_186 ();
 sg13g2_fill_1 FILLER_49_200 ();
 sg13g2_decap_4 FILLER_49_219 ();
 sg13g2_fill_1 FILLER_49_223 ();
 sg13g2_fill_1 FILLER_49_232 ();
 sg13g2_fill_1 FILLER_49_285 ();
 sg13g2_fill_2 FILLER_49_290 ();
 sg13g2_fill_1 FILLER_49_292 ();
 sg13g2_fill_2 FILLER_49_319 ();
 sg13g2_fill_1 FILLER_49_352 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_fill_2 FILLER_49_371 ();
 sg13g2_fill_1 FILLER_50_26 ();
 sg13g2_fill_2 FILLER_50_61 ();
 sg13g2_fill_1 FILLER_50_132 ();
 sg13g2_fill_2 FILLER_50_164 ();
 sg13g2_fill_2 FILLER_50_180 ();
 sg13g2_fill_1 FILLER_50_182 ();
 sg13g2_decap_8 FILLER_50_187 ();
 sg13g2_fill_2 FILLER_50_194 ();
 sg13g2_decap_8 FILLER_50_211 ();
 sg13g2_decap_8 FILLER_50_218 ();
 sg13g2_decap_4 FILLER_50_225 ();
 sg13g2_fill_2 FILLER_50_247 ();
 sg13g2_fill_1 FILLER_50_249 ();
 sg13g2_fill_1 FILLER_50_274 ();
 sg13g2_fill_2 FILLER_50_347 ();
 sg13g2_fill_1 FILLER_50_349 ();
 sg13g2_fill_1 FILLER_50_392 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_1 FILLER_51_35 ();
 sg13g2_fill_1 FILLER_51_48 ();
 sg13g2_decap_4 FILLER_51_61 ();
 sg13g2_fill_1 FILLER_51_65 ();
 sg13g2_decap_8 FILLER_51_214 ();
 sg13g2_fill_2 FILLER_51_221 ();
 sg13g2_fill_1 FILLER_51_223 ();
 sg13g2_fill_1 FILLER_51_256 ();
 sg13g2_decap_8 FILLER_51_281 ();
 sg13g2_fill_1 FILLER_51_347 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_fill_1 FILLER_52_40 ();
 sg13g2_fill_2 FILLER_52_103 ();
 sg13g2_fill_1 FILLER_52_136 ();
 sg13g2_fill_1 FILLER_52_197 ();
 sg13g2_fill_1 FILLER_52_250 ();
 sg13g2_fill_2 FILLER_52_271 ();
 sg13g2_fill_1 FILLER_52_273 ();
 sg13g2_decap_4 FILLER_52_279 ();
 sg13g2_fill_2 FILLER_52_283 ();
 sg13g2_fill_2 FILLER_52_316 ();
 sg13g2_fill_2 FILLER_52_360 ();
 sg13g2_fill_1 FILLER_52_383 ();
 sg13g2_fill_2 FILLER_52_389 ();
 sg13g2_fill_2 FILLER_53_18 ();
 sg13g2_fill_2 FILLER_53_34 ();
 sg13g2_fill_2 FILLER_53_85 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_fill_1 FILLER_53_92 ();
 sg13g2_fill_2 FILLER_53_124 ();
 sg13g2_fill_1 FILLER_53_126 ();
 sg13g2_fill_2 FILLER_53_161 ();
 sg13g2_fill_1 FILLER_53_163 ();
 sg13g2_fill_2 FILLER_53_174 ();
 sg13g2_fill_2 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_187 ();
 sg13g2_fill_1 FILLER_53_224 ();
 sg13g2_fill_2 FILLER_53_250 ();
 sg13g2_fill_1 FILLER_53_252 ();
 sg13g2_fill_1 FILLER_53_279 ();
 sg13g2_fill_2 FILLER_53_381 ();
 sg13g2_fill_2 FILLER_54_26 ();
 sg13g2_fill_2 FILLER_54_58 ();
 sg13g2_fill_2 FILLER_54_70 ();
 sg13g2_fill_2 FILLER_54_109 ();
 sg13g2_fill_1 FILLER_54_121 ();
 sg13g2_fill_2 FILLER_54_228 ();
 sg13g2_fill_1 FILLER_54_230 ();
 sg13g2_fill_2 FILLER_54_244 ();
 sg13g2_fill_2 FILLER_54_272 ();
 sg13g2_fill_1 FILLER_54_274 ();
 sg13g2_fill_1 FILLER_54_306 ();
 sg13g2_fill_2 FILLER_54_312 ();
 sg13g2_fill_1 FILLER_54_359 ();
 sg13g2_fill_2 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_16 ();
 sg13g2_decap_4 FILLER_55_85 ();
 sg13g2_fill_1 FILLER_55_89 ();
 sg13g2_fill_1 FILLER_55_118 ();
 sg13g2_fill_2 FILLER_55_124 ();
 sg13g2_fill_2 FILLER_55_136 ();
 sg13g2_fill_1 FILLER_55_138 ();
 sg13g2_decap_4 FILLER_55_154 ();
 sg13g2_fill_2 FILLER_55_162 ();
 sg13g2_fill_1 FILLER_55_164 ();
 sg13g2_fill_2 FILLER_55_178 ();
 sg13g2_fill_1 FILLER_55_180 ();
 sg13g2_fill_2 FILLER_55_242 ();
 sg13g2_fill_2 FILLER_55_288 ();
 sg13g2_fill_1 FILLER_55_290 ();
 sg13g2_fill_1 FILLER_55_332 ();
 sg13g2_fill_1 FILLER_55_358 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_fill_2 FILLER_56_36 ();
 sg13g2_fill_1 FILLER_56_38 ();
 sg13g2_fill_2 FILLER_56_145 ();
 sg13g2_fill_2 FILLER_56_173 ();
 sg13g2_fill_1 FILLER_56_175 ();
 sg13g2_decap_4 FILLER_56_200 ();
 sg13g2_fill_1 FILLER_56_230 ();
 sg13g2_fill_1 FILLER_56_276 ();
 sg13g2_fill_1 FILLER_56_312 ();
 sg13g2_fill_1 FILLER_56_346 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_1 FILLER_57_25 ();
 sg13g2_fill_2 FILLER_57_35 ();
 sg13g2_fill_1 FILLER_57_46 ();
 sg13g2_fill_2 FILLER_57_106 ();
 sg13g2_fill_1 FILLER_57_144 ();
 sg13g2_fill_2 FILLER_57_186 ();
 sg13g2_fill_1 FILLER_57_188 ();
 sg13g2_decap_8 FILLER_57_193 ();
 sg13g2_decap_8 FILLER_57_200 ();
 sg13g2_decap_4 FILLER_57_207 ();
 sg13g2_fill_1 FILLER_57_211 ();
 sg13g2_fill_1 FILLER_57_229 ();
 sg13g2_fill_2 FILLER_57_237 ();
 sg13g2_fill_1 FILLER_57_244 ();
 sg13g2_fill_2 FILLER_57_256 ();
 sg13g2_fill_1 FILLER_57_263 ();
 sg13g2_fill_2 FILLER_57_284 ();
 sg13g2_fill_2 FILLER_57_362 ();
 sg13g2_fill_1 FILLER_57_372 ();
 sg13g2_fill_2 FILLER_57_378 ();
 sg13g2_fill_2 FILLER_57_389 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_15 ();
 sg13g2_fill_2 FILLER_58_67 ();
 sg13g2_fill_2 FILLER_58_83 ();
 sg13g2_fill_1 FILLER_58_85 ();
 sg13g2_fill_1 FILLER_58_90 ();
 sg13g2_decap_8 FILLER_58_95 ();
 sg13g2_decap_8 FILLER_58_102 ();
 sg13g2_fill_1 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_198 ();
 sg13g2_decap_8 FILLER_58_205 ();
 sg13g2_decap_4 FILLER_58_212 ();
 sg13g2_fill_1 FILLER_58_216 ();
 sg13g2_fill_2 FILLER_58_271 ();
 sg13g2_fill_1 FILLER_58_312 ();
 sg13g2_fill_1 FILLER_58_372 ();
 sg13g2_fill_2 FILLER_58_387 ();
 sg13g2_fill_1 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_59_50 ();
 sg13g2_fill_2 FILLER_59_69 ();
 sg13g2_fill_1 FILLER_59_107 ();
 sg13g2_fill_1 FILLER_59_124 ();
 sg13g2_fill_1 FILLER_59_150 ();
 sg13g2_fill_2 FILLER_59_164 ();
 sg13g2_decap_4 FILLER_59_202 ();
 sg13g2_fill_1 FILLER_59_206 ();
 sg13g2_fill_1 FILLER_59_229 ();
 sg13g2_fill_1 FILLER_59_246 ();
 sg13g2_fill_2 FILLER_59_321 ();
 sg13g2_fill_1 FILLER_59_326 ();
 sg13g2_fill_1 FILLER_59_357 ();
 sg13g2_fill_1 FILLER_59_398 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_fill_1 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_52 ();
 sg13g2_fill_1 FILLER_60_54 ();
 sg13g2_fill_2 FILLER_60_81 ();
 sg13g2_fill_1 FILLER_60_83 ();
 sg13g2_fill_1 FILLER_60_117 ();
 sg13g2_fill_2 FILLER_60_162 ();
 sg13g2_fill_1 FILLER_60_164 ();
 sg13g2_fill_2 FILLER_60_200 ();
 sg13g2_fill_2 FILLER_60_277 ();
 sg13g2_fill_1 FILLER_60_298 ();
 sg13g2_fill_2 FILLER_60_360 ();
 sg13g2_fill_2 FILLER_60_367 ();
 sg13g2_fill_1 FILLER_61_22 ();
 sg13g2_fill_2 FILLER_61_49 ();
 sg13g2_fill_2 FILLER_61_64 ();
 sg13g2_fill_1 FILLER_61_92 ();
 sg13g2_fill_2 FILLER_61_183 ();
 sg13g2_fill_1 FILLER_61_262 ();
 sg13g2_fill_1 FILLER_61_355 ();
 sg13g2_fill_2 FILLER_61_380 ();
 sg13g2_fill_1 FILLER_61_382 ();
 sg13g2_fill_2 FILLER_62_26 ();
 sg13g2_fill_2 FILLER_62_54 ();
 sg13g2_fill_2 FILLER_62_64 ();
 sg13g2_fill_1 FILLER_62_66 ();
 sg13g2_fill_2 FILLER_62_95 ();
 sg13g2_fill_1 FILLER_62_97 ();
 sg13g2_fill_2 FILLER_62_135 ();
 sg13g2_fill_1 FILLER_62_137 ();
 sg13g2_fill_1 FILLER_62_245 ();
 sg13g2_fill_1 FILLER_62_273 ();
 sg13g2_fill_1 FILLER_62_279 ();
 sg13g2_fill_2 FILLER_62_293 ();
 sg13g2_fill_2 FILLER_62_305 ();
 sg13g2_fill_1 FILLER_62_307 ();
 sg13g2_fill_2 FILLER_62_351 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_27 ();
 sg13g2_fill_2 FILLER_63_49 ();
 sg13g2_fill_1 FILLER_63_63 ();
 sg13g2_fill_1 FILLER_63_108 ();
 sg13g2_fill_1 FILLER_63_141 ();
 sg13g2_fill_1 FILLER_63_151 ();
 sg13g2_fill_1 FILLER_63_171 ();
 sg13g2_decap_4 FILLER_63_209 ();
 sg13g2_fill_1 FILLER_63_213 ();
 sg13g2_decap_8 FILLER_63_222 ();
 sg13g2_decap_8 FILLER_63_229 ();
 sg13g2_fill_2 FILLER_63_236 ();
 sg13g2_fill_1 FILLER_63_238 ();
 sg13g2_fill_2 FILLER_63_257 ();
 sg13g2_fill_1 FILLER_63_259 ();
 sg13g2_fill_2 FILLER_63_310 ();
 sg13g2_fill_1 FILLER_63_312 ();
 sg13g2_fill_1 FILLER_63_318 ();
 sg13g2_fill_1 FILLER_63_377 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_43 ();
 sg13g2_fill_1 FILLER_64_57 ();
 sg13g2_fill_1 FILLER_64_75 ();
 sg13g2_fill_2 FILLER_64_81 ();
 sg13g2_fill_1 FILLER_64_83 ();
 sg13g2_fill_2 FILLER_64_167 ();
 sg13g2_decap_8 FILLER_64_192 ();
 sg13g2_fill_1 FILLER_64_199 ();
 sg13g2_fill_2 FILLER_64_230 ();
 sg13g2_fill_2 FILLER_64_367 ();
 sg13g2_fill_1 FILLER_64_369 ();
 sg13g2_fill_2 FILLER_64_391 ();
 sg13g2_fill_1 FILLER_64_393 ();
 sg13g2_fill_2 FILLER_64_398 ();
 sg13g2_fill_1 FILLER_64_400 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_33 ();
 sg13g2_fill_1 FILLER_65_35 ();
 sg13g2_fill_2 FILLER_65_44 ();
 sg13g2_fill_1 FILLER_65_46 ();
 sg13g2_fill_2 FILLER_65_164 ();
 sg13g2_fill_1 FILLER_65_166 ();
 sg13g2_fill_1 FILLER_65_171 ();
 sg13g2_fill_1 FILLER_65_231 ();
 sg13g2_fill_2 FILLER_65_264 ();
 sg13g2_fill_2 FILLER_65_284 ();
 sg13g2_fill_1 FILLER_65_286 ();
 sg13g2_fill_2 FILLER_65_296 ();
 sg13g2_fill_1 FILLER_65_323 ();
 sg13g2_fill_1 FILLER_65_336 ();
 sg13g2_fill_2 FILLER_65_371 ();
 sg13g2_fill_1 FILLER_65_373 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_55 ();
 sg13g2_fill_1 FILLER_66_57 ();
 sg13g2_fill_2 FILLER_66_73 ();
 sg13g2_fill_2 FILLER_66_173 ();
 sg13g2_decap_8 FILLER_66_204 ();
 sg13g2_fill_1 FILLER_66_229 ();
 sg13g2_fill_2 FILLER_66_339 ();
 sg13g2_fill_1 FILLER_66_341 ();
 sg13g2_fill_2 FILLER_66_375 ();
 sg13g2_fill_1 FILLER_66_377 ();
 sg13g2_fill_1 FILLER_66_382 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_19 ();
 sg13g2_fill_2 FILLER_67_62 ();
 sg13g2_fill_2 FILLER_67_88 ();
 sg13g2_fill_1 FILLER_67_99 ();
 sg13g2_fill_2 FILLER_67_105 ();
 sg13g2_fill_2 FILLER_67_127 ();
 sg13g2_fill_2 FILLER_67_138 ();
 sg13g2_fill_1 FILLER_67_140 ();
 sg13g2_fill_2 FILLER_67_146 ();
 sg13g2_fill_2 FILLER_67_156 ();
 sg13g2_fill_1 FILLER_67_158 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_fill_2 FILLER_67_217 ();
 sg13g2_fill_2 FILLER_67_227 ();
 sg13g2_fill_1 FILLER_67_271 ();
 sg13g2_fill_1 FILLER_67_313 ();
 sg13g2_fill_1 FILLER_67_336 ();
 sg13g2_fill_2 FILLER_67_357 ();
 sg13g2_fill_1 FILLER_67_359 ();
 sg13g2_fill_2 FILLER_67_381 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_1 FILLER_68_44 ();
 sg13g2_fill_1 FILLER_68_70 ();
 sg13g2_fill_1 FILLER_68_80 ();
 sg13g2_fill_1 FILLER_68_115 ();
 sg13g2_decap_4 FILLER_68_158 ();
 sg13g2_decap_8 FILLER_68_185 ();
 sg13g2_decap_4 FILLER_68_192 ();
 sg13g2_fill_1 FILLER_68_196 ();
 sg13g2_decap_8 FILLER_68_200 ();
 sg13g2_decap_4 FILLER_68_207 ();
 sg13g2_fill_1 FILLER_68_281 ();
 sg13g2_fill_1 FILLER_68_291 ();
 sg13g2_fill_2 FILLER_68_381 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_2 ();
 sg13g2_fill_2 FILLER_69_29 ();
 sg13g2_fill_2 FILLER_69_131 ();
 sg13g2_fill_2 FILLER_69_164 ();
 sg13g2_fill_2 FILLER_69_186 ();
 sg13g2_fill_2 FILLER_69_343 ();
 sg13g2_fill_1 FILLER_69_345 ();
 sg13g2_fill_2 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_23 ();
 sg13g2_fill_2 FILLER_70_103 ();
 sg13g2_fill_1 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_183 ();
 sg13g2_decap_8 FILLER_70_190 ();
 sg13g2_fill_2 FILLER_70_197 ();
 sg13g2_decap_4 FILLER_70_203 ();
 sg13g2_fill_1 FILLER_70_207 ();
 sg13g2_fill_1 FILLER_70_213 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_4 ();
 sg13g2_fill_1 FILLER_71_31 ();
 sg13g2_fill_2 FILLER_71_36 ();
 sg13g2_fill_1 FILLER_71_46 ();
 sg13g2_fill_2 FILLER_71_71 ();
 sg13g2_fill_1 FILLER_71_73 ();
 sg13g2_fill_1 FILLER_71_82 ();
 sg13g2_fill_1 FILLER_71_87 ();
 sg13g2_fill_2 FILLER_71_106 ();
 sg13g2_fill_1 FILLER_71_108 ();
 sg13g2_fill_2 FILLER_71_158 ();
 sg13g2_fill_1 FILLER_71_165 ();
 sg13g2_decap_4 FILLER_71_194 ();
 sg13g2_decap_4 FILLER_71_236 ();
 sg13g2_fill_2 FILLER_71_240 ();
 sg13g2_decap_8 FILLER_71_247 ();
 sg13g2_decap_4 FILLER_71_254 ();
 sg13g2_fill_2 FILLER_71_258 ();
 sg13g2_fill_2 FILLER_71_264 ();
 sg13g2_fill_1 FILLER_71_266 ();
 sg13g2_fill_1 FILLER_71_292 ();
 sg13g2_fill_2 FILLER_71_305 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_4 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_11 ();
 sg13g2_fill_2 FILLER_72_41 ();
 sg13g2_fill_1 FILLER_72_60 ();
 sg13g2_fill_2 FILLER_72_75 ();
 sg13g2_fill_2 FILLER_72_116 ();
 sg13g2_fill_1 FILLER_72_118 ();
 sg13g2_fill_2 FILLER_72_128 ();
 sg13g2_decap_4 FILLER_72_203 ();
 sg13g2_fill_2 FILLER_72_207 ();
 sg13g2_fill_2 FILLER_72_213 ();
 sg13g2_fill_1 FILLER_72_215 ();
 sg13g2_fill_2 FILLER_72_228 ();
 sg13g2_fill_1 FILLER_72_230 ();
 sg13g2_fill_2 FILLER_72_239 ();
 sg13g2_fill_1 FILLER_72_252 ();
 sg13g2_fill_1 FILLER_72_282 ();
 sg13g2_fill_2 FILLER_72_292 ();
 sg13g2_fill_1 FILLER_72_294 ();
 sg13g2_fill_1 FILLER_72_347 ();
 sg13g2_decap_4 FILLER_73_26 ();
 sg13g2_fill_2 FILLER_73_77 ();
 sg13g2_fill_1 FILLER_73_79 ();
 sg13g2_fill_2 FILLER_73_123 ();
 sg13g2_fill_1 FILLER_73_125 ();
 sg13g2_fill_2 FILLER_73_159 ();
 sg13g2_fill_1 FILLER_73_166 ();
 sg13g2_fill_1 FILLER_73_177 ();
 sg13g2_fill_2 FILLER_73_188 ();
 sg13g2_fill_1 FILLER_73_190 ();
 sg13g2_decap_8 FILLER_73_201 ();
 sg13g2_fill_2 FILLER_73_208 ();
 sg13g2_fill_1 FILLER_73_210 ();
 sg13g2_fill_1 FILLER_73_253 ();
 sg13g2_fill_2 FILLER_73_270 ();
 sg13g2_fill_1 FILLER_73_303 ();
 sg13g2_fill_2 FILLER_73_325 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_4 ();
 sg13g2_fill_1 FILLER_74_49 ();
 sg13g2_fill_2 FILLER_74_132 ();
 sg13g2_fill_1 FILLER_74_134 ();
 sg13g2_fill_2 FILLER_74_159 ();
 sg13g2_decap_4 FILLER_74_165 ();
 sg13g2_fill_1 FILLER_74_169 ();
 sg13g2_fill_1 FILLER_74_191 ();
 sg13g2_decap_8 FILLER_74_200 ();
 sg13g2_decap_8 FILLER_74_207 ();
 sg13g2_fill_2 FILLER_74_214 ();
 sg13g2_fill_2 FILLER_74_234 ();
 sg13g2_fill_1 FILLER_74_236 ();
 sg13g2_fill_2 FILLER_74_242 ();
 sg13g2_fill_1 FILLER_74_257 ();
 sg13g2_fill_2 FILLER_74_281 ();
 sg13g2_fill_1 FILLER_74_283 ();
 sg13g2_fill_1 FILLER_74_370 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_28 ();
 sg13g2_fill_2 FILLER_75_40 ();
 sg13g2_fill_1 FILLER_75_42 ();
 sg13g2_fill_2 FILLER_75_52 ();
 sg13g2_fill_1 FILLER_75_54 ();
 sg13g2_fill_2 FILLER_75_156 ();
 sg13g2_fill_1 FILLER_75_158 ();
 sg13g2_decap_4 FILLER_75_222 ();
 sg13g2_fill_1 FILLER_75_234 ();
 sg13g2_fill_2 FILLER_75_259 ();
 sg13g2_fill_1 FILLER_75_266 ();
 sg13g2_fill_2 FILLER_75_272 ();
 sg13g2_fill_1 FILLER_75_284 ();
 sg13g2_fill_1 FILLER_75_317 ();
 sg13g2_fill_2 FILLER_75_364 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_4 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_4 ();
 sg13g2_fill_2 FILLER_76_45 ();
 sg13g2_fill_1 FILLER_76_112 ();
 sg13g2_fill_1 FILLER_76_138 ();
 sg13g2_fill_2 FILLER_76_159 ();
 sg13g2_fill_1 FILLER_76_161 ();
 sg13g2_fill_2 FILLER_76_189 ();
 sg13g2_fill_2 FILLER_76_204 ();
 sg13g2_fill_1 FILLER_76_206 ();
 sg13g2_decap_8 FILLER_76_211 ();
 sg13g2_decap_4 FILLER_76_218 ();
 sg13g2_fill_2 FILLER_76_222 ();
 sg13g2_fill_2 FILLER_76_236 ();
 sg13g2_fill_1 FILLER_76_238 ();
 sg13g2_fill_2 FILLER_76_272 ();
 sg13g2_fill_1 FILLER_76_274 ();
 sg13g2_fill_2 FILLER_76_338 ();
 sg13g2_fill_2 FILLER_76_349 ();
 sg13g2_fill_2 FILLER_76_360 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_4 FILLER_77_14 ();
 sg13g2_fill_1 FILLER_77_67 ();
 sg13g2_fill_2 FILLER_77_151 ();
 sg13g2_fill_1 FILLER_77_153 ();
 sg13g2_fill_2 FILLER_77_184 ();
 sg13g2_decap_8 FILLER_77_208 ();
 sg13g2_decap_4 FILLER_77_215 ();
 sg13g2_fill_1 FILLER_77_240 ();
 sg13g2_fill_2 FILLER_77_273 ();
 sg13g2_fill_2 FILLER_77_368 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_7 ();
 sg13g2_fill_2 FILLER_78_154 ();
 sg13g2_fill_1 FILLER_78_156 ();
 sg13g2_fill_2 FILLER_78_172 ();
 sg13g2_fill_1 FILLER_78_174 ();
 sg13g2_fill_2 FILLER_78_294 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_36 ();
 sg13g2_fill_1 FILLER_79_38 ();
 sg13g2_fill_2 FILLER_79_80 ();
 sg13g2_fill_2 FILLER_79_115 ();
 sg13g2_fill_1 FILLER_79_117 ();
 sg13g2_fill_2 FILLER_79_147 ();
 sg13g2_fill_1 FILLER_79_149 ();
 sg13g2_fill_2 FILLER_79_181 ();
 sg13g2_fill_2 FILLER_79_225 ();
 sg13g2_fill_1 FILLER_79_227 ();
 sg13g2_fill_2 FILLER_79_232 ();
 sg13g2_fill_1 FILLER_79_246 ();
 sg13g2_fill_2 FILLER_79_343 ();
 sg13g2_fill_2 FILLER_80_40 ();
 sg13g2_fill_1 FILLER_80_42 ();
 sg13g2_fill_2 FILLER_80_99 ();
 sg13g2_fill_1 FILLER_80_119 ();
 sg13g2_decap_4 FILLER_80_177 ();
 sg13g2_decap_8 FILLER_80_185 ();
 sg13g2_decap_8 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_199 ();
 sg13g2_decap_8 FILLER_80_210 ();
 sg13g2_fill_2 FILLER_80_292 ();
 sg13g2_fill_1 FILLER_80_294 ();
 sg13g2_fill_2 FILLER_80_313 ();
 sg13g2_fill_1 FILLER_80_315 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_2 FILLER_80_393 ();
 assign uio_oe[0] = net376;
 assign uio_oe[1] = net377;
 assign uio_oe[2] = net378;
 assign uio_oe[3] = net379;
 assign uio_oe[4] = net2;
 assign uio_oe[5] = net3;
 assign uio_oe[6] = net4;
 assign uio_oe[7] = net5;
 assign uio_out[4] = net6;
 assign uio_out[5] = net7;
 assign uio_out[6] = net8;
 assign uio_out[7] = net9;
endmodule

module tt_um_rejunity_vga_logo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \grad1.acc[0] ;
 wire \grad1.acc[1] ;
 wire \grad1.acc[2] ;
 wire \grad1.acc[3] ;
 wire \grad1.acc[4] ;
 wire \grad1.acc[5] ;
 wire \grad1.acc[6] ;
 wire \grad1.acc[7] ;
 wire \grad1.acc[8] ;
 wire \grad1.lfsr[0] ;
 wire \grad1.lfsr[10] ;
 wire \grad1.lfsr[11] ;
 wire \grad1.lfsr[12] ;
 wire \grad1.lfsr[13] ;
 wire \grad1.lfsr[14] ;
 wire \grad1.lfsr[15] ;
 wire \grad1.lfsr[16] ;
 wire \grad1.lfsr[17] ;
 wire \grad1.lfsr[18] ;
 wire \grad1.lfsr[19] ;
 wire \grad1.lfsr[1] ;
 wire \grad1.lfsr[2] ;
 wire \grad1.lfsr[3] ;
 wire \grad1.lfsr[4] ;
 wire \grad1.lfsr[5] ;
 wire \grad1.lfsr[6] ;
 wire \grad1.lfsr[7] ;
 wire \grad1.lfsr[8] ;
 wire \grad1.lfsr[9] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \r[0] ;
 wire \r[10] ;
 wire \r[11] ;
 wire \r[12] ;
 wire \r[13] ;
 wire \r[14] ;
 wire \r[15] ;
 wire \r[16] ;
 wire \r[1] ;
 wire \r[2] ;
 wire \r[3] ;
 wire \r[4] ;
 wire \r[5] ;
 wire \r[6] ;
 wire \r[7] ;
 wire \r[8] ;
 wire \r[9] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire vsync_prev;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net1;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;

 sg13g2_inv_1 _0970_ (.Y(_0105_),
    .A(net105));
 sg13g2_inv_2 _0971_ (.Y(_0106_),
    .A(net156));
 sg13g2_inv_1 _0972_ (.Y(_0107_),
    .A(\r[13] ));
 sg13g2_inv_1 _0973_ (.Y(_0108_),
    .A(\counter[5] ));
 sg13g2_inv_1 _0974_ (.Y(_0109_),
    .A(\counter[3] ));
 sg13g2_inv_1 _0975_ (.Y(_0110_),
    .A(\counter[1] ));
 sg13g2_inv_1 _0976_ (.Y(_0111_),
    .A(net124));
 sg13g2_inv_2 _0977_ (.Y(_0112_),
    .A(net195));
 sg13g2_inv_2 _0978_ (.Y(_0113_),
    .A(\hvsync_gen.hpos[7] ));
 sg13g2_inv_2 _0979_ (.Y(_0114_),
    .A(net175));
 sg13g2_inv_1 _0980_ (.Y(_0115_),
    .A(net183));
 sg13g2_inv_1 _0981_ (.Y(_0116_),
    .A(_0009_));
 sg13g2_inv_1 _0982_ (.Y(_0117_),
    .A(net185));
 sg13g2_inv_2 _0983_ (.Y(_0118_),
    .A(net190));
 sg13g2_inv_2 _0984_ (.Y(_0119_),
    .A(net188));
 sg13g2_inv_2 _0985_ (.Y(_0120_),
    .A(net226));
 sg13g2_inv_1 _0986_ (.Y(_0121_),
    .A(\hvsync_gen.vpos[0] ));
 sg13g2_inv_1 _0987_ (.Y(_0122_),
    .A(net200));
 sg13g2_inv_2 _0988_ (.Y(_0123_),
    .A(net193));
 sg13g2_inv_2 _0989_ (.Y(_0124_),
    .A(net215));
 sg13g2_inv_1 _0990_ (.Y(_0125_),
    .A(\grad1.acc[6] ));
 sg13g2_inv_1 _0991_ (.Y(_0126_),
    .A(\grad1.acc[4] ));
 sg13g2_inv_1 _0992_ (.Y(_0127_),
    .A(\grad1.acc[3] ));
 sg13g2_inv_1 _0993_ (.Y(_0128_),
    .A(\grad1.acc[0] ));
 sg13g2_inv_1 _0994_ (.Y(_0129_),
    .A(_0022_));
 sg13g2_nand2_2 _0995_ (.Y(_0130_),
    .A(net179),
    .B(\hvsync_gen.vpos[6] ));
 sg13g2_nor2_1 _0996_ (.A(_0009_),
    .B(_0130_),
    .Y(_0131_));
 sg13g2_nand2_1 _0997_ (.Y(_0132_),
    .A(net183),
    .B(_0117_));
 sg13g2_nor2_1 _0998_ (.A(_0130_),
    .B(_0132_),
    .Y(_0133_));
 sg13g2_nor2_2 _0999_ (.A(_0118_),
    .B(_0119_),
    .Y(_0134_));
 sg13g2_nor2_2 _1000_ (.A(_0120_),
    .B(_0121_),
    .Y(_0135_));
 sg13g2_o21ai_1 _1001_ (.B1(net187),
    .Y(_0136_),
    .A1(net189),
    .A2(_0135_));
 sg13g2_nand2_1 _1002_ (.Y(_0137_),
    .A(_0133_),
    .B(_0136_));
 sg13g2_nor2_1 _1003_ (.A(_0120_),
    .B(\hvsync_gen.vpos[0] ),
    .Y(_0138_));
 sg13g2_nor4_1 _1004_ (.A(net189),
    .B(_0119_),
    .C(_0120_),
    .D(\hvsync_gen.vpos[0] ),
    .Y(_0139_));
 sg13g2_a22oi_1 _1005_ (.Y(_0140_),
    .B1(_0139_),
    .B2(_0133_),
    .A2(_0137_),
    .A1(_0131_));
 sg13g2_nand2_1 _1006_ (.Y(_0141_),
    .A(net177),
    .B(_0114_));
 sg13g2_nand2_2 _1007_ (.Y(_0142_),
    .A(net176),
    .B(net178));
 sg13g2_nand3_1 _1008_ (.B(net178),
    .C(net180),
    .A(net176),
    .Y(_0143_));
 sg13g2_o21ai_1 _1009_ (.B1(net131),
    .Y(_0144_),
    .A1(net184),
    .A2(_0134_));
 sg13g2_inv_1 _1010_ (.Y(_0145_),
    .A(_0144_));
 sg13g2_nor4_1 _1011_ (.A(_0130_),
    .B(_0140_),
    .C(_0141_),
    .D(_0145_),
    .Y(_0001_));
 sg13g2_nand2_2 _1012_ (.Y(_0146_),
    .A(\hvsync_gen.hpos[7] ),
    .B(net197));
 sg13g2_nand2_1 _1013_ (.Y(_0147_),
    .A(net200),
    .B(net198));
 sg13g2_or2_1 _1014_ (.X(_0148_),
    .B(_0147_),
    .A(_0146_));
 sg13g2_a21oi_1 _1015_ (.A1(_0112_),
    .A2(_0148_),
    .Y(_0149_),
    .B1(net149));
 sg13g2_or2_2 _1016_ (.X(_0150_),
    .B(net198),
    .A(net200));
 sg13g2_o21ai_1 _1017_ (.B1(\hvsync_gen.hpos[7] ),
    .Y(_0151_),
    .A1(net196),
    .A2(_0150_));
 sg13g2_and2_1 _1018_ (.A(_0112_),
    .B(_0151_),
    .X(_0152_));
 sg13g2_nor3_1 _1019_ (.A(_0123_),
    .B(_0149_),
    .C(_0152_),
    .Y(_0000_));
 sg13g2_nor2b_2 _1020_ (.A(vsync_prev),
    .B_N(net101),
    .Y(_0153_));
 sg13g2_o21ai_1 _1021_ (.B1(net215),
    .Y(_0154_),
    .A1(\counter[0] ),
    .A2(_0153_));
 sg13g2_a21oi_1 _1022_ (.A1(_0111_),
    .A2(_0153_),
    .Y(_0027_),
    .B1(_0154_));
 sg13g2_a21oi_1 _1023_ (.A1(net134),
    .A2(_0153_),
    .Y(_0155_),
    .B1(\counter[1] ));
 sg13g2_nand3_1 _1024_ (.B(net134),
    .C(_0153_),
    .A(\counter[1] ),
    .Y(_0156_));
 sg13g2_inv_1 _1025_ (.Y(_0157_),
    .A(_0156_));
 sg13g2_nor3_1 _1026_ (.A(net208),
    .B(net135),
    .C(_0157_),
    .Y(_0028_));
 sg13g2_o21ai_1 _1027_ (.B1(net215),
    .Y(_0158_),
    .A1(net129),
    .A2(_0157_));
 sg13g2_a21oi_1 _1028_ (.A1(net129),
    .A2(_0157_),
    .Y(_0029_),
    .B1(_0158_));
 sg13g2_nor2_1 _1029_ (.A(_0022_),
    .B(_0156_),
    .Y(_0159_));
 sg13g2_o21ai_1 _1030_ (.B1(net215),
    .Y(_0160_),
    .A1(net142),
    .A2(_0159_));
 sg13g2_a21oi_1 _1031_ (.A1(net142),
    .A2(_0159_),
    .Y(_0030_),
    .B1(_0160_));
 sg13g2_nand3_1 _1032_ (.B(\counter[2] ),
    .C(_0157_),
    .A(\counter[3] ),
    .Y(_0161_));
 sg13g2_xor2_1 _1033_ (.B(_0161_),
    .A(net138),
    .X(_0162_));
 sg13g2_nor2_1 _1034_ (.A(_0124_),
    .B(net139),
    .Y(_0031_));
 sg13g2_nor2_1 _1035_ (.A(_0021_),
    .B(_0161_),
    .Y(_0163_));
 sg13g2_o21ai_1 _1036_ (.B1(net215),
    .Y(_0164_),
    .A1(net116),
    .A2(_0163_));
 sg13g2_a21oi_1 _1037_ (.A1(net116),
    .A2(_0163_),
    .Y(_0032_),
    .B1(_0164_));
 sg13g2_and2_2 _1038_ (.A(net219),
    .B(\hvsync_gen.hpos[0] ),
    .X(_0165_));
 sg13g2_nand2_1 _1039_ (.Y(_0166_),
    .A(net206),
    .B(net204));
 sg13g2_nand3_1 _1040_ (.B(net205),
    .C(_0165_),
    .A(net203),
    .Y(_0167_));
 sg13g2_nand3b_1 _1041_ (.B(net200),
    .C(net195),
    .Y(_0168_),
    .A_N(net198));
 sg13g2_or2_2 _1042_ (.X(_0169_),
    .B(net196),
    .A(\hvsync_gen.hpos[7] ));
 sg13g2_nor4_2 _1043_ (.A(_0123_),
    .B(_0167_),
    .C(_0168_),
    .Y(_0170_),
    .D(_0169_));
 sg13g2_nor2_2 _1044_ (.A(net208),
    .B(_0170_),
    .Y(_0171_));
 sg13g2_nand2b_1 _1045_ (.Y(_0172_),
    .B(net210),
    .A_N(_0170_));
 sg13g2_and2_1 _1046_ (.A(net100),
    .B(_0171_),
    .X(_0033_));
 sg13g2_nor2_1 _1047_ (.A(net206),
    .B(net207),
    .Y(_0173_));
 sg13g2_nor3_1 _1048_ (.A(_0124_),
    .B(net220),
    .C(_0173_),
    .Y(_0034_));
 sg13g2_o21ai_1 _1049_ (.B1(net214),
    .Y(_0174_),
    .A1(net205),
    .A2(_0165_));
 sg13g2_a21oi_1 _1050_ (.A1(net204),
    .A2(_0165_),
    .Y(_0035_),
    .B1(_0174_));
 sg13g2_a21oi_2 _1051_ (.B1(net203),
    .Y(_0175_),
    .A2(net220),
    .A1(net205));
 sg13g2_nand2_1 _1052_ (.Y(_0176_),
    .A(net215),
    .B(_0167_));
 sg13g2_nor2_1 _1053_ (.A(_0175_),
    .B(_0176_),
    .Y(_0036_));
 sg13g2_and2_1 _1054_ (.A(_0122_),
    .B(_0167_),
    .X(_0177_));
 sg13g2_nor2_1 _1055_ (.A(_0122_),
    .B(_0167_),
    .Y(_0178_));
 sg13g2_nor3_1 _1056_ (.A(_0172_),
    .B(_0177_),
    .C(_0178_),
    .Y(_0037_));
 sg13g2_nor2_1 _1057_ (.A(net198),
    .B(_0178_),
    .Y(_0179_));
 sg13g2_nor2_1 _1058_ (.A(_0147_),
    .B(_0167_),
    .Y(_0180_));
 sg13g2_nor3_1 _1059_ (.A(net171),
    .B(_0179_),
    .C(_0180_),
    .Y(_0038_));
 sg13g2_xnor2_1 _1060_ (.Y(_0181_),
    .A(net196),
    .B(_0180_));
 sg13g2_nor2_1 _1061_ (.A(_0172_),
    .B(_0181_),
    .Y(_0039_));
 sg13g2_a21oi_1 _1062_ (.A1(net196),
    .A2(_0180_),
    .Y(_0182_),
    .B1(net218));
 sg13g2_nor3_1 _1063_ (.A(_0146_),
    .B(_0147_),
    .C(_0167_),
    .Y(_0183_));
 sg13g2_nor3_1 _1064_ (.A(net171),
    .B(_0182_),
    .C(_0183_),
    .Y(_0040_));
 sg13g2_nor2_1 _1065_ (.A(net195),
    .B(_0183_),
    .Y(_0184_));
 sg13g2_nand3_1 _1066_ (.B(\hvsync_gen.hpos[7] ),
    .C(net196),
    .A(net195),
    .Y(_0185_));
 sg13g2_nor3_1 _1067_ (.A(_0112_),
    .B(_0148_),
    .C(_0167_),
    .Y(_0186_));
 sg13g2_nor3_1 _1068_ (.A(net171),
    .B(_0184_),
    .C(_0186_),
    .Y(_0041_));
 sg13g2_xnor2_1 _1069_ (.Y(_0187_),
    .A(net193),
    .B(_0186_));
 sg13g2_nor2_1 _1070_ (.A(net171),
    .B(_0187_),
    .Y(_0042_));
 sg13g2_nor2_1 _1071_ (.A(net189),
    .B(net187),
    .Y(_0188_));
 sg13g2_nor2_1 _1072_ (.A(\hvsync_gen.vpos[1] ),
    .B(\hvsync_gen.vpos[0] ),
    .Y(_0189_));
 sg13g2_nand2_1 _1073_ (.Y(_0190_),
    .A(_0120_),
    .B(_0121_));
 sg13g2_nor4_1 _1074_ (.A(net189),
    .B(net187),
    .C(_0141_),
    .D(_0190_),
    .Y(_0191_));
 sg13g2_nor2_1 _1075_ (.A(net177),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_0192_));
 sg13g2_a221oi_1 _1076_ (.B2(_0191_),
    .C1(net175),
    .B1(_0133_),
    .A1(net177),
    .Y(_0193_),
    .A2(_0131_));
 sg13g2_a21oi_1 _1077_ (.A1(_0112_),
    .A2(_0113_),
    .Y(_0194_),
    .B1(_0008_));
 sg13g2_nor2b_2 _1078_ (.A(_0194_),
    .B_N(_0193_),
    .Y(_0195_));
 sg13g2_nand2b_1 _1079_ (.Y(_0196_),
    .B(_0193_),
    .A_N(_0194_));
 sg13g2_nor2_2 _1080_ (.A(net101),
    .B(_0195_),
    .Y(_0197_));
 sg13g2_nand2b_1 _1081_ (.Y(_0198_),
    .B(net170),
    .A_N(\hvsync_gen.vsync ));
 sg13g2_o21ai_1 _1082_ (.B1(net209),
    .Y(_0199_),
    .A1(net137),
    .A2(_0195_));
 sg13g2_a21oi_1 _1083_ (.A1(net137),
    .A2(net167),
    .Y(_0043_),
    .B1(_0199_));
 sg13g2_and2_1 _1084_ (.A(\r[1] ),
    .B(net207),
    .X(_0200_));
 sg13g2_xor2_1 _1085_ (.B(net207),
    .A(\r[1] ),
    .X(_0201_));
 sg13g2_xor2_1 _1086_ (.B(_0201_),
    .A(\r[0] ),
    .X(_0202_));
 sg13g2_or4_1 _1087_ (.A(net206),
    .B(net207),
    .C(net202),
    .D(net204),
    .X(_0203_));
 sg13g2_nor2_1 _1088_ (.A(net195),
    .B(net194),
    .Y(_0204_));
 sg13g2_nand2_2 _1089_ (.Y(_0205_),
    .A(_0112_),
    .B(_0123_));
 sg13g2_nor4_2 _1090_ (.A(_0150_),
    .B(_0169_),
    .C(_0203_),
    .Y(_0206_),
    .D(_0205_));
 sg13g2_or4_2 _1091_ (.A(_0150_),
    .B(_0169_),
    .C(_0203_),
    .D(_0205_),
    .X(_0207_));
 sg13g2_nand2_1 _1092_ (.Y(_0208_),
    .A(\hvsync_gen.vpos[0] ),
    .B(_0206_));
 sg13g2_xnor2_1 _1093_ (.Y(_0209_),
    .A(_0202_),
    .B(_0208_));
 sg13g2_a21oi_1 _1094_ (.A1(_0195_),
    .A2(_0209_),
    .Y(_0210_),
    .B1(net169));
 sg13g2_o21ai_1 _1095_ (.B1(net209),
    .Y(_0211_),
    .A1(net145),
    .A2(net167));
 sg13g2_nor2_1 _1096_ (.A(_0210_),
    .B(_0211_),
    .Y(_0044_));
 sg13g2_nor2_1 _1097_ (.A(net170),
    .B(_0206_),
    .Y(_0212_));
 sg13g2_nand2_2 _1098_ (.Y(_0213_),
    .A(_0195_),
    .B(_0207_));
 sg13g2_nand2_1 _1099_ (.Y(_0214_),
    .A(\r[2] ),
    .B(net206));
 sg13g2_xnor2_1 _1100_ (.Y(_0215_),
    .A(\r[2] ),
    .B(net206));
 sg13g2_a21oi_1 _1101_ (.A1(\r[0] ),
    .A2(_0201_),
    .Y(_0216_),
    .B1(_0200_));
 sg13g2_xor2_1 _1102_ (.B(_0216_),
    .A(_0215_),
    .X(_0217_));
 sg13g2_nor2_1 _1103_ (.A(net170),
    .B(_0207_),
    .Y(_0218_));
 sg13g2_nand2_2 _1104_ (.Y(_0219_),
    .A(_0195_),
    .B(_0206_));
 sg13g2_nand2_1 _1105_ (.Y(_0220_),
    .A(\r[2] ),
    .B(\hvsync_gen.vpos[1] ));
 sg13g2_xnor2_1 _1106_ (.Y(_0221_),
    .A(\r[2] ),
    .B(\hvsync_gen.vpos[1] ));
 sg13g2_nor2_2 _1107_ (.A(\r[1] ),
    .B(\r[0] ),
    .Y(_0222_));
 sg13g2_a21oi_1 _1108_ (.A1(\r[1] ),
    .A2(\r[0] ),
    .Y(_0223_),
    .B1(\hvsync_gen.vpos[0] ));
 sg13g2_o21ai_1 _1109_ (.B1(_0221_),
    .Y(_0224_),
    .A1(_0222_),
    .A2(_0223_));
 sg13g2_or3_1 _1110_ (.A(_0221_),
    .B(_0222_),
    .C(_0223_),
    .X(_0225_));
 sg13g2_and2_1 _1111_ (.A(_0224_),
    .B(_0225_),
    .X(_0226_));
 sg13g2_a22oi_1 _1112_ (.Y(_0227_),
    .B1(net164),
    .B2(_0226_),
    .A2(_0217_),
    .A1(net165));
 sg13g2_o21ai_1 _1113_ (.B1(net209),
    .Y(_0228_),
    .A1(net163),
    .A2(net166));
 sg13g2_a21oi_1 _1114_ (.A1(net166),
    .A2(_0227_),
    .Y(_0045_),
    .B1(_0228_));
 sg13g2_and2_1 _1115_ (.A(\r[3] ),
    .B(net204),
    .X(_0229_));
 sg13g2_xor2_1 _1116_ (.B(net204),
    .A(\r[3] ),
    .X(_0230_));
 sg13g2_o21ai_1 _1117_ (.B1(_0214_),
    .Y(_0231_),
    .A1(_0215_),
    .A2(_0216_));
 sg13g2_a21oi_1 _1118_ (.A1(_0230_),
    .A2(_0231_),
    .Y(_0232_),
    .B1(_0213_));
 sg13g2_o21ai_1 _1119_ (.B1(_0232_),
    .Y(_0233_),
    .A1(_0230_),
    .A2(_0231_));
 sg13g2_nand2_1 _1120_ (.Y(_0234_),
    .A(\r[3] ),
    .B(net191));
 sg13g2_xnor2_1 _1121_ (.Y(_0235_),
    .A(\r[3] ),
    .B(net191));
 sg13g2_and3_1 _1122_ (.X(_0236_),
    .A(_0220_),
    .B(_0225_),
    .C(_0235_));
 sg13g2_a21oi_1 _1123_ (.A1(_0220_),
    .A2(_0225_),
    .Y(_0237_),
    .B1(_0235_));
 sg13g2_nor2_1 _1124_ (.A(_0236_),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_a21oi_1 _1125_ (.A1(net164),
    .A2(_0238_),
    .Y(_0239_),
    .B1(net169));
 sg13g2_o21ai_1 _1126_ (.B1(net209),
    .Y(_0240_),
    .A1(net152),
    .A2(net167));
 sg13g2_a21oi_1 _1127_ (.A1(_0233_),
    .A2(_0239_),
    .Y(_0046_),
    .B1(_0240_));
 sg13g2_and2_1 _1128_ (.A(\r[4] ),
    .B(net202),
    .X(_0241_));
 sg13g2_xor2_1 _1129_ (.B(net202),
    .A(\r[4] ),
    .X(_0242_));
 sg13g2_a21o_1 _1130_ (.A2(_0231_),
    .A1(_0230_),
    .B1(_0229_),
    .X(_0243_));
 sg13g2_o21ai_1 _1131_ (.B1(net165),
    .Y(_0244_),
    .A1(_0242_),
    .A2(_0243_));
 sg13g2_a21o_1 _1132_ (.A2(_0243_),
    .A1(_0242_),
    .B1(_0244_),
    .X(_0245_));
 sg13g2_nand2_1 _1133_ (.Y(_0246_),
    .A(\r[4] ),
    .B(net188));
 sg13g2_xor2_1 _1134_ (.B(net188),
    .A(\r[4] ),
    .X(_0247_));
 sg13g2_nor2b_1 _1135_ (.A(_0234_),
    .B_N(_0247_),
    .Y(_0248_));
 sg13g2_or2_1 _1136_ (.X(_0249_),
    .B(_0247_),
    .A(_0234_));
 sg13g2_nand2_1 _1137_ (.Y(_0250_),
    .A(_0234_),
    .B(_0247_));
 sg13g2_nand2_1 _1138_ (.Y(_0251_),
    .A(_0249_),
    .B(_0250_));
 sg13g2_nor2_1 _1139_ (.A(_0237_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_a221oi_1 _1140_ (.B2(_0250_),
    .C1(_0235_),
    .B1(_0249_),
    .A1(_0220_),
    .Y(_0253_),
    .A2(_0225_));
 sg13g2_nand2_1 _1141_ (.Y(_0254_),
    .A(_0237_),
    .B(_0251_));
 sg13g2_nor2_1 _1142_ (.A(_0219_),
    .B(_0252_),
    .Y(_0255_));
 sg13g2_a21oi_1 _1143_ (.A1(_0254_),
    .A2(_0255_),
    .Y(_0256_),
    .B1(net169));
 sg13g2_o21ai_1 _1144_ (.B1(net209),
    .Y(_0257_),
    .A1(net216),
    .A2(net166));
 sg13g2_a21oi_1 _1145_ (.A1(_0245_),
    .A2(_0256_),
    .Y(_0047_),
    .B1(_0257_));
 sg13g2_a21oi_1 _1146_ (.A1(_0242_),
    .A2(_0243_),
    .Y(_0258_),
    .B1(_0241_));
 sg13g2_nor2_1 _1147_ (.A(net192),
    .B(net200),
    .Y(_0259_));
 sg13g2_xor2_1 _1148_ (.B(net200),
    .A(net192),
    .X(_0260_));
 sg13g2_xnor2_1 _1149_ (.Y(_0261_),
    .A(_0258_),
    .B(_0260_));
 sg13g2_nor2b_1 _1150_ (.A(net186),
    .B_N(net192),
    .Y(_0262_));
 sg13g2_xnor2_1 _1151_ (.Y(_0263_),
    .A(net192),
    .B(net186));
 sg13g2_nand2b_1 _1152_ (.Y(_0264_),
    .B(_0263_),
    .A_N(_0246_));
 sg13g2_xnor2_1 _1153_ (.Y(_0265_),
    .A(_0246_),
    .B(_0263_));
 sg13g2_o21ai_1 _1154_ (.B1(_0265_),
    .Y(_0266_),
    .A1(_0248_),
    .A2(_0253_));
 sg13g2_nor3_1 _1155_ (.A(_0248_),
    .B(_0253_),
    .C(_0265_),
    .Y(_0267_));
 sg13g2_nand2_1 _1156_ (.Y(_0268_),
    .A(net164),
    .B(_0266_));
 sg13g2_o21ai_1 _1157_ (.B1(net166),
    .Y(_0269_),
    .A1(_0267_),
    .A2(_0268_));
 sg13g2_a21oi_1 _1158_ (.A1(net165),
    .A2(_0261_),
    .Y(_0270_),
    .B1(_0269_));
 sg13g2_o21ai_1 _1159_ (.B1(net209),
    .Y(_0271_),
    .A1(net192),
    .A2(net166));
 sg13g2_nor2_1 _1160_ (.A(_0270_),
    .B(_0271_),
    .Y(_0048_));
 sg13g2_and2_1 _1161_ (.A(\r[6] ),
    .B(net198),
    .X(_0272_));
 sg13g2_xnor2_1 _1162_ (.Y(_0273_),
    .A(\r[6] ),
    .B(net198));
 sg13g2_a221oi_1 _1163_ (.B2(_0243_),
    .C1(_0241_),
    .B1(_0242_),
    .A1(\r[5] ),
    .Y(_0274_),
    .A2(net200));
 sg13g2_o21ai_1 _1164_ (.B1(_0273_),
    .Y(_0275_),
    .A1(_0259_),
    .A2(_0274_));
 sg13g2_nor3_1 _1165_ (.A(_0259_),
    .B(_0273_),
    .C(_0274_),
    .Y(_0276_));
 sg13g2_nand3b_1 _1166_ (.B(net165),
    .C(_0275_),
    .Y(_0277_),
    .A_N(_0276_));
 sg13g2_nor2_1 _1167_ (.A(net183),
    .B(_0117_),
    .Y(_0278_));
 sg13g2_xnor2_1 _1168_ (.Y(_0279_),
    .A(net182),
    .B(net186));
 sg13g2_nand2b_1 _1169_ (.Y(_0280_),
    .B(\r[6] ),
    .A_N(_0279_));
 sg13g2_xnor2_1 _1170_ (.Y(_0281_),
    .A(\r[6] ),
    .B(_0279_));
 sg13g2_nand2_1 _1171_ (.Y(_0282_),
    .A(_0262_),
    .B(_0281_));
 sg13g2_xnor2_1 _1172_ (.Y(_0283_),
    .A(_0262_),
    .B(_0281_));
 sg13g2_a21o_1 _1173_ (.A2(_0266_),
    .A1(_0264_),
    .B1(_0283_),
    .X(_0284_));
 sg13g2_nand3_1 _1174_ (.B(_0266_),
    .C(_0283_),
    .A(_0264_),
    .Y(_0285_));
 sg13g2_nand3_1 _1175_ (.B(_0284_),
    .C(_0285_),
    .A(net164),
    .Y(_0286_));
 sg13g2_nand3_1 _1176_ (.B(_0277_),
    .C(_0286_),
    .A(net166),
    .Y(_0287_));
 sg13g2_o21ai_1 _1177_ (.B1(_0287_),
    .Y(_0288_),
    .A1(net223),
    .A2(net166));
 sg13g2_nor2_1 _1178_ (.A(net208),
    .B(_0288_),
    .Y(_0049_));
 sg13g2_nand2b_1 _1179_ (.Y(_0289_),
    .B(\r[7] ),
    .A_N(net197));
 sg13g2_xnor2_1 _1180_ (.Y(_0290_),
    .A(\r[7] ),
    .B(net197));
 sg13g2_o21ai_1 _1181_ (.B1(_0290_),
    .Y(_0291_),
    .A1(_0272_),
    .A2(_0276_));
 sg13g2_or3_1 _1182_ (.A(_0272_),
    .B(_0276_),
    .C(_0290_),
    .X(_0292_));
 sg13g2_nand3_1 _1183_ (.B(_0291_),
    .C(_0292_),
    .A(net165),
    .Y(_0293_));
 sg13g2_nand2_1 _1184_ (.Y(_0294_),
    .A(_0282_),
    .B(_0284_));
 sg13g2_nand3_1 _1185_ (.B(net182),
    .C(net186),
    .A(net180),
    .Y(_0295_));
 sg13g2_a21o_1 _1186_ (.A2(net186),
    .A1(net182),
    .B1(net180),
    .X(_0296_));
 sg13g2_a21oi_1 _1187_ (.A1(_0295_),
    .A2(_0296_),
    .Y(_0297_),
    .B1(\r[7] ));
 sg13g2_nand3_1 _1188_ (.B(_0295_),
    .C(_0296_),
    .A(\r[7] ),
    .Y(_0298_));
 sg13g2_nand2b_1 _1189_ (.Y(_0299_),
    .B(_0298_),
    .A_N(_0297_));
 sg13g2_nor2b_1 _1190_ (.A(_0280_),
    .B_N(_0299_),
    .Y(_0300_));
 sg13g2_xor2_1 _1191_ (.B(_0299_),
    .A(_0280_),
    .X(_0301_));
 sg13g2_a21oi_1 _1192_ (.A1(_0282_),
    .A2(_0284_),
    .Y(_0302_),
    .B1(_0301_));
 sg13g2_xnor2_1 _1193_ (.Y(_0303_),
    .A(_0294_),
    .B(_0301_));
 sg13g2_a21oi_1 _1194_ (.A1(net164),
    .A2(_0303_),
    .Y(_0304_),
    .B1(net169));
 sg13g2_o21ai_1 _1195_ (.B1(net209),
    .Y(_0305_),
    .A1(net162),
    .A2(net166));
 sg13g2_a21oi_1 _1196_ (.A1(_0293_),
    .A2(_0304_),
    .Y(_0050_),
    .B1(_0305_));
 sg13g2_nand2_1 _1197_ (.Y(_0306_),
    .A(_0289_),
    .B(_0291_));
 sg13g2_nand2_1 _1198_ (.Y(_0307_),
    .A(_0146_),
    .B(_0169_));
 sg13g2_nand2b_1 _1199_ (.Y(_0308_),
    .B(_0307_),
    .A_N(\r[8] ));
 sg13g2_nand3_1 _1200_ (.B(_0146_),
    .C(_0169_),
    .A(\r[8] ),
    .Y(_0309_));
 sg13g2_nand2_1 _1201_ (.Y(_0310_),
    .A(_0308_),
    .B(_0309_));
 sg13g2_nand2_1 _1202_ (.Y(_0311_),
    .A(_0306_),
    .B(_0310_));
 sg13g2_xor2_1 _1203_ (.B(_0310_),
    .A(_0306_),
    .X(_0312_));
 sg13g2_xor2_1 _1204_ (.B(_0295_),
    .A(_0012_),
    .X(_0313_));
 sg13g2_xor2_1 _1205_ (.B(_0313_),
    .A(_0023_),
    .X(_0314_));
 sg13g2_nand2b_1 _1206_ (.Y(_0315_),
    .B(_0314_),
    .A_N(_0297_));
 sg13g2_xnor2_1 _1207_ (.Y(_0316_),
    .A(_0297_),
    .B(_0314_));
 sg13g2_o21ai_1 _1208_ (.B1(_0316_),
    .Y(_0317_),
    .A1(_0300_),
    .A2(_0302_));
 sg13g2_nor3_1 _1209_ (.A(_0300_),
    .B(_0302_),
    .C(_0316_),
    .Y(_0318_));
 sg13g2_nor2_1 _1210_ (.A(_0219_),
    .B(_0318_),
    .Y(_0319_));
 sg13g2_a221oi_1 _1211_ (.B2(_0319_),
    .C1(net170),
    .B1(_0317_),
    .A1(_0207_),
    .Y(_0320_),
    .A2(_0312_));
 sg13g2_o21ai_1 _1212_ (.B1(net209),
    .Y(_0321_),
    .A1(net224),
    .A2(net167));
 sg13g2_nor2_1 _1213_ (.A(_0320_),
    .B(_0321_),
    .Y(_0051_));
 sg13g2_nand2_2 _1214_ (.Y(_0322_),
    .A(net195),
    .B(_0169_));
 sg13g2_xnor2_1 _1215_ (.Y(_0323_),
    .A(_0112_),
    .B(_0169_));
 sg13g2_nand2_1 _1216_ (.Y(_0324_),
    .A(\r[9] ),
    .B(_0323_));
 sg13g2_xnor2_1 _1217_ (.Y(_0325_),
    .A(\r[9] ),
    .B(_0323_));
 sg13g2_a221oi_1 _1218_ (.B2(_0309_),
    .C1(_0325_),
    .B1(_0308_),
    .A1(_0289_),
    .Y(_0326_),
    .A2(_0291_));
 sg13g2_or2_1 _1219_ (.X(_0327_),
    .B(_0325_),
    .A(_0311_));
 sg13g2_nand2b_1 _1220_ (.Y(_0328_),
    .B(_0307_),
    .A_N(_0023_));
 sg13g2_and2_1 _1221_ (.A(_0325_),
    .B(_0328_),
    .X(_0329_));
 sg13g2_o21ai_1 _1222_ (.B1(_0212_),
    .Y(_0330_),
    .A1(_0325_),
    .A2(_0328_));
 sg13g2_a21oi_1 _1223_ (.A1(_0311_),
    .A2(_0329_),
    .Y(_0331_),
    .B1(_0330_));
 sg13g2_nand2_1 _1224_ (.Y(_0332_),
    .A(_0315_),
    .B(_0317_));
 sg13g2_nand2_1 _1225_ (.Y(_0333_),
    .A(net178),
    .B(net182));
 sg13g2_nand4_1 _1226_ (.B(net180),
    .C(net182),
    .A(net178),
    .Y(_0334_),
    .D(net186));
 sg13g2_nand2b_1 _1227_ (.Y(_0335_),
    .B(_0334_),
    .A_N(net176));
 sg13g2_o21ai_1 _1228_ (.B1(_0335_),
    .Y(_0336_),
    .A1(_0142_),
    .A2(_0295_));
 sg13g2_nand2_1 _1229_ (.Y(_0337_),
    .A(\r[9] ),
    .B(_0336_));
 sg13g2_xor2_1 _1230_ (.B(_0336_),
    .A(\r[9] ),
    .X(_0338_));
 sg13g2_o21ai_1 _1231_ (.B1(_0338_),
    .Y(_0339_),
    .A1(\r[8] ),
    .A2(_0313_));
 sg13g2_or3_1 _1232_ (.A(\r[8] ),
    .B(_0313_),
    .C(_0338_),
    .X(_0340_));
 sg13g2_inv_1 _1233_ (.Y(_0341_),
    .A(_0340_));
 sg13g2_nand2_1 _1234_ (.Y(_0342_),
    .A(_0339_),
    .B(_0340_));
 sg13g2_xnor2_1 _1235_ (.Y(_0343_),
    .A(_0332_),
    .B(_0342_));
 sg13g2_a221oi_1 _1236_ (.B2(net164),
    .C1(_0197_),
    .B1(_0343_),
    .A1(_0327_),
    .Y(_0344_),
    .A2(_0331_));
 sg13g2_o21ai_1 _1237_ (.B1(net210),
    .Y(_0345_),
    .A1(net230),
    .A2(net168));
 sg13g2_nor2_1 _1238_ (.A(_0344_),
    .B(_0345_),
    .Y(_0052_));
 sg13g2_o21ai_1 _1239_ (.B1(_0324_),
    .Y(_0346_),
    .A1(_0325_),
    .A2(_0328_));
 sg13g2_nor2_1 _1240_ (.A(net193),
    .B(_0322_),
    .Y(_0347_));
 sg13g2_xnor2_1 _1241_ (.Y(_0348_),
    .A(net193),
    .B(_0322_));
 sg13g2_xor2_1 _1242_ (.B(_0348_),
    .A(\r[10] ),
    .X(_0349_));
 sg13g2_inv_1 _1243_ (.Y(_0350_),
    .A(_0349_));
 sg13g2_or3_1 _1244_ (.A(_0326_),
    .B(_0346_),
    .C(_0350_),
    .X(_0351_));
 sg13g2_o21ai_1 _1245_ (.B1(_0350_),
    .Y(_0352_),
    .A1(_0326_),
    .A2(_0346_));
 sg13g2_and2_1 _1246_ (.A(_0212_),
    .B(_0352_),
    .X(_0353_));
 sg13g2_nand2_1 _1247_ (.Y(_0354_),
    .A(_0013_),
    .B(_0334_));
 sg13g2_xnor2_1 _1248_ (.Y(_0355_),
    .A(_0114_),
    .B(_0354_));
 sg13g2_xor2_1 _1249_ (.B(_0355_),
    .A(_0002_),
    .X(_0356_));
 sg13g2_nor2_1 _1250_ (.A(_0337_),
    .B(_0356_),
    .Y(_0357_));
 sg13g2_xnor2_1 _1251_ (.Y(_0358_),
    .A(_0337_),
    .B(_0356_));
 sg13g2_a21o_1 _1252_ (.A2(_0317_),
    .A1(_0315_),
    .B1(_0341_),
    .X(_0359_));
 sg13g2_nand3_1 _1253_ (.B(_0358_),
    .C(_0359_),
    .A(_0339_),
    .Y(_0360_));
 sg13g2_a21o_1 _1254_ (.A2(_0359_),
    .A1(_0339_),
    .B1(_0358_),
    .X(_0361_));
 sg13g2_and2_1 _1255_ (.A(net164),
    .B(_0360_),
    .X(_0362_));
 sg13g2_a221oi_1 _1256_ (.B2(_0362_),
    .C1(_0197_),
    .B1(_0361_),
    .A1(_0351_),
    .Y(_0363_),
    .A2(_0353_));
 sg13g2_o21ai_1 _1257_ (.B1(net210),
    .Y(_0364_),
    .A1(net144),
    .A2(net168));
 sg13g2_nor2_1 _1258_ (.A(_0363_),
    .B(_0364_),
    .Y(_0053_));
 sg13g2_nor2b_1 _1259_ (.A(_0347_),
    .B_N(_0008_),
    .Y(_0365_));
 sg13g2_o21ai_1 _1260_ (.B1(_0008_),
    .Y(_0366_),
    .A1(net193),
    .A2(_0322_));
 sg13g2_nor2_1 _1261_ (.A(_0003_),
    .B(net174),
    .Y(_0367_));
 sg13g2_nand2_1 _1262_ (.Y(_0368_),
    .A(_0003_),
    .B(net174));
 sg13g2_nand2b_1 _1263_ (.Y(_0369_),
    .B(_0368_),
    .A_N(_0367_));
 sg13g2_nor2_1 _1264_ (.A(_0002_),
    .B(_0348_),
    .Y(_0370_));
 sg13g2_o21ai_1 _1265_ (.B1(_0352_),
    .Y(_0371_),
    .A1(_0002_),
    .A2(_0348_));
 sg13g2_xnor2_1 _1266_ (.Y(_0372_),
    .A(_0369_),
    .B(_0371_));
 sg13g2_nand2b_1 _1267_ (.Y(_0373_),
    .B(_0361_),
    .A_N(_0357_));
 sg13g2_nor2b_1 _1268_ (.A(\r[10] ),
    .B_N(_0355_),
    .Y(_0374_));
 sg13g2_nor2_1 _1269_ (.A(net175),
    .B(_0335_),
    .Y(_0375_));
 sg13g2_xor2_1 _1270_ (.B(net172),
    .A(\r[11] ),
    .X(_0376_));
 sg13g2_nor2_1 _1271_ (.A(_0374_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_nand2_1 _1272_ (.Y(_0378_),
    .A(_0374_),
    .B(_0376_));
 sg13g2_nor2b_1 _1273_ (.A(_0377_),
    .B_N(_0378_),
    .Y(_0379_));
 sg13g2_or2_1 _1274_ (.X(_0380_),
    .B(_0379_),
    .A(_0373_));
 sg13g2_a21oi_1 _1275_ (.A1(_0373_),
    .A2(_0379_),
    .Y(_0381_),
    .B1(_0219_));
 sg13g2_a221oi_1 _1276_ (.B2(_0381_),
    .C1(_0197_),
    .B1(_0380_),
    .A1(net165),
    .Y(_0382_),
    .A2(_0372_));
 sg13g2_o21ai_1 _1277_ (.B1(net210),
    .Y(_0383_),
    .A1(net136),
    .A2(net168));
 sg13g2_nor2_1 _1278_ (.A(_0382_),
    .B(_0383_),
    .Y(_0054_));
 sg13g2_nor2_1 _1279_ (.A(_0367_),
    .B(_0370_),
    .Y(_0384_));
 sg13g2_a21oi_1 _1280_ (.A1(_0368_),
    .A2(_0371_),
    .Y(_0385_),
    .B1(_0367_));
 sg13g2_xnor2_1 _1281_ (.Y(_0386_),
    .A(_0004_),
    .B(net174));
 sg13g2_a221oi_1 _1282_ (.B2(_0352_),
    .C1(_0386_),
    .B1(_0384_),
    .A1(_0003_),
    .Y(_0387_),
    .A2(net174));
 sg13g2_xor2_1 _1283_ (.B(_0386_),
    .A(_0385_),
    .X(_0388_));
 sg13g2_nor2_1 _1284_ (.A(_0003_),
    .B(net172),
    .Y(_0389_));
 sg13g2_xnor2_1 _1285_ (.Y(_0390_),
    .A(\r[12] ),
    .B(_0389_));
 sg13g2_inv_1 _1286_ (.Y(_0391_),
    .A(_0390_));
 sg13g2_nor2_1 _1287_ (.A(_0357_),
    .B(_0377_),
    .Y(_0392_));
 sg13g2_a21oi_1 _1288_ (.A1(_0373_),
    .A2(_0378_),
    .Y(_0393_),
    .B1(_0377_));
 sg13g2_a221oi_1 _1289_ (.B2(_0361_),
    .C1(_0391_),
    .B1(_0392_),
    .A1(_0374_),
    .Y(_0394_),
    .A2(_0376_));
 sg13g2_nand2b_1 _1290_ (.Y(_0395_),
    .B(_0390_),
    .A_N(_0393_));
 sg13g2_a21oi_1 _1291_ (.A1(_0391_),
    .A2(_0393_),
    .Y(_0396_),
    .B1(_0219_));
 sg13g2_a221oi_1 _1292_ (.B2(_0396_),
    .C1(net170),
    .B1(_0395_),
    .A1(_0207_),
    .Y(_0397_),
    .A2(_0388_));
 sg13g2_o21ai_1 _1293_ (.B1(net210),
    .Y(_0398_),
    .A1(net217),
    .A2(net168));
 sg13g2_nor2_1 _1294_ (.A(_0397_),
    .B(_0398_),
    .Y(_0055_));
 sg13g2_and2_1 _1295_ (.A(\r[12] ),
    .B(_0365_),
    .X(_0399_));
 sg13g2_nor2_1 _1296_ (.A(_0387_),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_nand2_1 _1297_ (.Y(_0401_),
    .A(net234),
    .B(net174));
 sg13g2_or2_1 _1298_ (.X(_0402_),
    .B(net174),
    .A(_0005_));
 sg13g2_nand2_1 _1299_ (.Y(_0403_),
    .A(_0401_),
    .B(_0402_));
 sg13g2_xnor2_1 _1300_ (.Y(_0404_),
    .A(_0400_),
    .B(_0403_));
 sg13g2_a21oi_1 _1301_ (.A1(_0107_),
    .A2(net169),
    .Y(_0405_),
    .B1(net208));
 sg13g2_mux2_1 _1302_ (.A0(_0389_),
    .A1(net172),
    .S(\r[12] ),
    .X(_0406_));
 sg13g2_nor3_1 _1303_ (.A(\r[13] ),
    .B(_0004_),
    .C(net172),
    .Y(_0407_));
 sg13g2_o21ai_1 _1304_ (.B1(\r[13] ),
    .Y(_0408_),
    .A1(_0004_),
    .A2(net172));
 sg13g2_nor2b_1 _1305_ (.A(_0407_),
    .B_N(_0408_),
    .Y(_0409_));
 sg13g2_nor3_1 _1306_ (.A(_0394_),
    .B(_0406_),
    .C(_0409_),
    .Y(_0410_));
 sg13g2_o21ai_1 _1307_ (.B1(_0409_),
    .Y(_0411_),
    .A1(_0394_),
    .A2(_0406_));
 sg13g2_nor2b_1 _1308_ (.A(_0410_),
    .B_N(_0411_),
    .Y(_0412_));
 sg13g2_o21ai_1 _1309_ (.B1(_0405_),
    .Y(_0413_),
    .A1(_0219_),
    .A2(_0412_));
 sg13g2_a21oi_1 _1310_ (.A1(net165),
    .A2(_0404_),
    .Y(_0056_),
    .B1(_0413_));
 sg13g2_o21ai_1 _1311_ (.B1(_0401_),
    .Y(_0414_),
    .A1(_0387_),
    .A2(_0399_));
 sg13g2_xnor2_1 _1312_ (.Y(_0415_),
    .A(_0006_),
    .B(net174));
 sg13g2_a21oi_2 _1313_ (.B1(_0415_),
    .Y(_0416_),
    .A2(_0414_),
    .A1(_0402_));
 sg13g2_nand3_1 _1314_ (.B(_0414_),
    .C(_0415_),
    .A(_0402_),
    .Y(_0417_));
 sg13g2_nor2_1 _1315_ (.A(_0206_),
    .B(_0416_),
    .Y(_0418_));
 sg13g2_nand2_1 _1316_ (.Y(_0419_),
    .A(_0417_),
    .B(_0418_));
 sg13g2_a21oi_1 _1317_ (.A1(\r[13] ),
    .A2(net172),
    .Y(_0420_),
    .B1(_0407_));
 sg13g2_nor2_1 _1318_ (.A(_0005_),
    .B(net173),
    .Y(_0421_));
 sg13g2_xnor2_1 _1319_ (.Y(_0422_),
    .A(_0106_),
    .B(_0421_));
 sg13g2_a21oi_2 _1320_ (.B1(_0422_),
    .Y(_0423_),
    .A2(_0420_),
    .A1(_0411_));
 sg13g2_and3_1 _1321_ (.X(_0424_),
    .A(_0411_),
    .B(_0420_),
    .C(_0422_));
 sg13g2_nor3_1 _1322_ (.A(_0207_),
    .B(_0423_),
    .C(_0424_),
    .Y(_0425_));
 sg13g2_nor2_1 _1323_ (.A(net170),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_a221oi_1 _1324_ (.B2(_0426_),
    .C1(net208),
    .B1(_0419_),
    .A1(_0106_),
    .Y(_0057_),
    .A2(net169));
 sg13g2_mux2_1 _1325_ (.A0(net173),
    .A1(_0421_),
    .S(_0106_),
    .X(_0427_));
 sg13g2_nor3_1 _1326_ (.A(\r[15] ),
    .B(_0006_),
    .C(net173),
    .Y(_0428_));
 sg13g2_o21ai_1 _1327_ (.B1(\r[15] ),
    .Y(_0429_),
    .A1(_0006_),
    .A2(net173));
 sg13g2_nor2b_1 _1328_ (.A(_0428_),
    .B_N(_0429_),
    .Y(_0430_));
 sg13g2_nor3_1 _1329_ (.A(_0423_),
    .B(_0427_),
    .C(_0430_),
    .Y(_0431_));
 sg13g2_o21ai_1 _1330_ (.B1(_0430_),
    .Y(_0432_),
    .A1(_0423_),
    .A2(_0427_));
 sg13g2_nand3b_1 _1331_ (.B(_0432_),
    .C(_0218_),
    .Y(_0433_),
    .A_N(_0431_));
 sg13g2_xor2_1 _1332_ (.B(net174),
    .A(_0007_),
    .X(_0434_));
 sg13g2_nand2_1 _1333_ (.Y(_0435_),
    .A(_0416_),
    .B(_0434_));
 sg13g2_nor2_1 _1334_ (.A(_0106_),
    .B(_0366_),
    .Y(_0436_));
 sg13g2_nor3_1 _1335_ (.A(_0416_),
    .B(_0434_),
    .C(_0436_),
    .Y(_0437_));
 sg13g2_and3_1 _1336_ (.X(_0438_),
    .A(\r[14] ),
    .B(_0007_),
    .C(_0365_));
 sg13g2_nor3_1 _1337_ (.A(_0213_),
    .B(_0437_),
    .C(_0438_),
    .Y(_0439_));
 sg13g2_a21oi_1 _1338_ (.A1(_0435_),
    .A2(_0439_),
    .Y(_0440_),
    .B1(net169));
 sg13g2_o21ai_1 _1339_ (.B1(net210),
    .Y(_0441_),
    .A1(net155),
    .A2(net168));
 sg13g2_a21oi_1 _1340_ (.A1(_0433_),
    .A2(_0440_),
    .Y(_0058_),
    .B1(_0441_));
 sg13g2_a221oi_1 _1341_ (.B2(_0434_),
    .C1(_0438_),
    .B1(_0416_),
    .A1(\r[15] ),
    .Y(_0442_),
    .A2(_0365_));
 sg13g2_xnor2_1 _1342_ (.Y(_0443_),
    .A(\r[16] ),
    .B(_0366_));
 sg13g2_xnor2_1 _1343_ (.Y(_0444_),
    .A(_0442_),
    .B(_0443_));
 sg13g2_a21oi_1 _1344_ (.A1(\r[15] ),
    .A2(net172),
    .Y(_0445_),
    .B1(_0428_));
 sg13g2_nand2_1 _1345_ (.Y(_0446_),
    .A(_0432_),
    .B(_0445_));
 sg13g2_nor2_1 _1346_ (.A(_0007_),
    .B(net172),
    .Y(_0447_));
 sg13g2_xnor2_1 _1347_ (.Y(_0448_),
    .A(_0010_),
    .B(_0447_));
 sg13g2_xnor2_1 _1348_ (.Y(_0449_),
    .A(_0446_),
    .B(_0448_));
 sg13g2_a221oi_1 _1349_ (.B2(net164),
    .C1(net169),
    .B1(_0449_),
    .A1(net165),
    .Y(_0450_),
    .A2(_0444_));
 sg13g2_o21ai_1 _1350_ (.B1(net210),
    .Y(_0451_),
    .A1(net140),
    .A2(net168));
 sg13g2_nor2_1 _1351_ (.A(_0450_),
    .B(_0451_),
    .Y(_0059_));
 sg13g2_nand2_1 _1352_ (.Y(_0452_),
    .A(net133),
    .B(net122));
 sg13g2_o21ai_1 _1353_ (.B1(net214),
    .Y(_0453_),
    .A1(net133),
    .A2(net122));
 sg13g2_nor2b_1 _1354_ (.A(_0453_),
    .B_N(_0452_),
    .Y(_0060_));
 sg13g2_xnor2_1 _1355_ (.Y(_0454_),
    .A(net222),
    .B(net119));
 sg13g2_and2_1 _1356_ (.A(_0452_),
    .B(_0454_),
    .X(_0455_));
 sg13g2_nor2_1 _1357_ (.A(_0452_),
    .B(_0454_),
    .Y(_0456_));
 sg13g2_nor3_1 _1358_ (.A(net208),
    .B(_0455_),
    .C(_0456_),
    .Y(_0061_));
 sg13g2_xnor2_1 _1359_ (.Y(_0457_),
    .A(net147),
    .B(net120));
 sg13g2_a21oi_1 _1360_ (.A1(net222),
    .A2(net119),
    .Y(_0458_),
    .B1(_0456_));
 sg13g2_and2_1 _1361_ (.A(_0457_),
    .B(_0458_),
    .X(_0459_));
 sg13g2_nor2_1 _1362_ (.A(_0457_),
    .B(_0458_),
    .Y(_0460_));
 sg13g2_nor3_1 _1363_ (.A(net208),
    .B(_0459_),
    .C(_0460_),
    .Y(_0062_));
 sg13g2_xnor2_1 _1364_ (.Y(_0461_),
    .A(\grad1.acc[3] ),
    .B(net127));
 sg13g2_a21oi_1 _1365_ (.A1(net147),
    .A2(net120),
    .Y(_0462_),
    .B1(_0460_));
 sg13g2_or2_1 _1366_ (.X(_0463_),
    .B(_0462_),
    .A(_0461_));
 sg13g2_inv_1 _1367_ (.Y(_0464_),
    .A(_0463_));
 sg13g2_nand2_1 _1368_ (.Y(_0465_),
    .A(net212),
    .B(_0463_));
 sg13g2_a21oi_1 _1369_ (.A1(_0461_),
    .A2(_0462_),
    .Y(_0063_),
    .B1(_0465_));
 sg13g2_nand2_1 _1370_ (.Y(_0466_),
    .A(net150),
    .B(net126));
 sg13g2_xnor2_1 _1371_ (.Y(_0467_),
    .A(net150),
    .B(net126));
 sg13g2_a21oi_1 _1372_ (.A1(\grad1.acc[3] ),
    .A2(net127),
    .Y(_0468_),
    .B1(_0464_));
 sg13g2_or2_1 _1373_ (.X(_0469_),
    .B(_0468_),
    .A(_0467_));
 sg13g2_nand2_1 _1374_ (.Y(_0470_),
    .A(net212),
    .B(_0469_));
 sg13g2_a21oi_1 _1375_ (.A1(_0467_),
    .A2(_0468_),
    .Y(_0064_),
    .B1(_0470_));
 sg13g2_and2_1 _1376_ (.A(_0466_),
    .B(_0469_),
    .X(_0471_));
 sg13g2_nor2_1 _1377_ (.A(net232),
    .B(net128),
    .Y(_0472_));
 sg13g2_nand2_1 _1378_ (.Y(_0473_),
    .A(net232),
    .B(net128));
 sg13g2_nand2b_1 _1379_ (.Y(_0474_),
    .B(_0473_),
    .A_N(_0472_));
 sg13g2_o21ai_1 _1380_ (.B1(net213),
    .Y(_0475_),
    .A1(_0471_),
    .A2(_0474_));
 sg13g2_a21oi_1 _1381_ (.A1(_0471_),
    .A2(_0474_),
    .Y(_0065_),
    .B1(_0475_));
 sg13g2_xor2_1 _1382_ (.B(net118),
    .A(net227),
    .X(_0476_));
 sg13g2_o21ai_1 _1383_ (.B1(_0473_),
    .Y(_0477_),
    .A1(_0471_),
    .A2(_0472_));
 sg13g2_and2_1 _1384_ (.A(_0476_),
    .B(_0477_),
    .X(_0478_));
 sg13g2_o21ai_1 _1385_ (.B1(net213),
    .Y(_0479_),
    .A1(_0476_),
    .A2(_0477_));
 sg13g2_nor2_1 _1386_ (.A(_0478_),
    .B(_0479_),
    .Y(_0066_));
 sg13g2_xnor2_1 _1387_ (.Y(_0480_),
    .A(\grad1.acc[7] ),
    .B(net123));
 sg13g2_a21oi_1 _1388_ (.A1(net227),
    .A2(net118),
    .Y(_0481_),
    .B1(_0478_));
 sg13g2_nor2_1 _1389_ (.A(_0480_),
    .B(_0481_),
    .Y(_0482_));
 sg13g2_a21oi_1 _1390_ (.A1(_0480_),
    .A2(_0481_),
    .Y(_0483_),
    .B1(_0124_));
 sg13g2_nor2b_1 _1391_ (.A(net228),
    .B_N(_0483_),
    .Y(_0067_));
 sg13g2_a21oi_1 _1392_ (.A1(\grad1.acc[7] ),
    .A2(\grad1.lfsr[7] ),
    .Y(_0484_),
    .B1(_0482_));
 sg13g2_o21ai_1 _1393_ (.B1(net215),
    .Y(_0485_),
    .A1(net112),
    .A2(_0484_));
 sg13g2_a21oi_1 _1394_ (.A1(net112),
    .A2(_0484_),
    .Y(_0068_),
    .B1(_0485_));
 sg13g2_xor2_1 _1395_ (.B(net128),
    .A(net121),
    .X(_0486_));
 sg13g2_xor2_1 _1396_ (.B(\grad1.lfsr[3] ),
    .A(\grad1.lfsr[4] ),
    .X(_0487_));
 sg13g2_xor2_1 _1397_ (.B(net153),
    .A(net115),
    .X(_0488_));
 sg13g2_xnor2_1 _1398_ (.Y(_0489_),
    .A(_0487_),
    .B(_0488_));
 sg13g2_o21ai_1 _1399_ (.B1(net211),
    .Y(_0490_),
    .A1(_0486_),
    .A2(_0489_));
 sg13g2_a21oi_1 _1400_ (.A1(_0486_),
    .A2(net154),
    .Y(_0069_),
    .B1(_0490_));
 sg13g2_and2_1 _1401_ (.A(net214),
    .B(net122),
    .X(_0070_));
 sg13g2_and2_1 _1402_ (.A(net214),
    .B(net119),
    .X(_0071_));
 sg13g2_and2_1 _1403_ (.A(net214),
    .B(net120),
    .X(_0072_));
 sg13g2_and2_1 _1404_ (.A(net212),
    .B(net127),
    .X(_0073_));
 sg13g2_and2_1 _1405_ (.A(net212),
    .B(net126),
    .X(_0074_));
 sg13g2_and2_1 _1406_ (.A(net213),
    .B(net128),
    .X(_0075_));
 sg13g2_and2_1 _1407_ (.A(net213),
    .B(net118),
    .X(_0076_));
 sg13g2_and2_1 _1408_ (.A(net213),
    .B(net123),
    .X(_0077_));
 sg13g2_and2_1 _1409_ (.A(net213),
    .B(net109),
    .X(_0078_));
 sg13g2_and2_1 _1410_ (.A(net213),
    .B(net104),
    .X(_0079_));
 sg13g2_and2_1 _1411_ (.A(net214),
    .B(net103),
    .X(_0080_));
 sg13g2_and2_1 _1412_ (.A(net212),
    .B(net121),
    .X(_0081_));
 sg13g2_and2_1 _1413_ (.A(net211),
    .B(net102),
    .X(_0082_));
 sg13g2_and2_1 _1414_ (.A(net211),
    .B(net111),
    .X(_0083_));
 sg13g2_and2_1 _1415_ (.A(net211),
    .B(net110),
    .X(_0084_));
 sg13g2_and2_1 _1416_ (.A(net211),
    .B(net115),
    .X(_0085_));
 sg13g2_and2_1 _1417_ (.A(net211),
    .B(net114),
    .X(_0086_));
 sg13g2_and2_1 _1418_ (.A(net211),
    .B(net108),
    .X(_0087_));
 sg13g2_and2_1 _1419_ (.A(net211),
    .B(net107),
    .X(_0088_));
 sg13g2_nand2_1 _1420_ (.Y(_0491_),
    .A(\hvsync_gen.vpos[0] ),
    .B(_0171_));
 sg13g2_nand2_1 _1421_ (.Y(_0492_),
    .A(net175),
    .B(_0134_));
 sg13g2_nor2_1 _1422_ (.A(net182),
    .B(net184),
    .Y(_0493_));
 sg13g2_nor4_1 _1423_ (.A(net178),
    .B(net180),
    .C(net182),
    .D(net184),
    .Y(_0494_));
 sg13g2_nor3_1 _1424_ (.A(net176),
    .B(_0190_),
    .C(_0492_),
    .Y(_0495_));
 sg13g2_a21oi_2 _1425_ (.B1(net208),
    .Y(_0496_),
    .A2(_0495_),
    .A1(_0494_));
 sg13g2_nand2_2 _1426_ (.Y(_0497_),
    .A(_0170_),
    .B(_0496_));
 sg13g2_o21ai_1 _1427_ (.B1(_0491_),
    .Y(_0089_),
    .A1(_0105_),
    .A2(_0497_));
 sg13g2_or3_1 _1428_ (.A(_0135_),
    .B(_0189_),
    .C(_0497_),
    .X(_0498_));
 sg13g2_o21ai_1 _1429_ (.B1(_0498_),
    .Y(_0090_),
    .A1(_0120_),
    .A2(net171));
 sg13g2_nand2_1 _1430_ (.Y(_0499_),
    .A(net189),
    .B(_0135_));
 sg13g2_nand2_1 _1431_ (.Y(_0500_),
    .A(_0496_),
    .B(_0499_));
 sg13g2_a21oi_1 _1432_ (.A1(_0135_),
    .A2(net171),
    .Y(_0501_),
    .B1(net189));
 sg13g2_a21oi_1 _1433_ (.A1(net171),
    .A2(_0500_),
    .Y(_0091_),
    .B1(_0501_));
 sg13g2_a21oi_1 _1434_ (.A1(net171),
    .A2(_0500_),
    .Y(_0502_),
    .B1(_0119_));
 sg13g2_nor3_1 _1435_ (.A(net187),
    .B(_0497_),
    .C(_0499_),
    .Y(_0503_));
 sg13g2_or2_1 _1436_ (.X(_0092_),
    .B(_0503_),
    .A(_0502_));
 sg13g2_nand2_2 _1437_ (.Y(_0504_),
    .A(_0134_),
    .B(_0135_));
 sg13g2_nand3_1 _1438_ (.B(_0134_),
    .C(_0135_),
    .A(net184),
    .Y(_0505_));
 sg13g2_a21oi_1 _1439_ (.A1(_0496_),
    .A2(_0505_),
    .Y(_0506_),
    .B1(_0171_));
 sg13g2_nor2_2 _1440_ (.A(_0171_),
    .B(_0504_),
    .Y(_0507_));
 sg13g2_nor2_1 _1441_ (.A(net184),
    .B(_0507_),
    .Y(_0508_));
 sg13g2_nor2_1 _1442_ (.A(_0506_),
    .B(_0508_),
    .Y(_0093_));
 sg13g2_nand3_1 _1443_ (.B(_0496_),
    .C(_0507_),
    .A(_0278_),
    .Y(_0509_));
 sg13g2_o21ai_1 _1444_ (.B1(_0509_),
    .Y(_0094_),
    .A1(_0115_),
    .A2(_0506_));
 sg13g2_or2_1 _1445_ (.X(_0510_),
    .B(_0504_),
    .A(_0295_));
 sg13g2_a21o_1 _1446_ (.A2(_0510_),
    .A1(_0496_),
    .B1(_0171_),
    .X(_0511_));
 sg13g2_o21ai_1 _1447_ (.B1(_0296_),
    .Y(_0512_),
    .A1(net180),
    .A2(_0507_));
 sg13g2_nor2b_1 _1448_ (.A(_0512_),
    .B_N(_0511_),
    .Y(_0095_));
 sg13g2_nor3_1 _1449_ (.A(net178),
    .B(_0497_),
    .C(_0510_),
    .Y(_0513_));
 sg13g2_a21o_1 _1450_ (.A2(_0511_),
    .A1(net178),
    .B1(_0513_),
    .X(_0096_));
 sg13g2_or3_1 _1451_ (.A(_0142_),
    .B(_0295_),
    .C(_0504_),
    .X(_0514_));
 sg13g2_a21oi_1 _1452_ (.A1(_0496_),
    .A2(_0514_),
    .Y(_0515_),
    .B1(_0171_));
 sg13g2_o21ai_1 _1453_ (.B1(_0335_),
    .Y(_0516_),
    .A1(net176),
    .A2(_0507_));
 sg13g2_nor2_1 _1454_ (.A(_0515_),
    .B(_0516_),
    .Y(_0097_));
 sg13g2_nand2_1 _1455_ (.Y(_0517_),
    .A(net175),
    .B(_0171_));
 sg13g2_nor3_1 _1456_ (.A(net157),
    .B(_0334_),
    .C(_0504_),
    .Y(_0518_));
 sg13g2_xnor2_1 _1457_ (.Y(_0519_),
    .A(net175),
    .B(_0518_));
 sg13g2_o21ai_1 _1458_ (.B1(_0517_),
    .Y(_0098_),
    .A1(_0497_),
    .A2(net158));
 sg13g2_and2_1 _1459_ (.A(net177),
    .B(net197),
    .X(_0520_));
 sg13g2_xor2_1 _1460_ (.B(net197),
    .A(net177),
    .X(_0521_));
 sg13g2_nor2_1 _1461_ (.A(net183),
    .B(net202),
    .Y(_0522_));
 sg13g2_and2_1 _1462_ (.A(net184),
    .B(net204),
    .X(_0523_));
 sg13g2_nand2_1 _1463_ (.Y(_0524_),
    .A(net188),
    .B(net206));
 sg13g2_nand2_1 _1464_ (.Y(_0525_),
    .A(net190),
    .B(net207));
 sg13g2_nor2_1 _1465_ (.A(net188),
    .B(net206),
    .Y(_0526_));
 sg13g2_xor2_1 _1466_ (.B(net206),
    .A(net187),
    .X(_0527_));
 sg13g2_o21ai_1 _1467_ (.B1(_0524_),
    .Y(_0528_),
    .A1(_0525_),
    .A2(_0526_));
 sg13g2_or2_1 _1468_ (.X(_0529_),
    .B(net204),
    .A(net185));
 sg13g2_xnor2_1 _1469_ (.Y(_0530_),
    .A(net185),
    .B(net204));
 sg13g2_a21oi_2 _1470_ (.B1(_0523_),
    .Y(_0531_),
    .A2(_0529_),
    .A1(_0528_));
 sg13g2_nor2b_1 _1471_ (.A(_0522_),
    .B_N(_0523_),
    .Y(_0532_));
 sg13g2_xnor2_1 _1472_ (.Y(_0533_),
    .A(net183),
    .B(net202));
 sg13g2_nor2_1 _1473_ (.A(_0530_),
    .B(_0533_),
    .Y(_0534_));
 sg13g2_a221oi_1 _1474_ (.B2(_0534_),
    .C1(_0532_),
    .B1(_0528_),
    .A1(net183),
    .Y(_0535_),
    .A2(net202));
 sg13g2_nor2_1 _1475_ (.A(net179),
    .B(net199),
    .Y(_0536_));
 sg13g2_xor2_1 _1476_ (.B(net199),
    .A(net179),
    .X(_0537_));
 sg13g2_nand2_1 _1477_ (.Y(_0538_),
    .A(net181),
    .B(net201));
 sg13g2_nor2_1 _1478_ (.A(net181),
    .B(net201),
    .Y(_0539_));
 sg13g2_xor2_1 _1479_ (.B(net201),
    .A(net181),
    .X(_0540_));
 sg13g2_nand2_1 _1480_ (.Y(_0541_),
    .A(_0537_),
    .B(_0540_));
 sg13g2_nor2_1 _1481_ (.A(_0536_),
    .B(_0538_),
    .Y(_0542_));
 sg13g2_a21oi_1 _1482_ (.A1(net179),
    .A2(net199),
    .Y(_0543_),
    .B1(_0542_));
 sg13g2_o21ai_1 _1483_ (.B1(_0543_),
    .Y(_0544_),
    .A1(_0535_),
    .A2(_0541_));
 sg13g2_nand2_1 _1484_ (.Y(_0545_),
    .A(\hvsync_gen.hpos[7] ),
    .B(net175));
 sg13g2_nand2b_1 _1485_ (.Y(_0546_),
    .B(_0545_),
    .A_N(_0520_));
 sg13g2_a21o_1 _1486_ (.A2(_0544_),
    .A1(_0521_),
    .B1(_0546_),
    .X(_0547_));
 sg13g2_nand2_2 _1487_ (.Y(_0548_),
    .A(_0113_),
    .B(_0114_));
 sg13g2_and3_1 _1488_ (.X(_0549_),
    .A(\hvsync_gen.hpos[8] ),
    .B(_0547_),
    .C(_0548_));
 sg13g2_nand3_1 _1489_ (.B(_0547_),
    .C(_0548_),
    .A(\hvsync_gen.hpos[8] ),
    .Y(_0550_));
 sg13g2_xnor2_1 _1490_ (.Y(_0551_),
    .A(_0008_),
    .B(_0549_));
 sg13g2_xnor2_1 _1491_ (.Y(_0552_),
    .A(_0008_),
    .B(_0550_));
 sg13g2_a21o_1 _1492_ (.A2(_0548_),
    .A1(_0547_),
    .B1(\hvsync_gen.hpos[8] ),
    .X(_0553_));
 sg13g2_nand2_2 _1493_ (.Y(_0554_),
    .A(_0550_),
    .B(_0553_));
 sg13g2_nand2_1 _1494_ (.Y(_0555_),
    .A(_0545_),
    .B(_0548_));
 sg13g2_a21oi_1 _1495_ (.A1(_0521_),
    .A2(_0544_),
    .Y(_0556_),
    .B1(_0520_));
 sg13g2_xor2_1 _1496_ (.B(_0556_),
    .A(_0555_),
    .X(_0557_));
 sg13g2_xnor2_1 _1497_ (.Y(_0558_),
    .A(_0555_),
    .B(_0556_));
 sg13g2_xor2_1 _1498_ (.B(_0544_),
    .A(_0521_),
    .X(_0559_));
 sg13g2_o21ai_1 _1499_ (.B1(_0538_),
    .Y(_0560_),
    .A1(_0535_),
    .A2(_0539_));
 sg13g2_xnor2_1 _1500_ (.Y(_0561_),
    .A(_0537_),
    .B(_0560_));
 sg13g2_xor2_1 _1501_ (.B(_0560_),
    .A(_0537_),
    .X(_0562_));
 sg13g2_xnor2_1 _1502_ (.Y(_0563_),
    .A(_0535_),
    .B(_0540_));
 sg13g2_xnor2_1 _1503_ (.Y(_0564_),
    .A(_0531_),
    .B(_0533_));
 sg13g2_xor2_1 _1504_ (.B(_0533_),
    .A(_0531_),
    .X(_0565_));
 sg13g2_nand2b_1 _1505_ (.Y(_0566_),
    .B(_0564_),
    .A_N(_0563_));
 sg13g2_and2_1 _1506_ (.A(_0562_),
    .B(_0566_),
    .X(_0567_));
 sg13g2_and3_1 _1507_ (.X(_0568_),
    .A(_0559_),
    .B(_0562_),
    .C(_0566_));
 sg13g2_nor2_1 _1508_ (.A(_0557_),
    .B(_0568_),
    .Y(_0569_));
 sg13g2_a221oi_1 _1509_ (.B2(_0567_),
    .C1(_0557_),
    .B1(_0559_),
    .A1(_0550_),
    .Y(_0570_),
    .A2(_0553_));
 sg13g2_xnor2_1 _1510_ (.Y(_0571_),
    .A(_0551_),
    .B(_0570_));
 sg13g2_nand2_1 _1511_ (.Y(_0572_),
    .A(\counter[3] ),
    .B(_0571_));
 sg13g2_nor2_1 _1512_ (.A(\counter[3] ),
    .B(_0571_),
    .Y(_0573_));
 sg13g2_xor2_1 _1513_ (.B(_0569_),
    .A(_0554_),
    .X(_0574_));
 sg13g2_nor2_1 _1514_ (.A(\counter[2] ),
    .B(_0574_),
    .Y(_0575_));
 sg13g2_xnor2_1 _1515_ (.Y(_0576_),
    .A(_0022_),
    .B(_0574_));
 sg13g2_xnor2_1 _1516_ (.Y(_0577_),
    .A(_0558_),
    .B(_0568_));
 sg13g2_and2_1 _1517_ (.A(\counter[1] ),
    .B(_0577_),
    .X(_0578_));
 sg13g2_or2_1 _1518_ (.X(_0579_),
    .B(_0577_),
    .A(\counter[1] ));
 sg13g2_xnor2_1 _1519_ (.Y(_0580_),
    .A(_0559_),
    .B(_0567_));
 sg13g2_xnor2_1 _1520_ (.Y(_0581_),
    .A(_0528_),
    .B(_0530_));
 sg13g2_xor2_1 _1521_ (.B(net207),
    .A(net190),
    .X(_0582_));
 sg13g2_xnor2_1 _1522_ (.Y(_0583_),
    .A(_0525_),
    .B(_0527_));
 sg13g2_nor4_1 _1523_ (.A(_0563_),
    .B(_0581_),
    .C(_0582_),
    .D(_0583_),
    .Y(_0584_));
 sg13g2_nand4_1 _1524_ (.B(_0562_),
    .C(_0565_),
    .A(_0026_),
    .Y(_0585_),
    .D(_0584_));
 sg13g2_and3_1 _1525_ (.X(_0586_),
    .A(\counter[0] ),
    .B(_0580_),
    .C(_0585_));
 sg13g2_a221oi_1 _1526_ (.B2(_0586_),
    .C1(_0578_),
    .B1(_0579_),
    .A1(\counter[3] ),
    .Y(_0587_),
    .A2(_0571_));
 sg13g2_a221oi_1 _1527_ (.B2(_0587_),
    .C1(_0573_),
    .B1(_0576_),
    .A1(_0572_),
    .Y(_0588_),
    .A2(_0575_));
 sg13g2_nand2_2 _1528_ (.Y(_0589_),
    .A(net194),
    .B(_0549_));
 sg13g2_inv_1 _1529_ (.Y(_0590_),
    .A(_0589_));
 sg13g2_nand3_1 _1530_ (.B(_0570_),
    .C(_0589_),
    .A(_0552_),
    .Y(_0591_));
 sg13g2_and2_1 _1531_ (.A(_0108_),
    .B(_0591_),
    .X(_0592_));
 sg13g2_a21oi_2 _1532_ (.B1(_0589_),
    .Y(_0593_),
    .A2(_0570_),
    .A1(_0552_));
 sg13g2_a21o_1 _1533_ (.A2(_0021_),
    .A1(_0108_),
    .B1(_0593_),
    .X(_0594_));
 sg13g2_o21ai_1 _1534_ (.B1(_0021_),
    .Y(_0595_),
    .A1(_0108_),
    .A2(_0593_));
 sg13g2_mux2_1 _1535_ (.A0(_0595_),
    .A1(_0594_),
    .S(_0592_),
    .X(_0596_));
 sg13g2_nor2_1 _1536_ (.A(\counter[4] ),
    .B(_0593_),
    .Y(_0597_));
 sg13g2_a22oi_1 _1537_ (.Y(_0598_),
    .B1(_0597_),
    .B2(_0592_),
    .A2(_0593_),
    .A1(_0020_));
 sg13g2_o21ai_1 _1538_ (.B1(_0598_),
    .Y(_0599_),
    .A1(_0588_),
    .A2(_0596_));
 sg13g2_a21oi_1 _1539_ (.A1(_0562_),
    .A2(_0563_),
    .Y(_0600_),
    .B1(_0559_));
 sg13g2_and2_1 _1540_ (.A(_0558_),
    .B(_0600_),
    .X(_0601_));
 sg13g2_nor2_1 _1541_ (.A(_0554_),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_o21ai_1 _1542_ (.B1(_0552_),
    .Y(_0603_),
    .A1(_0554_),
    .A2(_0601_));
 sg13g2_nand3_1 _1543_ (.B(net194),
    .C(_0549_),
    .A(_0008_),
    .Y(_0604_));
 sg13g2_nand2_1 _1544_ (.Y(_0605_),
    .A(_0020_),
    .B(_0021_));
 sg13g2_nand2_1 _1545_ (.Y(_0606_),
    .A(_0604_),
    .B(_0605_));
 sg13g2_o21ai_1 _1546_ (.B1(_0020_),
    .Y(_0607_),
    .A1(_0590_),
    .A2(_0603_));
 sg13g2_nand2_1 _1547_ (.Y(_0608_),
    .A(_0021_),
    .B(_0606_));
 sg13g2_mux2_1 _1548_ (.A0(_0606_),
    .A1(_0608_),
    .S(_0607_),
    .X(_0609_));
 sg13g2_xnor2_1 _1549_ (.Y(_0610_),
    .A(_0551_),
    .B(_0602_));
 sg13g2_nor2_1 _1550_ (.A(_0109_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_xnor2_1 _1551_ (.Y(_0612_),
    .A(_0554_),
    .B(_0601_));
 sg13g2_or2_1 _1552_ (.X(_0613_),
    .B(_0612_),
    .A(_0129_));
 sg13g2_nand3_1 _1553_ (.B(_0562_),
    .C(_0563_),
    .A(_0559_),
    .Y(_0614_));
 sg13g2_a221oi_1 _1554_ (.B2(\counter[0] ),
    .C1(_0600_),
    .B1(_0614_),
    .A1(\counter[1] ),
    .Y(_0615_),
    .A2(_0558_));
 sg13g2_nor2_1 _1555_ (.A(\counter[1] ),
    .B(_0558_),
    .Y(_0616_));
 sg13g2_nor3_1 _1556_ (.A(_0601_),
    .B(_0615_),
    .C(_0616_),
    .Y(_0617_));
 sg13g2_a21oi_1 _1557_ (.A1(_0129_),
    .A2(_0612_),
    .Y(_0618_),
    .B1(_0617_));
 sg13g2_nor2_1 _1558_ (.A(\counter[2] ),
    .B(_0612_),
    .Y(_0619_));
 sg13g2_a221oi_1 _1559_ (.B2(_0618_),
    .C1(_0619_),
    .B1(_0613_),
    .A1(_0109_),
    .Y(_0620_),
    .A2(_0610_));
 sg13g2_or3_1 _1560_ (.A(_0609_),
    .B(_0611_),
    .C(_0620_),
    .X(_0621_));
 sg13g2_a21o_1 _1561_ (.A2(_0604_),
    .A1(\counter[4] ),
    .B1(_0607_),
    .X(_0622_));
 sg13g2_and3_1 _1562_ (.X(_0623_),
    .A(_0599_),
    .B(_0621_),
    .C(_0622_));
 sg13g2_nand3_1 _1563_ (.B(_0621_),
    .C(_0622_),
    .A(_0599_),
    .Y(_0624_));
 sg13g2_o21ai_1 _1564_ (.B1(net176),
    .Y(_0625_),
    .A1(net179),
    .A2(net181));
 sg13g2_nand2_1 _1565_ (.Y(_0626_),
    .A(_0114_),
    .B(_0625_));
 sg13g2_nand2_1 _1566_ (.Y(_0627_),
    .A(\hvsync_gen.vpos[1] ),
    .B(_0134_));
 sg13g2_nand3_1 _1567_ (.B(_0138_),
    .C(_0278_),
    .A(_0134_),
    .Y(_0628_));
 sg13g2_nand3_1 _1568_ (.B(_0505_),
    .C(_0628_),
    .A(_0115_),
    .Y(_0629_));
 sg13g2_a21oi_1 _1569_ (.A1(net176),
    .A2(_0629_),
    .Y(_0630_),
    .B1(_0626_));
 sg13g2_nor2_1 _1570_ (.A(net207),
    .B(_0166_),
    .Y(_0631_));
 sg13g2_nand3_1 _1571_ (.B(net201),
    .C(_0631_),
    .A(net202),
    .Y(_0632_));
 sg13g2_a21oi_1 _1572_ (.A1(_0179_),
    .A2(_0632_),
    .Y(_0633_),
    .B1(_0185_));
 sg13g2_nor2b_1 _1573_ (.A(net200),
    .B_N(net198),
    .Y(_0634_));
 sg13g2_nand2b_1 _1574_ (.Y(_0635_),
    .B(_0634_),
    .A_N(_0203_));
 sg13g2_a21oi_1 _1575_ (.A1(_0011_),
    .A2(_0635_),
    .Y(_0636_),
    .B1(_0146_));
 sg13g2_nor2_1 _1576_ (.A(_0205_),
    .B(_0636_),
    .Y(_0637_));
 sg13g2_nor3_1 _1577_ (.A(net193),
    .B(_0633_),
    .C(_0637_),
    .Y(_0638_));
 sg13g2_nor4_2 _1578_ (.A(_0113_),
    .B(net196),
    .C(net193),
    .Y(_0639_),
    .D(_0168_));
 sg13g2_a22oi_1 _1579_ (.Y(_0640_),
    .B1(_0175_),
    .B2(_0639_),
    .A2(_0151_),
    .A1(_0123_));
 sg13g2_nor3_1 _1580_ (.A(net207),
    .B(net202),
    .C(_0166_),
    .Y(_0641_));
 sg13g2_a22oi_1 _1581_ (.Y(_0642_),
    .B1(_0641_),
    .B2(_0639_),
    .A2(_0640_),
    .A1(_0205_));
 sg13g2_a21o_1 _1582_ (.A2(_0150_),
    .A1(net196),
    .B1(\hvsync_gen.hpos[7] ),
    .X(_0643_));
 sg13g2_nor3_1 _1583_ (.A(_0112_),
    .B(net193),
    .C(_0643_),
    .Y(_0644_));
 sg13g2_a21oi_1 _1584_ (.A1(_0493_),
    .A2(_0627_),
    .Y(_0645_),
    .B1(_0143_));
 sg13g2_nor4_1 _1585_ (.A(net175),
    .B(_0204_),
    .C(_0644_),
    .D(_0645_),
    .Y(_0646_));
 sg13g2_a22oi_1 _1586_ (.Y(_0647_),
    .B1(_0642_),
    .B2(_0646_),
    .A2(_0638_),
    .A1(_0630_));
 sg13g2_nand2b_1 _1587_ (.Y(_0648_),
    .B(_0629_),
    .A_N(_0130_));
 sg13g2_a21oi_1 _1588_ (.A1(_0192_),
    .A2(_0648_),
    .Y(_0649_),
    .B1(_0647_));
 sg13g2_nand3_1 _1589_ (.B(net198),
    .C(net196),
    .A(_0113_),
    .Y(_0650_));
 sg13g2_or2_1 _1590_ (.X(_0651_),
    .B(_0650_),
    .A(_0632_));
 sg13g2_nand3_1 _1591_ (.B(_0204_),
    .C(_0651_),
    .A(_0182_),
    .Y(_0652_));
 sg13g2_nor2_1 _1592_ (.A(net201),
    .B(_0650_),
    .Y(_0653_));
 sg13g2_a221oi_1 _1593_ (.B2(_0653_),
    .C1(_0322_),
    .B1(_0167_),
    .A1(_0113_),
    .Y(_0654_),
    .A2(_0011_));
 sg13g2_and3_1 _1594_ (.X(_0655_),
    .A(net203),
    .B(_0631_),
    .C(_0653_));
 sg13g2_nor2_1 _1595_ (.A(net180),
    .B(net184),
    .Y(_0656_));
 sg13g2_a21oi_1 _1596_ (.A1(_0188_),
    .A2(_0656_),
    .Y(_0657_),
    .B1(_0333_));
 sg13g2_nor3_1 _1597_ (.A(net176),
    .B(\hvsync_gen.vpos[9] ),
    .C(net194),
    .Y(_0658_));
 sg13g2_o21ai_1 _1598_ (.B1(_0658_),
    .Y(_0659_),
    .A1(net183),
    .A2(_0130_));
 sg13g2_nor4_1 _1599_ (.A(_0654_),
    .B(_0655_),
    .C(_0657_),
    .D(_0659_),
    .Y(_0660_));
 sg13g2_nand3b_1 _1600_ (.B(_0634_),
    .C(_0641_),
    .Y(_0661_),
    .A_N(_0169_));
 sg13g2_nand2b_1 _1601_ (.Y(_0662_),
    .B(\hvsync_gen.vpos[6] ),
    .A_N(net178));
 sg13g2_nor4_1 _1602_ (.A(net182),
    .B(net184),
    .C(_0141_),
    .D(_0662_),
    .Y(_0663_));
 sg13g2_nand4_1 _1603_ (.B(net187),
    .C(_0189_),
    .A(_0118_),
    .Y(_0664_),
    .D(_0663_));
 sg13g2_nand4_1 _1604_ (.B(_0322_),
    .C(_0661_),
    .A(_0123_),
    .Y(_0665_),
    .D(_0664_));
 sg13g2_nand2_1 _1605_ (.Y(_0666_),
    .A(_0119_),
    .B(_0663_));
 sg13g2_nand2_1 _1606_ (.Y(_0667_),
    .A(_0626_),
    .B(_0666_));
 sg13g2_nand2b_1 _1607_ (.Y(_0668_),
    .B(net195),
    .A_N(_0011_));
 sg13g2_a21oi_1 _1608_ (.A1(_0175_),
    .A2(_0634_),
    .Y(_0669_),
    .B1(_0668_));
 sg13g2_nor3_1 _1609_ (.A(_0637_),
    .B(_0665_),
    .C(_0669_),
    .Y(_0670_));
 sg13g2_a22oi_1 _1610_ (.Y(_0671_),
    .B1(_0667_),
    .B2(_0670_),
    .A2(_0660_),
    .A1(_0652_));
 sg13g2_nor2_1 _1611_ (.A(_0132_),
    .B(_0662_),
    .Y(_0672_));
 sg13g2_a21oi_1 _1612_ (.A1(net181),
    .A2(_0116_),
    .Y(_0673_),
    .B1(net179));
 sg13g2_a21oi_1 _1613_ (.A1(_0188_),
    .A2(_0672_),
    .Y(_0674_),
    .B1(_0673_));
 sg13g2_nand4_1 _1614_ (.B(_0119_),
    .C(_0189_),
    .A(net189),
    .Y(_0675_),
    .D(_0672_));
 sg13g2_nor2b_1 _1615_ (.A(_0674_),
    .B_N(_0192_),
    .Y(_0676_));
 sg13g2_a21oi_1 _1616_ (.A1(_0675_),
    .A2(_0676_),
    .Y(_0677_),
    .B1(_0671_));
 sg13g2_nand2b_1 _1617_ (.Y(_0678_),
    .B(\r[6] ),
    .A_N(\r[7] ));
 sg13g2_or3_1 _1618_ (.A(\r[4] ),
    .B(\r[3] ),
    .C(_0678_),
    .X(_0679_));
 sg13g2_nor2b_1 _1619_ (.A(_0222_),
    .B_N(\r[2] ),
    .Y(_0680_));
 sg13g2_nor2_1 _1620_ (.A(_0679_),
    .B(_0680_),
    .Y(_0681_));
 sg13g2_nor2_1 _1621_ (.A(net192),
    .B(_0678_),
    .Y(_0682_));
 sg13g2_nand3_1 _1622_ (.B(\r[9] ),
    .C(\r[8] ),
    .A(\r[12] ),
    .Y(_0683_));
 sg13g2_nor2_1 _1623_ (.A(\r[7] ),
    .B(\r[6] ),
    .Y(_0684_));
 sg13g2_and2_1 _1624_ (.A(\r[11] ),
    .B(\r[10] ),
    .X(_0685_));
 sg13g2_nand2b_1 _1625_ (.Y(_0686_),
    .B(_0685_),
    .A_N(_0684_));
 sg13g2_nor4_1 _1626_ (.A(_0681_),
    .B(_0682_),
    .C(_0683_),
    .D(_0686_),
    .Y(_0687_));
 sg13g2_nand2_1 _1627_ (.Y(_0688_),
    .A(\r[2] ),
    .B(_0222_));
 sg13g2_nor3_1 _1628_ (.A(net192),
    .B(_0679_),
    .C(_0688_),
    .Y(_0689_));
 sg13g2_nand2_1 _1629_ (.Y(_0690_),
    .A(\r[12] ),
    .B(_0685_));
 sg13g2_nor2_1 _1630_ (.A(\r[13] ),
    .B(\r[9] ),
    .Y(_0691_));
 sg13g2_nand4_1 _1631_ (.B(\r[14] ),
    .C(\r[8] ),
    .A(\r[15] ),
    .Y(_0692_),
    .D(_0691_));
 sg13g2_nor2_1 _1632_ (.A(_0690_),
    .B(_0692_),
    .Y(_0693_));
 sg13g2_a22oi_1 _1633_ (.Y(_0694_),
    .B1(_0689_),
    .B2(_0693_),
    .A2(_0107_),
    .A1(_0106_));
 sg13g2_o21ai_1 _1634_ (.B1(\r[15] ),
    .Y(_0695_),
    .A1(_0687_),
    .A2(_0694_));
 sg13g2_and2_1 _1635_ (.A(_0010_),
    .B(_0695_),
    .X(_0696_));
 sg13g2_nor2_1 _1636_ (.A(net180),
    .B(_0118_),
    .Y(_0697_));
 sg13g2_a221oi_1 _1637_ (.B2(_0697_),
    .C1(net187),
    .B1(_0138_),
    .A1(net189),
    .Y(_0698_),
    .A2(_0135_));
 sg13g2_or3_1 _1638_ (.A(_0117_),
    .B(_0333_),
    .C(_0698_),
    .X(_0699_));
 sg13g2_nand4_1 _1639_ (.B(_0192_),
    .C(_0643_),
    .A(_0130_),
    .Y(_0700_),
    .D(_0657_));
 sg13g2_nor2b_1 _1640_ (.A(_0700_),
    .B_N(_0699_),
    .Y(_0701_));
 sg13g2_nor2_1 _1641_ (.A(\r[9] ),
    .B(\r[8] ),
    .Y(_0702_));
 sg13g2_o21ai_1 _1642_ (.B1(_0107_),
    .Y(_0703_),
    .A1(_0690_),
    .A2(_0702_));
 sg13g2_nor3_1 _1643_ (.A(net192),
    .B(_0679_),
    .C(_0680_),
    .Y(_0704_));
 sg13g2_o21ai_1 _1644_ (.B1(_0693_),
    .Y(_0705_),
    .A1(_0684_),
    .A2(_0704_));
 sg13g2_nand4_1 _1645_ (.B(\r[14] ),
    .C(_0703_),
    .A(\r[15] ),
    .Y(_0706_),
    .D(_0705_));
 sg13g2_a21oi_1 _1646_ (.A1(_0637_),
    .A2(_0701_),
    .Y(_0707_),
    .B1(\r[16] ));
 sg13g2_nand2_1 _1647_ (.Y(_0708_),
    .A(_0706_),
    .B(_0707_));
 sg13g2_a21oi_1 _1648_ (.A1(net201),
    .A2(net199),
    .Y(_0709_),
    .B1(net197));
 sg13g2_nand3_1 _1649_ (.B(net205),
    .C(net199),
    .A(net203),
    .Y(_0710_));
 sg13g2_a21oi_1 _1650_ (.A1(_0709_),
    .A2(_0710_),
    .Y(_0711_),
    .B1(_0113_));
 sg13g2_nand3_1 _1651_ (.B(_0123_),
    .C(_0193_),
    .A(net195),
    .Y(_0712_));
 sg13g2_nor4_1 _1652_ (.A(_0630_),
    .B(_0642_),
    .C(_0711_),
    .D(_0712_),
    .Y(_0713_));
 sg13g2_nor3_1 _1653_ (.A(_0696_),
    .B(_0708_),
    .C(_0713_),
    .Y(_0714_));
 sg13g2_or3_2 _1654_ (.A(_0649_),
    .B(_0677_),
    .C(_0714_),
    .X(_0715_));
 sg13g2_nand2_1 _1655_ (.Y(_0716_),
    .A(_0563_),
    .B(_0565_));
 sg13g2_nor2_1 _1656_ (.A(_0561_),
    .B(_0716_),
    .Y(_0717_));
 sg13g2_nor2_1 _1657_ (.A(_0564_),
    .B(_0614_),
    .Y(_0718_));
 sg13g2_nor2_1 _1658_ (.A(_0557_),
    .B(_0718_),
    .Y(_0719_));
 sg13g2_nand2_1 _1659_ (.Y(_0720_),
    .A(_0554_),
    .B(_0719_));
 sg13g2_xor2_1 _1660_ (.B(_0719_),
    .A(_0554_),
    .X(_0721_));
 sg13g2_nand2_1 _1661_ (.Y(_0722_),
    .A(\grad1.acc[8] ),
    .B(_0721_));
 sg13g2_xnor2_1 _1662_ (.Y(_0723_),
    .A(_0561_),
    .B(_0716_));
 sg13g2_and2_1 _1663_ (.A(_0566_),
    .B(_0716_),
    .X(_0724_));
 sg13g2_or2_1 _1664_ (.X(_0725_),
    .B(_0581_),
    .A(_0018_));
 sg13g2_and2_1 _1665_ (.A(_0018_),
    .B(_0581_),
    .X(_0726_));
 sg13g2_nor2_1 _1666_ (.A(_0019_),
    .B(_0583_),
    .Y(_0727_));
 sg13g2_nand2_1 _1667_ (.Y(_0728_),
    .A(_0128_),
    .B(_0582_));
 sg13g2_xor2_1 _1668_ (.B(_0583_),
    .A(_0019_),
    .X(_0729_));
 sg13g2_a21oi_1 _1669_ (.A1(_0728_),
    .A2(_0729_),
    .Y(_0730_),
    .B1(_0727_));
 sg13g2_a21oi_1 _1670_ (.A1(_0725_),
    .A2(_0730_),
    .Y(_0731_),
    .B1(_0726_));
 sg13g2_nor2_1 _1671_ (.A(_0017_),
    .B(_0724_),
    .Y(_0732_));
 sg13g2_o21ai_1 _1672_ (.B1(_0731_),
    .Y(_0733_),
    .A1(\grad1.acc[3] ),
    .A2(_0565_));
 sg13g2_a21oi_1 _1673_ (.A1(\grad1.acc[3] ),
    .A2(_0565_),
    .Y(_0734_),
    .B1(_0732_));
 sg13g2_a22oi_1 _1674_ (.Y(_0735_),
    .B1(_0733_),
    .B2(_0734_),
    .A2(_0724_),
    .A1(_0017_));
 sg13g2_xnor2_1 _1675_ (.Y(_0736_),
    .A(_0016_),
    .B(_0723_));
 sg13g2_a22oi_1 _1676_ (.Y(_0737_),
    .B1(_0735_),
    .B2(_0736_),
    .A2(_0723_),
    .A1(\grad1.acc[5] ));
 sg13g2_xnor2_1 _1677_ (.Y(_0738_),
    .A(_0559_),
    .B(_0717_));
 sg13g2_xor2_1 _1678_ (.B(_0738_),
    .A(_0015_),
    .X(_0739_));
 sg13g2_nor2_1 _1679_ (.A(_0737_),
    .B(_0739_),
    .Y(_0740_));
 sg13g2_xnor2_1 _1680_ (.Y(_0741_),
    .A(_0558_),
    .B(_0718_));
 sg13g2_a221oi_1 _1681_ (.B2(\grad1.acc[7] ),
    .C1(_0740_),
    .B1(_0741_),
    .A1(\grad1.acc[6] ),
    .Y(_0742_),
    .A2(_0738_));
 sg13g2_xnor2_1 _1682_ (.Y(_0743_),
    .A(_0014_),
    .B(_0721_));
 sg13g2_o21ai_1 _1683_ (.B1(_0743_),
    .Y(_0744_),
    .A1(\grad1.acc[7] ),
    .A2(_0741_));
 sg13g2_o21ai_1 _1684_ (.B1(_0722_),
    .Y(_0745_),
    .A1(_0742_),
    .A2(_0744_));
 sg13g2_xnor2_1 _1685_ (.Y(_0746_),
    .A(_0552_),
    .B(_0720_));
 sg13g2_nand3_1 _1686_ (.B(_0745_),
    .C(_0746_),
    .A(_0589_),
    .Y(_0747_));
 sg13g2_nand2_1 _1687_ (.Y(_0748_),
    .A(_0715_),
    .B(_0747_));
 sg13g2_nor2_1 _1688_ (.A(_0623_),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_nor2_1 _1689_ (.A(_0026_),
    .B(_0562_),
    .Y(_0750_));
 sg13g2_xnor2_1 _1690_ (.Y(_0751_),
    .A(\counter[1] ),
    .B(_0559_));
 sg13g2_nor2b_1 _1691_ (.A(_0750_),
    .B_N(_0751_),
    .Y(_0752_));
 sg13g2_xnor2_1 _1692_ (.Y(_0753_),
    .A(_0750_),
    .B(_0751_));
 sg13g2_xnor2_1 _1693_ (.Y(_0754_),
    .A(_0111_),
    .B(_0561_));
 sg13g2_nor2_1 _1694_ (.A(_0016_),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_a22oi_1 _1695_ (.Y(_0756_),
    .B1(_0565_),
    .B2(_0127_),
    .A2(_0563_),
    .A1(_0017_));
 sg13g2_o21ai_1 _1696_ (.B1(_0756_),
    .Y(_0757_),
    .A1(_0017_),
    .A2(_0563_));
 sg13g2_nor2_1 _1697_ (.A(_0127_),
    .B(_0565_),
    .Y(_0758_));
 sg13g2_nor2_1 _1698_ (.A(_0731_),
    .B(_0758_),
    .Y(_0759_));
 sg13g2_or2_1 _1699_ (.X(_0760_),
    .B(_0759_),
    .A(_0757_));
 sg13g2_nand2b_1 _1700_ (.Y(_0761_),
    .B(\grad1.acc[4] ),
    .A_N(_0563_));
 sg13g2_o21ai_1 _1701_ (.B1(_0725_),
    .Y(_0762_),
    .A1(_0128_),
    .A2(_0582_));
 sg13g2_nor4_1 _1702_ (.A(_0726_),
    .B(_0757_),
    .C(_0758_),
    .D(_0762_),
    .Y(_0763_));
 sg13g2_nand3_1 _1703_ (.B(_0729_),
    .C(_0763_),
    .A(_0728_),
    .Y(_0764_));
 sg13g2_a22oi_1 _1704_ (.Y(_0765_),
    .B1(_0760_),
    .B2(_0761_),
    .A2(_0754_),
    .A1(_0016_));
 sg13g2_a21oi_1 _1705_ (.A1(_0764_),
    .A2(_0765_),
    .Y(_0766_),
    .B1(_0755_));
 sg13g2_a21o_1 _1706_ (.A2(_0753_),
    .A1(_0015_),
    .B1(_0766_),
    .X(_0767_));
 sg13g2_or2_1 _1707_ (.X(_0768_),
    .B(_0753_),
    .A(_0015_));
 sg13g2_and3_1 _1708_ (.X(_0769_),
    .A(_0715_),
    .B(_0767_),
    .C(_0768_));
 sg13g2_and2_1 _1709_ (.A(_0624_),
    .B(_0769_),
    .X(_0770_));
 sg13g2_a21oi_1 _1710_ (.A1(_0110_),
    .A2(_0559_),
    .Y(_0771_),
    .B1(_0752_));
 sg13g2_xnor2_1 _1711_ (.Y(_0772_),
    .A(_0022_),
    .B(_0557_));
 sg13g2_xnor2_1 _1712_ (.Y(_0773_),
    .A(_0771_),
    .B(_0772_));
 sg13g2_inv_1 _1713_ (.Y(_0774_),
    .A(_0773_));
 sg13g2_nand3_1 _1714_ (.B(_0769_),
    .C(_0774_),
    .A(_0624_),
    .Y(_0775_));
 sg13g2_nor2_1 _1715_ (.A(\counter[3] ),
    .B(_0554_),
    .Y(_0776_));
 sg13g2_xnor2_1 _1716_ (.Y(_0777_),
    .A(_0109_),
    .B(_0554_));
 sg13g2_nand2b_1 _1717_ (.Y(_0778_),
    .B(_0557_),
    .A_N(\counter[2] ));
 sg13g2_o21ai_1 _1718_ (.B1(_0778_),
    .Y(_0779_),
    .A1(_0771_),
    .A2(_0772_));
 sg13g2_xor2_1 _1719_ (.B(_0779_),
    .A(_0777_),
    .X(_0780_));
 sg13g2_inv_1 _1720_ (.Y(_0781_),
    .A(_0780_));
 sg13g2_nand4_1 _1721_ (.B(_0769_),
    .C(_0774_),
    .A(_0624_),
    .Y(_0782_),
    .D(_0780_));
 sg13g2_a21oi_2 _1722_ (.B1(_0776_),
    .Y(_0783_),
    .A2(_0779_),
    .A1(_0777_));
 sg13g2_xnor2_1 _1723_ (.Y(_0784_),
    .A(_0021_),
    .B(_0551_));
 sg13g2_xnor2_1 _1724_ (.Y(_0785_),
    .A(_0783_),
    .B(_0784_));
 sg13g2_nand2b_1 _1725_ (.Y(_0786_),
    .B(_0551_),
    .A_N(\counter[4] ));
 sg13g2_o21ai_1 _1726_ (.B1(_0786_),
    .Y(_0787_),
    .A1(_0783_),
    .A2(_0784_));
 sg13g2_xor2_1 _1727_ (.B(_0589_),
    .A(_0020_),
    .X(_0788_));
 sg13g2_xnor2_1 _1728_ (.Y(_0789_),
    .A(_0787_),
    .B(_0788_));
 sg13g2_o21ai_1 _1729_ (.B1(_0789_),
    .Y(_0790_),
    .A1(_0782_),
    .A2(_0785_));
 sg13g2_and2_1 _1730_ (.A(_0782_),
    .B(_0785_),
    .X(_0791_));
 sg13g2_nor2_1 _1731_ (.A(_0790_),
    .B(_0791_),
    .Y(_0792_));
 sg13g2_xnor2_1 _1732_ (.Y(_0793_),
    .A(_0775_),
    .B(_0780_));
 sg13g2_xnor2_1 _1733_ (.Y(_0794_),
    .A(_0775_),
    .B(_0781_));
 sg13g2_xnor2_1 _1734_ (.Y(_0795_),
    .A(_0770_),
    .B(_0773_));
 sg13g2_xnor2_1 _1735_ (.Y(_0796_),
    .A(_0770_),
    .B(_0774_));
 sg13g2_o21ai_1 _1736_ (.B1(_0792_),
    .Y(_0797_),
    .A1(_0793_),
    .A2(_0795_));
 sg13g2_a22oi_1 _1737_ (.Y(_0798_),
    .B1(\grad1.acc[0] ),
    .B2(_0121_),
    .A2(\grad1.acc[1] ),
    .A1(_0120_));
 sg13g2_nand2b_1 _1738_ (.Y(_0799_),
    .B(net190),
    .A_N(\grad1.acc[2] ));
 sg13g2_o21ai_1 _1739_ (.B1(_0799_),
    .Y(_0800_),
    .A1(_0120_),
    .A2(\grad1.acc[1] ));
 sg13g2_nor2_1 _1740_ (.A(_0798_),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_a221oi_1 _1741_ (.B2(_0118_),
    .C1(_0801_),
    .B1(\grad1.acc[2] ),
    .A1(_0119_),
    .Y(_0802_),
    .A2(\grad1.acc[3] ));
 sg13g2_a221oi_1 _1742_ (.B2(net187),
    .C1(_0802_),
    .B1(_0127_),
    .A1(net185),
    .Y(_0803_),
    .A2(_0126_));
 sg13g2_a221oi_1 _1743_ (.B2(_0117_),
    .C1(_0803_),
    .B1(\grad1.acc[4] ),
    .A1(_0115_),
    .Y(_0804_),
    .A2(\grad1.acc[5] ));
 sg13g2_a21oi_1 _1744_ (.A1(net181),
    .A2(_0125_),
    .Y(_0805_),
    .B1(_0804_));
 sg13g2_o21ai_1 _1745_ (.B1(_0805_),
    .Y(_0806_),
    .A1(_0115_),
    .A2(\grad1.acc[5] ));
 sg13g2_nor2b_1 _1746_ (.A(_0715_),
    .B_N(_0806_),
    .Y(_0807_));
 sg13g2_o21ai_1 _1747_ (.B1(_0807_),
    .Y(_0808_),
    .A1(net181),
    .A2(_0125_));
 sg13g2_nor2_1 _1748_ (.A(_0142_),
    .B(_0808_),
    .Y(_0809_));
 sg13g2_o21ai_1 _1749_ (.B1(_0195_),
    .Y(_0810_),
    .A1(_0142_),
    .A2(_0808_));
 sg13g2_a21oi_1 _1750_ (.A1(_0749_),
    .A2(_0797_),
    .Y(_0099_),
    .B1(_0810_));
 sg13g2_or2_1 _1751_ (.X(_0811_),
    .B(net179),
    .A(net177));
 sg13g2_a21oi_1 _1752_ (.A1(_0142_),
    .A2(_0811_),
    .Y(_0812_),
    .B1(_0808_));
 sg13g2_a21o_1 _1753_ (.A2(_0808_),
    .A1(net157),
    .B1(_0812_),
    .X(_0813_));
 sg13g2_xor2_1 _1754_ (.B(_0808_),
    .A(_0012_),
    .X(_0814_));
 sg13g2_inv_1 _1755_ (.Y(_0815_),
    .A(_0814_));
 sg13g2_nand2b_1 _1756_ (.Y(_0816_),
    .B(_0814_),
    .A_N(_0813_));
 sg13g2_nor2_1 _1757_ (.A(_0715_),
    .B(_0809_),
    .Y(_0817_));
 sg13g2_nand2_1 _1758_ (.Y(_0818_),
    .A(_0816_),
    .B(_0817_));
 sg13g2_nor4_1 _1759_ (.A(_0781_),
    .B(_0790_),
    .C(_0791_),
    .D(_0796_),
    .Y(_0819_));
 sg13g2_nor2_1 _1760_ (.A(_0623_),
    .B(_0819_),
    .Y(_0820_));
 sg13g2_o21ai_1 _1761_ (.B1(_0715_),
    .Y(_0821_),
    .A1(_0623_),
    .A2(_0819_));
 sg13g2_a21oi_1 _1762_ (.A1(_0818_),
    .A2(_0821_),
    .Y(_0100_),
    .B1(_0196_));
 sg13g2_nor2_1 _1763_ (.A(_0196_),
    .B(_0749_),
    .Y(_0101_));
 sg13g2_a21oi_1 _1764_ (.A1(_0782_),
    .A2(_0785_),
    .Y(_0822_),
    .B1(_0789_));
 sg13g2_nor3_1 _1765_ (.A(_0793_),
    .B(_0795_),
    .C(_0822_),
    .Y(_0823_));
 sg13g2_nand2b_1 _1766_ (.Y(_0824_),
    .B(_0715_),
    .A_N(_0747_));
 sg13g2_a21oi_1 _1767_ (.A1(_0790_),
    .A2(_0823_),
    .Y(_0825_),
    .B1(_0824_));
 sg13g2_o21ai_1 _1768_ (.B1(_0195_),
    .Y(_0826_),
    .A1(_0715_),
    .A2(_0816_));
 sg13g2_a21oi_1 _1769_ (.A1(_0820_),
    .A2(_0825_),
    .Y(_0102_),
    .B1(_0826_));
 sg13g2_nor4_1 _1770_ (.A(_0790_),
    .B(_0791_),
    .C(_0794_),
    .D(_0795_),
    .Y(_0827_));
 sg13g2_o21ai_1 _1771_ (.B1(_0715_),
    .Y(_0828_),
    .A1(_0623_),
    .A2(_0827_));
 sg13g2_o21ai_1 _1772_ (.B1(_0817_),
    .Y(_0829_),
    .A1(_0813_),
    .A2(_0814_));
 sg13g2_a21oi_1 _1773_ (.A1(_0828_),
    .A2(_0829_),
    .Y(_0103_),
    .B1(net170));
 sg13g2_nand3_1 _1774_ (.B(_0815_),
    .C(_0817_),
    .A(_0813_),
    .Y(_0830_));
 sg13g2_a21oi_1 _1775_ (.A1(_0748_),
    .A2(_0830_),
    .Y(_0104_),
    .B1(net170));
 sg13g2_dfrbp_1 _1776_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net81),
    .D(net101),
    .Q_N(_0885_),
    .Q(vsync_prev));
 sg13g2_dfrbp_1 _1777_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net18),
    .D(net99),
    .Q_N(_0884_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _1778_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net74),
    .D(net125),
    .Q_N(_0026_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net72),
    .D(_0028_),
    .Q_N(_0883_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _1780_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net70),
    .D(net130),
    .Q_N(_0022_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _1781_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net68),
    .D(net143),
    .Q_N(_0882_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net66),
    .D(_0031_),
    .Q_N(_0021_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net64),
    .D(net117),
    .Q_N(_0020_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net62),
    .D(_0033_),
    .Q_N(_0025_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net61),
    .D(net221),
    .Q_N(_0881_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _1786_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net60),
    .D(net161),
    .Q_N(_0880_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _1787_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net59),
    .D(_0036_),
    .Q_N(_0879_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _1788_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net58),
    .D(_0037_),
    .Q_N(_0878_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _1789_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net57),
    .D(_0038_),
    .Q_N(_0011_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _1790_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net56),
    .D(_0039_),
    .Q_N(_0877_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _1791_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net55),
    .D(_0040_),
    .Q_N(_0876_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _1792_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net54),
    .D(_0041_),
    .Q_N(_0875_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _1793_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net53),
    .D(_0042_),
    .Q_N(_0008_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _1794_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net52),
    .D(_0043_),
    .Q_N(_0874_),
    .Q(\r[0] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net50),
    .D(net146),
    .Q_N(_0873_),
    .Q(\r[1] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net48),
    .D(_0045_),
    .Q_N(_0872_),
    .Q(\r[2] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net46),
    .D(_0046_),
    .Q_N(_0871_),
    .Q(\r[3] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net44),
    .D(_0047_),
    .Q_N(_0870_),
    .Q(\r[4] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net42),
    .D(_0048_),
    .Q_N(_0869_),
    .Q(\r[5] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net40),
    .D(_0049_),
    .Q_N(_0868_),
    .Q(\r[6] ));
 sg13g2_dfrbp_1 _1801_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net38),
    .D(_0050_),
    .Q_N(_0867_),
    .Q(\r[7] ));
 sg13g2_dfrbp_1 _1802_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net36),
    .D(_0051_),
    .Q_N(_0023_),
    .Q(\r[8] ));
 sg13g2_dfrbp_1 _1803_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net34),
    .D(_0052_),
    .Q_N(_0866_),
    .Q(\r[9] ));
 sg13g2_dfrbp_1 _1804_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net32),
    .D(_0053_),
    .Q_N(_0002_),
    .Q(\r[10] ));
 sg13g2_dfrbp_1 _1805_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net30),
    .D(_0054_),
    .Q_N(_0003_),
    .Q(\r[11] ));
 sg13g2_dfrbp_1 _1806_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net28),
    .D(_0055_),
    .Q_N(_0004_),
    .Q(\r[12] ));
 sg13g2_dfrbp_1 _1807_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net26),
    .D(net235),
    .Q_N(_0005_),
    .Q(\r[13] ));
 sg13g2_dfrbp_1 _1808_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net24),
    .D(_0057_),
    .Q_N(_0006_),
    .Q(\r[14] ));
 sg13g2_dfrbp_1 _1809_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net22),
    .D(_0058_),
    .Q_N(_0007_),
    .Q(\r[15] ));
 sg13g2_dfrbp_1 _1810_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net20),
    .D(net141),
    .Q_N(_0010_),
    .Q(\r[16] ));
 sg13g2_dfrbp_1 _1811_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net17),
    .D(_0060_),
    .Q_N(_0865_),
    .Q(\grad1.acc[0] ));
 sg13g2_dfrbp_1 _1812_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net98),
    .D(_0061_),
    .Q_N(_0019_),
    .Q(\grad1.acc[1] ));
 sg13g2_dfrbp_1 _1813_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net97),
    .D(_0062_),
    .Q_N(_0018_),
    .Q(\grad1.acc[2] ));
 sg13g2_dfrbp_1 _1814_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net96),
    .D(net148),
    .Q_N(_0864_),
    .Q(\grad1.acc[3] ));
 sg13g2_dfrbp_1 _1815_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net95),
    .D(net151),
    .Q_N(_0017_),
    .Q(\grad1.acc[4] ));
 sg13g2_dfrbp_1 _1816_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net94),
    .D(_0065_),
    .Q_N(_0016_),
    .Q(\grad1.acc[5] ));
 sg13g2_dfrbp_1 _1817_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net93),
    .D(_0066_),
    .Q_N(_0015_),
    .Q(\grad1.acc[6] ));
 sg13g2_dfrbp_1 _1818_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net91),
    .D(net229),
    .Q_N(_0863_),
    .Q(\grad1.acc[7] ));
 sg13g2_dfrbp_1 _1819_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net90),
    .D(net113),
    .Q_N(_0014_),
    .Q(\grad1.acc[8] ));
 sg13g2_dfrbp_1 _1820_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net89),
    .D(_0069_),
    .Q_N(_0862_),
    .Q(\grad1.lfsr[0] ));
 sg13g2_dfrbp_1 _1821_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net88),
    .D(_0070_),
    .Q_N(_0861_),
    .Q(\grad1.lfsr[1] ));
 sg13g2_dfrbp_1 _1822_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net87),
    .D(_0071_),
    .Q_N(_0860_),
    .Q(\grad1.lfsr[2] ));
 sg13g2_dfrbp_1 _1823_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net86),
    .D(_0072_),
    .Q_N(_0859_),
    .Q(\grad1.lfsr[3] ));
 sg13g2_dfrbp_1 _1824_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net85),
    .D(_0073_),
    .Q_N(_0858_),
    .Q(\grad1.lfsr[4] ));
 sg13g2_dfrbp_1 _1825_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net84),
    .D(_0074_),
    .Q_N(_0857_),
    .Q(\grad1.lfsr[5] ));
 sg13g2_dfrbp_1 _1826_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net83),
    .D(_0075_),
    .Q_N(_0856_),
    .Q(\grad1.lfsr[6] ));
 sg13g2_dfrbp_1 _1827_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net82),
    .D(_0076_),
    .Q_N(_0855_),
    .Q(\grad1.lfsr[7] ));
 sg13g2_dfrbp_1 _1828_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net80),
    .D(_0077_),
    .Q_N(_0854_),
    .Q(\grad1.lfsr[8] ));
 sg13g2_dfrbp_1 _1829_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net79),
    .D(_0078_),
    .Q_N(_0853_),
    .Q(\grad1.lfsr[9] ));
 sg13g2_dfrbp_1 _1830_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net78),
    .D(_0079_),
    .Q_N(_0852_),
    .Q(\grad1.lfsr[10] ));
 sg13g2_dfrbp_1 _1831_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net77),
    .D(_0080_),
    .Q_N(_0851_),
    .Q(\grad1.lfsr[11] ));
 sg13g2_dfrbp_1 _1832_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net76),
    .D(_0081_),
    .Q_N(_0850_),
    .Q(\grad1.lfsr[12] ));
 sg13g2_dfrbp_1 _1833_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net75),
    .D(_0082_),
    .Q_N(_0849_),
    .Q(\grad1.lfsr[13] ));
 sg13g2_dfrbp_1 _1834_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net73),
    .D(_0083_),
    .Q_N(_0848_),
    .Q(\grad1.lfsr[14] ));
 sg13g2_dfrbp_1 _1835_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net71),
    .D(_0084_),
    .Q_N(_0847_),
    .Q(\grad1.lfsr[15] ));
 sg13g2_dfrbp_1 _1836_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net69),
    .D(_0085_),
    .Q_N(_0846_),
    .Q(\grad1.lfsr[16] ));
 sg13g2_dfrbp_1 _1837_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net67),
    .D(_0086_),
    .Q_N(_0845_),
    .Q(\grad1.lfsr[17] ));
 sg13g2_dfrbp_1 _1838_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net65),
    .D(_0087_),
    .Q_N(_0844_),
    .Q(\grad1.lfsr[18] ));
 sg13g2_dfrbp_1 _1839_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net92),
    .D(_0088_),
    .Q_N(_0886_),
    .Q(\grad1.lfsr[19] ));
 sg13g2_dfrbp_1 _1840_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net63),
    .D(_0000_),
    .Q_N(_0843_),
    .Q(hsync));
 sg13g2_dfrbp_1 _1841_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net51),
    .D(net106),
    .Q_N(_0024_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _1842_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net47),
    .D(_0090_),
    .Q_N(_0842_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _1843_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net43),
    .D(_0091_),
    .Q_N(_0841_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _1844_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net39),
    .D(_0092_),
    .Q_N(_0840_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _1845_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net35),
    .D(_0093_),
    .Q_N(_0839_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _1846_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net31),
    .D(_0094_),
    .Q_N(_0009_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _1847_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net27),
    .D(_0095_),
    .Q_N(_0838_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _1848_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net23),
    .D(_0096_),
    .Q_N(_0012_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _1849_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net19),
    .D(_0097_),
    .Q_N(_0013_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _1850_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net41),
    .D(net159),
    .Q_N(_0887_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _1851_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net45),
    .D(net132),
    .Q_N(_0837_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _1852_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net37),
    .D(_0099_),
    .Q_N(_0836_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1853_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net33),
    .D(_0100_),
    .Q_N(_0835_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1854_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net29),
    .D(_0101_),
    .Q_N(_0834_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1855_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net25),
    .D(_0102_),
    .Q_N(_0833_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1856_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net21),
    .D(_0103_),
    .Q_N(_0832_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1857_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net49),
    .D(_0104_),
    .Q_N(_0831_),
    .Q(uo_out[6]));
 sg13g2_tiehi _1777__18 (.L_HI(net18));
 sg13g2_tiehi _1849__19 (.L_HI(net19));
 sg13g2_tiehi _1810__20 (.L_HI(net20));
 sg13g2_tiehi _1856__21 (.L_HI(net21));
 sg13g2_tiehi _1809__22 (.L_HI(net22));
 sg13g2_tiehi _1848__23 (.L_HI(net23));
 sg13g2_tiehi _1808__24 (.L_HI(net24));
 sg13g2_tiehi _1855__25 (.L_HI(net25));
 sg13g2_tiehi _1807__26 (.L_HI(net26));
 sg13g2_tiehi _1847__27 (.L_HI(net27));
 sg13g2_tiehi _1806__28 (.L_HI(net28));
 sg13g2_tiehi _1854__29 (.L_HI(net29));
 sg13g2_tiehi _1805__30 (.L_HI(net30));
 sg13g2_tiehi _1846__31 (.L_HI(net31));
 sg13g2_tiehi _1804__32 (.L_HI(net32));
 sg13g2_tiehi _1853__33 (.L_HI(net33));
 sg13g2_tiehi _1803__34 (.L_HI(net34));
 sg13g2_tiehi _1845__35 (.L_HI(net35));
 sg13g2_tiehi _1802__36 (.L_HI(net36));
 sg13g2_tiehi _1852__37 (.L_HI(net37));
 sg13g2_tiehi _1801__38 (.L_HI(net38));
 sg13g2_tiehi _1844__39 (.L_HI(net39));
 sg13g2_tiehi _1800__40 (.L_HI(net40));
 sg13g2_tiehi _1850__41 (.L_HI(net41));
 sg13g2_tiehi _1799__42 (.L_HI(net42));
 sg13g2_tiehi _1843__43 (.L_HI(net43));
 sg13g2_tiehi _1798__44 (.L_HI(net44));
 sg13g2_tiehi _1851__45 (.L_HI(net45));
 sg13g2_tiehi _1797__46 (.L_HI(net46));
 sg13g2_tiehi _1842__47 (.L_HI(net47));
 sg13g2_tiehi _1796__48 (.L_HI(net48));
 sg13g2_tiehi _1857__49 (.L_HI(net49));
 sg13g2_tiehi _1795__50 (.L_HI(net50));
 sg13g2_tiehi _1841__51 (.L_HI(net51));
 sg13g2_tiehi _1794__52 (.L_HI(net52));
 sg13g2_tiehi _1793__53 (.L_HI(net53));
 sg13g2_tiehi _1792__54 (.L_HI(net54));
 sg13g2_tiehi _1791__55 (.L_HI(net55));
 sg13g2_tiehi _1790__56 (.L_HI(net56));
 sg13g2_tiehi _1789__57 (.L_HI(net57));
 sg13g2_tiehi _1788__58 (.L_HI(net58));
 sg13g2_tiehi _1787__59 (.L_HI(net59));
 sg13g2_tiehi _1786__60 (.L_HI(net60));
 sg13g2_tiehi _1785__61 (.L_HI(net61));
 sg13g2_tiehi _1784__62 (.L_HI(net62));
 sg13g2_tiehi _1840__63 (.L_HI(net63));
 sg13g2_tiehi _1783__64 (.L_HI(net64));
 sg13g2_tiehi _1838__65 (.L_HI(net65));
 sg13g2_tiehi _1782__66 (.L_HI(net66));
 sg13g2_tiehi _1837__67 (.L_HI(net67));
 sg13g2_tiehi _1781__68 (.L_HI(net68));
 sg13g2_tiehi _1836__69 (.L_HI(net69));
 sg13g2_tiehi _1780__70 (.L_HI(net70));
 sg13g2_tiehi _1835__71 (.L_HI(net71));
 sg13g2_tiehi _1779__72 (.L_HI(net72));
 sg13g2_tiehi _1834__73 (.L_HI(net73));
 sg13g2_tiehi _1778__74 (.L_HI(net74));
 sg13g2_tiehi _1833__75 (.L_HI(net75));
 sg13g2_tiehi _1832__76 (.L_HI(net76));
 sg13g2_tiehi _1831__77 (.L_HI(net77));
 sg13g2_tiehi _1830__78 (.L_HI(net78));
 sg13g2_tiehi _1829__79 (.L_HI(net79));
 sg13g2_tiehi _1828__80 (.L_HI(net80));
 sg13g2_tiehi _1776__81 (.L_HI(net81));
 sg13g2_tiehi _1827__82 (.L_HI(net82));
 sg13g2_tiehi _1826__83 (.L_HI(net83));
 sg13g2_tiehi _1825__84 (.L_HI(net84));
 sg13g2_tiehi _1824__85 (.L_HI(net85));
 sg13g2_tiehi _1823__86 (.L_HI(net86));
 sg13g2_tiehi _1822__87 (.L_HI(net87));
 sg13g2_tiehi _1821__88 (.L_HI(net88));
 sg13g2_tiehi _1820__89 (.L_HI(net89));
 sg13g2_tiehi _1819__90 (.L_HI(net90));
 sg13g2_tiehi _1818__91 (.L_HI(net91));
 sg13g2_tiehi _1839__92 (.L_HI(net92));
 sg13g2_tiehi _1817__93 (.L_HI(net93));
 sg13g2_tiehi _1816__94 (.L_HI(net94));
 sg13g2_tiehi _1815__95 (.L_HI(net95));
 sg13g2_tiehi _1814__96 (.L_HI(net96));
 sg13g2_tiehi _1813__97 (.L_HI(net97));
 sg13g2_tiehi _1812__98 (.L_HI(net98));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_rejunity_vga_logo_2 (.L_LO(net2));
 sg13g2_tielo tt_um_rejunity_vga_logo_3 (.L_LO(net3));
 sg13g2_tielo tt_um_rejunity_vga_logo_4 (.L_LO(net4));
 sg13g2_tielo tt_um_rejunity_vga_logo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_rejunity_vga_logo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_rejunity_vga_logo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_rejunity_vga_logo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_rejunity_vga_logo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_rejunity_vga_logo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_rejunity_vga_logo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_rejunity_vga_logo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rejunity_vga_logo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rejunity_vga_logo_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rejunity_vga_logo_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rejunity_vga_logo_16 (.L_LO(net16));
 sg13g2_tiehi _1811__17 (.L_HI(net17));
 sg13g2_buf_1 _1956_ (.A(vsync_prev),
    .X(uo_out[3]));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(_0218_));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(_0212_));
 sg13g2_buf_2 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_0198_),
    .X(net168));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(_0197_));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(_0196_));
 sg13g2_buf_2 fanout171 (.A(_0172_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_0375_),
    .X(net172));
 sg13g2_buf_1 fanout173 (.A(_0375_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_0366_),
    .X(net174));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(\hvsync_gen.vpos[9] ));
 sg13g2_buf_2 fanout176 (.A(net233),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(\hvsync_gen.vpos[8] ),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(net179),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(\hvsync_gen.vpos[7] ),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(\hvsync_gen.vpos[6] ),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(net183),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(net131),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(net186),
    .X(net184));
 sg13g2_buf_1 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(\hvsync_gen.vpos[4] ));
 sg13g2_buf_2 fanout187 (.A(net188),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(\hvsync_gen.vpos[3] ),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(net191),
    .X(net189));
 sg13g2_buf_1 fanout190 (.A(net191),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(\hvsync_gen.vpos[2] ),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(net236),
    .X(net192));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(net194));
 sg13g2_buf_2 fanout194 (.A(\hvsync_gen.hpos[9] ),
    .X(net194));
 sg13g2_buf_4 fanout195 (.X(net195),
    .A(net231));
 sg13g2_buf_2 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_buf_2 fanout198 (.A(net237),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(\hvsync_gen.hpos[5] ),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(\hvsync_gen.hpos[4] ),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(\hvsync_gen.hpos[4] ),
    .X(net201));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(\hvsync_gen.hpos[3] ));
 sg13g2_buf_1 fanout203 (.A(net225),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(net160),
    .X(net204));
 sg13g2_buf_1 fanout205 (.A(net160),
    .X(net205));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(net219));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(\hvsync_gen.hpos[0] ));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(_0124_));
 sg13g2_buf_2 fanout209 (.A(net210),
    .X(net209));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(rst_n));
 sg13g2_buf_2 fanout211 (.A(net212),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(net213),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(net214),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(net215),
    .X(net214));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(rst_n));
 sg13g2_tielo tt_um_rejunity_vga_logo_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(hsync),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0025_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold3 (.A(\hvsync_gen.vsync ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold4 (.A(\grad1.lfsr[12] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold5 (.A(\grad1.lfsr[10] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold6 (.A(\grad1.lfsr[9] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0024_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0089_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold9 (.A(\grad1.lfsr[18] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold10 (.A(\grad1.lfsr[17] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold11 (.A(\grad1.lfsr[8] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold12 (.A(\grad1.lfsr[14] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold13 (.A(\grad1.lfsr[13] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0014_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0068_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold16 (.A(\grad1.lfsr[16] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold17 (.A(\grad1.lfsr[15] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold18 (.A(\counter[5] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0032_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold20 (.A(\grad1.lfsr[6] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold21 (.A(\grad1.lfsr[1] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold22 (.A(\grad1.lfsr[2] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold23 (.A(\grad1.lfsr[11] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold24 (.A(\grad1.lfsr[0] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold25 (.A(\grad1.lfsr[7] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0026_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0027_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold28 (.A(\grad1.lfsr[4] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold29 (.A(\grad1.lfsr[3] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold30 (.A(\grad1.lfsr[5] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold31 (.A(\counter[2] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0029_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold33 (.A(\hvsync_gen.vpos[5] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0001_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold35 (.A(\grad1.acc[0] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold36 (.A(\counter[0] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0155_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold38 (.A(\r[11] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold39 (.A(\r[0] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold40 (.A(\counter[4] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0162_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold42 (.A(\r[16] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0059_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold44 (.A(\counter[3] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0030_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold46 (.A(\r[10] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold47 (.A(\r[1] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0044_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold49 (.A(\grad1.acc[2] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0063_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0008_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold52 (.A(\grad1.acc[4] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0064_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold54 (.A(\r[3] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold55 (.A(\grad1.lfsr[19] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0489_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold57 (.A(\r[15] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold58 (.A(\r[14] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0013_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0519_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0098_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold62 (.A(\hvsync_gen.hpos[2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0035_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold64 (.A(\r[7] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold65 (.A(\r[2] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold66 (.A(\r[4] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold67 (.A(\r[12] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold68 (.A(\hvsync_gen.hpos[7] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold69 (.A(\hvsync_gen.hpos[1] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0165_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0034_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold72 (.A(\grad1.acc[1] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold73 (.A(\r[6] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold74 (.A(\r[8] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold75 (.A(\hvsync_gen.hpos[3] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold76 (.A(\hvsync_gen.vpos[1] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold77 (.A(\grad1.acc[6] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0482_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0067_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold80 (.A(\r[9] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold81 (.A(\hvsync_gen.hpos[8] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold82 (.A(\grad1.acc[5] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold83 (.A(\hvsync_gen.vpos[8] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0005_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0056_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold86 (.A(\r[5] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold87 (.A(\hvsync_gen.hpos[5] ),
    .X(net237));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_fill_1 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_351 ();
 sg13g2_decap_4 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_380 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_fill_2 FILLER_8_315 ();
 sg13g2_fill_1 FILLER_8_317 ();
 sg13g2_fill_2 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_fill_1 FILLER_9_315 ();
 sg13g2_fill_2 FILLER_9_339 ();
 sg13g2_fill_2 FILLER_9_359 ();
 sg13g2_fill_1 FILLER_9_366 ();
 sg13g2_fill_2 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_fill_2 FILLER_10_294 ();
 sg13g2_fill_2 FILLER_10_322 ();
 sg13g2_fill_1 FILLER_10_324 ();
 sg13g2_fill_2 FILLER_10_377 ();
 sg13g2_fill_1 FILLER_10_379 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_fill_2 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_265 ();
 sg13g2_decap_8 FILLER_11_272 ();
 sg13g2_fill_2 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_281 ();
 sg13g2_decap_8 FILLER_11_286 ();
 sg13g2_fill_2 FILLER_11_334 ();
 sg13g2_fill_1 FILLER_11_340 ();
 sg13g2_fill_2 FILLER_11_365 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_fill_1 FILLER_12_245 ();
 sg13g2_fill_1 FILLER_12_303 ();
 sg13g2_fill_2 FILLER_12_312 ();
 sg13g2_fill_2 FILLER_12_349 ();
 sg13g2_fill_1 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_4 FILLER_13_224 ();
 sg13g2_fill_2 FILLER_13_228 ();
 sg13g2_fill_2 FILLER_13_266 ();
 sg13g2_fill_1 FILLER_13_268 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_fill_1 FILLER_13_297 ();
 sg13g2_fill_2 FILLER_13_321 ();
 sg13g2_fill_1 FILLER_13_323 ();
 sg13g2_fill_2 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_337 ();
 sg13g2_fill_1 FILLER_13_358 ();
 sg13g2_decap_4 FILLER_13_390 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_4 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_106 ();
 sg13g2_decap_8 FILLER_14_113 ();
 sg13g2_decap_8 FILLER_14_120 ();
 sg13g2_decap_8 FILLER_14_127 ();
 sg13g2_decap_4 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_150 ();
 sg13g2_decap_8 FILLER_14_157 ();
 sg13g2_decap_8 FILLER_14_164 ();
 sg13g2_decap_8 FILLER_14_171 ();
 sg13g2_decap_8 FILLER_14_178 ();
 sg13g2_decap_8 FILLER_14_185 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_4 FILLER_14_210 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_2 FILLER_14_246 ();
 sg13g2_fill_2 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_decap_4 FILLER_14_378 ();
 sg13g2_fill_1 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_4 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_153 ();
 sg13g2_fill_2 FILLER_15_160 ();
 sg13g2_fill_2 FILLER_15_224 ();
 sg13g2_fill_2 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_257 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_fill_2 FILLER_15_301 ();
 sg13g2_fill_2 FILLER_15_308 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_fill_2 FILLER_15_348 ();
 sg13g2_decap_4 FILLER_15_359 ();
 sg13g2_fill_2 FILLER_15_367 ();
 sg13g2_fill_1 FILLER_15_369 ();
 sg13g2_fill_2 FILLER_15_375 ();
 sg13g2_fill_1 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_4 FILLER_16_68 ();
 sg13g2_fill_1 FILLER_16_72 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_fill_2 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_177 ();
 sg13g2_fill_2 FILLER_16_182 ();
 sg13g2_fill_1 FILLER_16_184 ();
 sg13g2_decap_4 FILLER_16_200 ();
 sg13g2_fill_1 FILLER_16_204 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_4 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_276 ();
 sg13g2_fill_2 FILLER_16_290 ();
 sg13g2_fill_2 FILLER_16_318 ();
 sg13g2_fill_2 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_42 ();
 sg13g2_fill_2 FILLER_17_101 ();
 sg13g2_fill_1 FILLER_17_103 ();
 sg13g2_fill_2 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_decap_4 FILLER_17_171 ();
 sg13g2_fill_1 FILLER_17_175 ();
 sg13g2_fill_2 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_199 ();
 sg13g2_decap_4 FILLER_17_210 ();
 sg13g2_fill_1 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_219 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_241 ();
 sg13g2_decap_8 FILLER_17_282 ();
 sg13g2_decap_4 FILLER_17_289 ();
 sg13g2_fill_2 FILLER_17_293 ();
 sg13g2_decap_4 FILLER_17_298 ();
 sg13g2_fill_2 FILLER_17_302 ();
 sg13g2_fill_1 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_314 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_56 ();
 sg13g2_fill_2 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_71 ();
 sg13g2_fill_1 FILLER_18_83 ();
 sg13g2_decap_4 FILLER_18_105 ();
 sg13g2_fill_2 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_decap_4 FILLER_18_180 ();
 sg13g2_decap_4 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_fill_2 FILLER_18_216 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_4 FILLER_18_252 ();
 sg13g2_fill_2 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_365 ();
 sg13g2_fill_2 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_69 ();
 sg13g2_decap_8 FILLER_19_75 ();
 sg13g2_decap_4 FILLER_19_82 ();
 sg13g2_decap_4 FILLER_19_123 ();
 sg13g2_fill_1 FILLER_19_127 ();
 sg13g2_fill_2 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_137 ();
 sg13g2_fill_2 FILLER_19_145 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_193 ();
 sg13g2_decap_4 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_223 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_decap_4 FILLER_19_287 ();
 sg13g2_decap_4 FILLER_19_294 ();
 sg13g2_fill_2 FILLER_19_298 ();
 sg13g2_fill_2 FILLER_19_306 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_335 ();
 sg13g2_fill_1 FILLER_19_342 ();
 sg13g2_fill_1 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_366 ();
 sg13g2_fill_2 FILLER_19_384 ();
 sg13g2_fill_1 FILLER_19_386 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_58 ();
 sg13g2_decap_8 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_decap_8 FILLER_20_124 ();
 sg13g2_decap_4 FILLER_20_131 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_decap_4 FILLER_20_155 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_202 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_220 ();
 sg13g2_fill_2 FILLER_20_247 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_fill_1 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_323 ();
 sg13g2_fill_2 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_19 ();
 sg13g2_fill_2 FILLER_21_47 ();
 sg13g2_fill_2 FILLER_21_58 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_decap_4 FILLER_21_66 ();
 sg13g2_fill_2 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_78 ();
 sg13g2_fill_2 FILLER_21_92 ();
 sg13g2_fill_1 FILLER_21_94 ();
 sg13g2_decap_4 FILLER_21_99 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_decap_4 FILLER_21_114 ();
 sg13g2_fill_2 FILLER_21_130 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_1 FILLER_21_176 ();
 sg13g2_fill_2 FILLER_21_194 ();
 sg13g2_fill_2 FILLER_21_202 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_decap_4 FILLER_21_218 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_267 ();
 sg13g2_decap_4 FILLER_21_288 ();
 sg13g2_fill_1 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_decap_4 FILLER_21_313 ();
 sg13g2_fill_2 FILLER_21_317 ();
 sg13g2_fill_2 FILLER_21_324 ();
 sg13g2_fill_2 FILLER_21_337 ();
 sg13g2_fill_1 FILLER_21_339 ();
 sg13g2_fill_1 FILLER_21_354 ();
 sg13g2_decap_4 FILLER_21_358 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_decap_4 FILLER_21_371 ();
 sg13g2_fill_2 FILLER_21_375 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_41 ();
 sg13g2_fill_1 FILLER_22_43 ();
 sg13g2_fill_1 FILLER_22_100 ();
 sg13g2_decap_8 FILLER_22_121 ();
 sg13g2_fill_1 FILLER_22_140 ();
 sg13g2_fill_2 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_fill_2 FILLER_22_237 ();
 sg13g2_fill_1 FILLER_22_242 ();
 sg13g2_decap_4 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_251 ();
 sg13g2_fill_2 FILLER_22_287 ();
 sg13g2_fill_1 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_302 ();
 sg13g2_fill_2 FILLER_22_330 ();
 sg13g2_fill_1 FILLER_22_332 ();
 sg13g2_decap_4 FILLER_22_341 ();
 sg13g2_decap_4 FILLER_22_365 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_11 ();
 sg13g2_decap_4 FILLER_23_20 ();
 sg13g2_fill_2 FILLER_23_24 ();
 sg13g2_fill_1 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_59 ();
 sg13g2_fill_2 FILLER_23_66 ();
 sg13g2_decap_8 FILLER_23_90 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_fill_1 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_145 ();
 sg13g2_fill_2 FILLER_23_152 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_160 ();
 sg13g2_decap_8 FILLER_23_187 ();
 sg13g2_decap_8 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_2 FILLER_23_217 ();
 sg13g2_fill_2 FILLER_23_243 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_260 ();
 sg13g2_decap_4 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_fill_2 FILLER_23_283 ();
 sg13g2_decap_4 FILLER_23_289 ();
 sg13g2_decap_8 FILLER_23_310 ();
 sg13g2_fill_2 FILLER_23_317 ();
 sg13g2_fill_1 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_decap_4 FILLER_23_353 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_fill_2 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_55 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_121 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_fill_2 FILLER_24_194 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_216 ();
 sg13g2_fill_2 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_230 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_fill_2 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_decap_4 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_27 ();
 sg13g2_decap_4 FILLER_25_44 ();
 sg13g2_decap_4 FILLER_25_76 ();
 sg13g2_fill_2 FILLER_25_80 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_decap_8 FILLER_25_102 ();
 sg13g2_fill_1 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_136 ();
 sg13g2_fill_1 FILLER_25_138 ();
 sg13g2_decap_8 FILLER_25_149 ();
 sg13g2_fill_2 FILLER_25_156 ();
 sg13g2_fill_2 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_fill_2 FILLER_25_187 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_fill_2 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_4 FILLER_25_252 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_decap_8 FILLER_25_261 ();
 sg13g2_decap_8 FILLER_25_268 ();
 sg13g2_fill_2 FILLER_25_275 ();
 sg13g2_fill_2 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_288 ();
 sg13g2_decap_4 FILLER_25_306 ();
 sg13g2_fill_2 FILLER_25_310 ();
 sg13g2_decap_4 FILLER_25_320 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_11 ();
 sg13g2_decap_8 FILLER_26_16 ();
 sg13g2_decap_4 FILLER_26_23 ();
 sg13g2_decap_8 FILLER_26_58 ();
 sg13g2_decap_8 FILLER_26_65 ();
 sg13g2_decap_8 FILLER_26_72 ();
 sg13g2_decap_8 FILLER_26_103 ();
 sg13g2_decap_4 FILLER_26_110 ();
 sg13g2_fill_2 FILLER_26_114 ();
 sg13g2_fill_2 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_fill_2 FILLER_26_137 ();
 sg13g2_fill_1 FILLER_26_139 ();
 sg13g2_decap_4 FILLER_26_172 ();
 sg13g2_fill_2 FILLER_26_194 ();
 sg13g2_fill_1 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_fill_2 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_284 ();
 sg13g2_fill_2 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_309 ();
 sg13g2_fill_1 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_fill_1 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_fill_2 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_54 ();
 sg13g2_fill_2 FILLER_27_69 ();
 sg13g2_fill_2 FILLER_27_79 ();
 sg13g2_fill_1 FILLER_27_81 ();
 sg13g2_decap_8 FILLER_27_96 ();
 sg13g2_decap_8 FILLER_27_103 ();
 sg13g2_decap_4 FILLER_27_110 ();
 sg13g2_decap_4 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_decap_8 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_fill_1 FILLER_27_176 ();
 sg13g2_decap_8 FILLER_27_192 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_293 ();
 sg13g2_decap_4 FILLER_27_319 ();
 sg13g2_fill_2 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_365 ();
 sg13g2_fill_1 FILLER_27_367 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_9 ();
 sg13g2_fill_1 FILLER_28_23 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_decap_4 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_64 ();
 sg13g2_fill_2 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_103 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_4 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_decap_4 FILLER_28_146 ();
 sg13g2_decap_4 FILLER_28_156 ();
 sg13g2_fill_2 FILLER_28_167 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_182 ();
 sg13g2_fill_1 FILLER_28_184 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_fill_2 FILLER_28_196 ();
 sg13g2_decap_4 FILLER_28_208 ();
 sg13g2_decap_8 FILLER_28_260 ();
 sg13g2_decap_4 FILLER_28_267 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_fill_1 FILLER_28_290 ();
 sg13g2_decap_8 FILLER_28_296 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_decap_4 FILLER_28_318 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_343 ();
 sg13g2_fill_2 FILLER_28_370 ();
 sg13g2_fill_2 FILLER_28_395 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_29_26 ();
 sg13g2_fill_1 FILLER_29_43 ();
 sg13g2_fill_2 FILLER_29_52 ();
 sg13g2_fill_1 FILLER_29_54 ();
 sg13g2_fill_1 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_74 ();
 sg13g2_fill_1 FILLER_29_76 ();
 sg13g2_fill_2 FILLER_29_82 ();
 sg13g2_decap_8 FILLER_29_101 ();
 sg13g2_fill_2 FILLER_29_108 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_182 ();
 sg13g2_fill_2 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_212 ();
 sg13g2_fill_2 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_decap_8 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_decap_4 FILLER_29_348 ();
 sg13g2_fill_2 FILLER_29_352 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_55 ();
 sg13g2_fill_2 FILLER_30_62 ();
 sg13g2_fill_2 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_90 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_146 ();
 sg13g2_fill_2 FILLER_30_153 ();
 sg13g2_fill_1 FILLER_30_155 ();
 sg13g2_fill_2 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_fill_2 FILLER_30_189 ();
 sg13g2_fill_2 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_242 ();
 sg13g2_decap_4 FILLER_30_249 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_decap_4 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_decap_4 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_fill_2 FILLER_30_311 ();
 sg13g2_decap_8 FILLER_30_318 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_4 FILLER_30_349 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_31_52 ();
 sg13g2_fill_1 FILLER_31_54 ();
 sg13g2_decap_4 FILLER_31_68 ();
 sg13g2_fill_2 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_89 ();
 sg13g2_decap_4 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_173 ();
 sg13g2_fill_1 FILLER_31_183 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_fill_1 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_278 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_fill_2 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_15 ();
 sg13g2_fill_1 FILLER_32_17 ();
 sg13g2_decap_8 FILLER_32_22 ();
 sg13g2_fill_2 FILLER_32_29 ();
 sg13g2_fill_1 FILLER_32_31 ();
 sg13g2_fill_2 FILLER_32_45 ();
 sg13g2_fill_1 FILLER_32_47 ();
 sg13g2_fill_1 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_155 ();
 sg13g2_fill_1 FILLER_32_206 ();
 sg13g2_fill_2 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_233 ();
 sg13g2_fill_2 FILLER_32_244 ();
 sg13g2_decap_4 FILLER_32_251 ();
 sg13g2_decap_8 FILLER_32_281 ();
 sg13g2_fill_2 FILLER_32_288 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_decap_4 FILLER_32_302 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_decap_4 FILLER_32_352 ();
 sg13g2_fill_2 FILLER_32_361 ();
 sg13g2_fill_1 FILLER_32_363 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_15 ();
 sg13g2_decap_4 FILLER_33_25 ();
 sg13g2_fill_1 FILLER_33_29 ();
 sg13g2_fill_2 FILLER_33_43 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_1 FILLER_33_72 ();
 sg13g2_fill_1 FILLER_33_82 ();
 sg13g2_fill_1 FILLER_33_92 ();
 sg13g2_decap_4 FILLER_33_97 ();
 sg13g2_fill_2 FILLER_33_101 ();
 sg13g2_fill_2 FILLER_33_111 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_fill_2 FILLER_33_123 ();
 sg13g2_fill_1 FILLER_33_125 ();
 sg13g2_decap_4 FILLER_33_146 ();
 sg13g2_fill_2 FILLER_33_166 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_decap_4 FILLER_33_184 ();
 sg13g2_fill_1 FILLER_33_188 ();
 sg13g2_decap_4 FILLER_33_215 ();
 sg13g2_decap_4 FILLER_33_223 ();
 sg13g2_fill_2 FILLER_33_246 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_258 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_decap_8 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_356 ();
 sg13g2_fill_1 FILLER_33_375 ();
 sg13g2_fill_2 FILLER_33_394 ();
 sg13g2_fill_2 FILLER_34_48 ();
 sg13g2_fill_1 FILLER_34_50 ();
 sg13g2_fill_2 FILLER_34_73 ();
 sg13g2_fill_1 FILLER_34_75 ();
 sg13g2_fill_2 FILLER_34_89 ();
 sg13g2_fill_1 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_113 ();
 sg13g2_fill_2 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_156 ();
 sg13g2_fill_1 FILLER_34_158 ();
 sg13g2_fill_2 FILLER_34_163 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_decap_4 FILLER_34_171 ();
 sg13g2_decap_8 FILLER_34_230 ();
 sg13g2_fill_1 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_fill_1 FILLER_35_30 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_fill_2 FILLER_35_74 ();
 sg13g2_fill_2 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_116 ();
 sg13g2_decap_8 FILLER_35_174 ();
 sg13g2_decap_8 FILLER_35_181 ();
 sg13g2_decap_4 FILLER_35_188 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_decap_4 FILLER_35_198 ();
 sg13g2_fill_1 FILLER_35_202 ();
 sg13g2_decap_4 FILLER_35_212 ();
 sg13g2_decap_8 FILLER_35_268 ();
 sg13g2_decap_4 FILLER_35_275 ();
 sg13g2_fill_1 FILLER_35_279 ();
 sg13g2_decap_8 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_decap_4 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_decap_4 FILLER_35_354 ();
 sg13g2_fill_2 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_decap_4 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_38 ();
 sg13g2_decap_4 FILLER_36_43 ();
 sg13g2_fill_2 FILLER_36_47 ();
 sg13g2_fill_1 FILLER_36_53 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_117 ();
 sg13g2_fill_2 FILLER_36_135 ();
 sg13g2_fill_2 FILLER_36_162 ();
 sg13g2_fill_1 FILLER_36_164 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_230 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_decap_4 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_248 ();
 sg13g2_decap_8 FILLER_36_253 ();
 sg13g2_decap_4 FILLER_36_260 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_decap_8 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_299 ();
 sg13g2_decap_8 FILLER_36_306 ();
 sg13g2_decap_8 FILLER_36_313 ();
 sg13g2_decap_8 FILLER_36_320 ();
 sg13g2_decap_8 FILLER_36_327 ();
 sg13g2_decap_8 FILLER_36_334 ();
 sg13g2_decap_8 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_362 ();
 sg13g2_decap_8 FILLER_36_369 ();
 sg13g2_decap_8 FILLER_36_376 ();
 sg13g2_decap_8 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_fill_2 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_79 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_fill_2 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_104 ();
 sg13g2_fill_1 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_118 ();
 sg13g2_fill_1 FILLER_37_120 ();
 sg13g2_fill_2 FILLER_37_146 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_decap_8 FILLER_37_163 ();
 sg13g2_decap_8 FILLER_37_170 ();
 sg13g2_fill_1 FILLER_37_177 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_4 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_200 ();
 sg13g2_decap_8 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_265 ();
 sg13g2_decap_4 FILLER_37_272 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_101 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_fill_2 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_149 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_254 ();
 sg13g2_decap_8 FILLER_38_261 ();
 sg13g2_decap_8 FILLER_38_268 ();
 sg13g2_decap_8 FILLER_38_275 ();
 sg13g2_decap_8 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_310 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule

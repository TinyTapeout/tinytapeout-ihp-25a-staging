module tt_um_daosvik_aesinvsbox (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire \sbox_aesinv_inst.x0 ;
 wire \sbox_aesinv_inst.x00000008 ;
 wire \sbox_aesinv_inst.x00000013 ;
 wire \sbox_aesinv_inst.x00000054 ;
 wire \sbox_aesinv_inst.x00000080 ;
 wire \sbox_aesinv_inst.x00000117 ;
 wire \sbox_aesinv_inst.x00000550 ;
 wire \sbox_aesinv_inst.x00001011 ;
 wire \sbox_aesinv_inst.x0000101a ;
 wire \sbox_aesinv_inst.x000010dc ;
 wire \sbox_aesinv_inst.x00001110 ;
 wire \sbox_aesinv_inst.x00001175 ;
 wire \sbox_aesinv_inst.x00001355 ;
 wire \sbox_aesinv_inst.x00008000 ;
 wire \sbox_aesinv_inst.x00008880 ;
 wire \sbox_aesinv_inst.x0000a000 ;
 wire \sbox_aesinv_inst.x00010005 ;
 wire \sbox_aesinv_inst.x00010031 ;
 wire \sbox_aesinv_inst.x00050011 ;
 wire \sbox_aesinv_inst.x00050022 ;
 wire \sbox_aesinv_inst.x00050300 ;
 wire \sbox_aesinv_inst.x00060006 ;
 wire \sbox_aesinv_inst.x00070013 ;
 wire \sbox_aesinv_inst.x0007173f ;
 wire \sbox_aesinv_inst.x000a022a ;
 wire \sbox_aesinv_inst.x000a0808 ;
 wire \sbox_aesinv_inst.x000aaaab ;
 wire \sbox_aesinv_inst.x000c0e5e ;
 wire \sbox_aesinv_inst.x000ccc00 ;
 wire \sbox_aesinv_inst.x000f023f ;
 wire \sbox_aesinv_inst.x00113035 ;
 wire \sbox_aesinv_inst.x00130f0f ;
 wire \sbox_aesinv_inst.x00330404 ;
 wire \sbox_aesinv_inst.x004000c0 ;
 wire \sbox_aesinv_inst.x005dccdd ;
 wire \sbox_aesinv_inst.x007fabff ;
 wire \sbox_aesinv_inst.x01 ;
 wire \sbox_aesinv_inst.x0100011f ;
 wire \sbox_aesinv_inst.x01010003 ;
 wire \sbox_aesinv_inst.x01011010 ;
 wire \sbox_aesinv_inst.x01155fff ;
 wire \sbox_aesinv_inst.x0133273f ;
 wire \sbox_aesinv_inst.x0137133f ;
 wire \sbox_aesinv_inst.x01f731f7 ;
 wire \sbox_aesinv_inst.x02 ;
 wire \sbox_aesinv_inst.x03fc03fc ;
 wire \sbox_aesinv_inst.x04 ;
 wire \sbox_aesinv_inst.x04044447 ;
 wire \sbox_aesinv_inst.x040c0000 ;
 wire \sbox_aesinv_inst.x05500000 ;
 wire \sbox_aesinv_inst.x055f0557 ;
 wire \sbox_aesinv_inst.x08 ;
 wire \sbox_aesinv_inst.x08000000 ;
 wire \sbox_aesinv_inst.x0a ;
 wire \sbox_aesinv_inst.x0a000000 ;
 wire \sbox_aesinv_inst.x0a080000 ;
 wire \sbox_aesinv_inst.x0abf1bbf ;
 wire \sbox_aesinv_inst.x0b ;
 wire \sbox_aesinv_inst.x0b1fafbf ;
 wire \sbox_aesinv_inst.x0c ;
 wire \sbox_aesinv_inst.x0cd37660 ;
 wire \sbox_aesinv_inst.x0d ;
 wire \sbox_aesinv_inst.x0e0a0000 ;
 wire \sbox_aesinv_inst.x0eb6ef2f ;
 wire \sbox_aesinv_inst.x0f5f0a5f ;
 wire \sbox_aesinv_inst.x0ff7ffff ;
 wire \sbox_aesinv_inst.x1 ;
 wire \sbox_aesinv_inst.x10 ;
 wire \sbox_aesinv_inst.x10104040 ;
 wire \sbox_aesinv_inst.x11004400 ;
 wire \sbox_aesinv_inst.x11131313 ;
 wire \sbox_aesinv_inst.x11771333 ;
 wire \sbox_aesinv_inst.x11aa0000 ;
 wire \sbox_aesinv_inst.x12bf5b4f ;
 wire \sbox_aesinv_inst.x131317df ;
 wire \sbox_aesinv_inst.x1333131f ;
 wire \sbox_aesinv_inst.x135f5fdf ;
 wire \sbox_aesinv_inst.x13bfbfbf ;
 wire \sbox_aesinv_inst.x15000400 ;
 wire \sbox_aesinv_inst.x151d777f ;
 wire \sbox_aesinv_inst.x15555050 ;
 wire \sbox_aesinv_inst.x169287dc ;
 wire \sbox_aesinv_inst.x175f333f ;
 wire \sbox_aesinv_inst.x17ff555f ;
 wire \sbox_aesinv_inst.x1a ;
 wire \sbox_aesinv_inst.x1a10b72b ;
 wire \sbox_aesinv_inst.x1b ;
 wire \sbox_aesinv_inst.x1c ;
 wire \sbox_aesinv_inst.x1d ;
 wire \sbox_aesinv_inst.x1d7f5dff ;
 wire \sbox_aesinv_inst.x1f7b28d7 ;
 wire \sbox_aesinv_inst.x1f7f55ff ;
 wire \sbox_aesinv_inst.x2 ;
 wire \sbox_aesinv_inst.x20 ;
 wire \sbox_aesinv_inst.x229616fd ;
 wire \sbox_aesinv_inst.x23369e29 ;
 wire \sbox_aesinv_inst.x23853f57 ;
 wire \sbox_aesinv_inst.x24cc4461 ;
 wire \sbox_aesinv_inst.x2a ;
 wire \sbox_aesinv_inst.x2a000000 ;
 wire \sbox_aesinv_inst.x2aeeaaee ;
 wire \sbox_aesinv_inst.x2b ;
 wire \sbox_aesinv_inst.x2bffafff ;
 wire \sbox_aesinv_inst.x2c ;
 wire \sbox_aesinv_inst.x2c6cdf10 ;
 wire \sbox_aesinv_inst.x2ca62526 ;
 wire \sbox_aesinv_inst.x2d ;
 wire \sbox_aesinv_inst.x2d9fb2de ;
 wire \sbox_aesinv_inst.x2fa5e682 ;
 wire \sbox_aesinv_inst.x2fafffff ;
 wire \sbox_aesinv_inst.x3 ;
 wire \sbox_aesinv_inst.x30307000 ;
 wire \sbox_aesinv_inst.x3030f1f0 ;
 wire \sbox_aesinv_inst.x30c030c0 ;
 wire \sbox_aesinv_inst.x318ab4e1 ;
 wire \sbox_aesinv_inst.x32220000 ;
 wire \sbox_aesinv_inst.x32302020 ;
 wire \sbox_aesinv_inst.x323233fb ;
 wire \sbox_aesinv_inst.x326fc4dd ;
 wire \sbox_aesinv_inst.x333300cf ;
 wire \sbox_aesinv_inst.x33cfffff ;
 wire \sbox_aesinv_inst.x33ffff0f ;
 wire \sbox_aesinv_inst.x37303733 ;
 wire \sbox_aesinv_inst.x3777053f ;
 wire \sbox_aesinv_inst.x37ff5577 ;
 wire \sbox_aesinv_inst.x39fe8cff ;
 wire \sbox_aesinv_inst.x3a ;
 wire \sbox_aesinv_inst.x3b ;
 wire \sbox_aesinv_inst.x3c ;
 wire \sbox_aesinv_inst.x3c3ffdff ;
 wire \sbox_aesinv_inst.x3cf25843 ;
 wire \sbox_aesinv_inst.x3d ;
 wire \sbox_aesinv_inst.x3f00ff05 ;
 wire \sbox_aesinv_inst.x3f0fffcf ;
 wire \sbox_aesinv_inst.x3f557fff ;
 wire \sbox_aesinv_inst.x3fff2faf ;
 wire \sbox_aesinv_inst.x3fffffff ;
 wire \sbox_aesinv_inst.x4 ;
 wire \sbox_aesinv_inst.x40 ;
 wire \sbox_aesinv_inst.x40484048 ;
 wire \sbox_aesinv_inst.x40c00000 ;
 wire \sbox_aesinv_inst.x41d5cc5c ;
 wire \sbox_aesinv_inst.x4213e265 ;
 wire \sbox_aesinv_inst.x42e28881 ;
 wire \sbox_aesinv_inst.x4332245f ;
 wire \sbox_aesinv_inst.x434a8cf5 ;
 wire \sbox_aesinv_inst.x43fecdd2 ;
 wire \sbox_aesinv_inst.x4638af86 ;
 wire \sbox_aesinv_inst.x4a ;
 wire \sbox_aesinv_inst.x4b ;
 wire \sbox_aesinv_inst.x4c ;
 wire \sbox_aesinv_inst.x4d ;
 wire \sbox_aesinv_inst.x4e5feeff ;
 wire \sbox_aesinv_inst.x5 ;
 wire \sbox_aesinv_inst.x50004000 ;
 wire \sbox_aesinv_inst.x52af6f23 ;
 wire \sbox_aesinv_inst.x52c516d9 ;
 wire \sbox_aesinv_inst.x54eaa319 ;
 wire \sbox_aesinv_inst.x55556666 ;
 wire \sbox_aesinv_inst.x55775071 ;
 wire \sbox_aesinv_inst.x557f00ff ;
 wire \sbox_aesinv_inst.x571fff3f ;
 wire \sbox_aesinv_inst.x57ffff00 ;
 wire \sbox_aesinv_inst.x5a ;
 wire \sbox_aesinv_inst.x5a5f5b5f ;
 wire \sbox_aesinv_inst.x5aaa5aaa ;
 wire \sbox_aesinv_inst.x5b ;
 wire \sbox_aesinv_inst.x5b847ba9 ;
 wire \sbox_aesinv_inst.x5c ;
 wire \sbox_aesinv_inst.x5d ;
 wire \sbox_aesinv_inst.x5e9f51e4 ;
 wire \sbox_aesinv_inst.x5f5ffafa ;
 wire \sbox_aesinv_inst.x5fff0faf ;
 wire \sbox_aesinv_inst.x6 ;
 wire \sbox_aesinv_inst.x6191ae47 ;
 wire \sbox_aesinv_inst.x6a ;
 wire \sbox_aesinv_inst.x6a86145f ;
 wire \sbox_aesinv_inst.x6ad30f0f ;
 wire \sbox_aesinv_inst.x6b ;
 wire \sbox_aesinv_inst.x6c ;
 wire \sbox_aesinv_inst.x6d ;
 wire \sbox_aesinv_inst.x6d287e63 ;
 wire \sbox_aesinv_inst.x7 ;
 wire \sbox_aesinv_inst.x7077f7ff ;
 wire \sbox_aesinv_inst.x777717ff ;
 wire \sbox_aesinv_inst.x77cd77ff ;
 wire \sbox_aesinv_inst.x77fc77fc ;
 wire \sbox_aesinv_inst.x77ff3337 ;
 wire \sbox_aesinv_inst.x7847e6db ;
 wire \sbox_aesinv_inst.x7a ;
 wire \sbox_aesinv_inst.x7b ;
 wire \sbox_aesinv_inst.x7c ;
 wire \sbox_aesinv_inst.x7c7c7c7d ;
 wire \sbox_aesinv_inst.x7ca10f66 ;
 wire \sbox_aesinv_inst.x7d ;
 wire \sbox_aesinv_inst.x7f5f3300 ;
 wire \sbox_aesinv_inst.x80 ;
 wire \sbox_aesinv_inst.x80000000 ;
 wire \sbox_aesinv_inst.x80808080 ;
 wire \sbox_aesinv_inst.x854f7ef5 ;
 wire \sbox_aesinv_inst.x88000000 ;
 wire \sbox_aesinv_inst.x88008800 ;
 wire \sbox_aesinv_inst.x88880000 ;
 wire \sbox_aesinv_inst.x88888888 ;
 wire \sbox_aesinv_inst.x8ad2e815 ;
 wire \sbox_aesinv_inst.x8b30445b ;
 wire \sbox_aesinv_inst.x8df398a3 ;
 wire \sbox_aesinv_inst.x8fdfffff ;
 wire \sbox_aesinv_inst.x96492239 ;
 wire \sbox_aesinv_inst.x9d97aa84 ;
 wire \sbox_aesinv_inst.xa0008000 ;
 wire \sbox_aesinv_inst.xa000a000 ;
 wire \sbox_aesinv_inst.xa0a00000 ;
 wire \sbox_aesinv_inst.xa0a0a0a0 ;
 wire \sbox_aesinv_inst.xa0a0a1a1 ;
 wire \sbox_aesinv_inst.xa0fb7cd2 ;
 wire \sbox_aesinv_inst.xa1b3a5bf ;
 wire \sbox_aesinv_inst.xa4b75f65 ;
 wire \sbox_aesinv_inst.xa8000000 ;
 wire \sbox_aesinv_inst.xa8008000 ;
 wire \sbox_aesinv_inst.xa8800000 ;
 wire \sbox_aesinv_inst.xa8a8a8a8 ;
 wire \sbox_aesinv_inst.xa90301b8 ;
 wire \sbox_aesinv_inst.xa9e15289 ;
 wire \sbox_aesinv_inst.xaa000000 ;
 wire \sbox_aesinv_inst.xaa0faf5f ;
 wire \sbox_aesinv_inst.xaa88aa88 ;
 wire \sbox_aesinv_inst.xaaa0aaa0 ;
 wire \sbox_aesinv_inst.xaaaa0000 ;
 wire \sbox_aesinv_inst.xaaaa8888 ;
 wire \sbox_aesinv_inst.xaaaaa0a0 ;
 wire \sbox_aesinv_inst.xaaaaaa00 ;
 wire \sbox_aesinv_inst.xaaaf153f ;
 wire \sbox_aesinv_inst.xadffadff ;
 wire \sbox_aesinv_inst.xaf7faf7f ;
 wire \sbox_aesinv_inst.xafa5ffff ;
 wire \sbox_aesinv_inst.xb047c23f ;
 wire \sbox_aesinv_inst.xb1b1f5f7 ;
 wire \sbox_aesinv_inst.xbb3333ff ;
 wire \sbox_aesinv_inst.xbb77ffff ;
 wire \sbox_aesinv_inst.xbbbbf5f5 ;
 wire \sbox_aesinv_inst.xbfbf373f ;
 wire \sbox_aesinv_inst.xbfffffff ;
 wire \sbox_aesinv_inst.xc0008000 ;
 wire \sbox_aesinv_inst.xc000c000 ;
 wire \sbox_aesinv_inst.xc011c011 ;
 wire \sbox_aesinv_inst.xc0c00000 ;
 wire \sbox_aesinv_inst.xc0c0c0c0 ;
 wire \sbox_aesinv_inst.xc3c3c3cf ;
 wire \sbox_aesinv_inst.xc4cf14da ;
 wire \sbox_aesinv_inst.xc5cfc5df ;
 wire \sbox_aesinv_inst.xc60b25d3 ;
 wire \sbox_aesinv_inst.xc6aca424 ;
 wire \sbox_aesinv_inst.xc800c000 ;
 wire \sbox_aesinv_inst.xc8c8c8c8 ;
 wire \sbox_aesinv_inst.xcbea0a80 ;
 wire \sbox_aesinv_inst.xcbffcbff ;
 wire \sbox_aesinv_inst.xcc000000 ;
 wire \sbox_aesinv_inst.xcc00cc00 ;
 wire \sbox_aesinv_inst.xcc880000 ;
 wire \sbox_aesinv_inst.xcc88cc88 ;
 wire \sbox_aesinv_inst.xccc0ccc0 ;
 wire \sbox_aesinv_inst.xcccc0000 ;
 wire \sbox_aesinv_inst.xcccc8888 ;
 wire \sbox_aesinv_inst.xccccc0c0 ;
 wire \sbox_aesinv_inst.xcccccc00 ;
 wire \sbox_aesinv_inst.xcccf030f ;
 wire \sbox_aesinv_inst.xd1f16c3a ;
 wire \sbox_aesinv_inst.xd2a0de7f ;
 wire \sbox_aesinv_inst.xd7997ddd ;
 wire \sbox_aesinv_inst.xdd11cc00 ;
 wire \sbox_aesinv_inst.xdd5555ff ;
 wire \sbox_aesinv_inst.xdd7fff7f ;
 wire \sbox_aesinv_inst.xddf7ddf7 ;
 wire \sbox_aesinv_inst.xdf77df77 ;
 wire \sbox_aesinv_inst.xdfc11244 ;
 wire \sbox_aesinv_inst.xdfdf77ff ;
 wire \sbox_aesinv_inst.xe080c000 ;
 wire \sbox_aesinv_inst.xe0e0e0e0 ;
 wire \sbox_aesinv_inst.xe2cda26e ;
 wire \sbox_aesinv_inst.xe3ab5bd2 ;
 wire \sbox_aesinv_inst.xe8133bb7 ;
 wire \sbox_aesinv_inst.xe8e8e800 ;
 wire \sbox_aesinv_inst.xeaeaeaea ;
 wire \sbox_aesinv_inst.xeaefffff ;
 wire \sbox_aesinv_inst.xee00ee00 ;
 wire \sbox_aesinv_inst.xeeaaeeaa ;
 wire \sbox_aesinv_inst.xeecc98e2 ;
 wire \sbox_aesinv_inst.xeeee0000 ;
 wire \sbox_aesinv_inst.xeeee8080 ;
 wire \sbox_aesinv_inst.xeeeeaaaa ;
 wire \sbox_aesinv_inst.xeeeeeeee ;
 wire \sbox_aesinv_inst.xef715dd5 ;
 wire \sbox_aesinv_inst.xefefcf8f ;
 wire \sbox_aesinv_inst.xf0000000 ;
 wire \sbox_aesinv_inst.xf000f000 ;
 wire \sbox_aesinv_inst.xf003f003 ;
 wire \sbox_aesinv_inst.xf0a0a0a0 ;
 wire \sbox_aesinv_inst.xf0a0f0a0 ;
 wire \sbox_aesinv_inst.xf0a0f3a3 ;
 wire \sbox_aesinv_inst.xf0c0c000 ;
 wire \sbox_aesinv_inst.xf0c0f0c0 ;
 wire \sbox_aesinv_inst.xf0c0f5d5 ;
 wire \sbox_aesinv_inst.xf0f00000 ;
 wire \sbox_aesinv_inst.xf0f0a0a0 ;
 wire \sbox_aesinv_inst.xf0f0c0c0 ;
 wire \sbox_aesinv_inst.xf0f0f000 ;
 wire \sbox_aesinv_inst.xf0f0f0f0 ;
 wire \sbox_aesinv_inst.xf12405c2 ;
 wire \sbox_aesinv_inst.xf1a1f1a1 ;
 wire \sbox_aesinv_inst.xf1f1ffff ;
 wire \sbox_aesinv_inst.xf1f5f5f7 ;
 wire \sbox_aesinv_inst.xf333f377 ;
 wire \sbox_aesinv_inst.xf33fffff ;
 wire \sbox_aesinv_inst.xf35ff3ff ;
 wire \sbox_aesinv_inst.xf3f37f7f ;
 wire \sbox_aesinv_inst.xf446ce08 ;
 wire \sbox_aesinv_inst.xf4bcfdb0 ;
 wire \sbox_aesinv_inst.xf555f57f ;
 wire \sbox_aesinv_inst.xf5a5ffff ;
 wire \sbox_aesinv_inst.xf5ff5fff ;
 wire \sbox_aesinv_inst.xf8008000 ;
 wire \sbox_aesinv_inst.xf8f0c800 ;
 wire \sbox_aesinv_inst.xf8f8c8c8 ;
 wire \sbox_aesinv_inst.xfa00fa00 ;
 wire \sbox_aesinv_inst.xfaaafaaa ;
 wire \sbox_aesinv_inst.xfac8a080 ;
 wire \sbox_aesinv_inst.xfaf8fa00 ;
 wire \sbox_aesinv_inst.xfafa0000 ;
 wire \sbox_aesinv_inst.xfafaaaaa ;
 wire \sbox_aesinv_inst.xfafafafa ;
 wire \sbox_aesinv_inst.xfc00fc00 ;
 wire \sbox_aesinv_inst.xfccca000 ;
 wire \sbox_aesinv_inst.xfcccfccc ;
 wire \sbox_aesinv_inst.xfccfffff ;
 wire \sbox_aesinv_inst.xfcecf8a0 ;
 wire \sbox_aesinv_inst.xfcfc0000 ;
 wire \sbox_aesinv_inst.xfcfccccc ;
 wire \sbox_aesinv_inst.xfcfcccff ;
 wire \sbox_aesinv_inst.xfcfcf8a0 ;
 wire \sbox_aesinv_inst.xfcfcfcfc ;
 wire \sbox_aesinv_inst.xfd11ffff ;
 wire \sbox_aesinv_inst.xfec8eec8 ;
 wire \sbox_aesinv_inst.xfecccc00 ;
 wire \sbox_aesinv_inst.xfeccfec8 ;
 wire \sbox_aesinv_inst.xfeecfaa8 ;
 wire \sbox_aesinv_inst.xfeeef8a8 ;
 wire \sbox_aesinv_inst.xfefaeca8 ;
 wire \sbox_aesinv_inst.xfefafefa ;
 wire \sbox_aesinv_inst.xfefea8a0 ;
 wire \sbox_aesinv_inst.xfefefefe ;
 wire \sbox_aesinv_inst.xff000000 ;
 wire \sbox_aesinv_inst.xff00aa00 ;
 wire \sbox_aesinv_inst.xff00cc00 ;
 wire \sbox_aesinv_inst.xff00f000 ;
 wire \sbox_aesinv_inst.xff00ff00 ;
 wire \sbox_aesinv_inst.xff010103 ;
 wire \sbox_aesinv_inst.xff05333f ;
 wire \sbox_aesinv_inst.xff3f05ff ;
 wire \sbox_aesinv_inst.xff7f7f7f ;
 wire \sbox_aesinv_inst.xffaa0000 ;
 wire \sbox_aesinv_inst.xffaaaaaa ;
 wire \sbox_aesinv_inst.xffaaffaa ;
 wire \sbox_aesinv_inst.xffb3ffb3 ;
 wire \sbox_aesinv_inst.xffcc0000 ;
 wire \sbox_aesinv_inst.xffcccccc ;
 wire \sbox_aesinv_inst.xffcceec8 ;
 wire \sbox_aesinv_inst.xffccffcc ;
 wire \sbox_aesinv_inst.xffddddff ;
 wire \sbox_aesinv_inst.xffec8888 ;
 wire \sbox_aesinv_inst.xffecece8 ;
 wire \sbox_aesinv_inst.xffecffa8 ;
 wire \sbox_aesinv_inst.xffeeee88 ;
 wire \sbox_aesinv_inst.xffeeffee ;
 wire \sbox_aesinv_inst.xfff00000 ;
 wire \sbox_aesinv_inst.xfff0f0f0 ;
 wire \sbox_aesinv_inst.xfff0fff0 ;
 wire \sbox_aesinv_inst.xfff30000 ;
 wire \sbox_aesinv_inst.xfff5f5ff ;
 wire \sbox_aesinv_inst.xfff8fac8 ;
 wire \sbox_aesinv_inst.xfff8ffa0 ;
 wire \sbox_aesinv_inst.xfffafffa ;
 wire \sbox_aesinv_inst.xfffcfeec ;
 wire \sbox_aesinv_inst.xfffcfffc ;
 wire \sbox_aesinv_inst.xfffcfffd ;
 wire \sbox_aesinv_inst.xfffef888 ;
 wire \sbox_aesinv_inst.xffff0000 ;
 wire \sbox_aesinv_inst.xffff8f0f ;
 wire \sbox_aesinv_inst.xffffaaaa ;
 wire \sbox_aesinv_inst.xffffcccc ;
 wire \sbox_aesinv_inst.xffffeeee ;
 wire \sbox_aesinv_inst.xfffff0f0 ;
 wire \sbox_aesinv_inst.xfffff8a0 ;
 wire \sbox_aesinv_inst.xfffffafa ;
 wire \sbox_aesinv_inst.xfffffcfc ;
 wire \sbox_aesinv_inst.xfffffeee ;
 wire \sbox_aesinv_inst.xffffff00 ;
 wire \sbox_aesinv_inst.xffffffaa ;
 wire \sbox_aesinv_inst.xffffffcc ;
 wire \sbox_aesinv_inst.xffffffdd ;
 wire \sbox_aesinv_inst.xffffffea ;
 wire \sbox_aesinv_inst.xffffffec ;
 wire \sbox_aesinv_inst.xfffffff0 ;
 wire \sbox_aesinv_inst.xfffffffc ;
 wire \sbox_aesinv_inst.xfffffffe ;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire \sbox_aesinv_inst.m00000550/_0_ ;
 wire \sbox_aesinv_inst.m0000101a/_0_ ;
 wire \sbox_aesinv_inst.m000010dc/_0_ ;
 wire \sbox_aesinv_inst.m00001175/_0_ ;
 wire \sbox_aesinv_inst.m00001355/_0_ ;
 wire \sbox_aesinv_inst.m00010031/_0_ ;
 wire \sbox_aesinv_inst.m00050011/_0_ ;
 wire \sbox_aesinv_inst.m00050022/_0_ ;
 wire \sbox_aesinv_inst.m00050300/_0_ ;
 wire \sbox_aesinv_inst.m00060006/_0_ ;
 wire \sbox_aesinv_inst.m00070013/_0_ ;
 wire \sbox_aesinv_inst.m0007173f/_0_ ;
 wire \sbox_aesinv_inst.m000a022a/_0_ ;
 wire \sbox_aesinv_inst.m000aaaab/_0_ ;
 wire \sbox_aesinv_inst.m000f023f/_0_ ;
 wire \sbox_aesinv_inst.m00113035/_0_ ;
 wire \sbox_aesinv_inst.m00130f0f/_0_ ;
 wire \sbox_aesinv_inst.m00330404/_0_ ;
 wire \sbox_aesinv_inst.m007fabff/_0_ ;
 wire \sbox_aesinv_inst.m0100011f/_0_ ;
 wire \sbox_aesinv_inst.m01010003/_0_ ;
 wire \sbox_aesinv_inst.m01011010/_0_ ;
 wire \sbox_aesinv_inst.m01155fff/_0_ ;
 wire \sbox_aesinv_inst.m0133273f/_0_ ;
 wire \sbox_aesinv_inst.m0137133f/_0_ ;
 wire \sbox_aesinv_inst.m01f731f7/_0_ ;
 wire \sbox_aesinv_inst.m02/_0_ ;
 wire \sbox_aesinv_inst.m04/_0_ ;
 wire \sbox_aesinv_inst.m04044447/_0_ ;
 wire \sbox_aesinv_inst.m055f0557/_0_ ;
 wire \sbox_aesinv_inst.m08/_0_ ;
 wire \sbox_aesinv_inst.m0abf1bbf/_0_ ;
 wire \sbox_aesinv_inst.m0b1fafbf/_0_ ;
 wire \sbox_aesinv_inst.m0eb6ef2f/_0_ ;
 wire \sbox_aesinv_inst.m0f5f0a5f/_0_ ;
 wire \sbox_aesinv_inst.m0ff7ffff/_0_ ;
 wire \sbox_aesinv_inst.m10/_0_ ;
 wire \sbox_aesinv_inst.m11771333/_0_ ;
 wire \sbox_aesinv_inst.m131317df/_0_ ;
 wire \sbox_aesinv_inst.m1333131f/_0_ ;
 wire \sbox_aesinv_inst.m135f5fdf/_0_ ;
 wire \sbox_aesinv_inst.m13bfbfbf/_0_ ;
 wire \sbox_aesinv_inst.m151d777f/_0_ ;
 wire \sbox_aesinv_inst.m15555050/_0_ ;
 wire \sbox_aesinv_inst.m169287dc/_0_ ;
 wire \sbox_aesinv_inst.m175f333f/_0_ ;
 wire \sbox_aesinv_inst.m17ff555f/_0_ ;
 wire \sbox_aesinv_inst.m1a10b72b/_0_ ;
 wire \sbox_aesinv_inst.m1d7f5dff/_0_ ;
 wire \sbox_aesinv_inst.m1f7f55ff/_0_ ;
 wire \sbox_aesinv_inst.m20/_0_ ;
 wire \sbox_aesinv_inst.m229616fd/_0_ ;
 wire \sbox_aesinv_inst.m24cc4461/_0_ ;
 wire \sbox_aesinv_inst.m2aeeaaee/_0_ ;
 wire \sbox_aesinv_inst.m2bffafff/_0_ ;
 wire \sbox_aesinv_inst.m2d9fb2de/_0_ ;
 wire \sbox_aesinv_inst.m2fa5e682/_0_ ;
 wire \sbox_aesinv_inst.m3030f1f0/_0_ ;
 wire \sbox_aesinv_inst.m318ab4e1/_0_ ;
 wire \sbox_aesinv_inst.m323233fb/_0_ ;
 wire \sbox_aesinv_inst.m333300cf/_0_ ;
 wire \sbox_aesinv_inst.m33cfffff/_0_ ;
 wire \sbox_aesinv_inst.m33ffff0f/_0_ ;
 wire \sbox_aesinv_inst.m37303733/_0_ ;
 wire \sbox_aesinv_inst.m3777053f/_0_ ;
 wire \sbox_aesinv_inst.m37ff5577/_0_ ;
 wire \sbox_aesinv_inst.m3c3ffdff/_0_ ;
 wire \sbox_aesinv_inst.m3cf25843/_0_ ;
 wire \sbox_aesinv_inst.m3f0fffcf/_0_ ;
 wire \sbox_aesinv_inst.m3f557fff/_0_ ;
 wire \sbox_aesinv_inst.m3fff2faf/_0_ ;
 wire \sbox_aesinv_inst.m40/_0_ ;
 wire \sbox_aesinv_inst.m4213e265/_0_ ;
 wire \sbox_aesinv_inst.m4332245f/_0_ ;
 wire \sbox_aesinv_inst.m434a8cf5/_0_ ;
 wire \sbox_aesinv_inst.m43fecdd2/_0_ ;
 wire \sbox_aesinv_inst.m4638af86/_0_ ;
 wire \sbox_aesinv_inst.m4e5feeff/_0_ ;
 wire \sbox_aesinv_inst.m52c516d9/_0_ ;
 wire \sbox_aesinv_inst.m54eaa319/_0_ ;
 wire \sbox_aesinv_inst.m55775071/_0_ ;
 wire \sbox_aesinv_inst.m557f00ff/_0_ ;
 wire \sbox_aesinv_inst.m571fff3f/_0_ ;
 wire \sbox_aesinv_inst.m57ffff00/_0_ ;
 wire \sbox_aesinv_inst.m5a5f5b5f/_0_ ;
 wire \sbox_aesinv_inst.m5b847ba9/_0_ ;
 wire \sbox_aesinv_inst.m5e9f51e4/_0_ ;
 wire \sbox_aesinv_inst.m5fff0faf/_0_ ;
 wire \sbox_aesinv_inst.m6191ae47/_0_ ;
 wire \sbox_aesinv_inst.m6d287e63/_0_ ;
 wire \sbox_aesinv_inst.m7077f7ff/_0_ ;
 wire \sbox_aesinv_inst.m777717ff/_0_ ;
 wire \sbox_aesinv_inst.m77cd77ff/_0_ ;
 wire \sbox_aesinv_inst.m77ff3337/_0_ ;
 wire \sbox_aesinv_inst.m7847e6db/_0_ ;
 wire \sbox_aesinv_inst.m7c7c7c7d/_0_ ;
 wire \sbox_aesinv_inst.m7ca10f66/_0_ ;
 wire \sbox_aesinv_inst.m7f5f3300/_0_ ;
 wire \sbox_aesinv_inst.m854f7ef5/_0_ ;
 wire \sbox_aesinv_inst.m8ad2e815/_0_ ;
 wire \sbox_aesinv_inst.m8b30445b/_0_ ;
 wire \sbox_aesinv_inst.m8fdfffff/_0_ ;
 wire \sbox_aesinv_inst.m96492239/_0_ ;
 wire \sbox_aesinv_inst.ma0a0a1a1/_0_ ;
 wire \sbox_aesinv_inst.ma0fb7cd2/_0_ ;
 wire \sbox_aesinv_inst.ma1b3a5bf/_0_ ;
 wire \sbox_aesinv_inst.ma9e15289/_0_ ;
 wire \sbox_aesinv_inst.maa0faf5f/_0_ ;
 wire \sbox_aesinv_inst.maaaf153f/_0_ ;
 wire \sbox_aesinv_inst.maf7faf7f/_0_ ;
 wire \sbox_aesinv_inst.mb047c23f/_0_ ;
 wire \sbox_aesinv_inst.mb1b1f5f7/_0_ ;
 wire \sbox_aesinv_inst.mbb77ffff/_0_ ;
 wire \sbox_aesinv_inst.mbfbf373f/_0_ ;
 wire \sbox_aesinv_inst.mc3c3c3cf/_0_ ;
 wire \sbox_aesinv_inst.mc5cfc5df/_0_ ;
 wire \sbox_aesinv_inst.mc60b25d3/_0_ ;
 wire \sbox_aesinv_inst.mcccf030f/_0_ ;
 wire \sbox_aesinv_inst.mdd11cc00/_0_ ;
 wire \sbox_aesinv_inst.mdd7fff7f/_0_ ;
 wire \sbox_aesinv_inst.mdf77df77/_0_ ;
 wire \sbox_aesinv_inst.mdfdf77ff/_0_ ;
 wire \sbox_aesinv_inst.me3ab5bd2/_0_ ;
 wire \sbox_aesinv_inst.mf12405c2/_0_ ;
 wire \sbox_aesinv_inst.mf333f377/_0_ ;
 wire \sbox_aesinv_inst.mf33fffff/_0_ ;
 wire \sbox_aesinv_inst.mf35ff3ff/_0_ ;
 wire \sbox_aesinv_inst.mf3f37f7f/_0_ ;
 wire \sbox_aesinv_inst.mf555f57f/_0_ ;
 wire \sbox_aesinv_inst.mf5ff5fff/_0_ ;
 wire \sbox_aesinv_inst.mff010103/_0_ ;
 wire \sbox_aesinv_inst.mff05333f/_0_ ;
 wire \sbox_aesinv_inst.mff3f05ff/_0_ ;
 wire \sbox_aesinv_inst.mfff30000/_0_ ;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sg13g2_dfrbp_1 _16_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net6),
    .D(\sbox_aesinv_inst.x0 ),
    .Q_N(_01_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _17_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net7),
    .D(\sbox_aesinv_inst.x1 ),
    .Q_N(_02_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _18_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net8),
    .D(\sbox_aesinv_inst.x2 ),
    .Q_N(_03_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _19_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net9),
    .D(\sbox_aesinv_inst.x3 ),
    .Q_N(_04_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _20_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net10),
    .D(\sbox_aesinv_inst.x4 ),
    .Q_N(_05_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _21_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net11),
    .D(\sbox_aesinv_inst.x5 ),
    .Q_N(_06_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _22_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net4),
    .D(\sbox_aesinv_inst.x6 ),
    .Q_N(_07_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _23_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net5),
    .D(\sbox_aesinv_inst.x7 ),
    .Q_N(_00_),
    .Q(uio_out[7]));
 sg13g2_tiehi _23__5 (.L_HI(net5));
 sg13g2_tiehi _16__6 (.L_HI(net6));
 sg13g2_tiehi _17__7 (.L_HI(net7));
 sg13g2_tiehi _18__8 (.L_HI(net8));
 sg13g2_tiehi _19__9 (.L_HI(net9));
 sg13g2_tiehi _20__10 (.L_HI(net10));
 sg13g2_tiehi _21__11 (.L_HI(net11));
 sg13g2_tiehi tt_um_daosvik_aesinvsbox_12 (.L_HI(net12));
 sg13g2_tiehi tt_um_daosvik_aesinvsbox_13 (.L_HI(net13));
 sg13g2_tiehi tt_um_daosvik_aesinvsbox_14 (.L_HI(net14));
 sg13g2_tiehi tt_um_daosvik_aesinvsbox_15 (.L_HI(net15));
 sg13g2_tiehi tt_um_daosvik_aesinvsbox_16 (.L_HI(net16));
 sg13g2_tiehi tt_um_daosvik_aesinvsbox_17 (.L_HI(net17));
 sg13g2_tiehi tt_um_daosvik_aesinvsbox_18 (.L_HI(net18));
 sg13g2_tiehi tt_um_daosvik_aesinvsbox_19 (.L_HI(net19));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _40_ (.A(\sbox_aesinv_inst.x0 ),
    .X(uo_out[0]));
 sg13g2_buf_1 _41_ (.A(\sbox_aesinv_inst.x1 ),
    .X(uo_out[1]));
 sg13g2_buf_1 _42_ (.A(\sbox_aesinv_inst.x2 ),
    .X(uo_out[2]));
 sg13g2_buf_1 _43_ (.A(\sbox_aesinv_inst.x3 ),
    .X(uo_out[3]));
 sg13g2_buf_1 _44_ (.A(\sbox_aesinv_inst.x4 ),
    .X(uo_out[4]));
 sg13g2_buf_1 _45_ (.A(\sbox_aesinv_inst.x5 ),
    .X(uo_out[5]));
 sg13g2_buf_1 _46_ (.A(\sbox_aesinv_inst.x6 ),
    .X(uo_out[6]));
 sg13g2_buf_1 _47_ (.A(\sbox_aesinv_inst.x7 ),
    .X(uo_out[7]));
 sg13g2_nand4_1 \sbox_aesinv_inst.m0/_0_  (.B(\sbox_aesinv_inst.x0a ),
    .C(\sbox_aesinv_inst.x0c ),
    .A(\sbox_aesinv_inst.x0b ),
    .Y(\sbox_aesinv_inst.x0 ),
    .D(\sbox_aesinv_inst.x0d ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m00000008/_0_  (.A(\sbox_aesinv_inst.xfffffff0 ),
    .B_N(\sbox_aesinv_inst.xcc88cc88 ),
    .Y(\sbox_aesinv_inst.x00000008 ));
 sg13g2_nor2_1 \sbox_aesinv_inst.m00000013/_0_  (.A(\sbox_aesinv_inst.xffffffcc ),
    .B(\sbox_aesinv_inst.xf0f0a0a0 ),
    .Y(\sbox_aesinv_inst.x00000013 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m00000054/_0_  (.A(\sbox_aesinv_inst.xffffffaa ),
    .B_N(\sbox_aesinv_inst.xfffffcfc ),
    .Y(\sbox_aesinv_inst.x00000054 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m00000080/_0_  (.A(\sbox_aesinv_inst.xf0f0f000 ),
    .B_N(\sbox_aesinv_inst.x80808080 ),
    .Y(\sbox_aesinv_inst.x00000080 ));
 sg13g2_nor4_1 \sbox_aesinv_inst.m00000117/_0_  (.A(\sbox_aesinv_inst.xfc00fc00 ),
    .B(\sbox_aesinv_inst.xffff0000 ),
    .C(\sbox_aesinv_inst.xc8c8c8c8 ),
    .D(\sbox_aesinv_inst.xaaa0aaa0 ),
    .Y(\sbox_aesinv_inst.x00000117 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m00000550/_1_  (.X(\sbox_aesinv_inst.m00000550/_0_ ),
    .B(net296),
    .A(\sbox_aesinv_inst.xfffffafa ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00000550/_2_  (.B1(\sbox_aesinv_inst.m00000550/_0_ ),
    .Y(\sbox_aesinv_inst.x00000550 ),
    .A1(\sbox_aesinv_inst.xffffffaa ),
    .A2(net309));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m00001011/_0_  (.A1(net312),
    .A2(\sbox_aesinv_inst.xff00ff00 ),
    .Y(\sbox_aesinv_inst.x00001011 ),
    .B1(\sbox_aesinv_inst.xffffeeee ));
 sg13g2_or2_1 \sbox_aesinv_inst.m0000101a/_1_  (.X(\sbox_aesinv_inst.m0000101a/_0_ ),
    .B(net308),
    .A(\sbox_aesinv_inst.xffffeeee ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m0000101a/_2_  (.B1(\sbox_aesinv_inst.m0000101a/_0_ ),
    .Y(\sbox_aesinv_inst.x0000101a ),
    .A1(\sbox_aesinv_inst.xfffffff0 ),
    .A2(net333));
 sg13g2_or2_1 \sbox_aesinv_inst.m000010dc/_1_  (.X(\sbox_aesinv_inst.m000010dc/_0_ ),
    .B(net312),
    .A(\sbox_aesinv_inst.xffffeeee ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m000010dc/_2_  (.B1(\sbox_aesinv_inst.m000010dc/_0_ ),
    .Y(\sbox_aesinv_inst.x000010dc ),
    .A1(net261),
    .A2(net328));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m00001110/_0_  (.A(\sbox_aesinv_inst.xffffeeee ),
    .B_N(\sbox_aesinv_inst.xfff0fff0 ),
    .Y(\sbox_aesinv_inst.x00001110 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m00001175/_1_  (.X(\sbox_aesinv_inst.m00001175/_0_ ),
    .B(net304),
    .A(\sbox_aesinv_inst.xffffffcc ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00001175/_2_  (.B1(\sbox_aesinv_inst.m00001175/_0_ ),
    .Y(\sbox_aesinv_inst.x00001175 ),
    .A1(\sbox_aesinv_inst.xffffaaaa ),
    .A2(net262));
 sg13g2_or2_1 \sbox_aesinv_inst.m00001355/_1_  (.X(\sbox_aesinv_inst.m00001355/_0_ ),
    .B(net294),
    .A(\sbox_aesinv_inst.xfffffcfc ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00001355/_2_  (.B1(\sbox_aesinv_inst.m00001355/_0_ ),
    .Y(\sbox_aesinv_inst.x00001355 ),
    .A1(\sbox_aesinv_inst.xffffaaaa ),
    .A2(net262));
 sg13g2_and3_1 \sbox_aesinv_inst.m00008000/_0_  (.X(\sbox_aesinv_inst.x00008000 ),
    .A(net272),
    .B(\sbox_aesinv_inst.xf0f0f000 ),
    .C(net276));
 sg13g2_and3_1 \sbox_aesinv_inst.m00008880/_0_  (.X(\sbox_aesinv_inst.x00008880 ),
    .A(\sbox_aesinv_inst.xccc0ccc0 ),
    .B(\sbox_aesinv_inst.x88888888 ),
    .C(net285));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m0000a000/_0_  (.A(net259),
    .B_N(net269),
    .Y(\sbox_aesinv_inst.x0000a000 ));
 sg13g2_nor2_1 \sbox_aesinv_inst.m00010005/_0_  (.A(\sbox_aesinv_inst.xfffafffa ),
    .B(net260),
    .Y(\sbox_aesinv_inst.x00010005 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m00010031/_1_  (.X(\sbox_aesinv_inst.m00010031/_0_ ),
    .B(net313),
    .A(\sbox_aesinv_inst.xffffffcc ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00010031/_2_  (.B1(\sbox_aesinv_inst.m00010031/_0_ ),
    .Y(\sbox_aesinv_inst.x00010031 ),
    .A1(\sbox_aesinv_inst.xffeeffee ),
    .A2(net260));
 sg13g2_or2_1 \sbox_aesinv_inst.m00050011/_1_  (.X(\sbox_aesinv_inst.m00050011/_0_ ),
    .B(net281),
    .A(\sbox_aesinv_inst.xfffafffa ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00050011/_2_  (.B1(\sbox_aesinv_inst.m00050011/_0_ ),
    .Y(\sbox_aesinv_inst.x00050011 ),
    .A1(\sbox_aesinv_inst.xffeeffee ),
    .A2(net260));
 sg13g2_or2_1 \sbox_aesinv_inst.m00050022/_1_  (.X(\sbox_aesinv_inst.m00050022/_0_ ),
    .B(net281),
    .A(\sbox_aesinv_inst.xfffafffa ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00050022/_2_  (.B1(\sbox_aesinv_inst.m00050022/_0_ ),
    .Y(\sbox_aesinv_inst.x00050022 ),
    .A1(\sbox_aesinv_inst.xffffffcc ),
    .A2(net336));
 sg13g2_or2_1 \sbox_aesinv_inst.m00050300/_1_  (.X(\sbox_aesinv_inst.m00050300/_0_ ),
    .B(net278),
    .A(\sbox_aesinv_inst.xfffafffa ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00050300/_2_  (.B1(\sbox_aesinv_inst.m00050300/_0_ ),
    .Y(\sbox_aesinv_inst.x00050300 ),
    .A1(\sbox_aesinv_inst.xfffffcfc ),
    .A2(net294));
 sg13g2_or2_1 \sbox_aesinv_inst.m00060006/_1_  (.X(\sbox_aesinv_inst.m00060006/_0_ ),
    .B(net326),
    .A(\sbox_aesinv_inst.xfffafffa ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00060006/_2_  (.B1(\sbox_aesinv_inst.m00060006/_0_ ),
    .Y(\sbox_aesinv_inst.x00060006 ),
    .A1(\sbox_aesinv_inst.xfffcfffc ),
    .A2(net338));
 sg13g2_or2_1 \sbox_aesinv_inst.m00070013/_1_  (.X(\sbox_aesinv_inst.m00070013/_0_ ),
    .B(net281),
    .A(\sbox_aesinv_inst.xfffafffa ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00070013/_2_  (.B1(\sbox_aesinv_inst.m00070013/_0_ ),
    .Y(\sbox_aesinv_inst.x00070013 ),
    .A1(\sbox_aesinv_inst.xffccffcc ),
    .A2(\sbox_aesinv_inst.xf0f0a0a0 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m0007173f/_1_  (.B(\sbox_aesinv_inst.xfcccfccc ),
    .C(\sbox_aesinv_inst.xfffffff0 ),
    .A(\sbox_aesinv_inst.xeaeaeaea ),
    .Y(\sbox_aesinv_inst.m0007173f/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m0007173f/_2_  (.A(\sbox_aesinv_inst.xfff00000 ),
    .B_N(\sbox_aesinv_inst.m0007173f/_0_ ),
    .Y(\sbox_aesinv_inst.x0007173f ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m000a022a/_1_  (.B(\sbox_aesinv_inst.xfffffcfc ),
    .C(\sbox_aesinv_inst.xffffffcc ),
    .A(\sbox_aesinv_inst.xaaa0aaa0 ),
    .Y(\sbox_aesinv_inst.m000a022a/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m000a022a/_2_  (.A(net334),
    .B_N(\sbox_aesinv_inst.m000a022a/_0_ ),
    .Y(\sbox_aesinv_inst.x000a022a ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m000a0808/_0_  (.A(\sbox_aesinv_inst.xfff0f0f0 ),
    .B_N(\sbox_aesinv_inst.xaaaa8888 ),
    .Y(\sbox_aesinv_inst.x000a0808 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m000aaaab/_1_  (.X(\sbox_aesinv_inst.m000aaaab/_0_ ),
    .B(net333),
    .A(net257));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m000aaaab/_2_  (.B1(\sbox_aesinv_inst.m000aaaab/_0_ ),
    .Y(\sbox_aesinv_inst.x000aaaab ),
    .A1(\sbox_aesinv_inst.xfffffff0 ),
    .A2(\sbox_aesinv_inst.xfcfccccc ));
 sg13g2_nor2_1 \sbox_aesinv_inst.m000c0e5e/_0_  (.A(\sbox_aesinv_inst.xf1a1f1a1 ),
    .B(\sbox_aesinv_inst.xfff30000 ),
    .Y(\sbox_aesinv_inst.x000c0e5e ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m000ccc00/_0_  (.A(net257),
    .B_N(\sbox_aesinv_inst.xcccccc00 ),
    .Y(\sbox_aesinv_inst.x000ccc00 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m000f023f/_1_  (.X(\sbox_aesinv_inst.m000f023f/_0_ ),
    .B(net334),
    .A(\sbox_aesinv_inst.xfffffcfc ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m000f023f/_2_  (.B1(\sbox_aesinv_inst.m000f023f/_0_ ),
    .Y(\sbox_aesinv_inst.x000f023f ),
    .A1(\sbox_aesinv_inst.xff00ff00 ),
    .A2(\sbox_aesinv_inst.xf0f0c0c0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m00113035/_1_  (.X(\sbox_aesinv_inst.m00113035/_0_ ),
    .B(net312),
    .A(\sbox_aesinv_inst.xf0f0c0c0 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00113035/_2_  (.B1(\sbox_aesinv_inst.m00113035/_0_ ),
    .Y(\sbox_aesinv_inst.x00113035 ),
    .A1(\sbox_aesinv_inst.xffaaffaa ),
    .A2(\sbox_aesinv_inst.xccccc0c0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m00130f0f/_1_  (.X(\sbox_aesinv_inst.m00130f0f/_0_ ),
    .B(net281),
    .A(\sbox_aesinv_inst.xffeeffee ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00130f0f/_2_  (.B1(\sbox_aesinv_inst.m00130f0f/_0_ ),
    .Y(\sbox_aesinv_inst.x00130f0f ),
    .A1(\sbox_aesinv_inst.xfff0f0f0 ),
    .A2(net259));
 sg13g2_or2_1 \sbox_aesinv_inst.m00330404/_1_  (.X(\sbox_aesinv_inst.m00330404/_0_ ),
    .B(net282),
    .A(\sbox_aesinv_inst.xffcc0000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m00330404/_2_  (.B1(\sbox_aesinv_inst.m00330404/_0_ ),
    .Y(\sbox_aesinv_inst.x00330404 ),
    .A1(\sbox_aesinv_inst.xfffffafa ),
    .A2(net326));
 sg13g2_nor4_1 \sbox_aesinv_inst.m004000c0/_0_  (.A(\sbox_aesinv_inst.xf000f000 ),
    .B(net271),
    .C(net308),
    .D(net324),
    .Y(\sbox_aesinv_inst.x004000c0 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m005dccdd/_0_  (.B1(\sbox_aesinv_inst.xffaaffaa ),
    .Y(\sbox_aesinv_inst.x005dccdd ),
    .A1(net327),
    .A2(net257));
 sg13g2_or2_1 \sbox_aesinv_inst.m007fabff/_1_  (.X(\sbox_aesinv_inst.m007fabff/_0_ ),
    .B(net340),
    .A(net257));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m007fabff/_2_  (.B1(\sbox_aesinv_inst.m007fabff/_0_ ),
    .Y(\sbox_aesinv_inst.x007fabff ),
    .A1(\sbox_aesinv_inst.xff00f000 ),
    .A2(\sbox_aesinv_inst.xcc88cc88 ));
 sg13g2_and3_2 \sbox_aesinv_inst.m01/_0_  (.X(\sbox_aesinv_inst.x01 ),
    .A(net2),
    .B(net1),
    .C(net3));
 sg13g2_or2_1 \sbox_aesinv_inst.m0100011f/_1_  (.X(\sbox_aesinv_inst.m0100011f/_0_ ),
    .B(net293),
    .A(\sbox_aesinv_inst.xfefefefe ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m0100011f/_2_  (.B1(\sbox_aesinv_inst.m0100011f/_0_ ),
    .Y(\sbox_aesinv_inst.x0100011f ),
    .A1(\sbox_aesinv_inst.xffffff00 ),
    .A2(\sbox_aesinv_inst.xe0e0e0e0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m01010003/_1_  (.X(\sbox_aesinv_inst.m01010003/_0_ ),
    .B(net278),
    .A(\sbox_aesinv_inst.xfefefefe ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m01010003/_2_  (.B1(\sbox_aesinv_inst.m01010003/_0_ ),
    .Y(\sbox_aesinv_inst.x01010003 ),
    .A1(\sbox_aesinv_inst.xfffcfffc ),
    .A2(\sbox_aesinv_inst.xffaa0000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m01011010/_1_  (.X(\sbox_aesinv_inst.m01011010/_0_ ),
    .B(net278),
    .A(\sbox_aesinv_inst.xfefefefe ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m01011010/_2_  (.B1(\sbox_aesinv_inst.m01011010/_0_ ),
    .Y(\sbox_aesinv_inst.x01011010 ),
    .A1(\sbox_aesinv_inst.xffffeeee ),
    .A2(net308));
 sg13g2_or2_1 \sbox_aesinv_inst.m01155fff/_1_  (.X(\sbox_aesinv_inst.m01155fff/_0_ ),
    .B(\sbox_aesinv_inst.xeeee0000 ),
    .A(\sbox_aesinv_inst.xf000f000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m01155fff/_2_  (.B1(\sbox_aesinv_inst.m01155fff/_0_ ),
    .Y(\sbox_aesinv_inst.x01155fff ),
    .A1(\sbox_aesinv_inst.xff00aa00 ),
    .A2(\sbox_aesinv_inst.xfafa0000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m0133273f/_1_  (.X(\sbox_aesinv_inst.m0133273f/_0_ ),
    .B(net340),
    .A(\sbox_aesinv_inst.xaaaa8888 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m0133273f/_2_  (.B1(\sbox_aesinv_inst.m0133273f/_0_ ),
    .Y(\sbox_aesinv_inst.x0133273f ),
    .A1(\sbox_aesinv_inst.xfa00fa00 ),
    .A2(\sbox_aesinv_inst.xccccc0c0 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m0137133f/_1_  (.B(\sbox_aesinv_inst.xfffff0f0 ),
    .C(\sbox_aesinv_inst.xffccffcc ),
    .A(\sbox_aesinv_inst.xfafaaaaa ),
    .Y(\sbox_aesinv_inst.m0137133f/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m0137133f/_2_  (.A(\sbox_aesinv_inst.xccc0ccc0 ),
    .B_N(\sbox_aesinv_inst.m0137133f/_0_ ),
    .Y(\sbox_aesinv_inst.x0137133f ));
 sg13g2_or2_1 \sbox_aesinv_inst.m01f731f7/_1_  (.X(\sbox_aesinv_inst.m01f731f7/_0_ ),
    .B(net309),
    .A(net258));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m01f731f7/_2_  (.B1(\sbox_aesinv_inst.m01f731f7/_0_ ),
    .Y(\sbox_aesinv_inst.x01f731f7 ),
    .A1(\sbox_aesinv_inst.xfa00fa00 ),
    .A2(\sbox_aesinv_inst.xcc88cc88 ));
 sg13g2_nand2_1 \sbox_aesinv_inst.m02/_1_  (.Y(\sbox_aesinv_inst.m02/_0_ ),
    .A(net2),
    .B(net3));
 sg13g2_nor2_2 \sbox_aesinv_inst.m02/_2_  (.A(net1),
    .B(\sbox_aesinv_inst.m02/_0_ ),
    .Y(\sbox_aesinv_inst.x02 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m03fc03fc/_0_  (.A(\sbox_aesinv_inst.xfc00fc00 ),
    .B_N(\sbox_aesinv_inst.xfffcfffc ),
    .Y(\sbox_aesinv_inst.x03fc03fc ));
 sg13g2_nand2_1 \sbox_aesinv_inst.m04/_1_  (.Y(\sbox_aesinv_inst.m04/_0_ ),
    .A(net1),
    .B(net3));
 sg13g2_nor2_2 \sbox_aesinv_inst.m04/_2_  (.A(net2),
    .B(\sbox_aesinv_inst.m04/_0_ ),
    .Y(\sbox_aesinv_inst.x04 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m04044447/_1_  (.X(\sbox_aesinv_inst.m04044447/_0_ ),
    .B(net326),
    .A(\sbox_aesinv_inst.xfafaaaaa ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m04044447/_2_  (.B1(\sbox_aesinv_inst.m04044447/_0_ ),
    .Y(\sbox_aesinv_inst.x04044447 ),
    .A1(\sbox_aesinv_inst.xfffffff0 ),
    .A2(\sbox_aesinv_inst.xcc88cc88 ));
 sg13g2_nor4_1 \sbox_aesinv_inst.m040c0000/_0_  (.A(net267),
    .B(net265),
    .C(net322),
    .D(net279),
    .Y(\sbox_aesinv_inst.x040c0000 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m05500000/_0_  (.A(\sbox_aesinv_inst.xfaaafaaa ),
    .B_N(net257),
    .Y(\sbox_aesinv_inst.x05500000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m055f0557/_1_  (.X(\sbox_aesinv_inst.m055f0557/_0_ ),
    .B(net284),
    .A(\sbox_aesinv_inst.xfff00000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m055f0557/_2_  (.B1(\sbox_aesinv_inst.m055f0557/_0_ ),
    .Y(\sbox_aesinv_inst.x055f0557 ),
    .A1(\sbox_aesinv_inst.xfa00fa00 ),
    .A2(\sbox_aesinv_inst.xa8a8a8a8 ));
 sg13g2_inv_1 \sbox_aesinv_inst.m08/_1_  (.Y(\sbox_aesinv_inst.m08/_0_ ),
    .A(net3));
 sg13g2_nor3_2 \sbox_aesinv_inst.m08/_2_  (.A(\sbox_aesinv_inst.m08/_0_ ),
    .B(net1),
    .C(net2),
    .Y(\sbox_aesinv_inst.x08 ));
 sg13g2_and3_1 \sbox_aesinv_inst.m08000000/_0_  (.X(\sbox_aesinv_inst.x08000000 ),
    .A(net267),
    .B(net260),
    .C(net315));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m0a/_0_  (.Y(\sbox_aesinv_inst.x0a ),
    .B1(\sbox_aesinv_inst.x4332245f ),
    .B2(\sbox_aesinv_inst.x40 ),
    .A2(\sbox_aesinv_inst.x80 ),
    .A1(\sbox_aesinv_inst.x52af6f23 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m0a000000/_0_  (.A(\sbox_aesinv_inst.xf0f00000 ),
    .B_N(net267),
    .Y(\sbox_aesinv_inst.x0a000000 ));
 sg13g2_and3_1 \sbox_aesinv_inst.m0a080000/_0_  (.X(\sbox_aesinv_inst.x0a080000 ),
    .A(\sbox_aesinv_inst.xffcc0000 ),
    .B(\sbox_aesinv_inst.xaaaa0000 ),
    .C(net311));
 sg13g2_nand3_1 \sbox_aesinv_inst.m0abf1bbf/_1_  (.B(\sbox_aesinv_inst.xffcccccc ),
    .C(\sbox_aesinv_inst.xfff0fff0 ),
    .A(net342),
    .Y(\sbox_aesinv_inst.m0abf1bbf/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m0abf1bbf/_2_  (.A(net270),
    .B_N(\sbox_aesinv_inst.m0abf1bbf/_0_ ),
    .Y(\sbox_aesinv_inst.x0abf1bbf ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m0b/_0_  (.Y(\sbox_aesinv_inst.x0b ),
    .B1(\sbox_aesinv_inst.x229616fd ),
    .B2(\sbox_aesinv_inst.x10 ),
    .A2(\sbox_aesinv_inst.x20 ),
    .A1(\sbox_aesinv_inst.x000c0e5e ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m0b1fafbf/_1_  (.B(\sbox_aesinv_inst.xfcccfccc ),
    .C(net332),
    .A(\sbox_aesinv_inst.xfff0f0f0 ),
    .Y(\sbox_aesinv_inst.m0b1fafbf/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m0b1fafbf/_2_  (.A(net268),
    .B_N(\sbox_aesinv_inst.m0b1fafbf/_0_ ),
    .Y(\sbox_aesinv_inst.x0b1fafbf ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m0c/_0_  (.Y(\sbox_aesinv_inst.x0c ),
    .B1(\sbox_aesinv_inst.xdfc11244 ),
    .B2(\sbox_aesinv_inst.x04 ),
    .A2(\sbox_aesinv_inst.x08 ),
    .A1(\sbox_aesinv_inst.x7ca10f66 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m0cd37660/_0_  (.A1(\sbox_aesinv_inst.xf33fffff ),
    .A2(\sbox_aesinv_inst.xffec8888 ),
    .Y(\sbox_aesinv_inst.x0cd37660 ),
    .B1(\sbox_aesinv_inst.x00000117 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m0d/_0_  (.Y(\sbox_aesinv_inst.x0d ),
    .B1(\sbox_aesinv_inst.x326fc4dd ),
    .B2(\sbox_aesinv_inst.x01 ),
    .A2(\sbox_aesinv_inst.x02 ),
    .A1(\sbox_aesinv_inst.xd7997ddd ));
 sg13g2_and3_1 \sbox_aesinv_inst.m0e0a0000/_0_  (.X(\sbox_aesinv_inst.x0e0a0000 ),
    .A(\sbox_aesinv_inst.xeeee0000 ),
    .B(\sbox_aesinv_inst.xffaa0000 ),
    .C(net308));
 sg13g2_inv_1 \sbox_aesinv_inst.m0eb6ef2f/_1_  (.Y(\sbox_aesinv_inst.m0eb6ef2f/_0_ ),
    .A(\sbox_aesinv_inst.x0ff7ffff ));
 sg13g2_nor3_1 \sbox_aesinv_inst.m0eb6ef2f/_2_  (.A(\sbox_aesinv_inst.m0eb6ef2f/_0_ ),
    .B(\sbox_aesinv_inst.x01011010 ),
    .C(\sbox_aesinv_inst.x004000c0 ),
    .Y(\sbox_aesinv_inst.x0eb6ef2f ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m0f5f0a5f/_1_  (.B(net332),
    .C(net276),
    .A(\sbox_aesinv_inst.xff00ff00 ),
    .Y(\sbox_aesinv_inst.m0f5f0a5f/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m0f5f0a5f/_2_  (.A(\sbox_aesinv_inst.xf0a0f0a0 ),
    .B_N(\sbox_aesinv_inst.m0f5f0a5f/_0_ ),
    .Y(\sbox_aesinv_inst.x0f5f0a5f ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m0ff7ffff/_1_  (.B(net271),
    .C(net308),
    .A(net295),
    .Y(\sbox_aesinv_inst.m0ff7ffff/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m0ff7ffff/_2_  (.A(\sbox_aesinv_inst.xf0000000 ),
    .B_N(\sbox_aesinv_inst.m0ff7ffff/_0_ ),
    .Y(\sbox_aesinv_inst.x0ff7ffff ));
 sg13g2_nand4_1 \sbox_aesinv_inst.m1/_0_  (.B(\sbox_aesinv_inst.x1a ),
    .C(\sbox_aesinv_inst.x1c ),
    .A(\sbox_aesinv_inst.x1b ),
    .Y(\sbox_aesinv_inst.x1 ),
    .D(\sbox_aesinv_inst.x1d ));
 sg13g2_nand2_1 \sbox_aesinv_inst.m10/_1_  (.Y(\sbox_aesinv_inst.m10/_0_ ),
    .A(net1),
    .B(net2));
 sg13g2_nor2_2 \sbox_aesinv_inst.m10/_2_  (.A(net3),
    .B(\sbox_aesinv_inst.m10/_0_ ),
    .Y(\sbox_aesinv_inst.x10 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m10104040/_0_  (.A(\sbox_aesinv_inst.xeeeeaaaa ),
    .B_N(\sbox_aesinv_inst.xf0f0c0c0 ),
    .Y(\sbox_aesinv_inst.x10104040 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m11004400/_0_  (.A(\sbox_aesinv_inst.xeeeeaaaa ),
    .B_N(net258),
    .Y(\sbox_aesinv_inst.x11004400 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m11131313/_0_  (.A1(\sbox_aesinv_inst.xeeeeeeee ),
    .A2(\sbox_aesinv_inst.xfcfcfcfc ),
    .Y(\sbox_aesinv_inst.x11131313 ),
    .B1(\sbox_aesinv_inst.xaa000000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m11771333/_1_  (.X(\sbox_aesinv_inst.m11771333/_0_ ),
    .B(net285),
    .A(\sbox_aesinv_inst.xeeaaeeaa ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m11771333/_2_  (.B1(\sbox_aesinv_inst.m11771333/_0_ ),
    .Y(\sbox_aesinv_inst.x11771333 ),
    .A1(\sbox_aesinv_inst.xffcccccc ),
    .A2(net270));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m11aa0000/_0_  (.A(\sbox_aesinv_inst.xee00ee00 ),
    .B_N(\sbox_aesinv_inst.xffaa0000 ),
    .Y(\sbox_aesinv_inst.x11aa0000 ));
 sg13g2_a21o_1 \sbox_aesinv_inst.m12bf5b4f/_0_  (.A2(\sbox_aesinv_inst.x33ffff0f ),
    .A1(\sbox_aesinv_inst.x0abf1bbf ),
    .B1(\sbox_aesinv_inst.x10104040 ),
    .X(\sbox_aesinv_inst.x12bf5b4f ));
 sg13g2_or2_1 \sbox_aesinv_inst.m131317df/_1_  (.X(\sbox_aesinv_inst.m131317df/_0_ ),
    .B(net324),
    .A(\sbox_aesinv_inst.xcccccc00 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m131317df/_2_  (.B1(\sbox_aesinv_inst.m131317df/_0_ ),
    .Y(\sbox_aesinv_inst.x131317df ),
    .A1(\sbox_aesinv_inst.xe0e0e0e0 ),
    .A2(\sbox_aesinv_inst.xcccc8888 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m1333131f/_1_  (.X(\sbox_aesinv_inst.m1333131f/_0_ ),
    .B(net282),
    .A(\sbox_aesinv_inst.xffcc0000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m1333131f/_2_  (.B1(\sbox_aesinv_inst.m1333131f/_0_ ),
    .Y(\sbox_aesinv_inst.x1333131f ),
    .A1(\sbox_aesinv_inst.xe0e0e0e0 ),
    .A2(net261));
 sg13g2_or2_1 \sbox_aesinv_inst.m135f5fdf/_1_  (.X(\sbox_aesinv_inst.m135f5fdf/_0_ ),
    .B(net319),
    .A(net261));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m135f5fdf/_2_  (.B1(\sbox_aesinv_inst.m135f5fdf/_0_ ),
    .Y(\sbox_aesinv_inst.x135f5fdf ),
    .A1(net263),
    .A2(\sbox_aesinv_inst.xa0a0a0a0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m13bfbfbf/_1_  (.X(\sbox_aesinv_inst.m13bfbfbf/_0_ ),
    .B(net335),
    .A(\sbox_aesinv_inst.xff000000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m13bfbfbf/_2_  (.B1(\sbox_aesinv_inst.m13bfbfbf/_0_ ),
    .Y(\sbox_aesinv_inst.x13bfbfbf ),
    .A1(\sbox_aesinv_inst.xe0e0e0e0 ),
    .A2(net264));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m15000400/_0_  (.A(\sbox_aesinv_inst.xeaeaeaea ),
    .B_N(net258),
    .Y(\sbox_aesinv_inst.x15000400 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m151d777f/_1_  (.X(\sbox_aesinv_inst.m151d777f/_0_ ),
    .B(net326),
    .A(\sbox_aesinv_inst.xccc0ccc0 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m151d777f/_2_  (.B1(\sbox_aesinv_inst.m151d777f/_0_ ),
    .Y(\sbox_aesinv_inst.x151d777f ),
    .A1(net266),
    .A2(\sbox_aesinv_inst.xaaaa8888 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m15555050/_1_  (.X(\sbox_aesinv_inst.m15555050/_0_ ),
    .B(net286),
    .A(\sbox_aesinv_inst.xfaaafaaa ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m15555050/_2_  (.B1(\sbox_aesinv_inst.m15555050/_0_ ),
    .Y(\sbox_aesinv_inst.x15555050 ),
    .A1(\sbox_aesinv_inst.xeeeeaaaa ),
    .A2(net313));
 sg13g2_nand3_1 \sbox_aesinv_inst.m169287dc/_1_  (.B(\sbox_aesinv_inst.xfcfcf8a0 ),
    .C(\sbox_aesinv_inst.xeaefffff ),
    .A(\sbox_aesinv_inst.xff7f7f7f ),
    .Y(\sbox_aesinv_inst.m169287dc/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m169287dc/_2_  (.A(\sbox_aesinv_inst.x01010003 ),
    .B_N(\sbox_aesinv_inst.m169287dc/_0_ ),
    .Y(\sbox_aesinv_inst.x169287dc ));
 sg13g2_or2_1 \sbox_aesinv_inst.m175f333f/_1_  (.X(\sbox_aesinv_inst.m175f333f/_0_ ),
    .B(net286),
    .A(\sbox_aesinv_inst.xfaaafaaa ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m175f333f/_2_  (.B1(\sbox_aesinv_inst.m175f333f/_0_ ),
    .Y(\sbox_aesinv_inst.x175f333f ),
    .A1(\sbox_aesinv_inst.xccc0ccc0 ),
    .A2(\sbox_aesinv_inst.xa0a00000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m17ff555f/_1_  (.X(\sbox_aesinv_inst.m17ff555f/_0_ ),
    .B(net280),
    .A(\sbox_aesinv_inst.xfc00fc00 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m17ff555f/_2_  (.B1(\sbox_aesinv_inst.m17ff555f/_0_ ),
    .Y(\sbox_aesinv_inst.x17ff555f ),
    .A1(net265),
    .A2(\sbox_aesinv_inst.xaaa0aaa0 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m1a/_0_  (.Y(\sbox_aesinv_inst.x1a ),
    .B1(\sbox_aesinv_inst.x5e9f51e4 ),
    .B2(\sbox_aesinv_inst.x40 ),
    .A2(\sbox_aesinv_inst.x80 ),
    .A1(\sbox_aesinv_inst.xa4b75f65 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m1a10b72b/_1_  (.B(\sbox_aesinv_inst.xfffff8a0 ),
    .C(\sbox_aesinv_inst.xf5ff5fff ),
    .A(\sbox_aesinv_inst.xefefcf8f ),
    .Y(\sbox_aesinv_inst.m1a10b72b/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m1a10b72b/_2_  (.A(\sbox_aesinv_inst.x00000054 ),
    .B_N(\sbox_aesinv_inst.m1a10b72b/_0_ ),
    .Y(\sbox_aesinv_inst.x1a10b72b ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m1b/_0_  (.Y(\sbox_aesinv_inst.x1b ),
    .B1(\sbox_aesinv_inst.x23853f57 ),
    .B2(\sbox_aesinv_inst.x10 ),
    .A2(\sbox_aesinv_inst.x20 ),
    .A1(\sbox_aesinv_inst.xa90301b8 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m1c/_0_  (.Y(\sbox_aesinv_inst.x1c ),
    .B1(\sbox_aesinv_inst.xa0fb7cd2 ),
    .B2(\sbox_aesinv_inst.x04 ),
    .A2(\sbox_aesinv_inst.x08 ),
    .A1(\sbox_aesinv_inst.x8df398a3 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m1d/_0_  (.Y(\sbox_aesinv_inst.x1d ),
    .B1(\sbox_aesinv_inst.x2c6cdf10 ),
    .B2(\sbox_aesinv_inst.x01 ),
    .A2(\sbox_aesinv_inst.x02 ),
    .A1(\sbox_aesinv_inst.x96492239 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m1d7f5dff/_1_  (.X(\sbox_aesinv_inst.m1d7f5dff/_0_ ),
    .B(net324),
    .A(\sbox_aesinv_inst.xf0f0a0a0 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m1d7f5dff/_2_  (.B1(\sbox_aesinv_inst.m1d7f5dff/_0_ ),
    .Y(\sbox_aesinv_inst.x1d7f5dff ),
    .A1(\sbox_aesinv_inst.xee00ee00 ),
    .A2(net271));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m1f7b28d7/_0_  (.A1(\sbox_aesinv_inst.xffecffa8 ),
    .A2(\sbox_aesinv_inst.x0007173f ),
    .Y(\sbox_aesinv_inst.x1f7b28d7 ),
    .B1(\sbox_aesinv_inst.xe080c000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m1f7f55ff/_1_  (.X(\sbox_aesinv_inst.m1f7f55ff/_0_ ),
    .B(net288),
    .A(\sbox_aesinv_inst.xe0e0e0e0 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m1f7f55ff/_2_  (.B1(\sbox_aesinv_inst.m1f7f55ff/_0_ ),
    .Y(\sbox_aesinv_inst.x1f7f55ff ),
    .A1(\sbox_aesinv_inst.xff00aa00 ),
    .A2(\sbox_aesinv_inst.x88880000 ));
 sg13g2_nand4_1 \sbox_aesinv_inst.m2/_0_  (.B(\sbox_aesinv_inst.x2a ),
    .C(\sbox_aesinv_inst.x2c ),
    .A(\sbox_aesinv_inst.x2b ),
    .Y(\sbox_aesinv_inst.x2 ),
    .D(\sbox_aesinv_inst.x2d ));
 sg13g2_inv_1 \sbox_aesinv_inst.m20/_1_  (.Y(\sbox_aesinv_inst.m20/_0_ ),
    .A(net2));
 sg13g2_nor3_2 \sbox_aesinv_inst.m20/_2_  (.A(\sbox_aesinv_inst.m20/_0_ ),
    .B(net1),
    .C(net3),
    .Y(\sbox_aesinv_inst.x20 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m229616fd/_1_  (.X(\sbox_aesinv_inst.m229616fd/_0_ ),
    .B(\sbox_aesinv_inst.xe8e8e800 ),
    .A(\sbox_aesinv_inst.xff010103 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m229616fd/_2_  (.B(\sbox_aesinv_inst.xffffffaa ),
    .C(\sbox_aesinv_inst.m229616fd/_0_ ),
    .A(\sbox_aesinv_inst.xdd7fff7f ),
    .Y(\sbox_aesinv_inst.x229616fd ));
 sg13g2_a221oi_1 \sbox_aesinv_inst.m23369e29/_0_  (.B2(\sbox_aesinv_inst.xf0c0f5d5 ),
    .C1(\sbox_aesinv_inst.xcc880000 ),
    .B1(\sbox_aesinv_inst.x03fc03fc ),
    .A1(\sbox_aesinv_inst.x55556666 ),
    .Y(\sbox_aesinv_inst.x23369e29 ),
    .A2(\sbox_aesinv_inst.xf003f003 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m23853f57/_0_  (.A1(\sbox_aesinv_inst.x557f00ff ),
    .A2(\sbox_aesinv_inst.xfefaeca8 ),
    .Y(\sbox_aesinv_inst.x23853f57 ),
    .B1(\sbox_aesinv_inst.xc800c000 ));
 sg13g2_inv_1 \sbox_aesinv_inst.m24cc4461/_1_  (.Y(\sbox_aesinv_inst.m24cc4461/_0_ ),
    .A(\sbox_aesinv_inst.x37ff5577 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m24cc4461/_2_  (.A1(\sbox_aesinv_inst.xfffffffe ),
    .A2(\sbox_aesinv_inst.x1333131f ),
    .Y(\sbox_aesinv_inst.x24cc4461 ),
    .B1(\sbox_aesinv_inst.m24cc4461/_0_ ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m2a/_0_  (.Y(\sbox_aesinv_inst.x2a ),
    .B1(\sbox_aesinv_inst.xa9e15289 ),
    .B2(\sbox_aesinv_inst.x40 ),
    .A2(\sbox_aesinv_inst.x80 ),
    .A1(\sbox_aesinv_inst.x169287dc ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m2a000000/_0_  (.A(net266),
    .B_N(net267),
    .Y(\sbox_aesinv_inst.x2a000000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m2aeeaaee/_1_  (.X(\sbox_aesinv_inst.m2aeeaaee/_0_ ),
    .B(net329),
    .A(\sbox_aesinv_inst.xcc00cc00 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m2aeeaaee/_2_  (.B1(\sbox_aesinv_inst.m2aeeaaee/_0_ ),
    .Y(\sbox_aesinv_inst.x2aeeaaee ),
    .A1(\sbox_aesinv_inst.xc0c00000 ),
    .A2(net338));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m2b/_0_  (.Y(\sbox_aesinv_inst.x2b ),
    .B1(\sbox_aesinv_inst.x0cd37660 ),
    .B2(\sbox_aesinv_inst.x10 ),
    .A2(\sbox_aesinv_inst.x20 ),
    .A1(\sbox_aesinv_inst.x39fe8cff ));
 sg13g2_or2_1 \sbox_aesinv_inst.m2bffafff/_1_  (.X(\sbox_aesinv_inst.m2bffafff/_0_ ),
    .B(net336),
    .A(net266));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m2bffafff/_2_  (.B1(\sbox_aesinv_inst.m2bffafff/_0_ ),
    .Y(\sbox_aesinv_inst.x2bffafff ),
    .A1(\sbox_aesinv_inst.xf000f000 ),
    .A2(net264));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m2c/_0_  (.Y(\sbox_aesinv_inst.x2c ),
    .B1(\sbox_aesinv_inst.x8ad2e815 ),
    .B2(\sbox_aesinv_inst.x04 ),
    .A2(\sbox_aesinv_inst.x08 ),
    .A1(\sbox_aesinv_inst.x0eb6ef2f ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m2c6cdf10/_0_  (.B1(\sbox_aesinv_inst.xdfdf77ff ),
    .Y(\sbox_aesinv_inst.x2c6cdf10 ),
    .A1(\sbox_aesinv_inst.x333300cf ),
    .A2(\sbox_aesinv_inst.xf0a0a0a0 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m2ca62526/_0_  (.A1(\sbox_aesinv_inst.x135f5fdf ),
    .A2(\sbox_aesinv_inst.xfff8fac8 ),
    .Y(\sbox_aesinv_inst.x2ca62526 ),
    .B1(\sbox_aesinv_inst.xc011c011 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m2d/_0_  (.Y(\sbox_aesinv_inst.x2d ),
    .B1(\sbox_aesinv_inst.x1a10b72b ),
    .B2(\sbox_aesinv_inst.x01 ),
    .A2(\sbox_aesinv_inst.x02 ),
    .A1(\sbox_aesinv_inst.xc60b25d3 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m2d9fb2de/_1_  (.X(\sbox_aesinv_inst.m2d9fb2de/_0_ ),
    .B(\sbox_aesinv_inst.xfecccc00 ),
    .A(\sbox_aesinv_inst.xa0a0a1a1 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m2d9fb2de/_2_  (.B(\sbox_aesinv_inst.xf3f37f7f ),
    .C(\sbox_aesinv_inst.m2d9fb2de/_0_ ),
    .A(\sbox_aesinv_inst.xdf77df77 ),
    .Y(\sbox_aesinv_inst.x2d9fb2de ));
 sg13g2_inv_1 \sbox_aesinv_inst.m2fa5e682/_1_  (.Y(\sbox_aesinv_inst.m2fa5e682/_0_ ),
    .A(\sbox_aesinv_inst.x2fafffff ));
 sg13g2_nor3_1 \sbox_aesinv_inst.m2fa5e682/_2_  (.A(\sbox_aesinv_inst.m2fa5e682/_0_ ),
    .B(\sbox_aesinv_inst.x000a0808 ),
    .C(\sbox_aesinv_inst.x00001175 ),
    .Y(\sbox_aesinv_inst.x2fa5e682 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m2fafffff/_0_  (.B1(\sbox_aesinv_inst.xf0f00000 ),
    .Y(\sbox_aesinv_inst.x2fafffff ),
    .A1(net331),
    .A2(net263));
 sg13g2_nand4_1 \sbox_aesinv_inst.m3/_0_  (.B(\sbox_aesinv_inst.x3a ),
    .C(\sbox_aesinv_inst.x3c ),
    .A(\sbox_aesinv_inst.x3b ),
    .Y(\sbox_aesinv_inst.x3 ),
    .D(\sbox_aesinv_inst.x3d ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m30307000/_0_  (.A(\sbox_aesinv_inst.xcccc8888 ),
    .B_N(\sbox_aesinv_inst.xf0f0f000 ),
    .Y(\sbox_aesinv_inst.x30307000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m3030f1f0/_1_  (.X(\sbox_aesinv_inst.m3030f1f0/_0_ ),
    .B(net301),
    .A(\sbox_aesinv_inst.xffffeeee ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m3030f1f0/_2_  (.B1(\sbox_aesinv_inst.m3030f1f0/_0_ ),
    .Y(\sbox_aesinv_inst.x3030f1f0 ),
    .A1(\sbox_aesinv_inst.xc0c00000 ),
    .A2(net312));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m30c030c0/_0_  (.A(net262),
    .B_N(\sbox_aesinv_inst.xf0c0f0c0 ),
    .Y(\sbox_aesinv_inst.x30c030c0 ));
 sg13g2_nor3_1 \sbox_aesinv_inst.m318ab4e1/_1_  (.A(\sbox_aesinv_inst.x30c030c0 ),
    .B(\sbox_aesinv_inst.x15000400 ),
    .C(\sbox_aesinv_inst.x000aaaab ),
    .Y(\sbox_aesinv_inst.m318ab4e1/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m318ab4e1/_2_  (.A(\sbox_aesinv_inst.m318ab4e1/_0_ ),
    .B_N(\sbox_aesinv_inst.xbbbbf5f5 ),
    .Y(\sbox_aesinv_inst.x318ab4e1 ));
 sg13g2_and3_1 \sbox_aesinv_inst.m32220000/_0_  (.X(\sbox_aesinv_inst.x32220000 ),
    .A(\sbox_aesinv_inst.xfafa0000 ),
    .B(\sbox_aesinv_inst.xffaa0000 ),
    .C(net328));
 sg13g2_and3_1 \sbox_aesinv_inst.m32302020/_0_  (.X(\sbox_aesinv_inst.x32302020 ),
    .A(\sbox_aesinv_inst.xfafaaaaa ),
    .B(\sbox_aesinv_inst.xfff0f0f0 ),
    .C(net320));
 sg13g2_nand3_1 \sbox_aesinv_inst.m323233fb/_1_  (.B(\sbox_aesinv_inst.xffffcccc ),
    .C(net312),
    .A(net342),
    .Y(\sbox_aesinv_inst.m323233fb/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m323233fb/_2_  (.A(net261),
    .B_N(\sbox_aesinv_inst.m323233fb/_0_ ),
    .Y(\sbox_aesinv_inst.x323233fb ));
 sg13g2_a21o_1 \sbox_aesinv_inst.m326fc4dd/_0_  (.A2(\sbox_aesinv_inst.x005dccdd ),
    .A1(\sbox_aesinv_inst.xc5cfc5df ),
    .B1(\sbox_aesinv_inst.x32220000 ),
    .X(\sbox_aesinv_inst.x326fc4dd ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m333300cf/_1_  (.B(net327),
    .C(net286),
    .A(\sbox_aesinv_inst.xfff0fff0 ),
    .Y(\sbox_aesinv_inst.m333300cf/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m333300cf/_2_  (.A(net261),
    .B_N(\sbox_aesinv_inst.m333300cf/_0_ ),
    .Y(\sbox_aesinv_inst.x333300cf ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m33cfffff/_1_  (.B(net259),
    .C(net326),
    .A(net296),
    .Y(\sbox_aesinv_inst.m33cfffff/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m33cfffff/_2_  (.A(net263),
    .B_N(\sbox_aesinv_inst.m33cfffff/_0_ ),
    .Y(\sbox_aesinv_inst.x33cfffff ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m33ffff0f/_1_  (.B(\sbox_aesinv_inst.xfffff0f0 ),
    .C(net283),
    .A(net299),
    .Y(\sbox_aesinv_inst.m33ffff0f/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m33ffff0f/_2_  (.A(net263),
    .B_N(\sbox_aesinv_inst.m33ffff0f/_0_ ),
    .Y(\sbox_aesinv_inst.x33ffff0f ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m37303733/_1_  (.B(\sbox_aesinv_inst.xffffcccc ),
    .C(net312),
    .A(net301),
    .Y(\sbox_aesinv_inst.m37303733/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m37303733/_2_  (.A(\sbox_aesinv_inst.xc8c8c8c8 ),
    .B_N(\sbox_aesinv_inst.m37303733/_0_ ),
    .Y(\sbox_aesinv_inst.x37303733 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m3777053f/_1_  (.X(\sbox_aesinv_inst.m3777053f/_0_ ),
    .B(net275),
    .A(\sbox_aesinv_inst.xcc88cc88 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m3777053f/_2_  (.B1(\sbox_aesinv_inst.m3777053f/_0_ ),
    .Y(\sbox_aesinv_inst.x3777053f ),
    .A1(\sbox_aesinv_inst.xf0c0f0c0 ),
    .A2(\sbox_aesinv_inst.xaaaaaa00 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m37ff5577/_1_  (.X(\sbox_aesinv_inst.m37ff5577/_0_ ),
    .B(net283),
    .A(net263));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m37ff5577/_2_  (.B1(\sbox_aesinv_inst.m37ff5577/_0_ ),
    .Y(\sbox_aesinv_inst.x37ff5577 ),
    .A1(\sbox_aesinv_inst.xc0c00000 ),
    .A2(\sbox_aesinv_inst.xaa88aa88 ));
 sg13g2_a21o_1 \sbox_aesinv_inst.m39fe8cff/_0_  (.A2(\sbox_aesinv_inst.xfcfcccff ),
    .A1(\sbox_aesinv_inst.x2bffafff ),
    .B1(\sbox_aesinv_inst.x11aa0000 ),
    .X(\sbox_aesinv_inst.x39fe8cff ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m3a/_0_  (.Y(\sbox_aesinv_inst.x3a ),
    .B1(\sbox_aesinv_inst.x41d5cc5c ),
    .B2(\sbox_aesinv_inst.x40 ),
    .A2(\sbox_aesinv_inst.x80 ),
    .A1(\sbox_aesinv_inst.x6191ae47 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m3b/_0_  (.Y(\sbox_aesinv_inst.x3b ),
    .B1(\sbox_aesinv_inst.x6d287e63 ),
    .B2(\sbox_aesinv_inst.x10 ),
    .A2(\sbox_aesinv_inst.x20 ),
    .A1(\sbox_aesinv_inst.x4638af86 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m3c/_0_  (.Y(\sbox_aesinv_inst.x3c ),
    .B1(\sbox_aesinv_inst.x2d9fb2de ),
    .B2(\sbox_aesinv_inst.x04 ),
    .A2(\sbox_aesinv_inst.x08 ),
    .A1(\sbox_aesinv_inst.x8b30445b ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m3c3ffdff/_1_  (.B(\sbox_aesinv_inst.xff00aa00 ),
    .C(net322),
    .A(net307),
    .Y(\sbox_aesinv_inst.m3c3ffdff/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m3c3ffdff/_2_  (.A(net265),
    .B_N(\sbox_aesinv_inst.m3c3ffdff/_0_ ),
    .Y(\sbox_aesinv_inst.x3c3ffdff ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m3cf25843/_1_  (.B(\sbox_aesinv_inst.x0b1fafbf ),
    .C(\sbox_aesinv_inst.x77cd77ff ),
    .A(\sbox_aesinv_inst.xfffffffc ),
    .Y(\sbox_aesinv_inst.m3cf25843/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m3cf25843/_2_  (.A(\sbox_aesinv_inst.xc0008000 ),
    .B_N(\sbox_aesinv_inst.m3cf25843/_0_ ),
    .Y(\sbox_aesinv_inst.x3cf25843 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m3d/_0_  (.Y(\sbox_aesinv_inst.x3d ),
    .B1(\sbox_aesinv_inst.x3cf25843 ),
    .B2(\sbox_aesinv_inst.x01 ),
    .A2(\sbox_aesinv_inst.x02 ),
    .A1(\sbox_aesinv_inst.xe8133bb7 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m3f00ff05/_0_  (.A1(\sbox_aesinv_inst.xfffffafa ),
    .A2(net296),
    .Y(\sbox_aesinv_inst.x3f00ff05 ),
    .B1(net266));
 sg13g2_nand3_1 \sbox_aesinv_inst.m3f0fffcf/_1_  (.B(\sbox_aesinv_inst.xf0f0f0f0 ),
    .C(net319),
    .A(net292),
    .Y(\sbox_aesinv_inst.m3f0fffcf/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m3f0fffcf/_2_  (.A(net265),
    .B_N(\sbox_aesinv_inst.m3f0fffcf/_0_ ),
    .Y(\sbox_aesinv_inst.x3f0fffcf ));
 sg13g2_or2_1 \sbox_aesinv_inst.m3f557fff/_1_  (.X(\sbox_aesinv_inst.m3f557fff/_0_ ),
    .B(net291),
    .A(\sbox_aesinv_inst.xc000c000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m3f557fff/_2_  (.B1(\sbox_aesinv_inst.m3f557fff/_0_ ),
    .Y(\sbox_aesinv_inst.x3f557fff ),
    .A1(\sbox_aesinv_inst.xffaa0000 ),
    .A2(net269));
 sg13g2_nand3_1 \sbox_aesinv_inst.m3fff2faf/_1_  (.B(\sbox_aesinv_inst.xfffff0f0 ),
    .C(net276),
    .A(net331),
    .Y(\sbox_aesinv_inst.m3fff2faf/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m3fff2faf/_2_  (.A(\sbox_aesinv_inst.xc000c000 ),
    .B_N(\sbox_aesinv_inst.m3fff2faf/_0_ ),
    .Y(\sbox_aesinv_inst.x3fff2faf ));
 sg13g2_nand2_1 \sbox_aesinv_inst.m3fffffff/_0_  (.Y(\sbox_aesinv_inst.x3fffffff ),
    .A(net263),
    .B(net265));
 sg13g2_nand4_1 \sbox_aesinv_inst.m4/_0_  (.B(\sbox_aesinv_inst.x4a ),
    .C(\sbox_aesinv_inst.x4c ),
    .A(\sbox_aesinv_inst.x4b ),
    .Y(\sbox_aesinv_inst.x4 ),
    .D(\sbox_aesinv_inst.x4d ));
 sg13g2_inv_1 \sbox_aesinv_inst.m40/_1_  (.Y(\sbox_aesinv_inst.m40/_0_ ),
    .A(net1));
 sg13g2_nor3_2 \sbox_aesinv_inst.m40/_2_  (.A(\sbox_aesinv_inst.m40/_0_ ),
    .B(net2),
    .C(net3),
    .Y(\sbox_aesinv_inst.x40 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m40484048/_0_  (.A(\sbox_aesinv_inst.xaaa0aaa0 ),
    .B_N(\sbox_aesinv_inst.xc8c8c8c8 ),
    .Y(\sbox_aesinv_inst.x40484048 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m40c00000/_0_  (.A(net270),
    .B_N(net265),
    .Y(\sbox_aesinv_inst.x40c00000 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m41d5cc5c/_0_  (.A1(\sbox_aesinv_inst.xbb3333ff ),
    .A2(\sbox_aesinv_inst.xf0a0f3a3 ),
    .Y(\sbox_aesinv_inst.x41d5cc5c ),
    .B1(\sbox_aesinv_inst.x0e0a0000 ));
 sg13g2_nand2_1 \sbox_aesinv_inst.m4213e265/_1_  (.Y(\sbox_aesinv_inst.m4213e265/_0_ ),
    .A(\sbox_aesinv_inst.x4e5feeff ),
    .B(\sbox_aesinv_inst.xf333f377 ));
 sg13g2_nor2_1 \sbox_aesinv_inst.m4213e265/_2_  (.A(\sbox_aesinv_inst.x0000101a ),
    .B(\sbox_aesinv_inst.m4213e265/_0_ ),
    .Y(\sbox_aesinv_inst.x4213e265 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m42e28881/_0_  (.A1(\sbox_aesinv_inst.xfffffffe ),
    .A2(\sbox_aesinv_inst.x151d777f ),
    .Y(\sbox_aesinv_inst.x42e28881 ),
    .B1(\sbox_aesinv_inst.xa8000000 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m4332245f/_1_  (.B(\sbox_aesinv_inst.xfcecf8a0 ),
    .C(\sbox_aesinv_inst.xbfffffff ),
    .A(\sbox_aesinv_inst.xffddddff ),
    .Y(\sbox_aesinv_inst.m4332245f/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m4332245f/_2_  (.A(\sbox_aesinv_inst.x00050300 ),
    .B_N(\sbox_aesinv_inst.m4332245f/_0_ ),
    .Y(\sbox_aesinv_inst.x4332245f ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m434a8cf5/_1_  (.B(\sbox_aesinv_inst.xcccf030f ),
    .C(\sbox_aesinv_inst.xafa5ffff ),
    .A(\sbox_aesinv_inst.xffffffaa ),
    .Y(\sbox_aesinv_inst.m434a8cf5/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m434a8cf5/_2_  (.A(\sbox_aesinv_inst.x30307000 ),
    .B_N(\sbox_aesinv_inst.m434a8cf5/_0_ ),
    .Y(\sbox_aesinv_inst.x434a8cf5 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m43fecdd2/_1_  (.B(\sbox_aesinv_inst.xfeecfaa8 ),
    .C(\sbox_aesinv_inst.xfd11ffff ),
    .A(\sbox_aesinv_inst.xbfbf373f ),
    .Y(\sbox_aesinv_inst.m43fecdd2/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m43fecdd2/_2_  (.A(\sbox_aesinv_inst.x00010005 ),
    .B_N(\sbox_aesinv_inst.m43fecdd2/_0_ ),
    .Y(\sbox_aesinv_inst.x43fecdd2 ));
 sg13g2_and2_1 \sbox_aesinv_inst.m4638af86/_1_  (.A(\sbox_aesinv_inst.x33cfffff ),
    .B(\sbox_aesinv_inst.x55775071 ),
    .X(\sbox_aesinv_inst.m4638af86/_0_ ));
 sg13g2_nor3_1 \sbox_aesinv_inst.m4638af86/_2_  (.A(\sbox_aesinv_inst.xa8800000 ),
    .B(\sbox_aesinv_inst.x00000008 ),
    .C(\sbox_aesinv_inst.m4638af86/_0_ ),
    .Y(\sbox_aesinv_inst.x4638af86 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m4a/_0_  (.Y(\sbox_aesinv_inst.x4a ),
    .B1(\sbox_aesinv_inst.xf12405c2 ),
    .B2(\sbox_aesinv_inst.x40 ),
    .A2(\sbox_aesinv_inst.x80 ),
    .A1(\sbox_aesinv_inst.x9d97aa84 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m4b/_0_  (.Y(\sbox_aesinv_inst.x4b ),
    .B1(\sbox_aesinv_inst.xc6aca424 ),
    .B2(\sbox_aesinv_inst.x10 ),
    .A2(\sbox_aesinv_inst.x20 ),
    .A1(\sbox_aesinv_inst.xe3ab5bd2 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m4c/_0_  (.Y(\sbox_aesinv_inst.x4c ),
    .B1(\sbox_aesinv_inst.x7847e6db ),
    .B2(\sbox_aesinv_inst.x04 ),
    .A2(\sbox_aesinv_inst.x08 ),
    .A1(\sbox_aesinv_inst.xe2cda26e ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m4d/_0_  (.Y(\sbox_aesinv_inst.x4d ),
    .B1(\sbox_aesinv_inst.x23369e29 ),
    .B2(\sbox_aesinv_inst.x01 ),
    .A2(\sbox_aesinv_inst.x02 ),
    .A1(\sbox_aesinv_inst.xd1f16c3a ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m4e5feeff/_1_  (.B(net333),
    .C(net320),
    .A(\sbox_aesinv_inst.xff00ff00 ),
    .Y(\sbox_aesinv_inst.m4e5feeff/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m4e5feeff/_2_  (.A(net268),
    .B_N(\sbox_aesinv_inst.m4e5feeff/_0_ ),
    .Y(\sbox_aesinv_inst.x4e5feeff ));
 sg13g2_nand4_1 \sbox_aesinv_inst.m5/_0_  (.B(\sbox_aesinv_inst.x5a ),
    .C(\sbox_aesinv_inst.x5c ),
    .A(\sbox_aesinv_inst.x5b ),
    .Y(\sbox_aesinv_inst.x5 ),
    .D(\sbox_aesinv_inst.x5d ));
 sg13g2_and3_1 \sbox_aesinv_inst.m50004000/_0_  (.X(\sbox_aesinv_inst.x50004000 ),
    .A(net258),
    .B(\sbox_aesinv_inst.xf0f0f000 ),
    .C(net338));
 sg13g2_nor3_1 \sbox_aesinv_inst.m52af6f23/_0_  (.A(\sbox_aesinv_inst.x05500000 ),
    .B(\sbox_aesinv_inst.xa8008000 ),
    .C(\sbox_aesinv_inst.x000010dc ),
    .Y(\sbox_aesinv_inst.x52af6f23 ));
 sg13g2_and2_1 \sbox_aesinv_inst.m52c516d9/_1_  (.A(\sbox_aesinv_inst.x131317df ),
    .B(\sbox_aesinv_inst.xfeccfec8 ),
    .X(\sbox_aesinv_inst.m52c516d9/_0_ ));
 sg13g2_or3_1 \sbox_aesinv_inst.m52c516d9/_2_  (.A(\sbox_aesinv_inst.x40c00000 ),
    .B(\sbox_aesinv_inst.x00050011 ),
    .C(\sbox_aesinv_inst.m52c516d9/_0_ ),
    .X(\sbox_aesinv_inst.x52c516d9 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m54eaa319/_1_  (.B(\sbox_aesinv_inst.xddf7ddf7 ),
    .C(\sbox_aesinv_inst.x01155fff ),
    .A(\sbox_aesinv_inst.xfffffeee ),
    .Y(\sbox_aesinv_inst.m54eaa319/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m54eaa319/_2_  (.A(net267),
    .B_N(\sbox_aesinv_inst.m54eaa319/_0_ ),
    .Y(\sbox_aesinv_inst.x54eaa319 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m55556666/_0_  (.A(\sbox_aesinv_inst.xaaaa8888 ),
    .B_N(\sbox_aesinv_inst.xffffeeee ),
    .Y(\sbox_aesinv_inst.x55556666 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m55775071/_1_  (.B(net311),
    .C(net282),
    .A(\sbox_aesinv_inst.xffeeffee ),
    .Y(\sbox_aesinv_inst.m55775071/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m55775071/_2_  (.A(\sbox_aesinv_inst.xaa88aa88 ),
    .B_N(\sbox_aesinv_inst.m55775071/_0_ ),
    .Y(\sbox_aesinv_inst.x55775071 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m557f00ff/_1_  (.X(\sbox_aesinv_inst.m557f00ff/_0_ ),
    .B(net283),
    .A(\sbox_aesinv_inst.xaaaa0000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m557f00ff/_2_  (.B1(\sbox_aesinv_inst.m557f00ff/_0_ ),
    .Y(\sbox_aesinv_inst.x557f00ff ),
    .A1(\sbox_aesinv_inst.xff00ff00 ),
    .A2(net266));
 sg13g2_or2_1 \sbox_aesinv_inst.m571fff3f/_1_  (.X(\sbox_aesinv_inst.m571fff3f/_0_ ),
    .B(net297),
    .A(\sbox_aesinv_inst.xaaaa0000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m571fff3f/_2_  (.B1(\sbox_aesinv_inst.m571fff3f/_0_ ),
    .Y(\sbox_aesinv_inst.x571fff3f ),
    .A1(\sbox_aesinv_inst.xccc0ccc0 ),
    .A2(\sbox_aesinv_inst.xa0a00000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m57ffff00/_1_  (.X(\sbox_aesinv_inst.m57ffff00/_0_ ),
    .B(net282),
    .A(\sbox_aesinv_inst.xaa000000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m57ffff00/_2_  (.B1(\sbox_aesinv_inst.m57ffff00/_0_ ),
    .Y(\sbox_aesinv_inst.x57ffff00 ),
    .A1(net259),
    .A2(net296));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m5a/_0_  (.Y(\sbox_aesinv_inst.x5a ),
    .B1(\sbox_aesinv_inst.x5b847ba9 ),
    .B2(\sbox_aesinv_inst.x40 ),
    .A2(\sbox_aesinv_inst.x80 ),
    .A1(\sbox_aesinv_inst.x2fa5e682 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m5a5f5b5f/_1_  (.B(net258),
    .C(net303),
    .A(net330),
    .Y(\sbox_aesinv_inst.m5a5f5b5f/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m5a5f5b5f/_2_  (.A(\sbox_aesinv_inst.xa0a0a0a0 ),
    .B_N(\sbox_aesinv_inst.m5a5f5b5f/_0_ ),
    .Y(\sbox_aesinv_inst.x5a5f5b5f ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m5aaa5aaa/_0_  (.A(net270),
    .B_N(\sbox_aesinv_inst.xfaaafaaa ),
    .Y(\sbox_aesinv_inst.x5aaa5aaa ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m5b/_0_  (.Y(\sbox_aesinv_inst.x5b ),
    .B1(\sbox_aesinv_inst.x24cc4461 ),
    .B2(\sbox_aesinv_inst.x10 ),
    .A2(\sbox_aesinv_inst.x20 ),
    .A1(\sbox_aesinv_inst.xf446ce08 ));
 sg13g2_and2_1 \sbox_aesinv_inst.m5b847ba9/_1_  (.A(\sbox_aesinv_inst.xfefafefa ),
    .B(\sbox_aesinv_inst.x055f0557 ),
    .X(\sbox_aesinv_inst.m5b847ba9/_0_ ));
 sg13g2_nor3_1 \sbox_aesinv_inst.m5b847ba9/_2_  (.A(\sbox_aesinv_inst.xa0008000 ),
    .B(\sbox_aesinv_inst.x00330404 ),
    .C(\sbox_aesinv_inst.m5b847ba9/_0_ ),
    .Y(\sbox_aesinv_inst.x5b847ba9 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m5c/_0_  (.Y(\sbox_aesinv_inst.x5c ),
    .B1(\sbox_aesinv_inst.x54eaa319 ),
    .B2(\sbox_aesinv_inst.x04 ),
    .A2(\sbox_aesinv_inst.x08 ),
    .A1(\sbox_aesinv_inst.x854f7ef5 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m5d/_0_  (.Y(\sbox_aesinv_inst.x5d ),
    .B1(\sbox_aesinv_inst.xef715dd5 ),
    .B2(\sbox_aesinv_inst.x01 ),
    .A2(\sbox_aesinv_inst.x02 ),
    .A1(\sbox_aesinv_inst.x318ab4e1 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m5e9f51e4/_1_  (.B(\sbox_aesinv_inst.xffeeee88 ),
    .C(\sbox_aesinv_inst.xf1f1ffff ),
    .A(\sbox_aesinv_inst.xaf7faf7f ),
    .Y(\sbox_aesinv_inst.m5e9f51e4/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m5e9f51e4/_2_  (.A(\sbox_aesinv_inst.x00000013 ),
    .B_N(\sbox_aesinv_inst.m5e9f51e4/_0_ ),
    .Y(\sbox_aesinv_inst.x5e9f51e4 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m5f5ffafa/_0_  (.A(net268),
    .B_N(\sbox_aesinv_inst.xfffffafa ),
    .Y(\sbox_aesinv_inst.x5f5ffafa ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m5fff0faf/_1_  (.B(\sbox_aesinv_inst.xfffff0f0 ),
    .C(net275),
    .A(net331),
    .Y(\sbox_aesinv_inst.m5fff0faf/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m5fff0faf/_2_  (.A(net269),
    .B_N(\sbox_aesinv_inst.m5fff0faf/_0_ ),
    .Y(\sbox_aesinv_inst.x5fff0faf ));
 sg13g2_nand4_1 \sbox_aesinv_inst.m6/_0_  (.B(\sbox_aesinv_inst.x6a ),
    .C(\sbox_aesinv_inst.x6c ),
    .A(\sbox_aesinv_inst.x6b ),
    .Y(\sbox_aesinv_inst.x6 ),
    .D(\sbox_aesinv_inst.x6d ));
 sg13g2_and2_1 \sbox_aesinv_inst.m6191ae47/_1_  (.A(\sbox_aesinv_inst.x1f7f55ff ),
    .B(\sbox_aesinv_inst.xfeeef8a8 ),
    .X(\sbox_aesinv_inst.m6191ae47/_0_ ));
 sg13g2_nor3_1 \sbox_aesinv_inst.m6191ae47/_2_  (.A(\sbox_aesinv_inst.x88000000 ),
    .B(\sbox_aesinv_inst.x00001110 ),
    .C(\sbox_aesinv_inst.m6191ae47/_0_ ),
    .Y(\sbox_aesinv_inst.x6191ae47 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m6a/_0_  (.Y(\sbox_aesinv_inst.x6a ),
    .B1(\sbox_aesinv_inst.xc4cf14da ),
    .B2(\sbox_aesinv_inst.x40 ),
    .A2(\sbox_aesinv_inst.x80 ),
    .A1(\sbox_aesinv_inst.xb047c23f ));
 sg13g2_a221oi_1 \sbox_aesinv_inst.m6a86145f/_0_  (.B2(\sbox_aesinv_inst.xfff8ffa0 ),
    .C1(\sbox_aesinv_inst.x80000000 ),
    .B1(\sbox_aesinv_inst.x007fabff ),
    .A1(\sbox_aesinv_inst.x15555050 ),
    .Y(\sbox_aesinv_inst.x6a86145f ),
    .A2(\sbox_aesinv_inst.xdd11cc00 ));
 sg13g2_or3_1 \sbox_aesinv_inst.m6ad30f0f/_0_  (.A(\sbox_aesinv_inst.x40c00000 ),
    .B(\sbox_aesinv_inst.x2a000000 ),
    .C(\sbox_aesinv_inst.x00130f0f ),
    .X(\sbox_aesinv_inst.x6ad30f0f ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m6b/_0_  (.Y(\sbox_aesinv_inst.x6b ),
    .B1(\sbox_aesinv_inst.x42e28881 ),
    .B2(\sbox_aesinv_inst.x10 ),
    .A2(\sbox_aesinv_inst.x20 ),
    .A1(\sbox_aesinv_inst.xf4bcfdb0 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m6c/_0_  (.Y(\sbox_aesinv_inst.x6c ),
    .B1(\sbox_aesinv_inst.xd2a0de7f ),
    .B2(\sbox_aesinv_inst.x04 ),
    .A2(\sbox_aesinv_inst.x08 ),
    .A1(\sbox_aesinv_inst.x1f7b28d7 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m6d/_0_  (.Y(\sbox_aesinv_inst.x6d ),
    .B1(\sbox_aesinv_inst.x52c516d9 ),
    .B2(\sbox_aesinv_inst.x01 ),
    .A2(\sbox_aesinv_inst.x02 ),
    .A1(\sbox_aesinv_inst.x4213e265 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m6d287e63/_1_  (.B(\sbox_aesinv_inst.x3777053f ),
    .C(\sbox_aesinv_inst.xfffffffc ),
    .A(\sbox_aesinv_inst.x5a5f5b5f ),
    .Y(\sbox_aesinv_inst.m6d287e63/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m6d287e63/_2_  (.A(net274),
    .B_N(\sbox_aesinv_inst.m6d287e63/_0_ ),
    .Y(\sbox_aesinv_inst.x6d287e63 ));
 sg13g2_nand4_1 \sbox_aesinv_inst.m7/_0_  (.B(\sbox_aesinv_inst.x7a ),
    .C(\sbox_aesinv_inst.x7c ),
    .A(\sbox_aesinv_inst.x7b ),
    .Y(\sbox_aesinv_inst.x7 ),
    .D(\sbox_aesinv_inst.x7d ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m7077f7ff/_1_  (.B(\sbox_aesinv_inst.xff00cc00 ),
    .C(net315),
    .A(\sbox_aesinv_inst.xff00aa00 ),
    .Y(\sbox_aesinv_inst.m7077f7ff/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m7077f7ff/_2_  (.A(net271),
    .B_N(\sbox_aesinv_inst.m7077f7ff/_0_ ),
    .Y(\sbox_aesinv_inst.x7077f7ff ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m777717ff/_1_  (.B(\sbox_aesinv_inst.xfc00fc00 ),
    .C(net281),
    .A(\sbox_aesinv_inst.xeaeaeaea ),
    .Y(\sbox_aesinv_inst.m777717ff/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m777717ff/_2_  (.A(net271),
    .B_N(\sbox_aesinv_inst.m777717ff/_0_ ),
    .Y(\sbox_aesinv_inst.x777717ff ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m77cd77ff/_1_  (.B(\sbox_aesinv_inst.xfafa0000 ),
    .C(net319),
    .A(net292),
    .Y(\sbox_aesinv_inst.m77cd77ff/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m77cd77ff/_2_  (.A(net272),
    .B_N(\sbox_aesinv_inst.m77cd77ff/_0_ ),
    .Y(\sbox_aesinv_inst.x77cd77ff ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m77fc77fc/_0_  (.A(net273),
    .B_N(\sbox_aesinv_inst.xfffcfffc ),
    .Y(\sbox_aesinv_inst.x77fc77fc ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m77ff3337/_1_  (.B(\sbox_aesinv_inst.xfcfccccc ),
    .C(net283),
    .A(\sbox_aesinv_inst.xfffafffa ),
    .Y(\sbox_aesinv_inst.m77ff3337/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m77ff3337/_2_  (.A(net273),
    .B_N(\sbox_aesinv_inst.m77ff3337/_0_ ),
    .Y(\sbox_aesinv_inst.x77ff3337 ));
 sg13g2_and2_1 \sbox_aesinv_inst.m7847e6db/_1_  (.A(\sbox_aesinv_inst.x7077f7ff ),
    .B(\sbox_aesinv_inst.xffcceec8 ),
    .X(\sbox_aesinv_inst.m7847e6db/_0_ ));
 sg13g2_or3_1 \sbox_aesinv_inst.m7847e6db/_2_  (.A(\sbox_aesinv_inst.x08000000 ),
    .B(\sbox_aesinv_inst.x00070013 ),
    .C(\sbox_aesinv_inst.m7847e6db/_0_ ),
    .X(\sbox_aesinv_inst.x7847e6db ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m7a/_0_  (.Y(\sbox_aesinv_inst.x7a ),
    .B1(\sbox_aesinv_inst.x2ca62526 ),
    .B2(\sbox_aesinv_inst.x40 ),
    .A2(\sbox_aesinv_inst.x80 ),
    .A1(\sbox_aesinv_inst.x12bf5b4f ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m7b/_0_  (.Y(\sbox_aesinv_inst.x7b ),
    .B1(\sbox_aesinv_inst.xeecc98e2 ),
    .B2(\sbox_aesinv_inst.x10 ),
    .A2(\sbox_aesinv_inst.x20 ),
    .A1(\sbox_aesinv_inst.x6ad30f0f ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m7c/_0_  (.Y(\sbox_aesinv_inst.x7c ),
    .B1(\sbox_aesinv_inst.x434a8cf5 ),
    .B2(\sbox_aesinv_inst.x04 ),
    .A2(\sbox_aesinv_inst.x08 ),
    .A1(\sbox_aesinv_inst.x43fecdd2 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m7c7c7c7d/_1_  (.B(net304),
    .C(\sbox_aesinv_inst.xffffffaa ),
    .A(net318),
    .Y(\sbox_aesinv_inst.m7c7c7c7d/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m7c7c7c7d/_2_  (.A(net274),
    .B_N(\sbox_aesinv_inst.m7c7c7c7d/_0_ ),
    .Y(\sbox_aesinv_inst.x7c7c7c7d ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m7ca10f66/_1_  (.B(\sbox_aesinv_inst.xfffef888 ),
    .C(\sbox_aesinv_inst.xf35ff3ff ),
    .A(\sbox_aesinv_inst.x8fdfffff ),
    .Y(\sbox_aesinv_inst.m7ca10f66/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m7ca10f66/_2_  (.A(\sbox_aesinv_inst.x00001011 ),
    .B_N(\sbox_aesinv_inst.m7ca10f66/_0_ ),
    .Y(\sbox_aesinv_inst.x7ca10f66 ));
 sg13g2_a22oi_1 \sbox_aesinv_inst.m7d/_0_  (.Y(\sbox_aesinv_inst.x7d ),
    .B1(\sbox_aesinv_inst.xcbea0a80 ),
    .B2(\sbox_aesinv_inst.x01 ),
    .A2(\sbox_aesinv_inst.x02 ),
    .A1(\sbox_aesinv_inst.x6a86145f ));
 sg13g2_or2_1 \sbox_aesinv_inst.m7f5f3300/_1_  (.X(\sbox_aesinv_inst.m7f5f3300/_0_ ),
    .B(net285),
    .A(net268));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m7f5f3300/_2_  (.B1(\sbox_aesinv_inst.m7f5f3300/_0_ ),
    .Y(\sbox_aesinv_inst.x7f5f3300 ),
    .A1(\sbox_aesinv_inst.xcc00cc00 ),
    .A2(net298));
 sg13g2_nor3_2 \sbox_aesinv_inst.m80/_0_  (.A(net2),
    .B(net1),
    .C(net3),
    .Y(\sbox_aesinv_inst.x80 ));
 sg13g2_and2_1 \sbox_aesinv_inst.m80000000/_0_  (.A(net269),
    .B(net266),
    .X(\sbox_aesinv_inst.x80000000 ));
 sg13g2_nor3_2 \sbox_aesinv_inst.m80808080/_0_  (.A(net303),
    .B(net330),
    .C(net318),
    .Y(\sbox_aesinv_inst.x80808080 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m854f7ef5/_1_  (.X(\sbox_aesinv_inst.m854f7ef5/_0_ ),
    .B(\sbox_aesinv_inst.x3030f1f0 ),
    .A(\sbox_aesinv_inst.x5aaa5aaa ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m854f7ef5/_2_  (.B(\sbox_aesinv_inst.xffff8f0f ),
    .C(\sbox_aesinv_inst.m854f7ef5/_0_ ),
    .A(\sbox_aesinv_inst.xfff5f5ff ),
    .Y(\sbox_aesinv_inst.x854f7ef5 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m88000000/_0_  (.A(net301),
    .B_N(net271),
    .Y(\sbox_aesinv_inst.x88000000 ));
 sg13g2_nor3_2 \sbox_aesinv_inst.m88008800/_0_  (.A(net330),
    .B(net291),
    .C(net318),
    .Y(\sbox_aesinv_inst.x88008800 ));
 sg13g2_nor3_1 \sbox_aesinv_inst.m88880000/_0_  (.A(net328),
    .B(net342),
    .C(net288),
    .Y(\sbox_aesinv_inst.x88880000 ));
 sg13g2_nor2_1 \sbox_aesinv_inst.m88888888/_0_  (.A(net325),
    .B(net338),
    .Y(\sbox_aesinv_inst.x88888888 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m8ad2e815/_1_  (.B(\sbox_aesinv_inst.xffffffea ),
    .C(\sbox_aesinv_inst.x777717ff ),
    .A(\sbox_aesinv_inst.xf5a5ffff ),
    .Y(\sbox_aesinv_inst.m8ad2e815/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m8ad2e815/_2_  (.A(\sbox_aesinv_inst.x040c0000 ),
    .B_N(\sbox_aesinv_inst.m8ad2e815/_0_ ),
    .Y(\sbox_aesinv_inst.x8ad2e815 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.m8b30445b/_1_  (.B(\sbox_aesinv_inst.x77ff3337 ),
    .C(\sbox_aesinv_inst.xfccfffff ),
    .A(\sbox_aesinv_inst.xffffffec ),
    .Y(\sbox_aesinv_inst.m8b30445b/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.m8b30445b/_2_  (.A(\sbox_aesinv_inst.x00008880 ),
    .B_N(\sbox_aesinv_inst.m8b30445b/_0_ ),
    .Y(\sbox_aesinv_inst.x8b30445b ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m8df398a3/_0_  (.A1(\sbox_aesinv_inst.x77fc77fc ),
    .A2(\sbox_aesinv_inst.xaa0faf5f ),
    .Y(\sbox_aesinv_inst.x8df398a3 ),
    .B1(\sbox_aesinv_inst.x50004000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.m8fdfffff/_1_  (.X(\sbox_aesinv_inst.m8fdfffff/_0_ ),
    .B(net327),
    .A(net340));
 sg13g2_o21ai_1 \sbox_aesinv_inst.m8fdfffff/_2_  (.B1(\sbox_aesinv_inst.m8fdfffff/_0_ ),
    .Y(\sbox_aesinv_inst.x8fdfffff ),
    .A1(\sbox_aesinv_inst.xf0000000 ),
    .A2(net268));
 sg13g2_and2_1 \sbox_aesinv_inst.m96492239/_1_  (.A(\sbox_aesinv_inst.x175f333f ),
    .B(\sbox_aesinv_inst.xfec8eec8 ),
    .X(\sbox_aesinv_inst.m96492239/_0_ ));
 sg13g2_or3_1 \sbox_aesinv_inst.m96492239/_2_  (.A(\sbox_aesinv_inst.x80000000 ),
    .B(\sbox_aesinv_inst.x00010031 ),
    .C(\sbox_aesinv_inst.m96492239/_0_ ),
    .X(\sbox_aesinv_inst.x96492239 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.m9d97aa84/_0_  (.A1(\sbox_aesinv_inst.x37303733 ),
    .A2(\sbox_aesinv_inst.xaaaf153f ),
    .Y(\sbox_aesinv_inst.x9d97aa84 ),
    .B1(\sbox_aesinv_inst.x40484048 ));
 sg13g2_and2_1 \sbox_aesinv_inst.ma0008000/_0_  (.A(net269),
    .B(net258),
    .X(\sbox_aesinv_inst.xa0008000 ));
 sg13g2_nor3_1 \sbox_aesinv_inst.ma000a000/_0_  (.A(net338),
    .B(net297),
    .C(net309),
    .Y(\sbox_aesinv_inst.xa000a000 ));
 sg13g2_nor3_2 \sbox_aesinv_inst.ma0a00000/_0_  (.A(net310),
    .B(net339),
    .C(net284),
    .Y(\sbox_aesinv_inst.xa0a00000 ));
 sg13g2_nor2_1 \sbox_aesinv_inst.ma0a0a0a0/_0_  (.A(net303),
    .B(net330),
    .Y(\sbox_aesinv_inst.xa0a0a0a0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.ma0a0a1a1/_1_  (.X(\sbox_aesinv_inst.ma0a0a1a1/_0_ ),
    .B(net311),
    .A(net339));
 sg13g2_o21ai_1 \sbox_aesinv_inst.ma0a0a1a1/_2_  (.B1(\sbox_aesinv_inst.ma0a0a1a1/_0_ ),
    .Y(\sbox_aesinv_inst.xa0a0a1a1 ),
    .A1(\sbox_aesinv_inst.xfffffafa ),
    .A2(\sbox_aesinv_inst.xfcfccccc ));
 sg13g2_nand3_1 \sbox_aesinv_inst.ma0fb7cd2/_1_  (.B(\sbox_aesinv_inst.xff05333f ),
    .C(\sbox_aesinv_inst.xfffcfffd ),
    .A(\sbox_aesinv_inst.x5fff0faf ),
    .Y(\sbox_aesinv_inst.ma0fb7cd2/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.ma0fb7cd2/_2_  (.A(\sbox_aesinv_inst.x00008000 ),
    .B_N(\sbox_aesinv_inst.ma0fb7cd2/_0_ ),
    .Y(\sbox_aesinv_inst.xa0fb7cd2 ));
 sg13g2_or2_1 \sbox_aesinv_inst.ma1b3a5bf/_1_  (.X(\sbox_aesinv_inst.ma1b3a5bf/_0_ ),
    .B(net314),
    .A(net341));
 sg13g2_o21ai_1 \sbox_aesinv_inst.ma1b3a5bf/_2_  (.B1(\sbox_aesinv_inst.ma1b3a5bf/_0_ ),
    .Y(\sbox_aesinv_inst.xa1b3a5bf ),
    .A1(\sbox_aesinv_inst.xfa00fa00 ),
    .A2(\sbox_aesinv_inst.xccccc0c0 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.ma4b75f65/_0_  (.B1(\sbox_aesinv_inst.x5f5ffafa ),
    .Y(\sbox_aesinv_inst.xa4b75f65 ),
    .A1(\sbox_aesinv_inst.x0100011f ),
    .A2(\sbox_aesinv_inst.xfac8a080 ));
 sg13g2_and2_1 \sbox_aesinv_inst.ma8000000/_0_  (.A(net267),
    .B(net259),
    .X(\sbox_aesinv_inst.xa8000000 ));
 sg13g2_and3_1 \sbox_aesinv_inst.ma8008000/_0_  (.X(\sbox_aesinv_inst.xa8008000 ),
    .A(\sbox_aesinv_inst.xff00f000 ),
    .B(\sbox_aesinv_inst.xfc00fc00 ),
    .C(\sbox_aesinv_inst.xaaaa8888 ));
 sg13g2_and3_1 \sbox_aesinv_inst.ma8800000/_0_  (.X(\sbox_aesinv_inst.xa8800000 ),
    .A(\sbox_aesinv_inst.xffcc0000 ),
    .B(net257),
    .C(\sbox_aesinv_inst.xa8a8a8a8 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.ma8a8a8a8/_0_  (.B1(net338),
    .Y(\sbox_aesinv_inst.xa8a8a8a8 ),
    .A2(net309),
    .A1(net325));
 sg13g2_a21oi_1 \sbox_aesinv_inst.ma90301b8/_0_  (.A1(\sbox_aesinv_inst.x57ffff00 ),
    .A2(\sbox_aesinv_inst.xfaf8fa00 ),
    .Y(\sbox_aesinv_inst.xa90301b8 ),
    .B1(\sbox_aesinv_inst.x04044447 ));
 sg13g2_and2_1 \sbox_aesinv_inst.ma9e15289/_1_  (.A(\sbox_aesinv_inst.x571fff3f ),
    .B(\sbox_aesinv_inst.xfefea8a0 ),
    .X(\sbox_aesinv_inst.ma9e15289/_0_ ));
 sg13g2_nor3_1 \sbox_aesinv_inst.ma9e15289/_2_  (.A(\sbox_aesinv_inst.x00060006 ),
    .B(\sbox_aesinv_inst.x00000550 ),
    .C(\sbox_aesinv_inst.ma9e15289/_0_ ),
    .Y(\sbox_aesinv_inst.xa9e15289 ));
 sg13g2_nor3_2 \sbox_aesinv_inst.maa000000/_0_  (.A(net330),
    .B(net290),
    .C(net275),
    .Y(\sbox_aesinv_inst.xaa000000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.maa0faf5f/_1_  (.X(\sbox_aesinv_inst.maa0faf5f/_0_ ),
    .B(net300),
    .A(net340));
 sg13g2_o21ai_1 \sbox_aesinv_inst.maa0faf5f/_2_  (.B1(\sbox_aesinv_inst.maa0faf5f/_0_ ),
    .Y(\sbox_aesinv_inst.xaa0faf5f ),
    .A1(\sbox_aesinv_inst.xff00f000 ),
    .A2(\sbox_aesinv_inst.xf0f0a0a0 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.maa88aa88/_0_  (.B1(net336),
    .Y(\sbox_aesinv_inst.xaa88aa88 ),
    .A2(net295),
    .A1(net324));
 sg13g2_a21oi_2 \sbox_aesinv_inst.maaa0aaa0/_0_  (.B1(net335),
    .Y(\sbox_aesinv_inst.xaaa0aaa0 ),
    .A2(net294),
    .A1(net306));
 sg13g2_nor2_2 \sbox_aesinv_inst.maaaa0000/_0_  (.A(net284),
    .B(net338),
    .Y(\sbox_aesinv_inst.xaaaa0000 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.maaaa8888/_0_  (.B1(net340),
    .Y(\sbox_aesinv_inst.xaaaa8888 ),
    .A2(net327),
    .A1(net286));
 sg13g2_a21oi_1 \sbox_aesinv_inst.maaaaa0a0/_0_  (.A1(net285),
    .A2(net310),
    .Y(\sbox_aesinv_inst.xaaaaa0a0 ),
    .B1(net339));
 sg13g2_a21oi_2 \sbox_aesinv_inst.maaaaaa00/_0_  (.B1(net331),
    .Y(\sbox_aesinv_inst.xaaaaaa00 ),
    .A2(net290),
    .A1(net275));
 sg13g2_or2_1 \sbox_aesinv_inst.maaaf153f/_1_  (.X(\sbox_aesinv_inst.maaaf153f/_0_ ),
    .B(net281),
    .A(net336));
 sg13g2_o21ai_1 \sbox_aesinv_inst.maaaf153f/_2_  (.B1(\sbox_aesinv_inst.maaaf153f/_0_ ),
    .Y(\sbox_aesinv_inst.xaaaf153f ),
    .A1(\sbox_aesinv_inst.xff00aa00 ),
    .A2(\sbox_aesinv_inst.xf0f0c0c0 ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.madffadff/_0_  (.Y(\sbox_aesinv_inst.xadffadff ),
    .B(\sbox_aesinv_inst.xfa00fa00 ),
    .A_N(\sbox_aesinv_inst.xa8a8a8a8 ));
 sg13g2_or2_1 \sbox_aesinv_inst.maf7faf7f/_1_  (.X(\sbox_aesinv_inst.maf7faf7f/_0_ ),
    .B(net294),
    .A(net334));
 sg13g2_o21ai_1 \sbox_aesinv_inst.maf7faf7f/_2_  (.B1(\sbox_aesinv_inst.maf7faf7f/_0_ ),
    .Y(\sbox_aesinv_inst.xaf7faf7f ),
    .A1(\sbox_aesinv_inst.xf000f000 ),
    .A2(net274));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mafa5ffff/_0_  (.Y(\sbox_aesinv_inst.xafa5ffff ),
    .B(\sbox_aesinv_inst.xfafa0000 ),
    .A_N(\sbox_aesinv_inst.xaaa0aaa0 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mb047c23f/_1_  (.B1(\sbox_aesinv_inst.xbb77ffff ),
    .Y(\sbox_aesinv_inst.mb047c23f/_0_ ),
    .A1(\sbox_aesinv_inst.x000f023f ),
    .A2(\sbox_aesinv_inst.xf0c0c000 ));
 sg13g2_inv_1 \sbox_aesinv_inst.mb047c23f/_2_  (.Y(\sbox_aesinv_inst.xb047c23f ),
    .A(\sbox_aesinv_inst.mb047c23f/_0_ ));
 sg13g2_or2_1 \sbox_aesinv_inst.mb1b1f5f7/_1_  (.X(\sbox_aesinv_inst.mb1b1f5f7/_0_ ),
    .B(net305),
    .A(net337));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mb1b1f5f7/_2_  (.B1(\sbox_aesinv_inst.mb1b1f5f7/_0_ ),
    .Y(\sbox_aesinv_inst.xb1b1f5f7 ),
    .A1(\sbox_aesinv_inst.xcccc8888 ),
    .A2(\sbox_aesinv_inst.xaaaaaa00 ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mbb3333ff/_0_  (.Y(\sbox_aesinv_inst.xbb3333ff ),
    .B(net261),
    .A_N(net267));
 sg13g2_or2_1 \sbox_aesinv_inst.mbb77ffff/_1_  (.X(\sbox_aesinv_inst.mbb77ffff/_0_ ),
    .B(net295),
    .A(net336));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mbb77ffff/_2_  (.B1(\sbox_aesinv_inst.mbb77ffff/_0_ ),
    .Y(\sbox_aesinv_inst.xbb77ffff ),
    .A1(net264),
    .A2(net271));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mbbbbf5f5/_0_  (.Y(\sbox_aesinv_inst.xbbbbf5f5 ),
    .B(\sbox_aesinv_inst.xeeeeaaaa ),
    .A_N(\sbox_aesinv_inst.xaaaaa0a0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mbfbf373f/_1_  (.X(\sbox_aesinv_inst.mbfbf373f/_0_ ),
    .B(net279),
    .A(net334));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mbfbf373f/_2_  (.B1(\sbox_aesinv_inst.mbfbf373f/_0_ ),
    .Y(\sbox_aesinv_inst.xbfbf373f ),
    .A1(\sbox_aesinv_inst.xc0c0c0c0 ),
    .A2(net272));
 sg13g2_nand3_1 \sbox_aesinv_inst.mbfffffff/_0_  (.B(net265),
    .C(net334),
    .A(net264),
    .Y(\sbox_aesinv_inst.xbfffffff ));
 sg13g2_and2_1 \sbox_aesinv_inst.mc0008000/_0_  (.A(\sbox_aesinv_inst.xcccc8888 ),
    .B(\sbox_aesinv_inst.xf000f000 ),
    .X(\sbox_aesinv_inst.xc0008000 ));
 sg13g2_nor3_2 \sbox_aesinv_inst.mc000c000/_0_  (.A(net304),
    .B(net291),
    .C(net318),
    .Y(\sbox_aesinv_inst.xc000c000 ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mc011c011/_0_  (.Y(\sbox_aesinv_inst.xc011c011 ),
    .B(\sbox_aesinv_inst.xffeeffee ),
    .A_N(\sbox_aesinv_inst.xc000c000 ));
 sg13g2_nor3_2 \sbox_aesinv_inst.mc0c00000/_0_  (.A(net323),
    .B(net307),
    .C(net280),
    .Y(\sbox_aesinv_inst.xc0c00000 ));
 sg13g2_nor2_1 \sbox_aesinv_inst.mc0c0c0c0/_0_  (.A(net323),
    .B(net306),
    .Y(\sbox_aesinv_inst.xc0c0c0c0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mc3c3c3cf/_1_  (.X(\sbox_aesinv_inst.mc3c3c3cf/_0_ ),
    .B(net304),
    .A(net319));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mc3c3c3cf/_2_  (.B1(\sbox_aesinv_inst.mc3c3c3cf/_0_ ),
    .Y(\sbox_aesinv_inst.xc3c3c3cf ),
    .A1(\sbox_aesinv_inst.xf0f0f0f0 ),
    .A2(net261));
 sg13g2_a21oi_1 \sbox_aesinv_inst.mc4cf14da/_0_  (.A1(\sbox_aesinv_inst.xcbffcbff ),
    .A2(\sbox_aesinv_inst.x3f00ff05 ),
    .Y(\sbox_aesinv_inst.xc4cf14da ),
    .B1(\sbox_aesinv_inst.x32302020 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mc5cfc5df/_1_  (.X(\sbox_aesinv_inst.mc5cfc5df/_0_ ),
    .B(net313),
    .A(net327));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mc5cfc5df/_2_  (.B1(\sbox_aesinv_inst.mc5cfc5df/_0_ ),
    .Y(\sbox_aesinv_inst.xc5cfc5df ),
    .A1(\sbox_aesinv_inst.xfa00fa00 ),
    .A2(\sbox_aesinv_inst.xf0f0a0a0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mc60b25d3/_1_  (.X(\sbox_aesinv_inst.mc60b25d3/_0_ ),
    .B(\sbox_aesinv_inst.xf8f0c800 ),
    .A(\sbox_aesinv_inst.x0137133f ));
 sg13g2_nand3_1 \sbox_aesinv_inst.mc60b25d3/_2_  (.B(\sbox_aesinv_inst.x3fffffff ),
    .C(\sbox_aesinv_inst.mc60b25d3/_0_ ),
    .A(\sbox_aesinv_inst.xfffcfeec ),
    .Y(\sbox_aesinv_inst.xc60b25d3 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.mc6aca424/_0_  (.A1(\sbox_aesinv_inst.x3f557fff ),
    .A2(\sbox_aesinv_inst.xf8f8c8c8 ),
    .Y(\sbox_aesinv_inst.xc6aca424 ),
    .B1(\sbox_aesinv_inst.x11131313 ));
 sg13g2_and2_1 \sbox_aesinv_inst.mc800c000/_0_  (.A(\sbox_aesinv_inst.xc8c8c8c8 ),
    .B(\sbox_aesinv_inst.xff00f000 ),
    .X(\sbox_aesinv_inst.xc800c000 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mc8c8c8c8/_0_  (.B1(net322),
    .Y(\sbox_aesinv_inst.xc8c8c8c8 ),
    .A2(net334),
    .A1(net306));
 sg13g2_nand2_1 \sbox_aesinv_inst.mcbea0a80/_0_  (.Y(\sbox_aesinv_inst.xcbea0a80 ),
    .A(\sbox_aesinv_inst.x3c3ffdff ),
    .B(\sbox_aesinv_inst.xf555f57f ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mcbffcbff/_0_  (.Y(\sbox_aesinv_inst.xcbffcbff ),
    .B(\sbox_aesinv_inst.xfc00fc00 ),
    .A_N(\sbox_aesinv_inst.xc8c8c8c8 ));
 sg13g2_nor3_1 \sbox_aesinv_inst.mcc000000/_0_  (.A(net318),
    .B(net290),
    .C(net276),
    .Y(\sbox_aesinv_inst.xcc000000 ));
 sg13g2_nor2_1 \sbox_aesinv_inst.mcc00cc00/_0_  (.A(net325),
    .B(net298),
    .Y(\sbox_aesinv_inst.xcc00cc00 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.mcc880000/_0_  (.A(net322),
    .B_N(\sbox_aesinv_inst.xffaa0000 ),
    .Y(\sbox_aesinv_inst.xcc880000 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mcc88cc88/_0_  (.B1(net325),
    .Y(\sbox_aesinv_inst.xcc88cc88 ),
    .A2(net297),
    .A1(net339));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mccc0ccc0/_0_  (.B1(net329),
    .Y(\sbox_aesinv_inst.xccc0ccc0 ),
    .A2(net298),
    .A1(net310));
 sg13g2_nor2_1 \sbox_aesinv_inst.mcccc0000/_0_  (.A(net280),
    .B(net322),
    .Y(\sbox_aesinv_inst.xcccc0000 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mcccc8888/_0_  (.B1(net322),
    .Y(\sbox_aesinv_inst.xcccc8888 ),
    .A2(net334),
    .A1(net276));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mccccc0c0/_0_  (.B1(net329),
    .Y(\sbox_aesinv_inst.xccccc0c0 ),
    .A2(net314),
    .A1(net286));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mcccccc00/_0_  (.B1(net323),
    .Y(\sbox_aesinv_inst.xcccccc00 ),
    .A2(net294),
    .A1(net279));
 sg13g2_or2_1 \sbox_aesinv_inst.mcccf030f/_1_  (.X(\sbox_aesinv_inst.mcccf030f/_0_ ),
    .B(net280),
    .A(net322));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mcccf030f/_2_  (.B1(\sbox_aesinv_inst.mcccf030f/_0_ ),
    .Y(\sbox_aesinv_inst.xcccf030f ),
    .A1(\sbox_aesinv_inst.xfff0f0f0 ),
    .A2(net262));
 sg13g2_o21ai_1 \sbox_aesinv_inst.md1f16c3a/_0_  (.B1(\sbox_aesinv_inst.x3f0fffcf ),
    .Y(\sbox_aesinv_inst.xd1f16c3a ),
    .A1(\sbox_aesinv_inst.x00001355 ),
    .A2(\sbox_aesinv_inst.xeeee8080 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.md2a0de7f/_0_  (.A1(\sbox_aesinv_inst.x7f5f3300 ),
    .A2(\sbox_aesinv_inst.xadffadff ),
    .Y(\sbox_aesinv_inst.xd2a0de7f ),
    .B1(\sbox_aesinv_inst.x00000080 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.md7997ddd/_0_  (.B1(\sbox_aesinv_inst.x2aeeaaee ),
    .Y(\sbox_aesinv_inst.xd7997ddd ),
    .A1(\sbox_aesinv_inst.x11771333 ),
    .A2(\sbox_aesinv_inst.xf8008000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mdd11cc00/_1_  (.X(\sbox_aesinv_inst.mdd11cc00/_0_ ),
    .B(net288),
    .A(\sbox_aesinv_inst.xeeee0000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mdd11cc00/_2_  (.B1(\sbox_aesinv_inst.mdd11cc00/_0_ ),
    .Y(\sbox_aesinv_inst.xdd11cc00 ),
    .A1(net328),
    .A2(net300));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mdd5555ff/_0_  (.Y(\sbox_aesinv_inst.xdd5555ff ),
    .B(\sbox_aesinv_inst.xaaaaaa00 ),
    .A_N(net263));
 sg13g2_or2_1 \sbox_aesinv_inst.mdd7fff7f/_1_  (.X(\sbox_aesinv_inst.mdd7fff7f/_0_ ),
    .B(net293),
    .A(net320));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mdd7fff7f/_2_  (.B1(\sbox_aesinv_inst.mdd7fff7f/_0_ ),
    .Y(\sbox_aesinv_inst.xdd7fff7f ),
    .A1(\sbox_aesinv_inst.xaa000000 ),
    .A2(\sbox_aesinv_inst.x80808080 ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mddf7ddf7/_0_  (.Y(\sbox_aesinv_inst.xddf7ddf7 ),
    .B(\sbox_aesinv_inst.xaa88aa88 ),
    .A_N(\sbox_aesinv_inst.xccc0ccc0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mdf77df77/_1_  (.X(\sbox_aesinv_inst.mdf77df77/_0_ ),
    .B(net297),
    .A(net325));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mdf77df77/_2_  (.B1(\sbox_aesinv_inst.mdf77df77/_0_ ),
    .Y(\sbox_aesinv_inst.xdf77df77 ),
    .A1(\sbox_aesinv_inst.xcc88cc88 ),
    .A2(net269));
 sg13g2_a21oi_1 \sbox_aesinv_inst.mdfc11244/_0_  (.A1(\sbox_aesinv_inst.x323233fb ),
    .A2(\sbox_aesinv_inst.xa1b3a5bf ),
    .Y(\sbox_aesinv_inst.xdfc11244 ),
    .B1(\sbox_aesinv_inst.x000ccc00 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mdfdf77ff/_1_  (.X(\sbox_aesinv_inst.mdfdf77ff/_0_ ),
    .B(net287),
    .A(net327));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mdfdf77ff/_2_  (.B1(\sbox_aesinv_inst.mdfdf77ff/_0_ ),
    .Y(\sbox_aesinv_inst.xdfdf77ff ),
    .A1(net268),
    .A2(net273));
 sg13g2_and3_1 \sbox_aesinv_inst.me080c000/_0_  (.X(\sbox_aesinv_inst.xe080c000 ),
    .A(\sbox_aesinv_inst.xffcccccc ),
    .B(\sbox_aesinv_inst.xf0f0f000 ),
    .C(\sbox_aesinv_inst.xeeaaeeaa ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.me0e0e0e0/_0_  (.B1(net306),
    .Y(\sbox_aesinv_inst.xe0e0e0e0 ),
    .A2(net335),
    .A1(net323));
 sg13g2_nand3b_1 \sbox_aesinv_inst.me2cda26e/_0_  (.B(\sbox_aesinv_inst.xffb3ffb3 ),
    .C(\sbox_aesinv_inst.x1d7f5dff ),
    .Y(\sbox_aesinv_inst.xe2cda26e ),
    .A_N(\sbox_aesinv_inst.x00050022 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.me3ab5bd2/_1_  (.B(\sbox_aesinv_inst.x7c7c7c7d ),
    .C(\sbox_aesinv_inst.x3fff2faf ),
    .A(\sbox_aesinv_inst.xdd5555ff ),
    .Y(\sbox_aesinv_inst.me3ab5bd2/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.me3ab5bd2/_2_  (.A(\sbox_aesinv_inst.x0000a000 ),
    .B_N(\sbox_aesinv_inst.me3ab5bd2/_0_ ),
    .Y(\sbox_aesinv_inst.xe3ab5bd2 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.me8133bb7/_0_  (.A1(\sbox_aesinv_inst.x17ff555f ),
    .A2(\sbox_aesinv_inst.xffecece8 ),
    .Y(\sbox_aesinv_inst.xe8133bb7 ),
    .B1(\sbox_aesinv_inst.x00008000 ));
 sg13g2_and3_1 \sbox_aesinv_inst.me8e8e800/_0_  (.X(\sbox_aesinv_inst.xe8e8e800 ),
    .A(\sbox_aesinv_inst.xeaeaeaea ),
    .B(\sbox_aesinv_inst.xfcfcfcfc ),
    .C(\sbox_aesinv_inst.xffffff00 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.meaeaeaea/_0_  (.B1(net333),
    .Y(\sbox_aesinv_inst.xeaeaeaea ),
    .A1(net320),
    .A2(net317));
 sg13g2_nand2b_1 \sbox_aesinv_inst.meaefffff/_0_  (.Y(\sbox_aesinv_inst.xeaefffff ),
    .B(net257),
    .A_N(\sbox_aesinv_inst.xeaeaeaea ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.mee00ee00/_0_  (.A1(net324),
    .A2(net336),
    .Y(\sbox_aesinv_inst.xee00ee00 ),
    .B1(net295));
 sg13g2_o21ai_1 \sbox_aesinv_inst.meeaaeeaa/_0_  (.B1(net338),
    .Y(\sbox_aesinv_inst.xeeaaeeaa ),
    .A1(net325),
    .A2(net297));
 sg13g2_a21oi_1 \sbox_aesinv_inst.meecc98e2/_0_  (.A1(\sbox_aesinv_inst.xffffffdd ),
    .A2(\sbox_aesinv_inst.x0133273f ),
    .Y(\sbox_aesinv_inst.xeecc98e2 ),
    .B1(\sbox_aesinv_inst.x11004400 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.meeee0000/_0_  (.B1(net279),
    .Y(\sbox_aesinv_inst.xeeee0000 ),
    .A2(net335),
    .A1(net323));
 sg13g2_or2_1 \sbox_aesinv_inst.meeee8080/_0_  (.X(\sbox_aesinv_inst.xeeee8080 ),
    .B(\sbox_aesinv_inst.xeeee0000 ),
    .A(net274));
 sg13g2_o21ai_1 \sbox_aesinv_inst.meeeeaaaa/_0_  (.B1(net341),
    .Y(\sbox_aesinv_inst.xeeeeaaaa ),
    .A1(net286),
    .A2(net327));
 sg13g2_nand2_1 \sbox_aesinv_inst.meeeeeeee/_0_  (.Y(\sbox_aesinv_inst.xeeeeeeee ),
    .A(net320),
    .B(net333));
 sg13g2_a21oi_1 \sbox_aesinv_inst.mef715dd5/_0_  (.A1(\sbox_aesinv_inst.x13bfbfbf ),
    .A2(\sbox_aesinv_inst.xfccca000 ),
    .Y(\sbox_aesinv_inst.xef715dd5 ),
    .B1(\sbox_aesinv_inst.x000a022a ));
 sg13g2_or3_1 \sbox_aesinv_inst.mefefcf8f/_0_  (.A(\sbox_aesinv_inst.xcc88cc88 ),
    .B(\sbox_aesinv_inst.xeeee0000 ),
    .C(net308),
    .X(\sbox_aesinv_inst.xefefcf8f ));
 sg13g2_nor3_2 \sbox_aesinv_inst.mf0000000/_0_  (.A(net314),
    .B(net301),
    .C(net287),
    .Y(\sbox_aesinv_inst.xf0000000 ));
 sg13g2_nor2_2 \sbox_aesinv_inst.mf000f000/_0_  (.A(net306),
    .B(net294),
    .Y(\sbox_aesinv_inst.xf000f000 ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mf003f003/_0_  (.Y(\sbox_aesinv_inst.xf003f003 ),
    .B(\sbox_aesinv_inst.xfffcfffc ),
    .A_N(\sbox_aesinv_inst.xf000f000 ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.mf0a0a0a0/_0_  (.A(net314),
    .B_N(\sbox_aesinv_inst.xffaaaaaa ),
    .Y(\sbox_aesinv_inst.xf0a0a0a0 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mf0a0f0a0/_0_  (.B1(net303),
    .Y(\sbox_aesinv_inst.xf0a0f0a0 ),
    .A2(net291),
    .A1(net330));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mf0a0f3a3/_0_  (.Y(\sbox_aesinv_inst.xf0a0f3a3 ),
    .B(\sbox_aesinv_inst.xfffffcfc ),
    .A_N(\sbox_aesinv_inst.xf0a0f0a0 ));
 sg13g2_and2_1 \sbox_aesinv_inst.mf0c0c000/_0_  (.A(\sbox_aesinv_inst.xffcccccc ),
    .B(\sbox_aesinv_inst.xf0f0f000 ),
    .X(\sbox_aesinv_inst.xf0c0c000 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mf0c0f0c0/_0_  (.B1(net303),
    .Y(\sbox_aesinv_inst.xf0c0f0c0 ),
    .A2(net290),
    .A1(net318));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mf0c0f5d5/_0_  (.Y(\sbox_aesinv_inst.xf0c0f5d5 ),
    .B(\sbox_aesinv_inst.xffffaaaa ),
    .A_N(\sbox_aesinv_inst.xf0c0f0c0 ));
 sg13g2_nor2_1 \sbox_aesinv_inst.mf0f00000/_0_  (.A(net275),
    .B(net303),
    .Y(\sbox_aesinv_inst.xf0f00000 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mf0f0a0a0/_0_  (.B1(net313),
    .Y(\sbox_aesinv_inst.xf0f0a0a0 ),
    .A2(net340),
    .A1(net287));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mf0f0c0c0/_0_  (.B1(net315),
    .Y(\sbox_aesinv_inst.xf0f0c0c0 ),
    .A2(net328),
    .A1(net288));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mf0f0f000/_0_  (.B1(net310),
    .Y(\sbox_aesinv_inst.xf0f0f000 ),
    .A2(net298),
    .A1(net285));
 sg13g2_inv_1 \sbox_aesinv_inst.mf0f0f0f0/_0_  (.Y(\sbox_aesinv_inst.xf0f0f0f0 ),
    .A(net304));
 sg13g2_nand2_1 \sbox_aesinv_inst.mf12405c2/_1_  (.Y(\sbox_aesinv_inst.mf12405c2/_0_ ),
    .A(\sbox_aesinv_inst.xf1f5f5f7 ),
    .B(\sbox_aesinv_inst.xff3f05ff ));
 sg13g2_nor2_1 \sbox_aesinv_inst.mf12405c2/_2_  (.A(\sbox_aesinv_inst.x00113035 ),
    .B(\sbox_aesinv_inst.mf12405c2/_0_ ),
    .Y(\sbox_aesinv_inst.xf12405c2 ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mf1a1f1a1/_0_  (.Y(\sbox_aesinv_inst.xf1a1f1a1 ),
    .B(\sbox_aesinv_inst.xfefefefe ),
    .A_N(\sbox_aesinv_inst.xf0a0f0a0 ));
 sg13g2_nand2_1 \sbox_aesinv_inst.mf1f1ffff/_0_  (.Y(\sbox_aesinv_inst.xf1f1ffff ),
    .A(net308),
    .B(\sbox_aesinv_inst.xeeee0000 ));
 sg13g2_nand4_1 \sbox_aesinv_inst.mf1f5f5f7/_0_  (.B(\sbox_aesinv_inst.xeeeeaaaa ),
    .C(net313),
    .A(\sbox_aesinv_inst.xffaaaaaa ),
    .Y(\sbox_aesinv_inst.xf1f5f5f7 ),
    .D(\sbox_aesinv_inst.xffffffcc ));
 sg13g2_or2_1 \sbox_aesinv_inst.mf333f377/_1_  (.X(\sbox_aesinv_inst.mf333f377/_0_ ),
    .B(net293),
    .A(net305));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mf333f377/_2_  (.B1(\sbox_aesinv_inst.mf333f377/_0_ ),
    .Y(\sbox_aesinv_inst.xf333f377 ),
    .A1(\sbox_aesinv_inst.xcccc8888 ),
    .A2(net262));
 sg13g2_or2_1 \sbox_aesinv_inst.mf33fffff/_1_  (.X(\sbox_aesinv_inst.mf33fffff/_0_ ),
    .B(net295),
    .A(net307));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mf33fffff/_2_  (.B1(\sbox_aesinv_inst.mf33fffff/_0_ ),
    .Y(\sbox_aesinv_inst.xf33fffff ),
    .A1(net264),
    .A2(net265));
 sg13g2_or2_1 \sbox_aesinv_inst.mf35ff3ff/_1_  (.X(\sbox_aesinv_inst.mf35ff3ff/_0_ ),
    .B(net300),
    .A(net313));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mf35ff3ff/_2_  (.B1(\sbox_aesinv_inst.mf35ff3ff/_0_ ),
    .Y(\sbox_aesinv_inst.xf35ff3ff ),
    .A1(net262),
    .A2(net268));
 sg13g2_or2_1 \sbox_aesinv_inst.mf3f37f7f/_1_  (.X(\sbox_aesinv_inst.mf3f37f7f/_0_ ),
    .B(net284),
    .A(net309));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mf3f37f7f/_2_  (.B1(\sbox_aesinv_inst.mf3f37f7f/_0_ ),
    .Y(\sbox_aesinv_inst.xf3f37f7f ),
    .A1(net260),
    .A2(net274));
 sg13g2_a21oi_1 \sbox_aesinv_inst.mf446ce08/_0_  (.A1(\sbox_aesinv_inst.xb1b1f5f7 ),
    .A2(\sbox_aesinv_inst.x01f731f7 ),
    .Y(\sbox_aesinv_inst.xf446ce08 ),
    .B1(\sbox_aesinv_inst.x0a080000 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.mf4bcfdb0/_0_  (.A1(\sbox_aesinv_inst.xc3c3c3cf ),
    .A2(\sbox_aesinv_inst.x0f5f0a5f ),
    .Y(\sbox_aesinv_inst.xf4bcfdb0 ),
    .B1(\sbox_aesinv_inst.x0a000000 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mf555f57f/_1_  (.X(\sbox_aesinv_inst.mf555f57f/_0_ ),
    .B(net294),
    .A(net306));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mf555f57f/_2_  (.B1(\sbox_aesinv_inst.mf555f57f/_0_ ),
    .Y(\sbox_aesinv_inst.xf555f57f ),
    .A1(\sbox_aesinv_inst.xaaaaaa00 ),
    .A2(net274));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mf5a5ffff/_0_  (.Y(\sbox_aesinv_inst.xf5a5ffff ),
    .B(\sbox_aesinv_inst.xfafa0000 ),
    .A_N(\sbox_aesinv_inst.xf0a0f0a0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mf5ff5fff/_1_  (.X(\sbox_aesinv_inst.mf5ff5fff/_0_ ),
    .B(net279),
    .A(net306));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mf5ff5fff/_2_  (.B1(\sbox_aesinv_inst.mf5ff5fff/_0_ ),
    .Y(\sbox_aesinv_inst.xf5ff5fff ),
    .A1(net267),
    .A2(net269));
 sg13g2_and3_1 \sbox_aesinv_inst.mf8008000/_0_  (.X(\sbox_aesinv_inst.xf8008000 ),
    .A(\sbox_aesinv_inst.xfcfccccc ),
    .B(\sbox_aesinv_inst.xff00f000 ),
    .C(\sbox_aesinv_inst.xfafaaaaa ));
 sg13g2_or3_1 \sbox_aesinv_inst.mf8f0c800/_0_  (.A(net272),
    .B(\sbox_aesinv_inst.xf0f00000 ),
    .C(\sbox_aesinv_inst.xc000c000 ),
    .X(\sbox_aesinv_inst.xf8f0c800 ));
 sg13g2_and2_1 \sbox_aesinv_inst.mf8f8c8c8/_0_  (.A(\sbox_aesinv_inst.xfafafafa ),
    .B(\sbox_aesinv_inst.xfcfccccc ),
    .X(\sbox_aesinv_inst.xf8f8c8c8 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mfa00fa00/_0_  (.B1(net300),
    .Y(\sbox_aesinv_inst.xfa00fa00 ),
    .A2(net341),
    .A1(net314));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mfaaafaaa/_0_  (.B1(net340),
    .Y(\sbox_aesinv_inst.xfaaafaaa ),
    .A1(net313),
    .A2(net300));
 sg13g2_and3_1 \sbox_aesinv_inst.mfac8a080/_0_  (.X(\sbox_aesinv_inst.xfac8a080 ),
    .A(\sbox_aesinv_inst.xfafaaaaa ),
    .B(\sbox_aesinv_inst.xfffff0f0 ),
    .C(\sbox_aesinv_inst.xffccffcc ));
 sg13g2_and3_1 \sbox_aesinv_inst.mfaf8fa00/_0_  (.X(\sbox_aesinv_inst.xfaf8fa00 ),
    .A(\sbox_aesinv_inst.xffffff00 ),
    .B(\sbox_aesinv_inst.xfafafafa ),
    .C(\sbox_aesinv_inst.xfffcfffc ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mfafa0000/_0_  (.B1(net277),
    .Y(\sbox_aesinv_inst.xfafa0000 ),
    .A2(net332),
    .A1(net305));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mfafaaaaa/_0_  (.B1(net339),
    .Y(\sbox_aesinv_inst.xfafaaaaa ),
    .A1(net283),
    .A2(net311));
 sg13g2_nand2_1 \sbox_aesinv_inst.mfafafafa/_0_  (.Y(\sbox_aesinv_inst.xfafafafa ),
    .A(net305),
    .B(net333));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mfc00fc00/_0_  (.B1(net294),
    .Y(\sbox_aesinv_inst.xfc00fc00 ),
    .A2(net306),
    .A1(net322));
 sg13g2_or3_1 \sbox_aesinv_inst.mfccca000/_0_  (.A(net269),
    .B(\sbox_aesinv_inst.xcccc0000 ),
    .C(\sbox_aesinv_inst.xf0000000 ),
    .X(\sbox_aesinv_inst.xfccca000 ));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mfcccfccc/_0_  (.B1(net326),
    .Y(\sbox_aesinv_inst.xfcccfccc ),
    .A1(net311),
    .A2(net296));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mfccfffff/_0_  (.Y(\sbox_aesinv_inst.xfccfffff ),
    .B(\sbox_aesinv_inst.xfff00000 ),
    .A_N(\sbox_aesinv_inst.xfcccfccc ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfcecf8a0/_0_  (.A(net272),
    .B(\sbox_aesinv_inst.xcccc0000 ),
    .C(\sbox_aesinv_inst.xf0a0f0a0 ),
    .X(\sbox_aesinv_inst.xfcecf8a0 ));
 sg13g2_a21oi_1 \sbox_aesinv_inst.mfcfc0000/_0_  (.A1(net325),
    .A2(net309),
    .Y(\sbox_aesinv_inst.xfcfc0000 ),
    .B1(net284));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mfcfccccc/_0_  (.B1(net326),
    .Y(\sbox_aesinv_inst.xfcfccccc ),
    .A1(net282),
    .A2(net311));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mfcfcccff/_0_  (.Y(\sbox_aesinv_inst.xfcfcccff ),
    .B(\sbox_aesinv_inst.xffffff00 ),
    .A_N(\sbox_aesinv_inst.xfcfccccc ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfcfcf8a0/_0_  (.A(net272),
    .B(net259),
    .C(\sbox_aesinv_inst.xf0a0f0a0 ),
    .X(\sbox_aesinv_inst.xfcfcf8a0 ));
 sg13g2_nand2_1 \sbox_aesinv_inst.mfcfcfcfc/_0_  (.Y(\sbox_aesinv_inst.xfcfcfcfc ),
    .A(net320),
    .B(net305));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mfd11ffff/_0_  (.Y(\sbox_aesinv_inst.xfd11ffff ),
    .B(\sbox_aesinv_inst.xeeee0000 ),
    .A_N(\sbox_aesinv_inst.xfc00fc00 ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfec8eec8/_0_  (.A(\sbox_aesinv_inst.xccc0ccc0 ),
    .B(\sbox_aesinv_inst.xf0000000 ),
    .C(\sbox_aesinv_inst.xaa88aa88 ),
    .X(\sbox_aesinv_inst.xfec8eec8 ));
 sg13g2_and3_1 \sbox_aesinv_inst.mfecccc00/_0_  (.X(\sbox_aesinv_inst.xfecccc00 ),
    .A(\sbox_aesinv_inst.xfefefefe ),
    .B(\sbox_aesinv_inst.xffcccccc ),
    .C(\sbox_aesinv_inst.xffffff00 ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfeccfec8/_0_  (.A(\sbox_aesinv_inst.xccccc0c0 ),
    .B(\sbox_aesinv_inst.xfc00fc00 ),
    .C(\sbox_aesinv_inst.xaa88aa88 ),
    .X(\sbox_aesinv_inst.xfeccfec8 ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfeecfaa8/_0_  (.A(\sbox_aesinv_inst.xcccc8888 ),
    .B(\sbox_aesinv_inst.xf000f000 ),
    .C(\sbox_aesinv_inst.xaaa0aaa0 ),
    .X(\sbox_aesinv_inst.xfeecfaa8 ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfeeef8a8/_0_  (.A(\sbox_aesinv_inst.xeeee0000 ),
    .B(\sbox_aesinv_inst.xf000f000 ),
    .C(\sbox_aesinv_inst.xa8a8a8a8 ),
    .X(\sbox_aesinv_inst.xfeeef8a8 ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfefaeca8/_0_  (.A(\sbox_aesinv_inst.xfafa0000 ),
    .B(net262),
    .C(\sbox_aesinv_inst.xa8a8a8a8 ),
    .X(\sbox_aesinv_inst.xfefaeca8 ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mfefafefa/_0_  (.Y(\sbox_aesinv_inst.xfefafefa ),
    .B(net309),
    .A_N(\sbox_aesinv_inst.xeeaaeeaa ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfefea8a0/_0_  (.A(net273),
    .B(net260),
    .C(\sbox_aesinv_inst.xaaaaa0a0 ),
    .X(\sbox_aesinv_inst.xfefea8a0 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.mfefefefe/_0_  (.B(net333),
    .C(net320),
    .A(net305),
    .Y(\sbox_aesinv_inst.xfefefefe ));
 sg13g2_nor2_1 \sbox_aesinv_inst.mff000000/_0_  (.A(net279),
    .B(net295),
    .Y(\sbox_aesinv_inst.xff000000 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mff00aa00/_0_  (.B1(net295),
    .Y(\sbox_aesinv_inst.xff00aa00 ),
    .A2(net334),
    .A1(net279));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mff00cc00/_0_  (.B1(net290),
    .Y(\sbox_aesinv_inst.xff00cc00 ),
    .A2(net318),
    .A1(net275));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mff00f000/_0_  (.B1(net297),
    .Y(\sbox_aesinv_inst.xff00f000 ),
    .A2(net310),
    .A1(net284));
 sg13g2_inv_2 \sbox_aesinv_inst.mff00ff00/_0_  (.Y(\sbox_aesinv_inst.xff00ff00 ),
    .A(net296));
 sg13g2_or2_1 \sbox_aesinv_inst.mff010103/_1_  (.X(\sbox_aesinv_inst.mff010103/_0_ ),
    .B(net278),
    .A(net293));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mff010103/_2_  (.B1(\sbox_aesinv_inst.mff010103/_0_ ),
    .Y(\sbox_aesinv_inst.xff010103 ),
    .A1(\sbox_aesinv_inst.xfcfcfcfc ),
    .A2(\sbox_aesinv_inst.xaaaaaa00 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mff05333f/_1_  (.X(\sbox_aesinv_inst.mff05333f/_0_ ),
    .B(net277),
    .A(net292));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mff05333f/_2_  (.B1(\sbox_aesinv_inst.mff05333f/_0_ ),
    .Y(\sbox_aesinv_inst.xff05333f ),
    .A1(\sbox_aesinv_inst.xfafa0000 ),
    .A2(\sbox_aesinv_inst.xccc0ccc0 ));
 sg13g2_or2_1 \sbox_aesinv_inst.mff3f05ff/_1_  (.X(\sbox_aesinv_inst.mff3f05ff/_0_ ),
    .B(net286),
    .A(net301));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mff3f05ff/_2_  (.B1(\sbox_aesinv_inst.mff3f05ff/_0_ ),
    .Y(\sbox_aesinv_inst.xff3f05ff ),
    .A1(\sbox_aesinv_inst.xfa00fa00 ),
    .A2(net266));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mff7f7f7f/_0_  (.Y(\sbox_aesinv_inst.xff7f7f7f ),
    .B(net274),
    .A_N(net263));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mffaa0000/_0_  (.B1(net275),
    .Y(\sbox_aesinv_inst.xffaa0000 ),
    .A2(net290),
    .A1(net330));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mffaaaaaa/_0_  (.B1(net341),
    .Y(\sbox_aesinv_inst.xffaaaaaa ),
    .A1(net286),
    .A2(net300));
 sg13g2_nand2_1 \sbox_aesinv_inst.mffaaffaa/_0_  (.Y(\sbox_aesinv_inst.xffaaffaa ),
    .A(net340),
    .B(net301));
 sg13g2_or3_1 \sbox_aesinv_inst.mffb3ffb3/_0_  (.A(net274),
    .B(net262),
    .C(net324),
    .X(\sbox_aesinv_inst.xffb3ffb3 ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mffcc0000/_0_  (.B1(net282),
    .Y(\sbox_aesinv_inst.xffcc0000 ),
    .A2(net296),
    .A1(net326));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mffcccccc/_0_  (.B1(net325),
    .Y(\sbox_aesinv_inst.xffcccccc ),
    .A1(net284),
    .A2(net297));
 sg13g2_or3_1 \sbox_aesinv_inst.mffcceec8/_0_  (.A(\sbox_aesinv_inst.xccccc0c0 ),
    .B(net258),
    .C(\sbox_aesinv_inst.xaa88aa88 ),
    .X(\sbox_aesinv_inst.xffcceec8 ));
 sg13g2_nand2_2 \sbox_aesinv_inst.mffccffcc/_0_  (.Y(\sbox_aesinv_inst.xffccffcc ),
    .A(net321),
    .B(net293));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mffddddff/_0_  (.Y(\sbox_aesinv_inst.xffddddff ),
    .B(\sbox_aesinv_inst.xaaaaaa00 ),
    .A_N(\sbox_aesinv_inst.xffcccccc ));
 sg13g2_or3_1 \sbox_aesinv_inst.mffec8888/_0_  (.A(net268),
    .B(\sbox_aesinv_inst.xff000000 ),
    .C(\sbox_aesinv_inst.xcccc8888 ),
    .X(\sbox_aesinv_inst.xffec8888 ));
 sg13g2_or3_1 \sbox_aesinv_inst.mffecece8/_0_  (.A(\sbox_aesinv_inst.xcccc8888 ),
    .B(net258),
    .C(\sbox_aesinv_inst.xe0e0e0e0 ),
    .X(\sbox_aesinv_inst.xffecece8 ));
 sg13g2_and3_1 \sbox_aesinv_inst.mffecffa8/_0_  (.X(\sbox_aesinv_inst.xffecffa8 ),
    .A(\sbox_aesinv_inst.xffeeffee ),
    .B(\sbox_aesinv_inst.xffffffaa ),
    .C(\sbox_aesinv_inst.xfffcfffc ));
 sg13g2_or3_1 \sbox_aesinv_inst.mffeeee88/_0_  (.A(net261),
    .B(\sbox_aesinv_inst.xffaa0000 ),
    .C(\sbox_aesinv_inst.xaa88aa88 ),
    .X(\sbox_aesinv_inst.xffeeee88 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.mffeeffee/_0_  (.B(net302),
    .C(net320),
    .A(net333),
    .Y(\sbox_aesinv_inst.xffeeffee ));
 sg13g2_a21oi_2 \sbox_aesinv_inst.mfff00000/_0_  (.B1(net284),
    .Y(\sbox_aesinv_inst.xfff00000 ),
    .A2(net297),
    .A1(net309));
 sg13g2_o21ai_1 \sbox_aesinv_inst.mfff0f0f0/_0_  (.B1(net304),
    .Y(\sbox_aesinv_inst.xfff0f0f0 ),
    .A1(net277),
    .A2(net292));
 sg13g2_nand2_1 \sbox_aesinv_inst.mfff0fff0/_0_  (.Y(\sbox_aesinv_inst.xfff0fff0 ),
    .A(net313),
    .B(net300));
 sg13g2_nand3_1 \sbox_aesinv_inst.mfff30000/_1_  (.B(net259),
    .C(net305),
    .A(net293),
    .Y(\sbox_aesinv_inst.mfff30000/_0_ ));
 sg13g2_nor2b_1 \sbox_aesinv_inst.mfff30000/_2_  (.A(net278),
    .B_N(\sbox_aesinv_inst.mfff30000/_0_ ),
    .Y(\sbox_aesinv_inst.xfff30000 ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mfff5f5ff/_0_  (.Y(\sbox_aesinv_inst.xfff5f5ff ),
    .B(\sbox_aesinv_inst.xaaaaaa00 ),
    .A_N(\sbox_aesinv_inst.xfff0f0f0 ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfff8fac8/_0_  (.A(\sbox_aesinv_inst.xf0c0f0c0 ),
    .B(net257),
    .C(\sbox_aesinv_inst.xaa88aa88 ),
    .X(\sbox_aesinv_inst.xfff8fac8 ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfff8ffa0/_0_  (.A(\sbox_aesinv_inst.xf0f0a0a0 ),
    .B(net271),
    .C(\sbox_aesinv_inst.xff00ff00 ),
    .X(\sbox_aesinv_inst.xfff8ffa0 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.mfffafffa/_0_  (.B(net301),
    .C(net312),
    .A(net342),
    .Y(\sbox_aesinv_inst.xfffafffa ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfffcfeec/_0_  (.A(\sbox_aesinv_inst.xffcccccc ),
    .B(\sbox_aesinv_inst.xf0f0f000 ),
    .C(\sbox_aesinv_inst.xaaa0aaa0 ),
    .X(\sbox_aesinv_inst.xfffcfeec ));
 sg13g2_nand3_1 \sbox_aesinv_inst.mfffcfffc/_0_  (.B(net290),
    .C(net318),
    .A(net303),
    .Y(\sbox_aesinv_inst.xfffcfffc ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mfffcfffd/_0_  (.Y(\sbox_aesinv_inst.xfffcfffd ),
    .B(\sbox_aesinv_inst.xffffaaaa ),
    .A_N(\sbox_aesinv_inst.xfffcfffc ));
 sg13g2_or3_1 \sbox_aesinv_inst.mfffef888/_0_  (.A(\sbox_aesinv_inst.xff00f000 ),
    .B(net260),
    .C(\sbox_aesinv_inst.xaaaa8888 ),
    .X(\sbox_aesinv_inst.xfffef888 ));
 sg13g2_inv_1 \sbox_aesinv_inst.mffff0000/_0_  (.Y(\sbox_aesinv_inst.xffff0000 ),
    .A(net279));
 sg13g2_or3_1 \sbox_aesinv_inst.mffff8f0f/_0_  (.A(net272),
    .B(net259),
    .C(net312),
    .X(\sbox_aesinv_inst.xffff8f0f ));
 sg13g2_nand2_2 \sbox_aesinv_inst.mffffaaaa/_0_  (.Y(\sbox_aesinv_inst.xffffaaaa ),
    .A(net277),
    .B(net332));
 sg13g2_nand2_1 \sbox_aesinv_inst.mffffcccc/_0_  (.Y(\sbox_aesinv_inst.xffffcccc ),
    .A(net288),
    .B(net328));
 sg13g2_nand3_1 \sbox_aesinv_inst.mffffeeee/_0_  (.B(net342),
    .C(net288),
    .A(net328),
    .Y(\sbox_aesinv_inst.xffffeeee ));
 sg13g2_nand2_2 \sbox_aesinv_inst.mfffff0f0/_0_  (.Y(\sbox_aesinv_inst.xfffff0f0 ),
    .A(net276),
    .B(net303));
 sg13g2_or3_1 \sbox_aesinv_inst.mfffff8a0/_0_  (.A(net272),
    .B(\sbox_aesinv_inst.xffff0000 ),
    .C(\sbox_aesinv_inst.xf0a0f0a0 ),
    .X(\sbox_aesinv_inst.xfffff8a0 ));
 sg13g2_nand3_1 \sbox_aesinv_inst.mfffffafa/_0_  (.B(net339),
    .C(net282),
    .A(net311),
    .Y(\sbox_aesinv_inst.xfffffafa ));
 sg13g2_nand3_1 \sbox_aesinv_inst.mfffffcfc/_0_  (.B(net304),
    .C(net276),
    .A(net319),
    .Y(\sbox_aesinv_inst.xfffffcfc ));
 sg13g2_or2_1 \sbox_aesinv_inst.mfffffeee/_0_  (.X(\sbox_aesinv_inst.xfffffeee ),
    .B(\sbox_aesinv_inst.xf0f0f000 ),
    .A(\sbox_aesinv_inst.xffffeeee ));
 sg13g2_nand2_2 \sbox_aesinv_inst.mffffff00/_0_  (.Y(\sbox_aesinv_inst.xffffff00 ),
    .A(net278),
    .B(net293));
 sg13g2_nand3_1 \sbox_aesinv_inst.mffffffaa/_0_  (.B(net290),
    .C(net275),
    .A(net330),
    .Y(\sbox_aesinv_inst.xffffffaa ));
 sg13g2_nand3_1 \sbox_aesinv_inst.mffffffcc/_0_  (.B(net300),
    .C(net287),
    .A(net327),
    .Y(\sbox_aesinv_inst.xffffffcc ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mffffffdd/_0_  (.Y(\sbox_aesinv_inst.xffffffdd ),
    .B(\sbox_aesinv_inst.xeeeeaaaa ),
    .A_N(\sbox_aesinv_inst.xffffffcc ));
 sg13g2_or2_1 \sbox_aesinv_inst.mffffffea/_0_  (.X(\sbox_aesinv_inst.xffffffea ),
    .B(\sbox_aesinv_inst.xf0f0c0c0 ),
    .A(\sbox_aesinv_inst.xffffffaa ));
 sg13g2_or2_1 \sbox_aesinv_inst.mffffffec/_0_  (.X(\sbox_aesinv_inst.xffffffec ),
    .B(\sbox_aesinv_inst.xf0f0a0a0 ),
    .A(\sbox_aesinv_inst.xffffffcc ));
 sg13g2_nand3_1 \sbox_aesinv_inst.mfffffff0/_0_  (.B(net296),
    .C(net282),
    .A(net311),
    .Y(\sbox_aesinv_inst.xfffffff0 ));
 sg13g2_nand2b_1 \sbox_aesinv_inst.mfffffffc/_0_  (.Y(\sbox_aesinv_inst.xfffffffc ),
    .B(net292),
    .A_N(\sbox_aesinv_inst.xfffffcfc ));
 sg13g2_or2_1 \sbox_aesinv_inst.mfffffffe/_0_  (.X(\sbox_aesinv_inst.xfffffffe ),
    .B(\sbox_aesinv_inst.xffffcccc ),
    .A(\sbox_aesinv_inst.xfffafffa ));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(\sbox_aesinv_inst.xfff00000 ));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(\sbox_aesinv_inst.xff00cc00 ));
 sg13g2_buf_2 fanout259 (.A(net260),
    .X(net259));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(\sbox_aesinv_inst.xfcfc0000 ));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(\sbox_aesinv_inst.xcccccc00 ));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(\sbox_aesinv_inst.xcc00cc00 ));
 sg13g2_buf_2 fanout263 (.A(\sbox_aesinv_inst.xcc000000 ),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(\sbox_aesinv_inst.xcc000000 ),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(net266),
    .X(net265));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(\sbox_aesinv_inst.xc0c00000 ));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(\sbox_aesinv_inst.xaa000000 ));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(\sbox_aesinv_inst.xa0a00000 ));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(\sbox_aesinv_inst.xa000a000 ));
 sg13g2_buf_2 fanout270 (.A(\sbox_aesinv_inst.xa000a000 ),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(\sbox_aesinv_inst.x88880000 ),
    .X(net271));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(\sbox_aesinv_inst.x88008800 ));
 sg13g2_buf_1 fanout273 (.A(\sbox_aesinv_inst.x88008800 ),
    .X(net273));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(\sbox_aesinv_inst.x80808080 ));
 sg13g2_buf_2 fanout275 (.A(net276),
    .X(net275));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(net278));
 sg13g2_buf_1 fanout277 (.A(net278),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(ui_in[4]),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(ui_in[4]),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(net283),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(net289),
    .X(net283));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(net289));
 sg13g2_buf_1 fanout285 (.A(net289),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(net288),
    .X(net286));
 sg13g2_buf_1 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_1 fanout289 (.A(ui_in[4]),
    .X(net289));
 sg13g2_buf_4 fanout290 (.X(net290),
    .A(net291));
 sg13g2_buf_2 fanout291 (.A(net292),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(net293),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net302),
    .X(net293));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(net295));
 sg13g2_buf_2 fanout295 (.A(net302),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(net299),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(net299),
    .X(net297));
 sg13g2_buf_1 fanout298 (.A(net299),
    .X(net298));
 sg13g2_buf_1 fanout299 (.A(net302),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(net301),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(net302),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(ui_in[3]),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(net304),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(net305),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(net317),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(net307),
    .X(net306));
 sg13g2_buf_1 fanout307 (.A(net308),
    .X(net307));
 sg13g2_buf_4 fanout308 (.X(net308),
    .A(net317));
 sg13g2_buf_2 fanout309 (.A(net316),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(net316),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(net316),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net315),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net315),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(net315),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(net316),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(ui_in[2]),
    .X(net317));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(net321));
 sg13g2_buf_1 fanout319 (.A(net321),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(net321),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(ui_in[1]),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(net324),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(ui_in[1]),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(net329),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(net329),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(net329),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(ui_in[1]),
    .X(net329));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(net332));
 sg13g2_buf_1 fanout331 (.A(net332),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(net337),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(net337),
    .X(net333));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(net336));
 sg13g2_buf_2 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(net337),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(ui_in[0]),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(net339),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(ui_in[0]),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(net342),
    .X(net340));
 sg13g2_buf_1 fanout341 (.A(net342),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(ui_in[0]),
    .X(net342));
 sg13g2_buf_4 input1 (.X(net1),
    .A(ui_in[5]));
 sg13g2_buf_2 input2 (.A(ui_in[6]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[7]),
    .X(net3));
 sg13g2_tiehi _22__4 (.L_HI(net4));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_250 ();
 sg13g2_decap_4 FILLER_16_257 ();
 sg13g2_fill_2 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_282 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_decap_8 FILLER_16_296 ();
 sg13g2_decap_8 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_155 ();
 sg13g2_decap_8 FILLER_17_162 ();
 sg13g2_decap_4 FILLER_17_169 ();
 sg13g2_fill_1 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_187 ();
 sg13g2_decap_4 FILLER_17_194 ();
 sg13g2_fill_1 FILLER_17_208 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_decap_4 FILLER_17_221 ();
 sg13g2_fill_1 FILLER_17_225 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_280 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_fill_2 FILLER_17_288 ();
 sg13g2_decap_4 FILLER_17_295 ();
 sg13g2_fill_2 FILLER_17_304 ();
 sg13g2_fill_1 FILLER_17_306 ();
 sg13g2_decap_4 FILLER_17_312 ();
 sg13g2_fill_1 FILLER_17_316 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_4 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_144 ();
 sg13g2_fill_2 FILLER_18_184 ();
 sg13g2_fill_1 FILLER_18_186 ();
 sg13g2_fill_2 FILLER_18_210 ();
 sg13g2_fill_1 FILLER_18_217 ();
 sg13g2_decap_4 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_242 ();
 sg13g2_fill_2 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_279 ();
 sg13g2_decap_4 FILLER_18_300 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_decap_4 FILLER_18_334 ();
 sg13g2_fill_2 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_4 FILLER_19_145 ();
 sg13g2_fill_1 FILLER_19_149 ();
 sg13g2_decap_8 FILLER_19_159 ();
 sg13g2_fill_2 FILLER_19_166 ();
 sg13g2_fill_2 FILLER_19_176 ();
 sg13g2_fill_1 FILLER_19_178 ();
 sg13g2_decap_4 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_232 ();
 sg13g2_decap_4 FILLER_19_239 ();
 sg13g2_fill_2 FILLER_19_253 ();
 sg13g2_decap_4 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_4 FILLER_19_302 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_decap_4 FILLER_19_317 ();
 sg13g2_decap_4 FILLER_19_345 ();
 sg13g2_fill_2 FILLER_19_362 ();
 sg13g2_fill_2 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_fill_2 FILLER_20_149 ();
 sg13g2_fill_2 FILLER_20_156 ();
 sg13g2_fill_2 FILLER_20_171 ();
 sg13g2_decap_4 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_211 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_220 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_decap_4 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_268 ();
 sg13g2_decap_4 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_306 ();
 sg13g2_decap_4 FILLER_20_327 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_fill_1 FILLER_20_340 ();
 sg13g2_decap_4 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_4 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_130 ();
 sg13g2_fill_2 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_147 ();
 sg13g2_fill_1 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_192 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_decap_4 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_decap_4 FILLER_21_239 ();
 sg13g2_fill_1 FILLER_21_258 ();
 sg13g2_fill_2 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_292 ();
 sg13g2_decap_4 FILLER_21_306 ();
 sg13g2_fill_2 FILLER_21_310 ();
 sg13g2_fill_1 FILLER_21_317 ();
 sg13g2_fill_2 FILLER_21_323 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_fill_1 FILLER_21_337 ();
 sg13g2_decap_4 FILLER_21_346 ();
 sg13g2_fill_2 FILLER_21_350 ();
 sg13g2_decap_4 FILLER_21_357 ();
 sg13g2_decap_4 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_163 ();
 sg13g2_fill_2 FILLER_22_170 ();
 sg13g2_decap_8 FILLER_22_177 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_decap_4 FILLER_22_191 ();
 sg13g2_fill_1 FILLER_22_195 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_decap_4 FILLER_22_211 ();
 sg13g2_fill_2 FILLER_22_215 ();
 sg13g2_fill_1 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_239 ();
 sg13g2_fill_1 FILLER_22_241 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_4 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_285 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_fill_1 FILLER_22_294 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_2 FILLER_22_321 ();
 sg13g2_fill_1 FILLER_22_323 ();
 sg13g2_decap_4 FILLER_22_341 ();
 sg13g2_fill_2 FILLER_22_357 ();
 sg13g2_fill_1 FILLER_22_359 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_fill_2 FILLER_23_133 ();
 sg13g2_fill_1 FILLER_23_164 ();
 sg13g2_decap_4 FILLER_23_185 ();
 sg13g2_fill_2 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_fill_2 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_229 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_261 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_decap_4 FILLER_23_284 ();
 sg13g2_fill_2 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_324 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_fill_2 FILLER_23_341 ();
 sg13g2_fill_2 FILLER_23_348 ();
 sg13g2_fill_2 FILLER_23_365 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_4 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_decap_4 FILLER_24_166 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_fill_1 FILLER_24_181 ();
 sg13g2_decap_4 FILLER_24_207 ();
 sg13g2_fill_2 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_218 ();
 sg13g2_decap_4 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_240 ();
 sg13g2_fill_1 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_decap_4 FILLER_24_262 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_fill_2 FILLER_24_280 ();
 sg13g2_fill_1 FILLER_24_282 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_decap_4 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_326 ();
 sg13g2_fill_1 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_334 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_347 ();
 sg13g2_fill_2 FILLER_24_363 ();
 sg13g2_fill_2 FILLER_24_370 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_133 ();
 sg13g2_fill_1 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_152 ();
 sg13g2_fill_1 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_187 ();
 sg13g2_decap_8 FILLER_25_201 ();
 sg13g2_fill_2 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_214 ();
 sg13g2_fill_1 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_fill_1 FILLER_25_289 ();
 sg13g2_decap_4 FILLER_25_307 ();
 sg13g2_decap_4 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_decap_4 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_fill_1 FILLER_25_351 ();
 sg13g2_fill_2 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_153 ();
 sg13g2_fill_2 FILLER_26_160 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_decap_4 FILLER_26_193 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_decap_4 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_223 ();
 sg13g2_decap_4 FILLER_26_230 ();
 sg13g2_fill_2 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_246 ();
 sg13g2_decap_4 FILLER_26_254 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_decap_4 FILLER_26_279 ();
 sg13g2_fill_1 FILLER_26_289 ();
 sg13g2_decap_4 FILLER_26_301 ();
 sg13g2_decap_4 FILLER_26_317 ();
 sg13g2_fill_1 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_fill_2 FILLER_26_376 ();
 sg13g2_fill_1 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_fill_2 FILLER_27_148 ();
 sg13g2_fill_2 FILLER_27_167 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_2 FILLER_27_190 ();
 sg13g2_fill_2 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_decap_4 FILLER_27_232 ();
 sg13g2_fill_1 FILLER_27_236 ();
 sg13g2_decap_4 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_277 ();
 sg13g2_decap_4 FILLER_27_291 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_303 ();
 sg13g2_decap_4 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_314 ();
 sg13g2_decap_4 FILLER_27_333 ();
 sg13g2_fill_1 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_348 ();
 sg13g2_fill_1 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_4 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_137 ();
 sg13g2_fill_1 FILLER_28_144 ();
 sg13g2_decap_4 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_171 ();
 sg13g2_fill_2 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_decap_4 FILLER_28_217 ();
 sg13g2_decap_4 FILLER_28_236 ();
 sg13g2_fill_2 FILLER_28_245 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_decap_8 FILLER_28_288 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_decap_4 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_decap_4 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_decap_4 FILLER_29_151 ();
 sg13g2_fill_2 FILLER_29_155 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_decap_4 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_206 ();
 sg13g2_decap_4 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_240 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_decap_4 FILLER_29_261 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_fill_2 FILLER_29_294 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_fill_2 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_4 FILLER_29_331 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_166 ();
 sg13g2_decap_4 FILLER_30_185 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_decap_4 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_220 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_239 ();
 sg13g2_fill_2 FILLER_30_243 ();
 sg13g2_decap_4 FILLER_30_250 ();
 sg13g2_decap_8 FILLER_30_281 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_2 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_324 ();
 sg13g2_fill_2 FILLER_30_350 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_decap_4 FILLER_30_365 ();
 sg13g2_fill_2 FILLER_30_369 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_150 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_194 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_decap_4 FILLER_31_257 ();
 sg13g2_fill_2 FILLER_31_261 ();
 sg13g2_decap_4 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_271 ();
 sg13g2_fill_2 FILLER_31_290 ();
 sg13g2_fill_1 FILLER_31_292 ();
 sg13g2_decap_8 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_330 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_367 ();
 sg13g2_fill_1 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_133 ();
 sg13g2_decap_4 FILLER_32_201 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_fill_2 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_decap_4 FILLER_32_230 ();
 sg13g2_decap_4 FILLER_32_241 ();
 sg13g2_fill_2 FILLER_32_245 ();
 sg13g2_fill_1 FILLER_32_257 ();
 sg13g2_fill_2 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_289 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_decap_8 FILLER_32_313 ();
 sg13g2_fill_2 FILLER_32_320 ();
 sg13g2_decap_4 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_334 ();
 sg13g2_fill_1 FILLER_32_341 ();
 sg13g2_decap_4 FILLER_32_347 ();
 sg13g2_fill_2 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_362 ();
 sg13g2_fill_2 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_4 FILLER_33_133 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_decap_8 FILLER_33_156 ();
 sg13g2_fill_1 FILLER_33_163 ();
 sg13g2_fill_2 FILLER_33_191 ();
 sg13g2_decap_4 FILLER_33_208 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_fill_2 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_260 ();
 sg13g2_decap_4 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_271 ();
 sg13g2_decap_4 FILLER_33_276 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_291 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_352 ();
 sg13g2_fill_2 FILLER_33_359 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_decap_4 FILLER_34_172 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_decap_4 FILLER_34_185 ();
 sg13g2_decap_8 FILLER_34_197 ();
 sg13g2_decap_4 FILLER_34_214 ();
 sg13g2_fill_2 FILLER_34_234 ();
 sg13g2_fill_2 FILLER_34_242 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_257 ();
 sg13g2_decap_4 FILLER_34_267 ();
 sg13g2_fill_1 FILLER_34_271 ();
 sg13g2_decap_4 FILLER_34_295 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_fill_2 FILLER_34_305 ();
 sg13g2_decap_4 FILLER_34_317 ();
 sg13g2_fill_2 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_343 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_217 ();
 sg13g2_fill_1 FILLER_35_219 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_235 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_249 ();
 sg13g2_fill_2 FILLER_35_275 ();
 sg13g2_fill_1 FILLER_35_277 ();
 sg13g2_fill_2 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_342 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_decap_8 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_379 ();
 sg13g2_decap_8 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_fill_2 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_decap_4 FILLER_36_319 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_decap_8 FILLER_36_367 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_4 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_278 ();
 sg13g2_fill_2 FILLER_37_285 ();
 sg13g2_fill_2 FILLER_37_308 ();
 sg13g2_fill_1 FILLER_37_310 ();
 sg13g2_decap_8 FILLER_37_337 ();
 sg13g2_decap_8 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_123 ();
 sg13g2_decap_8 FILLER_38_130 ();
 sg13g2_decap_8 FILLER_38_137 ();
 sg13g2_decap_8 FILLER_38_144 ();
 sg13g2_decap_8 FILLER_38_151 ();
 sg13g2_decap_8 FILLER_38_158 ();
 sg13g2_decap_8 FILLER_38_165 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_decap_8 FILLER_38_186 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_decap_8 FILLER_38_228 ();
 sg13g2_fill_2 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_248 ();
 sg13g2_fill_2 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_262 ();
 sg13g2_decap_8 FILLER_38_267 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_285 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net12;
 assign uio_oe[1] = net13;
 assign uio_oe[2] = net14;
 assign uio_oe[3] = net15;
 assign uio_oe[4] = net16;
 assign uio_oe[5] = net17;
 assign uio_oe[6] = net18;
 assign uio_oe[7] = net19;
endmodule

module tt_um_obriensp_jtag (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire \bsr.reset_i ;
 wire \bsr.update_data_i[0] ;
 wire \bsr.update_data_i[10] ;
 wire \bsr.update_data_i[11] ;
 wire \bsr.update_data_i[12] ;
 wire \bsr.update_data_i[13] ;
 wire \bsr.update_data_i[14] ;
 wire \bsr.update_data_i[15] ;
 wire \bsr.update_data_i[16] ;
 wire \bsr.update_data_i[17] ;
 wire \bsr.update_data_i[18] ;
 wire \bsr.update_data_i[19] ;
 wire \bsr.update_data_i[1] ;
 wire \bsr.update_data_i[20] ;
 wire \bsr.update_data_i[21] ;
 wire \bsr.update_data_i[22] ;
 wire \bsr.update_data_i[23] ;
 wire \bsr.update_data_i[24] ;
 wire \bsr.update_data_i[25] ;
 wire \bsr.update_data_i[2] ;
 wire \bsr.update_data_i[3] ;
 wire \bsr.update_data_i[4] ;
 wire \bsr.update_data_i[5] ;
 wire \bsr.update_data_i[6] ;
 wire \bsr.update_data_i[7] ;
 wire \bsr.update_data_i[8] ;
 wire \bsr.update_data_i[9] ;
 wire \bsr.values[10] ;
 wire \bsr.values[11] ;
 wire \bsr.values[12] ;
 wire \bsr.values[13] ;
 wire \bsr.values[14] ;
 wire \bsr.values[15] ;
 wire \bsr.values[16] ;
 wire \bsr.values[17] ;
 wire \bsr.values[18] ;
 wire \bsr.values[19] ;
 wire \bsr.values[20] ;
 wire \bsr.values[21] ;
 wire \bsr.values[22] ;
 wire \bsr.values[23] ;
 wire \bsr.values[24] ;
 wire \bsr.values[25] ;
 wire \bsr.values[2] ;
 wire \bsr.values[3] ;
 wire \bsr.values[4] ;
 wire \bsr.values[5] ;
 wire \bsr.values[6] ;
 wire \inner.counter[0] ;
 wire \inner.counter[1] ;
 wire \inner.counter[2] ;
 wire \inner.counter[3] ;
 wire \ir[0] ;
 wire \ir[1] ;
 wire \ir[2] ;
 wire \ir[3] ;
 wire \shift_q[26] ;
 wire \shift_q[27] ;
 wire \shift_q[28] ;
 wire \shift_q[29] ;
 wire \shift_q[30] ;
 wire \shift_q[31] ;
 wire \tap_sm.bypass_shift_q ;
 wire \tap_sm.ir_shift_q[0] ;
 wire \tap_sm.ir_shift_q[1] ;
 wire \tap_sm.ir_shift_q[2] ;
 wire \tap_sm.ir_shift_q[3] ;
 wire \tap_sm.state_d[0] ;
 wire \tap_sm.state_d[1] ;
 wire \tap_sm.state_d[2] ;
 wire \tap_sm.state_d[3] ;
 wire \tap_sm.state_q[0] ;
 wire \tap_sm.state_q[1] ;
 wire \tap_sm.state_q[2] ;
 wire \tap_sm.state_q[3] ;
 wire \tap_sm.tdo_o ;
 wire \tap_sm.tdo_oe_o ;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;

 sg13g2_inv_1 _461_ (.Y(_084_),
    .A(net184));
 sg13g2_inv_1 _462_ (.Y(_150_),
    .A(\bsr.values[24] ));
 sg13g2_inv_1 _463_ (.Y(_151_),
    .A(\bsr.update_data_i[24] ));
 sg13g2_inv_1 _464_ (.Y(_152_),
    .A(\bsr.values[23] ));
 sg13g2_inv_1 _465_ (.Y(_153_),
    .A(\bsr.update_data_i[23] ));
 sg13g2_inv_1 _466_ (.Y(_154_),
    .A(\bsr.values[22] ));
 sg13g2_inv_1 _467_ (.Y(_155_),
    .A(\bsr.update_data_i[22] ));
 sg13g2_inv_1 _468_ (.Y(_156_),
    .A(\bsr.update_data_i[21] ));
 sg13g2_inv_1 _469_ (.Y(_157_),
    .A(\bsr.values[20] ));
 sg13g2_inv_1 _470_ (.Y(_158_),
    .A(\bsr.update_data_i[20] ));
 sg13g2_inv_1 _471_ (.Y(_159_),
    .A(\bsr.update_data_i[18] ));
 sg13g2_inv_1 _472_ (.Y(_160_),
    .A(\bsr.update_data_i[13] ));
 sg13g2_inv_1 _473_ (.Y(_161_),
    .A(\bsr.update_data_i[11] ));
 sg13g2_inv_1 _474_ (.Y(_162_),
    .A(\bsr.update_data_i[10] ));
 sg13g2_inv_1 _475_ (.Y(_163_),
    .A(\bsr.update_data_i[6] ));
 sg13g2_inv_1 _476_ (.Y(_164_),
    .A(\bsr.values[5] ));
 sg13g2_inv_1 _477_ (.Y(_165_),
    .A(\bsr.update_data_i[5] ));
 sg13g2_inv_1 _478_ (.Y(_166_),
    .A(\bsr.update_data_i[4] ));
 sg13g2_inv_1 _479_ (.Y(_167_),
    .A(\bsr.update_data_i[8] ));
 sg13g2_inv_1 _480_ (.Y(_168_),
    .A(net1));
 sg13g2_inv_1 _481_ (.Y(_169_),
    .A(net2));
 sg13g2_inv_1 _482_ (.Y(_170_),
    .A(net3));
 sg13g2_inv_1 _483_ (.Y(_171_),
    .A(net6));
 sg13g2_inv_1 _484_ (.Y(_172_),
    .A(net8));
 sg13g2_inv_1 _485_ (.Y(_173_),
    .A(_004_));
 sg13g2_inv_1 _486_ (.Y(_174_),
    .A(\tap_sm.bypass_shift_q ));
 sg13g2_inv_1 _487_ (.Y(_045_),
    .A(net200));
 sg13g2_nor2_2 _488_ (.A(\tap_sm.state_q[3] ),
    .B(\tap_sm.state_q[2] ),
    .Y(_175_));
 sg13g2_inv_1 _489_ (.Y(_176_),
    .A(_175_));
 sg13g2_nor2b_1 _490_ (.A(net180),
    .B_N(net181),
    .Y(_177_));
 sg13g2_nor2_2 _491_ (.A(net180),
    .B(net181),
    .Y(_178_));
 sg13g2_nor2b_2 _492_ (.A(\tap_sm.state_q[2] ),
    .B_N(\tap_sm.state_q[3] ),
    .Y(_179_));
 sg13g2_and2_1 _493_ (.A(_178_),
    .B(_179_),
    .X(_180_));
 sg13g2_nand2_2 _494_ (.Y(_181_),
    .A(\tap_sm.state_q[3] ),
    .B(\tap_sm.state_q[2] ));
 sg13g2_o21ai_1 _495_ (.B1(_181_),
    .Y(_182_),
    .A1(net180),
    .A2(_176_));
 sg13g2_a21oi_1 _496_ (.A1(\tap_sm.state_q[0] ),
    .A2(_182_),
    .Y(_183_),
    .B1(_180_));
 sg13g2_or2_1 _497_ (.X(_184_),
    .B(_181_),
    .A(net180));
 sg13g2_nand2_1 _498_ (.Y(_185_),
    .A(_183_),
    .B(_184_));
 sg13g2_nand2_1 _499_ (.Y(_186_),
    .A(net191),
    .B(_185_));
 sg13g2_nor2b_2 _500_ (.A(net181),
    .B_N(net180),
    .Y(_187_));
 sg13g2_nor2b_2 _501_ (.A(\tap_sm.state_q[3] ),
    .B_N(\tap_sm.state_q[2] ),
    .Y(_188_));
 sg13g2_a22oi_1 _502_ (.Y(_189_),
    .B1(_188_),
    .B2(_177_),
    .A2(_187_),
    .A1(_175_));
 sg13g2_nor2_1 _503_ (.A(net191),
    .B(_189_),
    .Y(_190_));
 sg13g2_and2_1 _504_ (.A(net180),
    .B(_179_),
    .X(_191_));
 sg13g2_nand2_1 _505_ (.Y(_192_),
    .A(\tap_sm.state_q[1] ),
    .B(_179_));
 sg13g2_nor2_1 _506_ (.A(net191),
    .B(_192_),
    .Y(_193_));
 sg13g2_and2_1 _507_ (.A(_187_),
    .B(_188_),
    .X(_194_));
 sg13g2_a21oi_1 _508_ (.A1(net13),
    .A2(_194_),
    .Y(_195_),
    .B1(_193_));
 sg13g2_nand3b_1 _509_ (.B(_177_),
    .C(_179_),
    .Y(_196_),
    .A_N(net191));
 sg13g2_a21oi_1 _510_ (.A1(\tap_sm.state_q[2] ),
    .A2(_187_),
    .Y(_197_),
    .B1(_190_));
 sg13g2_nand4_1 _511_ (.B(_195_),
    .C(_196_),
    .A(_186_),
    .Y(\tap_sm.state_d[1] ),
    .D(_197_));
 sg13g2_and2_1 _512_ (.A(_175_),
    .B(_178_),
    .X(_198_));
 sg13g2_nor2b_1 _513_ (.A(_198_),
    .B_N(_183_),
    .Y(_199_));
 sg13g2_nand2_2 _514_ (.Y(_200_),
    .A(\tap_sm.state_q[1] ),
    .B(\tap_sm.state_q[0] ));
 sg13g2_nor2_2 _515_ (.A(_176_),
    .B(_200_),
    .Y(_201_));
 sg13g2_nand3_1 _516_ (.B(net181),
    .C(_175_),
    .A(net180),
    .Y(_202_));
 sg13g2_and2_1 _517_ (.A(_178_),
    .B(_188_),
    .X(_203_));
 sg13g2_nand2_2 _518_ (.Y(_204_),
    .A(_178_),
    .B(_188_));
 sg13g2_nor2_1 _519_ (.A(_201_),
    .B(_203_),
    .Y(_205_));
 sg13g2_nand2_1 _520_ (.Y(_206_),
    .A(_202_),
    .B(_204_));
 sg13g2_nor2_1 _521_ (.A(net181),
    .B(_181_),
    .Y(_207_));
 sg13g2_a221oi_1 _522_ (.B2(net191),
    .C1(_207_),
    .B1(net175),
    .A1(_175_),
    .Y(_208_),
    .A2(_187_));
 sg13g2_and2_1 _523_ (.A(_195_),
    .B(_208_),
    .X(_209_));
 sg13g2_o21ai_1 _524_ (.B1(_209_),
    .Y(\tap_sm.state_d[0] ),
    .A1(net13),
    .A2(_199_));
 sg13g2_a22oi_1 _525_ (.Y(_210_),
    .B1(_188_),
    .B2(net181),
    .A2(_187_),
    .A1(_175_));
 sg13g2_nand2b_1 _526_ (.Y(_211_),
    .B(net191),
    .A_N(_210_));
 sg13g2_a21oi_1 _527_ (.A1(net180),
    .A2(_207_),
    .Y(_212_),
    .B1(_191_));
 sg13g2_nand4_1 _528_ (.B(_196_),
    .C(_211_),
    .A(_184_),
    .Y(\tap_sm.state_d[3] ),
    .D(_212_));
 sg13g2_nand2b_1 _529_ (.Y(_213_),
    .B(net191),
    .A_N(_212_));
 sg13g2_nand3b_1 _530_ (.B(_188_),
    .C(net181),
    .Y(_214_),
    .A_N(net191));
 sg13g2_nand2_1 _531_ (.Y(_215_),
    .A(_184_),
    .B(net165));
 sg13g2_nor2_1 _532_ (.A(_194_),
    .B(_215_),
    .Y(_216_));
 sg13g2_nand3_1 _533_ (.B(_214_),
    .C(_216_),
    .A(_213_),
    .Y(\tap_sm.state_d[2] ));
 sg13g2_or4_1 _534_ (.A(\tap_sm.state_d[1] ),
    .B(\tap_sm.state_d[0] ),
    .C(\tap_sm.state_d[3] ),
    .D(\tap_sm.state_d[2] ),
    .X(_087_));
 sg13g2_nor2_1 _535_ (.A(\ir[3] ),
    .B(\ir[2] ),
    .Y(_217_));
 sg13g2_or2_1 _536_ (.X(_218_),
    .B(\ir[2] ),
    .A(\ir[3] ));
 sg13g2_nor2_2 _537_ (.A(\ir[1] ),
    .B(\ir[0] ),
    .Y(_219_));
 sg13g2_inv_1 _538_ (.Y(_220_),
    .A(_219_));
 sg13g2_nand3_1 _539_ (.B(net178),
    .C(_220_),
    .A(_180_),
    .Y(_221_));
 sg13g2_mux2_1 _540_ (.A0(\bsr.update_data_i[25] ),
    .A1(\bsr.values[25] ),
    .S(net169),
    .X(_149_));
 sg13g2_nor2_1 _541_ (.A(\bsr.update_data_i[24] ),
    .B(net168),
    .Y(_222_));
 sg13g2_a21oi_1 _542_ (.A1(_150_),
    .A2(net169),
    .Y(_148_),
    .B1(_222_));
 sg13g2_nor2_1 _543_ (.A(\bsr.update_data_i[23] ),
    .B(net170),
    .Y(_223_));
 sg13g2_a21oi_1 _544_ (.A1(_152_),
    .A2(net171),
    .Y(_147_),
    .B1(_223_));
 sg13g2_nor2_1 _545_ (.A(\bsr.update_data_i[22] ),
    .B(net170),
    .Y(_224_));
 sg13g2_a21oi_1 _546_ (.A1(_154_),
    .A2(net170),
    .Y(_146_),
    .B1(_224_));
 sg13g2_nand2_1 _547_ (.Y(_225_),
    .A(\bsr.values[21] ),
    .B(net170));
 sg13g2_o21ai_1 _548_ (.B1(_225_),
    .Y(_145_),
    .A1(_156_),
    .A2(net170));
 sg13g2_nor2_1 _549_ (.A(\bsr.update_data_i[20] ),
    .B(net170),
    .Y(_226_));
 sg13g2_a21oi_1 _550_ (.A1(_157_),
    .A2(net171),
    .Y(_144_),
    .B1(_226_));
 sg13g2_mux2_1 _551_ (.A0(\bsr.update_data_i[19] ),
    .A1(\bsr.values[19] ),
    .S(net170),
    .X(_143_));
 sg13g2_nand2_1 _552_ (.Y(_227_),
    .A(\bsr.values[18] ),
    .B(net172));
 sg13g2_o21ai_1 _553_ (.B1(_227_),
    .Y(_142_),
    .A1(_159_),
    .A2(net172));
 sg13g2_mux2_1 _554_ (.A0(\bsr.update_data_i[17] ),
    .A1(\bsr.values[17] ),
    .S(net168),
    .X(_141_));
 sg13g2_mux2_1 _555_ (.A0(\bsr.update_data_i[16] ),
    .A1(\bsr.values[16] ),
    .S(net169),
    .X(_140_));
 sg13g2_mux2_1 _556_ (.A0(\bsr.update_data_i[15] ),
    .A1(\bsr.values[15] ),
    .S(net170),
    .X(_139_));
 sg13g2_mux2_1 _557_ (.A0(\bsr.update_data_i[14] ),
    .A1(\bsr.values[14] ),
    .S(net169),
    .X(_138_));
 sg13g2_nand2_1 _558_ (.Y(_228_),
    .A(\bsr.values[13] ),
    .B(net168));
 sg13g2_o21ai_1 _559_ (.B1(_228_),
    .Y(_137_),
    .A1(_160_),
    .A2(net168));
 sg13g2_mux2_1 _560_ (.A0(\bsr.update_data_i[12] ),
    .A1(\bsr.values[12] ),
    .S(net169),
    .X(_136_));
 sg13g2_nand2_1 _561_ (.Y(_229_),
    .A(\bsr.values[11] ),
    .B(net168));
 sg13g2_o21ai_1 _562_ (.B1(_229_),
    .Y(_135_),
    .A1(_161_),
    .A2(net168));
 sg13g2_nand2_1 _563_ (.Y(_230_),
    .A(\bsr.values[10] ),
    .B(net168));
 sg13g2_o21ai_1 _564_ (.B1(_230_),
    .Y(_134_),
    .A1(_162_),
    .A2(net168));
 sg13g2_nand2_1 _565_ (.Y(_231_),
    .A(\bsr.values[6] ),
    .B(net173));
 sg13g2_o21ai_1 _566_ (.B1(_231_),
    .Y(_133_),
    .A1(_163_),
    .A2(net173));
 sg13g2_nor2_1 _567_ (.A(\bsr.update_data_i[5] ),
    .B(net172),
    .Y(_232_));
 sg13g2_a21oi_1 _568_ (.A1(_164_),
    .A2(net172),
    .Y(_132_),
    .B1(_232_));
 sg13g2_nand2_1 _569_ (.Y(_233_),
    .A(\bsr.values[4] ),
    .B(net172));
 sg13g2_o21ai_1 _570_ (.B1(_233_),
    .Y(_131_),
    .A1(_166_),
    .A2(net172));
 sg13g2_mux2_1 _571_ (.A0(\bsr.update_data_i[3] ),
    .A1(\bsr.values[3] ),
    .S(net172),
    .X(_130_));
 sg13g2_mux2_1 _572_ (.A0(\bsr.update_data_i[2] ),
    .A1(\bsr.values[2] ),
    .S(net172),
    .X(_129_));
 sg13g2_nand2_1 _573_ (.Y(_234_),
    .A(\shift_q[31] ),
    .B(net162));
 sg13g2_nand2_2 _574_ (.Y(_235_),
    .A(net178),
    .B(_219_));
 sg13g2_nand2_1 _575_ (.Y(_236_),
    .A(net14),
    .B(_203_));
 sg13g2_o21ai_1 _576_ (.B1(_234_),
    .Y(_123_),
    .A1(_235_),
    .A2(_236_));
 sg13g2_nor2_2 _577_ (.A(_204_),
    .B(net176),
    .Y(_237_));
 sg13g2_nor3_2 _578_ (.A(_204_),
    .B(net176),
    .C(_220_),
    .Y(_238_));
 sg13g2_a22oi_1 _579_ (.Y(_239_),
    .B1(_238_),
    .B2(\shift_q[31] ),
    .A2(net162),
    .A1(\shift_q[30] ));
 sg13g2_inv_1 _580_ (.Y(_122_),
    .A(_239_));
 sg13g2_nor2_1 _581_ (.A(_202_),
    .B(_235_),
    .Y(_240_));
 sg13g2_a221oi_1 _582_ (.B2(\shift_q[30] ),
    .C1(_240_),
    .B1(_238_),
    .A1(\shift_q[29] ),
    .Y(_241_),
    .A2(net162));
 sg13g2_inv_1 _583_ (.Y(_121_),
    .A(_241_));
 sg13g2_a221oi_1 _584_ (.B2(\shift_q[29] ),
    .C1(_240_),
    .B1(_238_),
    .A1(\shift_q[28] ),
    .Y(_242_),
    .A2(net162));
 sg13g2_inv_1 _585_ (.Y(_120_),
    .A(_242_));
 sg13g2_a22oi_1 _586_ (.Y(_243_),
    .B1(_238_),
    .B2(\shift_q[28] ),
    .A2(net162),
    .A1(\shift_q[27] ));
 sg13g2_inv_1 _587_ (.Y(_119_),
    .A(_243_));
 sg13g2_a22oi_1 _588_ (.Y(_244_),
    .B1(_238_),
    .B2(\shift_q[27] ),
    .A2(net162),
    .A1(\shift_q[26] ));
 sg13g2_inv_1 _589_ (.Y(_118_),
    .A(_244_));
 sg13g2_nor3_1 _590_ (.A(net176),
    .B(_219_),
    .C(_236_),
    .Y(_245_));
 sg13g2_a221oi_1 _591_ (.B2(\shift_q[26] ),
    .C1(_245_),
    .B1(_238_),
    .A1(\bsr.update_data_i[25] ),
    .Y(_246_),
    .A2(net162));
 sg13g2_inv_1 _592_ (.Y(_117_),
    .A(_246_));
 sg13g2_nor2_1 _593_ (.A(_202_),
    .B(net176),
    .Y(_247_));
 sg13g2_nand2_1 _594_ (.Y(_248_),
    .A(_201_),
    .B(net178));
 sg13g2_and2_2 _595_ (.A(\ir[0] ),
    .B(net167),
    .X(_249_));
 sg13g2_and2_2 _596_ (.A(\ir[1] ),
    .B(\ir[0] ),
    .X(_250_));
 sg13g2_nand2_2 _597_ (.Y(_251_),
    .A(\ir[1] ),
    .B(\ir[0] ));
 sg13g2_nor2_2 _598_ (.A(net177),
    .B(_251_),
    .Y(_252_));
 sg13g2_nand2_2 _599_ (.Y(_253_),
    .A(net179),
    .B(_250_));
 sg13g2_a21oi_2 _600_ (.B1(_168_),
    .Y(_254_),
    .A2(_250_),
    .A1(net179));
 sg13g2_o21ai_1 _601_ (.B1(net1),
    .Y(_255_),
    .A1(net177),
    .A2(_251_));
 sg13g2_nor3_2 _602_ (.A(_002_),
    .B(net177),
    .C(_251_),
    .Y(_256_));
 sg13g2_nand3b_1 _603_ (.B(net179),
    .C(_250_),
    .Y(_257_),
    .A_N(_002_));
 sg13g2_nor2_1 _604_ (.A(_254_),
    .B(_256_),
    .Y(_258_));
 sg13g2_nand2_2 _605_ (.Y(_259_),
    .A(_255_),
    .B(_257_));
 sg13g2_nor3_1 _606_ (.A(_007_),
    .B(net177),
    .C(_251_),
    .Y(_260_));
 sg13g2_a221oi_1 _607_ (.B2(_257_),
    .C1(_260_),
    .B1(_255_),
    .A1(net5),
    .Y(_261_),
    .A2(_253_));
 sg13g2_a21oi_1 _608_ (.A1(_006_),
    .A2(_258_),
    .Y(_262_),
    .B1(_261_));
 sg13g2_a21o_2 _609_ (.A2(_258_),
    .A1(_006_),
    .B1(_261_),
    .X(_263_));
 sg13g2_a21oi_1 _610_ (.A1(net178),
    .A2(_250_),
    .Y(_264_),
    .B1(_170_));
 sg13g2_o21ai_1 _611_ (.B1(net3),
    .Y(_265_),
    .A1(net177),
    .A2(_251_));
 sg13g2_a21oi_1 _612_ (.A1(\bsr.values[4] ),
    .A2(_252_),
    .Y(_266_),
    .B1(_264_));
 sg13g2_nor3_1 _613_ (.A(\inner.counter[1] ),
    .B(_254_),
    .C(_256_),
    .Y(_267_));
 sg13g2_a21o_1 _614_ (.A2(_266_),
    .A1(_259_),
    .B1(_267_),
    .X(_268_));
 sg13g2_a21oi_1 _615_ (.A1(_259_),
    .A2(_266_),
    .Y(_269_),
    .B1(_267_));
 sg13g2_a21oi_1 _616_ (.A1(net178),
    .A2(_250_),
    .Y(_270_),
    .B1(_169_));
 sg13g2_a221oi_1 _617_ (.B2(_257_),
    .C1(_270_),
    .B1(_255_),
    .A1(\bsr.values[3] ),
    .Y(_271_),
    .A2(_252_));
 sg13g2_nor3_2 _618_ (.A(\inner.counter[0] ),
    .B(_254_),
    .C(_256_),
    .Y(_272_));
 sg13g2_nor2_2 _619_ (.A(_271_),
    .B(_272_),
    .Y(_273_));
 sg13g2_or2_1 _620_ (.X(_274_),
    .B(_272_),
    .A(_271_));
 sg13g2_nand3_1 _621_ (.B(_255_),
    .C(_257_),
    .A(_004_),
    .Y(_275_));
 sg13g2_o21ai_1 _622_ (.B1(net4),
    .Y(_276_),
    .A1(net176),
    .A2(_251_));
 sg13g2_o21ai_1 _623_ (.B1(_276_),
    .Y(_277_),
    .A1(_005_),
    .A2(_253_));
 sg13g2_mux2_2 _624_ (.A0(_173_),
    .A1(_277_),
    .S(_259_),
    .X(_278_));
 sg13g2_o21ai_1 _625_ (.B1(_275_),
    .Y(_279_),
    .A1(_258_),
    .A2(_277_));
 sg13g2_a21oi_1 _626_ (.A1(_269_),
    .A2(_273_),
    .Y(_280_),
    .B1(_279_));
 sg13g2_nor2_1 _627_ (.A(_262_),
    .B(_279_),
    .Y(_281_));
 sg13g2_and2_1 _628_ (.A(_263_),
    .B(_280_),
    .X(_282_));
 sg13g2_nand2_1 _629_ (.Y(_283_),
    .A(_268_),
    .B(_274_));
 sg13g2_a21oi_1 _630_ (.A1(_263_),
    .A2(_268_),
    .Y(_284_),
    .B1(_278_));
 sg13g2_a21o_1 _631_ (.A2(_283_),
    .A1(_262_),
    .B1(_284_),
    .X(_285_));
 sg13g2_o21ai_1 _632_ (.B1(_249_),
    .Y(_286_),
    .A1(_282_),
    .A2(_285_));
 sg13g2_nor2_1 _633_ (.A(_201_),
    .B(net176),
    .Y(_287_));
 sg13g2_a21oi_1 _634_ (.A1(\bsr.update_data_i[25] ),
    .A2(net160),
    .Y(_288_),
    .B1(net161));
 sg13g2_a22oi_1 _635_ (.Y(_116_),
    .B1(_286_),
    .B2(_288_),
    .A2(net161),
    .A1(_151_));
 sg13g2_nor2_1 _636_ (.A(_263_),
    .B(_278_),
    .Y(_289_));
 sg13g2_nand3b_1 _637_ (.B(net178),
    .C(_250_),
    .Y(_290_),
    .A_N(_003_));
 sg13g2_a22oi_1 _638_ (.Y(_291_),
    .B1(_265_),
    .B2(_290_),
    .A2(_257_),
    .A1(_255_));
 sg13g2_nor3_2 _639_ (.A(_001_),
    .B(_254_),
    .C(_256_),
    .Y(_292_));
 sg13g2_nor2_2 _640_ (.A(_291_),
    .B(_292_),
    .Y(_293_));
 sg13g2_nor4_2 _641_ (.A(_271_),
    .B(_272_),
    .C(_291_),
    .Y(_294_),
    .D(_292_));
 sg13g2_a21oi_1 _642_ (.A1(_278_),
    .A2(_294_),
    .Y(_295_),
    .B1(_263_));
 sg13g2_nand3_1 _643_ (.B(_274_),
    .C(_293_),
    .A(_263_),
    .Y(_296_));
 sg13g2_nand2b_1 _644_ (.Y(_297_),
    .B(_296_),
    .A_N(_295_));
 sg13g2_o21ai_1 _645_ (.B1(_249_),
    .Y(_298_),
    .A1(_282_),
    .A2(_297_));
 sg13g2_a21oi_1 _646_ (.A1(\bsr.update_data_i[24] ),
    .A2(net160),
    .Y(_299_),
    .B1(net164));
 sg13g2_a22oi_1 _647_ (.Y(_115_),
    .B1(_298_),
    .B2(_299_),
    .A2(net161),
    .A1(_153_));
 sg13g2_nand2_1 _648_ (.Y(_300_),
    .A(_268_),
    .B(_281_));
 sg13g2_o21ai_1 _649_ (.B1(_276_),
    .Y(_301_),
    .A1(_164_),
    .A2(_253_));
 sg13g2_mux2_1 _650_ (.A0(\inner.counter[2] ),
    .A1(_301_),
    .S(_259_),
    .X(_302_));
 sg13g2_nand2b_1 _651_ (.Y(_303_),
    .B(_294_),
    .A_N(_302_));
 sg13g2_nand2_1 _652_ (.Y(_304_),
    .A(_263_),
    .B(_273_));
 sg13g2_nand4_1 _653_ (.B(_300_),
    .C(_303_),
    .A(_249_),
    .Y(_305_),
    .D(_304_));
 sg13g2_a21oi_1 _654_ (.A1(\bsr.update_data_i[23] ),
    .A2(net160),
    .Y(_306_),
    .B1(net161));
 sg13g2_a22oi_1 _655_ (.Y(_114_),
    .B1(_305_),
    .B2(_306_),
    .A2(net163),
    .A1(_155_));
 sg13g2_nor3_1 _656_ (.A(_262_),
    .B(_278_),
    .C(_294_),
    .Y(_307_));
 sg13g2_nand2b_1 _657_ (.Y(_308_),
    .B(_274_),
    .A_N(_293_));
 sg13g2_a221oi_1 _658_ (.B2(_289_),
    .C1(_307_),
    .B1(_308_),
    .A1(_280_),
    .Y(_309_),
    .A2(_296_));
 sg13g2_nand2b_1 _659_ (.Y(_310_),
    .B(_249_),
    .A_N(_309_));
 sg13g2_a21oi_1 _660_ (.A1(\bsr.update_data_i[22] ),
    .A2(net160),
    .Y(_311_),
    .B1(net163));
 sg13g2_a22oi_1 _661_ (.Y(_113_),
    .B1(_310_),
    .B2(_311_),
    .A2(net163),
    .A1(_156_));
 sg13g2_a21oi_1 _662_ (.A1(_268_),
    .A2(_273_),
    .Y(_312_),
    .B1(_263_));
 sg13g2_nor3_1 _663_ (.A(_273_),
    .B(_278_),
    .C(_293_),
    .Y(_313_));
 sg13g2_nor2_1 _664_ (.A(_312_),
    .B(_313_),
    .Y(_314_));
 sg13g2_o21ai_1 _665_ (.B1(_249_),
    .Y(_315_),
    .A1(_289_),
    .A2(_314_));
 sg13g2_a21oi_1 _666_ (.A1(\bsr.update_data_i[21] ),
    .A2(net160),
    .Y(_316_),
    .B1(net163));
 sg13g2_a22oi_1 _667_ (.Y(_112_),
    .B1(_315_),
    .B2(_316_),
    .A2(net163),
    .A1(_158_));
 sg13g2_xnor2_1 _668_ (.Y(_317_),
    .A(_273_),
    .B(_293_));
 sg13g2_or2_1 _669_ (.X(_318_),
    .B(_302_),
    .A(_273_));
 sg13g2_a22oi_1 _670_ (.Y(_319_),
    .B1(_318_),
    .B2(_312_),
    .A2(_317_),
    .A1(_281_));
 sg13g2_a22oi_1 _671_ (.Y(_320_),
    .B1(_319_),
    .B2(_249_),
    .A2(net158),
    .A1(\bsr.update_data_i[20] ));
 sg13g2_nor2_1 _672_ (.A(\bsr.update_data_i[19] ),
    .B(net174),
    .Y(_321_));
 sg13g2_a21oi_1 _673_ (.A1(net174),
    .A2(_320_),
    .Y(_111_),
    .B1(_321_));
 sg13g2_nand3_1 _674_ (.B(_273_),
    .C(_279_),
    .A(_269_),
    .Y(_322_));
 sg13g2_a221oi_1 _675_ (.B2(_322_),
    .C1(_307_),
    .B1(_295_),
    .A1(_281_),
    .Y(_323_),
    .A2(_283_));
 sg13g2_nand2b_1 _676_ (.Y(_324_),
    .B(_249_),
    .A_N(_323_));
 sg13g2_a21oi_1 _677_ (.A1(\bsr.update_data_i[19] ),
    .A2(net158),
    .Y(_325_),
    .B1(net165));
 sg13g2_a22oi_1 _678_ (.Y(_110_),
    .B1(_324_),
    .B2(_325_),
    .A2(net165),
    .A1(_159_));
 sg13g2_nor2_2 _679_ (.A(net162),
    .B(_240_),
    .Y(_326_));
 sg13g2_o21ai_1 _680_ (.B1(net174),
    .Y(_327_),
    .A1(_202_),
    .A2(_235_));
 sg13g2_a21oi_1 _681_ (.A1(\bsr.update_data_i[18] ),
    .A2(net158),
    .Y(_328_),
    .B1(_327_));
 sg13g2_nor2_1 _682_ (.A(\bsr.update_data_i[17] ),
    .B(net175),
    .Y(_329_));
 sg13g2_nand2_1 _683_ (.Y(_330_),
    .A(\ir[1] ),
    .B(net178));
 sg13g2_nor3_2 _684_ (.A(\ir[0] ),
    .B(_202_),
    .C(_330_),
    .Y(_331_));
 sg13g2_nand2_1 _685_ (.Y(_332_),
    .A(net12),
    .B(_331_));
 sg13g2_o21ai_1 _686_ (.B1(_332_),
    .Y(_109_),
    .A1(_328_),
    .A2(_329_));
 sg13g2_a22oi_1 _687_ (.Y(_333_),
    .B1(_331_),
    .B2(net11),
    .A2(net158),
    .A1(\bsr.update_data_i[17] ));
 sg13g2_nor2_1 _688_ (.A(\bsr.update_data_i[16] ),
    .B(net174),
    .Y(_334_));
 sg13g2_a21oi_1 _689_ (.A1(net174),
    .A2(_333_),
    .Y(_108_),
    .B1(_334_));
 sg13g2_a21oi_1 _690_ (.A1(\bsr.update_data_i[16] ),
    .A2(net158),
    .Y(_335_),
    .B1(_327_));
 sg13g2_nor2_1 _691_ (.A(\bsr.update_data_i[15] ),
    .B(net174),
    .Y(_336_));
 sg13g2_nand2_1 _692_ (.Y(_337_),
    .A(net10),
    .B(_331_));
 sg13g2_o21ai_1 _693_ (.B1(_337_),
    .Y(_107_),
    .A1(_335_),
    .A2(_336_));
 sg13g2_a22oi_1 _694_ (.Y(_338_),
    .B1(_331_),
    .B2(net9),
    .A2(net158),
    .A1(\bsr.update_data_i[15] ));
 sg13g2_nor2_1 _695_ (.A(\bsr.update_data_i[14] ),
    .B(net174),
    .Y(_339_));
 sg13g2_a21oi_1 _696_ (.A1(net174),
    .A2(_338_),
    .Y(_106_),
    .B1(_339_));
 sg13g2_nand2_1 _697_ (.Y(_340_),
    .A(\bsr.update_data_i[14] ),
    .B(net160));
 sg13g2_a22oi_1 _698_ (.Y(_105_),
    .B1(_326_),
    .B2(_340_),
    .A2(net161),
    .A1(_160_));
 sg13g2_a22oi_1 _699_ (.Y(_341_),
    .B1(_237_),
    .B2(\bsr.update_data_i[13] ),
    .A2(net161),
    .A1(\bsr.update_data_i[12] ));
 sg13g2_inv_1 _700_ (.Y(_104_),
    .A(_341_));
 sg13g2_nand2_1 _701_ (.Y(_342_),
    .A(\bsr.update_data_i[12] ),
    .B(net160));
 sg13g2_a22oi_1 _702_ (.Y(_103_),
    .B1(_326_),
    .B2(_342_),
    .A2(net161),
    .A1(_161_));
 sg13g2_nand2_1 _703_ (.Y(_343_),
    .A(\bsr.update_data_i[11] ),
    .B(net160));
 sg13g2_a22oi_1 _704_ (.Y(_102_),
    .B1(_326_),
    .B2(_343_),
    .A2(net161),
    .A1(_162_));
 sg13g2_o21ai_1 _705_ (.B1(_235_),
    .Y(_344_),
    .A1(_172_),
    .A2(_252_));
 sg13g2_a22oi_1 _706_ (.Y(_345_),
    .B1(_344_),
    .B2(net167),
    .A2(net159),
    .A1(\bsr.update_data_i[10] ));
 sg13g2_nor2_1 _707_ (.A(\bsr.update_data_i[9] ),
    .B(net175),
    .Y(_346_));
 sg13g2_a21oi_1 _708_ (.A1(net175),
    .A2(_345_),
    .Y(_101_),
    .B1(_346_));
 sg13g2_nand4_1 _709_ (.B(_220_),
    .C(net167),
    .A(net7),
    .Y(_347_),
    .D(_253_));
 sg13g2_a21oi_1 _710_ (.A1(\bsr.update_data_i[9] ),
    .A2(net159),
    .Y(_348_),
    .B1(net166));
 sg13g2_a22oi_1 _711_ (.Y(_100_),
    .B1(_347_),
    .B2(_348_),
    .A2(net166),
    .A1(_167_));
 sg13g2_o21ai_1 _712_ (.B1(_235_),
    .Y(_349_),
    .A1(_171_),
    .A2(_252_));
 sg13g2_nand3_1 _713_ (.B(_202_),
    .C(_204_),
    .A(\bsr.update_data_i[7] ),
    .Y(_350_));
 sg13g2_a22oi_1 _714_ (.Y(_351_),
    .B1(_349_),
    .B2(net167),
    .A2(net159),
    .A1(\bsr.update_data_i[8] ));
 sg13g2_o21ai_1 _715_ (.B1(_350_),
    .Y(_099_),
    .A1(net166),
    .A2(_351_));
 sg13g2_nand3_1 _716_ (.B(net167),
    .C(_253_),
    .A(net5),
    .Y(_352_));
 sg13g2_a21oi_1 _717_ (.A1(\bsr.update_data_i[7] ),
    .A2(net159),
    .Y(_353_),
    .B1(_327_));
 sg13g2_a22oi_1 _718_ (.Y(_098_),
    .B1(_352_),
    .B2(_353_),
    .A2(net166),
    .A1(_163_));
 sg13g2_nand3_1 _719_ (.B(net167),
    .C(_253_),
    .A(net4),
    .Y(_354_));
 sg13g2_a21oi_1 _720_ (.A1(\bsr.update_data_i[6] ),
    .A2(net159),
    .Y(_355_),
    .B1(_327_));
 sg13g2_a22oi_1 _721_ (.Y(_097_),
    .B1(_354_),
    .B2(_355_),
    .A2(net165),
    .A1(_165_));
 sg13g2_a22oi_1 _722_ (.Y(_356_),
    .B1(net159),
    .B2(\bsr.update_data_i[5] ),
    .A2(_264_),
    .A1(net167));
 sg13g2_a22oi_1 _723_ (.Y(_096_),
    .B1(_326_),
    .B2(_356_),
    .A2(net166),
    .A1(_166_));
 sg13g2_o21ai_1 _724_ (.B1(_235_),
    .Y(_357_),
    .A1(_169_),
    .A2(_252_));
 sg13g2_nand2_1 _725_ (.Y(_358_),
    .A(\bsr.update_data_i[3] ),
    .B(net165));
 sg13g2_a22oi_1 _726_ (.Y(_359_),
    .B1(_357_),
    .B2(_247_),
    .A2(net158),
    .A1(\bsr.update_data_i[4] ));
 sg13g2_o21ai_1 _727_ (.B1(_358_),
    .Y(_095_),
    .A1(net165),
    .A2(_359_));
 sg13g2_nor2_1 _728_ (.A(\bsr.update_data_i[2] ),
    .B(net175),
    .Y(_360_));
 sg13g2_nand2_1 _729_ (.Y(_361_),
    .A(_235_),
    .B(_255_));
 sg13g2_a22oi_1 _730_ (.Y(_362_),
    .B1(_361_),
    .B2(net167),
    .A2(net158),
    .A1(\bsr.update_data_i[3] ));
 sg13g2_a21oi_1 _731_ (.A1(net175),
    .A2(_362_),
    .Y(_094_),
    .B1(_360_));
 sg13g2_nand2_1 _732_ (.Y(_363_),
    .A(_203_),
    .B(net176));
 sg13g2_nor2_1 _733_ (.A(net178),
    .B(_236_),
    .Y(_364_));
 sg13g2_a221oi_1 _734_ (.B2(\bsr.update_data_i[2] ),
    .C1(_364_),
    .B1(_237_),
    .A1(\bsr.update_data_i[1] ),
    .Y(_365_),
    .A2(net165));
 sg13g2_o21ai_1 _735_ (.B1(_365_),
    .Y(_093_),
    .A1(_219_),
    .A2(_248_));
 sg13g2_a22oi_1 _736_ (.Y(_366_),
    .B1(net165),
    .B2(\bsr.update_data_i[0] ),
    .A2(_203_),
    .A1(\bsr.update_data_i[1] ));
 sg13g2_nand2_1 _737_ (.Y(_092_),
    .A(_248_),
    .B(_366_));
 sg13g2_and2_2 _738_ (.A(\tap_sm.state_q[0] ),
    .B(_191_),
    .X(_367_));
 sg13g2_or2_1 _739_ (.X(\tap_sm.tdo_oe_o ),
    .B(_367_),
    .A(_203_));
 sg13g2_a22oi_1 _740_ (.Y(_368_),
    .B1(_367_),
    .B2(\tap_sm.ir_shift_q[0] ),
    .A2(_237_),
    .A1(\bsr.update_data_i[0] ));
 sg13g2_o21ai_1 _741_ (.B1(_368_),
    .Y(_000_),
    .A1(_174_),
    .A2(_363_));
 sg13g2_nor2_1 _742_ (.A(\ir[3] ),
    .B(_220_),
    .Y(_369_));
 sg13g2_a22oi_1 _743_ (.Y(_370_),
    .B1(_369_),
    .B2(\ir[2] ),
    .A2(net179),
    .A1(\ir[1] ));
 sg13g2_nor2b_2 _744_ (.A(net155),
    .B_N(\bsr.values[10] ),
    .Y(uio_oe[0]));
 sg13g2_nor2b_1 _745_ (.A(net155),
    .B_N(\bsr.values[11] ),
    .Y(uio_oe[1]));
 sg13g2_nor2b_2 _746_ (.A(net155),
    .B_N(\bsr.values[12] ),
    .Y(uio_oe[2]));
 sg13g2_nor2b_2 _747_ (.A(net155),
    .B_N(\bsr.values[13] ),
    .Y(uio_oe[3]));
 sg13g2_nor2b_1 _748_ (.A(_370_),
    .B_N(\bsr.values[14] ),
    .Y(uio_out[0]));
 sg13g2_nor2b_1 _749_ (.A(net155),
    .B_N(\bsr.values[15] ),
    .Y(uio_out[1]));
 sg13g2_nor2b_1 _750_ (.A(net155),
    .B_N(\bsr.values[16] ),
    .Y(uio_out[2]));
 sg13g2_nor2b_1 _751_ (.A(net155),
    .B_N(\bsr.values[17] ),
    .Y(uio_out[3]));
 sg13g2_nor2_1 _752_ (.A(\bsr.values[18] ),
    .B(net156),
    .Y(_371_));
 sg13g2_a21oi_2 _753_ (.B1(_371_),
    .Y(uo_out[0]),
    .A2(net156),
    .A1(_323_));
 sg13g2_mux2_1 _754_ (.A0(\bsr.values[19] ),
    .A1(_319_),
    .S(net157),
    .X(uo_out[1]));
 sg13g2_o21ai_1 _755_ (.B1(net156),
    .Y(_372_),
    .A1(_289_),
    .A2(_314_));
 sg13g2_o21ai_1 _756_ (.B1(_372_),
    .Y(uo_out[2]),
    .A1(_157_),
    .A2(net156));
 sg13g2_nor2_1 _757_ (.A(\bsr.values[21] ),
    .B(net157),
    .Y(_373_));
 sg13g2_a21oi_1 _758_ (.A1(_309_),
    .A2(net156),
    .Y(uo_out[3]),
    .B1(_373_));
 sg13g2_nand4_1 _759_ (.B(_303_),
    .C(_304_),
    .A(_300_),
    .Y(_374_),
    .D(net156));
 sg13g2_o21ai_1 _760_ (.B1(_374_),
    .Y(uo_out[4]),
    .A1(_154_),
    .A2(net157));
 sg13g2_o21ai_1 _761_ (.B1(net156),
    .Y(_375_),
    .A1(_282_),
    .A2(_297_));
 sg13g2_o21ai_1 _762_ (.B1(_375_),
    .Y(uo_out[5]),
    .A1(_152_),
    .A2(net157));
 sg13g2_o21ai_1 _763_ (.B1(net156),
    .Y(_376_),
    .A1(_282_),
    .A2(_285_));
 sg13g2_o21ai_1 _764_ (.B1(_376_),
    .Y(uo_out[6]),
    .A1(_150_),
    .A2(net157));
 sg13g2_nor2b_2 _765_ (.A(net155),
    .B_N(\bsr.values[25] ),
    .Y(uo_out[7]));
 sg13g2_nand2_1 _766_ (.Y(_377_),
    .A(\inner.counter[1] ),
    .B(\inner.counter[0] ));
 sg13g2_xor2_1 _767_ (.B(\inner.counter[0] ),
    .A(net26),
    .X(_008_));
 sg13g2_xnor2_1 _768_ (.Y(_009_),
    .A(net24),
    .B(_377_));
 sg13g2_nor2_1 _769_ (.A(_004_),
    .B(_377_),
    .Y(_378_));
 sg13g2_xor2_1 _770_ (.B(_378_),
    .A(net22),
    .X(_010_));
 sg13g2_nor2_2 _771_ (.A(_181_),
    .B(_200_),
    .Y(_379_));
 sg13g2_or2_1 _772_ (.X(_380_),
    .B(_200_),
    .A(_181_));
 sg13g2_nor2_1 _773_ (.A(_198_),
    .B(_379_),
    .Y(_381_));
 sg13g2_a22oi_1 _774_ (.Y(_382_),
    .B1(_381_),
    .B2(\ir[0] ),
    .A2(_379_),
    .A1(\tap_sm.ir_shift_q[0] ));
 sg13g2_inv_1 _775_ (.Y(_088_),
    .A(_382_));
 sg13g2_nand2_1 _776_ (.Y(_383_),
    .A(\ir[1] ),
    .B(_381_));
 sg13g2_nor2_1 _777_ (.A(net181),
    .B(_192_),
    .Y(_384_));
 sg13g2_nor2_1 _778_ (.A(\tap_sm.ir_shift_q[1] ),
    .B(_384_),
    .Y(_385_));
 sg13g2_o21ai_1 _779_ (.B1(_383_),
    .Y(_089_),
    .A1(_380_),
    .A2(_385_));
 sg13g2_a22oi_1 _780_ (.Y(_386_),
    .B1(_381_),
    .B2(\ir[2] ),
    .A2(_379_),
    .A1(\tap_sm.ir_shift_q[2] ));
 sg13g2_inv_1 _781_ (.Y(_090_),
    .A(_386_));
 sg13g2_nor2_1 _782_ (.A(\tap_sm.ir_shift_q[3] ),
    .B(_380_),
    .Y(_387_));
 sg13g2_nor2_1 _783_ (.A(\ir[3] ),
    .B(_379_),
    .Y(_388_));
 sg13g2_nor3_1 _784_ (.A(_198_),
    .B(_387_),
    .C(_388_),
    .Y(_091_));
 sg13g2_a21oi_1 _785_ (.A1(\tap_sm.bypass_shift_q ),
    .A2(_363_),
    .Y(_389_),
    .B1(_364_));
 sg13g2_a221oi_1 _786_ (.B2(net176),
    .C1(_389_),
    .B1(_201_),
    .A1(_175_),
    .Y(_124_),
    .A2(_178_));
 sg13g2_nor2_2 _787_ (.A(_191_),
    .B(_198_),
    .Y(_390_));
 sg13g2_nand2_1 _788_ (.Y(_391_),
    .A(\tap_sm.ir_shift_q[0] ),
    .B(_390_));
 sg13g2_o21ai_1 _789_ (.B1(_391_),
    .Y(_125_),
    .A1(_192_),
    .A2(_385_));
 sg13g2_a22oi_1 _790_ (.Y(_392_),
    .B1(_390_),
    .B2(\tap_sm.ir_shift_q[1] ),
    .A2(_367_),
    .A1(\tap_sm.ir_shift_q[2] ));
 sg13g2_inv_1 _791_ (.Y(_126_),
    .A(_392_));
 sg13g2_nand2_1 _792_ (.Y(_393_),
    .A(\tap_sm.ir_shift_q[3] ),
    .B(_367_));
 sg13g2_a22oi_1 _793_ (.Y(_394_),
    .B1(_390_),
    .B2(\tap_sm.ir_shift_q[2] ),
    .A2(_384_),
    .A1(\ir[2] ));
 sg13g2_nand2_1 _794_ (.Y(_127_),
    .A(_393_),
    .B(_394_));
 sg13g2_nand2_1 _795_ (.Y(_395_),
    .A(net14),
    .B(_367_));
 sg13g2_a22oi_1 _796_ (.Y(_396_),
    .B1(_390_),
    .B2(\tap_sm.ir_shift_q[3] ),
    .A2(_384_),
    .A1(\ir[3] ));
 sg13g2_nand2_1 _797_ (.Y(_128_),
    .A(_395_),
    .B(_396_));
 sg13g2_inv_1 _798_ (.Y(_082_),
    .A(net183));
 sg13g2_inv_1 _799_ (.Y(_080_),
    .A(net186));
 sg13g2_inv_1 _800_ (.Y(_078_),
    .A(net186));
 sg13g2_inv_1 _801_ (.Y(_076_),
    .A(net185));
 sg13g2_inv_1 _802_ (.Y(_074_),
    .A(net186));
 sg13g2_inv_1 _803_ (.Y(_072_),
    .A(net185));
 sg13g2_inv_1 _804_ (.Y(_070_),
    .A(net189));
 sg13g2_inv_1 _805_ (.Y(_068_),
    .A(net182));
 sg13g2_inv_1 _806_ (.Y(_066_),
    .A(net183));
 sg13g2_inv_1 _807_ (.Y(_064_),
    .A(net186));
 sg13g2_inv_1 _808_ (.Y(_062_),
    .A(net183));
 sg13g2_inv_1 _809_ (.Y(_060_),
    .A(net182));
 sg13g2_inv_1 _810_ (.Y(_058_),
    .A(net182));
 sg13g2_inv_1 _811_ (.Y(_056_),
    .A(net182));
 sg13g2_inv_1 _812_ (.Y(_054_),
    .A(net182));
 sg13g2_inv_1 _813_ (.Y(_052_),
    .A(net188));
 sg13g2_inv_1 _814_ (.Y(_050_),
    .A(net188));
 sg13g2_inv_1 _815_ (.Y(_048_),
    .A(net188));
 sg13g2_inv_1 _816_ (.Y(_046_),
    .A(net187));
 sg13g2_inv_1 _817_ (.Y(_044_),
    .A(net187));
 sg13g2_inv_1 _818_ (.Y(_012_),
    .A(net189));
 sg13g2_inv_1 _819_ (.Y(_013_),
    .A(net189));
 sg13g2_inv_1 _820_ (.Y(_014_),
    .A(net187));
 sg13g2_inv_1 _821_ (.Y(_015_),
    .A(net187));
 sg13g2_inv_1 _822_ (.Y(_016_),
    .A(net187));
 sg13g2_inv_1 _823_ (.Y(_017_),
    .A(net187));
 sg13g2_inv_1 _824_ (.Y(_018_),
    .A(net188));
 sg13g2_inv_1 _825_ (.Y(_019_),
    .A(net187));
 sg13g2_inv_1 _826_ (.Y(_020_),
    .A(net187));
 sg13g2_inv_1 _827_ (.Y(_021_),
    .A(net189));
 sg13g2_inv_1 _828_ (.Y(_022_),
    .A(net182));
 sg13g2_inv_1 _829_ (.Y(_023_),
    .A(net182));
 sg13g2_inv_1 _830_ (.Y(_024_),
    .A(net184));
 sg13g2_inv_1 _831_ (.Y(_025_),
    .A(net184));
 sg13g2_inv_1 _832_ (.Y(_026_),
    .A(net186));
 sg13g2_inv_1 _833_ (.Y(_027_),
    .A(net189));
 sg13g2_inv_1 _834_ (.Y(_028_),
    .A(net189));
 sg13g2_inv_1 _835_ (.Y(_029_),
    .A(net189));
 sg13g2_inv_1 _836_ (.Y(_030_),
    .A(net189));
 sg13g2_inv_1 _837_ (.Y(_031_),
    .A(net185));
 sg13g2_inv_1 _838_ (.Y(_032_),
    .A(net186));
 sg13g2_inv_1 _839_ (.Y(_033_),
    .A(net186));
 sg13g2_inv_1 _840_ (.Y(_034_),
    .A(net186));
 sg13g2_inv_1 _841_ (.Y(_035_),
    .A(net183));
 sg13g2_inv_1 _842_ (.Y(_036_),
    .A(net182));
 sg13g2_inv_1 _843_ (.Y(_037_),
    .A(net184));
 sg13g2_inv_1 _844_ (.Y(_038_),
    .A(net184));
 sg13g2_inv_1 _845_ (.Y(_039_),
    .A(net185));
 sg13g2_inv_1 _846_ (.Y(_040_),
    .A(net185));
 sg13g2_inv_1 _847_ (.Y(_041_),
    .A(net185));
 sg13g2_inv_1 _848_ (.Y(_042_),
    .A(net185));
 sg13g2_inv_1 _849_ (.Y(_043_),
    .A(net185));
 sg13g2_inv_1 _850_ (.Y(_047_),
    .A(net202));
 sg13g2_inv_1 _851_ (.Y(_049_),
    .A(net201));
 sg13g2_inv_1 _852_ (.Y(_051_),
    .A(net201));
 sg13g2_inv_1 _853_ (.Y(_053_),
    .A(net201));
 sg13g2_inv_1 _854_ (.Y(_055_),
    .A(net192));
 sg13g2_inv_1 _855_ (.Y(_057_),
    .A(net192));
 sg13g2_inv_1 _856_ (.Y(_059_),
    .A(net192));
 sg13g2_inv_1 _857_ (.Y(_061_),
    .A(net192));
 sg13g2_inv_1 _858_ (.Y(_063_),
    .A(net193));
 sg13g2_inv_1 _859_ (.Y(_065_),
    .A(net195));
 sg13g2_inv_1 _860_ (.Y(_067_),
    .A(net193));
 sg13g2_inv_1 _861_ (.Y(_069_),
    .A(net193));
 sg13g2_inv_1 _862_ (.Y(_071_),
    .A(net198));
 sg13g2_inv_1 _863_ (.Y(_073_),
    .A(net196));
 sg13g2_inv_1 _864_ (.Y(_075_),
    .A(net196));
 sg13g2_inv_1 _865_ (.Y(_077_),
    .A(net195));
 sg13g2_inv_1 _866_ (.Y(_079_),
    .A(net195));
 sg13g2_inv_1 _867_ (.Y(_081_),
    .A(net195));
 sg13g2_inv_1 _868_ (.Y(_083_),
    .A(net193));
 sg13g2_inv_1 _869_ (.Y(_085_),
    .A(net194));
 sg13g2_inv_1 _870_ (.Y(_086_),
    .A(net197));
 sg13g2_dfrbp_1 _871_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net206),
    .D(net21),
    .Q_N(_397_),
    .Q(\inner.counter[0] ));
 sg13g2_dfrbp_1 _872_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net206),
    .D(net27),
    .Q_N(_001_),
    .Q(\inner.counter[1] ));
 sg13g2_dfrbp_1 _873_ (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net206),
    .D(net25),
    .Q_N(_004_),
    .Q(\inner.counter[2] ));
 sg13g2_dfrbp_1 _874_ (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net206),
    .D(net23),
    .Q_N(_006_),
    .Q(\inner.counter[3] ));
 sg13g2_dfrbp_1 _875_ (.CLK(net199),
    .RESET_B(net205),
    .D(_088_),
    .Q_N(_457_),
    .Q(\ir[0] ));
 sg13g2_dfrbp_1 _876_ (.CLK(net199),
    .RESET_B(net205),
    .D(_089_),
    .Q_N(_456_),
    .Q(\ir[1] ));
 sg13g2_dfrbp_1 _877_ (.CLK(net200),
    .RESET_B(net205),
    .D(_090_),
    .Q_N(_455_),
    .Q(\ir[2] ));
 sg13g2_dfrbp_1 _878_ (.CLK(net199),
    .RESET_B(net205),
    .D(_091_),
    .Q_N(_454_),
    .Q(\ir[3] ));
 sg13g2_dfrbp_1 _879_ (.CLK(net197),
    .RESET_B(_012_),
    .D(_092_),
    .Q_N(_453_),
    .Q(\bsr.update_data_i[0] ));
 sg13g2_dfrbp_1 _880_ (.CLK(net197),
    .RESET_B(_013_),
    .D(_093_),
    .Q_N(_452_),
    .Q(\bsr.update_data_i[1] ));
 sg13g2_dfrbp_1 _881_ (.CLK(net200),
    .RESET_B(_014_),
    .D(_094_),
    .Q_N(_451_),
    .Q(\bsr.update_data_i[2] ));
 sg13g2_dfrbp_1 _882_ (.CLK(net200),
    .RESET_B(_015_),
    .D(_095_),
    .Q_N(_450_),
    .Q(\bsr.update_data_i[3] ));
 sg13g2_dfrbp_1 _883_ (.CLK(net202),
    .RESET_B(_016_),
    .D(_096_),
    .Q_N(_449_),
    .Q(\bsr.update_data_i[4] ));
 sg13g2_dfrbp_1 _884_ (.CLK(net201),
    .RESET_B(_017_),
    .D(_097_),
    .Q_N(_448_),
    .Q(\bsr.update_data_i[5] ));
 sg13g2_dfrbp_1 _885_ (.CLK(net201),
    .RESET_B(_018_),
    .D(_098_),
    .Q_N(_447_),
    .Q(\bsr.update_data_i[6] ));
 sg13g2_dfrbp_1 _886_ (.CLK(net199),
    .RESET_B(_019_),
    .D(_099_),
    .Q_N(_446_),
    .Q(\bsr.update_data_i[7] ));
 sg13g2_dfrbp_1 _887_ (.CLK(net201),
    .RESET_B(_020_),
    .D(_100_),
    .Q_N(_445_),
    .Q(\bsr.update_data_i[8] ));
 sg13g2_dfrbp_1 _888_ (.CLK(net198),
    .RESET_B(_021_),
    .D(_101_),
    .Q_N(_444_),
    .Q(\bsr.update_data_i[9] ));
 sg13g2_dfrbp_1 _889_ (.CLK(net192),
    .RESET_B(_022_),
    .D(_102_),
    .Q_N(_443_),
    .Q(\bsr.update_data_i[10] ));
 sg13g2_dfrbp_1 _890_ (.CLK(net192),
    .RESET_B(_023_),
    .D(_103_),
    .Q_N(_442_),
    .Q(\bsr.update_data_i[11] ));
 sg13g2_dfrbp_1 _891_ (.CLK(net192),
    .RESET_B(_024_),
    .D(_104_),
    .Q_N(_441_),
    .Q(\bsr.update_data_i[12] ));
 sg13g2_dfrbp_1 _892_ (.CLK(net192),
    .RESET_B(_025_),
    .D(_105_),
    .Q_N(_440_),
    .Q(\bsr.update_data_i[13] ));
 sg13g2_dfrbp_1 _893_ (.CLK(net203),
    .RESET_B(_026_),
    .D(_106_),
    .Q_N(_439_),
    .Q(\bsr.update_data_i[14] ));
 sg13g2_dfrbp_1 _894_ (.CLK(net198),
    .RESET_B(_027_),
    .D(_107_),
    .Q_N(_438_),
    .Q(\bsr.update_data_i[15] ));
 sg13g2_dfrbp_1 _895_ (.CLK(net198),
    .RESET_B(_028_),
    .D(_108_),
    .Q_N(_437_),
    .Q(\bsr.update_data_i[16] ));
 sg13g2_dfrbp_1 _896_ (.CLK(net198),
    .RESET_B(_029_),
    .D(_109_),
    .Q_N(_436_),
    .Q(\bsr.update_data_i[17] ));
 sg13g2_dfrbp_1 _897_ (.CLK(net198),
    .RESET_B(_030_),
    .D(_110_),
    .Q_N(_435_),
    .Q(\bsr.update_data_i[18] ));
 sg13g2_dfrbp_1 _898_ (.CLK(net195),
    .RESET_B(_031_),
    .D(_111_),
    .Q_N(_434_),
    .Q(\bsr.update_data_i[19] ));
 sg13g2_dfrbp_1 _899_ (.CLK(net195),
    .RESET_B(_032_),
    .D(_112_),
    .Q_N(_433_),
    .Q(\bsr.update_data_i[20] ));
 sg13g2_dfrbp_1 _900_ (.CLK(net195),
    .RESET_B(_033_),
    .D(_113_),
    .Q_N(_432_),
    .Q(\bsr.update_data_i[21] ));
 sg13g2_dfrbp_1 _901_ (.CLK(net195),
    .RESET_B(_034_),
    .D(_114_),
    .Q_N(_431_),
    .Q(\bsr.update_data_i[22] ));
 sg13g2_dfrbp_1 _902_ (.CLK(net193),
    .RESET_B(_035_),
    .D(_115_),
    .Q_N(_430_),
    .Q(\bsr.update_data_i[23] ));
 sg13g2_dfrbp_1 _903_ (.CLK(net193),
    .RESET_B(_036_),
    .D(_116_),
    .Q_N(_429_),
    .Q(\bsr.update_data_i[24] ));
 sg13g2_dfrbp_1 _904_ (.CLK(net194),
    .RESET_B(_037_),
    .D(_117_),
    .Q_N(_428_),
    .Q(\bsr.update_data_i[25] ));
 sg13g2_dfrbp_1 _905_ (.CLK(net194),
    .RESET_B(_038_),
    .D(_118_),
    .Q_N(_427_),
    .Q(\shift_q[26] ));
 sg13g2_dfrbp_1 _906_ (.CLK(net196),
    .RESET_B(_039_),
    .D(_119_),
    .Q_N(_426_),
    .Q(\shift_q[27] ));
 sg13g2_dfrbp_1 _907_ (.CLK(net196),
    .RESET_B(_040_),
    .D(_120_),
    .Q_N(_425_),
    .Q(\shift_q[28] ));
 sg13g2_dfrbp_1 _908_ (.CLK(net196),
    .RESET_B(_041_),
    .D(_121_),
    .Q_N(_424_),
    .Q(\shift_q[29] ));
 sg13g2_dfrbp_1 _909_ (.CLK(net196),
    .RESET_B(_042_),
    .D(_122_),
    .Q_N(_423_),
    .Q(\shift_q[30] ));
 sg13g2_dfrbp_1 _910_ (.CLK(net196),
    .RESET_B(_043_),
    .D(_123_),
    .Q_N(_422_),
    .Q(\shift_q[31] ));
 sg13g2_dfrbp_1 _911_ (.CLK(net197),
    .RESET_B(net204),
    .D(_124_),
    .Q_N(_421_),
    .Q(\tap_sm.bypass_shift_q ));
 sg13g2_dfrbp_1 _912_ (.CLK(net199),
    .RESET_B(net205),
    .D(_125_),
    .Q_N(_420_),
    .Q(\tap_sm.ir_shift_q[0] ));
 sg13g2_dfrbp_1 _913_ (.CLK(net199),
    .RESET_B(net205),
    .D(_126_),
    .Q_N(_419_),
    .Q(\tap_sm.ir_shift_q[1] ));
 sg13g2_dfrbp_1 _914_ (.CLK(net199),
    .RESET_B(net205),
    .D(_127_),
    .Q_N(_418_),
    .Q(\tap_sm.ir_shift_q[2] ));
 sg13g2_dfrbp_1 _915_ (.CLK(net199),
    .RESET_B(net204),
    .D(_128_),
    .Q_N(_417_),
    .Q(\tap_sm.ir_shift_q[3] ));
 sg13g2_dfrbp_1 _916_ (.CLK(_045_),
    .RESET_B(_044_),
    .D(_129_),
    .Q_N(_002_),
    .Q(\bsr.values[2] ));
 sg13g2_dfrbp_1 _917_ (.CLK(_047_),
    .RESET_B(_046_),
    .D(_130_),
    .Q_N(_416_),
    .Q(\bsr.values[3] ));
 sg13g2_dfrbp_1 _918_ (.CLK(_049_),
    .RESET_B(_048_),
    .D(_131_),
    .Q_N(_003_),
    .Q(\bsr.values[4] ));
 sg13g2_dfrbp_1 _919_ (.CLK(_051_),
    .RESET_B(_050_),
    .D(_132_),
    .Q_N(_005_),
    .Q(\bsr.values[5] ));
 sg13g2_dfrbp_1 _920_ (.CLK(_053_),
    .RESET_B(_052_),
    .D(_133_),
    .Q_N(_007_),
    .Q(\bsr.values[6] ));
 sg13g2_dfrbp_1 _921_ (.CLK(_055_),
    .RESET_B(_054_),
    .D(_134_),
    .Q_N(_415_),
    .Q(\bsr.values[10] ));
 sg13g2_dfrbp_1 _922_ (.CLK(_057_),
    .RESET_B(_056_),
    .D(_135_),
    .Q_N(_414_),
    .Q(\bsr.values[11] ));
 sg13g2_dfrbp_1 _923_ (.CLK(_059_),
    .RESET_B(_058_),
    .D(_136_),
    .Q_N(_413_),
    .Q(\bsr.values[12] ));
 sg13g2_dfrbp_1 _924_ (.CLK(_061_),
    .RESET_B(_060_),
    .D(_137_),
    .Q_N(_412_),
    .Q(\bsr.values[13] ));
 sg13g2_dfrbp_1 _925_ (.CLK(_063_),
    .RESET_B(_062_),
    .D(_138_),
    .Q_N(_411_),
    .Q(\bsr.values[14] ));
 sg13g2_dfrbp_1 _926_ (.CLK(_065_),
    .RESET_B(_064_),
    .D(_139_),
    .Q_N(_410_),
    .Q(\bsr.values[15] ));
 sg13g2_dfrbp_1 _927_ (.CLK(_067_),
    .RESET_B(_066_),
    .D(_140_),
    .Q_N(_409_),
    .Q(\bsr.values[16] ));
 sg13g2_dfrbp_1 _928_ (.CLK(_069_),
    .RESET_B(_068_),
    .D(_141_),
    .Q_N(_408_),
    .Q(\bsr.values[17] ));
 sg13g2_dfrbp_1 _929_ (.CLK(_071_),
    .RESET_B(_070_),
    .D(_142_),
    .Q_N(_407_),
    .Q(\bsr.values[18] ));
 sg13g2_dfrbp_1 _930_ (.CLK(_073_),
    .RESET_B(_072_),
    .D(_143_),
    .Q_N(_406_),
    .Q(\bsr.values[19] ));
 sg13g2_dfrbp_1 _931_ (.CLK(_075_),
    .RESET_B(_074_),
    .D(_144_),
    .Q_N(_405_),
    .Q(\bsr.values[20] ));
 sg13g2_dfrbp_1 _932_ (.CLK(_077_),
    .RESET_B(_076_),
    .D(_145_),
    .Q_N(_404_),
    .Q(\bsr.values[21] ));
 sg13g2_dfrbp_1 _933_ (.CLK(_079_),
    .RESET_B(_078_),
    .D(_146_),
    .Q_N(_403_),
    .Q(\bsr.values[22] ));
 sg13g2_dfrbp_1 _934_ (.CLK(_081_),
    .RESET_B(_080_),
    .D(_147_),
    .Q_N(_402_),
    .Q(\bsr.values[23] ));
 sg13g2_dfrbp_1 _935_ (.CLK(_083_),
    .RESET_B(_082_),
    .D(_148_),
    .Q_N(_401_),
    .Q(\bsr.values[24] ));
 sg13g2_dfrbp_1 _936_ (.CLK(_085_),
    .RESET_B(_084_),
    .D(_149_),
    .Q_N(_400_),
    .Q(\bsr.values[25] ));
 sg13g2_dfrbp_1 _937_ (.CLK(_086_),
    .RESET_B(net204),
    .D(_000_),
    .Q_N(_399_),
    .Q(\tap_sm.tdo_o ));
 sg13g2_dfrbp_1 _938_ (.CLK(net197),
    .RESET_B(net204),
    .D(_087_),
    .Q_N(\bsr.reset_i ),
    .Q(_011_));
 sg13g2_dfrbp_1 _939_ (.CLK(net198),
    .RESET_B(net204),
    .D(\tap_sm.state_d[0] ),
    .Q_N(_458_),
    .Q(\tap_sm.state_q[0] ));
 sg13g2_dfrbp_1 _940_ (.CLK(net197),
    .RESET_B(net204),
    .D(\tap_sm.state_d[1] ),
    .Q_N(_459_),
    .Q(\tap_sm.state_q[1] ));
 sg13g2_dfrbp_1 _941_ (.CLK(net197),
    .RESET_B(net204),
    .D(\tap_sm.state_d[2] ),
    .Q_N(_460_),
    .Q(\tap_sm.state_q[2] ));
 sg13g2_dfrbp_1 _942_ (.CLK(net197),
    .RESET_B(net204),
    .D(\tap_sm.state_d[3] ),
    .Q_N(_398_),
    .Q(\tap_sm.state_q[3] ));
 sg13g2_tielo tt_um_obriensp_jtag_16 (.L_LO(net16));
 sg13g2_tielo tt_um_obriensp_jtag_17 (.L_LO(net17));
 sg13g2_tielo tt_um_obriensp_jtag_18 (.L_LO(net18));
 sg13g2_tielo tt_um_obriensp_jtag_19 (.L_LO(net19));
 sg13g2_tielo tt_um_obriensp_jtag_20 (.L_LO(net20));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 _949_ (.A(\tap_sm.tdo_oe_o ),
    .X(uio_oe[7]));
 sg13g2_buf_2 _950_ (.A(\tap_sm.tdo_o ),
    .X(uio_out[7]));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(_370_));
 sg13g2_buf_2 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_370_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_287_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_287_),
    .X(net159));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(_287_));
 sg13g2_buf_2 fanout161 (.A(net164),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(net164),
    .X(net162));
 sg13g2_buf_1 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_205_),
    .X(net164));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(_205_));
 sg13g2_buf_1 fanout166 (.A(_205_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_247_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(net171));
 sg13g2_buf_2 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_1 fanout171 (.A(net173),
    .X(net171));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(net173));
 sg13g2_buf_2 fanout173 (.A(_221_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_206_),
    .X(net175));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(_218_));
 sg13g2_buf_2 fanout177 (.A(_218_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_217_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_217_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(\tap_sm.state_q[1] ),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(\tap_sm.state_q[0] ),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(net184),
    .X(net182));
 sg13g2_buf_1 fanout183 (.A(net184),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(net190),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(net190),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(net190),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(net190),
    .X(net187));
 sg13g2_buf_1 fanout188 (.A(net190),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(net190),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(\bsr.reset_i ),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(net13),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net194),
    .X(net193));
 sg13g2_buf_1 fanout194 (.A(net203),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(net203),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(net202),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(net201),
    .X(net199));
 sg13g2_buf_1 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(net202),
    .X(net201));
 sg13g2_buf_1 fanout202 (.A(net203),
    .X(net202));
 sg13g2_buf_1 fanout203 (.A(uio_in[4]),
    .X(net203));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(net206));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(net206));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[6]),
    .X(net14));
 sg13g2_tielo tt_um_obriensp_jtag_15 (.L_LO(net15));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_397_),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold2 (.A(\inner.counter[3] ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold3 (.A(_010_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold4 (.A(\inner.counter[2] ),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold5 (.A(_009_),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold6 (.A(\inner.counter[1] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold7 (.A(_008_),
    .X(net27));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_fill_2 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_4 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_263 ();
 sg13g2_fill_2 FILLER_16_290 ();
 sg13g2_fill_1 FILLER_16_292 ();
 sg13g2_decap_8 FILLER_16_327 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_355 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_fill_1 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_fill_2 FILLER_17_237 ();
 sg13g2_fill_1 FILLER_17_239 ();
 sg13g2_decap_8 FILLER_17_248 ();
 sg13g2_decap_8 FILLER_17_255 ();
 sg13g2_decap_8 FILLER_17_262 ();
 sg13g2_fill_1 FILLER_17_269 ();
 sg13g2_fill_1 FILLER_17_274 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_4 FILLER_17_315 ();
 sg13g2_fill_2 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_fill_1 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_248 ();
 sg13g2_fill_2 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_258 ();
 sg13g2_fill_1 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_284 ();
 sg13g2_fill_2 FILLER_18_295 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_fill_1 FILLER_18_322 ();
 sg13g2_fill_2 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_4 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_decap_4 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_238 ();
 sg13g2_fill_1 FILLER_19_261 ();
 sg13g2_decap_4 FILLER_19_275 ();
 sg13g2_fill_2 FILLER_19_279 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_308 ();
 sg13g2_fill_2 FILLER_19_333 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_264 ();
 sg13g2_decap_4 FILLER_20_279 ();
 sg13g2_fill_2 FILLER_20_283 ();
 sg13g2_decap_4 FILLER_20_304 ();
 sg13g2_fill_2 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_decap_4 FILLER_20_346 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_fill_2 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_215 ();
 sg13g2_decap_4 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_226 ();
 sg13g2_decap_4 FILLER_21_237 ();
 sg13g2_fill_2 FILLER_21_246 ();
 sg13g2_decap_4 FILLER_21_258 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_decap_8 FILLER_21_272 ();
 sg13g2_decap_8 FILLER_21_279 ();
 sg13g2_fill_1 FILLER_21_286 ();
 sg13g2_fill_2 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_300 ();
 sg13g2_fill_2 FILLER_21_307 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_316 ();
 sg13g2_decap_4 FILLER_21_358 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_4 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_247 ();
 sg13g2_fill_2 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_281 ();
 sg13g2_fill_1 FILLER_22_305 ();
 sg13g2_fill_2 FILLER_22_320 ();
 sg13g2_fill_1 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_fill_2 FILLER_22_350 ();
 sg13g2_decap_4 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_fill_2 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_145 ();
 sg13g2_decap_8 FILLER_23_152 ();
 sg13g2_fill_1 FILLER_23_159 ();
 sg13g2_decap_8 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_4 FILLER_23_203 ();
 sg13g2_fill_1 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_fill_2 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_fill_2 FILLER_23_227 ();
 sg13g2_decap_8 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_250 ();
 sg13g2_decap_4 FILLER_23_257 ();
 sg13g2_fill_1 FILLER_23_261 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_decap_4 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_317 ();
 sg13g2_decap_4 FILLER_23_327 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_decap_4 FILLER_23_363 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_decap_4 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_4 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_157 ();
 sg13g2_fill_2 FILLER_24_170 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_fill_2 FILLER_24_216 ();
 sg13g2_fill_1 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_279 ();
 sg13g2_decap_8 FILLER_24_304 ();
 sg13g2_decap_8 FILLER_24_311 ();
 sg13g2_decap_4 FILLER_24_318 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_fill_2 FILLER_24_332 ();
 sg13g2_decap_4 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_351 ();
 sg13g2_fill_2 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_91 ();
 sg13g2_fill_2 FILLER_25_131 ();
 sg13g2_fill_1 FILLER_25_133 ();
 sg13g2_decap_4 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_141 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_decap_4 FILLER_25_172 ();
 sg13g2_decap_4 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_192 ();
 sg13g2_fill_2 FILLER_25_200 ();
 sg13g2_fill_2 FILLER_25_240 ();
 sg13g2_fill_1 FILLER_25_242 ();
 sg13g2_decap_8 FILLER_25_247 ();
 sg13g2_decap_4 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_decap_4 FILLER_25_263 ();
 sg13g2_fill_2 FILLER_25_267 ();
 sg13g2_decap_8 FILLER_25_272 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_291 ();
 sg13g2_decap_4 FILLER_25_300 ();
 sg13g2_decap_4 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_314 ();
 sg13g2_decap_4 FILLER_25_344 ();
 sg13g2_fill_2 FILLER_25_351 ();
 sg13g2_fill_2 FILLER_25_358 ();
 sg13g2_fill_1 FILLER_25_360 ();
 sg13g2_fill_2 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_4 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_94 ();
 sg13g2_fill_2 FILLER_26_99 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_fill_2 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_fill_2 FILLER_26_204 ();
 sg13g2_fill_1 FILLER_26_209 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_decap_4 FILLER_26_225 ();
 sg13g2_fill_1 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_261 ();
 sg13g2_fill_1 FILLER_26_268 ();
 sg13g2_decap_4 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_313 ();
 sg13g2_fill_2 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_fill_2 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_124 ();
 sg13g2_fill_1 FILLER_27_131 ();
 sg13g2_decap_4 FILLER_27_142 ();
 sg13g2_fill_1 FILLER_27_146 ();
 sg13g2_decap_4 FILLER_27_156 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_188 ();
 sg13g2_decap_8 FILLER_27_195 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_decap_4 FILLER_27_213 ();
 sg13g2_decap_8 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_229 ();
 sg13g2_fill_2 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_decap_4 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_264 ();
 sg13g2_decap_4 FILLER_27_271 ();
 sg13g2_fill_1 FILLER_27_275 ();
 sg13g2_decap_4 FILLER_27_279 ();
 sg13g2_fill_2 FILLER_27_283 ();
 sg13g2_decap_4 FILLER_27_290 ();
 sg13g2_decap_8 FILLER_27_307 ();
 sg13g2_decap_4 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_decap_4 FILLER_27_340 ();
 sg13g2_fill_2 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_4 FILLER_27_372 ();
 sg13g2_fill_1 FILLER_27_376 ();
 sg13g2_decap_4 FILLER_27_385 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_134 ();
 sg13g2_fill_2 FILLER_28_170 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_258 ();
 sg13g2_fill_2 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_267 ();
 sg13g2_fill_2 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_103 ();
 sg13g2_fill_1 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_decap_4 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_134 ();
 sg13g2_fill_1 FILLER_29_139 ();
 sg13g2_decap_4 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_149 ();
 sg13g2_decap_8 FILLER_29_153 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_182 ();
 sg13g2_fill_2 FILLER_29_188 ();
 sg13g2_decap_8 FILLER_29_193 ();
 sg13g2_decap_4 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_4 FILLER_29_291 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_4 FILLER_29_315 ();
 sg13g2_fill_2 FILLER_29_319 ();
 sg13g2_decap_8 FILLER_29_330 ();
 sg13g2_decap_8 FILLER_29_337 ();
 sg13g2_fill_1 FILLER_29_344 ();
 sg13g2_decap_4 FILLER_29_356 ();
 sg13g2_fill_2 FILLER_29_360 ();
 sg13g2_fill_1 FILLER_29_366 ();
 sg13g2_fill_1 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_374 ();
 sg13g2_decap_4 FILLER_29_381 ();
 sg13g2_fill_2 FILLER_29_388 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_88 ();
 sg13g2_fill_2 FILLER_30_155 ();
 sg13g2_decap_4 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_264 ();
 sg13g2_decap_4 FILLER_30_271 ();
 sg13g2_decap_4 FILLER_30_290 ();
 sg13g2_fill_1 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_fill_1 FILLER_30_309 ();
 sg13g2_fill_2 FILLER_30_334 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_fill_2 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_103 ();
 sg13g2_decap_8 FILLER_31_110 ();
 sg13g2_fill_2 FILLER_31_127 ();
 sg13g2_fill_1 FILLER_31_129 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_145 ();
 sg13g2_decap_8 FILLER_31_170 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_decap_8 FILLER_31_216 ();
 sg13g2_fill_2 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_228 ();
 sg13g2_fill_2 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_243 ();
 sg13g2_fill_1 FILLER_31_245 ();
 sg13g2_decap_4 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_decap_4 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_fill_2 FILLER_31_338 ();
 sg13g2_fill_1 FILLER_31_340 ();
 sg13g2_decap_8 FILLER_31_356 ();
 sg13g2_decap_4 FILLER_31_363 ();
 sg13g2_fill_2 FILLER_31_367 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_decap_4 FILLER_32_195 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_fill_2 FILLER_32_211 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_decap_4 FILLER_32_227 ();
 sg13g2_decap_8 FILLER_32_261 ();
 sg13g2_decap_8 FILLER_32_268 ();
 sg13g2_fill_2 FILLER_32_275 ();
 sg13g2_decap_8 FILLER_32_282 ();
 sg13g2_fill_2 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_295 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_312 ();
 sg13g2_decap_4 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_116 ();
 sg13g2_decap_8 FILLER_33_122 ();
 sg13g2_fill_1 FILLER_33_129 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_137 ();
 sg13g2_fill_1 FILLER_33_142 ();
 sg13g2_decap_4 FILLER_33_152 ();
 sg13g2_fill_2 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_165 ();
 sg13g2_decap_4 FILLER_33_172 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_195 ();
 sg13g2_fill_2 FILLER_33_201 ();
 sg13g2_decap_8 FILLER_33_232 ();
 sg13g2_decap_4 FILLER_33_245 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_decap_8 FILLER_33_253 ();
 sg13g2_decap_4 FILLER_33_260 ();
 sg13g2_decap_4 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_289 ();
 sg13g2_decap_8 FILLER_33_303 ();
 sg13g2_fill_2 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_335 ();
 sg13g2_fill_2 FILLER_33_342 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_decap_4 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_128 ();
 sg13g2_fill_2 FILLER_34_197 ();
 sg13g2_decap_4 FILLER_34_207 ();
 sg13g2_fill_1 FILLER_34_211 ();
 sg13g2_decap_8 FILLER_34_215 ();
 sg13g2_decap_4 FILLER_34_222 ();
 sg13g2_fill_1 FILLER_34_226 ();
 sg13g2_fill_1 FILLER_34_234 ();
 sg13g2_fill_1 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_269 ();
 sg13g2_decap_4 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_308 ();
 sg13g2_fill_2 FILLER_34_319 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_decap_8 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_decap_4 FILLER_34_391 ();
 sg13g2_fill_2 FILLER_34_395 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_144 ();
 sg13g2_decap_8 FILLER_35_151 ();
 sg13g2_decap_8 FILLER_35_158 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_fill_2 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_174 ();
 sg13g2_fill_2 FILLER_35_270 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_fill_2 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_decap_4 FILLER_36_199 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_208 ();
 sg13g2_decap_4 FILLER_36_215 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_fill_2 FILLER_36_320 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_fill_2 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_fill_2 FILLER_37_189 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_270 ();
 sg13g2_fill_1 FILLER_37_274 ();
 sg13g2_fill_2 FILLER_37_355 ();
 sg13g2_fill_1 FILLER_37_357 ();
 sg13g2_fill_2 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_fill_1 FILLER_38_63 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_126 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_148 ();
 sg13g2_decap_8 FILLER_38_155 ();
 sg13g2_decap_8 FILLER_38_162 ();
 sg13g2_decap_8 FILLER_38_169 ();
 sg13g2_decap_8 FILLER_38_176 ();
 sg13g2_decap_8 FILLER_38_183 ();
 sg13g2_decap_8 FILLER_38_190 ();
 sg13g2_decap_8 FILLER_38_197 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_211 ();
 sg13g2_decap_4 FILLER_38_218 ();
 sg13g2_fill_1 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_4 FILLER_38_243 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_decap_4 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_fill_1 FILLER_38_312 ();
 sg13g2_fill_1 FILLER_38_318 ();
 sg13g2_fill_1 FILLER_38_340 ();
 sg13g2_fill_1 FILLER_38_384 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[4] = net15;
 assign uio_oe[5] = net16;
 assign uio_oe[6] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
endmodule

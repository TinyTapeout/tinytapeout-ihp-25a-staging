module tt_um_riscv_mini (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire \reg_file.registers[0][0] ;
 wire \reg_file.registers[0][1] ;
 wire \reg_file.registers[0][2] ;
 wire \reg_file.registers[0][3] ;
 wire \reg_file.registers[0][4] ;
 wire \reg_file.registers[0][5] ;
 wire \reg_file.registers[0][6] ;
 wire \reg_file.registers[0][7] ;
 wire \reg_file.registers[1][0] ;
 wire \reg_file.registers[1][1] ;
 wire \reg_file.registers[1][2] ;
 wire \reg_file.registers[1][3] ;
 wire \reg_file.registers[1][4] ;
 wire \reg_file.registers[1][5] ;
 wire \reg_file.registers[1][6] ;
 wire \reg_file.registers[1][7] ;
 wire \reg_file.registers[2][0] ;
 wire \reg_file.registers[2][1] ;
 wire \reg_file.registers[2][2] ;
 wire \reg_file.registers[2][3] ;
 wire \reg_file.registers[2][4] ;
 wire \reg_file.registers[2][5] ;
 wire \reg_file.registers[2][6] ;
 wire \reg_file.registers[2][7] ;
 wire \reg_file.registers[3][0] ;
 wire \reg_file.registers[3][1] ;
 wire \reg_file.registers[3][2] ;
 wire \reg_file.registers[3][3] ;
 wire \reg_file.registers[3][4] ;
 wire \reg_file.registers[3][5] ;
 wire \reg_file.registers[3][6] ;
 wire \reg_file.registers[3][7] ;
 wire \reg_file.registers[4][0] ;
 wire \reg_file.registers[4][1] ;
 wire \reg_file.registers[4][2] ;
 wire \reg_file.registers[4][3] ;
 wire \reg_file.registers[4][4] ;
 wire \reg_file.registers[4][5] ;
 wire \reg_file.registers[4][6] ;
 wire \reg_file.registers[4][7] ;
 wire \reg_file.registers[5][0] ;
 wire \reg_file.registers[5][1] ;
 wire \reg_file.registers[5][2] ;
 wire \reg_file.registers[5][3] ;
 wire \reg_file.registers[5][4] ;
 wire \reg_file.registers[5][5] ;
 wire \reg_file.registers[5][6] ;
 wire \reg_file.registers[5][7] ;
 wire \reg_file.registers[6][0] ;
 wire \reg_file.registers[6][1] ;
 wire \reg_file.registers[6][2] ;
 wire \reg_file.registers[6][3] ;
 wire \reg_file.registers[6][4] ;
 wire \reg_file.registers[6][5] ;
 wire \reg_file.registers[6][6] ;
 wire \reg_file.registers[6][7] ;
 wire \reg_file.registers[7][0] ;
 wire \reg_file.registers[7][1] ;
 wire \reg_file.registers[7][2] ;
 wire \reg_file.registers[7][3] ;
 wire \reg_file.registers[7][4] ;
 wire \reg_file.registers[7][5] ;
 wire \reg_file.registers[7][6] ;
 wire \reg_file.registers[7][7] ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire clknet_0_clk;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;

 sg13g2_inv_1 _0618_ (.Y(_0074_),
    .A(net217));
 sg13g2_inv_1 _0619_ (.Y(_0075_),
    .A(\reg_file.registers[6][0] ));
 sg13g2_inv_1 _0620_ (.Y(_0076_),
    .A(\reg_file.registers[5][0] ));
 sg13g2_inv_1 _0621_ (.Y(_0077_),
    .A(\reg_file.registers[3][0] ));
 sg13g2_inv_1 _0622_ (.Y(_0078_),
    .A(\reg_file.registers[2][0] ));
 sg13g2_inv_2 _0623_ (.Y(_0079_),
    .A(net222));
 sg13g2_inv_1 _0624_ (.Y(_0080_),
    .A(net224));
 sg13g2_inv_1 _0625_ (.Y(_0081_),
    .A(\reg_file.registers[6][1] ));
 sg13g2_inv_1 _0626_ (.Y(_0082_),
    .A(\reg_file.registers[5][1] ));
 sg13g2_inv_1 _0627_ (.Y(_0083_),
    .A(\reg_file.registers[3][1] ));
 sg13g2_inv_1 _0628_ (.Y(_0084_),
    .A(\reg_file.registers[2][1] ));
 sg13g2_inv_1 _0629_ (.Y(_0085_),
    .A(_0002_));
 sg13g2_inv_1 _0630_ (.Y(_0086_),
    .A(\reg_file.registers[0][5] ));
 sg13g2_inv_1 _0631_ (.Y(_0087_),
    .A(\reg_file.registers[0][6] ));
 sg13g2_nor2_2 _0632_ (.A(net216),
    .B(net12),
    .Y(_0088_));
 sg13g2_nor2b_2 _0633_ (.A(net2),
    .B_N(net1),
    .Y(_0089_));
 sg13g2_nand2b_2 _0634_ (.Y(_0090_),
    .B(net1),
    .A_N(net2));
 sg13g2_nand2_1 _0635_ (.Y(_0091_),
    .A(net10),
    .B(_0090_));
 sg13g2_a21oi_2 _0636_ (.B1(net212),
    .Y(_0092_),
    .A2(_0090_),
    .A1(net10));
 sg13g2_and2_1 _0637_ (.A(_0088_),
    .B(_0092_),
    .X(_0093_));
 sg13g2_nand2_2 _0638_ (.Y(_0094_),
    .A(_0088_),
    .B(_0092_));
 sg13g2_and3_2 _0639_ (.X(_0095_),
    .A(net220),
    .B(net218),
    .C(_0074_));
 sg13g2_nand3b_1 _0640_ (.B(net219),
    .C(net221),
    .Y(_0096_),
    .A_N(net9));
 sg13g2_nand2b_2 _0641_ (.Y(_0097_),
    .B(net218),
    .A_N(net220));
 sg13g2_nor2_2 _0642_ (.A(net217),
    .B(_0097_),
    .Y(_0098_));
 sg13g2_nor2_2 _0643_ (.A(_0074_),
    .B(_0097_),
    .Y(_0099_));
 sg13g2_nand3b_1 _0644_ (.B(net219),
    .C(net9),
    .Y(_0100_),
    .A_N(net221));
 sg13g2_and3_2 _0645_ (.X(_0101_),
    .A(net220),
    .B(net218),
    .C(net217));
 sg13g2_nor2_2 _0646_ (.A(net220),
    .B(net218),
    .Y(_0102_));
 sg13g2_nor3_1 _0647_ (.A(net220),
    .B(net218),
    .C(net217),
    .Y(_0103_));
 sg13g2_inv_1 _0648_ (.Y(_0104_),
    .A(net210));
 sg13g2_a21o_1 _0649_ (.A2(_0102_),
    .A1(\reg_file.registers[4][7] ),
    .B1(net210),
    .X(_0105_));
 sg13g2_nor2b_1 _0650_ (.A(net218),
    .B_N(net220),
    .Y(_0106_));
 sg13g2_and2_2 _0651_ (.A(net217),
    .B(_0106_),
    .X(_0107_));
 sg13g2_nand3b_1 _0652_ (.B(net9),
    .C(net220),
    .Y(_0108_),
    .A_N(net218));
 sg13g2_and2_2 _0653_ (.A(_0074_),
    .B(_0106_),
    .X(_0109_));
 sg13g2_a221oi_1 _0654_ (.B2(\reg_file.registers[1][7] ),
    .C1(_0105_),
    .B1(_0109_),
    .A1(\reg_file.registers[5][7] ),
    .Y(_0110_),
    .A2(_0107_));
 sg13g2_a22oi_1 _0655_ (.Y(_0111_),
    .B1(_0099_),
    .B2(\reg_file.registers[6][7] ),
    .A2(_0095_),
    .A1(\reg_file.registers[3][7] ));
 sg13g2_a22oi_1 _0656_ (.Y(_0112_),
    .B1(_0101_),
    .B2(\reg_file.registers[7][7] ),
    .A2(_0098_),
    .A1(\reg_file.registers[2][7] ));
 sg13g2_nand3_1 _0657_ (.B(_0111_),
    .C(_0112_),
    .A(_0110_),
    .Y(_0113_));
 sg13g2_a21oi_1 _0658_ (.A1(_0005_),
    .A2(net209),
    .Y(_0114_),
    .B1(net211));
 sg13g2_nand2_1 _0659_ (.Y(_0115_),
    .A(_0113_),
    .B(_0114_));
 sg13g2_nor2_2 _0660_ (.A(net223),
    .B(net224),
    .Y(_0116_));
 sg13g2_and2_1 _0661_ (.A(net222),
    .B(_0116_),
    .X(_0117_));
 sg13g2_nand2b_2 _0662_ (.Y(_0118_),
    .B(net223),
    .A_N(net224));
 sg13g2_nor2_2 _0663_ (.A(net222),
    .B(_0118_),
    .Y(_0119_));
 sg13g2_nor2_2 _0664_ (.A(_0079_),
    .B(_0118_),
    .Y(_0120_));
 sg13g2_nand3b_1 _0665_ (.B(net7),
    .C(net222),
    .Y(_0121_),
    .A_N(net6));
 sg13g2_and3_2 _0666_ (.X(_0122_),
    .A(_0079_),
    .B(net223),
    .C(net224));
 sg13g2_nand3b_1 _0667_ (.B(net7),
    .C(net224),
    .Y(_0123_),
    .A_N(net222));
 sg13g2_and3_2 _0668_ (.X(_0124_),
    .A(net222),
    .B(net223),
    .C(net224));
 sg13g2_nor3_2 _0669_ (.A(net8),
    .B(net223),
    .C(net224),
    .Y(_0125_));
 sg13g2_nand2_2 _0670_ (.Y(_0126_),
    .A(_0079_),
    .B(_0116_));
 sg13g2_nor3_2 _0671_ (.A(net8),
    .B(net223),
    .C(_0080_),
    .Y(_0127_));
 sg13g2_nor3_2 _0672_ (.A(_0079_),
    .B(net223),
    .C(_0080_),
    .Y(_0128_));
 sg13g2_a22oi_1 _0673_ (.Y(_0129_),
    .B1(_0120_),
    .B2(\reg_file.registers[6][7] ),
    .A2(_0117_),
    .A1(\reg_file.registers[4][7] ));
 sg13g2_a22oi_1 _0674_ (.Y(_0130_),
    .B1(_0128_),
    .B2(\reg_file.registers[5][7] ),
    .A2(_0122_),
    .A1(\reg_file.registers[3][7] ));
 sg13g2_a22oi_1 _0675_ (.Y(_0131_),
    .B1(_0127_),
    .B2(\reg_file.registers[1][7] ),
    .A2(_0124_),
    .A1(\reg_file.registers[7][7] ));
 sg13g2_a21oi_1 _0676_ (.A1(\reg_file.registers[2][7] ),
    .A2(_0119_),
    .Y(_0132_),
    .B1(net208));
 sg13g2_nand4_1 _0677_ (.B(_0130_),
    .C(_0131_),
    .A(_0129_),
    .Y(_0133_),
    .D(_0132_));
 sg13g2_o21ai_1 _0678_ (.B1(_0133_),
    .Y(_0134_),
    .A1(\reg_file.registers[0][7] ),
    .A2(_0126_));
 sg13g2_inv_1 _0679_ (.Y(_0135_),
    .A(_0134_));
 sg13g2_nor2_1 _0680_ (.A(_0115_),
    .B(_0134_),
    .Y(_0136_));
 sg13g2_and2_1 _0681_ (.A(_0115_),
    .B(_0134_),
    .X(_0137_));
 sg13g2_nor2_2 _0682_ (.A(_0136_),
    .B(_0137_),
    .Y(_0138_));
 sg13g2_inv_1 _0683_ (.Y(_0139_),
    .A(_0138_));
 sg13g2_nand2_1 _0684_ (.Y(_0140_),
    .A(\reg_file.registers[3][6] ),
    .B(_0095_));
 sg13g2_a22oi_1 _0685_ (.Y(_0141_),
    .B1(_0101_),
    .B2(\reg_file.registers[7][6] ),
    .A2(_0098_),
    .A1(\reg_file.registers[2][6] ));
 sg13g2_a22oi_1 _0686_ (.Y(_0142_),
    .B1(_0107_),
    .B2(\reg_file.registers[5][6] ),
    .A2(_0099_),
    .A1(\reg_file.registers[6][6] ));
 sg13g2_a221oi_1 _0687_ (.B2(\reg_file.registers[1][6] ),
    .C1(net209),
    .B1(_0109_),
    .A1(\reg_file.registers[4][6] ),
    .Y(_0143_),
    .A2(_0102_));
 sg13g2_nand4_1 _0688_ (.B(_0141_),
    .C(_0142_),
    .A(_0140_),
    .Y(_0144_),
    .D(_0143_));
 sg13g2_a21oi_1 _0689_ (.A1(_0006_),
    .A2(net209),
    .Y(_0145_),
    .B1(net211));
 sg13g2_nand2_2 _0690_ (.Y(_0146_),
    .A(_0144_),
    .B(_0145_));
 sg13g2_a22oi_1 _0691_ (.Y(_0147_),
    .B1(_0120_),
    .B2(\reg_file.registers[6][6] ),
    .A2(_0119_),
    .A1(\reg_file.registers[2][6] ));
 sg13g2_a21oi_1 _0692_ (.A1(\reg_file.registers[3][6] ),
    .A2(_0122_),
    .Y(_0148_),
    .B1(net208));
 sg13g2_a22oi_1 _0693_ (.Y(_0149_),
    .B1(_0128_),
    .B2(\reg_file.registers[5][6] ),
    .A2(_0124_),
    .A1(\reg_file.registers[7][6] ));
 sg13g2_a22oi_1 _0694_ (.Y(_0150_),
    .B1(_0127_),
    .B2(\reg_file.registers[1][6] ),
    .A2(_0117_),
    .A1(\reg_file.registers[4][6] ));
 sg13g2_and3_1 _0695_ (.X(_0151_),
    .A(_0148_),
    .B(_0149_),
    .C(_0150_));
 sg13g2_a22oi_1 _0696_ (.Y(_0152_),
    .B1(_0147_),
    .B2(_0151_),
    .A2(net208),
    .A1(_0087_));
 sg13g2_inv_1 _0697_ (.Y(_0153_),
    .A(_0152_));
 sg13g2_nand2_2 _0698_ (.Y(_0154_),
    .A(_0146_),
    .B(_0152_));
 sg13g2_nor2_1 _0699_ (.A(_0146_),
    .B(_0153_),
    .Y(_0155_));
 sg13g2_nor2_1 _0700_ (.A(_0146_),
    .B(_0152_),
    .Y(_0156_));
 sg13g2_inv_1 _0701_ (.Y(_0157_),
    .A(_0156_));
 sg13g2_nand2_2 _0702_ (.Y(_0158_),
    .A(_0154_),
    .B(_0157_));
 sg13g2_nand2_1 _0703_ (.Y(_0159_),
    .A(\reg_file.registers[2][5] ),
    .B(_0098_));
 sg13g2_a22oi_1 _0704_ (.Y(_0160_),
    .B1(_0107_),
    .B2(\reg_file.registers[5][5] ),
    .A2(_0095_),
    .A1(\reg_file.registers[3][5] ));
 sg13g2_a22oi_1 _0705_ (.Y(_0161_),
    .B1(_0109_),
    .B2(\reg_file.registers[1][5] ),
    .A2(_0099_),
    .A1(\reg_file.registers[6][5] ));
 sg13g2_a221oi_1 _0706_ (.B2(\reg_file.registers[4][5] ),
    .C1(net210),
    .B1(_0102_),
    .A1(\reg_file.registers[7][5] ),
    .Y(_0162_),
    .A2(_0101_));
 sg13g2_nand4_1 _0707_ (.B(_0160_),
    .C(_0161_),
    .A(_0159_),
    .Y(_0163_),
    .D(_0162_));
 sg13g2_a21oi_1 _0708_ (.A1(_0007_),
    .A2(net209),
    .Y(_0164_),
    .B1(net211));
 sg13g2_nand2_2 _0709_ (.Y(_0165_),
    .A(_0163_),
    .B(_0164_));
 sg13g2_a22oi_1 _0710_ (.Y(_0166_),
    .B1(_0124_),
    .B2(\reg_file.registers[7][5] ),
    .A2(_0120_),
    .A1(\reg_file.registers[6][5] ));
 sg13g2_a22oi_1 _0711_ (.Y(_0167_),
    .B1(_0128_),
    .B2(\reg_file.registers[5][5] ),
    .A2(_0119_),
    .A1(\reg_file.registers[2][5] ));
 sg13g2_o21ai_1 _0712_ (.B1(_0116_),
    .Y(_0168_),
    .A1(_0079_),
    .A2(\reg_file.registers[4][5] ));
 sg13g2_nand2_1 _0713_ (.Y(_0169_),
    .A(_0166_),
    .B(_0168_));
 sg13g2_a221oi_1 _0714_ (.B2(\reg_file.registers[1][5] ),
    .C1(_0169_),
    .B1(_0127_),
    .A1(\reg_file.registers[3][5] ),
    .Y(_0170_),
    .A2(_0122_));
 sg13g2_a22oi_1 _0715_ (.Y(_0171_),
    .B1(_0167_),
    .B2(_0170_),
    .A2(net208),
    .A1(_0086_));
 sg13g2_inv_1 _0716_ (.Y(_0172_),
    .A(_0171_));
 sg13g2_nand2_1 _0717_ (.Y(_0173_),
    .A(_0165_),
    .B(_0171_));
 sg13g2_inv_1 _0718_ (.Y(_0174_),
    .A(_0173_));
 sg13g2_or2_1 _0719_ (.X(_0175_),
    .B(_0171_),
    .A(_0165_));
 sg13g2_inv_1 _0720_ (.Y(_0176_),
    .A(_0175_));
 sg13g2_nand2_1 _0721_ (.Y(_0177_),
    .A(\reg_file.registers[1][4] ),
    .B(_0109_));
 sg13g2_a22oi_1 _0722_ (.Y(_0178_),
    .B1(_0101_),
    .B2(\reg_file.registers[7][4] ),
    .A2(_0098_),
    .A1(\reg_file.registers[2][4] ));
 sg13g2_a22oi_1 _0723_ (.Y(_0179_),
    .B1(_0099_),
    .B2(\reg_file.registers[6][4] ),
    .A2(_0095_),
    .A1(\reg_file.registers[3][4] ));
 sg13g2_a22oi_1 _0724_ (.Y(_0180_),
    .B1(_0107_),
    .B2(\reg_file.registers[5][4] ),
    .A2(_0102_),
    .A1(\reg_file.registers[4][4] ));
 sg13g2_and4_1 _0725_ (.A(_0104_),
    .B(_0177_),
    .C(_0178_),
    .D(_0180_),
    .X(_0181_));
 sg13g2_a221oi_1 _0726_ (.B2(_0181_),
    .C1(_0089_),
    .B1(_0179_),
    .A1(_0008_),
    .Y(_0182_),
    .A2(net210));
 sg13g2_a21o_2 _0727_ (.A2(_0089_),
    .A1(net11),
    .B1(_0182_),
    .X(_0183_));
 sg13g2_nand2_1 _0728_ (.Y(_0184_),
    .A(\reg_file.registers[2][4] ),
    .B(_0119_));
 sg13g2_a22oi_1 _0729_ (.Y(_0185_),
    .B1(_0127_),
    .B2(\reg_file.registers[1][4] ),
    .A2(_0120_),
    .A1(\reg_file.registers[6][4] ));
 sg13g2_a221oi_1 _0730_ (.B2(\reg_file.registers[5][4] ),
    .C1(_0125_),
    .B1(_0128_),
    .A1(\reg_file.registers[4][4] ),
    .Y(_0186_),
    .A2(_0116_));
 sg13g2_a22oi_1 _0731_ (.Y(_0187_),
    .B1(_0124_),
    .B2(\reg_file.registers[7][4] ),
    .A2(_0122_),
    .A1(\reg_file.registers[3][4] ));
 sg13g2_nand4_1 _0732_ (.B(_0185_),
    .C(_0186_),
    .A(_0184_),
    .Y(_0188_),
    .D(_0187_));
 sg13g2_o21ai_1 _0733_ (.B1(_0188_),
    .Y(_0189_),
    .A1(\reg_file.registers[0][4] ),
    .A2(_0126_));
 sg13g2_or2_1 _0734_ (.X(_0190_),
    .B(net187),
    .A(_0183_));
 sg13g2_inv_1 _0735_ (.Y(_0191_),
    .A(_0190_));
 sg13g2_and2_1 _0736_ (.A(net10),
    .B(net211),
    .X(_0192_));
 sg13g2_nand2_1 _0737_ (.Y(_0193_),
    .A(\reg_file.registers[1][3] ),
    .B(_0109_));
 sg13g2_a22oi_1 _0738_ (.Y(_0194_),
    .B1(_0098_),
    .B2(\reg_file.registers[2][3] ),
    .A2(_0095_),
    .A1(\reg_file.registers[3][3] ));
 sg13g2_a221oi_1 _0739_ (.B2(\reg_file.registers[4][3] ),
    .C1(net210),
    .B1(_0102_),
    .A1(\reg_file.registers[7][3] ),
    .Y(_0195_),
    .A2(_0101_));
 sg13g2_a22oi_1 _0740_ (.Y(_0196_),
    .B1(_0107_),
    .B2(\reg_file.registers[5][3] ),
    .A2(_0099_),
    .A1(\reg_file.registers[6][3] ));
 sg13g2_nand4_1 _0741_ (.B(_0194_),
    .C(_0195_),
    .A(_0193_),
    .Y(_0197_),
    .D(_0196_));
 sg13g2_a21oi_1 _0742_ (.A1(_0009_),
    .A2(net209),
    .Y(_0198_),
    .B1(net211));
 sg13g2_a21o_2 _0743_ (.A2(_0198_),
    .A1(_0197_),
    .B1(_0192_),
    .X(_0199_));
 sg13g2_a22oi_1 _0744_ (.Y(_0200_),
    .B1(_0120_),
    .B2(\reg_file.registers[6][3] ),
    .A2(_0117_),
    .A1(\reg_file.registers[4][3] ));
 sg13g2_a22oi_1 _0745_ (.Y(_0201_),
    .B1(_0127_),
    .B2(\reg_file.registers[1][3] ),
    .A2(_0124_),
    .A1(\reg_file.registers[7][3] ));
 sg13g2_and2_1 _0746_ (.A(_0200_),
    .B(_0201_),
    .X(_0202_));
 sg13g2_a21o_1 _0747_ (.A2(_0128_),
    .A1(\reg_file.registers[5][3] ),
    .B1(net208),
    .X(_0203_));
 sg13g2_a221oi_1 _0748_ (.B2(\reg_file.registers[3][3] ),
    .C1(_0203_),
    .B1(_0122_),
    .A1(\reg_file.registers[2][3] ),
    .Y(_0204_),
    .A2(_0119_));
 sg13g2_nor2_1 _0749_ (.A(\reg_file.registers[0][3] ),
    .B(_0126_),
    .Y(_0205_));
 sg13g2_a21oi_2 _0750_ (.B1(_0205_),
    .Y(_0206_),
    .A2(_0204_),
    .A1(_0202_));
 sg13g2_a21o_2 _0751_ (.A2(_0204_),
    .A1(_0202_),
    .B1(_0205_),
    .X(_0207_));
 sg13g2_nand2b_1 _0752_ (.Y(_0208_),
    .B(_0206_),
    .A_N(_0199_));
 sg13g2_and2_1 _0753_ (.A(_0199_),
    .B(_0207_),
    .X(_0209_));
 sg13g2_nor2_1 _0754_ (.A(_0074_),
    .B(_0090_),
    .Y(_0210_));
 sg13g2_nor2b_1 _0755_ (.A(_0003_),
    .B_N(_0101_),
    .Y(_0211_));
 sg13g2_a221oi_1 _0756_ (.B2(\reg_file.registers[5][2] ),
    .C1(_0211_),
    .B1(_0107_),
    .A1(\reg_file.registers[2][2] ),
    .Y(_0212_),
    .A2(_0098_));
 sg13g2_a221oi_1 _0757_ (.B2(\reg_file.registers[4][2] ),
    .C1(net210),
    .B1(_0102_),
    .A1(\reg_file.registers[3][2] ),
    .Y(_0213_),
    .A2(_0095_));
 sg13g2_a22oi_1 _0758_ (.Y(_0214_),
    .B1(_0109_),
    .B2(\reg_file.registers[1][2] ),
    .A2(_0099_),
    .A1(\reg_file.registers[6][2] ));
 sg13g2_nand3_1 _0759_ (.B(_0213_),
    .C(_0214_),
    .A(_0212_),
    .Y(_0215_));
 sg13g2_a21oi_1 _0760_ (.A1(_0002_),
    .A2(net209),
    .Y(_0216_),
    .B1(net211));
 sg13g2_a21oi_1 _0761_ (.A1(_0215_),
    .A2(_0216_),
    .Y(_0217_),
    .B1(_0210_));
 sg13g2_a21o_2 _0762_ (.A2(_0216_),
    .A1(_0215_),
    .B1(_0210_),
    .X(_0218_));
 sg13g2_nor2b_1 _0763_ (.A(_0003_),
    .B_N(_0124_),
    .Y(_0219_));
 sg13g2_a221oi_1 _0764_ (.B2(\reg_file.registers[3][2] ),
    .C1(_0219_),
    .B1(_0122_),
    .A1(\reg_file.registers[2][2] ),
    .Y(_0220_),
    .A2(_0119_));
 sg13g2_a22oi_1 _0765_ (.Y(_0221_),
    .B1(_0128_),
    .B2(\reg_file.registers[5][2] ),
    .A2(_0127_),
    .A1(\reg_file.registers[1][2] ));
 sg13g2_a221oi_1 _0766_ (.B2(\reg_file.registers[6][2] ),
    .C1(net208),
    .B1(_0120_),
    .A1(\reg_file.registers[4][2] ),
    .Y(_0222_),
    .A2(_0116_));
 sg13g2_nand3_1 _0767_ (.B(_0221_),
    .C(_0222_),
    .A(_0220_),
    .Y(_0223_));
 sg13g2_o21ai_1 _0768_ (.B1(_0223_),
    .Y(_0224_),
    .A1(_0085_),
    .A2(_0126_));
 sg13g2_nor2_1 _0769_ (.A(_0218_),
    .B(_0224_),
    .Y(_0225_));
 sg13g2_nor2_1 _0770_ (.A(net186),
    .B(_0224_),
    .Y(_0226_));
 sg13g2_nand2_1 _0771_ (.Y(_0227_),
    .A(net186),
    .B(_0224_));
 sg13g2_and2_1 _0772_ (.A(_0218_),
    .B(_0224_),
    .X(_0228_));
 sg13g2_nor2_2 _0773_ (.A(_0225_),
    .B(_0228_),
    .Y(_0229_));
 sg13g2_nor2_1 _0774_ (.A(_0082_),
    .B(_0108_),
    .Y(_0230_));
 sg13g2_and2_1 _0775_ (.A(\reg_file.registers[4][1] ),
    .B(_0102_),
    .X(_0231_));
 sg13g2_nor2_1 _0776_ (.A(_0083_),
    .B(_0096_),
    .Y(_0232_));
 sg13g2_nand4_1 _0777_ (.B(net219),
    .C(net217),
    .A(net220),
    .Y(_0233_),
    .D(\reg_file.registers[7][1] ));
 sg13g2_a221oi_1 _0778_ (.B2(\reg_file.registers[1][1] ),
    .C1(_0230_),
    .B1(_0109_),
    .A1(\reg_file.registers[2][1] ),
    .Y(_0234_),
    .A2(_0098_));
 sg13g2_o21ai_1 _0779_ (.B1(_0233_),
    .Y(_0235_),
    .A1(_0081_),
    .A2(_0100_));
 sg13g2_nor4_1 _0780_ (.A(net210),
    .B(_0231_),
    .C(_0232_),
    .D(_0235_),
    .Y(_0236_));
 sg13g2_o21ai_1 _0781_ (.B1(_0090_),
    .Y(_0237_),
    .A1(\reg_file.registers[0][1] ),
    .A2(_0104_));
 sg13g2_a21o_1 _0782_ (.A2(_0236_),
    .A1(_0234_),
    .B1(_0237_),
    .X(_0238_));
 sg13g2_nand2_1 _0783_ (.Y(_0239_),
    .A(net219),
    .B(net211));
 sg13g2_and2_1 _0784_ (.A(_0238_),
    .B(_0239_),
    .X(_0240_));
 sg13g2_and2_1 _0785_ (.A(_0004_),
    .B(net208),
    .X(_0241_));
 sg13g2_nor4_1 _0786_ (.A(_0079_),
    .B(net223),
    .C(_0080_),
    .D(_0082_),
    .Y(_0242_));
 sg13g2_nor3_1 _0787_ (.A(net8),
    .B(_0084_),
    .C(_0118_),
    .Y(_0243_));
 sg13g2_nand4_1 _0788_ (.B(net7),
    .C(net224),
    .A(net222),
    .Y(_0244_),
    .D(\reg_file.registers[7][1] ));
 sg13g2_nor2_1 _0789_ (.A(_0083_),
    .B(_0123_),
    .Y(_0245_));
 sg13g2_a221oi_1 _0790_ (.B2(\reg_file.registers[1][1] ),
    .C1(_0125_),
    .B1(_0127_),
    .A1(\reg_file.registers[4][1] ),
    .Y(_0246_),
    .A2(_0116_));
 sg13g2_o21ai_1 _0791_ (.B1(_0244_),
    .Y(_0247_),
    .A1(_0081_),
    .A2(_0121_));
 sg13g2_nor4_2 _0792_ (.A(_0242_),
    .B(_0243_),
    .C(_0245_),
    .Y(_0248_),
    .D(_0247_));
 sg13g2_a21oi_1 _0793_ (.A1(_0246_),
    .A2(_0248_),
    .Y(_0249_),
    .B1(_0241_));
 sg13g2_a21o_2 _0794_ (.A2(_0248_),
    .A1(_0246_),
    .B1(_0241_),
    .X(_0250_));
 sg13g2_a21oi_2 _0795_ (.B1(_0250_),
    .Y(_0251_),
    .A2(_0239_),
    .A1(_0238_));
 sg13g2_nand3_1 _0796_ (.B(_0239_),
    .C(_0250_),
    .A(_0238_),
    .Y(_0252_));
 sg13g2_nor2b_2 _0797_ (.A(_0251_),
    .B_N(_0252_),
    .Y(_0253_));
 sg13g2_nand2b_1 _0798_ (.Y(_0254_),
    .B(_0252_),
    .A_N(_0251_));
 sg13g2_nand2_2 _0799_ (.Y(_0255_),
    .A(net221),
    .B(net211));
 sg13g2_nor2b_1 _0800_ (.A(_0001_),
    .B_N(_0101_),
    .Y(_0256_));
 sg13g2_a221oi_1 _0801_ (.B2(\reg_file.registers[1][0] ),
    .C1(_0256_),
    .B1(_0109_),
    .A1(\reg_file.registers[6][0] ),
    .Y(_0257_),
    .A2(_0099_));
 sg13g2_nor2_1 _0802_ (.A(_0076_),
    .B(_0108_),
    .Y(_0258_));
 sg13g2_a21o_1 _0803_ (.A2(_0102_),
    .A1(\reg_file.registers[4][0] ),
    .B1(net209),
    .X(_0259_));
 sg13g2_nor3_1 _0804_ (.A(net217),
    .B(_0078_),
    .C(_0097_),
    .Y(_0260_));
 sg13g2_nor2_1 _0805_ (.A(_0077_),
    .B(_0096_),
    .Y(_0261_));
 sg13g2_nor4_1 _0806_ (.A(_0258_),
    .B(_0259_),
    .C(_0260_),
    .D(_0261_),
    .Y(_0262_));
 sg13g2_a21o_1 _0807_ (.A2(net209),
    .A1(_0000_),
    .B1(_0089_),
    .X(_0263_));
 sg13g2_a21o_1 _0808_ (.A2(_0262_),
    .A1(_0257_),
    .B1(_0263_),
    .X(_0264_));
 sg13g2_nand2_1 _0809_ (.Y(_0265_),
    .A(_0255_),
    .B(_0264_));
 sg13g2_inv_1 _0810_ (.Y(_0266_),
    .A(net178));
 sg13g2_nor2_1 _0811_ (.A(_0075_),
    .B(_0121_),
    .Y(_0267_));
 sg13g2_a221oi_1 _0812_ (.B2(\reg_file.registers[5][0] ),
    .C1(_0267_),
    .B1(_0128_),
    .A1(\reg_file.registers[1][0] ),
    .Y(_0268_),
    .A2(_0127_));
 sg13g2_nor2b_1 _0813_ (.A(_0001_),
    .B_N(_0124_),
    .Y(_0269_));
 sg13g2_a21o_1 _0814_ (.A2(_0116_),
    .A1(\reg_file.registers[4][0] ),
    .B1(_0125_),
    .X(_0270_));
 sg13g2_nor3_1 _0815_ (.A(_0078_),
    .B(net222),
    .C(_0118_),
    .Y(_0271_));
 sg13g2_nor2_1 _0816_ (.A(_0077_),
    .B(_0123_),
    .Y(_0272_));
 sg13g2_nor4_2 _0817_ (.A(_0269_),
    .B(_0270_),
    .C(_0271_),
    .Y(_0273_),
    .D(_0272_));
 sg13g2_and2_1 _0818_ (.A(_0000_),
    .B(net208),
    .X(_0274_));
 sg13g2_a21oi_1 _0819_ (.A1(_0268_),
    .A2(_0273_),
    .Y(_0275_),
    .B1(_0274_));
 sg13g2_a21o_1 _0820_ (.A2(_0273_),
    .A1(_0268_),
    .B1(_0274_),
    .X(_0276_));
 sg13g2_a21o_1 _0821_ (.A2(_0264_),
    .A1(_0255_),
    .B1(_0275_),
    .X(_0277_));
 sg13g2_and2_1 _0822_ (.A(net183),
    .B(_0249_),
    .X(_0278_));
 sg13g2_a21o_2 _0823_ (.A2(_0277_),
    .A1(_0254_),
    .B1(_0278_),
    .X(_0279_));
 sg13g2_a21oi_2 _0824_ (.B1(_0225_),
    .Y(_0280_),
    .A2(_0279_),
    .A1(_0229_));
 sg13g2_a21oi_1 _0825_ (.A1(_0208_),
    .A2(_0280_),
    .Y(_0281_),
    .B1(_0209_));
 sg13g2_a221oi_1 _0826_ (.B2(_0280_),
    .C1(_0209_),
    .B1(_0208_),
    .A1(_0183_),
    .Y(_0282_),
    .A2(net187));
 sg13g2_nor2b_2 _0827_ (.A(net187),
    .B_N(_0183_),
    .Y(_0283_));
 sg13g2_nand2b_1 _0828_ (.Y(_0284_),
    .B(net187),
    .A_N(_0183_));
 sg13g2_nand2b_1 _0829_ (.Y(_0285_),
    .B(_0284_),
    .A_N(_0283_));
 sg13g2_nor2b_2 _0830_ (.A(_0283_),
    .B_N(_0284_),
    .Y(_0286_));
 sg13g2_nor2_1 _0831_ (.A(_0191_),
    .B(_0282_),
    .Y(_0287_));
 sg13g2_or3_1 _0832_ (.A(_0174_),
    .B(_0191_),
    .C(_0282_),
    .X(_0288_));
 sg13g2_and2_1 _0833_ (.A(_0175_),
    .B(_0288_),
    .X(_0289_));
 sg13g2_nand4_1 _0834_ (.B(_0157_),
    .C(_0175_),
    .A(_0154_),
    .Y(_0290_),
    .D(_0288_));
 sg13g2_a21o_1 _0835_ (.A2(_0290_),
    .A1(_0154_),
    .B1(_0138_),
    .X(_0291_));
 sg13g2_nand3_1 _0836_ (.B(_0154_),
    .C(_0290_),
    .A(_0138_),
    .Y(_0292_));
 sg13g2_and2_2 _0837_ (.A(net213),
    .B(_0092_),
    .X(_0293_));
 sg13g2_nand2_1 _0838_ (.Y(_0294_),
    .A(net213),
    .B(_0092_));
 sg13g2_nand2_1 _0839_ (.Y(_0295_),
    .A(net216),
    .B(net12));
 sg13g2_and2_2 _0840_ (.A(net214),
    .B(_0293_),
    .X(_0296_));
 sg13g2_nand3_1 _0841_ (.B(_0292_),
    .C(_0296_),
    .A(_0291_),
    .Y(_0297_));
 sg13g2_nand2b_1 _0842_ (.Y(_0298_),
    .B(_0171_),
    .A_N(_0165_));
 sg13g2_nor2_2 _0843_ (.A(_0174_),
    .B(_0176_),
    .Y(_0299_));
 sg13g2_and2_1 _0844_ (.A(_0199_),
    .B(_0206_),
    .X(_0300_));
 sg13g2_inv_1 _0845_ (.Y(_0301_),
    .A(_0300_));
 sg13g2_a21oi_2 _0846_ (.B1(_0276_),
    .Y(_0302_),
    .A2(_0264_),
    .A1(_0255_));
 sg13g2_a21o_1 _0847_ (.A2(_0302_),
    .A1(_0252_),
    .B1(_0251_),
    .X(_0303_));
 sg13g2_a21oi_1 _0848_ (.A1(_0227_),
    .A2(_0303_),
    .Y(_0304_),
    .B1(_0226_));
 sg13g2_nand2b_1 _0849_ (.Y(_0305_),
    .B(_0207_),
    .A_N(_0199_));
 sg13g2_xnor2_1 _0850_ (.Y(_0306_),
    .A(_0199_),
    .B(_0206_));
 sg13g2_o21ai_1 _0851_ (.B1(_0301_),
    .Y(_0307_),
    .A1(_0304_),
    .A2(_0306_));
 sg13g2_a21oi_1 _0852_ (.A1(_0286_),
    .A2(_0307_),
    .Y(_0308_),
    .B1(_0283_));
 sg13g2_o21ai_1 _0853_ (.B1(_0298_),
    .Y(_0309_),
    .A1(_0299_),
    .A2(_0308_));
 sg13g2_a21oi_1 _0854_ (.A1(_0158_),
    .A2(_0309_),
    .Y(_0310_),
    .B1(_0155_));
 sg13g2_nand2b_1 _0855_ (.Y(_0311_),
    .B(net213),
    .A_N(net215));
 sg13g2_nor2_2 _0856_ (.A(net214),
    .B(_0294_),
    .Y(_0312_));
 sg13g2_nand2b_2 _0857_ (.Y(_0313_),
    .B(_0293_),
    .A_N(net214));
 sg13g2_xnor2_1 _0858_ (.Y(_0314_),
    .A(_0138_),
    .B(_0310_));
 sg13g2_nor2b_1 _0859_ (.A(net213),
    .B_N(net214),
    .Y(_0315_));
 sg13g2_nand2b_1 _0860_ (.Y(_0316_),
    .B(net215),
    .A_N(net213));
 sg13g2_and2_1 _0861_ (.A(_0092_),
    .B(_0315_),
    .X(_0317_));
 sg13g2_nand2_1 _0862_ (.Y(_0318_),
    .A(_0092_),
    .B(_0315_));
 sg13g2_nand2_2 _0863_ (.Y(_0319_),
    .A(net212),
    .B(_0091_));
 sg13g2_nor2_1 _0864_ (.A(net213),
    .B(_0319_),
    .Y(_0320_));
 sg13g2_nor3_2 _0865_ (.A(net215),
    .B(net213),
    .C(_0319_),
    .Y(_0321_));
 sg13g2_nand3_1 _0866_ (.B(_0088_),
    .C(_0091_),
    .A(net212),
    .Y(_0322_));
 sg13g2_nand2b_2 _0867_ (.Y(_0323_),
    .B(net184),
    .A_N(net182));
 sg13g2_inv_1 _0868_ (.Y(_0324_),
    .A(_0323_));
 sg13g2_nand2_1 _0869_ (.Y(_0325_),
    .A(net187),
    .B(net179));
 sg13g2_o21ai_1 _0870_ (.B1(_0325_),
    .Y(_0326_),
    .A1(_0171_),
    .A2(net179));
 sg13g2_nor2_1 _0871_ (.A(_0323_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_mux2_1 _0872_ (.A0(_0207_),
    .A1(_0224_),
    .S(net179),
    .X(_0328_));
 sg13g2_o21ai_1 _0873_ (.B1(_0277_),
    .Y(_0329_),
    .A1(_0249_),
    .A2(net180));
 sg13g2_mux2_1 _0874_ (.A0(_0329_),
    .A1(_0328_),
    .S(net183),
    .X(_0330_));
 sg13g2_nor2_1 _0875_ (.A(net186),
    .B(_0330_),
    .Y(_0331_));
 sg13g2_o21ai_1 _0876_ (.B1(_0321_),
    .Y(_0332_),
    .A1(_0327_),
    .A2(_0331_));
 sg13g2_nor2_2 _0877_ (.A(_0134_),
    .B(net179),
    .Y(_0333_));
 sg13g2_inv_1 _0878_ (.Y(_0334_),
    .A(_0333_));
 sg13g2_and2_1 _0879_ (.A(_0152_),
    .B(net178),
    .X(_0335_));
 sg13g2_and2_1 _0880_ (.A(net184),
    .B(net181),
    .X(_0336_));
 sg13g2_nand2_1 _0881_ (.Y(_0337_),
    .A(net184),
    .B(net182));
 sg13g2_a22oi_1 _0882_ (.Y(_0338_),
    .B1(_0335_),
    .B2(_0321_),
    .A2(_0333_),
    .A1(_0320_));
 sg13g2_nor2_1 _0883_ (.A(_0337_),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_nor3_1 _0884_ (.A(net212),
    .B(_0091_),
    .C(_0316_),
    .Y(_0340_));
 sg13g2_nor3_1 _0885_ (.A(_0134_),
    .B(_0311_),
    .C(_0319_),
    .Y(_0341_));
 sg13g2_nor3_1 _0886_ (.A(_0339_),
    .B(net189),
    .C(_0341_),
    .Y(_0342_));
 sg13g2_a221oi_1 _0887_ (.B2(_0332_),
    .C1(_0296_),
    .B1(_0342_),
    .A1(_0139_),
    .Y(_0343_),
    .A2(net189));
 sg13g2_a221oi_1 _0888_ (.B2(_0092_),
    .C1(_0343_),
    .B1(_0315_),
    .A1(_0312_),
    .Y(_0344_),
    .A2(_0314_));
 sg13g2_a221oi_1 _0889_ (.B2(_0297_),
    .C1(_0093_),
    .B1(_0344_),
    .A1(_0137_),
    .Y(_0345_),
    .A2(_0317_));
 sg13g2_a21oi_1 _0890_ (.A1(net191),
    .A2(_0136_),
    .Y(_0346_),
    .B1(_0345_));
 sg13g2_xor2_1 _0891_ (.B(_0309_),
    .A(_0158_),
    .X(_0347_));
 sg13g2_nor2_1 _0892_ (.A(_0313_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_xnor2_1 _0893_ (.Y(_0349_),
    .A(_0158_),
    .B(_0289_));
 sg13g2_nor2_1 _0894_ (.A(net180),
    .B(_0276_),
    .Y(_0350_));
 sg13g2_nor2_1 _0895_ (.A(net182),
    .B(_0350_),
    .Y(_0351_));
 sg13g2_nor2_1 _0896_ (.A(_0224_),
    .B(net178),
    .Y(_0352_));
 sg13g2_a21oi_1 _0897_ (.A1(_0255_),
    .A2(_0264_),
    .Y(_0353_),
    .B1(_0250_));
 sg13g2_nor2_1 _0898_ (.A(_0352_),
    .B(_0353_),
    .Y(_0354_));
 sg13g2_a21oi_1 _0899_ (.A1(net182),
    .A2(_0354_),
    .Y(_0355_),
    .B1(_0351_));
 sg13g2_and2_1 _0900_ (.A(_0218_),
    .B(_0355_),
    .X(_0356_));
 sg13g2_nand2_1 _0901_ (.Y(_0357_),
    .A(_0152_),
    .B(_0266_));
 sg13g2_o21ai_1 _0902_ (.B1(_0357_),
    .Y(_0358_),
    .A1(_0172_),
    .A2(_0266_));
 sg13g2_nand2_1 _0903_ (.Y(_0359_),
    .A(_0336_),
    .B(_0358_));
 sg13g2_nor2_1 _0904_ (.A(net187),
    .B(net178),
    .Y(_0360_));
 sg13g2_a21oi_1 _0905_ (.A1(_0206_),
    .A2(net178),
    .Y(_0361_),
    .B1(_0360_));
 sg13g2_o21ai_1 _0906_ (.B1(_0359_),
    .Y(_0362_),
    .A1(_0323_),
    .A2(_0361_));
 sg13g2_o21ai_1 _0907_ (.B1(_0321_),
    .Y(_0363_),
    .A1(_0356_),
    .A2(_0362_));
 sg13g2_a21oi_2 _0908_ (.B1(_0319_),
    .Y(_0364_),
    .A2(_0316_),
    .A1(_0311_));
 sg13g2_a21o_2 _0909_ (.A2(_0320_),
    .A1(net215),
    .B1(_0134_),
    .X(_0365_));
 sg13g2_inv_1 _0910_ (.Y(_0366_),
    .A(_0365_));
 sg13g2_mux2_1 _0911_ (.A0(_0135_),
    .A1(_0152_),
    .S(_0266_),
    .X(_0367_));
 sg13g2_nand3_1 _0912_ (.B(net181),
    .C(_0367_),
    .A(net185),
    .Y(_0368_));
 sg13g2_o21ai_1 _0913_ (.B1(_0368_),
    .Y(_0369_),
    .A1(_0336_),
    .A2(_0365_));
 sg13g2_a21oi_1 _0914_ (.A1(_0364_),
    .A2(_0369_),
    .Y(_0370_),
    .B1(net188));
 sg13g2_nand2_1 _0915_ (.Y(_0371_),
    .A(_0363_),
    .B(_0370_));
 sg13g2_nand3_1 _0916_ (.B(_0157_),
    .C(net189),
    .A(_0154_),
    .Y(_0372_));
 sg13g2_a221oi_1 _0917_ (.B2(_0372_),
    .C1(_0312_),
    .B1(_0371_),
    .A1(_0296_),
    .Y(_0373_),
    .A2(_0349_));
 sg13g2_o21ai_1 _0918_ (.B1(_0318_),
    .Y(_0374_),
    .A1(_0348_),
    .A2(_0373_));
 sg13g2_nand3_1 _0919_ (.B(_0153_),
    .C(net190),
    .A(_0146_),
    .Y(_0375_));
 sg13g2_a22oi_1 _0920_ (.Y(_0376_),
    .B1(_0374_),
    .B2(_0375_),
    .A2(_0155_),
    .A1(net191));
 sg13g2_a21oi_1 _0921_ (.A1(_0171_),
    .A2(_0266_),
    .Y(_0377_),
    .B1(_0335_));
 sg13g2_nor2_1 _0922_ (.A(net182),
    .B(_0333_),
    .Y(_0378_));
 sg13g2_a21oi_1 _0923_ (.A1(net181),
    .A2(_0377_),
    .Y(_0379_),
    .B1(_0378_));
 sg13g2_nand2_1 _0924_ (.Y(_0380_),
    .A(net184),
    .B(_0379_));
 sg13g2_o21ai_1 _0925_ (.B1(_0380_),
    .Y(_0381_),
    .A1(_0336_),
    .A2(_0365_));
 sg13g2_o21ai_1 _0926_ (.B1(net189),
    .Y(_0382_),
    .A1(_0174_),
    .A2(_0176_));
 sg13g2_nor2b_1 _0927_ (.A(_0329_),
    .B_N(net183),
    .Y(_0383_));
 sg13g2_or2_1 _0928_ (.X(_0384_),
    .B(_0328_),
    .A(_0323_));
 sg13g2_o21ai_1 _0929_ (.B1(_0384_),
    .Y(_0385_),
    .A1(_0326_),
    .A2(_0337_));
 sg13g2_a21oi_1 _0930_ (.A1(_0218_),
    .A2(_0383_),
    .Y(_0386_),
    .B1(_0385_));
 sg13g2_nor2_1 _0931_ (.A(_0322_),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_a221oi_1 _0932_ (.B2(_0381_),
    .C1(_0387_),
    .B1(_0364_),
    .A1(net214),
    .Y(_0388_),
    .A2(_0293_));
 sg13g2_xor2_1 _0933_ (.B(_0299_),
    .A(_0287_),
    .X(_0389_));
 sg13g2_a22oi_1 _0934_ (.Y(_0390_),
    .B1(_0389_),
    .B2(_0296_),
    .A2(_0388_),
    .A1(_0382_));
 sg13g2_xnor2_1 _0935_ (.Y(_0391_),
    .A(_0299_),
    .B(_0308_));
 sg13g2_o21ai_1 _0936_ (.B1(_0318_),
    .Y(_0392_),
    .A1(_0313_),
    .A2(_0391_));
 sg13g2_nand3_1 _0937_ (.B(_0172_),
    .C(net190),
    .A(_0165_),
    .Y(_0393_));
 sg13g2_o21ai_1 _0938_ (.B1(_0393_),
    .Y(_0394_),
    .A1(_0390_),
    .A2(_0392_));
 sg13g2_o21ai_1 _0939_ (.B1(_0394_),
    .Y(_0395_),
    .A1(_0094_),
    .A2(_0298_));
 sg13g2_nor2b_1 _0940_ (.A(_0138_),
    .B_N(_0154_),
    .Y(_0396_));
 sg13g2_nand2_1 _0941_ (.Y(_0397_),
    .A(_0229_),
    .B(_0306_));
 sg13g2_nand2_1 _0942_ (.Y(_0398_),
    .A(net182),
    .B(_0350_));
 sg13g2_a21oi_1 _0943_ (.A1(_0250_),
    .A2(_0398_),
    .Y(_0399_),
    .B1(_0351_));
 sg13g2_o21ai_1 _0944_ (.B1(_0208_),
    .Y(_0400_),
    .A1(_0209_),
    .A2(_0228_));
 sg13g2_o21ai_1 _0945_ (.B1(_0400_),
    .Y(_0401_),
    .A1(_0397_),
    .A2(_0399_));
 sg13g2_nand3_1 _0946_ (.B(_0299_),
    .C(_0401_),
    .A(_0285_),
    .Y(_0402_));
 sg13g2_nand3_1 _0947_ (.B(_0183_),
    .C(net187),
    .A(_0173_),
    .Y(_0403_));
 sg13g2_nand4_1 _0948_ (.B(_0175_),
    .C(_0402_),
    .A(_0157_),
    .Y(_0404_),
    .D(_0403_));
 sg13g2_a22oi_1 _0949_ (.Y(_0405_),
    .B1(_0396_),
    .B2(_0404_),
    .A2(_0135_),
    .A1(_0115_));
 sg13g2_nor2b_1 _0950_ (.A(net180),
    .B_N(_0276_),
    .Y(_0406_));
 sg13g2_o21ai_1 _0951_ (.B1(_0396_),
    .Y(_0407_),
    .A1(_0302_),
    .A2(_0406_));
 sg13g2_nand4_1 _0952_ (.B(_0285_),
    .C(_0299_),
    .A(_0229_),
    .Y(_0408_),
    .D(_0306_));
 sg13g2_nor4_1 _0953_ (.A(_0156_),
    .B(_0253_),
    .C(_0407_),
    .D(_0408_),
    .Y(_0409_));
 sg13g2_nor4_1 _0954_ (.A(_0295_),
    .B(_0319_),
    .C(_0405_),
    .D(_0409_),
    .Y(_0410_));
 sg13g2_nor2_1 _0955_ (.A(_0218_),
    .B(_0322_),
    .Y(_0411_));
 sg13g2_nand2_1 _0956_ (.Y(_0412_),
    .A(net185),
    .B(_0321_));
 sg13g2_a21o_1 _0957_ (.A2(net178),
    .A1(_0171_),
    .B1(_0360_),
    .X(_0413_));
 sg13g2_mux2_1 _0958_ (.A0(_0367_),
    .A1(_0413_),
    .S(net181),
    .X(_0414_));
 sg13g2_nor3_1 _0959_ (.A(_0337_),
    .B(_0350_),
    .C(_0353_),
    .Y(_0415_));
 sg13g2_a21o_1 _0960_ (.A2(net178),
    .A1(_0206_),
    .B1(_0352_),
    .X(_0416_));
 sg13g2_o21ai_1 _0961_ (.B1(_0364_),
    .Y(_0417_),
    .A1(_0323_),
    .A2(_0416_));
 sg13g2_nor2_1 _0962_ (.A(_0415_),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_o21ai_1 _0963_ (.B1(_0418_),
    .Y(_0419_),
    .A1(net185),
    .A2(_0414_));
 sg13g2_o21ai_1 _0964_ (.B1(_0419_),
    .Y(_0420_),
    .A1(_0398_),
    .A2(_0412_));
 sg13g2_nor2_1 _0965_ (.A(_0293_),
    .B(net188),
    .Y(_0421_));
 sg13g2_nor3_1 _0966_ (.A(_0302_),
    .B(_0406_),
    .C(_0421_),
    .Y(_0422_));
 sg13g2_or4_1 _0967_ (.A(net190),
    .B(_0410_),
    .C(_0420_),
    .D(_0422_),
    .X(_0423_));
 sg13g2_a21oi_1 _0968_ (.A1(net190),
    .A2(_0406_),
    .Y(_0424_),
    .B1(net191));
 sg13g2_a22oi_1 _0969_ (.Y(_0425_),
    .B1(_0423_),
    .B2(_0424_),
    .A2(_0302_),
    .A1(net191));
 sg13g2_nor2_1 _0970_ (.A(net214),
    .B(_0307_),
    .Y(_0426_));
 sg13g2_a21oi_1 _0971_ (.A1(net214),
    .A2(_0281_),
    .Y(_0427_),
    .B1(_0426_));
 sg13g2_o21ai_1 _0972_ (.B1(_0293_),
    .Y(_0428_),
    .A1(_0286_),
    .A2(_0427_));
 sg13g2_a21oi_1 _0973_ (.A1(_0286_),
    .A2(_0427_),
    .Y(_0429_),
    .B1(_0428_));
 sg13g2_a22oi_1 _0974_ (.Y(_0430_),
    .B1(_0284_),
    .B2(net190),
    .A2(_0283_),
    .A1(net191));
 sg13g2_nor2_1 _0975_ (.A(net184),
    .B(_0365_),
    .Y(_0431_));
 sg13g2_inv_1 _0976_ (.Y(_0432_),
    .A(_0431_));
 sg13g2_a21o_1 _0977_ (.A2(_0414_),
    .A1(net185),
    .B1(_0431_),
    .X(_0433_));
 sg13g2_nand2b_1 _0978_ (.Y(_0434_),
    .B(_0354_),
    .A_N(net181));
 sg13g2_nand2_1 _0979_ (.Y(_0435_),
    .A(net184),
    .B(_0434_));
 sg13g2_a221oi_1 _0980_ (.B2(_0435_),
    .C1(_0322_),
    .B1(_0398_),
    .A1(_0336_),
    .Y(_0436_),
    .A2(_0361_));
 sg13g2_a221oi_1 _0981_ (.B2(_0433_),
    .C1(_0436_),
    .B1(_0364_),
    .A1(_0286_),
    .Y(_0437_),
    .A2(net188));
 sg13g2_nand2_1 _0982_ (.Y(_0438_),
    .A(_0430_),
    .B(_0437_));
 sg13g2_nor2_1 _0983_ (.A(_0429_),
    .B(_0438_),
    .Y(_0439_));
 sg13g2_mux2_1 _0984_ (.A0(_0207_),
    .A1(net187),
    .S(net179),
    .X(_0440_));
 sg13g2_a21oi_1 _0985_ (.A1(net181),
    .A2(_0333_),
    .Y(_0441_),
    .B1(net184));
 sg13g2_a221oi_1 _0986_ (.B2(_0336_),
    .C1(_0441_),
    .B1(_0440_),
    .A1(_0324_),
    .Y(_0442_),
    .A2(_0377_));
 sg13g2_o21ai_1 _0987_ (.B1(_0364_),
    .Y(_0443_),
    .A1(_0431_),
    .A2(_0442_));
 sg13g2_nand2b_1 _0988_ (.Y(_0444_),
    .B(net188),
    .A_N(_0306_));
 sg13g2_o21ai_1 _0989_ (.B1(_0444_),
    .Y(_0445_),
    .A1(_0330_),
    .A2(_0412_));
 sg13g2_nor2_1 _0990_ (.A(_0296_),
    .B(_0445_),
    .Y(_0446_));
 sg13g2_xor2_1 _0991_ (.B(_0306_),
    .A(_0280_),
    .X(_0447_));
 sg13g2_a22oi_1 _0992_ (.Y(_0448_),
    .B1(_0447_),
    .B2(_0296_),
    .A2(_0446_),
    .A1(_0443_));
 sg13g2_nor2_1 _0993_ (.A(_0312_),
    .B(_0448_),
    .Y(_0449_));
 sg13g2_xnor2_1 _0994_ (.Y(_0450_),
    .A(_0304_),
    .B(_0306_));
 sg13g2_a21oi_1 _0995_ (.A1(_0312_),
    .A2(_0450_),
    .Y(_0451_),
    .B1(_0449_));
 sg13g2_a221oi_1 _0996_ (.B2(net190),
    .C1(_0451_),
    .B1(_0305_),
    .A1(net191),
    .Y(_0452_),
    .A2(_0300_));
 sg13g2_mux4_1 _0997_ (.S0(net181),
    .A0(_0366_),
    .A1(_0367_),
    .A2(_0413_),
    .A3(_0416_),
    .S1(net185),
    .X(_0453_));
 sg13g2_a221oi_1 _0998_ (.B2(_0364_),
    .C1(net188),
    .B1(_0453_),
    .A1(_0355_),
    .Y(_0454_),
    .A2(_0411_));
 sg13g2_a21oi_1 _0999_ (.A1(_0229_),
    .A2(net188),
    .Y(_0455_),
    .B1(_0454_));
 sg13g2_xnor2_1 _1000_ (.Y(_0456_),
    .A(_0229_),
    .B(_0279_));
 sg13g2_a21oi_1 _1001_ (.A1(net214),
    .A2(_0456_),
    .Y(_0457_),
    .B1(_0294_));
 sg13g2_nor2_1 _1002_ (.A(_0455_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_xnor2_1 _1003_ (.Y(_0459_),
    .A(_0229_),
    .B(_0303_));
 sg13g2_o21ai_1 _1004_ (.B1(_0318_),
    .Y(_0460_),
    .A1(_0313_),
    .A2(_0459_));
 sg13g2_a21oi_1 _1005_ (.A1(_0227_),
    .A2(net190),
    .Y(_0461_),
    .B1(net191));
 sg13g2_o21ai_1 _1006_ (.B1(_0461_),
    .Y(_0462_),
    .A1(_0458_),
    .A2(_0460_));
 sg13g2_o21ai_1 _1007_ (.B1(_0462_),
    .Y(_0463_),
    .A1(_0094_),
    .A2(_0226_));
 sg13g2_mux2_1 _1008_ (.A0(_0250_),
    .A1(_0224_),
    .S(net178),
    .X(_0464_));
 sg13g2_mux4_1 _1009_ (.S0(net181),
    .A0(_0334_),
    .A1(_0377_),
    .A2(_0440_),
    .A3(_0464_),
    .S1(net184),
    .X(_0465_));
 sg13g2_o21ai_1 _1010_ (.B1(_0465_),
    .Y(_0466_),
    .A1(net182),
    .A2(_0432_));
 sg13g2_a221oi_1 _1011_ (.B2(_0364_),
    .C1(net188),
    .B1(_0466_),
    .A1(_0383_),
    .Y(_0467_),
    .A2(_0411_));
 sg13g2_a21o_1 _1012_ (.A2(net188),
    .A1(_0254_),
    .B1(_0467_),
    .X(_0468_));
 sg13g2_xnor2_1 _1013_ (.Y(_0469_),
    .A(_0253_),
    .B(_0277_));
 sg13g2_a21oi_1 _1014_ (.A1(_0253_),
    .A2(_0302_),
    .Y(_0470_),
    .B1(_0313_));
 sg13g2_o21ai_1 _1015_ (.B1(_0470_),
    .Y(_0471_),
    .A1(_0253_),
    .A2(_0302_));
 sg13g2_a221oi_1 _1016_ (.B2(_0296_),
    .C1(net191),
    .B1(_0469_),
    .A1(_0252_),
    .Y(_0472_),
    .A2(net190));
 sg13g2_nand3_1 _1017_ (.B(_0471_),
    .C(_0472_),
    .A(_0468_),
    .Y(_0473_));
 sg13g2_o21ai_1 _1018_ (.B1(_0473_),
    .Y(_0474_),
    .A1(_0094_),
    .A2(_0251_));
 sg13g2_nand4_1 _1019_ (.B(_0452_),
    .C(_0463_),
    .A(_0439_),
    .Y(_0475_),
    .D(_0474_));
 sg13g2_nor2_1 _1020_ (.A(_0395_),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_nand4_1 _1021_ (.B(_0376_),
    .C(_0425_),
    .A(_0346_),
    .Y(_0477_),
    .D(_0476_));
 sg13g2_nand2_2 _1022_ (.Y(_0478_),
    .A(net1),
    .B(net2));
 sg13g2_nor3_1 _1023_ (.A(net212),
    .B(_0295_),
    .C(_0478_),
    .Y(_0479_));
 sg13g2_nand2_1 _1024_ (.Y(_0480_),
    .A(net212),
    .B(_0425_));
 sg13g2_nor3_1 _1025_ (.A(net11),
    .B(_0295_),
    .C(_0478_),
    .Y(_0481_));
 sg13g2_nor4_1 _1026_ (.A(net212),
    .B(net11),
    .C(_0295_),
    .D(_0478_),
    .Y(_0482_));
 sg13g2_a22oi_1 _1027_ (.Y(_0483_),
    .B1(_0480_),
    .B2(_0481_),
    .A2(_0479_),
    .A1(_0477_));
 sg13g2_or4_2 _1028_ (.A(net216),
    .B(net12),
    .C(net212),
    .D(_0478_),
    .X(_0484_));
 sg13g2_inv_1 _1029_ (.Y(_0485_),
    .A(_0484_));
 sg13g2_a21o_1 _1030_ (.A2(_0482_),
    .A1(_0477_),
    .B1(_0485_),
    .X(_0486_));
 sg13g2_nand2b_1 _1031_ (.Y(_0487_),
    .B(_0485_),
    .A_N(_0276_));
 sg13g2_o21ai_1 _1032_ (.B1(_0487_),
    .Y(uo_out[0]),
    .A1(_0483_),
    .A2(_0486_));
 sg13g2_nor2_1 _1033_ (.A(_0250_),
    .B(_0484_),
    .Y(uo_out[1]));
 sg13g2_nor2_1 _1034_ (.A(_0224_),
    .B(_0484_),
    .Y(uo_out[2]));
 sg13g2_nor2_1 _1035_ (.A(_0207_),
    .B(_0484_),
    .Y(uo_out[3]));
 sg13g2_nor2_2 _1036_ (.A(_0189_),
    .B(_0484_),
    .Y(uo_out[4]));
 sg13g2_nor2_2 _1037_ (.A(_0172_),
    .B(_0484_),
    .Y(uo_out[5]));
 sg13g2_nor2_2 _1038_ (.A(_0153_),
    .B(_0484_),
    .Y(uo_out[6]));
 sg13g2_nor2_1 _1039_ (.A(_0134_),
    .B(_0484_),
    .Y(uo_out[7]));
 sg13g2_nand4_1 _1040_ (.B(net3),
    .C(net5),
    .A(net4),
    .Y(_0488_),
    .D(_0478_));
 sg13g2_nand2b_1 _1041_ (.Y(_0489_),
    .B(net2),
    .A_N(net1));
 sg13g2_nand2_1 _1042_ (.Y(_0490_),
    .A(_0425_),
    .B(net207));
 sg13g2_o21ai_1 _1043_ (.B1(_0490_),
    .Y(_0491_),
    .A1(net221),
    .A2(net207));
 sg13g2_nand2_1 _1044_ (.Y(_0492_),
    .A(net38),
    .B(net205));
 sg13g2_o21ai_1 _1045_ (.B1(_0492_),
    .Y(_0010_),
    .A1(net205),
    .A2(_0491_));
 sg13g2_nand2_1 _1046_ (.Y(_0493_),
    .A(_0474_),
    .B(net207));
 sg13g2_o21ai_1 _1047_ (.B1(_0493_),
    .Y(_0494_),
    .A1(net218),
    .A2(net207));
 sg13g2_nand2_1 _1048_ (.Y(_0495_),
    .A(net53),
    .B(net205));
 sg13g2_o21ai_1 _1049_ (.B1(_0495_),
    .Y(_0011_),
    .A1(net205),
    .A2(_0494_));
 sg13g2_nand2_1 _1050_ (.Y(_0496_),
    .A(_0463_),
    .B(net206));
 sg13g2_o21ai_1 _1051_ (.B1(_0496_),
    .Y(_0497_),
    .A1(net217),
    .A2(net207));
 sg13g2_nand2_1 _1052_ (.Y(_0498_),
    .A(net39),
    .B(net205));
 sg13g2_o21ai_1 _1053_ (.B1(_0498_),
    .Y(_0012_),
    .A1(net204),
    .A2(_0497_));
 sg13g2_nand2_1 _1054_ (.Y(_0499_),
    .A(_0452_),
    .B(net206));
 sg13g2_o21ai_1 _1055_ (.B1(_0499_),
    .Y(_0500_),
    .A1(net10),
    .A2(net206));
 sg13g2_nand2_1 _1056_ (.Y(_0501_),
    .A(net47),
    .B(net204));
 sg13g2_o21ai_1 _1057_ (.B1(_0501_),
    .Y(_0013_),
    .A1(net204),
    .A2(_0500_));
 sg13g2_nand2_1 _1058_ (.Y(_0502_),
    .A(_0439_),
    .B(net206));
 sg13g2_o21ai_1 _1059_ (.B1(_0502_),
    .Y(_0503_),
    .A1(net11),
    .A2(net207));
 sg13g2_nand2_1 _1060_ (.Y(_0504_),
    .A(net63),
    .B(net205));
 sg13g2_o21ai_1 _1061_ (.B1(_0504_),
    .Y(_0014_),
    .A1(net205),
    .A2(_0503_));
 sg13g2_mux2_2 _1062_ (.A0(net216),
    .A1(_0395_),
    .S(net206),
    .X(_0505_));
 sg13g2_mux2_1 _1063_ (.A0(_0505_),
    .A1(net93),
    .S(net204),
    .X(_0015_));
 sg13g2_nand2_1 _1064_ (.Y(_0506_),
    .A(_0376_),
    .B(net206));
 sg13g2_o21ai_1 _1065_ (.B1(_0506_),
    .Y(_0507_),
    .A1(net213),
    .A2(net206));
 sg13g2_nand2_1 _1066_ (.Y(_0508_),
    .A(net59),
    .B(net204));
 sg13g2_o21ai_1 _1067_ (.B1(_0508_),
    .Y(_0016_),
    .A1(net204),
    .A2(_0507_));
 sg13g2_nand2_1 _1068_ (.Y(_0509_),
    .A(_0346_),
    .B(net206));
 sg13g2_o21ai_1 _1069_ (.B1(_0509_),
    .Y(_0510_),
    .A1(net13),
    .A2(net207));
 sg13g2_nand2_1 _1070_ (.Y(_0511_),
    .A(net60),
    .B(net204));
 sg13g2_o21ai_1 _1071_ (.B1(_0511_),
    .Y(_0017_),
    .A1(net204),
    .A2(_0510_));
 sg13g2_nor2b_1 _1072_ (.A(net3),
    .B_N(net4),
    .Y(_0512_));
 sg13g2_nand3_1 _1073_ (.B(_0478_),
    .C(_0512_),
    .A(net5),
    .Y(_0513_));
 sg13g2_nand2_1 _1074_ (.Y(_0514_),
    .A(net84),
    .B(net203));
 sg13g2_o21ai_1 _1075_ (.B1(_0514_),
    .Y(_0018_),
    .A1(_0491_),
    .A2(net203));
 sg13g2_nand2_1 _1076_ (.Y(_0515_),
    .A(net42),
    .B(net203));
 sg13g2_o21ai_1 _1077_ (.B1(_0515_),
    .Y(_0019_),
    .A1(_0494_),
    .A2(net203));
 sg13g2_nand2_1 _1078_ (.Y(_0516_),
    .A(net64),
    .B(net203));
 sg13g2_o21ai_1 _1079_ (.B1(_0516_),
    .Y(_0020_),
    .A1(_0497_),
    .A2(net203));
 sg13g2_nand2_1 _1080_ (.Y(_0517_),
    .A(net50),
    .B(net202));
 sg13g2_o21ai_1 _1081_ (.B1(_0517_),
    .Y(_0021_),
    .A1(_0500_),
    .A2(net202));
 sg13g2_nand2_1 _1082_ (.Y(_0518_),
    .A(net66),
    .B(net202));
 sg13g2_o21ai_1 _1083_ (.B1(_0518_),
    .Y(_0022_),
    .A1(_0503_),
    .A2(net203));
 sg13g2_mux2_1 _1084_ (.A0(_0505_),
    .A1(net89),
    .S(net202),
    .X(_0023_));
 sg13g2_nand2_1 _1085_ (.Y(_0519_),
    .A(net56),
    .B(net202));
 sg13g2_o21ai_1 _1086_ (.B1(_0519_),
    .Y(_0024_),
    .A1(_0507_),
    .A2(net202));
 sg13g2_nand2_1 _1087_ (.Y(_0520_),
    .A(net72),
    .B(net202));
 sg13g2_o21ai_1 _1088_ (.B1(_0520_),
    .Y(_0025_),
    .A1(_0510_),
    .A2(net202));
 sg13g2_nor2_1 _1089_ (.A(net4),
    .B(net3),
    .Y(_0521_));
 sg13g2_nand3_1 _1090_ (.B(_0478_),
    .C(_0521_),
    .A(net5),
    .Y(_0522_));
 sg13g2_nand2_1 _1091_ (.Y(_0523_),
    .A(net82),
    .B(net201));
 sg13g2_o21ai_1 _1092_ (.B1(_0523_),
    .Y(_0026_),
    .A1(_0491_),
    .A2(net201));
 sg13g2_nand2_1 _1093_ (.Y(_0524_),
    .A(net51),
    .B(net201));
 sg13g2_o21ai_1 _1094_ (.B1(_0524_),
    .Y(_0027_),
    .A1(_0494_),
    .A2(net201));
 sg13g2_nand2_1 _1095_ (.Y(_0525_),
    .A(net49),
    .B(net200));
 sg13g2_o21ai_1 _1096_ (.B1(_0525_),
    .Y(_0028_),
    .A1(_0497_),
    .A2(net201));
 sg13g2_nand2_1 _1097_ (.Y(_0526_),
    .A(net61),
    .B(net200));
 sg13g2_o21ai_1 _1098_ (.B1(_0526_),
    .Y(_0029_),
    .A1(_0500_),
    .A2(net200));
 sg13g2_nand2_1 _1099_ (.Y(_0527_),
    .A(net70),
    .B(net201));
 sg13g2_o21ai_1 _1100_ (.B1(_0527_),
    .Y(_0030_),
    .A1(_0503_),
    .A2(net201));
 sg13g2_mux2_1 _1101_ (.A0(_0505_),
    .A1(net88),
    .S(net200),
    .X(_0031_));
 sg13g2_nand2_1 _1102_ (.Y(_0528_),
    .A(net48),
    .B(net200));
 sg13g2_o21ai_1 _1103_ (.B1(_0528_),
    .Y(_0032_),
    .A1(_0507_),
    .A2(net200));
 sg13g2_nand2_1 _1104_ (.Y(_0529_),
    .A(net46),
    .B(net200));
 sg13g2_o21ai_1 _1105_ (.B1(_0529_),
    .Y(_0033_),
    .A1(_0510_),
    .A2(net200));
 sg13g2_a21oi_1 _1106_ (.A1(net1),
    .A2(net2),
    .Y(_0530_),
    .B1(net5));
 sg13g2_nand3_1 _1107_ (.B(net3),
    .C(_0530_),
    .A(net4),
    .Y(_0531_));
 sg13g2_nand2_1 _1108_ (.Y(_0532_),
    .A(net44),
    .B(net198));
 sg13g2_o21ai_1 _1109_ (.B1(_0532_),
    .Y(_0034_),
    .A1(_0491_),
    .A2(net198));
 sg13g2_nand2_1 _1110_ (.Y(_0533_),
    .A(net40),
    .B(net198));
 sg13g2_o21ai_1 _1111_ (.B1(_0533_),
    .Y(_0035_),
    .A1(_0494_),
    .A2(net198));
 sg13g2_nand2_1 _1112_ (.Y(_0534_),
    .A(net77),
    .B(net198));
 sg13g2_o21ai_1 _1113_ (.B1(_0534_),
    .Y(_0036_),
    .A1(_0497_),
    .A2(net198));
 sg13g2_nand2_1 _1114_ (.Y(_0535_),
    .A(net58),
    .B(net199));
 sg13g2_o21ai_1 _1115_ (.B1(_0535_),
    .Y(_0037_),
    .A1(_0500_),
    .A2(net199));
 sg13g2_nand2_1 _1116_ (.Y(_0536_),
    .A(net80),
    .B(net199));
 sg13g2_o21ai_1 _1117_ (.B1(_0536_),
    .Y(_0038_),
    .A1(_0503_),
    .A2(net198));
 sg13g2_mux2_1 _1118_ (.A0(_0505_),
    .A1(net91),
    .S(net198),
    .X(_0039_));
 sg13g2_nand2_1 _1119_ (.Y(_0537_),
    .A(net74),
    .B(net199));
 sg13g2_o21ai_1 _1120_ (.B1(_0537_),
    .Y(_0040_),
    .A1(_0507_),
    .A2(net199));
 sg13g2_nand2_1 _1121_ (.Y(_0538_),
    .A(net43),
    .B(net199));
 sg13g2_o21ai_1 _1122_ (.B1(_0538_),
    .Y(_0041_),
    .A1(_0510_),
    .A2(net199));
 sg13g2_nand2_1 _1123_ (.Y(_0539_),
    .A(_0512_),
    .B(_0530_));
 sg13g2_nand2_1 _1124_ (.Y(_0540_),
    .A(net45),
    .B(net197));
 sg13g2_o21ai_1 _1125_ (.B1(_0540_),
    .Y(_0042_),
    .A1(_0491_),
    .A2(net197));
 sg13g2_nand2_1 _1126_ (.Y(_0541_),
    .A(net76),
    .B(net197));
 sg13g2_o21ai_1 _1127_ (.B1(_0541_),
    .Y(_0043_),
    .A1(_0494_),
    .A2(net197));
 sg13g2_nand2_1 _1128_ (.Y(_0542_),
    .A(net67),
    .B(net196));
 sg13g2_o21ai_1 _1129_ (.B1(_0542_),
    .Y(_0044_),
    .A1(_0497_),
    .A2(net197));
 sg13g2_nand2_1 _1130_ (.Y(_0543_),
    .A(net57),
    .B(net196));
 sg13g2_o21ai_1 _1131_ (.B1(_0543_),
    .Y(_0045_),
    .A1(_0500_),
    .A2(net196));
 sg13g2_nand2_1 _1132_ (.Y(_0544_),
    .A(net52),
    .B(net197));
 sg13g2_o21ai_1 _1133_ (.B1(_0544_),
    .Y(_0046_),
    .A1(_0503_),
    .A2(net197));
 sg13g2_mux2_1 _1134_ (.A0(_0505_),
    .A1(net86),
    .S(net196),
    .X(_0047_));
 sg13g2_nand2_1 _1135_ (.Y(_0545_),
    .A(net68),
    .B(net196));
 sg13g2_o21ai_1 _1136_ (.B1(_0545_),
    .Y(_0048_),
    .A1(_0507_),
    .A2(net196));
 sg13g2_nand2_1 _1137_ (.Y(_0546_),
    .A(net65),
    .B(net196));
 sg13g2_o21ai_1 _1138_ (.B1(_0546_),
    .Y(_0049_),
    .A1(_0510_),
    .A2(net196));
 sg13g2_nor2b_1 _1139_ (.A(net4),
    .B_N(net3),
    .Y(_0547_));
 sg13g2_nand2_1 _1140_ (.Y(_0548_),
    .A(_0530_),
    .B(_0547_));
 sg13g2_nand2_1 _1141_ (.Y(_0549_),
    .A(net85),
    .B(net195));
 sg13g2_o21ai_1 _1142_ (.B1(_0549_),
    .Y(_0050_),
    .A1(_0491_),
    .A2(net195));
 sg13g2_nand2_1 _1143_ (.Y(_0550_),
    .A(net79),
    .B(net194));
 sg13g2_o21ai_1 _1144_ (.B1(_0550_),
    .Y(_0051_),
    .A1(_0494_),
    .A2(net194));
 sg13g2_nand2_1 _1145_ (.Y(_0551_),
    .A(net62),
    .B(net195));
 sg13g2_o21ai_1 _1146_ (.B1(_0551_),
    .Y(_0052_),
    .A1(_0497_),
    .A2(net195));
 sg13g2_nand2_1 _1147_ (.Y(_0552_),
    .A(net54),
    .B(net194));
 sg13g2_o21ai_1 _1148_ (.B1(_0552_),
    .Y(_0053_),
    .A1(_0500_),
    .A2(net194));
 sg13g2_nand2_1 _1149_ (.Y(_0553_),
    .A(net81),
    .B(net195));
 sg13g2_o21ai_1 _1150_ (.B1(_0553_),
    .Y(_0054_),
    .A1(_0503_),
    .A2(net195));
 sg13g2_mux2_1 _1151_ (.A0(_0505_),
    .A1(net92),
    .S(net195),
    .X(_0055_));
 sg13g2_nand2_1 _1152_ (.Y(_0554_),
    .A(net69),
    .B(net194));
 sg13g2_o21ai_1 _1153_ (.B1(_0554_),
    .Y(_0056_),
    .A1(_0507_),
    .A2(net194));
 sg13g2_nand2_1 _1154_ (.Y(_0555_),
    .A(net75),
    .B(net194));
 sg13g2_o21ai_1 _1155_ (.B1(_0555_),
    .Y(_0057_),
    .A1(_0510_),
    .A2(net194));
 sg13g2_nand3_1 _1156_ (.B(_0478_),
    .C(_0547_),
    .A(net5),
    .Y(_0556_));
 sg13g2_nand2_1 _1157_ (.Y(_0557_),
    .A(net87),
    .B(net193));
 sg13g2_o21ai_1 _1158_ (.B1(_0557_),
    .Y(_0066_),
    .A1(_0491_),
    .A2(net193));
 sg13g2_nand2_1 _1159_ (.Y(_0558_),
    .A(net41),
    .B(net193));
 sg13g2_o21ai_1 _1160_ (.B1(_0558_),
    .Y(_0067_),
    .A1(_0494_),
    .A2(net193));
 sg13g2_nand2_1 _1161_ (.Y(_0559_),
    .A(net78),
    .B(net192));
 sg13g2_o21ai_1 _1162_ (.B1(_0559_),
    .Y(_0068_),
    .A1(_0497_),
    .A2(net192));
 sg13g2_nand2_1 _1163_ (.Y(_0560_),
    .A(net73),
    .B(net192));
 sg13g2_o21ai_1 _1164_ (.B1(_0560_),
    .Y(_0069_),
    .A1(_0500_),
    .A2(net192));
 sg13g2_nand2_1 _1165_ (.Y(_0561_),
    .A(net71),
    .B(net193));
 sg13g2_o21ai_1 _1166_ (.B1(_0561_),
    .Y(_0070_),
    .A1(_0503_),
    .A2(net193));
 sg13g2_mux2_1 _1167_ (.A0(_0505_),
    .A1(net90),
    .S(net193),
    .X(_0071_));
 sg13g2_nand2_1 _1168_ (.Y(_0562_),
    .A(net55),
    .B(net192));
 sg13g2_o21ai_1 _1169_ (.B1(_0562_),
    .Y(_0072_),
    .A1(_0507_),
    .A2(net192));
 sg13g2_nand2_1 _1170_ (.Y(_0563_),
    .A(net83),
    .B(net192));
 sg13g2_o21ai_1 _1171_ (.B1(_0563_),
    .Y(_0073_),
    .A1(_0510_),
    .A2(net192));
 sg13g2_buf_1 _1172_ (.A(net31),
    .X(_0058_));
 sg13g2_buf_1 _1173_ (.A(net35),
    .X(_0059_));
 sg13g2_buf_1 _1174_ (.A(net30),
    .X(_0060_));
 sg13g2_buf_1 _1175_ (.A(net37),
    .X(_0061_));
 sg13g2_buf_1 _1176_ (.A(net36),
    .X(_0062_));
 sg13g2_buf_1 _1177_ (.A(net32),
    .X(_0063_));
 sg13g2_buf_1 _1178_ (.A(net33),
    .X(_0064_));
 sg13g2_buf_1 _1179_ (.A(net34),
    .X(_0065_));
 sg13g2_dfrbp_1 _1180_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net232),
    .D(_0010_),
    .Q_N(_0001_),
    .Q(\reg_file.registers[7][0] ));
 sg13g2_dfrbp_1 _1181_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net228),
    .D(_0011_),
    .Q_N(_0617_),
    .Q(\reg_file.registers[7][1] ));
 sg13g2_dfrbp_1 _1182_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net230),
    .D(_0012_),
    .Q_N(_0003_),
    .Q(\reg_file.registers[7][2] ));
 sg13g2_dfrbp_1 _1183_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net225),
    .D(_0013_),
    .Q_N(_0616_),
    .Q(\reg_file.registers[7][3] ));
 sg13g2_dfrbp_1 _1184_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net232),
    .D(_0014_),
    .Q_N(_0615_),
    .Q(\reg_file.registers[7][4] ));
 sg13g2_dfrbp_1 _1185_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net229),
    .D(_0015_),
    .Q_N(_0614_),
    .Q(\reg_file.registers[7][5] ));
 sg13g2_dfrbp_1 _1186_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net225),
    .D(_0016_),
    .Q_N(_0613_),
    .Q(\reg_file.registers[7][6] ));
 sg13g2_dfrbp_1 _1187_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net231),
    .D(_0017_),
    .Q_N(_0612_),
    .Q(\reg_file.registers[7][7] ));
 sg13g2_dfrbp_1 _1188_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net232),
    .D(_0018_),
    .Q_N(_0611_),
    .Q(\reg_file.registers[6][0] ));
 sg13g2_dfrbp_1 _1189_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net234),
    .D(_0019_),
    .Q_N(_0610_),
    .Q(\reg_file.registers[6][1] ));
 sg13g2_dfrbp_1 _1190_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net230),
    .D(_0020_),
    .Q_N(_0609_),
    .Q(\reg_file.registers[6][2] ));
 sg13g2_dfrbp_1 _1191_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net226),
    .D(_0021_),
    .Q_N(_0608_),
    .Q(\reg_file.registers[6][3] ));
 sg13g2_dfrbp_1 _1192_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net234),
    .D(_0022_),
    .Q_N(_0607_),
    .Q(\reg_file.registers[6][4] ));
 sg13g2_dfrbp_1 _1193_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net229),
    .D(_0023_),
    .Q_N(_0606_),
    .Q(\reg_file.registers[6][5] ));
 sg13g2_dfrbp_1 _1194_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net225),
    .D(_0024_),
    .Q_N(_0605_),
    .Q(\reg_file.registers[6][6] ));
 sg13g2_dfrbp_1 _1195_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net231),
    .D(_0025_),
    .Q_N(_0604_),
    .Q(\reg_file.registers[6][7] ));
 sg13g2_dfrbp_1 _1196_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net233),
    .D(_0026_),
    .Q_N(_0603_),
    .Q(\reg_file.registers[4][0] ));
 sg13g2_dfrbp_1 _1197_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net228),
    .D(_0027_),
    .Q_N(_0602_),
    .Q(\reg_file.registers[4][1] ));
 sg13g2_dfrbp_1 _1198_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net231),
    .D(_0028_),
    .Q_N(_0601_),
    .Q(\reg_file.registers[4][2] ));
 sg13g2_dfrbp_1 _1199_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net235),
    .D(_0029_),
    .Q_N(_0600_),
    .Q(\reg_file.registers[4][3] ));
 sg13g2_dfrbp_1 _1200_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net232),
    .D(_0030_),
    .Q_N(_0599_),
    .Q(\reg_file.registers[4][4] ));
 sg13g2_dfrbp_1 _1201_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net229),
    .D(_0031_),
    .Q_N(_0598_),
    .Q(\reg_file.registers[4][5] ));
 sg13g2_dfrbp_1 _1202_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net226),
    .D(_0032_),
    .Q_N(_0597_),
    .Q(\reg_file.registers[4][6] ));
 sg13g2_dfrbp_1 _1203_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net231),
    .D(_0033_),
    .Q_N(_0596_),
    .Q(\reg_file.registers[4][7] ));
 sg13g2_dfrbp_1 _1204_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net233),
    .D(_0034_),
    .Q_N(_0595_),
    .Q(\reg_file.registers[3][0] ));
 sg13g2_dfrbp_1 _1205_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net233),
    .D(_0035_),
    .Q_N(_0594_),
    .Q(\reg_file.registers[3][1] ));
 sg13g2_dfrbp_1 _1206_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net229),
    .D(_0036_),
    .Q_N(_0593_),
    .Q(\reg_file.registers[3][2] ));
 sg13g2_dfrbp_1 _1207_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net227),
    .D(_0037_),
    .Q_N(_0592_),
    .Q(\reg_file.registers[3][3] ));
 sg13g2_dfrbp_1 _1208_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net233),
    .D(_0038_),
    .Q_N(_0591_),
    .Q(\reg_file.registers[3][4] ));
 sg13g2_dfrbp_1 _1209_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net229),
    .D(_0039_),
    .Q_N(_0590_),
    .Q(\reg_file.registers[3][5] ));
 sg13g2_dfrbp_1 _1210_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net227),
    .D(_0040_),
    .Q_N(_0589_),
    .Q(\reg_file.registers[3][6] ));
 sg13g2_dfrbp_1 _1211_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net225),
    .D(_0041_),
    .Q_N(_0588_),
    .Q(\reg_file.registers[3][7] ));
 sg13g2_dfrbp_1 _1212_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net233),
    .D(_0042_),
    .Q_N(_0587_),
    .Q(\reg_file.registers[2][0] ));
 sg13g2_dfrbp_1 _1213_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net234),
    .D(_0043_),
    .Q_N(_0586_),
    .Q(\reg_file.registers[2][1] ));
 sg13g2_dfrbp_1 _1214_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net230),
    .D(_0044_),
    .Q_N(_0585_),
    .Q(\reg_file.registers[2][2] ));
 sg13g2_dfrbp_1 _1215_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net226),
    .D(_0045_),
    .Q_N(_0584_),
    .Q(\reg_file.registers[2][3] ));
 sg13g2_dfrbp_1 _1216_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net232),
    .D(_0046_),
    .Q_N(_0583_),
    .Q(\reg_file.registers[2][4] ));
 sg13g2_dfrbp_1 _1217_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net231),
    .D(_0047_),
    .Q_N(_0582_),
    .Q(\reg_file.registers[2][5] ));
 sg13g2_dfrbp_1 _1218_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net225),
    .D(_0048_),
    .Q_N(_0581_),
    .Q(\reg_file.registers[2][6] ));
 sg13g2_dfrbp_1 _1219_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net225),
    .D(_0049_),
    .Q_N(_0580_),
    .Q(\reg_file.registers[2][7] ));
 sg13g2_dfrbp_1 _1220_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net232),
    .D(_0050_),
    .Q_N(_0579_),
    .Q(\reg_file.registers[1][0] ));
 sg13g2_dfrbp_1 _1221_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net228),
    .D(_0051_),
    .Q_N(_0578_),
    .Q(\reg_file.registers[1][1] ));
 sg13g2_dfrbp_1 _1222_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net230),
    .D(_0052_),
    .Q_N(_0577_),
    .Q(\reg_file.registers[1][2] ));
 sg13g2_dfrbp_1 _1223_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net228),
    .D(_0053_),
    .Q_N(_0576_),
    .Q(\reg_file.registers[1][3] ));
 sg13g2_dfrbp_1 _1224_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net232),
    .D(_0054_),
    .Q_N(_0575_),
    .Q(\reg_file.registers[1][4] ));
 sg13g2_dfrbp_1 _1225_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net229),
    .D(_0055_),
    .Q_N(_0574_),
    .Q(\reg_file.registers[1][5] ));
 sg13g2_dfrbp_1 _1226_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net225),
    .D(_0056_),
    .Q_N(_0573_),
    .Q(\reg_file.registers[1][6] ));
 sg13g2_dfrbp_1 _1227_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net231),
    .D(_0057_),
    .Q_N(_0572_),
    .Q(\reg_file.registers[1][7] ));
 sg13g2_dfrbp_1 _1228_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net228),
    .D(_0058_),
    .Q_N(_0000_),
    .Q(\reg_file.registers[0][0] ));
 sg13g2_dfrbp_1 _1229_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net228),
    .D(_0059_),
    .Q_N(_0004_),
    .Q(\reg_file.registers[0][1] ));
 sg13g2_dfrbp_1 _1230_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net227),
    .D(_0060_),
    .Q_N(_0002_),
    .Q(\reg_file.registers[0][2] ));
 sg13g2_dfrbp_1 _1231_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net227),
    .D(_0061_),
    .Q_N(_0009_),
    .Q(\reg_file.registers[0][3] ));
 sg13g2_dfrbp_1 _1232_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net234),
    .D(_0062_),
    .Q_N(_0008_),
    .Q(\reg_file.registers[0][4] ));
 sg13g2_dfrbp_1 _1233_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net227),
    .D(_0063_),
    .Q_N(_0007_),
    .Q(\reg_file.registers[0][5] ));
 sg13g2_dfrbp_1 _1234_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net227),
    .D(_0064_),
    .Q_N(_0006_),
    .Q(\reg_file.registers[0][6] ));
 sg13g2_dfrbp_1 _1235_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net227),
    .D(_0065_),
    .Q_N(_0005_),
    .Q(\reg_file.registers[0][7] ));
 sg13g2_dfrbp_1 _1236_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net233),
    .D(_0066_),
    .Q_N(_0571_),
    .Q(\reg_file.registers[5][0] ));
 sg13g2_dfrbp_1 _1237_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net233),
    .D(_0067_),
    .Q_N(_0570_),
    .Q(\reg_file.registers[5][1] ));
 sg13g2_dfrbp_1 _1238_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net229),
    .D(_0068_),
    .Q_N(_0569_),
    .Q(\reg_file.registers[5][2] ));
 sg13g2_dfrbp_1 _1239_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net226),
    .D(_0069_),
    .Q_N(_0568_),
    .Q(\reg_file.registers[5][3] ));
 sg13g2_dfrbp_1 _1240_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net232),
    .D(_0070_),
    .Q_N(_0567_),
    .Q(\reg_file.registers[5][4] ));
 sg13g2_dfrbp_1 _1241_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net229),
    .D(_0071_),
    .Q_N(_0566_),
    .Q(\reg_file.registers[5][5] ));
 sg13g2_dfrbp_1 _1242_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net225),
    .D(_0072_),
    .Q_N(_0565_),
    .Q(\reg_file.registers[5][6] ));
 sg13g2_dfrbp_1 _1243_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net231),
    .D(_0073_),
    .Q_N(_0564_),
    .Q(\reg_file.registers[5][7] ));
 sg13g2_tielo tt_um_riscv_mini_15 (.L_LO(net15));
 sg13g2_tielo tt_um_riscv_mini_16 (.L_LO(net16));
 sg13g2_tielo tt_um_riscv_mini_17 (.L_LO(net17));
 sg13g2_tielo tt_um_riscv_mini_18 (.L_LO(net18));
 sg13g2_tielo tt_um_riscv_mini_19 (.L_LO(net19));
 sg13g2_tielo tt_um_riscv_mini_20 (.L_LO(net20));
 sg13g2_tielo tt_um_riscv_mini_21 (.L_LO(net21));
 sg13g2_tielo tt_um_riscv_mini_22 (.L_LO(net22));
 sg13g2_tielo tt_um_riscv_mini_23 (.L_LO(net23));
 sg13g2_tielo tt_um_riscv_mini_24 (.L_LO(net24));
 sg13g2_tielo tt_um_riscv_mini_25 (.L_LO(net25));
 sg13g2_tielo tt_um_riscv_mini_26 (.L_LO(net26));
 sg13g2_tielo tt_um_riscv_mini_27 (.L_LO(net27));
 sg13g2_tielo tt_um_riscv_mini_28 (.L_LO(net28));
 sg13g2_tielo tt_um_riscv_mini_29 (.L_LO(net29));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 fanout178 (.A(net179),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(_0265_),
    .X(net180));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(net182));
 sg13g2_buf_2 fanout182 (.A(net183),
    .X(net182));
 sg13g2_buf_1 fanout183 (.A(_0240_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(net185),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_1 fanout186 (.A(_0217_),
    .X(net186));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(_0189_));
 sg13g2_buf_2 fanout188 (.A(net189),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_0340_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_0317_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_0093_),
    .X(net191));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(net193));
 sg13g2_buf_2 fanout193 (.A(_0556_),
    .X(net193));
 sg13g2_buf_4 fanout194 (.X(net194),
    .A(_0548_));
 sg13g2_buf_2 fanout195 (.A(_0548_),
    .X(net195));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(net197));
 sg13g2_buf_2 fanout197 (.A(_0539_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(_0531_));
 sg13g2_buf_4 fanout200 (.X(net200),
    .A(net201));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(_0522_));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(net203));
 sg13g2_buf_2 fanout203 (.A(_0513_),
    .X(net203));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(net205));
 sg13g2_buf_2 fanout205 (.A(_0488_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(net207),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_0489_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_0125_),
    .X(net208));
 sg13g2_buf_4 fanout209 (.X(net209),
    .A(_0103_));
 sg13g2_buf_2 fanout210 (.A(_0103_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_0089_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(net13),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(net12),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(net216),
    .X(net214));
 sg13g2_buf_1 fanout215 (.A(net216),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(uio_in[5]),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(net9),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(uio_in[1]),
    .X(net218));
 sg13g2_buf_1 fanout219 (.A(uio_in[1]),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(net221),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(uio_in[0]),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(net8),
    .X(net222));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(net7));
 sg13g2_buf_2 fanout224 (.A(net6),
    .X(net224));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(net228));
 sg13g2_buf_2 fanout226 (.A(net227),
    .X(net226));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(net228));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(net235));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(net235));
 sg13g2_buf_2 fanout230 (.A(net231),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(net235));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(net233));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(net234));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(net235));
 sg13g2_buf_4 fanout235 (.X(net235),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[6]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_riscv_mini_14 (.L_LO(net14));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\reg_file.registers[0][2] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold2 (.A(\reg_file.registers[0][0] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold3 (.A(\reg_file.registers[0][5] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold4 (.A(\reg_file.registers[0][6] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold5 (.A(\reg_file.registers[0][7] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold6 (.A(\reg_file.registers[0][1] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold7 (.A(\reg_file.registers[0][4] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold8 (.A(\reg_file.registers[0][3] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold9 (.A(\reg_file.registers[7][0] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold10 (.A(\reg_file.registers[7][2] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold11 (.A(\reg_file.registers[3][1] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold12 (.A(\reg_file.registers[5][1] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold13 (.A(\reg_file.registers[6][1] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold14 (.A(\reg_file.registers[3][7] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold15 (.A(\reg_file.registers[3][0] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold16 (.A(\reg_file.registers[2][0] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold17 (.A(\reg_file.registers[4][7] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold18 (.A(\reg_file.registers[7][3] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold19 (.A(\reg_file.registers[4][6] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold20 (.A(\reg_file.registers[4][2] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold21 (.A(\reg_file.registers[6][3] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold22 (.A(\reg_file.registers[4][1] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold23 (.A(\reg_file.registers[2][4] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold24 (.A(\reg_file.registers[7][1] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold25 (.A(\reg_file.registers[1][3] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold26 (.A(\reg_file.registers[5][6] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold27 (.A(\reg_file.registers[6][6] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold28 (.A(\reg_file.registers[2][3] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold29 (.A(\reg_file.registers[3][3] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold30 (.A(\reg_file.registers[7][6] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold31 (.A(\reg_file.registers[7][7] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold32 (.A(\reg_file.registers[4][3] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold33 (.A(\reg_file.registers[1][2] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold34 (.A(\reg_file.registers[7][4] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold35 (.A(\reg_file.registers[6][2] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold36 (.A(\reg_file.registers[2][7] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold37 (.A(\reg_file.registers[6][4] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold38 (.A(\reg_file.registers[2][2] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold39 (.A(\reg_file.registers[2][6] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold40 (.A(\reg_file.registers[1][6] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold41 (.A(\reg_file.registers[4][4] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold42 (.A(\reg_file.registers[5][4] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold43 (.A(\reg_file.registers[6][7] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold44 (.A(\reg_file.registers[5][3] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold45 (.A(\reg_file.registers[3][6] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold46 (.A(\reg_file.registers[1][7] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold47 (.A(\reg_file.registers[2][1] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold48 (.A(\reg_file.registers[3][2] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold49 (.A(\reg_file.registers[5][2] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold50 (.A(\reg_file.registers[1][1] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold51 (.A(\reg_file.registers[3][4] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold52 (.A(\reg_file.registers[1][4] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold53 (.A(\reg_file.registers[4][0] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold54 (.A(\reg_file.registers[5][7] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold55 (.A(\reg_file.registers[6][0] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold56 (.A(\reg_file.registers[1][0] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold57 (.A(\reg_file.registers[2][5] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold58 (.A(\reg_file.registers[5][0] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold59 (.A(\reg_file.registers[4][5] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold60 (.A(\reg_file.registers[6][5] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold61 (.A(\reg_file.registers[5][5] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold62 (.A(\reg_file.registers[3][5] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold63 (.A(\reg_file.registers[1][5] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold64 (.A(\reg_file.registers[7][5] ),
    .X(net93));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_277 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_312 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_4 FILLER_17_189 ();
 sg13g2_fill_2 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_221 ();
 sg13g2_decap_8 FILLER_17_226 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_decap_4 FILLER_17_240 ();
 sg13g2_fill_2 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_250 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_4 FILLER_18_182 ();
 sg13g2_fill_2 FILLER_18_186 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_fill_2 FILLER_18_209 ();
 sg13g2_fill_2 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_decap_8 FILLER_19_172 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_187 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_fill_1 FILLER_19_204 ();
 sg13g2_fill_1 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_249 ();
 sg13g2_fill_2 FILLER_19_264 ();
 sg13g2_fill_1 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_140 ();
 sg13g2_fill_2 FILLER_20_171 ();
 sg13g2_fill_1 FILLER_20_173 ();
 sg13g2_decap_4 FILLER_20_200 ();
 sg13g2_decap_4 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_decap_4 FILLER_20_299 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_decap_4 FILLER_20_318 ();
 sg13g2_fill_2 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_342 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_decap_4 FILLER_21_157 ();
 sg13g2_decap_4 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_190 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_204 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_2 FILLER_21_221 ();
 sg13g2_decap_8 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_243 ();
 sg13g2_fill_2 FILLER_21_303 ();
 sg13g2_fill_1 FILLER_21_310 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_2 FILLER_22_151 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_fill_2 FILLER_22_216 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_228 ();
 sg13g2_fill_1 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_fill_2 FILLER_22_256 ();
 sg13g2_fill_1 FILLER_22_258 ();
 sg13g2_fill_2 FILLER_22_285 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_375 ();
 sg13g2_fill_2 FILLER_22_385 ();
 sg13g2_fill_1 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_103 ();
 sg13g2_fill_1 FILLER_23_110 ();
 sg13g2_decap_8 FILLER_23_117 ();
 sg13g2_fill_2 FILLER_23_124 ();
 sg13g2_fill_1 FILLER_23_126 ();
 sg13g2_decap_4 FILLER_23_172 ();
 sg13g2_fill_2 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_decap_4 FILLER_23_196 ();
 sg13g2_fill_2 FILLER_23_205 ();
 sg13g2_decap_4 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_215 ();
 sg13g2_fill_2 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_decap_4 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_decap_4 FILLER_23_350 ();
 sg13g2_fill_2 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_76 ();
 sg13g2_fill_2 FILLER_24_90 ();
 sg13g2_fill_2 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_128 ();
 sg13g2_fill_2 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_155 ();
 sg13g2_decap_8 FILLER_24_170 ();
 sg13g2_fill_2 FILLER_24_177 ();
 sg13g2_fill_1 FILLER_24_179 ();
 sg13g2_decap_4 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_192 ();
 sg13g2_decap_4 FILLER_24_254 ();
 sg13g2_fill_1 FILLER_24_258 ();
 sg13g2_decap_8 FILLER_24_276 ();
 sg13g2_fill_2 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_fill_2 FILLER_24_370 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_4 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_71 ();
 sg13g2_decap_8 FILLER_25_97 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_123 ();
 sg13g2_fill_2 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_165 ();
 sg13g2_fill_1 FILLER_25_167 ();
 sg13g2_decap_4 FILLER_25_207 ();
 sg13g2_fill_2 FILLER_25_211 ();
 sg13g2_decap_4 FILLER_25_218 ();
 sg13g2_fill_1 FILLER_25_222 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_330 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_2 FILLER_26_25 ();
 sg13g2_fill_2 FILLER_26_69 ();
 sg13g2_fill_1 FILLER_26_89 ();
 sg13g2_fill_2 FILLER_26_117 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_decap_4 FILLER_26_136 ();
 sg13g2_decap_4 FILLER_26_144 ();
 sg13g2_fill_2 FILLER_26_148 ();
 sg13g2_fill_2 FILLER_26_155 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_decap_4 FILLER_26_176 ();
 sg13g2_decap_8 FILLER_26_185 ();
 sg13g2_fill_2 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_194 ();
 sg13g2_fill_2 FILLER_26_221 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_269 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_312 ();
 sg13g2_fill_1 FILLER_26_314 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_fill_1 FILLER_26_350 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_30 ();
 sg13g2_decap_4 FILLER_27_41 ();
 sg13g2_decap_8 FILLER_27_50 ();
 sg13g2_fill_2 FILLER_27_57 ();
 sg13g2_decap_8 FILLER_27_69 ();
 sg13g2_decap_8 FILLER_27_76 ();
 sg13g2_fill_2 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_95 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_4 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_178 ();
 sg13g2_fill_1 FILLER_27_180 ();
 sg13g2_fill_2 FILLER_27_217 ();
 sg13g2_fill_1 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_229 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_decap_4 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_2 FILLER_27_321 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_fill_2 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_fill_1 FILLER_28_21 ();
 sg13g2_decap_4 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_46 ();
 sg13g2_decap_4 FILLER_28_52 ();
 sg13g2_fill_2 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_decap_4 FILLER_28_125 ();
 sg13g2_fill_1 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_163 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_260 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_346 ();
 sg13g2_fill_2 FILLER_28_378 ();
 sg13g2_fill_1 FILLER_28_380 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_14 ();
 sg13g2_fill_2 FILLER_29_18 ();
 sg13g2_fill_2 FILLER_29_54 ();
 sg13g2_decap_8 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_83 ();
 sg13g2_fill_2 FILLER_29_106 ();
 sg13g2_fill_1 FILLER_29_108 ();
 sg13g2_decap_8 FILLER_29_118 ();
 sg13g2_decap_8 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_132 ();
 sg13g2_fill_2 FILLER_29_138 ();
 sg13g2_fill_1 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_180 ();
 sg13g2_fill_1 FILLER_29_182 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_fill_1 FILLER_29_208 ();
 sg13g2_fill_2 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_262 ();
 sg13g2_fill_1 FILLER_29_289 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_fill_2 FILLER_29_312 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_381 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_25 ();
 sg13g2_decap_8 FILLER_30_47 ();
 sg13g2_decap_8 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_99 ();
 sg13g2_decap_8 FILLER_30_143 ();
 sg13g2_fill_2 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_152 ();
 sg13g2_decap_8 FILLER_30_165 ();
 sg13g2_decap_4 FILLER_30_172 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_decap_8 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_204 ();
 sg13g2_decap_8 FILLER_30_209 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_246 ();
 sg13g2_decap_4 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_277 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_fill_2 FILLER_30_369 ();
 sg13g2_fill_2 FILLER_30_395 ();
 sg13g2_fill_1 FILLER_30_397 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_28 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_fill_2 FILLER_31_73 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_81 ();
 sg13g2_fill_1 FILLER_31_83 ();
 sg13g2_decap_8 FILLER_31_92 ();
 sg13g2_fill_2 FILLER_31_99 ();
 sg13g2_fill_1 FILLER_31_101 ();
 sg13g2_fill_2 FILLER_31_125 ();
 sg13g2_fill_2 FILLER_31_151 ();
 sg13g2_fill_2 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_decap_4 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_249 ();
 sg13g2_decap_8 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_decap_8 FILLER_31_278 ();
 sg13g2_decap_8 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_317 ();
 sg13g2_fill_1 FILLER_31_319 ();
 sg13g2_fill_2 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_2 FILLER_32_32 ();
 sg13g2_decap_8 FILLER_32_44 ();
 sg13g2_decap_8 FILLER_32_51 ();
 sg13g2_fill_2 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_72 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_decap_8 FILLER_32_94 ();
 sg13g2_decap_4 FILLER_32_101 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_fill_2 FILLER_32_124 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_fill_2 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_146 ();
 sg13g2_fill_1 FILLER_32_157 ();
 sg13g2_decap_8 FILLER_32_162 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_decap_4 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_246 ();
 sg13g2_fill_1 FILLER_32_253 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_fill_1 FILLER_32_261 ();
 sg13g2_decap_4 FILLER_32_270 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_fill_2 FILLER_32_304 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_355 ();
 sg13g2_fill_1 FILLER_32_384 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_53 ();
 sg13g2_fill_2 FILLER_33_66 ();
 sg13g2_fill_2 FILLER_33_76 ();
 sg13g2_fill_1 FILLER_33_78 ();
 sg13g2_decap_4 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_102 ();
 sg13g2_fill_2 FILLER_33_121 ();
 sg13g2_fill_1 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_decap_8 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_decap_4 FILLER_33_174 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_fill_2 FILLER_33_184 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_decap_8 FILLER_33_218 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_4 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_4 FILLER_34_28 ();
 sg13g2_decap_4 FILLER_34_47 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_60 ();
 sg13g2_decap_4 FILLER_34_75 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_2 FILLER_34_97 ();
 sg13g2_decap_4 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_148 ();
 sg13g2_decap_4 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_183 ();
 sg13g2_fill_2 FILLER_34_195 ();
 sg13g2_fill_2 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_214 ();
 sg13g2_fill_2 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_fill_2 FILLER_34_236 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_fill_2 FILLER_34_257 ();
 sg13g2_fill_1 FILLER_34_259 ();
 sg13g2_decap_4 FILLER_34_265 ();
 sg13g2_decap_4 FILLER_34_273 ();
 sg13g2_fill_2 FILLER_34_277 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_23 ();
 sg13g2_fill_1 FILLER_35_44 ();
 sg13g2_fill_2 FILLER_35_68 ();
 sg13g2_fill_2 FILLER_35_75 ();
 sg13g2_fill_1 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_95 ();
 sg13g2_fill_1 FILLER_35_97 ();
 sg13g2_fill_1 FILLER_35_103 ();
 sg13g2_decap_8 FILLER_35_123 ();
 sg13g2_decap_4 FILLER_35_135 ();
 sg13g2_decap_4 FILLER_35_152 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_216 ();
 sg13g2_fill_1 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_255 ();
 sg13g2_decap_4 FILLER_35_268 ();
 sg13g2_fill_2 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_fill_2 FILLER_35_334 ();
 sg13g2_fill_1 FILLER_35_362 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_40 ();
 sg13g2_fill_1 FILLER_36_47 ();
 sg13g2_fill_2 FILLER_36_52 ();
 sg13g2_fill_1 FILLER_36_58 ();
 sg13g2_fill_2 FILLER_36_64 ();
 sg13g2_fill_1 FILLER_36_71 ();
 sg13g2_fill_2 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_83 ();
 sg13g2_decap_4 FILLER_36_111 ();
 sg13g2_fill_1 FILLER_36_125 ();
 sg13g2_decap_8 FILLER_36_151 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_168 ();
 sg13g2_fill_1 FILLER_36_204 ();
 sg13g2_decap_4 FILLER_36_210 ();
 sg13g2_fill_2 FILLER_36_227 ();
 sg13g2_fill_1 FILLER_36_229 ();
 sg13g2_fill_2 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_241 ();
 sg13g2_fill_2 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_108 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_decap_8 FILLER_37_137 ();
 sg13g2_decap_4 FILLER_37_144 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_167 ();
 sg13g2_fill_2 FILLER_37_174 ();
 sg13g2_decap_4 FILLER_37_180 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_decap_4 FILLER_37_200 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_fill_2 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_342 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_4 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_120 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_166 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_2 FILLER_38_237 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_2 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_286 ();
 sg13g2_fill_2 FILLER_38_318 ();
 sg13g2_fill_1 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_354 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net24;
 assign uio_out[3] = net25;
 assign uio_out[4] = net26;
 assign uio_out[5] = net27;
 assign uio_out[6] = net28;
 assign uio_out[7] = net29;
endmodule

module tt_um_jp_cd101_saw (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire clknet_0_clk;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire data;
 wire \stop.adsr_ai[0] ;
 wire \stop.adsr_ai[1] ;
 wire \stop.adsr_ai[2] ;
 wire \stop.adsr_ai[3] ;
 wire \stop.adsr_ai[4] ;
 wire \stop.adsr_ai[5] ;
 wire \stop.adsr_ai[6] ;
 wire \stop.adsr_ai[7] ;
 wire \stop.adsr_di[0] ;
 wire \stop.adsr_di[1] ;
 wire \stop.adsr_di[2] ;
 wire \stop.adsr_di[3] ;
 wire \stop.adsr_di[4] ;
 wire \stop.adsr_di[5] ;
 wire \stop.adsr_di[6] ;
 wire \stop.adsr_di[7] ;
 wire \stop.adsr_ri[0] ;
 wire \stop.adsr_ri[1] ;
 wire \stop.adsr_ri[2] ;
 wire \stop.adsr_ri[3] ;
 wire \stop.adsr_ri[4] ;
 wire \stop.adsr_ri[5] ;
 wire \stop.adsr_ri[6] ;
 wire \stop.adsr_ri[7] ;
 wire \stop.adsr_s[0] ;
 wire \stop.adsr_s[1] ;
 wire \stop.adsr_s[2] ;
 wire \stop.adsr_s[3] ;
 wire \stop.adsr_s[4] ;
 wire \stop.adsr_s[5] ;
 wire \stop.adsr_s[6] ;
 wire \stop.adsr_s[7] ;
 wire \stop.ctrl.cfg[32] ;
 wire \stop.ctrl.cfg[33] ;
 wire \stop.ctrl.cfg[34] ;
 wire \stop.ctrl.cfg[35] ;
 wire \stop.ctrl.cfg[36] ;
 wire \stop.ctrl.cfg[37] ;
 wire \stop.ctrl.cfg[38] ;
 wire \stop.ctrl.cfg[39] ;
 wire \stop.ctrl.cfg[40] ;
 wire \stop.ctrl.cfg[41] ;
 wire \stop.ctrl.cfg[42] ;
 wire \stop.ctrl.cfg[43] ;
 wire \stop.ctrl.cfg[44] ;
 wire \stop.ctrl.cfg[45] ;
 wire \stop.ctrl.cfg[46] ;
 wire \stop.ctrl.cfg[47] ;
 wire \stop.ctrl.cfg[48] ;
 wire \stop.ctrl.cfg[49] ;
 wire \stop.ctrl.cfg[50] ;
 wire \stop.ctrl.cfg[51] ;
 wire \stop.ctrl.cfg[52] ;
 wire \stop.ctrl.cfg[53] ;
 wire \stop.ctrl.cfg[54] ;
 wire \stop.ctrl.cfg[55] ;
 wire \stop.ctrl.cfg[56] ;
 wire \stop.ctrl.cfg[57] ;
 wire \stop.ctrl.cfg[58] ;
 wire \stop.ctrl.cfg[59] ;
 wire \stop.ctrl.first_bit ;
 wire \stop.ctrl.first_bit_reg ;
 wire \stop.ctrl.trig ;
 wire \stop.dbg_adsr0 ;
 wire \stop.dbg_adsr_filt0 ;
 wire \stop.dbg_adsr_reg0 ;
 wire \stop.dbg_clk_adsr ;
 wire \stop.dbg_clk_sample ;
 wire \stop.dbg_env0 ;
 wire \stop.dbg_osc0 ;
 wire \stop.dbg_rstn ;
 wire \stop.dbg_trig ;
 wire \stop.syn.adsr_data[10] ;
 wire \stop.syn.adsr_data[11] ;
 wire \stop.syn.adsr_data[12] ;
 wire \stop.syn.adsr_data[13] ;
 wire \stop.syn.adsr_data[14] ;
 wire \stop.syn.adsr_data[15] ;
 wire \stop.syn.adsr_data[1] ;
 wire \stop.syn.adsr_data[2] ;
 wire \stop.syn.adsr_data[3] ;
 wire \stop.syn.adsr_data[4] ;
 wire \stop.syn.adsr_data[5] ;
 wire \stop.syn.adsr_data[6] ;
 wire \stop.syn.adsr_data[7] ;
 wire \stop.syn.adsr_data[8] ;
 wire \stop.syn.adsr_data[9] ;
 wire \stop.syn.adsr_data_reg[10] ;
 wire \stop.syn.adsr_data_reg[11] ;
 wire \stop.syn.adsr_data_reg[12] ;
 wire \stop.syn.adsr_data_reg[13] ;
 wire \stop.syn.adsr_data_reg[14] ;
 wire \stop.syn.adsr_data_reg[15] ;
 wire \stop.syn.adsr_data_reg[1] ;
 wire \stop.syn.adsr_data_reg[2] ;
 wire \stop.syn.adsr_data_reg[3] ;
 wire \stop.syn.adsr_data_reg[4] ;
 wire \stop.syn.adsr_data_reg[5] ;
 wire \stop.syn.adsr_data_reg[6] ;
 wire \stop.syn.adsr_data_reg[7] ;
 wire \stop.syn.adsr_data_reg[8] ;
 wire \stop.syn.adsr_data_reg[9] ;
 wire \stop.syn.adsri.envelope[1] ;
 wire \stop.syn.adsri.envelope[2] ;
 wire \stop.syn.adsri.envelope[3] ;
 wire \stop.syn.adsri.envelope[4] ;
 wire \stop.syn.adsri.envelope[5] ;
 wire \stop.syn.adsri.envelope[6] ;
 wire \stop.syn.adsri.envelope[7] ;
 wire \stop.syn.adsri.rstn ;
 wire \stop.syn.adsri.state[0] ;
 wire \stop.syn.adsri.state[1] ;
 wire \stop.syn.adsri.state[2] ;
 wire \stop.syn.adsri.state[3] ;
 wire \stop.syn.adsri.state[4] ;
 wire \stop.syn.adsri.trig ;
 wire \stop.syn.clk_mult ;
 wire \stop.syn.clk_sample_x2 ;
 wire \stop.syn.clki.arstn ;
 wire \stop.syn.clki.gen[0].inst.q ;
 wire \stop.syn.clki.gen[10].inst.clk ;
 wire \stop.syn.clki.gen[10].inst.q ;
 wire \stop.syn.clki.gen[11].inst.q ;
 wire \stop.syn.clki.gen[12].inst.q ;
 wire \stop.syn.clki.gen[13].inst.q ;
 wire \stop.syn.clki.gen[14].inst.q ;
 wire \stop.syn.clki.gen[1].inst.q ;
 wire \stop.syn.clki.gen[2].inst.q ;
 wire \stop.syn.clki.gen[3].inst.q ;
 wire \stop.syn.clki.gen[5].inst.q ;
 wire \stop.syn.clki.gen[6].inst.q ;
 wire \stop.syn.daci.accumulator[0] ;
 wire \stop.syn.daci.accumulator[10] ;
 wire \stop.syn.daci.accumulator[11] ;
 wire \stop.syn.daci.accumulator[12] ;
 wire \stop.syn.daci.accumulator[13] ;
 wire \stop.syn.daci.accumulator[14] ;
 wire \stop.syn.daci.accumulator[15] ;
 wire \stop.syn.daci.accumulator[1] ;
 wire \stop.syn.daci.accumulator[2] ;
 wire \stop.syn.daci.accumulator[3] ;
 wire \stop.syn.daci.accumulator[4] ;
 wire \stop.syn.daci.accumulator[5] ;
 wire \stop.syn.daci.accumulator[6] ;
 wire \stop.syn.daci.accumulator[7] ;
 wire \stop.syn.daci.accumulator[8] ;
 wire \stop.syn.daci.accumulator[9] ;
 wire \stop.syn.daci.din[10] ;
 wire \stop.syn.daci.din[11] ;
 wire \stop.syn.daci.din[12] ;
 wire \stop.syn.daci.din[13] ;
 wire \stop.syn.daci.din[14] ;
 wire \stop.syn.daci.din[15] ;
 wire \stop.syn.daci.din[1] ;
 wire \stop.syn.daci.din[2] ;
 wire \stop.syn.daci.din[3] ;
 wire \stop.syn.daci.din[4] ;
 wire \stop.syn.daci.din[5] ;
 wire \stop.syn.daci.din[6] ;
 wire \stop.syn.daci.din[7] ;
 wire \stop.syn.daci.din[8] ;
 wire \stop.syn.daci.din[9] ;
 wire \stop.syn.filt.m1.b_bit ;
 wire \stop.syn.filt.m1.b_latched[1] ;
 wire \stop.syn.filt.m1.b_latched[2] ;
 wire \stop.syn.filt.m1.b_latched[3] ;
 wire \stop.syn.filt.m1.b_latched[4] ;
 wire \stop.syn.filt.m1.b_latched[5] ;
 wire \stop.syn.filt.m1.b_latched[6] ;
 wire \stop.syn.filt.m1.b_latched[7] ;
 wire \stop.syn.filt.m1.sum[10] ;
 wire \stop.syn.filt.m1.sum[11] ;
 wire \stop.syn.filt.m1.sum[12] ;
 wire \stop.syn.filt.m1.sum[13] ;
 wire \stop.syn.filt.m1.sum[14] ;
 wire \stop.syn.filt.m1.sum[15] ;
 wire \stop.syn.filt.m1.sum[16] ;
 wire \stop.syn.filt.m1.sum[1] ;
 wire \stop.syn.filt.m1.sum[2] ;
 wire \stop.syn.filt.m1.sum[3] ;
 wire \stop.syn.filt.m1.sum[4] ;
 wire \stop.syn.filt.m1.sum[5] ;
 wire \stop.syn.filt.m1.sum[6] ;
 wire \stop.syn.filt.m1.sum[7] ;
 wire \stop.syn.filt.m1.sum[8] ;
 wire \stop.syn.filt.m1.sum[9] ;
 wire \stop.syn.filt.m1.sum_in2[0] ;
 wire \stop.syn.filt.m1.sum_in2[10] ;
 wire \stop.syn.filt.m1.sum_in2[11] ;
 wire \stop.syn.filt.m1.sum_in2[12] ;
 wire \stop.syn.filt.m1.sum_in2[13] ;
 wire \stop.syn.filt.m1.sum_in2[14] ;
 wire \stop.syn.filt.m1.sum_in2[15] ;
 wire \stop.syn.filt.m1.sum_in2[1] ;
 wire \stop.syn.filt.m1.sum_in2[2] ;
 wire \stop.syn.filt.m1.sum_in2[3] ;
 wire \stop.syn.filt.m1.sum_in2[4] ;
 wire \stop.syn.filt.m1.sum_in2[5] ;
 wire \stop.syn.filt.m1.sum_in2[6] ;
 wire \stop.syn.filt.m1.sum_in2[7] ;
 wire \stop.syn.filt.m1.sum_in2[8] ;
 wire \stop.syn.filt.m1.sum_in2[9] ;
 wire \stop.syn.filt.m2.b_bit ;
 wire \stop.syn.filt.m2.b_latched[1] ;
 wire \stop.syn.filt.m2.b_latched[2] ;
 wire \stop.syn.filt.m2.b_latched[3] ;
 wire \stop.syn.filt.m2.b_latched[4] ;
 wire \stop.syn.filt.m2.b_latched[5] ;
 wire \stop.syn.filt.m2.b_latched[6] ;
 wire \stop.syn.filt.m2.b_latched[7] ;
 wire \stop.syn.filt.m2.sum[10] ;
 wire \stop.syn.filt.m2.sum[11] ;
 wire \stop.syn.filt.m2.sum[12] ;
 wire \stop.syn.filt.m2.sum[13] ;
 wire \stop.syn.filt.m2.sum[14] ;
 wire \stop.syn.filt.m2.sum[15] ;
 wire \stop.syn.filt.m2.sum[16] ;
 wire \stop.syn.filt.m2.sum[1] ;
 wire \stop.syn.filt.m2.sum[2] ;
 wire \stop.syn.filt.m2.sum[3] ;
 wire \stop.syn.filt.m2.sum[4] ;
 wire \stop.syn.filt.m2.sum[5] ;
 wire \stop.syn.filt.m2.sum[6] ;
 wire \stop.syn.filt.m2.sum[7] ;
 wire \stop.syn.filt.m2.sum[8] ;
 wire \stop.syn.filt.m2.sum[9] ;
 wire \stop.syn.filt.m2.sum_in2[0] ;
 wire \stop.syn.filt.m2.sum_in2[10] ;
 wire \stop.syn.filt.m2.sum_in2[11] ;
 wire \stop.syn.filt.m2.sum_in2[12] ;
 wire \stop.syn.filt.m2.sum_in2[13] ;
 wire \stop.syn.filt.m2.sum_in2[14] ;
 wire \stop.syn.filt.m2.sum_in2[15] ;
 wire \stop.syn.filt.m2.sum_in2[1] ;
 wire \stop.syn.filt.m2.sum_in2[2] ;
 wire \stop.syn.filt.m2.sum_in2[3] ;
 wire \stop.syn.filt.m2.sum_in2[4] ;
 wire \stop.syn.filt.m2.sum_in2[5] ;
 wire \stop.syn.filt.m2.sum_in2[6] ;
 wire \stop.syn.filt.m2.sum_in2[7] ;
 wire \stop.syn.filt.m2.sum_in2[8] ;
 wire \stop.syn.filt.m2.sum_in2[9] ;
 wire \stop.syn.osc_data[1] ;
 wire \stop.syn.osc_data[2] ;
 wire \stop.syn.osc_data[3] ;
 wire \stop.syn.osc_data[4] ;
 wire \stop.syn.osc_data[5] ;
 wire \stop.syn.osc_data[6] ;
 wire \stop.syn.osc_data[7] ;
 wire \stop.syn.osci.counter[0] ;
 wire \stop.syn.osci.counter[1] ;
 wire \stop.syn.osci.counter[2] ;
 wire \stop.syn.osci.counter[3] ;
 wire \stop.syn.rstn_fst_reg1 ;
 wire \stop.syn.rstn_fst_reg2 ;
 wire \stop.syn.rstn_reg1 ;
 wire \stop.syn.smul8.b_bit ;
 wire \stop.syn.smul8.b_latched[1] ;
 wire \stop.syn.smul8.b_latched[2] ;
 wire \stop.syn.smul8.b_latched[3] ;
 wire \stop.syn.smul8.b_latched[4] ;
 wire \stop.syn.smul8.b_latched[5] ;
 wire \stop.syn.smul8.b_latched[6] ;
 wire \stop.syn.smul8.b_latched[7] ;
 wire \stop.syn.trig_reg1 ;
 wire net105;
 wire net106;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;

 sg13g2_inv_1 _1011_ (.Y(_0315_),
    .A(\stop.syn.adsri.envelope[1] ));
 sg13g2_inv_1 _1012_ (.Y(_0316_),
    .A(\stop.dbg_env0 ));
 sg13g2_inv_1 _1013_ (.Y(_0080_),
    .A(\stop.ctrl.first_bit ));
 sg13g2_inv_2 _1014_ (.Y(_0317_),
    .A(\stop.syn.adsri.state[3] ));
 sg13g2_inv_1 _1015_ (.Y(_0318_),
    .A(\stop.syn.adsri.state[0] ));
 sg13g2_inv_1 _1016_ (.Y(_0319_),
    .A(\stop.syn.adsri.trig ));
 sg13g2_inv_4 _1017_ (.A(net277),
    .Y(_0320_));
 sg13g2_inv_1 _1018_ (.Y(_0321_),
    .A(\stop.adsr_ai[2] ));
 sg13g2_inv_1 _1019_ (.Y(_0322_),
    .A(\stop.adsr_ai[3] ));
 sg13g2_inv_1 _1020_ (.Y(_0323_),
    .A(\stop.adsr_ai[4] ));
 sg13g2_inv_1 _1021_ (.Y(_0324_),
    .A(\stop.adsr_ai[5] ));
 sg13g2_inv_1 _1022_ (.Y(_0325_),
    .A(\stop.adsr_ai[6] ));
 sg13g2_inv_1 _1023_ (.Y(_0326_),
    .A(\stop.adsr_ai[7] ));
 sg13g2_inv_1 _1024_ (.Y(_0081_),
    .A(net2));
 sg13g2_nor2b_1 _1025_ (.A(\stop.syn.clk_sample_x2 ),
    .B_N(net300),
    .Y(_0327_));
 sg13g2_inv_4 _1026_ (.A(net295),
    .Y(_0131_));
 sg13g2_and2_1 _1027_ (.A(\stop.ctrl.cfg[51] ),
    .B(net288),
    .X(_0155_));
 sg13g2_and2_1 _1028_ (.A(\stop.ctrl.cfg[59] ),
    .B(net289),
    .X(_0154_));
 sg13g2_and2_1 _1029_ (.A(\stop.syn.adsri.envelope[7] ),
    .B(net298),
    .X(_0132_));
 sg13g2_a22oi_1 _1030_ (.Y(_0328_),
    .B1(\stop.adsr_di[6] ),
    .B2(net282),
    .A2(\stop.adsr_ri[6] ),
    .A1(net283));
 sg13g2_o21ai_1 _1031_ (.B1(_0328_),
    .Y(_0329_),
    .A1(_0317_),
    .A2(_0325_));
 sg13g2_and2_1 _1032_ (.A(\stop.syn.adsri.envelope[6] ),
    .B(_0329_),
    .X(_0330_));
 sg13g2_xor2_1 _1033_ (.B(_0329_),
    .A(\stop.syn.adsri.envelope[6] ),
    .X(_0331_));
 sg13g2_a22oi_1 _1034_ (.Y(_0332_),
    .B1(\stop.adsr_di[5] ),
    .B2(net282),
    .A2(\stop.adsr_ri[5] ),
    .A1(net283));
 sg13g2_o21ai_1 _1035_ (.B1(_0332_),
    .Y(_0333_),
    .A1(_0317_),
    .A2(_0324_));
 sg13g2_and2_1 _1036_ (.A(\stop.syn.adsri.envelope[5] ),
    .B(_0333_),
    .X(_0334_));
 sg13g2_a22oi_1 _1037_ (.Y(_0335_),
    .B1(\stop.adsr_di[4] ),
    .B2(\stop.syn.adsri.state[2] ),
    .A2(\stop.adsr_ri[4] ),
    .A1(net284));
 sg13g2_o21ai_1 _1038_ (.B1(_0335_),
    .Y(_0336_),
    .A1(_0317_),
    .A2(_0323_));
 sg13g2_and2_1 _1039_ (.A(\stop.syn.adsri.envelope[4] ),
    .B(_0336_),
    .X(_0337_));
 sg13g2_a22oi_1 _1040_ (.Y(_0338_),
    .B1(\stop.adsr_di[3] ),
    .B2(\stop.syn.adsri.state[2] ),
    .A2(\stop.adsr_ri[3] ),
    .A1(net284));
 sg13g2_o21ai_1 _1041_ (.B1(_0338_),
    .Y(_0339_),
    .A1(_0317_),
    .A2(_0322_));
 sg13g2_nand2_1 _1042_ (.Y(_0340_),
    .A(\stop.syn.adsri.envelope[3] ),
    .B(_0339_));
 sg13g2_nor2_1 _1043_ (.A(\stop.syn.adsri.envelope[3] ),
    .B(_0339_),
    .Y(_0341_));
 sg13g2_a22oi_1 _1044_ (.Y(_0342_),
    .B1(\stop.adsr_di[2] ),
    .B2(\stop.syn.adsri.state[2] ),
    .A2(\stop.adsr_ri[2] ),
    .A1(net284));
 sg13g2_o21ai_1 _1045_ (.B1(_0342_),
    .Y(_0343_),
    .A1(_0317_),
    .A2(_0321_));
 sg13g2_and2_1 _1046_ (.A(\stop.syn.adsri.envelope[2] ),
    .B(_0343_),
    .X(_0344_));
 sg13g2_nand2_1 _1047_ (.Y(_0345_),
    .A(\stop.syn.adsri.state[3] ),
    .B(\stop.adsr_ai[1] ));
 sg13g2_a22oi_1 _1048_ (.Y(_0346_),
    .B1(\stop.adsr_di[1] ),
    .B2(net282),
    .A2(\stop.adsr_ri[1] ),
    .A1(net284));
 sg13g2_a21oi_1 _1049_ (.A1(_0345_),
    .A2(_0346_),
    .Y(_0347_),
    .B1(_0315_));
 sg13g2_a21o_1 _1050_ (.A2(_0346_),
    .A1(_0345_),
    .B1(_0315_),
    .X(_0348_));
 sg13g2_nand2_1 _1051_ (.Y(_0349_),
    .A(net283),
    .B(\stop.adsr_ri[0] ));
 sg13g2_a22oi_1 _1052_ (.Y(_0350_),
    .B1(\stop.adsr_ai[0] ),
    .B2(\stop.syn.adsri.state[3] ),
    .A2(\stop.adsr_di[0] ),
    .A1(net282));
 sg13g2_a21o_1 _1053_ (.A2(_0350_),
    .A1(_0349_),
    .B1(_0316_),
    .X(_0351_));
 sg13g2_and3_1 _1054_ (.X(_0352_),
    .A(_0315_),
    .B(_0345_),
    .C(_0346_));
 sg13g2_nor2_1 _1055_ (.A(_0347_),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_o21ai_1 _1056_ (.B1(_0348_),
    .Y(_0354_),
    .A1(_0351_),
    .A2(_0352_));
 sg13g2_xor2_1 _1057_ (.B(_0343_),
    .A(\stop.syn.adsri.envelope[2] ),
    .X(_0355_));
 sg13g2_a21oi_2 _1058_ (.B1(_0344_),
    .Y(_0356_),
    .A2(_0355_),
    .A1(_0354_));
 sg13g2_a21oi_2 _1059_ (.B1(_0341_),
    .Y(_0357_),
    .A2(_0356_),
    .A1(_0340_));
 sg13g2_xor2_1 _1060_ (.B(_0336_),
    .A(\stop.syn.adsri.envelope[4] ),
    .X(_0358_));
 sg13g2_a21oi_1 _1061_ (.A1(_0357_),
    .A2(_0358_),
    .Y(_0359_),
    .B1(_0337_));
 sg13g2_xor2_1 _1062_ (.B(_0333_),
    .A(\stop.syn.adsri.envelope[5] ),
    .X(_0360_));
 sg13g2_and2_1 _1063_ (.A(_0358_),
    .B(_0360_),
    .X(_0361_));
 sg13g2_a21o_1 _1064_ (.A2(_0360_),
    .A1(_0337_),
    .B1(_0334_),
    .X(_0362_));
 sg13g2_a21o_1 _1065_ (.A2(_0361_),
    .A1(_0357_),
    .B1(_0362_),
    .X(_0363_));
 sg13g2_a21oi_1 _1066_ (.A1(_0331_),
    .A2(_0363_),
    .Y(_0364_),
    .B1(_0330_));
 sg13g2_a22oi_1 _1067_ (.Y(_0365_),
    .B1(\stop.adsr_di[7] ),
    .B2(net282),
    .A2(\stop.adsr_ri[7] ),
    .A1(net283));
 sg13g2_o21ai_1 _1068_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_0317_),
    .A2(_0326_));
 sg13g2_xor2_1 _1069_ (.B(_0366_),
    .A(\stop.syn.adsri.envelope[7] ),
    .X(_0367_));
 sg13g2_nor2b_1 _1070_ (.A(_0364_),
    .B_N(_0367_),
    .Y(_0368_));
 sg13g2_xnor2_1 _1071_ (.Y(_0369_),
    .A(_0364_),
    .B(_0367_));
 sg13g2_inv_1 _1072_ (.Y(_0370_),
    .A(_0369_));
 sg13g2_xnor2_1 _1073_ (.Y(_0371_),
    .A(\stop.adsr_s[7] ),
    .B(_0369_));
 sg13g2_xnor2_1 _1074_ (.Y(_0372_),
    .A(_0331_),
    .B(_0363_));
 sg13g2_xor2_1 _1075_ (.B(_0360_),
    .A(_0359_),
    .X(_0373_));
 sg13g2_xnor2_1 _1076_ (.Y(_0374_),
    .A(_0357_),
    .B(_0358_));
 sg13g2_xnor2_1 _1077_ (.Y(_0375_),
    .A(\stop.syn.adsri.envelope[3] ),
    .B(_0339_));
 sg13g2_xnor2_1 _1078_ (.Y(_0376_),
    .A(_0356_),
    .B(_0375_));
 sg13g2_xnor2_1 _1079_ (.Y(_0377_),
    .A(_0354_),
    .B(_0355_));
 sg13g2_xor2_1 _1080_ (.B(_0377_),
    .A(\stop.adsr_s[2] ),
    .X(_0378_));
 sg13g2_xor2_1 _1081_ (.B(_0353_),
    .A(_0351_),
    .X(_0379_));
 sg13g2_xor2_1 _1082_ (.B(_0379_),
    .A(\stop.adsr_s[1] ),
    .X(_0380_));
 sg13g2_nand3_1 _1083_ (.B(_0349_),
    .C(_0350_),
    .A(_0316_),
    .Y(_0381_));
 sg13g2_nand2_1 _1084_ (.Y(_0382_),
    .A(_0351_),
    .B(_0381_));
 sg13g2_xor2_1 _1085_ (.B(_0382_),
    .A(\stop.adsr_s[0] ),
    .X(_0383_));
 sg13g2_xor2_1 _1086_ (.B(_0376_),
    .A(\stop.adsr_s[3] ),
    .X(_0384_));
 sg13g2_nand4_1 _1087_ (.B(_0380_),
    .C(_0383_),
    .A(_0378_),
    .Y(_0385_),
    .D(_0384_));
 sg13g2_xnor2_1 _1088_ (.Y(_0386_),
    .A(\stop.adsr_s[4] ),
    .B(_0374_));
 sg13g2_xnor2_1 _1089_ (.Y(_0387_),
    .A(\stop.adsr_s[5] ),
    .B(_0373_));
 sg13g2_nor3_1 _1090_ (.A(_0385_),
    .B(_0386_),
    .C(_0387_),
    .Y(_0388_));
 sg13g2_xor2_1 _1091_ (.B(_0372_),
    .A(\stop.adsr_s[6] ),
    .X(_0389_));
 sg13g2_nand3_1 _1092_ (.B(_0388_),
    .C(_0389_),
    .A(_0371_),
    .Y(_0390_));
 sg13g2_nor2b_1 _1093_ (.A(\stop.syn.adsri.state[4] ),
    .B_N(_0390_),
    .Y(_0391_));
 sg13g2_nand2_1 _1094_ (.Y(_0392_),
    .A(\stop.syn.adsri.trig ),
    .B(net281));
 sg13g2_nor2_1 _1095_ (.A(net282),
    .B(\stop.syn.adsri.state[4] ),
    .Y(_0393_));
 sg13g2_nor3_1 _1096_ (.A(_0391_),
    .B(_0392_),
    .C(_0393_),
    .Y(_0004_));
 sg13g2_a21oi_2 _1097_ (.B1(_0368_),
    .Y(_0394_),
    .A2(_0366_),
    .A1(\stop.syn.adsri.envelope[7] ));
 sg13g2_nor2_1 _1098_ (.A(net283),
    .B(net282),
    .Y(_0395_));
 sg13g2_xor2_1 _1099_ (.B(_0395_),
    .A(_0394_),
    .X(_0396_));
 sg13g2_o21ai_1 _1100_ (.B1(_0318_),
    .Y(_0397_),
    .A1(_0317_),
    .A2(_0396_));
 sg13g2_nor2b_1 _1101_ (.A(_0392_),
    .B_N(_0397_),
    .Y(_0003_));
 sg13g2_a22oi_1 _1102_ (.Y(_0398_),
    .B1(_0396_),
    .B2(\stop.syn.adsri.state[3] ),
    .A2(_0390_),
    .A1(net282));
 sg13g2_nor2_1 _1103_ (.A(_0392_),
    .B(_0398_),
    .Y(_0002_));
 sg13g2_nor2_1 _1104_ (.A(\stop.syn.adsri.trig ),
    .B(_0320_),
    .Y(_0399_));
 sg13g2_nand2_1 _1105_ (.Y(_0400_),
    .A(_0317_),
    .B(_0393_));
 sg13g2_nand2_1 _1106_ (.Y(_0401_),
    .A(_0399_),
    .B(_0400_));
 sg13g2_nand2_1 _1107_ (.Y(_0402_),
    .A(net283),
    .B(net281));
 sg13g2_o21ai_1 _1108_ (.B1(_0401_),
    .Y(_0001_),
    .A1(_0394_),
    .A2(_0402_));
 sg13g2_nand2_1 _1109_ (.Y(_0403_),
    .A(net283),
    .B(_0394_));
 sg13g2_a21oi_1 _1110_ (.A1(\stop.syn.adsri.state[0] ),
    .A2(_0399_),
    .Y(_0404_),
    .B1(_0045_));
 sg13g2_nand2_1 _1111_ (.Y(_0000_),
    .A(_0403_),
    .B(_0404_));
 sg13g2_nor2_1 _1112_ (.A(\stop.syn.smul8.b_latched[1] ),
    .B(net295),
    .Y(_0405_));
 sg13g2_a21oi_2 _1113_ (.B1(_0405_),
    .Y(_0019_),
    .A2(net295),
    .A1(_0316_));
 sg13g2_nand2_1 _1114_ (.Y(_0406_),
    .A(\stop.syn.smul8.b_latched[2] ),
    .B(_0131_));
 sg13g2_o21ai_1 _1115_ (.B1(_0406_),
    .Y(_0020_),
    .A1(_0315_),
    .A2(_0131_));
 sg13g2_mux2_1 _1116_ (.A0(\stop.syn.adsri.envelope[2] ),
    .A1(\stop.syn.smul8.b_latched[3] ),
    .S(_0131_),
    .X(_0021_));
 sg13g2_mux2_1 _1117_ (.A0(\stop.syn.adsri.envelope[3] ),
    .A1(\stop.syn.smul8.b_latched[4] ),
    .S(_0131_),
    .X(_0022_));
 sg13g2_mux2_1 _1118_ (.A0(\stop.syn.adsri.envelope[4] ),
    .A1(\stop.syn.smul8.b_latched[5] ),
    .S(_0131_),
    .X(_0023_));
 sg13g2_mux2_1 _1119_ (.A0(\stop.syn.adsri.envelope[5] ),
    .A1(\stop.syn.smul8.b_latched[6] ),
    .S(_0131_),
    .X(_0024_));
 sg13g2_mux2_1 _1120_ (.A0(\stop.syn.adsri.envelope[6] ),
    .A1(\stop.syn.smul8.b_latched[7] ),
    .S(_0131_),
    .X(_0025_));
 sg13g2_mux2_1 _1121_ (.A0(\stop.syn.filt.m2.b_latched[1] ),
    .A1(\stop.ctrl.cfg[52] ),
    .S(net289),
    .X(_0012_));
 sg13g2_mux2_1 _1122_ (.A0(\stop.syn.filt.m2.b_latched[2] ),
    .A1(\stop.ctrl.cfg[53] ),
    .S(net289),
    .X(_0013_));
 sg13g2_mux2_1 _1123_ (.A0(\stop.syn.filt.m2.b_latched[3] ),
    .A1(\stop.ctrl.cfg[54] ),
    .S(net289),
    .X(_0014_));
 sg13g2_mux2_1 _1124_ (.A0(\stop.syn.filt.m2.b_latched[4] ),
    .A1(\stop.ctrl.cfg[55] ),
    .S(net289),
    .X(_0015_));
 sg13g2_mux2_1 _1125_ (.A0(\stop.syn.filt.m2.b_latched[5] ),
    .A1(\stop.ctrl.cfg[56] ),
    .S(net294),
    .X(_0016_));
 sg13g2_mux2_1 _1126_ (.A0(\stop.syn.filt.m2.b_latched[6] ),
    .A1(\stop.ctrl.cfg[57] ),
    .S(net295),
    .X(_0017_));
 sg13g2_mux2_1 _1127_ (.A0(\stop.syn.filt.m2.b_latched[7] ),
    .A1(\stop.ctrl.cfg[58] ),
    .S(net295),
    .X(_0018_));
 sg13g2_mux2_1 _1128_ (.A0(\stop.syn.filt.m1.b_latched[1] ),
    .A1(\stop.ctrl.cfg[44] ),
    .S(net294),
    .X(_0005_));
 sg13g2_mux2_1 _1129_ (.A0(\stop.syn.filt.m1.b_latched[2] ),
    .A1(\stop.ctrl.cfg[45] ),
    .S(net288),
    .X(_0006_));
 sg13g2_mux2_1 _1130_ (.A0(\stop.syn.filt.m1.b_latched[3] ),
    .A1(\stop.ctrl.cfg[46] ),
    .S(net288),
    .X(_0007_));
 sg13g2_mux2_1 _1131_ (.A0(\stop.syn.filt.m1.b_latched[4] ),
    .A1(\stop.ctrl.cfg[47] ),
    .S(net288),
    .X(_0008_));
 sg13g2_mux2_1 _1132_ (.A0(\stop.syn.filt.m1.b_latched[5] ),
    .A1(\stop.ctrl.cfg[48] ),
    .S(net288),
    .X(_0009_));
 sg13g2_mux2_1 _1133_ (.A0(\stop.syn.filt.m1.b_latched[6] ),
    .A1(\stop.ctrl.cfg[49] ),
    .S(net288),
    .X(_0010_));
 sg13g2_mux2_1 _1134_ (.A0(\stop.syn.filt.m1.b_latched[7] ),
    .A1(\stop.ctrl.cfg[50] ),
    .S(net288),
    .X(_0011_));
 sg13g2_nand3_1 _1135_ (.B(\stop.dbg_adsr_filt0 ),
    .C(\stop.syn.filt.m1.sum_in2[0] ),
    .A(net312),
    .Y(_0407_));
 sg13g2_and3_1 _1136_ (.X(_0408_),
    .A(net312),
    .B(\stop.syn.daci.din[1] ),
    .C(\stop.syn.filt.m1.sum_in2[1] ));
 sg13g2_nand3_1 _1137_ (.B(\stop.syn.daci.din[1] ),
    .C(\stop.syn.filt.m1.sum_in2[1] ),
    .A(net312),
    .Y(_0409_));
 sg13g2_a21oi_1 _1138_ (.A1(net312),
    .A2(\stop.syn.daci.din[1] ),
    .Y(_0410_),
    .B1(\stop.syn.filt.m1.sum_in2[1] ));
 sg13g2_nor2_1 _1139_ (.A(_0408_),
    .B(_0410_),
    .Y(_0411_));
 sg13g2_xnor2_1 _1140_ (.Y(\stop.syn.filt.m1.sum[1] ),
    .A(_0407_),
    .B(_0411_));
 sg13g2_o21ai_1 _1141_ (.B1(_0409_),
    .Y(_0412_),
    .A1(_0407_),
    .A2(_0410_));
 sg13g2_and3_1 _1142_ (.X(_0413_),
    .A(net313),
    .B(\stop.syn.daci.din[2] ),
    .C(\stop.syn.filt.m1.sum_in2[2] ));
 sg13g2_a21o_1 _1143_ (.A2(\stop.syn.daci.din[2] ),
    .A1(net312),
    .B1(\stop.syn.filt.m1.sum_in2[2] ),
    .X(_0414_));
 sg13g2_nand2b_1 _1144_ (.Y(_0415_),
    .B(_0414_),
    .A_N(_0413_));
 sg13g2_xnor2_1 _1145_ (.Y(\stop.syn.filt.m1.sum[2] ),
    .A(_0412_),
    .B(_0415_));
 sg13g2_a21o_1 _1146_ (.A2(_0414_),
    .A1(_0412_),
    .B1(_0413_),
    .X(_0416_));
 sg13g2_nand2_1 _1147_ (.Y(_0417_),
    .A(net312),
    .B(\stop.syn.daci.din[3] ));
 sg13g2_nor2_1 _1148_ (.A(_0046_),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_xor2_1 _1149_ (.B(_0417_),
    .A(_0046_),
    .X(_0419_));
 sg13g2_xor2_1 _1150_ (.B(_0419_),
    .A(_0416_),
    .X(\stop.syn.filt.m1.sum[3] ));
 sg13g2_a21oi_1 _1151_ (.A1(_0416_),
    .A2(_0419_),
    .Y(_0420_),
    .B1(_0418_));
 sg13g2_nand3_1 _1152_ (.B(\stop.syn.daci.din[4] ),
    .C(\stop.syn.filt.m1.sum_in2[4] ),
    .A(net311),
    .Y(_0421_));
 sg13g2_a21o_1 _1153_ (.A2(\stop.syn.daci.din[4] ),
    .A1(net311),
    .B1(\stop.syn.filt.m1.sum_in2[4] ),
    .X(_0422_));
 sg13g2_nand2_1 _1154_ (.Y(_0423_),
    .A(_0421_),
    .B(_0422_));
 sg13g2_xor2_1 _1155_ (.B(_0423_),
    .A(_0420_),
    .X(\stop.syn.filt.m1.sum[4] ));
 sg13g2_o21ai_1 _1156_ (.B1(_0421_),
    .Y(_0424_),
    .A1(_0420_),
    .A2(_0423_));
 sg13g2_nand2_1 _1157_ (.Y(_0425_),
    .A(net311),
    .B(\stop.syn.daci.din[5] ));
 sg13g2_nor2_1 _1158_ (.A(_0047_),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_nand2_1 _1159_ (.Y(_0427_),
    .A(_0047_),
    .B(_0425_));
 sg13g2_nor2b_1 _1160_ (.A(_0426_),
    .B_N(_0427_),
    .Y(_0428_));
 sg13g2_xor2_1 _1161_ (.B(_0428_),
    .A(_0424_),
    .X(\stop.syn.filt.m1.sum[5] ));
 sg13g2_nand3_1 _1162_ (.B(\stop.syn.daci.din[6] ),
    .C(\stop.syn.filt.m1.sum_in2[6] ),
    .A(net312),
    .Y(_0429_));
 sg13g2_a21o_1 _1163_ (.A2(\stop.syn.daci.din[6] ),
    .A1(net311),
    .B1(\stop.syn.filt.m1.sum_in2[6] ),
    .X(_0430_));
 sg13g2_and2_1 _1164_ (.A(_0429_),
    .B(_0430_),
    .X(_0431_));
 sg13g2_inv_1 _1165_ (.Y(_0432_),
    .A(_0431_));
 sg13g2_o21ai_1 _1166_ (.B1(_0427_),
    .Y(_0433_),
    .A1(_0424_),
    .A2(_0426_));
 sg13g2_xnor2_1 _1167_ (.Y(\stop.syn.filt.m1.sum[6] ),
    .A(_0431_),
    .B(_0433_));
 sg13g2_o21ai_1 _1168_ (.B1(_0429_),
    .Y(_0434_),
    .A1(_0432_),
    .A2(_0433_));
 sg13g2_and3_1 _1169_ (.X(_0435_),
    .A(net311),
    .B(\stop.syn.daci.din[7] ),
    .C(\stop.syn.filt.m1.sum_in2[7] ));
 sg13g2_a21o_1 _1170_ (.A2(\stop.syn.daci.din[7] ),
    .A1(net311),
    .B1(\stop.syn.filt.m1.sum_in2[7] ),
    .X(_0436_));
 sg13g2_nand2b_1 _1171_ (.Y(_0437_),
    .B(_0436_),
    .A_N(_0435_));
 sg13g2_xnor2_1 _1172_ (.Y(\stop.syn.filt.m1.sum[7] ),
    .A(_0434_),
    .B(_0437_));
 sg13g2_a21o_1 _1173_ (.A2(_0436_),
    .A1(_0434_),
    .B1(_0435_),
    .X(_0438_));
 sg13g2_inv_1 _1174_ (.Y(_0439_),
    .A(_0438_));
 sg13g2_nand3_1 _1175_ (.B(\stop.syn.daci.din[8] ),
    .C(\stop.syn.filt.m1.sum_in2[8] ),
    .A(net311),
    .Y(_0440_));
 sg13g2_a21o_1 _1176_ (.A2(\stop.syn.daci.din[8] ),
    .A1(net311),
    .B1(\stop.syn.filt.m1.sum_in2[8] ),
    .X(_0441_));
 sg13g2_nand2_1 _1177_ (.Y(_0442_),
    .A(_0440_),
    .B(_0441_));
 sg13g2_xnor2_1 _1178_ (.Y(\stop.syn.filt.m1.sum[8] ),
    .A(_0438_),
    .B(_0442_));
 sg13g2_nand2_1 _1179_ (.Y(_0443_),
    .A(net309),
    .B(\stop.syn.daci.din[9] ));
 sg13g2_xor2_1 _1180_ (.B(_0443_),
    .A(_0048_),
    .X(_0444_));
 sg13g2_o21ai_1 _1181_ (.B1(_0440_),
    .Y(_0445_),
    .A1(_0439_),
    .A2(_0442_));
 sg13g2_xor2_1 _1182_ (.B(_0445_),
    .A(_0444_),
    .X(\stop.syn.filt.m1.sum[9] ));
 sg13g2_nand3_1 _1183_ (.B(\stop.syn.daci.din[10] ),
    .C(\stop.syn.filt.m1.sum_in2[10] ),
    .A(net309),
    .Y(_0446_));
 sg13g2_a21o_1 _1184_ (.A2(\stop.syn.daci.din[10] ),
    .A1(net309),
    .B1(\stop.syn.filt.m1.sum_in2[10] ),
    .X(_0447_));
 sg13g2_nand2_1 _1185_ (.Y(_0448_),
    .A(_0446_),
    .B(_0447_));
 sg13g2_a21o_1 _1186_ (.A2(_0443_),
    .A1(_0048_),
    .B1(_0440_),
    .X(_0449_));
 sg13g2_o21ai_1 _1187_ (.B1(_0449_),
    .Y(_0450_),
    .A1(_0048_),
    .A2(_0443_));
 sg13g2_nor2b_1 _1188_ (.A(_0442_),
    .B_N(_0444_),
    .Y(_0451_));
 sg13g2_a21oi_1 _1189_ (.A1(_0438_),
    .A2(_0451_),
    .Y(_0452_),
    .B1(_0450_));
 sg13g2_xor2_1 _1190_ (.B(_0452_),
    .A(_0448_),
    .X(\stop.syn.filt.m1.sum[10] ));
 sg13g2_a21oi_1 _1191_ (.A1(net309),
    .A2(\stop.syn.daci.din[11] ),
    .Y(_0453_),
    .B1(\stop.syn.filt.m1.sum_in2[11] ));
 sg13g2_nand3_1 _1192_ (.B(\stop.syn.daci.din[11] ),
    .C(\stop.syn.filt.m1.sum_in2[11] ),
    .A(net309),
    .Y(_0454_));
 sg13g2_nand2b_1 _1193_ (.Y(_0455_),
    .B(_0454_),
    .A_N(_0453_));
 sg13g2_o21ai_1 _1194_ (.B1(_0446_),
    .Y(_0456_),
    .A1(_0448_),
    .A2(_0452_));
 sg13g2_xnor2_1 _1195_ (.Y(\stop.syn.filt.m1.sum[11] ),
    .A(_0455_),
    .B(_0456_));
 sg13g2_nor2_1 _1196_ (.A(_0448_),
    .B(_0455_),
    .Y(_0457_));
 sg13g2_and2_1 _1197_ (.A(_0451_),
    .B(_0457_),
    .X(_0458_));
 sg13g2_o21ai_1 _1198_ (.B1(_0454_),
    .Y(_0459_),
    .A1(_0446_),
    .A2(_0453_));
 sg13g2_a221oi_1 _1199_ (.B2(_0438_),
    .C1(_0459_),
    .B1(_0458_),
    .A1(_0450_),
    .Y(_0460_),
    .A2(_0457_));
 sg13g2_nand3_1 _1200_ (.B(\stop.syn.daci.din[12] ),
    .C(\stop.syn.filt.m1.sum_in2[12] ),
    .A(net310),
    .Y(_0461_));
 sg13g2_a21o_1 _1201_ (.A2(\stop.syn.daci.din[12] ),
    .A1(net310),
    .B1(\stop.syn.filt.m1.sum_in2[12] ),
    .X(_0462_));
 sg13g2_nand2_1 _1202_ (.Y(_0463_),
    .A(_0461_),
    .B(_0462_));
 sg13g2_xor2_1 _1203_ (.B(_0463_),
    .A(_0460_),
    .X(\stop.syn.filt.m1.sum[12] ));
 sg13g2_o21ai_1 _1204_ (.B1(_0461_),
    .Y(_0464_),
    .A1(_0460_),
    .A2(_0463_));
 sg13g2_nand2_1 _1205_ (.Y(_0465_),
    .A(net310),
    .B(\stop.syn.daci.din[13] ));
 sg13g2_nor2_1 _1206_ (.A(_0049_),
    .B(_0465_),
    .Y(_0466_));
 sg13g2_xor2_1 _1207_ (.B(_0465_),
    .A(_0049_),
    .X(_0467_));
 sg13g2_xor2_1 _1208_ (.B(_0467_),
    .A(_0464_),
    .X(\stop.syn.filt.m1.sum[13] ));
 sg13g2_nand2b_1 _1209_ (.Y(_0468_),
    .B(_0467_),
    .A_N(_0463_));
 sg13g2_a21oi_1 _1210_ (.A1(_0049_),
    .A2(_0465_),
    .Y(_0469_),
    .B1(_0461_));
 sg13g2_nor2_1 _1211_ (.A(_0466_),
    .B(_0469_),
    .Y(_0470_));
 sg13g2_o21ai_1 _1212_ (.B1(_0470_),
    .Y(_0471_),
    .A1(_0460_),
    .A2(_0468_));
 sg13g2_and3_1 _1213_ (.X(_0472_),
    .A(net310),
    .B(\stop.syn.daci.din[14] ),
    .C(\stop.syn.filt.m1.sum_in2[14] ));
 sg13g2_a21o_1 _1214_ (.A2(\stop.syn.daci.din[14] ),
    .A1(net309),
    .B1(\stop.syn.filt.m1.sum_in2[14] ),
    .X(_0473_));
 sg13g2_nand2b_1 _1215_ (.Y(_0474_),
    .B(_0473_),
    .A_N(_0472_));
 sg13g2_xnor2_1 _1216_ (.Y(\stop.syn.filt.m1.sum[14] ),
    .A(_0471_),
    .B(_0474_));
 sg13g2_and3_1 _1217_ (.X(_0475_),
    .A(net310),
    .B(\stop.syn.daci.din[15] ),
    .C(\stop.syn.filt.m1.sum_in2[15] ));
 sg13g2_nand3_1 _1218_ (.B(\stop.syn.daci.din[15] ),
    .C(\stop.syn.filt.m1.sum_in2[15] ),
    .A(net309),
    .Y(_0476_));
 sg13g2_a21oi_1 _1219_ (.A1(net309),
    .A2(\stop.syn.daci.din[15] ),
    .Y(_0477_),
    .B1(\stop.syn.filt.m1.sum_in2[15] ));
 sg13g2_nor2_1 _1220_ (.A(_0475_),
    .B(_0477_),
    .Y(_0478_));
 sg13g2_a21oi_1 _1221_ (.A1(_0471_),
    .A2(_0473_),
    .Y(_0479_),
    .B1(_0472_));
 sg13g2_xnor2_1 _1222_ (.Y(\stop.syn.filt.m1.sum[15] ),
    .A(_0478_),
    .B(_0479_));
 sg13g2_nand2_1 _1223_ (.Y(_0480_),
    .A(\stop.syn.filt.m1.sum_in2[0] ),
    .B(\stop.syn.filt.m2.sum_in2[0] ));
 sg13g2_nand2_1 _1224_ (.Y(_0481_),
    .A(\stop.syn.filt.m1.sum_in2[1] ),
    .B(\stop.syn.filt.m2.sum_in2[1] ));
 sg13g2_nor2_1 _1225_ (.A(\stop.syn.filt.m1.sum_in2[1] ),
    .B(\stop.syn.filt.m2.sum_in2[1] ),
    .Y(_0482_));
 sg13g2_xor2_1 _1226_ (.B(\stop.syn.filt.m2.sum_in2[1] ),
    .A(\stop.syn.filt.m1.sum_in2[1] ),
    .X(_0483_));
 sg13g2_xnor2_1 _1227_ (.Y(_0060_),
    .A(_0480_),
    .B(_0483_));
 sg13g2_o21ai_1 _1228_ (.B1(_0481_),
    .Y(_0484_),
    .A1(_0480_),
    .A2(_0482_));
 sg13g2_and2_1 _1229_ (.A(\stop.syn.filt.m1.sum_in2[2] ),
    .B(\stop.syn.filt.m2.sum_in2[2] ),
    .X(_0485_));
 sg13g2_or2_1 _1230_ (.X(_0486_),
    .B(\stop.syn.filt.m2.sum_in2[2] ),
    .A(\stop.syn.filt.m1.sum_in2[2] ));
 sg13g2_nand2b_1 _1231_ (.Y(_0487_),
    .B(_0486_),
    .A_N(_0485_));
 sg13g2_xnor2_1 _1232_ (.Y(_0061_),
    .A(_0484_),
    .B(_0487_));
 sg13g2_a21o_1 _1233_ (.A2(_0486_),
    .A1(_0484_),
    .B1(_0485_),
    .X(_0488_));
 sg13g2_and2_1 _1234_ (.A(\stop.syn.filt.m1.sum_in2[3] ),
    .B(\stop.syn.filt.m2.sum_in2[3] ),
    .X(_0489_));
 sg13g2_or2_1 _1235_ (.X(_0490_),
    .B(\stop.syn.filt.m2.sum_in2[3] ),
    .A(\stop.syn.filt.m1.sum_in2[3] ));
 sg13g2_nand2b_1 _1236_ (.Y(_0491_),
    .B(_0490_),
    .A_N(_0489_));
 sg13g2_xnor2_1 _1237_ (.Y(_0062_),
    .A(_0488_),
    .B(_0491_));
 sg13g2_nand2_1 _1238_ (.Y(_0492_),
    .A(\stop.syn.filt.m1.sum_in2[4] ),
    .B(\stop.syn.filt.m2.sum_in2[4] ));
 sg13g2_xnor2_1 _1239_ (.Y(_0493_),
    .A(\stop.syn.filt.m1.sum_in2[4] ),
    .B(\stop.syn.filt.m2.sum_in2[4] ));
 sg13g2_a21oi_2 _1240_ (.B1(_0489_),
    .Y(_0494_),
    .A2(_0490_),
    .A1(_0488_));
 sg13g2_xor2_1 _1241_ (.B(_0494_),
    .A(_0493_),
    .X(_0063_));
 sg13g2_or2_1 _1242_ (.X(_0495_),
    .B(\stop.syn.filt.m2.sum_in2[5] ),
    .A(\stop.syn.filt.m1.sum_in2[5] ));
 sg13g2_xnor2_1 _1243_ (.Y(_0496_),
    .A(\stop.syn.filt.m1.sum_in2[5] ),
    .B(\stop.syn.filt.m2.sum_in2[5] ));
 sg13g2_o21ai_1 _1244_ (.B1(_0492_),
    .Y(_0497_),
    .A1(_0493_),
    .A2(_0494_));
 sg13g2_xnor2_1 _1245_ (.Y(_0064_),
    .A(_0496_),
    .B(_0497_));
 sg13g2_nand2_1 _1246_ (.Y(_0498_),
    .A(\stop.syn.filt.m1.sum_in2[6] ),
    .B(\stop.syn.filt.m2.sum_in2[6] ));
 sg13g2_xnor2_1 _1247_ (.Y(_0499_),
    .A(\stop.syn.filt.m1.sum_in2[6] ),
    .B(\stop.syn.filt.m2.sum_in2[6] ));
 sg13g2_inv_1 _1248_ (.Y(_0500_),
    .A(_0499_));
 sg13g2_a22oi_1 _1249_ (.Y(_0501_),
    .B1(\stop.syn.filt.m2.sum_in2[5] ),
    .B2(\stop.syn.filt.m1.sum_in2[5] ),
    .A2(\stop.syn.filt.m2.sum_in2[4] ),
    .A1(\stop.syn.filt.m1.sum_in2[4] ));
 sg13g2_o21ai_1 _1250_ (.B1(_0501_),
    .Y(_0502_),
    .A1(_0493_),
    .A2(_0494_));
 sg13g2_nand2_1 _1251_ (.Y(_0503_),
    .A(_0495_),
    .B(_0502_));
 sg13g2_nand3_1 _1252_ (.B(_0500_),
    .C(_0502_),
    .A(_0495_),
    .Y(_0504_));
 sg13g2_xnor2_1 _1253_ (.Y(_0065_),
    .A(_0500_),
    .B(_0503_));
 sg13g2_and2_1 _1254_ (.A(\stop.syn.filt.m1.sum_in2[7] ),
    .B(\stop.syn.filt.m2.sum_in2[7] ),
    .X(_0505_));
 sg13g2_xnor2_1 _1255_ (.Y(_0506_),
    .A(\stop.syn.filt.m1.sum_in2[7] ),
    .B(\stop.syn.filt.m2.sum_in2[7] ));
 sg13g2_a21oi_1 _1256_ (.A1(_0498_),
    .A2(_0504_),
    .Y(_0507_),
    .B1(_0506_));
 sg13g2_nand3_1 _1257_ (.B(_0504_),
    .C(_0506_),
    .A(_0498_),
    .Y(_0508_));
 sg13g2_nor2b_1 _1258_ (.A(_0507_),
    .B_N(_0508_),
    .Y(_0066_));
 sg13g2_nor2_1 _1259_ (.A(_0505_),
    .B(_0507_),
    .Y(_0509_));
 sg13g2_nand2_1 _1260_ (.Y(_0510_),
    .A(\stop.syn.filt.m1.sum_in2[8] ),
    .B(\stop.syn.filt.m2.sum_in2[8] ));
 sg13g2_xnor2_1 _1261_ (.Y(_0511_),
    .A(\stop.syn.filt.m1.sum_in2[8] ),
    .B(\stop.syn.filt.m2.sum_in2[8] ));
 sg13g2_xor2_1 _1262_ (.B(_0511_),
    .A(_0509_),
    .X(_0067_));
 sg13g2_xnor2_1 _1263_ (.Y(_0512_),
    .A(\stop.syn.filt.m1.sum_in2[9] ),
    .B(\stop.syn.filt.m2.sum_in2[9] ));
 sg13g2_o21ai_1 _1264_ (.B1(_0510_),
    .Y(_0513_),
    .A1(_0509_),
    .A2(_0511_));
 sg13g2_xnor2_1 _1265_ (.Y(_0068_),
    .A(_0512_),
    .B(_0513_));
 sg13g2_nand2_1 _1266_ (.Y(_0514_),
    .A(\stop.syn.filt.m1.sum_in2[10] ),
    .B(\stop.syn.filt.m2.sum_in2[10] ));
 sg13g2_nor2_1 _1267_ (.A(\stop.syn.filt.m1.sum_in2[10] ),
    .B(\stop.syn.filt.m2.sum_in2[10] ),
    .Y(_0515_));
 sg13g2_xor2_1 _1268_ (.B(\stop.syn.filt.m2.sum_in2[10] ),
    .A(\stop.syn.filt.m1.sum_in2[10] ),
    .X(_0516_));
 sg13g2_nor2_1 _1269_ (.A(_0511_),
    .B(_0512_),
    .Y(_0517_));
 sg13g2_o21ai_1 _1270_ (.B1(_0517_),
    .Y(_0518_),
    .A1(_0505_),
    .A2(_0507_));
 sg13g2_a22oi_1 _1271_ (.Y(_0519_),
    .B1(\stop.syn.filt.m2.sum_in2[9] ),
    .B2(\stop.syn.filt.m1.sum_in2[9] ),
    .A2(\stop.syn.filt.m2.sum_in2[8] ),
    .A1(\stop.syn.filt.m1.sum_in2[8] ));
 sg13g2_inv_1 _1272_ (.Y(_0520_),
    .A(_0519_));
 sg13g2_o21ai_1 _1273_ (.B1(_0520_),
    .Y(_0521_),
    .A1(\stop.syn.filt.m1.sum_in2[9] ),
    .A2(\stop.syn.filt.m2.sum_in2[9] ));
 sg13g2_and2_1 _1274_ (.A(_0518_),
    .B(_0521_),
    .X(_0522_));
 sg13g2_xnor2_1 _1275_ (.Y(_0054_),
    .A(_0516_),
    .B(_0522_));
 sg13g2_nor2_1 _1276_ (.A(\stop.syn.filt.m1.sum_in2[11] ),
    .B(\stop.syn.filt.m2.sum_in2[11] ),
    .Y(_0523_));
 sg13g2_nand2_1 _1277_ (.Y(_0524_),
    .A(\stop.syn.filt.m1.sum_in2[11] ),
    .B(\stop.syn.filt.m2.sum_in2[11] ));
 sg13g2_nand2b_1 _1278_ (.Y(_0525_),
    .B(_0524_),
    .A_N(_0523_));
 sg13g2_o21ai_1 _1279_ (.B1(_0514_),
    .Y(_0526_),
    .A1(_0515_),
    .A2(_0522_));
 sg13g2_xnor2_1 _1280_ (.Y(_0055_),
    .A(_0525_),
    .B(_0526_));
 sg13g2_and2_1 _1281_ (.A(\stop.syn.filt.m1.sum_in2[12] ),
    .B(\stop.syn.filt.m2.sum_in2[12] ),
    .X(_0527_));
 sg13g2_xor2_1 _1282_ (.B(\stop.syn.filt.m2.sum_in2[12] ),
    .A(\stop.syn.filt.m1.sum_in2[12] ),
    .X(_0528_));
 sg13g2_nand2_1 _1283_ (.Y(_0529_),
    .A(_0514_),
    .B(_0524_));
 sg13g2_nand2b_1 _1284_ (.Y(_0530_),
    .B(_0529_),
    .A_N(_0523_));
 sg13g2_and2_1 _1285_ (.A(_0521_),
    .B(_0530_),
    .X(_0531_));
 sg13g2_a221oi_1 _1286_ (.B2(_0518_),
    .C1(_0523_),
    .B1(_0531_),
    .A1(_0515_),
    .Y(_0532_),
    .A2(_0524_));
 sg13g2_xor2_1 _1287_ (.B(_0532_),
    .A(_0528_),
    .X(_0056_));
 sg13g2_nand2_1 _1288_ (.Y(_0533_),
    .A(\stop.syn.filt.m1.sum_in2[13] ),
    .B(\stop.syn.filt.m2.sum_in2[13] ));
 sg13g2_xor2_1 _1289_ (.B(\stop.syn.filt.m2.sum_in2[13] ),
    .A(\stop.syn.filt.m1.sum_in2[13] ),
    .X(_0534_));
 sg13g2_a21oi_1 _1290_ (.A1(_0528_),
    .A2(_0532_),
    .Y(_0535_),
    .B1(_0527_));
 sg13g2_xnor2_1 _1291_ (.Y(_0057_),
    .A(_0534_),
    .B(_0535_));
 sg13g2_and2_1 _1292_ (.A(_0528_),
    .B(_0534_),
    .X(_0536_));
 sg13g2_o21ai_1 _1293_ (.B1(_0527_),
    .Y(_0537_),
    .A1(\stop.syn.filt.m1.sum_in2[13] ),
    .A2(\stop.syn.filt.m2.sum_in2[13] ));
 sg13g2_nand2_1 _1294_ (.Y(_0538_),
    .A(_0533_),
    .B(_0537_));
 sg13g2_a21o_1 _1295_ (.A2(_0536_),
    .A1(_0532_),
    .B1(_0538_),
    .X(_0539_));
 sg13g2_and2_1 _1296_ (.A(\stop.syn.filt.m1.sum_in2[14] ),
    .B(\stop.syn.filt.m2.sum_in2[14] ),
    .X(_0540_));
 sg13g2_xor2_1 _1297_ (.B(\stop.syn.filt.m2.sum_in2[14] ),
    .A(\stop.syn.filt.m1.sum_in2[14] ),
    .X(_0541_));
 sg13g2_xor2_1 _1298_ (.B(_0541_),
    .A(_0539_),
    .X(_0058_));
 sg13g2_a21oi_1 _1299_ (.A1(_0539_),
    .A2(_0541_),
    .Y(_0542_),
    .B1(_0540_));
 sg13g2_xor2_1 _1300_ (.B(\stop.syn.filt.m2.sum_in2[15] ),
    .A(\stop.syn.filt.m1.sum_in2[15] ),
    .X(_0543_));
 sg13g2_xnor2_1 _1301_ (.Y(_0059_),
    .A(_0542_),
    .B(_0543_));
 sg13g2_xor2_1 _1302_ (.B(\stop.syn.filt.m2.sum_in2[0] ),
    .A(\stop.syn.filt.m1.sum_in2[0] ),
    .X(_0053_));
 sg13g2_nand3_1 _1303_ (.B(net317),
    .C(\stop.dbg_adsr_reg0 ),
    .A(\stop.syn.filt.m2.sum_in2[0] ),
    .Y(_0544_));
 sg13g2_and3_1 _1304_ (.X(_0545_),
    .A(\stop.syn.filt.m2.sum_in2[1] ),
    .B(\stop.syn.adsr_data_reg[1] ),
    .C(net317));
 sg13g2_nand3_1 _1305_ (.B(\stop.syn.adsr_data_reg[1] ),
    .C(net317),
    .A(\stop.syn.filt.m2.sum_in2[1] ),
    .Y(_0546_));
 sg13g2_a21oi_1 _1306_ (.A1(\stop.syn.adsr_data_reg[1] ),
    .A2(net317),
    .Y(_0547_),
    .B1(\stop.syn.filt.m2.sum_in2[1] ));
 sg13g2_nor2_1 _1307_ (.A(_0545_),
    .B(_0547_),
    .Y(_0548_));
 sg13g2_xnor2_1 _1308_ (.Y(\stop.syn.filt.m2.sum[1] ),
    .A(_0544_),
    .B(_0548_));
 sg13g2_o21ai_1 _1309_ (.B1(_0546_),
    .Y(_0549_),
    .A1(_0544_),
    .A2(_0547_));
 sg13g2_and3_1 _1310_ (.X(_0550_),
    .A(\stop.syn.filt.m2.sum_in2[2] ),
    .B(net317),
    .C(\stop.syn.adsr_data_reg[2] ));
 sg13g2_a21o_1 _1311_ (.A2(\stop.syn.adsr_data_reg[2] ),
    .A1(net317),
    .B1(\stop.syn.filt.m2.sum_in2[2] ),
    .X(_0551_));
 sg13g2_nand2b_1 _1312_ (.Y(_0552_),
    .B(_0551_),
    .A_N(_0550_));
 sg13g2_xnor2_1 _1313_ (.Y(\stop.syn.filt.m2.sum[2] ),
    .A(_0549_),
    .B(_0552_));
 sg13g2_nand2_1 _1314_ (.Y(_0553_),
    .A(net316),
    .B(\stop.syn.adsr_data_reg[3] ));
 sg13g2_nor2_1 _1315_ (.A(_0050_),
    .B(_0553_),
    .Y(_0554_));
 sg13g2_xor2_1 _1316_ (.B(_0553_),
    .A(_0050_),
    .X(_0555_));
 sg13g2_a21o_1 _1317_ (.A2(_0551_),
    .A1(_0549_),
    .B1(_0550_),
    .X(_0556_));
 sg13g2_xor2_1 _1318_ (.B(_0556_),
    .A(_0555_),
    .X(\stop.syn.filt.m2.sum[3] ));
 sg13g2_a21oi_2 _1319_ (.B1(_0554_),
    .Y(_0557_),
    .A2(_0556_),
    .A1(_0555_));
 sg13g2_nand3_1 _1320_ (.B(net316),
    .C(\stop.syn.adsr_data_reg[4] ),
    .A(\stop.syn.filt.m2.sum_in2[4] ),
    .Y(_0558_));
 sg13g2_a21o_1 _1321_ (.A2(\stop.syn.adsr_data_reg[4] ),
    .A1(net316),
    .B1(\stop.syn.filt.m2.sum_in2[4] ),
    .X(_0559_));
 sg13g2_nand2_1 _1322_ (.Y(_0560_),
    .A(_0558_),
    .B(_0559_));
 sg13g2_xor2_1 _1323_ (.B(_0560_),
    .A(_0557_),
    .X(\stop.syn.filt.m2.sum[4] ));
 sg13g2_nand2_1 _1324_ (.Y(_0561_),
    .A(net317),
    .B(\stop.syn.adsr_data_reg[5] ));
 sg13g2_nor2_1 _1325_ (.A(_0051_),
    .B(_0561_),
    .Y(_0562_));
 sg13g2_xor2_1 _1326_ (.B(_0561_),
    .A(_0051_),
    .X(_0563_));
 sg13g2_o21ai_1 _1327_ (.B1(_0558_),
    .Y(_0564_),
    .A1(_0557_),
    .A2(_0560_));
 sg13g2_xor2_1 _1328_ (.B(_0564_),
    .A(_0563_),
    .X(\stop.syn.filt.m2.sum[5] ));
 sg13g2_and3_1 _1329_ (.X(_0565_),
    .A(\stop.syn.filt.m2.sum_in2[6] ),
    .B(net316),
    .C(\stop.syn.adsr_data_reg[6] ));
 sg13g2_a21oi_1 _1330_ (.A1(net316),
    .A2(\stop.syn.adsr_data_reg[6] ),
    .Y(_0566_),
    .B1(\stop.syn.filt.m2.sum_in2[6] ));
 sg13g2_nor2_1 _1331_ (.A(_0565_),
    .B(_0566_),
    .Y(_0567_));
 sg13g2_a21oi_1 _1332_ (.A1(_0051_),
    .A2(_0561_),
    .Y(_0568_),
    .B1(_0558_));
 sg13g2_nor2_1 _1333_ (.A(_0562_),
    .B(_0568_),
    .Y(_0569_));
 sg13g2_nand2b_1 _1334_ (.Y(_0570_),
    .B(_0563_),
    .A_N(_0560_));
 sg13g2_o21ai_1 _1335_ (.B1(_0569_),
    .Y(_0571_),
    .A1(_0557_),
    .A2(_0570_));
 sg13g2_xor2_1 _1336_ (.B(_0571_),
    .A(_0567_),
    .X(\stop.syn.filt.m2.sum[6] ));
 sg13g2_a21oi_1 _1337_ (.A1(_0567_),
    .A2(_0571_),
    .Y(_0572_),
    .B1(_0565_));
 sg13g2_nand3_1 _1338_ (.B(net316),
    .C(\stop.syn.adsr_data_reg[7] ),
    .A(\stop.syn.filt.m2.sum_in2[7] ),
    .Y(_0573_));
 sg13g2_a21o_1 _1339_ (.A2(\stop.syn.adsr_data_reg[7] ),
    .A1(net316),
    .B1(\stop.syn.filt.m2.sum_in2[7] ),
    .X(_0574_));
 sg13g2_nand2_1 _1340_ (.Y(_0575_),
    .A(_0573_),
    .B(_0574_));
 sg13g2_xor2_1 _1341_ (.B(_0575_),
    .A(_0572_),
    .X(\stop.syn.filt.m2.sum[7] ));
 sg13g2_o21ai_1 _1342_ (.B1(_0573_),
    .Y(_0576_),
    .A1(_0572_),
    .A2(_0575_));
 sg13g2_inv_1 _1343_ (.Y(_0577_),
    .A(_0576_));
 sg13g2_nand3_1 _1344_ (.B(net318),
    .C(\stop.syn.adsr_data_reg[8] ),
    .A(\stop.syn.filt.m2.sum_in2[8] ),
    .Y(_0578_));
 sg13g2_a21o_1 _1345_ (.A2(\stop.syn.adsr_data_reg[8] ),
    .A1(net318),
    .B1(\stop.syn.filt.m2.sum_in2[8] ),
    .X(_0579_));
 sg13g2_nand2_1 _1346_ (.Y(_0580_),
    .A(_0578_),
    .B(_0579_));
 sg13g2_xnor2_1 _1347_ (.Y(\stop.syn.filt.m2.sum[8] ),
    .A(_0576_),
    .B(_0580_));
 sg13g2_nand2_1 _1348_ (.Y(_0581_),
    .A(net316),
    .B(\stop.syn.adsr_data_reg[9] ));
 sg13g2_xor2_1 _1349_ (.B(_0581_),
    .A(_0052_),
    .X(_0582_));
 sg13g2_o21ai_1 _1350_ (.B1(_0578_),
    .Y(_0583_),
    .A1(_0577_),
    .A2(_0580_));
 sg13g2_xor2_1 _1351_ (.B(_0583_),
    .A(_0582_),
    .X(\stop.syn.filt.m2.sum[9] ));
 sg13g2_nand3_1 _1352_ (.B(net315),
    .C(\stop.syn.adsr_data_reg[10] ),
    .A(\stop.syn.filt.m2.sum_in2[10] ),
    .Y(_0584_));
 sg13g2_a21o_1 _1353_ (.A2(\stop.syn.adsr_data_reg[10] ),
    .A1(net315),
    .B1(\stop.syn.filt.m2.sum_in2[10] ),
    .X(_0585_));
 sg13g2_nand2_1 _1354_ (.Y(_0586_),
    .A(_0584_),
    .B(_0585_));
 sg13g2_a21o_1 _1355_ (.A2(_0581_),
    .A1(_0052_),
    .B1(_0578_),
    .X(_0587_));
 sg13g2_o21ai_1 _1356_ (.B1(_0587_),
    .Y(_0588_),
    .A1(_0052_),
    .A2(_0581_));
 sg13g2_nor2b_1 _1357_ (.A(_0580_),
    .B_N(_0582_),
    .Y(_0589_));
 sg13g2_a21oi_1 _1358_ (.A1(_0576_),
    .A2(_0589_),
    .Y(_0590_),
    .B1(_0588_));
 sg13g2_xor2_1 _1359_ (.B(_0590_),
    .A(_0586_),
    .X(\stop.syn.filt.m2.sum[10] ));
 sg13g2_a21oi_1 _1360_ (.A1(net315),
    .A2(\stop.syn.adsr_data_reg[11] ),
    .Y(_0591_),
    .B1(\stop.syn.filt.m2.sum_in2[11] ));
 sg13g2_nand3_1 _1361_ (.B(net314),
    .C(\stop.syn.adsr_data_reg[11] ),
    .A(\stop.syn.filt.m2.sum_in2[11] ),
    .Y(_0592_));
 sg13g2_nand2b_1 _1362_ (.Y(_0593_),
    .B(_0592_),
    .A_N(_0591_));
 sg13g2_o21ai_1 _1363_ (.B1(_0584_),
    .Y(_0594_),
    .A1(_0586_),
    .A2(_0590_));
 sg13g2_xnor2_1 _1364_ (.Y(\stop.syn.filt.m2.sum[11] ),
    .A(_0593_),
    .B(_0594_));
 sg13g2_nor2_1 _1365_ (.A(_0586_),
    .B(_0593_),
    .Y(_0595_));
 sg13g2_and2_1 _1366_ (.A(_0589_),
    .B(_0595_),
    .X(_0596_));
 sg13g2_o21ai_1 _1367_ (.B1(_0592_),
    .Y(_0597_),
    .A1(_0584_),
    .A2(_0591_));
 sg13g2_a221oi_1 _1368_ (.B2(_0576_),
    .C1(_0597_),
    .B1(_0596_),
    .A1(_0588_),
    .Y(_0598_),
    .A2(_0595_));
 sg13g2_nand3_1 _1369_ (.B(net314),
    .C(\stop.syn.adsr_data_reg[12] ),
    .A(\stop.syn.filt.m2.sum_in2[12] ),
    .Y(_0599_));
 sg13g2_a21o_1 _1370_ (.A2(\stop.syn.adsr_data_reg[12] ),
    .A1(net314),
    .B1(\stop.syn.filt.m2.sum_in2[12] ),
    .X(_0600_));
 sg13g2_nand2_1 _1371_ (.Y(_0601_),
    .A(_0599_),
    .B(_0600_));
 sg13g2_xor2_1 _1372_ (.B(_0601_),
    .A(_0598_),
    .X(\stop.syn.filt.m2.sum[12] ));
 sg13g2_nand2_1 _1373_ (.Y(_0602_),
    .A(net314),
    .B(\stop.syn.adsr_data_reg[13] ));
 sg13g2_nor2_1 _1374_ (.A(_0042_),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_xor2_1 _1375_ (.B(_0602_),
    .A(_0042_),
    .X(_0604_));
 sg13g2_o21ai_1 _1376_ (.B1(_0599_),
    .Y(_0605_),
    .A1(_0598_),
    .A2(_0601_));
 sg13g2_xor2_1 _1377_ (.B(_0605_),
    .A(_0604_),
    .X(\stop.syn.filt.m2.sum[13] ));
 sg13g2_nand2b_1 _1378_ (.Y(_0606_),
    .B(_0604_),
    .A_N(_0601_));
 sg13g2_a21oi_1 _1379_ (.A1(_0042_),
    .A2(_0602_),
    .Y(_0607_),
    .B1(_0599_));
 sg13g2_nor2_1 _1380_ (.A(_0603_),
    .B(_0607_),
    .Y(_0608_));
 sg13g2_o21ai_1 _1381_ (.B1(_0608_),
    .Y(_0609_),
    .A1(_0598_),
    .A2(_0606_));
 sg13g2_nand3_1 _1382_ (.B(net314),
    .C(\stop.syn.adsr_data_reg[14] ),
    .A(\stop.syn.filt.m2.sum_in2[14] ),
    .Y(_0610_));
 sg13g2_a21o_1 _1383_ (.A2(\stop.syn.adsr_data_reg[14] ),
    .A1(net314),
    .B1(\stop.syn.filt.m2.sum_in2[14] ),
    .X(_0611_));
 sg13g2_nand2_1 _1384_ (.Y(_0612_),
    .A(_0610_),
    .B(_0611_));
 sg13g2_nand2b_1 _1385_ (.Y(_0613_),
    .B(_0609_),
    .A_N(_0612_));
 sg13g2_xnor2_1 _1386_ (.Y(\stop.syn.filt.m2.sum[14] ),
    .A(_0609_),
    .B(_0612_));
 sg13g2_and3_1 _1387_ (.X(_0614_),
    .A(\stop.syn.filt.m2.sum_in2[15] ),
    .B(net314),
    .C(\stop.syn.adsr_data_reg[15] ));
 sg13g2_a21oi_1 _1388_ (.A1(net314),
    .A2(\stop.syn.adsr_data_reg[15] ),
    .Y(_0615_),
    .B1(\stop.syn.filt.m2.sum_in2[15] ));
 sg13g2_nor2_1 _1389_ (.A(_0614_),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_nand2_1 _1390_ (.Y(_0617_),
    .A(_0610_),
    .B(_0613_));
 sg13g2_xor2_1 _1391_ (.B(_0617_),
    .A(_0616_),
    .X(\stop.syn.filt.m2.sum[15] ));
 sg13g2_nand3_1 _1392_ (.B(net308),
    .C(\stop.syn.adsr_data[8] ),
    .A(\stop.dbg_osc0 ),
    .Y(_0618_));
 sg13g2_a21o_1 _1393_ (.A2(net308),
    .A1(\stop.dbg_osc0 ),
    .B1(\stop.syn.adsr_data[8] ),
    .X(_0619_));
 sg13g2_and2_1 _1394_ (.A(_0618_),
    .B(_0619_),
    .X(_0070_));
 sg13g2_and3_1 _1395_ (.X(_0620_),
    .A(\stop.syn.osc_data[1] ),
    .B(net308),
    .C(\stop.syn.adsr_data[9] ));
 sg13g2_nand3_1 _1396_ (.B(net308),
    .C(\stop.syn.adsr_data[9] ),
    .A(\stop.syn.osc_data[1] ),
    .Y(_0621_));
 sg13g2_a21oi_1 _1397_ (.A1(\stop.syn.osc_data[1] ),
    .A2(net308),
    .Y(_0622_),
    .B1(\stop.syn.adsr_data[9] ));
 sg13g2_nor2_1 _1398_ (.A(_0620_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_xnor2_1 _1399_ (.Y(_0071_),
    .A(_0618_),
    .B(_0623_));
 sg13g2_o21ai_1 _1400_ (.B1(_0621_),
    .Y(_0624_),
    .A1(_0618_),
    .A2(_0622_));
 sg13g2_inv_1 _1401_ (.Y(_0625_),
    .A(_0624_));
 sg13g2_nand3_1 _1402_ (.B(net308),
    .C(\stop.syn.adsr_data[10] ),
    .A(\stop.syn.osc_data[2] ),
    .Y(_0626_));
 sg13g2_a21o_1 _1403_ (.A2(net308),
    .A1(\stop.syn.osc_data[2] ),
    .B1(\stop.syn.adsr_data[10] ),
    .X(_0627_));
 sg13g2_nand2_1 _1404_ (.Y(_0628_),
    .A(_0626_),
    .B(_0627_));
 sg13g2_xnor2_1 _1405_ (.Y(_0072_),
    .A(_0624_),
    .B(_0628_));
 sg13g2_o21ai_1 _1406_ (.B1(_0626_),
    .Y(_0629_),
    .A1(_0625_),
    .A2(_0628_));
 sg13g2_nand2_1 _1407_ (.Y(_0630_),
    .A(\stop.syn.osc_data[3] ),
    .B(net307));
 sg13g2_nor2_1 _1408_ (.A(_0043_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_xor2_1 _1409_ (.B(_0630_),
    .A(_0043_),
    .X(_0632_));
 sg13g2_xor2_1 _1410_ (.B(_0632_),
    .A(_0629_),
    .X(_0073_));
 sg13g2_a21oi_1 _1411_ (.A1(_0629_),
    .A2(_0632_),
    .Y(_0633_),
    .B1(_0631_));
 sg13g2_nand3_1 _1412_ (.B(net307),
    .C(\stop.syn.adsr_data[12] ),
    .A(\stop.syn.osc_data[4] ),
    .Y(_0634_));
 sg13g2_a21o_1 _1413_ (.A2(net307),
    .A1(\stop.syn.osc_data[4] ),
    .B1(\stop.syn.adsr_data[12] ),
    .X(_0635_));
 sg13g2_nand2_1 _1414_ (.Y(_0636_),
    .A(_0634_),
    .B(_0635_));
 sg13g2_xor2_1 _1415_ (.B(_0636_),
    .A(_0633_),
    .X(_0074_));
 sg13g2_o21ai_1 _1416_ (.B1(_0634_),
    .Y(_0637_),
    .A1(_0633_),
    .A2(_0636_));
 sg13g2_nand2_1 _1417_ (.Y(_0638_),
    .A(\stop.syn.osc_data[5] ),
    .B(net307));
 sg13g2_nor2_1 _1418_ (.A(_0044_),
    .B(_0638_),
    .Y(_0639_));
 sg13g2_xor2_1 _1419_ (.B(_0638_),
    .A(_0044_),
    .X(_0640_));
 sg13g2_xor2_1 _1420_ (.B(_0640_),
    .A(_0637_),
    .X(_0075_));
 sg13g2_a21oi_1 _1421_ (.A1(_0637_),
    .A2(_0640_),
    .Y(_0641_),
    .B1(_0639_));
 sg13g2_nand3_1 _1422_ (.B(net307),
    .C(\stop.syn.adsr_data[14] ),
    .A(\stop.syn.osc_data[6] ),
    .Y(_0642_));
 sg13g2_a21o_1 _1423_ (.A2(net307),
    .A1(\stop.syn.osc_data[6] ),
    .B1(\stop.syn.adsr_data[14] ),
    .X(_0643_));
 sg13g2_nand2_1 _1424_ (.Y(_0644_),
    .A(_0642_),
    .B(_0643_));
 sg13g2_xor2_1 _1425_ (.B(_0644_),
    .A(_0641_),
    .X(_0076_));
 sg13g2_o21ai_1 _1426_ (.B1(_0642_),
    .Y(_0645_),
    .A1(_0641_),
    .A2(_0644_));
 sg13g2_inv_1 _1427_ (.Y(_0646_),
    .A(_0645_));
 sg13g2_nand3_1 _1428_ (.B(net307),
    .C(\stop.syn.adsr_data[15] ),
    .A(\stop.syn.osc_data[7] ),
    .Y(_0647_));
 sg13g2_a21o_1 _1429_ (.A2(net307),
    .A1(\stop.syn.osc_data[7] ),
    .B1(\stop.syn.adsr_data[15] ),
    .X(_0648_));
 sg13g2_nand2_1 _1430_ (.Y(_0649_),
    .A(_0647_),
    .B(_0648_));
 sg13g2_xnor2_1 _1431_ (.Y(_0077_),
    .A(_0645_),
    .B(_0649_));
 sg13g2_a21oi_1 _1432_ (.A1(_0476_),
    .A2(_0479_),
    .Y(\stop.syn.filt.m1.sum[16] ),
    .B1(_0477_));
 sg13g2_a21oi_1 _1433_ (.A1(_0610_),
    .A2(_0613_),
    .Y(_0650_),
    .B1(_0615_));
 sg13g2_or2_1 _1434_ (.X(\stop.syn.filt.m2.sum[16] ),
    .B(_0650_),
    .A(_0614_));
 sg13g2_o21ai_1 _1435_ (.B1(_0647_),
    .Y(_0069_),
    .A1(_0646_),
    .A2(_0649_));
 sg13g2_nand2b_1 _1436_ (.Y(\stop.syn.clki.arstn ),
    .B(net134),
    .A_N(\stop.syn.rstn_fst_reg1 ));
 sg13g2_o21ai_1 _1437_ (.B1(net370),
    .Y(_0651_),
    .A1(net2),
    .A2(\stop.ctrl.first_bit_reg ));
 sg13g2_inv_1 _1438_ (.Y(\stop.dbg_rstn ),
    .A(_0651_));
 sg13g2_or2_1 _1439_ (.X(\stop.dbg_trig ),
    .B(net1),
    .A(\stop.ctrl.trig ));
 sg13g2_nor2_1 _1440_ (.A(_0080_),
    .B(net2),
    .Y(_0652_));
 sg13g2_mux2_1 _1441_ (.A0(\stop.ctrl.trig ),
    .A1(net3),
    .S(_0652_),
    .X(_0133_));
 sg13g2_or2_1 _1442_ (.X(_0653_),
    .B(\stop.syn.osci.counter[0] ),
    .A(\stop.ctrl.cfg[32] ));
 sg13g2_nand2_2 _1443_ (.Y(_0654_),
    .A(\stop.ctrl.cfg[32] ),
    .B(\stop.syn.osci.counter[0] ));
 sg13g2_and3_1 _1444_ (.X(_0134_),
    .A(\stop.syn.adsri.rstn ),
    .B(_0653_),
    .C(_0654_));
 sg13g2_nand2_1 _1445_ (.Y(_0655_),
    .A(\stop.ctrl.cfg[33] ),
    .B(\stop.syn.osci.counter[1] ));
 sg13g2_xnor2_1 _1446_ (.Y(_0656_),
    .A(\stop.ctrl.cfg[33] ),
    .B(\stop.syn.osci.counter[1] ));
 sg13g2_o21ai_1 _1447_ (.B1(net277),
    .Y(_0657_),
    .A1(_0654_),
    .A2(_0656_));
 sg13g2_a21oi_1 _1448_ (.A1(_0654_),
    .A2(_0656_),
    .Y(_0135_),
    .B1(_0657_));
 sg13g2_and2_1 _1449_ (.A(\stop.ctrl.cfg[34] ),
    .B(\stop.syn.osci.counter[2] ),
    .X(_0658_));
 sg13g2_xor2_1 _1450_ (.B(\stop.syn.osci.counter[2] ),
    .A(\stop.ctrl.cfg[34] ),
    .X(_0659_));
 sg13g2_o21ai_1 _1451_ (.B1(_0655_),
    .Y(_0660_),
    .A1(_0654_),
    .A2(_0656_));
 sg13g2_nor2_1 _1452_ (.A(_0659_),
    .B(_0660_),
    .Y(_0661_));
 sg13g2_a21oi_1 _1453_ (.A1(_0659_),
    .A2(_0660_),
    .Y(_0662_),
    .B1(_0320_));
 sg13g2_nor2b_1 _1454_ (.A(_0661_),
    .B_N(_0662_),
    .Y(_0136_));
 sg13g2_nand2_1 _1455_ (.Y(_0663_),
    .A(\stop.ctrl.cfg[35] ),
    .B(\stop.syn.osci.counter[3] ));
 sg13g2_xnor2_1 _1456_ (.Y(_0664_),
    .A(\stop.ctrl.cfg[35] ),
    .B(\stop.syn.osci.counter[3] ));
 sg13g2_a21oi_2 _1457_ (.B1(_0658_),
    .Y(_0665_),
    .A2(_0660_),
    .A1(_0659_));
 sg13g2_o21ai_1 _1458_ (.B1(net277),
    .Y(_0666_),
    .A1(_0664_),
    .A2(_0665_));
 sg13g2_a21oi_1 _1459_ (.A1(_0664_),
    .A2(_0665_),
    .Y(_0137_),
    .B1(_0666_));
 sg13g2_and2_1 _1460_ (.A(\stop.ctrl.cfg[36] ),
    .B(\stop.dbg_osc0 ),
    .X(_0667_));
 sg13g2_xor2_1 _1461_ (.B(\stop.dbg_osc0 ),
    .A(\stop.ctrl.cfg[36] ),
    .X(_0668_));
 sg13g2_o21ai_1 _1462_ (.B1(_0663_),
    .Y(_0669_),
    .A1(_0664_),
    .A2(_0665_));
 sg13g2_or2_1 _1463_ (.X(_0670_),
    .B(_0669_),
    .A(_0668_));
 sg13g2_a21oi_1 _1464_ (.A1(_0668_),
    .A2(_0669_),
    .Y(_0671_),
    .B1(_0320_));
 sg13g2_and2_1 _1465_ (.A(_0670_),
    .B(_0671_),
    .X(_0138_));
 sg13g2_a21oi_1 _1466_ (.A1(_0668_),
    .A2(_0669_),
    .Y(_0672_),
    .B1(_0667_));
 sg13g2_nor2_1 _1467_ (.A(\stop.ctrl.cfg[37] ),
    .B(\stop.syn.osc_data[1] ),
    .Y(_0673_));
 sg13g2_and2_1 _1468_ (.A(\stop.ctrl.cfg[37] ),
    .B(\stop.syn.osc_data[1] ),
    .X(_0674_));
 sg13g2_nor3_1 _1469_ (.A(_0672_),
    .B(_0673_),
    .C(_0674_),
    .Y(_0675_));
 sg13g2_o21ai_1 _1470_ (.B1(_0672_),
    .Y(_0676_),
    .A1(_0673_),
    .A2(_0674_));
 sg13g2_nand2_1 _1471_ (.Y(_0677_),
    .A(net277),
    .B(_0676_));
 sg13g2_nor2_1 _1472_ (.A(_0675_),
    .B(_0677_),
    .Y(_0139_));
 sg13g2_nand2_1 _1473_ (.Y(_0678_),
    .A(\stop.ctrl.cfg[38] ),
    .B(\stop.syn.osc_data[2] ));
 sg13g2_xnor2_1 _1474_ (.Y(_0679_),
    .A(\stop.ctrl.cfg[38] ),
    .B(\stop.syn.osc_data[2] ));
 sg13g2_a221oi_1 _1475_ (.B2(_0669_),
    .C1(_0667_),
    .B1(_0668_),
    .A1(\stop.ctrl.cfg[37] ),
    .Y(_0680_),
    .A2(\stop.syn.osc_data[1] ));
 sg13g2_o21ai_1 _1476_ (.B1(_0679_),
    .Y(_0681_),
    .A1(_0673_),
    .A2(_0680_));
 sg13g2_or3_1 _1477_ (.A(_0673_),
    .B(_0679_),
    .C(_0680_),
    .X(_0682_));
 sg13g2_and3_1 _1478_ (.X(_0140_),
    .A(net277),
    .B(_0681_),
    .C(_0682_));
 sg13g2_xnor2_1 _1479_ (.Y(_0683_),
    .A(\stop.ctrl.cfg[39] ),
    .B(\stop.syn.osc_data[3] ));
 sg13g2_and2_1 _1480_ (.A(_0678_),
    .B(_0682_),
    .X(_0684_));
 sg13g2_a21oi_1 _1481_ (.A1(_0678_),
    .A2(_0682_),
    .Y(_0685_),
    .B1(_0683_));
 sg13g2_a21oi_1 _1482_ (.A1(_0683_),
    .A2(_0684_),
    .Y(_0686_),
    .B1(_0320_));
 sg13g2_nor2b_1 _1483_ (.A(_0685_),
    .B_N(_0686_),
    .Y(_0141_));
 sg13g2_a21oi_2 _1484_ (.B1(_0685_),
    .Y(_0687_),
    .A2(\stop.syn.osc_data[3] ),
    .A1(\stop.ctrl.cfg[39] ));
 sg13g2_nand2_1 _1485_ (.Y(_0688_),
    .A(\stop.ctrl.cfg[40] ),
    .B(\stop.syn.osc_data[4] ));
 sg13g2_xnor2_1 _1486_ (.Y(_0689_),
    .A(\stop.ctrl.cfg[40] ),
    .B(\stop.syn.osc_data[4] ));
 sg13g2_o21ai_1 _1487_ (.B1(net277),
    .Y(_0690_),
    .A1(_0687_),
    .A2(_0689_));
 sg13g2_a21oi_1 _1488_ (.A1(_0687_),
    .A2(_0689_),
    .Y(_0142_),
    .B1(_0690_));
 sg13g2_nor2_1 _1489_ (.A(\stop.ctrl.cfg[41] ),
    .B(\stop.syn.osc_data[5] ),
    .Y(_0691_));
 sg13g2_nand2_1 _1490_ (.Y(_0692_),
    .A(\stop.ctrl.cfg[41] ),
    .B(\stop.syn.osc_data[5] ));
 sg13g2_nor2b_1 _1491_ (.A(_0691_),
    .B_N(_0692_),
    .Y(_0693_));
 sg13g2_inv_1 _1492_ (.Y(_0694_),
    .A(_0693_));
 sg13g2_o21ai_1 _1493_ (.B1(_0688_),
    .Y(_0695_),
    .A1(_0687_),
    .A2(_0689_));
 sg13g2_o21ai_1 _1494_ (.B1(net277),
    .Y(_0696_),
    .A1(_0693_),
    .A2(_0695_));
 sg13g2_a21oi_1 _1495_ (.A1(_0693_),
    .A2(_0695_),
    .Y(_0143_),
    .B1(_0696_));
 sg13g2_nand2_1 _1496_ (.Y(_0697_),
    .A(\stop.ctrl.cfg[42] ),
    .B(\stop.syn.osc_data[6] ));
 sg13g2_xor2_1 _1497_ (.B(\stop.syn.osc_data[6] ),
    .A(\stop.ctrl.cfg[42] ),
    .X(_0698_));
 sg13g2_o21ai_1 _1498_ (.B1(_0692_),
    .Y(_0699_),
    .A1(_0688_),
    .A2(_0691_));
 sg13g2_nor3_1 _1499_ (.A(_0687_),
    .B(_0689_),
    .C(_0694_),
    .Y(_0700_));
 sg13g2_nor3_1 _1500_ (.A(_0698_),
    .B(_0699_),
    .C(_0700_),
    .Y(_0701_));
 sg13g2_o21ai_1 _1501_ (.B1(_0698_),
    .Y(_0702_),
    .A1(_0699_),
    .A2(_0700_));
 sg13g2_nand2_1 _1502_ (.Y(_0703_),
    .A(net277),
    .B(_0702_));
 sg13g2_nor2_1 _1503_ (.A(_0701_),
    .B(_0703_),
    .Y(_0144_));
 sg13g2_xnor2_1 _1504_ (.Y(_0704_),
    .A(\stop.ctrl.cfg[43] ),
    .B(\stop.syn.osc_data[7] ));
 sg13g2_and3_1 _1505_ (.X(_0705_),
    .A(_0697_),
    .B(_0702_),
    .C(_0704_));
 sg13g2_a21oi_1 _1506_ (.A1(_0697_),
    .A2(_0702_),
    .Y(_0706_),
    .B1(_0704_));
 sg13g2_nor3_1 _1507_ (.A(_0320_),
    .B(_0705_),
    .C(_0706_),
    .Y(_0145_));
 sg13g2_nand2_1 _1508_ (.Y(_0707_),
    .A(_0318_),
    .B(_0393_));
 sg13g2_o21ai_1 _1509_ (.B1(net281),
    .Y(_0708_),
    .A1(_0403_),
    .A2(_0707_));
 sg13g2_or4_2 _1510_ (.A(net283),
    .B(_0319_),
    .C(_0394_),
    .D(_0707_),
    .X(_0709_));
 sg13g2_a21oi_1 _1511_ (.A1(_0382_),
    .A2(_0709_),
    .Y(_0146_),
    .B1(_0708_));
 sg13g2_a21oi_1 _1512_ (.A1(_0379_),
    .A2(_0709_),
    .Y(_0147_),
    .B1(_0708_));
 sg13g2_a21oi_1 _1513_ (.A1(_0377_),
    .A2(_0709_),
    .Y(_0148_),
    .B1(_0708_));
 sg13g2_a21oi_1 _1514_ (.A1(_0376_),
    .A2(_0709_),
    .Y(_0149_),
    .B1(_0708_));
 sg13g2_a21oi_1 _1515_ (.A1(_0374_),
    .A2(_0709_),
    .Y(_0150_),
    .B1(_0708_));
 sg13g2_a21oi_1 _1516_ (.A1(_0373_),
    .A2(_0709_),
    .Y(_0151_),
    .B1(_0708_));
 sg13g2_a21oi_1 _1517_ (.A1(_0372_),
    .A2(_0709_),
    .Y(_0152_),
    .B1(_0708_));
 sg13g2_a21oi_1 _1518_ (.A1(_0370_),
    .A2(_0709_),
    .Y(_0153_),
    .B1(_0708_));
 sg13g2_or2_1 _1519_ (.X(_0710_),
    .B(net109),
    .A(\stop.dbg_adsr_filt0 ));
 sg13g2_nand2_1 _1520_ (.Y(_0711_),
    .A(\stop.dbg_adsr_filt0 ),
    .B(net109));
 sg13g2_and3_1 _1521_ (.X(_0156_),
    .A(net278),
    .B(_0710_),
    .C(_0711_));
 sg13g2_nand2_1 _1522_ (.Y(_0712_),
    .A(\stop.syn.daci.din[1] ),
    .B(\stop.syn.daci.accumulator[1] ));
 sg13g2_xnor2_1 _1523_ (.Y(_0713_),
    .A(\stop.syn.daci.din[1] ),
    .B(\stop.syn.daci.accumulator[1] ));
 sg13g2_o21ai_1 _1524_ (.B1(net279),
    .Y(_0714_),
    .A1(_0711_),
    .A2(_0713_));
 sg13g2_a21oi_1 _1525_ (.A1(_0711_),
    .A2(_0713_),
    .Y(_0157_),
    .B1(_0714_));
 sg13g2_and2_1 _1526_ (.A(\stop.syn.daci.din[2] ),
    .B(net133),
    .X(_0715_));
 sg13g2_xor2_1 _1527_ (.B(net124),
    .A(\stop.syn.daci.din[2] ),
    .X(_0716_));
 sg13g2_o21ai_1 _1528_ (.B1(_0712_),
    .Y(_0717_),
    .A1(_0711_),
    .A2(_0713_));
 sg13g2_nor2_1 _1529_ (.A(_0716_),
    .B(_0717_),
    .Y(_0718_));
 sg13g2_a21oi_1 _1530_ (.A1(_0716_),
    .A2(_0717_),
    .Y(_0719_),
    .B1(_0320_));
 sg13g2_nor2b_1 _1531_ (.A(net125),
    .B_N(_0719_),
    .Y(_0158_));
 sg13g2_nand2_1 _1532_ (.Y(_0720_),
    .A(\stop.syn.daci.din[3] ),
    .B(\stop.syn.daci.accumulator[3] ));
 sg13g2_xnor2_1 _1533_ (.Y(_0233_),
    .A(\stop.syn.daci.din[3] ),
    .B(net128));
 sg13g2_a21oi_1 _1534_ (.A1(_0716_),
    .A2(_0717_),
    .Y(_0234_),
    .B1(_0715_));
 sg13g2_nor2_1 _1535_ (.A(_0233_),
    .B(_0234_),
    .Y(_0235_));
 sg13g2_a21oi_1 _1536_ (.A1(_0233_),
    .A2(_0234_),
    .Y(_0236_),
    .B1(_0320_));
 sg13g2_nor2b_1 _1537_ (.A(_0235_),
    .B_N(_0236_),
    .Y(_0159_));
 sg13g2_a21oi_1 _1538_ (.A1(\stop.syn.daci.din[3] ),
    .A2(net128),
    .Y(_0237_),
    .B1(_0235_));
 sg13g2_o21ai_1 _1539_ (.B1(_0720_),
    .Y(_0238_),
    .A1(_0233_),
    .A2(_0234_));
 sg13g2_xnor2_1 _1540_ (.Y(_0239_),
    .A(\stop.syn.daci.din[4] ),
    .B(\stop.syn.daci.accumulator[4] ));
 sg13g2_nor2_1 _1541_ (.A(_0237_),
    .B(_0239_),
    .Y(_0240_));
 sg13g2_a21oi_1 _1542_ (.A1(_0237_),
    .A2(_0239_),
    .Y(_0241_),
    .B1(_0320_));
 sg13g2_nor2b_1 _1543_ (.A(net129),
    .B_N(_0241_),
    .Y(_0160_));
 sg13g2_or2_1 _1544_ (.X(_0242_),
    .B(\stop.syn.daci.accumulator[5] ),
    .A(\stop.syn.daci.din[5] ));
 sg13g2_xnor2_1 _1545_ (.Y(_0243_),
    .A(\stop.syn.daci.din[5] ),
    .B(net121));
 sg13g2_a21oi_1 _1546_ (.A1(\stop.syn.daci.din[4] ),
    .A2(\stop.syn.daci.accumulator[4] ),
    .Y(_0244_),
    .B1(_0240_));
 sg13g2_o21ai_1 _1547_ (.B1(net279),
    .Y(_0245_),
    .A1(_0243_),
    .A2(_0244_));
 sg13g2_a21oi_1 _1548_ (.A1(_0243_),
    .A2(_0244_),
    .Y(_0161_),
    .B1(_0245_));
 sg13g2_nand2_1 _1549_ (.Y(_0246_),
    .A(\stop.syn.daci.din[6] ),
    .B(net123));
 sg13g2_xnor2_1 _1550_ (.Y(_0247_),
    .A(\stop.syn.daci.din[6] ),
    .B(net123));
 sg13g2_and3_1 _1551_ (.X(_0248_),
    .A(\stop.syn.daci.din[4] ),
    .B(\stop.syn.daci.accumulator[4] ),
    .C(_0242_));
 sg13g2_nor2_1 _1552_ (.A(_0239_),
    .B(_0243_),
    .Y(_0249_));
 sg13g2_a221oi_1 _1553_ (.B2(_0249_),
    .C1(_0248_),
    .B1(_0238_),
    .A1(\stop.syn.daci.din[5] ),
    .Y(_0250_),
    .A2(net121));
 sg13g2_o21ai_1 _1554_ (.B1(net279),
    .Y(_0251_),
    .A1(_0247_),
    .A2(_0250_));
 sg13g2_a21oi_1 _1555_ (.A1(_0247_),
    .A2(_0250_),
    .Y(_0162_),
    .B1(_0251_));
 sg13g2_o21ai_1 _1556_ (.B1(_0246_),
    .Y(_0252_),
    .A1(_0247_),
    .A2(_0250_));
 sg13g2_and2_1 _1557_ (.A(\stop.syn.daci.din[7] ),
    .B(\stop.syn.daci.accumulator[7] ),
    .X(_0253_));
 sg13g2_xor2_1 _1558_ (.B(net132),
    .A(\stop.syn.daci.din[7] ),
    .X(_0254_));
 sg13g2_o21ai_1 _1559_ (.B1(net278),
    .Y(_0255_),
    .A1(_0252_),
    .A2(_0254_));
 sg13g2_a21oi_1 _1560_ (.A1(_0252_),
    .A2(_0254_),
    .Y(_0163_),
    .B1(_0255_));
 sg13g2_a21oi_2 _1561_ (.B1(_0253_),
    .Y(_0256_),
    .A2(_0254_),
    .A1(_0252_));
 sg13g2_a21o_1 _1562_ (.A2(_0254_),
    .A1(_0252_),
    .B1(_0253_),
    .X(_0257_));
 sg13g2_nand2_1 _1563_ (.Y(_0258_),
    .A(\stop.syn.daci.din[8] ),
    .B(net117));
 sg13g2_xnor2_1 _1564_ (.Y(_0259_),
    .A(\stop.syn.daci.din[8] ),
    .B(net117));
 sg13g2_nand2b_1 _1565_ (.Y(_0260_),
    .B(_0257_),
    .A_N(_0259_));
 sg13g2_nand2_1 _1566_ (.Y(_0261_),
    .A(net278),
    .B(_0260_));
 sg13g2_a21oi_1 _1567_ (.A1(_0256_),
    .A2(_0259_),
    .Y(_0164_),
    .B1(_0261_));
 sg13g2_nor2_1 _1568_ (.A(\stop.syn.daci.din[9] ),
    .B(net131),
    .Y(_0262_));
 sg13g2_nand2_1 _1569_ (.Y(_0263_),
    .A(\stop.syn.daci.din[9] ),
    .B(net131));
 sg13g2_nand2b_1 _1570_ (.Y(_0264_),
    .B(_0263_),
    .A_N(_0262_));
 sg13g2_nand3_1 _1571_ (.B(_0260_),
    .C(_0264_),
    .A(_0258_),
    .Y(_0265_));
 sg13g2_a21oi_1 _1572_ (.A1(_0258_),
    .A2(_0260_),
    .Y(_0266_),
    .B1(_0264_));
 sg13g2_nand2_1 _1573_ (.Y(_0267_),
    .A(net278),
    .B(_0265_));
 sg13g2_nor2_1 _1574_ (.A(_0266_),
    .B(_0267_),
    .Y(_0165_));
 sg13g2_nand2_1 _1575_ (.Y(_0268_),
    .A(\stop.syn.daci.din[10] ),
    .B(net113));
 sg13g2_xnor2_1 _1576_ (.Y(_0269_),
    .A(\stop.syn.daci.din[10] ),
    .B(net113));
 sg13g2_o21ai_1 _1577_ (.B1(_0263_),
    .Y(_0270_),
    .A1(_0258_),
    .A2(_0262_));
 sg13g2_nor2_1 _1578_ (.A(_0259_),
    .B(_0264_),
    .Y(_0271_));
 sg13g2_a21oi_1 _1579_ (.A1(_0257_),
    .A2(_0271_),
    .Y(_0272_),
    .B1(_0270_));
 sg13g2_or2_1 _1580_ (.X(_0273_),
    .B(_0272_),
    .A(_0269_));
 sg13g2_nand2_1 _1581_ (.Y(_0274_),
    .A(net278),
    .B(_0273_));
 sg13g2_a21oi_1 _1582_ (.A1(_0269_),
    .A2(_0272_),
    .Y(_0166_),
    .B1(_0274_));
 sg13g2_nor2_1 _1583_ (.A(\stop.syn.daci.din[11] ),
    .B(\stop.syn.daci.accumulator[11] ),
    .Y(_0275_));
 sg13g2_xnor2_1 _1584_ (.Y(_0276_),
    .A(\stop.syn.daci.din[11] ),
    .B(net127));
 sg13g2_nand3_1 _1585_ (.B(_0273_),
    .C(_0276_),
    .A(_0268_),
    .Y(_0277_));
 sg13g2_a21oi_1 _1586_ (.A1(_0268_),
    .A2(_0273_),
    .Y(_0278_),
    .B1(_0276_));
 sg13g2_nand2_1 _1587_ (.Y(_0279_),
    .A(net278),
    .B(_0277_));
 sg13g2_nor2_1 _1588_ (.A(_0278_),
    .B(_0279_),
    .Y(_0167_));
 sg13g2_nor2_1 _1589_ (.A(_0269_),
    .B(_0276_),
    .Y(_0280_));
 sg13g2_nand2_1 _1590_ (.Y(_0281_),
    .A(_0271_),
    .B(_0280_));
 sg13g2_nor2_1 _1591_ (.A(_0256_),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_nor2_1 _1592_ (.A(_0268_),
    .B(_0275_),
    .Y(_0283_));
 sg13g2_a221oi_1 _1593_ (.B2(_0280_),
    .C1(_0283_),
    .B1(_0270_),
    .A1(\stop.syn.daci.din[11] ),
    .Y(_0284_),
    .A2(\stop.syn.daci.accumulator[11] ));
 sg13g2_nor2b_1 _1594_ (.A(_0282_),
    .B_N(_0284_),
    .Y(_0285_));
 sg13g2_o21ai_1 _1595_ (.B1(_0284_),
    .Y(_0286_),
    .A1(_0256_),
    .A2(_0281_));
 sg13g2_nand2_1 _1596_ (.Y(_0287_),
    .A(\stop.syn.daci.din[12] ),
    .B(net116));
 sg13g2_xnor2_1 _1597_ (.Y(_0288_),
    .A(\stop.syn.daci.din[12] ),
    .B(net116));
 sg13g2_nand2b_1 _1598_ (.Y(_0289_),
    .B(_0286_),
    .A_N(_0288_));
 sg13g2_nand2_1 _1599_ (.Y(_0290_),
    .A(net280),
    .B(_0289_));
 sg13g2_a21oi_1 _1600_ (.A1(_0285_),
    .A2(_0288_),
    .Y(_0168_),
    .B1(_0290_));
 sg13g2_nor2_1 _1601_ (.A(\stop.syn.daci.din[13] ),
    .B(\stop.syn.daci.accumulator[13] ),
    .Y(_0291_));
 sg13g2_xnor2_1 _1602_ (.Y(_0292_),
    .A(\stop.syn.daci.din[13] ),
    .B(net119));
 sg13g2_nand3_1 _1603_ (.B(_0289_),
    .C(_0292_),
    .A(_0287_),
    .Y(_0293_));
 sg13g2_a21oi_1 _1604_ (.A1(_0287_),
    .A2(_0289_),
    .Y(_0294_),
    .B1(_0292_));
 sg13g2_nand2_1 _1605_ (.Y(_0295_),
    .A(net280),
    .B(_0293_));
 sg13g2_nor2_1 _1606_ (.A(_0294_),
    .B(_0295_),
    .Y(_0169_));
 sg13g2_nor2_1 _1607_ (.A(_0288_),
    .B(_0292_),
    .Y(_0296_));
 sg13g2_nor2_1 _1608_ (.A(_0287_),
    .B(_0291_),
    .Y(_0297_));
 sg13g2_a221oi_1 _1609_ (.B2(_0296_),
    .C1(_0297_),
    .B1(_0286_),
    .A1(\stop.syn.daci.din[13] ),
    .Y(_0298_),
    .A2(net119));
 sg13g2_nand2_1 _1610_ (.Y(_0299_),
    .A(\stop.syn.daci.din[14] ),
    .B(net115));
 sg13g2_xnor2_1 _1611_ (.Y(_0300_),
    .A(\stop.syn.daci.din[14] ),
    .B(net115));
 sg13g2_o21ai_1 _1612_ (.B1(net280),
    .Y(_0301_),
    .A1(net120),
    .A2(_0300_));
 sg13g2_a21oi_1 _1613_ (.A1(net120),
    .A2(_0300_),
    .Y(_0170_),
    .B1(_0301_));
 sg13g2_xor2_1 _1614_ (.B(net111),
    .A(\stop.syn.daci.din[15] ),
    .X(_0302_));
 sg13g2_o21ai_1 _1615_ (.B1(_0299_),
    .Y(_0303_),
    .A1(_0298_),
    .A2(_0300_));
 sg13g2_o21ai_1 _1616_ (.B1(net278),
    .Y(_0304_),
    .A1(_0302_),
    .A2(_0303_));
 sg13g2_a21oi_1 _1617_ (.A1(_0302_),
    .A2(_0303_),
    .Y(_0171_),
    .B1(_0304_));
 sg13g2_a21oi_1 _1618_ (.A1(\stop.syn.daci.din[15] ),
    .A2(net111),
    .Y(_0305_),
    .B1(_0303_));
 sg13g2_o21ai_1 _1619_ (.B1(net278),
    .Y(_0306_),
    .A1(\stop.syn.daci.din[15] ),
    .A2(net111));
 sg13g2_nor2_1 _1620_ (.A(net112),
    .B(_0306_),
    .Y(_0172_));
 sg13g2_nor2_2 _1621_ (.A(\stop.ctrl.first_bit ),
    .B(net2),
    .Y(_0307_));
 sg13g2_mux2_1 _1622_ (.A0(\stop.adsr_ai[0] ),
    .A1(\stop.adsr_ai[1] ),
    .S(net342),
    .X(_0173_));
 sg13g2_nor2_1 _1623_ (.A(\stop.adsr_ai[1] ),
    .B(net343),
    .Y(_0308_));
 sg13g2_a21oi_1 _1624_ (.A1(_0321_),
    .A2(net343),
    .Y(_0174_),
    .B1(_0308_));
 sg13g2_nor2_1 _1625_ (.A(\stop.adsr_ai[2] ),
    .B(net341),
    .Y(_0309_));
 sg13g2_a21oi_1 _1626_ (.A1(_0322_),
    .A2(net341),
    .Y(_0175_),
    .B1(_0309_));
 sg13g2_nor2_1 _1627_ (.A(\stop.adsr_ai[3] ),
    .B(net341),
    .Y(_0310_));
 sg13g2_a21oi_1 _1628_ (.A1(_0323_),
    .A2(net341),
    .Y(_0176_),
    .B1(_0310_));
 sg13g2_nor2_1 _1629_ (.A(\stop.adsr_ai[4] ),
    .B(net341),
    .Y(_0311_));
 sg13g2_a21oi_1 _1630_ (.A1(_0324_),
    .A2(net342),
    .Y(_0177_),
    .B1(_0311_));
 sg13g2_nor2_1 _1631_ (.A(\stop.adsr_ai[5] ),
    .B(net339),
    .Y(_0312_));
 sg13g2_a21oi_1 _1632_ (.A1(_0325_),
    .A2(net339),
    .Y(_0178_),
    .B1(_0312_));
 sg13g2_nor2_1 _1633_ (.A(\stop.adsr_ai[6] ),
    .B(net339),
    .Y(_0313_));
 sg13g2_a21oi_1 _1634_ (.A1(_0326_),
    .A2(net339),
    .Y(_0179_),
    .B1(_0313_));
 sg13g2_nand2_1 _1635_ (.Y(_0314_),
    .A(\stop.adsr_di[0] ),
    .B(net340));
 sg13g2_o21ai_1 _1636_ (.B1(_0314_),
    .Y(_0180_),
    .A1(_0326_),
    .A2(net339));
 sg13g2_mux2_1 _1637_ (.A0(\stop.adsr_di[0] ),
    .A1(\stop.adsr_di[1] ),
    .S(net342),
    .X(_0181_));
 sg13g2_mux2_1 _1638_ (.A0(\stop.adsr_di[1] ),
    .A1(\stop.adsr_di[2] ),
    .S(net342),
    .X(_0182_));
 sg13g2_mux2_1 _1639_ (.A0(\stop.adsr_di[2] ),
    .A1(\stop.adsr_di[3] ),
    .S(net342),
    .X(_0183_));
 sg13g2_mux2_1 _1640_ (.A0(\stop.adsr_di[3] ),
    .A1(\stop.adsr_di[4] ),
    .S(net342),
    .X(_0184_));
 sg13g2_mux2_1 _1641_ (.A0(\stop.adsr_di[4] ),
    .A1(\stop.adsr_di[5] ),
    .S(net339),
    .X(_0185_));
 sg13g2_mux2_1 _1642_ (.A0(\stop.adsr_di[5] ),
    .A1(\stop.adsr_di[6] ),
    .S(net339),
    .X(_0186_));
 sg13g2_mux2_1 _1643_ (.A0(\stop.adsr_di[6] ),
    .A1(\stop.adsr_di[7] ),
    .S(net340),
    .X(_0187_));
 sg13g2_mux2_1 _1644_ (.A0(\stop.adsr_di[7] ),
    .A1(\stop.adsr_s[0] ),
    .S(net340),
    .X(_0188_));
 sg13g2_mux2_1 _1645_ (.A0(\stop.adsr_s[0] ),
    .A1(\stop.adsr_s[1] ),
    .S(net345),
    .X(_0189_));
 sg13g2_mux2_1 _1646_ (.A0(\stop.adsr_s[1] ),
    .A1(\stop.adsr_s[2] ),
    .S(net344),
    .X(_0190_));
 sg13g2_mux2_1 _1647_ (.A0(\stop.adsr_s[2] ),
    .A1(\stop.adsr_s[3] ),
    .S(net344),
    .X(_0191_));
 sg13g2_mux2_1 _1648_ (.A0(\stop.adsr_s[3] ),
    .A1(\stop.adsr_s[4] ),
    .S(net344),
    .X(_0192_));
 sg13g2_mux2_1 _1649_ (.A0(\stop.adsr_s[4] ),
    .A1(\stop.adsr_s[5] ),
    .S(net344),
    .X(_0193_));
 sg13g2_mux2_1 _1650_ (.A0(\stop.adsr_s[5] ),
    .A1(\stop.adsr_s[6] ),
    .S(net344),
    .X(_0194_));
 sg13g2_mux2_1 _1651_ (.A0(\stop.adsr_s[6] ),
    .A1(\stop.adsr_s[7] ),
    .S(net344),
    .X(_0195_));
 sg13g2_mux2_1 _1652_ (.A0(\stop.adsr_s[7] ),
    .A1(\stop.adsr_ri[0] ),
    .S(net341),
    .X(_0196_));
 sg13g2_mux2_1 _1653_ (.A0(\stop.adsr_ri[0] ),
    .A1(\stop.adsr_ri[1] ),
    .S(net343),
    .X(_0197_));
 sg13g2_mux2_1 _1654_ (.A0(\stop.adsr_ri[1] ),
    .A1(\stop.adsr_ri[2] ),
    .S(net341),
    .X(_0198_));
 sg13g2_mux2_1 _1655_ (.A0(\stop.adsr_ri[2] ),
    .A1(\stop.adsr_ri[3] ),
    .S(net341),
    .X(_0199_));
 sg13g2_mux2_1 _1656_ (.A0(\stop.adsr_ri[3] ),
    .A1(\stop.adsr_ri[4] ),
    .S(net342),
    .X(_0200_));
 sg13g2_mux2_1 _1657_ (.A0(\stop.adsr_ri[4] ),
    .A1(\stop.adsr_ri[5] ),
    .S(net342),
    .X(_0201_));
 sg13g2_mux2_1 _1658_ (.A0(\stop.adsr_ri[5] ),
    .A1(\stop.adsr_ri[6] ),
    .S(net339),
    .X(_0202_));
 sg13g2_mux2_1 _1659_ (.A0(\stop.adsr_ri[6] ),
    .A1(\stop.adsr_ri[7] ),
    .S(net340),
    .X(_0203_));
 sg13g2_mux2_1 _1660_ (.A0(\stop.adsr_ri[7] ),
    .A1(\stop.ctrl.cfg[32] ),
    .S(net336),
    .X(_0204_));
 sg13g2_mux2_1 _1661_ (.A0(\stop.ctrl.cfg[32] ),
    .A1(\stop.ctrl.cfg[33] ),
    .S(net337),
    .X(_0205_));
 sg13g2_mux2_1 _1662_ (.A0(\stop.ctrl.cfg[33] ),
    .A1(\stop.ctrl.cfg[34] ),
    .S(net346),
    .X(_0206_));
 sg13g2_mux2_1 _1663_ (.A0(\stop.ctrl.cfg[34] ),
    .A1(\stop.ctrl.cfg[35] ),
    .S(net338),
    .X(_0207_));
 sg13g2_mux2_1 _1664_ (.A0(\stop.ctrl.cfg[35] ),
    .A1(\stop.ctrl.cfg[36] ),
    .S(net338),
    .X(_0208_));
 sg13g2_mux2_1 _1665_ (.A0(\stop.ctrl.cfg[36] ),
    .A1(\stop.ctrl.cfg[37] ),
    .S(net338),
    .X(_0209_));
 sg13g2_mux2_1 _1666_ (.A0(\stop.ctrl.cfg[37] ),
    .A1(\stop.ctrl.cfg[38] ),
    .S(net338),
    .X(_0210_));
 sg13g2_mux2_1 _1667_ (.A0(\stop.ctrl.cfg[38] ),
    .A1(\stop.ctrl.cfg[39] ),
    .S(net338),
    .X(_0211_));
 sg13g2_mux2_1 _1668_ (.A0(\stop.ctrl.cfg[39] ),
    .A1(\stop.ctrl.cfg[40] ),
    .S(net338),
    .X(_0212_));
 sg13g2_mux2_1 _1669_ (.A0(\stop.ctrl.cfg[40] ),
    .A1(\stop.ctrl.cfg[41] ),
    .S(net338),
    .X(_0213_));
 sg13g2_mux2_1 _1670_ (.A0(\stop.ctrl.cfg[41] ),
    .A1(\stop.ctrl.cfg[42] ),
    .S(net338),
    .X(_0214_));
 sg13g2_mux2_1 _1671_ (.A0(\stop.ctrl.cfg[42] ),
    .A1(\stop.ctrl.cfg[43] ),
    .S(net335),
    .X(_0215_));
 sg13g2_mux2_1 _1672_ (.A0(\stop.ctrl.cfg[43] ),
    .A1(\stop.ctrl.cfg[44] ),
    .S(net335),
    .X(_0216_));
 sg13g2_mux2_1 _1673_ (.A0(\stop.ctrl.cfg[44] ),
    .A1(\stop.ctrl.cfg[45] ),
    .S(net337),
    .X(_0217_));
 sg13g2_mux2_1 _1674_ (.A0(\stop.ctrl.cfg[45] ),
    .A1(\stop.ctrl.cfg[46] ),
    .S(net337),
    .X(_0218_));
 sg13g2_mux2_1 _1675_ (.A0(\stop.ctrl.cfg[46] ),
    .A1(\stop.ctrl.cfg[47] ),
    .S(net335),
    .X(_0219_));
 sg13g2_mux2_1 _1676_ (.A0(\stop.ctrl.cfg[47] ),
    .A1(\stop.ctrl.cfg[48] ),
    .S(net335),
    .X(_0220_));
 sg13g2_mux2_1 _1677_ (.A0(\stop.ctrl.cfg[48] ),
    .A1(\stop.ctrl.cfg[49] ),
    .S(net335),
    .X(_0221_));
 sg13g2_mux2_1 _1678_ (.A0(\stop.ctrl.cfg[49] ),
    .A1(\stop.ctrl.cfg[50] ),
    .S(net335),
    .X(_0222_));
 sg13g2_mux2_1 _1679_ (.A0(\stop.ctrl.cfg[50] ),
    .A1(\stop.ctrl.cfg[51] ),
    .S(net335),
    .X(_0223_));
 sg13g2_mux2_1 _1680_ (.A0(\stop.ctrl.cfg[51] ),
    .A1(\stop.ctrl.cfg[52] ),
    .S(net335),
    .X(_0224_));
 sg13g2_mux2_1 _1681_ (.A0(\stop.ctrl.cfg[52] ),
    .A1(\stop.ctrl.cfg[53] ),
    .S(net336),
    .X(_0225_));
 sg13g2_mux2_1 _1682_ (.A0(\stop.ctrl.cfg[53] ),
    .A1(\stop.ctrl.cfg[54] ),
    .S(net336),
    .X(_0226_));
 sg13g2_mux2_1 _1683_ (.A0(\stop.ctrl.cfg[54] ),
    .A1(\stop.ctrl.cfg[55] ),
    .S(net336),
    .X(_0227_));
 sg13g2_mux2_1 _1684_ (.A0(\stop.ctrl.cfg[55] ),
    .A1(\stop.ctrl.cfg[56] ),
    .S(net336),
    .X(_0228_));
 sg13g2_mux2_1 _1685_ (.A0(\stop.ctrl.cfg[56] ),
    .A1(\stop.ctrl.cfg[57] ),
    .S(net336),
    .X(_0229_));
 sg13g2_mux2_1 _1686_ (.A0(\stop.ctrl.cfg[57] ),
    .A1(\stop.ctrl.cfg[58] ),
    .S(net336),
    .X(_0230_));
 sg13g2_mux2_1 _1687_ (.A0(\stop.ctrl.cfg[58] ),
    .A1(\stop.ctrl.cfg[59] ),
    .S(net336),
    .X(_0231_));
 sg13g2_mux2_1 _1688_ (.A0(\stop.ctrl.cfg[59] ),
    .A1(net3),
    .S(net345),
    .X(_0232_));
 sg13g2_inv_1 _1689_ (.Y(_0130_),
    .A(net295));
 sg13g2_inv_1 _1690_ (.Y(_0129_),
    .A(net298));
 sg13g2_inv_1 _1691_ (.Y(_0128_),
    .A(net297));
 sg13g2_inv_1 _1692_ (.Y(_0127_),
    .A(net297));
 sg13g2_inv_1 _1693_ (.Y(_0126_),
    .A(net296));
 sg13g2_inv_1 _1694_ (.Y(_0125_),
    .A(net296));
 sg13g2_inv_1 _1695_ (.Y(_0124_),
    .A(net296));
 sg13g2_inv_1 _1696_ (.Y(_0123_),
    .A(net296));
 sg13g2_inv_1 _1697_ (.Y(_0122_),
    .A(net296));
 sg13g2_inv_1 _1698_ (.Y(_0121_),
    .A(net296));
 sg13g2_inv_1 _1699_ (.Y(_0120_),
    .A(net297));
 sg13g2_inv_1 _1700_ (.Y(_0119_),
    .A(net297));
 sg13g2_inv_1 _1701_ (.Y(_0118_),
    .A(net297));
 sg13g2_inv_1 _1702_ (.Y(_0117_),
    .A(net297));
 sg13g2_inv_1 _1703_ (.Y(_0116_),
    .A(net297));
 sg13g2_inv_1 _1704_ (.Y(_0115_),
    .A(net295));
 sg13g2_inv_1 _1705_ (.Y(_0114_),
    .A(net295));
 sg13g2_inv_1 _1706_ (.Y(_0113_),
    .A(net296));
 sg13g2_inv_1 _1707_ (.Y(_0112_),
    .A(net292));
 sg13g2_inv_1 _1708_ (.Y(_0111_),
    .A(net292));
 sg13g2_inv_1 _1709_ (.Y(_0110_),
    .A(net292));
 sg13g2_inv_1 _1710_ (.Y(_0109_),
    .A(net292));
 sg13g2_inv_1 _1711_ (.Y(_0108_),
    .A(net293));
 sg13g2_inv_1 _1712_ (.Y(_0107_),
    .A(net293));
 sg13g2_inv_1 _1713_ (.Y(_0106_),
    .A(net293));
 sg13g2_inv_1 _1714_ (.Y(_0105_),
    .A(net291));
 sg13g2_inv_1 _1715_ (.Y(_0104_),
    .A(net290));
 sg13g2_inv_1 _1716_ (.Y(_0103_),
    .A(net293));
 sg13g2_inv_1 _1717_ (.Y(_0102_),
    .A(net292));
 sg13g2_inv_1 _1718_ (.Y(_0101_),
    .A(net292));
 sg13g2_inv_1 _1719_ (.Y(_0100_),
    .A(net296));
 sg13g2_inv_1 _1720_ (.Y(_0099_),
    .A(net289));
 sg13g2_inv_1 _1721_ (.Y(_0098_),
    .A(net289));
 sg13g2_inv_1 _1722_ (.Y(_0097_),
    .A(net288));
 sg13g2_inv_1 _1723_ (.Y(_0096_),
    .A(net291));
 sg13g2_inv_1 _1724_ (.Y(_0095_),
    .A(net291));
 sg13g2_inv_1 _1725_ (.Y(_0094_),
    .A(net291));
 sg13g2_inv_1 _1726_ (.Y(_0093_),
    .A(net290));
 sg13g2_inv_1 _1727_ (.Y(_0092_),
    .A(net290));
 sg13g2_inv_1 _1728_ (.Y(_0091_),
    .A(net290));
 sg13g2_inv_1 _1729_ (.Y(_0090_),
    .A(net290));
 sg13g2_inv_1 _1730_ (.Y(_0089_),
    .A(net290));
 sg13g2_inv_1 _1731_ (.Y(_0088_),
    .A(net290));
 sg13g2_inv_1 _1732_ (.Y(_0087_),
    .A(net290));
 sg13g2_inv_1 _1733_ (.Y(_0086_),
    .A(net291));
 sg13g2_inv_1 _1734_ (.Y(_0085_),
    .A(net292));
 sg13g2_inv_1 _1735_ (.Y(_0084_),
    .A(net292));
 sg13g2_inv_1 _1736_ (.Y(_0083_),
    .A(net2));
 sg13g2_dfrbp_1 _1737_ (.CLK(net321),
    .RESET_B(net23),
    .D(_0012_),
    .Q_N(_0879_),
    .Q(\stop.syn.filt.m2.b_bit ));
 sg13g2_dfrbp_1 _1738_ (.CLK(net321),
    .RESET_B(net28),
    .D(_0013_),
    .Q_N(_0878_),
    .Q(\stop.syn.filt.m2.b_latched[1] ));
 sg13g2_dfrbp_1 _1739_ (.CLK(net321),
    .RESET_B(net22),
    .D(_0014_),
    .Q_N(_0877_),
    .Q(\stop.syn.filt.m2.b_latched[2] ));
 sg13g2_dfrbp_1 _1740_ (.CLK(net321),
    .RESET_B(net21),
    .D(_0015_),
    .Q_N(_0876_),
    .Q(\stop.syn.filt.m2.b_latched[3] ));
 sg13g2_dfrbp_1 _1741_ (.CLK(net321),
    .RESET_B(net20),
    .D(_0016_),
    .Q_N(_0875_),
    .Q(\stop.syn.filt.m2.b_latched[4] ));
 sg13g2_dfrbp_1 _1742_ (.CLK(net327),
    .RESET_B(net19),
    .D(_0017_),
    .Q_N(_0874_),
    .Q(\stop.syn.filt.m2.b_latched[5] ));
 sg13g2_dfrbp_1 _1743_ (.CLK(net321),
    .RESET_B(net24),
    .D(_0018_),
    .Q_N(_0880_),
    .Q(\stop.syn.filt.m2.b_latched[6] ));
 sg13g2_dfrbp_1 _1744_ (.CLK(net285),
    .RESET_B(net25),
    .D(_0000_),
    .Q_N(_0881_),
    .Q(\stop.syn.adsri.state[0] ));
 sg13g2_dfrbp_1 _1745_ (.CLK(net285),
    .RESET_B(net26),
    .D(_0001_),
    .Q_N(_0882_),
    .Q(\stop.syn.adsri.state[1] ));
 sg13g2_dfrbp_1 _1746_ (.CLK(net285),
    .RESET_B(net27),
    .D(_0002_),
    .Q_N(_0883_),
    .Q(\stop.syn.adsri.state[2] ));
 sg13g2_dfrbp_1 _1747_ (.CLK(net285),
    .RESET_B(net45),
    .D(_0003_),
    .Q_N(_0884_),
    .Q(\stop.syn.adsri.state[3] ));
 sg13g2_dfrbp_1 _1748_ (.CLK(net285),
    .RESET_B(net18),
    .D(_0004_),
    .Q_N(_0873_),
    .Q(\stop.syn.adsri.state[4] ));
 sg13g2_dfrbp_1 _1749_ (.CLK(net327),
    .RESET_B(net17),
    .D(_0132_),
    .Q_N(_0872_),
    .Q(\stop.syn.smul8.b_latched[7] ));
 sg13g2_dfrbp_1 _1750_ (.CLK(net322),
    .RESET_B(net103),
    .D(_0005_),
    .Q_N(_0871_),
    .Q(\stop.syn.filt.m1.b_bit ));
 sg13g2_dfrbp_1 _1751_ (.CLK(net319),
    .RESET_B(net102),
    .D(_0006_),
    .Q_N(_0870_),
    .Q(\stop.syn.filt.m1.b_latched[1] ));
 sg13g2_dfrbp_1 _1752_ (.CLK(net319),
    .RESET_B(net101),
    .D(_0007_),
    .Q_N(_0869_),
    .Q(\stop.syn.filt.m1.b_latched[2] ));
 sg13g2_dfrbp_1 _1753_ (.CLK(net319),
    .RESET_B(net100),
    .D(_0008_),
    .Q_N(_0868_),
    .Q(\stop.syn.filt.m1.b_latched[3] ));
 sg13g2_dfrbp_1 _1754_ (.CLK(net319),
    .RESET_B(net99),
    .D(_0009_),
    .Q_N(_0867_),
    .Q(\stop.syn.filt.m1.b_latched[4] ));
 sg13g2_dfrbp_1 _1755_ (.CLK(net319),
    .RESET_B(net98),
    .D(_0010_),
    .Q_N(_0866_),
    .Q(\stop.syn.filt.m1.b_latched[5] ));
 sg13g2_dfrbp_1 _1756_ (.CLK(net319),
    .RESET_B(net97),
    .D(_0011_),
    .Q_N(_0865_),
    .Q(\stop.syn.filt.m1.b_latched[6] ));
 sg13g2_dfrbp_1 _1757_ (.CLK(net319),
    .RESET_B(net96),
    .D(_0019_),
    .Q_N(_0864_),
    .Q(\stop.syn.smul8.b_bit ));
 sg13g2_dfrbp_1 _1758_ (.CLK(net327),
    .RESET_B(net95),
    .D(_0020_),
    .Q_N(_0863_),
    .Q(\stop.syn.smul8.b_latched[1] ));
 sg13g2_dfrbp_1 _1759_ (.CLK(net330),
    .RESET_B(net94),
    .D(_0021_),
    .Q_N(_0862_),
    .Q(\stop.syn.smul8.b_latched[2] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(net327),
    .RESET_B(net93),
    .D(_0022_),
    .Q_N(_0861_),
    .Q(\stop.syn.smul8.b_latched[3] ));
 sg13g2_dfrbp_1 _1761_ (.CLK(net327),
    .RESET_B(net92),
    .D(_0023_),
    .Q_N(_0860_),
    .Q(\stop.syn.smul8.b_latched[4] ));
 sg13g2_dfrbp_1 _1762_ (.CLK(net327),
    .RESET_B(net91),
    .D(_0024_),
    .Q_N(_0859_),
    .Q(\stop.syn.smul8.b_latched[5] ));
 sg13g2_dfrbp_1 _1763_ (.CLK(net327),
    .RESET_B(net90),
    .D(_0025_),
    .Q_N(_0858_),
    .Q(\stop.syn.smul8.b_latched[6] ));
 sg13g2_dfrbp_1 _1764_ (.CLK(net359),
    .RESET_B(_0081_),
    .D(_0080_),
    .Q_N(\stop.ctrl.first_bit_reg ),
    .Q(_0078_));
 sg13g2_dfrbp_1 _1765_ (.CLK(net359),
    .RESET_B(net370),
    .D(_0133_),
    .Q_N(_0857_),
    .Q(\stop.ctrl.trig ));
 sg13g2_dfrbp_1 _1766_ (.CLK(net359),
    .RESET_B(_0083_),
    .D(net106),
    .Q_N(\stop.ctrl.first_bit ),
    .Q(_0079_));
 sg13g2_dfrbp_1 _1767_ (.CLK(net299),
    .RESET_B(net88),
    .D(_0134_),
    .Q_N(_0856_),
    .Q(\stop.syn.osci.counter[0] ));
 sg13g2_dfrbp_1 _1768_ (.CLK(net299),
    .RESET_B(net87),
    .D(_0135_),
    .Q_N(_0855_),
    .Q(\stop.syn.osci.counter[1] ));
 sg13g2_dfrbp_1 _1769_ (.CLK(net299),
    .RESET_B(net86),
    .D(_0136_),
    .Q_N(_0854_),
    .Q(\stop.syn.osci.counter[2] ));
 sg13g2_dfrbp_1 _1770_ (.CLK(net299),
    .RESET_B(net85),
    .D(_0137_),
    .Q_N(_0853_),
    .Q(\stop.syn.osci.counter[3] ));
 sg13g2_dfrbp_1 _1771_ (.CLK(net301),
    .RESET_B(net84),
    .D(_0138_),
    .Q_N(_0852_),
    .Q(\stop.dbg_osc0 ));
 sg13g2_dfrbp_1 _1772_ (.CLK(net301),
    .RESET_B(net83),
    .D(_0139_),
    .Q_N(_0851_),
    .Q(\stop.syn.osc_data[1] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(net301),
    .RESET_B(net82),
    .D(_0140_),
    .Q_N(_0850_),
    .Q(\stop.syn.osc_data[2] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(net300),
    .RESET_B(net81),
    .D(_0141_),
    .Q_N(_0849_),
    .Q(\stop.syn.osc_data[3] ));
 sg13g2_dfrbp_1 _1775_ (.CLK(net300),
    .RESET_B(net80),
    .D(_0142_),
    .Q_N(_0848_),
    .Q(\stop.syn.osc_data[4] ));
 sg13g2_dfrbp_1 _1776_ (.CLK(net300),
    .RESET_B(net79),
    .D(_0143_),
    .Q_N(_0847_),
    .Q(\stop.syn.osc_data[5] ));
 sg13g2_dfrbp_1 _1777_ (.CLK(net300),
    .RESET_B(net78),
    .D(_0144_),
    .Q_N(_0846_),
    .Q(\stop.syn.osc_data[6] ));
 sg13g2_dfrbp_1 _1778_ (.CLK(net300),
    .RESET_B(net46),
    .D(_0145_),
    .Q_N(_0885_),
    .Q(\stop.syn.osc_data[7] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(net303),
    .RESET_B(net47),
    .D(\stop.dbg_adsr0 ),
    .Q_N(_0886_),
    .Q(\stop.dbg_adsr_reg0 ));
 sg13g2_dfrbp_1 _1780_ (.CLK(net302),
    .RESET_B(net48),
    .D(\stop.syn.adsr_data[1] ),
    .Q_N(_0887_),
    .Q(\stop.syn.adsr_data_reg[1] ));
 sg13g2_dfrbp_1 _1781_ (.CLK(net302),
    .RESET_B(net49),
    .D(\stop.syn.adsr_data[2] ),
    .Q_N(_0888_),
    .Q(\stop.syn.adsr_data_reg[2] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(net301),
    .RESET_B(net50),
    .D(\stop.syn.adsr_data[3] ),
    .Q_N(_0889_),
    .Q(\stop.syn.adsr_data_reg[3] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(net301),
    .RESET_B(net51),
    .D(\stop.syn.adsr_data[4] ),
    .Q_N(_0890_),
    .Q(\stop.syn.adsr_data_reg[4] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(net301),
    .RESET_B(net52),
    .D(\stop.syn.adsr_data[5] ),
    .Q_N(_0891_),
    .Q(\stop.syn.adsr_data_reg[5] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(net302),
    .RESET_B(net53),
    .D(\stop.syn.adsr_data[6] ),
    .Q_N(_0892_),
    .Q(\stop.syn.adsr_data_reg[6] ));
 sg13g2_dfrbp_1 _1786_ (.CLK(net301),
    .RESET_B(net54),
    .D(\stop.syn.adsr_data[7] ),
    .Q_N(_0893_),
    .Q(\stop.syn.adsr_data_reg[7] ));
 sg13g2_dfrbp_1 _1787_ (.CLK(net302),
    .RESET_B(net55),
    .D(\stop.syn.adsr_data[8] ),
    .Q_N(_0894_),
    .Q(\stop.syn.adsr_data_reg[8] ));
 sg13g2_dfrbp_1 _1788_ (.CLK(net301),
    .RESET_B(net56),
    .D(\stop.syn.adsr_data[9] ),
    .Q_N(_0895_),
    .Q(\stop.syn.adsr_data_reg[9] ));
 sg13g2_dfrbp_1 _1789_ (.CLK(net302),
    .RESET_B(net57),
    .D(\stop.syn.adsr_data[10] ),
    .Q_N(_0896_),
    .Q(\stop.syn.adsr_data_reg[10] ));
 sg13g2_dfrbp_1 _1790_ (.CLK(net300),
    .RESET_B(net58),
    .D(\stop.syn.adsr_data[11] ),
    .Q_N(_0897_),
    .Q(\stop.syn.adsr_data_reg[11] ));
 sg13g2_dfrbp_1 _1791_ (.CLK(net299),
    .RESET_B(net59),
    .D(\stop.syn.adsr_data[12] ),
    .Q_N(_0898_),
    .Q(\stop.syn.adsr_data_reg[12] ));
 sg13g2_dfrbp_1 _1792_ (.CLK(net306),
    .RESET_B(net60),
    .D(\stop.syn.adsr_data[13] ),
    .Q_N(_0899_),
    .Q(\stop.syn.adsr_data_reg[13] ));
 sg13g2_dfrbp_1 _1793_ (.CLK(net299),
    .RESET_B(net61),
    .D(\stop.syn.adsr_data[14] ),
    .Q_N(_0900_),
    .Q(\stop.syn.adsr_data_reg[14] ));
 sg13g2_dfrbp_1 _1794_ (.CLK(net299),
    .RESET_B(net62),
    .D(\stop.syn.adsr_data[15] ),
    .Q_N(_0901_),
    .Q(\stop.syn.adsr_data_reg[15] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net63),
    .D(net333),
    .Q_N(_0902_),
    .Q(\stop.syn.rstn_fst_reg1 ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net64),
    .D(net108),
    .Q_N(_0903_),
    .Q(\stop.syn.rstn_fst_reg2 ));
 sg13g2_dfrbp_1 _1797_ (.CLK(net287),
    .RESET_B(net65),
    .D(\stop.dbg_trig ),
    .Q_N(_0904_),
    .Q(\stop.syn.trig_reg1 ));
 sg13g2_dfrbp_1 _1798_ (.CLK(net287),
    .RESET_B(net66),
    .D(\stop.syn.trig_reg1 ),
    .Q_N(_0905_),
    .Q(\stop.syn.adsri.trig ));
 sg13g2_dfrbp_1 _1799_ (.CLK(net286),
    .RESET_B(net67),
    .D(net333),
    .Q_N(_0906_),
    .Q(\stop.syn.rstn_reg1 ));
 sg13g2_dfrbp_1 _1800_ (.CLK(net286),
    .RESET_B(net68),
    .D(\stop.syn.rstn_reg1 ),
    .Q_N(_0045_),
    .Q(\stop.syn.adsri.rstn ));
 sg13g2_dfrbp_1 _1801_ (.CLK(\stop.syn.clki.gen[14].inst.q ),
    .RESET_B(net348),
    .D(_0033_),
    .Q_N(_0033_),
    .Q(\stop.dbg_clk_adsr ));
 sg13g2_dfrbp_1 _1802_ (.CLK(\stop.syn.clki.gen[13].inst.q ),
    .RESET_B(net348),
    .D(_0032_),
    .Q_N(_0032_),
    .Q(\stop.syn.clki.gen[14].inst.q ));
 sg13g2_dfrbp_1 _1803_ (.CLK(\stop.syn.clki.gen[12].inst.q ),
    .RESET_B(net348),
    .D(_0031_),
    .Q_N(_0031_),
    .Q(\stop.syn.clki.gen[13].inst.q ));
 sg13g2_dfrbp_1 _1804_ (.CLK(\stop.syn.clki.gen[11].inst.q ),
    .RESET_B(net348),
    .D(_0030_),
    .Q_N(_0030_),
    .Q(\stop.syn.clki.gen[12].inst.q ));
 sg13g2_dfrbp_1 _1805_ (.CLK(\stop.syn.clki.gen[10].inst.q ),
    .RESET_B(net348),
    .D(_0029_),
    .Q_N(_0029_),
    .Q(\stop.syn.clki.gen[11].inst.q ));
 sg13g2_dfrbp_1 _1806_ (.CLK(\stop.syn.clki.gen[10].inst.clk ),
    .RESET_B(net348),
    .D(_0028_),
    .Q_N(_0028_),
    .Q(\stop.syn.clki.gen[10].inst.q ));
 sg13g2_dfrbp_1 _1807_ (.CLK(net299),
    .RESET_B(net348),
    .D(_0041_),
    .Q_N(_0041_),
    .Q(\stop.syn.clki.gen[10].inst.clk ));
 sg13g2_dfrbp_1 _1808_ (.CLK(\stop.syn.clk_sample_x2 ),
    .RESET_B(net347),
    .D(_0040_),
    .Q_N(_0040_),
    .Q(\stop.dbg_clk_sample ));
 sg13g2_dfrbp_1 _1809_ (.CLK(\stop.syn.clki.gen[6].inst.q ),
    .RESET_B(net347),
    .D(_0026_),
    .Q_N(_0026_),
    .Q(\stop.syn.clk_sample_x2 ));
 sg13g2_dfrbp_1 _1810_ (.CLK(\stop.syn.clki.gen[5].inst.q ),
    .RESET_B(net347),
    .D(_0039_),
    .Q_N(_0039_),
    .Q(\stop.syn.clki.gen[6].inst.q ));
 sg13g2_dfrbp_1 _1811_ (.CLK(\stop.syn.clk_mult ),
    .RESET_B(net347),
    .D(_0038_),
    .Q_N(_0038_),
    .Q(\stop.syn.clki.gen[5].inst.q ));
 sg13g2_dfrbp_1 _1812_ (.CLK(\stop.syn.clki.gen[3].inst.q ),
    .RESET_B(net347),
    .D(net320),
    .Q_N(_0037_),
    .Q(\stop.syn.clk_mult ));
 sg13g2_dfrbp_1 _1813_ (.CLK(\stop.syn.clki.gen[2].inst.q ),
    .RESET_B(net347),
    .D(_0036_),
    .Q_N(_0036_),
    .Q(\stop.syn.clki.gen[3].inst.q ));
 sg13g2_dfrbp_1 _1814_ (.CLK(\stop.syn.clki.gen[1].inst.q ),
    .RESET_B(net347),
    .D(_0035_),
    .Q_N(_0035_),
    .Q(\stop.syn.clki.gen[2].inst.q ));
 sg13g2_dfrbp_1 _1815_ (.CLK(\stop.syn.clki.gen[0].inst.q ),
    .RESET_B(net347),
    .D(_0034_),
    .Q_N(_0034_),
    .Q(\stop.syn.clki.gen[1].inst.q ));
 sg13g2_dfrbp_1 _1816_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net348),
    .D(net107),
    .Q_N(_0027_),
    .Q(\stop.syn.clki.gen[0].inst.q ));
 sg13g2_dfrbp_1 _1817_ (.CLK(net285),
    .RESET_B(net77),
    .D(_0146_),
    .Q_N(_0845_),
    .Q(\stop.dbg_env0 ));
 sg13g2_dfrbp_1 _1818_ (.CLK(net286),
    .RESET_B(net76),
    .D(_0147_),
    .Q_N(_0844_),
    .Q(\stop.syn.adsri.envelope[1] ));
 sg13g2_dfrbp_1 _1819_ (.CLK(net286),
    .RESET_B(net75),
    .D(_0148_),
    .Q_N(_0843_),
    .Q(\stop.syn.adsri.envelope[2] ));
 sg13g2_dfrbp_1 _1820_ (.CLK(net286),
    .RESET_B(net74),
    .D(_0149_),
    .Q_N(_0842_),
    .Q(\stop.syn.adsri.envelope[3] ));
 sg13g2_dfrbp_1 _1821_ (.CLK(net286),
    .RESET_B(net73),
    .D(_0150_),
    .Q_N(_0841_),
    .Q(\stop.syn.adsri.envelope[4] ));
 sg13g2_dfrbp_1 _1822_ (.CLK(net286),
    .RESET_B(net72),
    .D(_0151_),
    .Q_N(_0840_),
    .Q(\stop.syn.adsri.envelope[5] ));
 sg13g2_dfrbp_1 _1823_ (.CLK(net285),
    .RESET_B(net71),
    .D(_0152_),
    .Q_N(_0839_),
    .Q(\stop.syn.adsri.envelope[6] ));
 sg13g2_dfrbp_1 _1824_ (.CLK(net285),
    .RESET_B(net70),
    .D(_0153_),
    .Q_N(_0838_),
    .Q(\stop.syn.adsri.envelope[7] ));
 sg13g2_dfrbp_1 _1825_ (.CLK(net321),
    .RESET_B(net69),
    .D(_0154_),
    .Q_N(_0837_),
    .Q(\stop.syn.filt.m2.b_latched[7] ));
 sg13g2_dfrbp_1 _1826_ (.CLK(net325),
    .RESET_B(_0084_),
    .D(\stop.syn.adsr_data[1] ),
    .Q_N(_0836_),
    .Q(\stop.dbg_adsr0 ));
 sg13g2_dfrbp_1 _1827_ (.CLK(net325),
    .RESET_B(_0085_),
    .D(\stop.syn.adsr_data[2] ),
    .Q_N(_0835_),
    .Q(\stop.syn.adsr_data[1] ));
 sg13g2_dfrbp_1 _1828_ (.CLK(net324),
    .RESET_B(_0086_),
    .D(\stop.syn.adsr_data[3] ),
    .Q_N(_0834_),
    .Q(\stop.syn.adsr_data[2] ));
 sg13g2_dfrbp_1 _1829_ (.CLK(net323),
    .RESET_B(_0087_),
    .D(\stop.syn.adsr_data[4] ),
    .Q_N(_0833_),
    .Q(\stop.syn.adsr_data[3] ));
 sg13g2_dfrbp_1 _1830_ (.CLK(net323),
    .RESET_B(_0088_),
    .D(\stop.syn.adsr_data[5] ),
    .Q_N(_0832_),
    .Q(\stop.syn.adsr_data[4] ));
 sg13g2_dfrbp_1 _1831_ (.CLK(net323),
    .RESET_B(_0089_),
    .D(\stop.syn.adsr_data[6] ),
    .Q_N(_0831_),
    .Q(\stop.syn.adsr_data[5] ));
 sg13g2_dfrbp_1 _1832_ (.CLK(net323),
    .RESET_B(_0090_),
    .D(\stop.syn.adsr_data[7] ),
    .Q_N(_0830_),
    .Q(\stop.syn.adsr_data[6] ));
 sg13g2_dfrbp_1 _1833_ (.CLK(net323),
    .RESET_B(_0091_),
    .D(_0070_),
    .Q_N(_0829_),
    .Q(\stop.syn.adsr_data[7] ));
 sg13g2_dfrbp_1 _1834_ (.CLK(net323),
    .RESET_B(_0092_),
    .D(_0071_),
    .Q_N(_0828_),
    .Q(\stop.syn.adsr_data[8] ));
 sg13g2_dfrbp_1 _1835_ (.CLK(net323),
    .RESET_B(_0093_),
    .D(_0072_),
    .Q_N(_0827_),
    .Q(\stop.syn.adsr_data[9] ));
 sg13g2_dfrbp_1 _1836_ (.CLK(net324),
    .RESET_B(_0094_),
    .D(_0073_),
    .Q_N(_0826_),
    .Q(\stop.syn.adsr_data[10] ));
 sg13g2_dfrbp_1 _1837_ (.CLK(net324),
    .RESET_B(_0095_),
    .D(_0074_),
    .Q_N(_0043_),
    .Q(\stop.syn.adsr_data[11] ));
 sg13g2_dfrbp_1 _1838_ (.CLK(net324),
    .RESET_B(_0096_),
    .D(_0075_),
    .Q_N(_0825_),
    .Q(\stop.syn.adsr_data[12] ));
 sg13g2_dfrbp_1 _1839_ (.CLK(net320),
    .RESET_B(_0097_),
    .D(_0076_),
    .Q_N(_0044_),
    .Q(\stop.syn.adsr_data[13] ));
 sg13g2_dfrbp_1 _1840_ (.CLK(net320),
    .RESET_B(_0098_),
    .D(_0077_),
    .Q_N(_0824_),
    .Q(\stop.syn.adsr_data[14] ));
 sg13g2_dfrbp_1 _1841_ (.CLK(net320),
    .RESET_B(_0099_),
    .D(_0069_),
    .Q_N(_0823_),
    .Q(\stop.syn.adsr_data[15] ));
 sg13g2_dfrbp_1 _1842_ (.CLK(net325),
    .RESET_B(_0100_),
    .D(\stop.syn.filt.m2.sum[1] ),
    .Q_N(_0822_),
    .Q(\stop.syn.filt.m2.sum_in2[0] ));
 sg13g2_dfrbp_1 _1843_ (.CLK(net326),
    .RESET_B(_0101_),
    .D(\stop.syn.filt.m2.sum[2] ),
    .Q_N(_0821_),
    .Q(\stop.syn.filt.m2.sum_in2[1] ));
 sg13g2_dfrbp_1 _1844_ (.CLK(net325),
    .RESET_B(_0102_),
    .D(\stop.syn.filt.m2.sum[3] ),
    .Q_N(_0820_),
    .Q(\stop.syn.filt.m2.sum_in2[2] ));
 sg13g2_dfrbp_1 _1845_ (.CLK(net324),
    .RESET_B(_0103_),
    .D(\stop.syn.filt.m2.sum[4] ),
    .Q_N(_0050_),
    .Q(\stop.syn.filt.m2.sum_in2[3] ));
 sg13g2_dfrbp_1 _1846_ (.CLK(net323),
    .RESET_B(_0104_),
    .D(\stop.syn.filt.m2.sum[5] ),
    .Q_N(_0819_),
    .Q(\stop.syn.filt.m2.sum_in2[4] ));
 sg13g2_dfrbp_1 _1847_ (.CLK(net324),
    .RESET_B(_0105_),
    .D(\stop.syn.filt.m2.sum[6] ),
    .Q_N(_0051_),
    .Q(\stop.syn.filt.m2.sum_in2[5] ));
 sg13g2_dfrbp_1 _1848_ (.CLK(net325),
    .RESET_B(_0106_),
    .D(\stop.syn.filt.m2.sum[7] ),
    .Q_N(_0818_),
    .Q(\stop.syn.filt.m2.sum_in2[6] ));
 sg13g2_dfrbp_1 _1849_ (.CLK(net325),
    .RESET_B(_0107_),
    .D(\stop.syn.filt.m2.sum[8] ),
    .Q_N(_0817_),
    .Q(\stop.syn.filt.m2.sum_in2[7] ));
 sg13g2_dfrbp_1 _1850_ (.CLK(net325),
    .RESET_B(_0108_),
    .D(\stop.syn.filt.m2.sum[9] ),
    .Q_N(_0816_),
    .Q(\stop.syn.filt.m2.sum_in2[8] ));
 sg13g2_dfrbp_1 _1851_ (.CLK(net326),
    .RESET_B(_0109_),
    .D(\stop.syn.filt.m2.sum[10] ),
    .Q_N(_0052_),
    .Q(\stop.syn.filt.m2.sum_in2[9] ));
 sg13g2_dfrbp_1 _1852_ (.CLK(net326),
    .RESET_B(_0110_),
    .D(\stop.syn.filt.m2.sum[11] ),
    .Q_N(_0815_),
    .Q(\stop.syn.filt.m2.sum_in2[10] ));
 sg13g2_dfrbp_1 _1853_ (.CLK(net326),
    .RESET_B(_0111_),
    .D(\stop.syn.filt.m2.sum[12] ),
    .Q_N(_0814_),
    .Q(\stop.syn.filt.m2.sum_in2[11] ));
 sg13g2_dfrbp_1 _1854_ (.CLK(net326),
    .RESET_B(_0112_),
    .D(\stop.syn.filt.m2.sum[13] ),
    .Q_N(_0813_),
    .Q(\stop.syn.filt.m2.sum_in2[12] ));
 sg13g2_dfrbp_1 _1855_ (.CLK(net326),
    .RESET_B(_0113_),
    .D(\stop.syn.filt.m2.sum[14] ),
    .Q_N(_0042_),
    .Q(\stop.syn.filt.m2.sum_in2[13] ));
 sg13g2_dfrbp_1 _1856_ (.CLK(net327),
    .RESET_B(_0114_),
    .D(\stop.syn.filt.m2.sum[15] ),
    .Q_N(_0812_),
    .Q(\stop.syn.filt.m2.sum_in2[14] ));
 sg13g2_dfrbp_1 _1857_ (.CLK(net321),
    .RESET_B(_0115_),
    .D(\stop.syn.filt.m2.sum[16] ),
    .Q_N(_0811_),
    .Q(\stop.syn.filt.m2.sum_in2[15] ));
 sg13g2_dfrbp_1 _1858_ (.CLK(net329),
    .RESET_B(_0116_),
    .D(\stop.syn.filt.m1.sum[1] ),
    .Q_N(_0810_),
    .Q(\stop.syn.filt.m1.sum_in2[0] ));
 sg13g2_dfrbp_1 _1859_ (.CLK(net329),
    .RESET_B(_0117_),
    .D(\stop.syn.filt.m1.sum[2] ),
    .Q_N(_0809_),
    .Q(\stop.syn.filt.m1.sum_in2[1] ));
 sg13g2_dfrbp_1 _1860_ (.CLK(net328),
    .RESET_B(_0118_),
    .D(\stop.syn.filt.m1.sum[3] ),
    .Q_N(_0808_),
    .Q(\stop.syn.filt.m1.sum_in2[2] ));
 sg13g2_dfrbp_1 _1861_ (.CLK(net328),
    .RESET_B(_0119_),
    .D(\stop.syn.filt.m1.sum[4] ),
    .Q_N(_0046_),
    .Q(\stop.syn.filt.m1.sum_in2[3] ));
 sg13g2_dfrbp_1 _1862_ (.CLK(net329),
    .RESET_B(_0120_),
    .D(\stop.syn.filt.m1.sum[5] ),
    .Q_N(_0807_),
    .Q(\stop.syn.filt.m1.sum_in2[4] ));
 sg13g2_dfrbp_1 _1863_ (.CLK(net328),
    .RESET_B(_0121_),
    .D(\stop.syn.filt.m1.sum[6] ),
    .Q_N(_0047_),
    .Q(\stop.syn.filt.m1.sum_in2[5] ));
 sg13g2_dfrbp_1 _1864_ (.CLK(net326),
    .RESET_B(_0122_),
    .D(\stop.syn.filt.m1.sum[7] ),
    .Q_N(_0806_),
    .Q(\stop.syn.filt.m1.sum_in2[6] ));
 sg13g2_dfrbp_1 _1865_ (.CLK(net325),
    .RESET_B(_0123_),
    .D(\stop.syn.filt.m1.sum[8] ),
    .Q_N(_0805_),
    .Q(\stop.syn.filt.m1.sum_in2[7] ));
 sg13g2_dfrbp_1 _1866_ (.CLK(net328),
    .RESET_B(_0124_),
    .D(\stop.syn.filt.m1.sum[9] ),
    .Q_N(_0804_),
    .Q(\stop.syn.filt.m1.sum_in2[8] ));
 sg13g2_dfrbp_1 _1867_ (.CLK(net328),
    .RESET_B(_0125_),
    .D(\stop.syn.filt.m1.sum[10] ),
    .Q_N(_0048_),
    .Q(\stop.syn.filt.m1.sum_in2[9] ));
 sg13g2_dfrbp_1 _1868_ (.CLK(net328),
    .RESET_B(_0126_),
    .D(\stop.syn.filt.m1.sum[11] ),
    .Q_N(_0803_),
    .Q(\stop.syn.filt.m1.sum_in2[10] ));
 sg13g2_dfrbp_1 _1869_ (.CLK(net328),
    .RESET_B(_0127_),
    .D(\stop.syn.filt.m1.sum[12] ),
    .Q_N(_0802_),
    .Q(\stop.syn.filt.m1.sum_in2[11] ));
 sg13g2_dfrbp_1 _1870_ (.CLK(net329),
    .RESET_B(_0128_),
    .D(\stop.syn.filt.m1.sum[13] ),
    .Q_N(_0801_),
    .Q(\stop.syn.filt.m1.sum_in2[12] ));
 sg13g2_dfrbp_1 _1871_ (.CLK(net328),
    .RESET_B(_0129_),
    .D(\stop.syn.filt.m1.sum[14] ),
    .Q_N(_0049_),
    .Q(\stop.syn.filt.m1.sum_in2[13] ));
 sg13g2_dfrbp_1 _1872_ (.CLK(net330),
    .RESET_B(_0130_),
    .D(\stop.syn.filt.m1.sum[15] ),
    .Q_N(_0800_),
    .Q(\stop.syn.filt.m1.sum_in2[14] ));
 sg13g2_dfrbp_1 _1873_ (.CLK(net330),
    .RESET_B(_0131_),
    .D(\stop.syn.filt.m1.sum[16] ),
    .Q_N(_0907_),
    .Q(\stop.syn.filt.m1.sum_in2[15] ));
 sg13g2_dfrbp_1 _1874_ (.CLK(net304),
    .RESET_B(net334),
    .D(_0053_),
    .Q_N(_0908_),
    .Q(\stop.dbg_adsr_filt0 ));
 sg13g2_dfrbp_1 _1875_ (.CLK(net304),
    .RESET_B(net332),
    .D(_0060_),
    .Q_N(_0909_),
    .Q(\stop.syn.daci.din[1] ));
 sg13g2_dfrbp_1 _1876_ (.CLK(net304),
    .RESET_B(net334),
    .D(_0061_),
    .Q_N(_0910_),
    .Q(\stop.syn.daci.din[2] ));
 sg13g2_dfrbp_1 _1877_ (.CLK(net304),
    .RESET_B(net334),
    .D(_0062_),
    .Q_N(_0911_),
    .Q(\stop.syn.daci.din[3] ));
 sg13g2_dfrbp_1 _1878_ (.CLK(net303),
    .RESET_B(net332),
    .D(_0063_),
    .Q_N(_0912_),
    .Q(\stop.syn.daci.din[4] ));
 sg13g2_dfrbp_1 _1879_ (.CLK(net303),
    .RESET_B(net332),
    .D(_0064_),
    .Q_N(_0913_),
    .Q(\stop.syn.daci.din[5] ));
 sg13g2_dfrbp_1 _1880_ (.CLK(net303),
    .RESET_B(net332),
    .D(_0065_),
    .Q_N(_0914_),
    .Q(\stop.syn.daci.din[6] ));
 sg13g2_dfrbp_1 _1881_ (.CLK(net303),
    .RESET_B(net332),
    .D(_0066_),
    .Q_N(_0915_),
    .Q(\stop.syn.daci.din[7] ));
 sg13g2_dfrbp_1 _1882_ (.CLK(net303),
    .RESET_B(net332),
    .D(_0067_),
    .Q_N(_0916_),
    .Q(\stop.syn.daci.din[8] ));
 sg13g2_dfrbp_1 _1883_ (.CLK(net303),
    .RESET_B(net332),
    .D(_0068_),
    .Q_N(_0917_),
    .Q(\stop.syn.daci.din[9] ));
 sg13g2_dfrbp_1 _1884_ (.CLK(net305),
    .RESET_B(net333),
    .D(_0054_),
    .Q_N(_0918_),
    .Q(\stop.syn.daci.din[10] ));
 sg13g2_dfrbp_1 _1885_ (.CLK(net305),
    .RESET_B(net333),
    .D(_0055_),
    .Q_N(_0919_),
    .Q(\stop.syn.daci.din[11] ));
 sg13g2_dfrbp_1 _1886_ (.CLK(net305),
    .RESET_B(net333),
    .D(_0056_),
    .Q_N(_0920_),
    .Q(\stop.syn.daci.din[12] ));
 sg13g2_dfrbp_1 _1887_ (.CLK(net305),
    .RESET_B(net333),
    .D(_0057_),
    .Q_N(_0921_),
    .Q(\stop.syn.daci.din[13] ));
 sg13g2_dfrbp_1 _1888_ (.CLK(net305),
    .RESET_B(net333),
    .D(_0058_),
    .Q_N(_0922_),
    .Q(\stop.syn.daci.din[14] ));
 sg13g2_dfrbp_1 _1889_ (.CLK(net305),
    .RESET_B(net333),
    .D(_0059_),
    .Q_N(_0799_),
    .Q(\stop.syn.daci.din[15] ));
 sg13g2_dfrbp_1 _1890_ (.CLK(net319),
    .RESET_B(net44),
    .D(_0155_),
    .Q_N(_0798_),
    .Q(\stop.syn.filt.m1.b_latched[7] ));
 sg13g2_dfrbp_1 _1891_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net43),
    .D(_0156_),
    .Q_N(_0797_),
    .Q(\stop.syn.daci.accumulator[0] ));
 sg13g2_dfrbp_1 _1892_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net42),
    .D(net110),
    .Q_N(_0796_),
    .Q(\stop.syn.daci.accumulator[1] ));
 sg13g2_dfrbp_1 _1893_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net41),
    .D(net126),
    .Q_N(_0795_),
    .Q(\stop.syn.daci.accumulator[2] ));
 sg13g2_dfrbp_1 _1894_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net40),
    .D(_0159_),
    .Q_N(_0794_),
    .Q(\stop.syn.daci.accumulator[3] ));
 sg13g2_dfrbp_1 _1895_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net39),
    .D(net130),
    .Q_N(_0793_),
    .Q(\stop.syn.daci.accumulator[4] ));
 sg13g2_dfrbp_1 _1896_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net38),
    .D(net122),
    .Q_N(_0792_),
    .Q(\stop.syn.daci.accumulator[5] ));
 sg13g2_dfrbp_1 _1897_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net37),
    .D(_0162_),
    .Q_N(_0791_),
    .Q(\stop.syn.daci.accumulator[6] ));
 sg13g2_dfrbp_1 _1898_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net36),
    .D(_0163_),
    .Q_N(_0790_),
    .Q(\stop.syn.daci.accumulator[7] ));
 sg13g2_dfrbp_1 _1899_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net35),
    .D(net118),
    .Q_N(_0789_),
    .Q(\stop.syn.daci.accumulator[8] ));
 sg13g2_dfrbp_1 _1900_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net34),
    .D(_0165_),
    .Q_N(_0788_),
    .Q(\stop.syn.daci.accumulator[9] ));
 sg13g2_dfrbp_1 _1901_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net33),
    .D(net114),
    .Q_N(_0787_),
    .Q(\stop.syn.daci.accumulator[10] ));
 sg13g2_dfrbp_1 _1902_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net32),
    .D(_0167_),
    .Q_N(_0786_),
    .Q(\stop.syn.daci.accumulator[11] ));
 sg13g2_dfrbp_1 _1903_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net31),
    .D(_0168_),
    .Q_N(_0785_),
    .Q(\stop.syn.daci.accumulator[12] ));
 sg13g2_dfrbp_1 _1904_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net30),
    .D(_0169_),
    .Q_N(_0784_),
    .Q(\stop.syn.daci.accumulator[13] ));
 sg13g2_dfrbp_1 _1905_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net29),
    .D(_0170_),
    .Q_N(_0783_),
    .Q(\stop.syn.daci.accumulator[14] ));
 sg13g2_dfrbp_1 _1906_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net16),
    .D(_0171_),
    .Q_N(_0782_),
    .Q(\stop.syn.daci.accumulator[15] ));
 sg13g2_dfrbp_1 _1907_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net89),
    .D(_0172_),
    .Q_N(_0781_),
    .Q(data));
 sg13g2_dfrbp_1 _1908_ (.CLK(net356),
    .RESET_B(net367),
    .D(_0173_),
    .Q_N(_0780_),
    .Q(\stop.adsr_ai[0] ));
 sg13g2_dfrbp_1 _1909_ (.CLK(net358),
    .RESET_B(net369),
    .D(_0174_),
    .Q_N(_0779_),
    .Q(\stop.adsr_ai[1] ));
 sg13g2_dfrbp_1 _1910_ (.CLK(net357),
    .RESET_B(net368),
    .D(_0175_),
    .Q_N(_0778_),
    .Q(\stop.adsr_ai[2] ));
 sg13g2_dfrbp_1 _1911_ (.CLK(net357),
    .RESET_B(net368),
    .D(_0176_),
    .Q_N(_0777_),
    .Q(\stop.adsr_ai[3] ));
 sg13g2_dfrbp_1 _1912_ (.CLK(net356),
    .RESET_B(net367),
    .D(_0177_),
    .Q_N(_0776_),
    .Q(\stop.adsr_ai[4] ));
 sg13g2_dfrbp_1 _1913_ (.CLK(net355),
    .RESET_B(net366),
    .D(_0178_),
    .Q_N(_0775_),
    .Q(\stop.adsr_ai[5] ));
 sg13g2_dfrbp_1 _1914_ (.CLK(net354),
    .RESET_B(net365),
    .D(_0179_),
    .Q_N(_0774_),
    .Q(\stop.adsr_ai[6] ));
 sg13g2_dfrbp_1 _1915_ (.CLK(net354),
    .RESET_B(net365),
    .D(_0180_),
    .Q_N(_0773_),
    .Q(\stop.adsr_ai[7] ));
 sg13g2_dfrbp_1 _1916_ (.CLK(net355),
    .RESET_B(net366),
    .D(_0181_),
    .Q_N(_0772_),
    .Q(\stop.adsr_di[0] ));
 sg13g2_dfrbp_1 _1917_ (.CLK(net356),
    .RESET_B(net367),
    .D(_0182_),
    .Q_N(_0771_),
    .Q(\stop.adsr_di[1] ));
 sg13g2_dfrbp_1 _1918_ (.CLK(net356),
    .RESET_B(net367),
    .D(_0183_),
    .Q_N(_0770_),
    .Q(\stop.adsr_di[2] ));
 sg13g2_dfrbp_1 _1919_ (.CLK(net356),
    .RESET_B(net367),
    .D(_0184_),
    .Q_N(_0769_),
    .Q(\stop.adsr_di[3] ));
 sg13g2_dfrbp_1 _1920_ (.CLK(net355),
    .RESET_B(net366),
    .D(_0185_),
    .Q_N(_0768_),
    .Q(\stop.adsr_di[4] ));
 sg13g2_dfrbp_1 _1921_ (.CLK(net354),
    .RESET_B(net365),
    .D(_0186_),
    .Q_N(_0767_),
    .Q(\stop.adsr_di[5] ));
 sg13g2_dfrbp_1 _1922_ (.CLK(net354),
    .RESET_B(net365),
    .D(_0187_),
    .Q_N(_0766_),
    .Q(\stop.adsr_di[6] ));
 sg13g2_dfrbp_1 _1923_ (.CLK(net354),
    .RESET_B(net365),
    .D(_0188_),
    .Q_N(_0765_),
    .Q(\stop.adsr_di[7] ));
 sg13g2_dfrbp_1 _1924_ (.CLK(net354),
    .RESET_B(net365),
    .D(_0189_),
    .Q_N(_0764_),
    .Q(\stop.adsr_s[0] ));
 sg13g2_dfrbp_1 _1925_ (.CLK(net356),
    .RESET_B(net367),
    .D(_0190_),
    .Q_N(_0763_),
    .Q(\stop.adsr_s[1] ));
 sg13g2_dfrbp_1 _1926_ (.CLK(net358),
    .RESET_B(net369),
    .D(_0191_),
    .Q_N(_0762_),
    .Q(\stop.adsr_s[2] ));
 sg13g2_dfrbp_1 _1927_ (.CLK(net358),
    .RESET_B(net369),
    .D(_0192_),
    .Q_N(_0761_),
    .Q(\stop.adsr_s[3] ));
 sg13g2_dfrbp_1 _1928_ (.CLK(net357),
    .RESET_B(net368),
    .D(_0193_),
    .Q_N(_0760_),
    .Q(\stop.adsr_s[4] ));
 sg13g2_dfrbp_1 _1929_ (.CLK(net357),
    .RESET_B(net368),
    .D(_0194_),
    .Q_N(_0759_),
    .Q(\stop.adsr_s[5] ));
 sg13g2_dfrbp_1 _1930_ (.CLK(net357),
    .RESET_B(net368),
    .D(_0195_),
    .Q_N(_0758_),
    .Q(\stop.adsr_s[6] ));
 sg13g2_dfrbp_1 _1931_ (.CLK(net357),
    .RESET_B(net368),
    .D(_0196_),
    .Q_N(_0757_),
    .Q(\stop.adsr_s[7] ));
 sg13g2_dfrbp_1 _1932_ (.CLK(net358),
    .RESET_B(net369),
    .D(_0197_),
    .Q_N(_0756_),
    .Q(\stop.adsr_ri[0] ));
 sg13g2_dfrbp_1 _1933_ (.CLK(net357),
    .RESET_B(net368),
    .D(_0198_),
    .Q_N(_0755_),
    .Q(\stop.adsr_ri[1] ));
 sg13g2_dfrbp_1 _1934_ (.CLK(net357),
    .RESET_B(net368),
    .D(_0199_),
    .Q_N(_0754_),
    .Q(\stop.adsr_ri[2] ));
 sg13g2_dfrbp_1 _1935_ (.CLK(net356),
    .RESET_B(net367),
    .D(_0200_),
    .Q_N(_0753_),
    .Q(\stop.adsr_ri[3] ));
 sg13g2_dfrbp_1 _1936_ (.CLK(net356),
    .RESET_B(net367),
    .D(_0201_),
    .Q_N(_0752_),
    .Q(\stop.adsr_ri[4] ));
 sg13g2_dfrbp_1 _1937_ (.CLK(net354),
    .RESET_B(net365),
    .D(_0202_),
    .Q_N(_0751_),
    .Q(\stop.adsr_ri[5] ));
 sg13g2_dfrbp_1 _1938_ (.CLK(net354),
    .RESET_B(net365),
    .D(_0203_),
    .Q_N(_0750_),
    .Q(\stop.adsr_ri[6] ));
 sg13g2_dfrbp_1 _1939_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0204_),
    .Q_N(_0749_),
    .Q(\stop.adsr_ri[7] ));
 sg13g2_dfrbp_1 _1940_ (.CLK(net352),
    .RESET_B(net363),
    .D(_0205_),
    .Q_N(_0748_),
    .Q(\stop.ctrl.cfg[32] ));
 sg13g2_dfrbp_1 _1941_ (.CLK(net352),
    .RESET_B(net363),
    .D(_0206_),
    .Q_N(_0747_),
    .Q(\stop.ctrl.cfg[33] ));
 sg13g2_dfrbp_1 _1942_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0207_),
    .Q_N(_0746_),
    .Q(\stop.ctrl.cfg[34] ));
 sg13g2_dfrbp_1 _1943_ (.CLK(net353),
    .RESET_B(net364),
    .D(_0208_),
    .Q_N(_0745_),
    .Q(\stop.ctrl.cfg[35] ));
 sg13g2_dfrbp_1 _1944_ (.CLK(net353),
    .RESET_B(net364),
    .D(_0209_),
    .Q_N(_0744_),
    .Q(\stop.ctrl.cfg[36] ));
 sg13g2_dfrbp_1 _1945_ (.CLK(net353),
    .RESET_B(net364),
    .D(_0210_),
    .Q_N(_0743_),
    .Q(\stop.ctrl.cfg[37] ));
 sg13g2_dfrbp_1 _1946_ (.CLK(net353),
    .RESET_B(net364),
    .D(_0211_),
    .Q_N(_0742_),
    .Q(\stop.ctrl.cfg[38] ));
 sg13g2_dfrbp_1 _1947_ (.CLK(net353),
    .RESET_B(net364),
    .D(_0212_),
    .Q_N(_0741_),
    .Q(\stop.ctrl.cfg[39] ));
 sg13g2_dfrbp_1 _1948_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0213_),
    .Q_N(_0740_),
    .Q(\stop.ctrl.cfg[40] ));
 sg13g2_dfrbp_1 _1949_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0214_),
    .Q_N(_0739_),
    .Q(\stop.ctrl.cfg[41] ));
 sg13g2_dfrbp_1 _1950_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0215_),
    .Q_N(_0738_),
    .Q(\stop.ctrl.cfg[42] ));
 sg13g2_dfrbp_1 _1951_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0216_),
    .Q_N(_0737_),
    .Q(\stop.ctrl.cfg[43] ));
 sg13g2_dfrbp_1 _1952_ (.CLK(net350),
    .RESET_B(net361),
    .D(_0217_),
    .Q_N(_0736_),
    .Q(\stop.ctrl.cfg[44] ));
 sg13g2_dfrbp_1 _1953_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0218_),
    .Q_N(_0735_),
    .Q(\stop.ctrl.cfg[45] ));
 sg13g2_dfrbp_1 _1954_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0219_),
    .Q_N(_0734_),
    .Q(\stop.ctrl.cfg[46] ));
 sg13g2_dfrbp_1 _1955_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0220_),
    .Q_N(_0733_),
    .Q(\stop.ctrl.cfg[47] ));
 sg13g2_dfrbp_1 _1956_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0221_),
    .Q_N(_0732_),
    .Q(\stop.ctrl.cfg[48] ));
 sg13g2_dfrbp_1 _1957_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0222_),
    .Q_N(_0731_),
    .Q(\stop.ctrl.cfg[49] ));
 sg13g2_dfrbp_1 _1958_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0223_),
    .Q_N(_0730_),
    .Q(\stop.ctrl.cfg[50] ));
 sg13g2_dfrbp_1 _1959_ (.CLK(net349),
    .RESET_B(net360),
    .D(_0224_),
    .Q_N(_0729_),
    .Q(\stop.ctrl.cfg[51] ));
 sg13g2_dfrbp_1 _1960_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0225_),
    .Q_N(_0728_),
    .Q(\stop.ctrl.cfg[52] ));
 sg13g2_dfrbp_1 _1961_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0226_),
    .Q_N(_0727_),
    .Q(\stop.ctrl.cfg[53] ));
 sg13g2_dfrbp_1 _1962_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0227_),
    .Q_N(_0726_),
    .Q(\stop.ctrl.cfg[54] ));
 sg13g2_dfrbp_1 _1963_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0228_),
    .Q_N(_0725_),
    .Q(\stop.ctrl.cfg[55] ));
 sg13g2_dfrbp_1 _1964_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0229_),
    .Q_N(_0724_),
    .Q(\stop.ctrl.cfg[56] ));
 sg13g2_dfrbp_1 _1965_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0230_),
    .Q_N(_0723_),
    .Q(\stop.ctrl.cfg[57] ));
 sg13g2_dfrbp_1 _1966_ (.CLK(net351),
    .RESET_B(net362),
    .D(_0231_),
    .Q_N(_0722_),
    .Q(\stop.ctrl.cfg[58] ));
 sg13g2_dfrbp_1 _1967_ (.CLK(net359),
    .RESET_B(net370),
    .D(_0232_),
    .Q_N(_0721_),
    .Q(\stop.ctrl.cfg[59] ));
 sg13g2_tiehi _1749__17 (.L_HI(net17));
 sg13g2_tiehi _1748__18 (.L_HI(net18));
 sg13g2_tiehi _1742__19 (.L_HI(net19));
 sg13g2_tiehi _1741__20 (.L_HI(net20));
 sg13g2_tiehi _1740__21 (.L_HI(net21));
 sg13g2_tiehi _1739__22 (.L_HI(net22));
 sg13g2_tiehi _1737__23 (.L_HI(net23));
 sg13g2_tiehi _1743__24 (.L_HI(net24));
 sg13g2_tiehi _1744__25 (.L_HI(net25));
 sg13g2_tiehi _1745__26 (.L_HI(net26));
 sg13g2_tiehi _1746__27 (.L_HI(net27));
 sg13g2_tiehi _1738__28 (.L_HI(net28));
 sg13g2_tiehi _1905__29 (.L_HI(net29));
 sg13g2_tiehi _1904__30 (.L_HI(net30));
 sg13g2_tiehi _1903__31 (.L_HI(net31));
 sg13g2_tiehi _1902__32 (.L_HI(net32));
 sg13g2_tiehi _1901__33 (.L_HI(net33));
 sg13g2_tiehi _1900__34 (.L_HI(net34));
 sg13g2_tiehi _1899__35 (.L_HI(net35));
 sg13g2_tiehi _1898__36 (.L_HI(net36));
 sg13g2_tiehi _1897__37 (.L_HI(net37));
 sg13g2_tiehi _1896__38 (.L_HI(net38));
 sg13g2_tiehi _1895__39 (.L_HI(net39));
 sg13g2_tiehi _1894__40 (.L_HI(net40));
 sg13g2_tiehi _1893__41 (.L_HI(net41));
 sg13g2_tiehi _1892__42 (.L_HI(net42));
 sg13g2_tiehi _1891__43 (.L_HI(net43));
 sg13g2_tiehi _1890__44 (.L_HI(net44));
 sg13g2_tiehi _1747__45 (.L_HI(net45));
 sg13g2_tiehi _1778__46 (.L_HI(net46));
 sg13g2_tiehi _1779__47 (.L_HI(net47));
 sg13g2_tiehi _1780__48 (.L_HI(net48));
 sg13g2_tiehi _1781__49 (.L_HI(net49));
 sg13g2_tiehi _1782__50 (.L_HI(net50));
 sg13g2_tiehi _1783__51 (.L_HI(net51));
 sg13g2_tiehi _1784__52 (.L_HI(net52));
 sg13g2_tiehi _1785__53 (.L_HI(net53));
 sg13g2_tiehi _1786__54 (.L_HI(net54));
 sg13g2_tiehi _1787__55 (.L_HI(net55));
 sg13g2_tiehi _1788__56 (.L_HI(net56));
 sg13g2_tiehi _1789__57 (.L_HI(net57));
 sg13g2_tiehi _1790__58 (.L_HI(net58));
 sg13g2_tiehi _1791__59 (.L_HI(net59));
 sg13g2_tiehi _1792__60 (.L_HI(net60));
 sg13g2_tiehi _1793__61 (.L_HI(net61));
 sg13g2_tiehi _1794__62 (.L_HI(net62));
 sg13g2_tiehi _1795__63 (.L_HI(net63));
 sg13g2_tiehi _1796__64 (.L_HI(net64));
 sg13g2_tiehi _1797__65 (.L_HI(net65));
 sg13g2_tiehi _1798__66 (.L_HI(net66));
 sg13g2_tiehi _1799__67 (.L_HI(net67));
 sg13g2_tiehi _1800__68 (.L_HI(net68));
 sg13g2_tiehi _1825__69 (.L_HI(net69));
 sg13g2_tiehi _1824__70 (.L_HI(net70));
 sg13g2_tiehi _1823__71 (.L_HI(net71));
 sg13g2_tiehi _1822__72 (.L_HI(net72));
 sg13g2_tiehi _1821__73 (.L_HI(net73));
 sg13g2_tiehi _1820__74 (.L_HI(net74));
 sg13g2_tiehi _1819__75 (.L_HI(net75));
 sg13g2_tiehi _1818__76 (.L_HI(net76));
 sg13g2_tiehi _1817__77 (.L_HI(net77));
 sg13g2_tiehi _1777__78 (.L_HI(net78));
 sg13g2_tiehi _1776__79 (.L_HI(net79));
 sg13g2_tiehi _1775__80 (.L_HI(net80));
 sg13g2_tiehi _1774__81 (.L_HI(net81));
 sg13g2_tiehi _1773__82 (.L_HI(net82));
 sg13g2_tiehi _1772__83 (.L_HI(net83));
 sg13g2_tiehi _1771__84 (.L_HI(net84));
 sg13g2_tiehi _1770__85 (.L_HI(net85));
 sg13g2_tiehi _1769__86 (.L_HI(net86));
 sg13g2_tiehi _1768__87 (.L_HI(net87));
 sg13g2_tiehi _1767__88 (.L_HI(net88));
 sg13g2_tiehi _1907__89 (.L_HI(net89));
 sg13g2_tiehi _1763__90 (.L_HI(net90));
 sg13g2_tiehi _1762__91 (.L_HI(net91));
 sg13g2_tiehi _1761__92 (.L_HI(net92));
 sg13g2_tiehi _1760__93 (.L_HI(net93));
 sg13g2_tiehi _1759__94 (.L_HI(net94));
 sg13g2_tiehi _1758__95 (.L_HI(net95));
 sg13g2_tiehi _1757__96 (.L_HI(net96));
 sg13g2_tiehi _1756__97 (.L_HI(net97));
 sg13g2_tiehi _1755__98 (.L_HI(net98));
 sg13g2_tiehi _1754__99 (.L_HI(net99));
 sg13g2_tiehi _1753__100 (.L_HI(net100));
 sg13g2_tiehi _1752__101 (.L_HI(net101));
 sg13g2_tiehi _1751__102 (.L_HI(net102));
 sg13g2_tiehi _1750__103 (.L_HI(net103));
 sg13g2_tiehi tt_um_jp_cd101_saw_104 (.L_HI(net104));
 sg13g2_tiehi tt_um_jp_cd101_saw_105 (.L_HI(net105));
 sg13g2_tiehi _1766__106 (.L_HI(net106));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_jp_cd101_saw_5 (.L_LO(net5));
 sg13g2_tielo tt_um_jp_cd101_saw_6 (.L_LO(net6));
 sg13g2_tielo tt_um_jp_cd101_saw_7 (.L_LO(net7));
 sg13g2_tielo tt_um_jp_cd101_saw_8 (.L_LO(net8));
 sg13g2_tielo tt_um_jp_cd101_saw_9 (.L_LO(net9));
 sg13g2_tielo tt_um_jp_cd101_saw_10 (.L_LO(net10));
 sg13g2_tielo tt_um_jp_cd101_saw_11 (.L_LO(net11));
 sg13g2_tielo tt_um_jp_cd101_saw_12 (.L_LO(net12));
 sg13g2_tielo tt_um_jp_cd101_saw_13 (.L_LO(net13));
 sg13g2_tielo tt_um_jp_cd101_saw_14 (.L_LO(net14));
 sg13g2_tielo tt_um_jp_cd101_saw_15 (.L_LO(net15));
 sg13g2_tiehi _1906__16 (.L_HI(net16));
 sg13g2_buf_1 _2071_ (.A(\stop.dbg_adsr_filt0 ),
    .X(uio_out[0]));
 sg13g2_buf_1 _2072_ (.A(\stop.dbg_adsr_reg0 ),
    .X(uio_out[1]));
 sg13g2_buf_1 _2073_ (.A(\stop.dbg_adsr0 ),
    .X(uo_out[0]));
 sg13g2_buf_2 _2074_ (.A(\stop.dbg_env0 ),
    .X(uo_out[1]));
 sg13g2_buf_2 _2075_ (.A(\stop.dbg_osc0 ),
    .X(uo_out[2]));
 sg13g2_buf_2 _2076_ (.A(net287),
    .X(uo_out[3]));
 sg13g2_buf_1 _2077_ (.A(net303),
    .X(uo_out[4]));
 sg13g2_buf_1 _2078_ (.A(\stop.dbg_trig ),
    .X(uo_out[5]));
 sg13g2_buf_1 _2079_ (.A(net332),
    .X(uo_out[6]));
 sg13g2_buf_2 _2080_ (.A(data),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(\stop.syn.adsri.rstn ));
 sg13g2_buf_2 fanout278 (.A(net279),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(\stop.syn.adsri.rstn ),
    .X(net281));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(\stop.syn.adsri.state[2] ));
 sg13g2_buf_2 fanout283 (.A(\stop.syn.adsri.state[1] ),
    .X(net283));
 sg13g2_buf_1 fanout284 (.A(\stop.syn.adsri.state[1] ),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(net286),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(net287),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(\stop.dbg_clk_adsr ),
    .X(net287));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(net289));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(net294));
 sg13g2_buf_2 fanout290 (.A(net291),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(net294),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(net294),
    .X(net292));
 sg13g2_buf_1 fanout293 (.A(net294),
    .X(net293));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(_0327_));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(net298));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(net297));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(net298));
 sg13g2_buf_2 fanout298 (.A(_0327_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(net300),
    .X(net299));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(net306));
 sg13g2_buf_2 fanout301 (.A(net302),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(net306),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(net305),
    .X(net303));
 sg13g2_buf_1 fanout304 (.A(net305),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(\stop.dbg_clk_sample ),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(\stop.syn.smul8.b_bit ),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(\stop.syn.smul8.b_bit ),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(net313),
    .X(net309));
 sg13g2_buf_1 fanout310 (.A(net313),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(net312),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net313),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(\stop.syn.filt.m1.b_bit ),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(net315),
    .X(net314));
 sg13g2_buf_1 fanout315 (.A(net318),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(\stop.syn.filt.m2.b_bit ),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net322),
    .X(net319));
 sg13g2_buf_1 fanout320 (.A(net322),
    .X(net320));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(net322));
 sg13g2_buf_2 fanout322 (.A(net331),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(net331),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(net326),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(net331),
    .X(net326));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(net330));
 sg13g2_buf_2 fanout328 (.A(net329),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(net330),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(net331),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_0037_),
    .X(net331));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(net334));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(\stop.dbg_rstn ));
 sg13g2_buf_2 fanout334 (.A(\stop.dbg_rstn ),
    .X(net334));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(net337));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(net337));
 sg13g2_buf_2 fanout337 (.A(net346),
    .X(net337));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(net346));
 sg13g2_buf_2 fanout339 (.A(net340),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(net345),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(net343),
    .X(net341));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(net344));
 sg13g2_buf_1 fanout343 (.A(net344),
    .X(net343));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(net345));
 sg13g2_buf_2 fanout345 (.A(net346),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_0307_),
    .X(net346));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(\stop.syn.clki.arstn ));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(\stop.syn.clki.arstn ));
 sg13g2_buf_2 fanout349 (.A(net352),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(net352),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(uio_in[3]),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(net355),
    .X(net354));
 sg13g2_buf_1 fanout355 (.A(net359),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(net358),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(net359),
    .X(net358));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(uio_in[3]));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(net363));
 sg13g2_buf_2 fanout361 (.A(net363),
    .X(net361));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(net363));
 sg13g2_buf_2 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(rst_n));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(net366));
 sg13g2_buf_2 fanout366 (.A(net370),
    .X(net366));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(net369));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(net369));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(net370));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(uio_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(uio_in[1]),
    .X(net3));
 sg13g2_tielo tt_um_jp_cd101_saw_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0027_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold2 (.A(\stop.syn.rstn_fst_reg1 ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold3 (.A(\stop.syn.daci.accumulator[0] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0157_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold5 (.A(\stop.syn.daci.accumulator[15] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0305_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold7 (.A(\stop.syn.daci.accumulator[10] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0166_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold9 (.A(\stop.syn.daci.accumulator[14] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold10 (.A(\stop.syn.daci.accumulator[12] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold11 (.A(\stop.syn.daci.accumulator[8] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0164_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold13 (.A(\stop.syn.daci.accumulator[13] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0298_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold15 (.A(\stop.syn.daci.accumulator[5] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0161_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold17 (.A(\stop.syn.daci.accumulator[6] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold18 (.A(\stop.syn.daci.accumulator[2] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0718_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0158_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold21 (.A(\stop.syn.daci.accumulator[11] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold22 (.A(\stop.syn.daci.accumulator[3] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0240_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0160_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold25 (.A(\stop.syn.daci.accumulator[9] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold26 (.A(\stop.syn.daci.accumulator[7] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold27 (.A(\stop.syn.daci.accumulator[2] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold28 (.A(\stop.syn.rstn_fst_reg2 ),
    .X(net134));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_4 FILLER_0_168 ();
 sg13g2_fill_2 FILLER_0_172 ();
 sg13g2_fill_2 FILLER_0_210 ();
 sg13g2_fill_1 FILLER_0_212 ();
 sg13g2_decap_8 FILLER_0_223 ();
 sg13g2_decap_8 FILLER_0_230 ();
 sg13g2_decap_4 FILLER_0_237 ();
 sg13g2_fill_2 FILLER_0_241 ();
 sg13g2_decap_8 FILLER_0_269 ();
 sg13g2_fill_2 FILLER_0_276 ();
 sg13g2_fill_2 FILLER_0_304 ();
 sg13g2_fill_1 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_4 FILLER_1_35 ();
 sg13g2_decap_4 FILLER_1_43 ();
 sg13g2_fill_2 FILLER_1_47 ();
 sg13g2_decap_8 FILLER_1_59 ();
 sg13g2_decap_8 FILLER_1_66 ();
 sg13g2_decap_8 FILLER_1_73 ();
 sg13g2_decap_8 FILLER_1_80 ();
 sg13g2_decap_8 FILLER_1_87 ();
 sg13g2_decap_8 FILLER_1_94 ();
 sg13g2_decap_8 FILLER_1_101 ();
 sg13g2_decap_8 FILLER_1_108 ();
 sg13g2_decap_8 FILLER_1_115 ();
 sg13g2_decap_8 FILLER_1_122 ();
 sg13g2_decap_8 FILLER_1_129 ();
 sg13g2_decap_8 FILLER_1_136 ();
 sg13g2_decap_8 FILLER_1_143 ();
 sg13g2_decap_8 FILLER_1_150 ();
 sg13g2_decap_8 FILLER_1_157 ();
 sg13g2_decap_8 FILLER_1_164 ();
 sg13g2_decap_8 FILLER_1_171 ();
 sg13g2_decap_8 FILLER_1_178 ();
 sg13g2_fill_2 FILLER_1_185 ();
 sg13g2_fill_1 FILLER_1_187 ();
 sg13g2_decap_8 FILLER_1_263 ();
 sg13g2_fill_2 FILLER_1_270 ();
 sg13g2_fill_1 FILLER_1_272 ();
 sg13g2_decap_8 FILLER_1_283 ();
 sg13g2_fill_1 FILLER_1_290 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_324 ();
 sg13g2_decap_8 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_338 ();
 sg13g2_decap_8 FILLER_1_345 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_21 ();
 sg13g2_fill_2 FILLER_2_54 ();
 sg13g2_fill_1 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_83 ();
 sg13g2_decap_8 FILLER_2_90 ();
 sg13g2_decap_8 FILLER_2_97 ();
 sg13g2_decap_8 FILLER_2_114 ();
 sg13g2_decap_8 FILLER_2_121 ();
 sg13g2_decap_8 FILLER_2_128 ();
 sg13g2_decap_8 FILLER_2_135 ();
 sg13g2_decap_8 FILLER_2_142 ();
 sg13g2_decap_8 FILLER_2_149 ();
 sg13g2_decap_8 FILLER_2_156 ();
 sg13g2_decap_8 FILLER_2_163 ();
 sg13g2_decap_8 FILLER_2_170 ();
 sg13g2_decap_8 FILLER_2_177 ();
 sg13g2_decap_4 FILLER_2_184 ();
 sg13g2_fill_1 FILLER_2_198 ();
 sg13g2_decap_8 FILLER_2_213 ();
 sg13g2_decap_4 FILLER_2_220 ();
 sg13g2_fill_1 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_fill_2 FILLER_2_235 ();
 sg13g2_fill_1 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_fill_1 FILLER_2_294 ();
 sg13g2_decap_4 FILLER_2_301 ();
 sg13g2_fill_1 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_4 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_16 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_4 FILLER_3_60 ();
 sg13g2_fill_2 FILLER_3_64 ();
 sg13g2_decap_8 FILLER_3_80 ();
 sg13g2_decap_4 FILLER_3_87 ();
 sg13g2_fill_2 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_157 ();
 sg13g2_decap_8 FILLER_3_164 ();
 sg13g2_fill_2 FILLER_3_171 ();
 sg13g2_fill_1 FILLER_3_173 ();
 sg13g2_fill_2 FILLER_3_205 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_fill_2 FILLER_3_326 ();
 sg13g2_fill_1 FILLER_3_340 ();
 sg13g2_fill_2 FILLER_3_351 ();
 sg13g2_decap_4 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_4_26 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_fill_2 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_4 FILLER_4_196 ();
 sg13g2_fill_2 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_216 ();
 sg13g2_fill_2 FILLER_4_223 ();
 sg13g2_fill_2 FILLER_4_236 ();
 sg13g2_decap_4 FILLER_4_242 ();
 sg13g2_fill_2 FILLER_4_246 ();
 sg13g2_decap_8 FILLER_4_292 ();
 sg13g2_fill_1 FILLER_4_345 ();
 sg13g2_decap_4 FILLER_4_365 ();
 sg13g2_fill_1 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_fill_2 FILLER_4_380 ();
 sg13g2_fill_1 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_9 ();
 sg13g2_decap_8 FILLER_5_40 ();
 sg13g2_decap_8 FILLER_5_47 ();
 sg13g2_fill_2 FILLER_5_54 ();
 sg13g2_fill_1 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_4 FILLER_5_74 ();
 sg13g2_fill_2 FILLER_5_78 ();
 sg13g2_fill_2 FILLER_5_84 ();
 sg13g2_fill_1 FILLER_5_86 ();
 sg13g2_decap_8 FILLER_5_97 ();
 sg13g2_fill_1 FILLER_5_104 ();
 sg13g2_decap_8 FILLER_5_115 ();
 sg13g2_decap_4 FILLER_5_122 ();
 sg13g2_decap_8 FILLER_5_146 ();
 sg13g2_decap_4 FILLER_5_153 ();
 sg13g2_fill_1 FILLER_5_157 ();
 sg13g2_fill_2 FILLER_5_184 ();
 sg13g2_fill_1 FILLER_5_212 ();
 sg13g2_decap_4 FILLER_5_239 ();
 sg13g2_decap_4 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_261 ();
 sg13g2_decap_8 FILLER_5_268 ();
 sg13g2_decap_8 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_282 ();
 sg13g2_fill_1 FILLER_5_289 ();
 sg13g2_fill_2 FILLER_5_304 ();
 sg13g2_fill_2 FILLER_5_314 ();
 sg13g2_fill_2 FILLER_5_321 ();
 sg13g2_decap_4 FILLER_5_331 ();
 sg13g2_fill_1 FILLER_5_335 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_fill_2 FILLER_5_346 ();
 sg13g2_decap_4 FILLER_5_363 ();
 sg13g2_fill_2 FILLER_5_367 ();
 sg13g2_fill_2 FILLER_5_381 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_27 ();
 sg13g2_fill_1 FILLER_6_31 ();
 sg13g2_decap_4 FILLER_6_136 ();
 sg13g2_decap_4 FILLER_6_186 ();
 sg13g2_fill_2 FILLER_6_190 ();
 sg13g2_decap_8 FILLER_6_197 ();
 sg13g2_decap_4 FILLER_6_204 ();
 sg13g2_decap_8 FILLER_6_218 ();
 sg13g2_decap_8 FILLER_6_225 ();
 sg13g2_decap_4 FILLER_6_232 ();
 sg13g2_fill_1 FILLER_6_236 ();
 sg13g2_fill_1 FILLER_6_241 ();
 sg13g2_decap_8 FILLER_6_247 ();
 sg13g2_decap_8 FILLER_6_254 ();
 sg13g2_fill_1 FILLER_6_261 ();
 sg13g2_fill_2 FILLER_6_270 ();
 sg13g2_fill_2 FILLER_6_306 ();
 sg13g2_fill_1 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_fill_2 FILLER_7_36 ();
 sg13g2_fill_1 FILLER_7_38 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_fill_2 FILLER_7_70 ();
 sg13g2_fill_1 FILLER_7_72 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_110 ();
 sg13g2_decap_4 FILLER_7_117 ();
 sg13g2_decap_8 FILLER_7_125 ();
 sg13g2_decap_8 FILLER_7_132 ();
 sg13g2_fill_1 FILLER_7_139 ();
 sg13g2_fill_1 FILLER_7_144 ();
 sg13g2_decap_8 FILLER_7_165 ();
 sg13g2_decap_8 FILLER_7_172 ();
 sg13g2_fill_2 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_181 ();
 sg13g2_decap_8 FILLER_7_208 ();
 sg13g2_decap_8 FILLER_7_215 ();
 sg13g2_decap_4 FILLER_7_222 ();
 sg13g2_fill_1 FILLER_7_226 ();
 sg13g2_decap_8 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_4 FILLER_7_326 ();
 sg13g2_decap_4 FILLER_7_340 ();
 sg13g2_fill_1 FILLER_7_344 ();
 sg13g2_fill_2 FILLER_7_363 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_fill_2 FILLER_7_380 ();
 sg13g2_fill_1 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_21 ();
 sg13g2_fill_2 FILLER_8_74 ();
 sg13g2_fill_1 FILLER_8_76 ();
 sg13g2_decap_8 FILLER_8_103 ();
 sg13g2_fill_1 FILLER_8_128 ();
 sg13g2_decap_8 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_198 ();
 sg13g2_fill_1 FILLER_8_245 ();
 sg13g2_fill_2 FILLER_8_256 ();
 sg13g2_fill_2 FILLER_8_284 ();
 sg13g2_decap_4 FILLER_8_298 ();
 sg13g2_decap_4 FILLER_8_324 ();
 sg13g2_fill_2 FILLER_8_328 ();
 sg13g2_fill_2 FILLER_8_356 ();
 sg13g2_fill_1 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_28 ();
 sg13g2_decap_4 FILLER_9_47 ();
 sg13g2_fill_2 FILLER_9_51 ();
 sg13g2_fill_1 FILLER_9_65 ();
 sg13g2_decap_4 FILLER_9_76 ();
 sg13g2_fill_1 FILLER_9_80 ();
 sg13g2_decap_4 FILLER_9_93 ();
 sg13g2_fill_1 FILLER_9_100 ();
 sg13g2_decap_4 FILLER_9_109 ();
 sg13g2_fill_1 FILLER_9_113 ();
 sg13g2_decap_4 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_172 ();
 sg13g2_decap_8 FILLER_9_179 ();
 sg13g2_fill_1 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_201 ();
 sg13g2_fill_2 FILLER_9_208 ();
 sg13g2_fill_1 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_215 ();
 sg13g2_fill_2 FILLER_9_222 ();
 sg13g2_fill_2 FILLER_9_237 ();
 sg13g2_fill_1 FILLER_9_260 ();
 sg13g2_decap_4 FILLER_9_265 ();
 sg13g2_decap_4 FILLER_9_273 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_fill_1 FILLER_9_286 ();
 sg13g2_decap_4 FILLER_9_291 ();
 sg13g2_fill_2 FILLER_9_295 ();
 sg13g2_decap_8 FILLER_9_325 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_4 FILLER_9_345 ();
 sg13g2_fill_2 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_fill_2 FILLER_10_66 ();
 sg13g2_decap_8 FILLER_10_72 ();
 sg13g2_fill_2 FILLER_10_79 ();
 sg13g2_decap_4 FILLER_10_96 ();
 sg13g2_fill_2 FILLER_10_100 ();
 sg13g2_fill_1 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_118 ();
 sg13g2_decap_4 FILLER_10_129 ();
 sg13g2_fill_1 FILLER_10_133 ();
 sg13g2_fill_2 FILLER_10_139 ();
 sg13g2_decap_4 FILLER_10_151 ();
 sg13g2_fill_2 FILLER_10_155 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_168 ();
 sg13g2_decap_4 FILLER_10_221 ();
 sg13g2_fill_2 FILLER_10_236 ();
 sg13g2_fill_2 FILLER_10_255 ();
 sg13g2_fill_1 FILLER_10_257 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_293 ();
 sg13g2_decap_4 FILLER_10_300 ();
 sg13g2_fill_1 FILLER_10_317 ();
 sg13g2_fill_1 FILLER_10_334 ();
 sg13g2_decap_4 FILLER_10_348 ();
 sg13g2_decap_4 FILLER_10_368 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_4 ();
 sg13g2_decap_4 FILLER_11_31 ();
 sg13g2_decap_8 FILLER_11_45 ();
 sg13g2_decap_4 FILLER_11_52 ();
 sg13g2_fill_2 FILLER_11_56 ();
 sg13g2_decap_4 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_114 ();
 sg13g2_fill_1 FILLER_11_116 ();
 sg13g2_fill_2 FILLER_11_143 ();
 sg13g2_fill_1 FILLER_11_145 ();
 sg13g2_decap_4 FILLER_11_172 ();
 sg13g2_fill_2 FILLER_11_200 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_fill_1 FILLER_11_233 ();
 sg13g2_fill_1 FILLER_11_239 ();
 sg13g2_decap_4 FILLER_11_248 ();
 sg13g2_fill_2 FILLER_11_252 ();
 sg13g2_decap_4 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_307 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_4 FILLER_11_329 ();
 sg13g2_fill_2 FILLER_11_333 ();
 sg13g2_fill_2 FILLER_11_343 ();
 sg13g2_decap_4 FILLER_11_353 ();
 sg13g2_fill_1 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_2 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_82 ();
 sg13g2_decap_8 FILLER_12_89 ();
 sg13g2_fill_1 FILLER_12_96 ();
 sg13g2_decap_8 FILLER_12_106 ();
 sg13g2_fill_1 FILLER_12_113 ();
 sg13g2_decap_4 FILLER_12_118 ();
 sg13g2_fill_2 FILLER_12_122 ();
 sg13g2_fill_2 FILLER_12_136 ();
 sg13g2_fill_2 FILLER_12_150 ();
 sg13g2_decap_8 FILLER_12_156 ();
 sg13g2_fill_1 FILLER_12_163 ();
 sg13g2_decap_8 FILLER_12_230 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_decap_4 FILLER_12_243 ();
 sg13g2_fill_1 FILLER_12_247 ();
 sg13g2_fill_1 FILLER_12_253 ();
 sg13g2_decap_8 FILLER_12_265 ();
 sg13g2_decap_4 FILLER_12_272 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_decap_8 FILLER_12_281 ();
 sg13g2_fill_2 FILLER_12_288 ();
 sg13g2_fill_1 FILLER_12_290 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_fill_2 FILLER_12_319 ();
 sg13g2_fill_2 FILLER_12_329 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_4 FILLER_12_349 ();
 sg13g2_fill_2 FILLER_12_353 ();
 sg13g2_decap_4 FILLER_12_373 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_38 ();
 sg13g2_fill_2 FILLER_13_45 ();
 sg13g2_fill_1 FILLER_13_52 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_188 ();
 sg13g2_decap_8 FILLER_13_195 ();
 sg13g2_fill_2 FILLER_13_202 ();
 sg13g2_fill_1 FILLER_13_204 ();
 sg13g2_decap_4 FILLER_13_210 ();
 sg13g2_fill_2 FILLER_13_214 ();
 sg13g2_fill_1 FILLER_13_242 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_decap_8 FILLER_13_310 ();
 sg13g2_fill_1 FILLER_13_317 ();
 sg13g2_fill_1 FILLER_13_359 ();
 sg13g2_fill_2 FILLER_13_376 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_4 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_4 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_87 ();
 sg13g2_fill_2 FILLER_14_97 ();
 sg13g2_fill_1 FILLER_14_99 ();
 sg13g2_decap_4 FILLER_14_136 ();
 sg13g2_decap_8 FILLER_14_146 ();
 sg13g2_decap_8 FILLER_14_153 ();
 sg13g2_decap_8 FILLER_14_160 ();
 sg13g2_decap_8 FILLER_14_167 ();
 sg13g2_decap_4 FILLER_14_174 ();
 sg13g2_fill_1 FILLER_14_178 ();
 sg13g2_decap_4 FILLER_14_205 ();
 sg13g2_fill_2 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_220 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_265 ();
 sg13g2_decap_8 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_278 ();
 sg13g2_decap_4 FILLER_14_284 ();
 sg13g2_decap_4 FILLER_14_321 ();
 sg13g2_fill_1 FILLER_14_337 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_fill_2 FILLER_14_350 ();
 sg13g2_fill_2 FILLER_14_365 ();
 sg13g2_fill_1 FILLER_14_367 ();
 sg13g2_fill_1 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_decap_4 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_48 ();
 sg13g2_decap_8 FILLER_15_55 ();
 sg13g2_fill_2 FILLER_15_62 ();
 sg13g2_fill_2 FILLER_15_74 ();
 sg13g2_fill_1 FILLER_15_76 ();
 sg13g2_fill_1 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_fill_2 FILLER_15_193 ();
 sg13g2_fill_1 FILLER_15_195 ();
 sg13g2_fill_1 FILLER_15_248 ();
 sg13g2_fill_2 FILLER_15_314 ();
 sg13g2_fill_2 FILLER_15_320 ();
 sg13g2_fill_1 FILLER_15_322 ();
 sg13g2_fill_2 FILLER_15_328 ();
 sg13g2_fill_1 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_9 ();
 sg13g2_decap_4 FILLER_16_16 ();
 sg13g2_fill_1 FILLER_16_20 ();
 sg13g2_fill_1 FILLER_16_29 ();
 sg13g2_fill_2 FILLER_16_54 ();
 sg13g2_fill_1 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_61 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_93 ();
 sg13g2_fill_2 FILLER_16_100 ();
 sg13g2_fill_1 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_fill_2 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_fill_2 FILLER_16_170 ();
 sg13g2_decap_8 FILLER_16_177 ();
 sg13g2_fill_2 FILLER_16_184 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_decap_8 FILLER_16_233 ();
 sg13g2_fill_1 FILLER_16_240 ();
 sg13g2_decap_4 FILLER_16_254 ();
 sg13g2_fill_2 FILLER_16_258 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_decap_4 FILLER_16_365 ();
 sg13g2_fill_1 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_4 FILLER_16_387 ();
 sg13g2_fill_1 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_1 FILLER_17_26 ();
 sg13g2_fill_1 FILLER_17_45 ();
 sg13g2_fill_2 FILLER_17_72 ();
 sg13g2_fill_1 FILLER_17_81 ();
 sg13g2_decap_4 FILLER_17_87 ();
 sg13g2_fill_1 FILLER_17_120 ();
 sg13g2_decap_8 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_137 ();
 sg13g2_fill_1 FILLER_17_139 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_fill_2 FILLER_17_275 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_294 ();
 sg13g2_decap_4 FILLER_17_304 ();
 sg13g2_fill_2 FILLER_17_347 ();
 sg13g2_fill_1 FILLER_17_349 ();
 sg13g2_decap_4 FILLER_17_376 ();
 sg13g2_fill_1 FILLER_17_380 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_15 ();
 sg13g2_fill_1 FILLER_18_31 ();
 sg13g2_decap_8 FILLER_18_41 ();
 sg13g2_decap_8 FILLER_18_48 ();
 sg13g2_decap_8 FILLER_18_55 ();
 sg13g2_fill_1 FILLER_18_62 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_decap_4 FILLER_18_91 ();
 sg13g2_fill_2 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_fill_1 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_157 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_decap_8 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_184 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_226 ();
 sg13g2_decap_4 FILLER_18_233 ();
 sg13g2_fill_2 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_247 ();
 sg13g2_fill_2 FILLER_18_254 ();
 sg13g2_fill_1 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_fill_1 FILLER_18_360 ();
 sg13g2_decap_4 FILLER_18_365 ();
 sg13g2_fill_1 FILLER_18_373 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_17 ();
 sg13g2_fill_1 FILLER_19_39 ();
 sg13g2_decap_4 FILLER_19_66 ();
 sg13g2_fill_1 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_88 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_116 ();
 sg13g2_decap_4 FILLER_19_123 ();
 sg13g2_fill_1 FILLER_19_127 ();
 sg13g2_fill_2 FILLER_19_166 ();
 sg13g2_decap_8 FILLER_19_194 ();
 sg13g2_decap_8 FILLER_19_227 ();
 sg13g2_decap_4 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_4 FILLER_19_284 ();
 sg13g2_fill_2 FILLER_19_295 ();
 sg13g2_decap_4 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_332 ();
 sg13g2_fill_2 FILLER_19_359 ();
 sg13g2_fill_1 FILLER_19_365 ();
 sg13g2_fill_2 FILLER_19_371 ();
 sg13g2_fill_1 FILLER_19_373 ();
 sg13g2_fill_1 FILLER_19_397 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_27 ();
 sg13g2_fill_2 FILLER_20_31 ();
 sg13g2_fill_1 FILLER_20_33 ();
 sg13g2_decap_8 FILLER_20_38 ();
 sg13g2_decap_4 FILLER_20_45 ();
 sg13g2_fill_2 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_55 ();
 sg13g2_fill_1 FILLER_20_62 ();
 sg13g2_fill_2 FILLER_20_84 ();
 sg13g2_fill_1 FILLER_20_86 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_decap_4 FILLER_20_152 ();
 sg13g2_fill_2 FILLER_20_156 ();
 sg13g2_fill_2 FILLER_20_170 ();
 sg13g2_decap_8 FILLER_20_180 ();
 sg13g2_decap_8 FILLER_20_187 ();
 sg13g2_decap_8 FILLER_20_199 ();
 sg13g2_decap_4 FILLER_20_206 ();
 sg13g2_decap_8 FILLER_20_213 ();
 sg13g2_decap_8 FILLER_20_220 ();
 sg13g2_decap_4 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_294 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_decap_4 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_17 ();
 sg13g2_fill_1 FILLER_21_24 ();
 sg13g2_fill_1 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_62 ();
 sg13g2_decap_4 FILLER_21_69 ();
 sg13g2_fill_2 FILLER_21_73 ();
 sg13g2_fill_2 FILLER_21_80 ();
 sg13g2_fill_2 FILLER_21_95 ();
 sg13g2_fill_1 FILLER_21_97 ();
 sg13g2_decap_4 FILLER_21_124 ();
 sg13g2_fill_2 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_decap_4 FILLER_21_176 ();
 sg13g2_fill_2 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_226 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_decap_8 FILLER_21_253 ();
 sg13g2_decap_8 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_278 ();
 sg13g2_decap_8 FILLER_21_285 ();
 sg13g2_fill_2 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_307 ();
 sg13g2_fill_1 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_4 FILLER_21_343 ();
 sg13g2_fill_2 FILLER_21_360 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_fill_1 FILLER_21_386 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_27 ();
 sg13g2_fill_1 FILLER_22_29 ();
 sg13g2_decap_4 FILLER_22_66 ();
 sg13g2_fill_1 FILLER_22_70 ();
 sg13g2_decap_4 FILLER_22_86 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_decap_8 FILLER_22_101 ();
 sg13g2_decap_4 FILLER_22_108 ();
 sg13g2_decap_4 FILLER_22_121 ();
 sg13g2_fill_1 FILLER_22_125 ();
 sg13g2_decap_4 FILLER_22_130 ();
 sg13g2_fill_2 FILLER_22_134 ();
 sg13g2_decap_8 FILLER_22_145 ();
 sg13g2_fill_2 FILLER_22_152 ();
 sg13g2_decap_4 FILLER_22_206 ();
 sg13g2_fill_2 FILLER_22_210 ();
 sg13g2_decap_4 FILLER_22_232 ();
 sg13g2_fill_1 FILLER_22_236 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_2 FILLER_22_295 ();
 sg13g2_fill_1 FILLER_22_302 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_fill_2 FILLER_22_347 ();
 sg13g2_fill_1 FILLER_22_358 ();
 sg13g2_fill_2 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_4 FILLER_23_30 ();
 sg13g2_fill_1 FILLER_23_34 ();
 sg13g2_fill_2 FILLER_23_87 ();
 sg13g2_fill_1 FILLER_23_89 ();
 sg13g2_decap_8 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_decap_8 FILLER_23_177 ();
 sg13g2_decap_8 FILLER_23_184 ();
 sg13g2_decap_8 FILLER_23_191 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_fill_1 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_264 ();
 sg13g2_decap_8 FILLER_23_274 ();
 sg13g2_decap_8 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_352 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_24 ();
 sg13g2_fill_1 FILLER_24_26 ();
 sg13g2_decap_8 FILLER_24_37 ();
 sg13g2_decap_8 FILLER_24_44 ();
 sg13g2_decap_8 FILLER_24_51 ();
 sg13g2_decap_4 FILLER_24_58 ();
 sg13g2_decap_8 FILLER_24_106 ();
 sg13g2_decap_8 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_120 ();
 sg13g2_decap_4 FILLER_24_131 ();
 sg13g2_decap_4 FILLER_24_143 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_210 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_236 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_decap_8 FILLER_24_276 ();
 sg13g2_decap_4 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_287 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_fill_2 FILLER_24_344 ();
 sg13g2_fill_1 FILLER_24_346 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_fill_1 FILLER_24_387 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_31 ();
 sg13g2_decap_4 FILLER_25_84 ();
 sg13g2_fill_2 FILLER_25_88 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_decap_4 FILLER_25_192 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_2 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_241 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_fill_2 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_fill_2 FILLER_25_368 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_fill_1 FILLER_26_17 ();
 sg13g2_fill_2 FILLER_26_33 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_decap_4 FILLER_26_72 ();
 sg13g2_decap_4 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_93 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_decap_8 FILLER_26_106 ();
 sg13g2_decap_4 FILLER_26_113 ();
 sg13g2_decap_8 FILLER_26_121 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_decap_8 FILLER_26_162 ();
 sg13g2_decap_8 FILLER_26_169 ();
 sg13g2_fill_2 FILLER_26_176 ();
 sg13g2_decap_4 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_decap_4 FILLER_26_207 ();
 sg13g2_fill_1 FILLER_26_211 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_fill_2 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_308 ();
 sg13g2_fill_2 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_368 ();
 sg13g2_fill_2 FILLER_26_391 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_27_26 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_44 ();
 sg13g2_fill_1 FILLER_27_58 ();
 sg13g2_decap_8 FILLER_27_132 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_fill_1 FILLER_27_141 ();
 sg13g2_decap_8 FILLER_27_163 ();
 sg13g2_decap_4 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_229 ();
 sg13g2_fill_2 FILLER_27_235 ();
 sg13g2_decap_4 FILLER_27_242 ();
 sg13g2_fill_1 FILLER_27_246 ();
 sg13g2_decap_8 FILLER_27_276 ();
 sg13g2_decap_8 FILLER_27_283 ();
 sg13g2_decap_4 FILLER_27_318 ();
 sg13g2_decap_8 FILLER_27_325 ();
 sg13g2_decap_8 FILLER_27_332 ();
 sg13g2_fill_1 FILLER_27_339 ();
 sg13g2_fill_2 FILLER_27_353 ();
 sg13g2_fill_2 FILLER_27_378 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_15 ();
 sg13g2_decap_8 FILLER_28_47 ();
 sg13g2_fill_2 FILLER_28_54 ();
 sg13g2_fill_1 FILLER_28_61 ();
 sg13g2_decap_4 FILLER_28_73 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_109 ();
 sg13g2_decap_4 FILLER_28_116 ();
 sg13g2_fill_2 FILLER_28_132 ();
 sg13g2_fill_1 FILLER_28_139 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_163 ();
 sg13g2_decap_8 FILLER_28_190 ();
 sg13g2_decap_4 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_4 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_284 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_2 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_342 ();
 sg13g2_fill_2 FILLER_28_360 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_29 ();
 sg13g2_fill_1 FILLER_29_31 ();
 sg13g2_decap_8 FILLER_29_36 ();
 sg13g2_decap_4 FILLER_29_43 ();
 sg13g2_decap_4 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_4 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_88 ();
 sg13g2_fill_1 FILLER_29_120 ();
 sg13g2_fill_1 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_165 ();
 sg13g2_fill_1 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_decap_8 FILLER_29_205 ();
 sg13g2_fill_1 FILLER_29_212 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_decap_8 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_256 ();
 sg13g2_decap_8 FILLER_29_262 ();
 sg13g2_decap_4 FILLER_29_269 ();
 sg13g2_fill_1 FILLER_29_273 ();
 sg13g2_decap_4 FILLER_29_288 ();
 sg13g2_fill_2 FILLER_29_300 ();
 sg13g2_decap_8 FILLER_29_314 ();
 sg13g2_decap_8 FILLER_29_321 ();
 sg13g2_fill_2 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_357 ();
 sg13g2_fill_2 FILLER_29_368 ();
 sg13g2_decap_8 FILLER_30_26 ();
 sg13g2_fill_2 FILLER_30_33 ();
 sg13g2_fill_1 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_60 ();
 sg13g2_fill_2 FILLER_30_64 ();
 sg13g2_decap_8 FILLER_30_92 ();
 sg13g2_decap_4 FILLER_30_99 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_134 ();
 sg13g2_decap_4 FILLER_30_141 ();
 sg13g2_decap_8 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_187 ();
 sg13g2_decap_8 FILLER_30_191 ();
 sg13g2_decap_4 FILLER_30_198 ();
 sg13g2_fill_2 FILLER_30_202 ();
 sg13g2_decap_4 FILLER_30_258 ();
 sg13g2_decap_4 FILLER_30_270 ();
 sg13g2_decap_8 FILLER_30_289 ();
 sg13g2_decap_4 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_319 ();
 sg13g2_fill_2 FILLER_30_325 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_decap_8 FILLER_30_331 ();
 sg13g2_decap_8 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_12 ();
 sg13g2_fill_2 FILLER_31_18 ();
 sg13g2_fill_1 FILLER_31_20 ();
 sg13g2_decap_4 FILLER_31_47 ();
 sg13g2_fill_2 FILLER_31_51 ();
 sg13g2_fill_2 FILLER_31_79 ();
 sg13g2_decap_8 FILLER_31_86 ();
 sg13g2_fill_2 FILLER_31_93 ();
 sg13g2_fill_1 FILLER_31_95 ();
 sg13g2_decap_4 FILLER_31_116 ();
 sg13g2_fill_2 FILLER_31_120 ();
 sg13g2_fill_2 FILLER_31_125 ();
 sg13g2_fill_1 FILLER_31_127 ();
 sg13g2_decap_4 FILLER_31_162 ();
 sg13g2_fill_2 FILLER_31_169 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_decap_4 FILLER_31_231 ();
 sg13g2_decap_4 FILLER_31_261 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_fill_2 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_31_356 ();
 sg13g2_fill_1 FILLER_31_358 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_37 ();
 sg13g2_decap_8 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_72 ();
 sg13g2_fill_2 FILLER_32_97 ();
 sg13g2_fill_1 FILLER_32_99 ();
 sg13g2_decap_4 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_111 ();
 sg13g2_decap_4 FILLER_32_138 ();
 sg13g2_fill_2 FILLER_32_142 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_184 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_fill_1 FILLER_32_208 ();
 sg13g2_decap_4 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_309 ();
 sg13g2_fill_1 FILLER_32_311 ();
 sg13g2_decap_4 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_332 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_33_26 ();
 sg13g2_decap_8 FILLER_33_33 ();
 sg13g2_decap_8 FILLER_33_40 ();
 sg13g2_fill_2 FILLER_33_47 ();
 sg13g2_fill_1 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_54 ();
 sg13g2_decap_8 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_68 ();
 sg13g2_decap_4 FILLER_33_87 ();
 sg13g2_fill_2 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_122 ();
 sg13g2_fill_2 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_decap_8 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_172 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_decap_4 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_decap_8 FILLER_33_200 ();
 sg13g2_decap_4 FILLER_33_207 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_decap_4 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_272 ();
 sg13g2_decap_4 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_4 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_330 ();
 sg13g2_decap_8 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_12 ();
 sg13g2_fill_2 FILLER_34_16 ();
 sg13g2_decap_8 FILLER_34_47 ();
 sg13g2_decap_8 FILLER_34_54 ();
 sg13g2_fill_1 FILLER_34_61 ();
 sg13g2_decap_4 FILLER_34_85 ();
 sg13g2_fill_1 FILLER_34_89 ();
 sg13g2_decap_4 FILLER_34_102 ();
 sg13g2_decap_4 FILLER_34_132 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_decap_4 FILLER_34_151 ();
 sg13g2_fill_1 FILLER_34_172 ();
 sg13g2_decap_8 FILLER_34_215 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_34_316 ();
 sg13g2_fill_1 FILLER_34_318 ();
 sg13g2_decap_4 FILLER_34_345 ();
 sg13g2_fill_2 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_16 ();
 sg13g2_decap_8 FILLER_35_20 ();
 sg13g2_fill_2 FILLER_35_27 ();
 sg13g2_fill_1 FILLER_35_66 ();
 sg13g2_decap_8 FILLER_35_79 ();
 sg13g2_fill_1 FILLER_35_110 ();
 sg13g2_fill_2 FILLER_35_137 ();
 sg13g2_decap_4 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_decap_4 FILLER_35_257 ();
 sg13g2_fill_2 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_fill_1 FILLER_35_348 ();
 sg13g2_fill_2 FILLER_35_390 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_87 ();
 sg13g2_fill_1 FILLER_36_89 ();
 sg13g2_fill_1 FILLER_36_94 ();
 sg13g2_decap_8 FILLER_36_124 ();
 sg13g2_decap_8 FILLER_36_165 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_fill_2 FILLER_36_200 ();
 sg13g2_fill_2 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_254 ();
 sg13g2_decap_8 FILLER_36_289 ();
 sg13g2_fill_1 FILLER_36_296 ();
 sg13g2_decap_4 FILLER_36_312 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_346 ();
 sg13g2_fill_2 FILLER_36_370 ();
 sg13g2_fill_1 FILLER_36_372 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_4 FILLER_37_35 ();
 sg13g2_fill_2 FILLER_37_39 ();
 sg13g2_fill_2 FILLER_37_53 ();
 sg13g2_decap_8 FILLER_37_97 ();
 sg13g2_fill_1 FILLER_37_104 ();
 sg13g2_decap_4 FILLER_37_131 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_decap_4 FILLER_37_140 ();
 sg13g2_decap_4 FILLER_37_156 ();
 sg13g2_fill_1 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_fill_2 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_317 ();
 sg13g2_decap_4 FILLER_37_321 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_32 ();
 sg13g2_fill_2 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_62 ();
 sg13g2_fill_2 FILLER_38_93 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_2 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_110 ();
 sg13g2_fill_1 FILLER_38_116 ();
 sg13g2_fill_2 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_186 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_4 FILLER_38_207 ();
 sg13g2_fill_2 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_4 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_decap_4 FILLER_38_260 ();
 sg13g2_fill_1 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_269 ();
 sg13g2_decap_8 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_283 ();
 sg13g2_fill_1 FILLER_38_285 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_fill_1 FILLER_38_308 ();
 sg13g2_fill_2 FILLER_38_335 ();
 sg13g2_fill_1 FILLER_38_337 ();
 assign uio_oe[0] = net104;
 assign uio_oe[1] = net105;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[2] = net10;
 assign uio_out[3] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
 assign uio_out[7] = net15;
endmodule

module tt_um_dmtd_arghunter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire \u_dmtd.async_reg1[0] ;
 wire \u_dmtd.async_reg1[1] ;
 wire \u_dmtd.async_reg1[2] ;
 wire \u_dmtd.async_reg2[0] ;
 wire \u_dmtd.async_reg2[1] ;
 wire \u_dmtd.async_reg2[2] ;
 wire \u_dmtd.dmtd_out ;
 wire \u_dmtd.shift_reg[0] ;
 wire \u_dmtd.shift_reg[100] ;
 wire \u_dmtd.shift_reg[101] ;
 wire \u_dmtd.shift_reg[102] ;
 wire \u_dmtd.shift_reg[103] ;
 wire \u_dmtd.shift_reg[104] ;
 wire \u_dmtd.shift_reg[105] ;
 wire \u_dmtd.shift_reg[106] ;
 wire \u_dmtd.shift_reg[107] ;
 wire \u_dmtd.shift_reg[108] ;
 wire \u_dmtd.shift_reg[109] ;
 wire \u_dmtd.shift_reg[10] ;
 wire \u_dmtd.shift_reg[110] ;
 wire \u_dmtd.shift_reg[111] ;
 wire \u_dmtd.shift_reg[112] ;
 wire \u_dmtd.shift_reg[113] ;
 wire \u_dmtd.shift_reg[114] ;
 wire \u_dmtd.shift_reg[115] ;
 wire \u_dmtd.shift_reg[116] ;
 wire \u_dmtd.shift_reg[117] ;
 wire \u_dmtd.shift_reg[118] ;
 wire \u_dmtd.shift_reg[119] ;
 wire \u_dmtd.shift_reg[11] ;
 wire \u_dmtd.shift_reg[120] ;
 wire \u_dmtd.shift_reg[121] ;
 wire \u_dmtd.shift_reg[122] ;
 wire \u_dmtd.shift_reg[123] ;
 wire \u_dmtd.shift_reg[124] ;
 wire \u_dmtd.shift_reg[125] ;
 wire \u_dmtd.shift_reg[126] ;
 wire \u_dmtd.shift_reg[127] ;
 wire \u_dmtd.shift_reg[12] ;
 wire \u_dmtd.shift_reg[13] ;
 wire \u_dmtd.shift_reg[14] ;
 wire \u_dmtd.shift_reg[15] ;
 wire \u_dmtd.shift_reg[16] ;
 wire \u_dmtd.shift_reg[17] ;
 wire \u_dmtd.shift_reg[18] ;
 wire \u_dmtd.shift_reg[19] ;
 wire \u_dmtd.shift_reg[1] ;
 wire \u_dmtd.shift_reg[20] ;
 wire \u_dmtd.shift_reg[21] ;
 wire \u_dmtd.shift_reg[22] ;
 wire \u_dmtd.shift_reg[23] ;
 wire \u_dmtd.shift_reg[24] ;
 wire \u_dmtd.shift_reg[25] ;
 wire \u_dmtd.shift_reg[26] ;
 wire \u_dmtd.shift_reg[27] ;
 wire \u_dmtd.shift_reg[28] ;
 wire \u_dmtd.shift_reg[29] ;
 wire \u_dmtd.shift_reg[2] ;
 wire \u_dmtd.shift_reg[30] ;
 wire \u_dmtd.shift_reg[31] ;
 wire \u_dmtd.shift_reg[32] ;
 wire \u_dmtd.shift_reg[33] ;
 wire \u_dmtd.shift_reg[34] ;
 wire \u_dmtd.shift_reg[35] ;
 wire \u_dmtd.shift_reg[36] ;
 wire \u_dmtd.shift_reg[37] ;
 wire \u_dmtd.shift_reg[38] ;
 wire \u_dmtd.shift_reg[39] ;
 wire \u_dmtd.shift_reg[3] ;
 wire \u_dmtd.shift_reg[40] ;
 wire \u_dmtd.shift_reg[41] ;
 wire \u_dmtd.shift_reg[42] ;
 wire \u_dmtd.shift_reg[43] ;
 wire \u_dmtd.shift_reg[44] ;
 wire \u_dmtd.shift_reg[45] ;
 wire \u_dmtd.shift_reg[46] ;
 wire \u_dmtd.shift_reg[47] ;
 wire \u_dmtd.shift_reg[48] ;
 wire \u_dmtd.shift_reg[49] ;
 wire \u_dmtd.shift_reg[4] ;
 wire \u_dmtd.shift_reg[50] ;
 wire \u_dmtd.shift_reg[51] ;
 wire \u_dmtd.shift_reg[52] ;
 wire \u_dmtd.shift_reg[53] ;
 wire \u_dmtd.shift_reg[54] ;
 wire \u_dmtd.shift_reg[55] ;
 wire \u_dmtd.shift_reg[56] ;
 wire \u_dmtd.shift_reg[57] ;
 wire \u_dmtd.shift_reg[58] ;
 wire \u_dmtd.shift_reg[59] ;
 wire \u_dmtd.shift_reg[5] ;
 wire \u_dmtd.shift_reg[60] ;
 wire \u_dmtd.shift_reg[61] ;
 wire \u_dmtd.shift_reg[62] ;
 wire \u_dmtd.shift_reg[63] ;
 wire \u_dmtd.shift_reg[64] ;
 wire \u_dmtd.shift_reg[65] ;
 wire \u_dmtd.shift_reg[66] ;
 wire \u_dmtd.shift_reg[67] ;
 wire \u_dmtd.shift_reg[68] ;
 wire \u_dmtd.shift_reg[69] ;
 wire \u_dmtd.shift_reg[6] ;
 wire \u_dmtd.shift_reg[70] ;
 wire \u_dmtd.shift_reg[71] ;
 wire \u_dmtd.shift_reg[72] ;
 wire \u_dmtd.shift_reg[73] ;
 wire \u_dmtd.shift_reg[74] ;
 wire \u_dmtd.shift_reg[75] ;
 wire \u_dmtd.shift_reg[76] ;
 wire \u_dmtd.shift_reg[77] ;
 wire \u_dmtd.shift_reg[78] ;
 wire \u_dmtd.shift_reg[79] ;
 wire \u_dmtd.shift_reg[7] ;
 wire \u_dmtd.shift_reg[80] ;
 wire \u_dmtd.shift_reg[81] ;
 wire \u_dmtd.shift_reg[82] ;
 wire \u_dmtd.shift_reg[83] ;
 wire \u_dmtd.shift_reg[84] ;
 wire \u_dmtd.shift_reg[85] ;
 wire \u_dmtd.shift_reg[86] ;
 wire \u_dmtd.shift_reg[87] ;
 wire \u_dmtd.shift_reg[88] ;
 wire \u_dmtd.shift_reg[89] ;
 wire \u_dmtd.shift_reg[8] ;
 wire \u_dmtd.shift_reg[90] ;
 wire \u_dmtd.shift_reg[91] ;
 wire \u_dmtd.shift_reg[92] ;
 wire \u_dmtd.shift_reg[93] ;
 wire \u_dmtd.shift_reg[94] ;
 wire \u_dmtd.shift_reg[95] ;
 wire \u_dmtd.shift_reg[96] ;
 wire \u_dmtd.shift_reg[97] ;
 wire \u_dmtd.shift_reg[98] ;
 wire \u_dmtd.shift_reg[99] ;
 wire \u_dmtd.shift_reg[9] ;
 wire \u_dmtd.sync_out2 ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;

 sg13g2_inv_2 _282_ (.Y(_000_),
    .A(net4));
 sg13g2_inv_2 _283_ (.Y(_001_),
    .A(net5));
 sg13g2_inv_1 _284_ (.Y(_002_),
    .A(net6));
 sg13g2_nor2b_1 _285_ (.A(net3),
    .B_N(\u_dmtd.async_reg1[2] ),
    .Y(_003_));
 sg13g2_a21oi_2 _286_ (.B1(_003_),
    .Y(_004_),
    .A2(net3),
    .A1(\u_dmtd.async_reg2[2] ));
 sg13g2_nor2b_1 _287_ (.A(net234),
    .B_N(\u_dmtd.shift_reg[30] ),
    .Y(_005_));
 sg13g2_a21oi_1 _288_ (.A1(net234),
    .A2(\u_dmtd.shift_reg[31] ),
    .Y(_006_),
    .B1(_005_));
 sg13g2_mux2_1 _289_ (.A0(\u_dmtd.shift_reg[28] ),
    .A1(\u_dmtd.shift_reg[29] ),
    .S(net234),
    .X(_007_));
 sg13g2_o21ai_1 _290_ (.B1(net216),
    .Y(_008_),
    .A1(net224),
    .A2(_007_));
 sg13g2_a21oi_1 _291_ (.A1(net224),
    .A2(_006_),
    .Y(_009_),
    .B1(_008_));
 sg13g2_mux4_1 _292_ (.S0(net230),
    .A0(\u_dmtd.shift_reg[24] ),
    .A1(\u_dmtd.shift_reg[25] ),
    .A2(\u_dmtd.shift_reg[26] ),
    .A3(\u_dmtd.shift_reg[27] ),
    .S1(net224),
    .X(_010_));
 sg13g2_nor2b_1 _293_ (.A(net216),
    .B_N(_010_),
    .Y(_011_));
 sg13g2_o21ai_1 _294_ (.B1(net4),
    .Y(_012_),
    .A1(_009_),
    .A2(_011_));
 sg13g2_nor2b_1 _295_ (.A(net238),
    .B_N(\u_dmtd.shift_reg[22] ),
    .Y(_013_));
 sg13g2_a21oi_1 _296_ (.A1(net232),
    .A2(\u_dmtd.shift_reg[23] ),
    .Y(_014_),
    .B1(_013_));
 sg13g2_mux2_1 _297_ (.A0(\u_dmtd.shift_reg[20] ),
    .A1(\u_dmtd.shift_reg[21] ),
    .S(net232),
    .X(_015_));
 sg13g2_o21ai_1 _298_ (.B1(net215),
    .Y(_016_),
    .A1(net222),
    .A2(_015_));
 sg13g2_a21oi_1 _299_ (.A1(net222),
    .A2(_014_),
    .Y(_017_),
    .B1(_016_));
 sg13g2_mux4_1 _300_ (.S0(net232),
    .A0(\u_dmtd.shift_reg[16] ),
    .A1(\u_dmtd.shift_reg[17] ),
    .A2(\u_dmtd.shift_reg[18] ),
    .A3(\u_dmtd.shift_reg[19] ),
    .S1(net222),
    .X(_018_));
 sg13g2_nor2b_1 _301_ (.A(net215),
    .B_N(_018_),
    .Y(_019_));
 sg13g2_o21ai_1 _302_ (.B1(_000_),
    .Y(_020_),
    .A1(_017_),
    .A2(_019_));
 sg13g2_a21o_1 _303_ (.A2(_020_),
    .A1(_012_),
    .B1(_001_),
    .X(_021_));
 sg13g2_nand2b_1 _304_ (.Y(_022_),
    .B(\u_dmtd.shift_reg[6] ),
    .A_N(net236));
 sg13g2_nand2_1 _305_ (.Y(_023_),
    .A(net236),
    .B(\u_dmtd.shift_reg[7] ));
 sg13g2_and3_1 _306_ (.X(_024_),
    .A(net227),
    .B(_022_),
    .C(_023_));
 sg13g2_mux2_1 _307_ (.A0(\u_dmtd.shift_reg[4] ),
    .A1(\u_dmtd.shift_reg[5] ),
    .S(net235),
    .X(_025_));
 sg13g2_o21ai_1 _308_ (.B1(net217),
    .Y(_026_),
    .A1(net227),
    .A2(_025_));
 sg13g2_mux4_1 _309_ (.S0(net236),
    .A0(\u_dmtd.shift_reg[0] ),
    .A1(\u_dmtd.shift_reg[1] ),
    .A2(\u_dmtd.shift_reg[2] ),
    .A3(\u_dmtd.shift_reg[3] ),
    .S1(net227),
    .X(_027_));
 sg13g2_nand2b_1 _310_ (.Y(_028_),
    .B(_027_),
    .A_N(net217));
 sg13g2_o21ai_1 _311_ (.B1(_028_),
    .Y(_029_),
    .A1(_024_),
    .A2(_026_));
 sg13g2_mux4_1 _312_ (.S0(net235),
    .A0(\u_dmtd.shift_reg[8] ),
    .A1(\u_dmtd.shift_reg[9] ),
    .A2(\u_dmtd.shift_reg[10] ),
    .A3(\u_dmtd.shift_reg[11] ),
    .S1(net226),
    .X(_030_));
 sg13g2_nand2b_1 _313_ (.Y(_031_),
    .B(_030_),
    .A_N(net217));
 sg13g2_nand2b_1 _314_ (.Y(_032_),
    .B(\u_dmtd.shift_reg[14] ),
    .A_N(net235));
 sg13g2_nand2_1 _315_ (.Y(_033_),
    .A(net235),
    .B(\u_dmtd.shift_reg[15] ));
 sg13g2_and3_1 _316_ (.X(_034_),
    .A(net226),
    .B(_032_),
    .C(_033_));
 sg13g2_mux2_1 _317_ (.A0(\u_dmtd.shift_reg[12] ),
    .A1(\u_dmtd.shift_reg[13] ),
    .S(net235),
    .X(_035_));
 sg13g2_o21ai_1 _318_ (.B1(net217),
    .Y(_036_),
    .A1(net226),
    .A2(_035_));
 sg13g2_o21ai_1 _319_ (.B1(_031_),
    .Y(_037_),
    .A1(_034_),
    .A2(_036_));
 sg13g2_mux2_1 _320_ (.A0(_029_),
    .A1(_037_),
    .S(net4),
    .X(_038_));
 sg13g2_a21oi_1 _321_ (.A1(_001_),
    .A2(_038_),
    .Y(_039_),
    .B1(net6));
 sg13g2_nor2b_1 _322_ (.A(net230),
    .B_N(\u_dmtd.shift_reg[54] ),
    .Y(_040_));
 sg13g2_a21oi_1 _323_ (.A1(net230),
    .A2(\u_dmtd.shift_reg[55] ),
    .Y(_041_),
    .B1(_040_));
 sg13g2_mux2_1 _324_ (.A0(\u_dmtd.shift_reg[52] ),
    .A1(\u_dmtd.shift_reg[53] ),
    .S(net230),
    .X(_042_));
 sg13g2_o21ai_1 _325_ (.B1(net214),
    .Y(_043_),
    .A1(net220),
    .A2(_042_));
 sg13g2_a21oi_1 _326_ (.A1(net220),
    .A2(_041_),
    .Y(_044_),
    .B1(_043_));
 sg13g2_mux4_1 _327_ (.S0(net230),
    .A0(\u_dmtd.shift_reg[48] ),
    .A1(\u_dmtd.shift_reg[49] ),
    .A2(\u_dmtd.shift_reg[50] ),
    .A3(\u_dmtd.shift_reg[51] ),
    .S1(net220),
    .X(_045_));
 sg13g2_nor2b_1 _328_ (.A(net214),
    .B_N(_045_),
    .Y(_046_));
 sg13g2_nor3_1 _329_ (.A(net4),
    .B(_044_),
    .C(_046_),
    .Y(_047_));
 sg13g2_mux4_1 _330_ (.S0(net229),
    .A0(\u_dmtd.shift_reg[56] ),
    .A1(\u_dmtd.shift_reg[57] ),
    .A2(\u_dmtd.shift_reg[58] ),
    .A3(\u_dmtd.shift_reg[59] ),
    .S1(net220),
    .X(_048_));
 sg13g2_nor2b_1 _331_ (.A(net214),
    .B_N(_048_),
    .Y(_049_));
 sg13g2_nor2b_1 _332_ (.A(net228),
    .B_N(\u_dmtd.shift_reg[62] ),
    .Y(_050_));
 sg13g2_a21oi_1 _333_ (.A1(net228),
    .A2(\u_dmtd.shift_reg[63] ),
    .Y(_051_),
    .B1(_050_));
 sg13g2_mux2_1 _334_ (.A0(\u_dmtd.shift_reg[60] ),
    .A1(\u_dmtd.shift_reg[61] ),
    .S(net229),
    .X(_052_));
 sg13g2_o21ai_1 _335_ (.B1(net214),
    .Y(_053_),
    .A1(net219),
    .A2(_052_));
 sg13g2_a21oi_1 _336_ (.A1(net219),
    .A2(_051_),
    .Y(_054_),
    .B1(_053_));
 sg13g2_nor3_1 _337_ (.A(_000_),
    .B(_049_),
    .C(_054_),
    .Y(_055_));
 sg13g2_or3_1 _338_ (.A(_001_),
    .B(_047_),
    .C(_055_),
    .X(_056_));
 sg13g2_nand2b_1 _339_ (.Y(_057_),
    .B(\u_dmtd.shift_reg[46] ),
    .A_N(net234));
 sg13g2_nand2_1 _340_ (.Y(_058_),
    .A(net234),
    .B(\u_dmtd.shift_reg[47] ));
 sg13g2_and3_1 _341_ (.X(_059_),
    .A(net224),
    .B(_057_),
    .C(_058_));
 sg13g2_mux2_1 _342_ (.A0(\u_dmtd.shift_reg[44] ),
    .A1(\u_dmtd.shift_reg[45] ),
    .S(net234),
    .X(_060_));
 sg13g2_o21ai_1 _343_ (.B1(net216),
    .Y(_061_),
    .A1(net224),
    .A2(_060_));
 sg13g2_mux4_1 _344_ (.S0(net234),
    .A0(\u_dmtd.shift_reg[40] ),
    .A1(\u_dmtd.shift_reg[41] ),
    .A2(\u_dmtd.shift_reg[42] ),
    .A3(\u_dmtd.shift_reg[43] ),
    .S1(net224),
    .X(_062_));
 sg13g2_nand2b_1 _345_ (.Y(_063_),
    .B(_062_),
    .A_N(net216));
 sg13g2_o21ai_1 _346_ (.B1(_063_),
    .Y(_064_),
    .A1(_059_),
    .A2(_061_));
 sg13g2_nand2b_1 _347_ (.Y(_065_),
    .B(\u_dmtd.shift_reg[38] ),
    .A_N(net233));
 sg13g2_nand2_1 _348_ (.Y(_066_),
    .A(net233),
    .B(\u_dmtd.shift_reg[39] ));
 sg13g2_and3_1 _349_ (.X(_067_),
    .A(net225),
    .B(_065_),
    .C(_066_));
 sg13g2_mux2_1 _350_ (.A0(\u_dmtd.shift_reg[36] ),
    .A1(\u_dmtd.shift_reg[37] ),
    .S(net233),
    .X(_068_));
 sg13g2_o21ai_1 _351_ (.B1(net216),
    .Y(_069_),
    .A1(net225),
    .A2(_068_));
 sg13g2_mux4_1 _352_ (.S0(net233),
    .A0(\u_dmtd.shift_reg[32] ),
    .A1(\u_dmtd.shift_reg[33] ),
    .A2(\u_dmtd.shift_reg[34] ),
    .A3(\u_dmtd.shift_reg[35] ),
    .S1(net225),
    .X(_070_));
 sg13g2_nand2b_1 _353_ (.Y(_071_),
    .B(_070_),
    .A_N(net216));
 sg13g2_o21ai_1 _354_ (.B1(_071_),
    .Y(_072_),
    .A1(_067_),
    .A2(_069_));
 sg13g2_mux2_1 _355_ (.A0(_064_),
    .A1(_072_),
    .S(_000_),
    .X(_073_));
 sg13g2_a21oi_1 _356_ (.A1(_001_),
    .A2(_073_),
    .Y(_074_),
    .B1(_002_));
 sg13g2_nand2b_1 _357_ (.Y(_075_),
    .B(\u_dmtd.shift_reg[126] ),
    .A_N(net233));
 sg13g2_nand2_1 _358_ (.Y(_076_),
    .A(net233),
    .B(\u_dmtd.shift_reg[127] ));
 sg13g2_and3_1 _359_ (.X(_077_),
    .A(net225),
    .B(_075_),
    .C(_076_));
 sg13g2_mux2_1 _360_ (.A0(\u_dmtd.shift_reg[124] ),
    .A1(\u_dmtd.shift_reg[125] ),
    .S(net233),
    .X(_078_));
 sg13g2_o21ai_1 _361_ (.B1(net216),
    .Y(_079_),
    .A1(net225),
    .A2(_078_));
 sg13g2_mux4_1 _362_ (.S0(net237),
    .A0(\u_dmtd.shift_reg[120] ),
    .A1(\u_dmtd.shift_reg[121] ),
    .A2(\u_dmtd.shift_reg[122] ),
    .A3(\u_dmtd.shift_reg[123] ),
    .S1(net224),
    .X(_080_));
 sg13g2_nand2b_1 _363_ (.Y(_081_),
    .B(_080_),
    .A_N(net216));
 sg13g2_o21ai_1 _364_ (.B1(_081_),
    .Y(_082_),
    .A1(_077_),
    .A2(_079_));
 sg13g2_nand2b_1 _365_ (.Y(_083_),
    .B(\u_dmtd.shift_reg[118] ),
    .A_N(net237));
 sg13g2_nand2_1 _366_ (.Y(_084_),
    .A(net233),
    .B(\u_dmtd.shift_reg[119] ));
 sg13g2_and3_1 _367_ (.X(_085_),
    .A(net224),
    .B(_083_),
    .C(_084_));
 sg13g2_mux2_1 _368_ (.A0(\u_dmtd.shift_reg[116] ),
    .A1(\u_dmtd.shift_reg[117] ),
    .S(net236),
    .X(_086_));
 sg13g2_o21ai_1 _369_ (.B1(net217),
    .Y(_087_),
    .A1(net226),
    .A2(_086_));
 sg13g2_mux4_1 _370_ (.S0(net235),
    .A0(\u_dmtd.shift_reg[112] ),
    .A1(\u_dmtd.shift_reg[113] ),
    .A2(\u_dmtd.shift_reg[114] ),
    .A3(\u_dmtd.shift_reg[115] ),
    .S1(net226),
    .X(_088_));
 sg13g2_nand2b_1 _371_ (.Y(_089_),
    .B(_088_),
    .A_N(net217));
 sg13g2_o21ai_1 _372_ (.B1(_089_),
    .Y(_090_),
    .A1(_085_),
    .A2(_087_));
 sg13g2_mux2_1 _373_ (.A0(_082_),
    .A1(_090_),
    .S(_000_),
    .X(_091_));
 sg13g2_nor2b_1 _374_ (.A(net232),
    .B_N(\u_dmtd.shift_reg[102] ),
    .Y(_092_));
 sg13g2_a21oi_1 _375_ (.A1(net232),
    .A2(\u_dmtd.shift_reg[103] ),
    .Y(_093_),
    .B1(_092_));
 sg13g2_mux2_1 _376_ (.A0(\u_dmtd.shift_reg[100] ),
    .A1(\u_dmtd.shift_reg[101] ),
    .S(net231),
    .X(_094_));
 sg13g2_o21ai_1 _377_ (.B1(net215),
    .Y(_095_),
    .A1(net221),
    .A2(_094_));
 sg13g2_a21oi_1 _378_ (.A1(net222),
    .A2(_093_),
    .Y(_096_),
    .B1(_095_));
 sg13g2_mux4_1 _379_ (.S0(net232),
    .A0(\u_dmtd.shift_reg[96] ),
    .A1(\u_dmtd.shift_reg[97] ),
    .A2(\u_dmtd.shift_reg[98] ),
    .A3(\u_dmtd.shift_reg[99] ),
    .S1(net221),
    .X(_097_));
 sg13g2_nor2b_1 _380_ (.A(net215),
    .B_N(_097_),
    .Y(_098_));
 sg13g2_nor3_1 _381_ (.A(net4),
    .B(_096_),
    .C(_098_),
    .Y(_099_));
 sg13g2_mux4_1 _382_ (.S0(net235),
    .A0(\u_dmtd.shift_reg[104] ),
    .A1(\u_dmtd.shift_reg[105] ),
    .A2(\u_dmtd.shift_reg[106] ),
    .A3(\u_dmtd.shift_reg[107] ),
    .S1(net226),
    .X(_100_));
 sg13g2_nor2b_1 _383_ (.A(net217),
    .B_N(_100_),
    .Y(_101_));
 sg13g2_nor2b_1 _384_ (.A(net236),
    .B_N(\u_dmtd.shift_reg[110] ),
    .Y(_102_));
 sg13g2_a21oi_1 _385_ (.A1(net236),
    .A2(\u_dmtd.shift_reg[111] ),
    .Y(_103_),
    .B1(_102_));
 sg13g2_mux2_1 _386_ (.A0(\u_dmtd.shift_reg[108] ),
    .A1(\u_dmtd.shift_reg[109] ),
    .S(net235),
    .X(_104_));
 sg13g2_o21ai_1 _387_ (.B1(net217),
    .Y(_105_),
    .A1(net226),
    .A2(_104_));
 sg13g2_a21oi_1 _388_ (.A1(net226),
    .A2(_103_),
    .Y(_106_),
    .B1(_105_));
 sg13g2_nor3_1 _389_ (.A(_000_),
    .B(_101_),
    .C(_106_),
    .Y(_107_));
 sg13g2_or3_1 _390_ (.A(net5),
    .B(_099_),
    .C(_107_),
    .X(_108_));
 sg13g2_a21oi_1 _391_ (.A1(net5),
    .A2(_091_),
    .Y(_109_),
    .B1(_002_));
 sg13g2_nor2b_1 _392_ (.A(net231),
    .B_N(\u_dmtd.shift_reg[94] ),
    .Y(_110_));
 sg13g2_a21oi_1 _393_ (.A1(net231),
    .A2(\u_dmtd.shift_reg[95] ),
    .Y(_111_),
    .B1(_110_));
 sg13g2_mux2_1 _394_ (.A0(\u_dmtd.shift_reg[92] ),
    .A1(\u_dmtd.shift_reg[93] ),
    .S(net231),
    .X(_112_));
 sg13g2_o21ai_1 _395_ (.B1(net215),
    .Y(_113_),
    .A1(net221),
    .A2(_112_));
 sg13g2_a21oi_1 _396_ (.A1(net221),
    .A2(_111_),
    .Y(_114_),
    .B1(_113_));
 sg13g2_mux4_1 _397_ (.S0(net232),
    .A0(\u_dmtd.shift_reg[88] ),
    .A1(\u_dmtd.shift_reg[89] ),
    .A2(\u_dmtd.shift_reg[90] ),
    .A3(\u_dmtd.shift_reg[91] ),
    .S1(net221),
    .X(_115_));
 sg13g2_nor2b_1 _398_ (.A(net215),
    .B_N(_115_),
    .Y(_116_));
 sg13g2_o21ai_1 _399_ (.B1(net4),
    .Y(_117_),
    .A1(_114_),
    .A2(_116_));
 sg13g2_nor2b_1 _400_ (.A(net231),
    .B_N(\u_dmtd.shift_reg[86] ),
    .Y(_118_));
 sg13g2_a21oi_1 _401_ (.A1(net231),
    .A2(\u_dmtd.shift_reg[87] ),
    .Y(_119_),
    .B1(_118_));
 sg13g2_mux2_1 _402_ (.A0(\u_dmtd.shift_reg[84] ),
    .A1(\u_dmtd.shift_reg[85] ),
    .S(net231),
    .X(_120_));
 sg13g2_o21ai_1 _403_ (.B1(net215),
    .Y(_121_),
    .A1(net221),
    .A2(_120_));
 sg13g2_a21oi_1 _404_ (.A1(net221),
    .A2(_119_),
    .Y(_122_),
    .B1(_121_));
 sg13g2_mux4_1 _405_ (.S0(net231),
    .A0(\u_dmtd.shift_reg[80] ),
    .A1(\u_dmtd.shift_reg[81] ),
    .A2(\u_dmtd.shift_reg[82] ),
    .A3(\u_dmtd.shift_reg[83] ),
    .S1(net221),
    .X(_123_));
 sg13g2_nor2b_1 _406_ (.A(net215),
    .B_N(_123_),
    .Y(_124_));
 sg13g2_o21ai_1 _407_ (.B1(_000_),
    .Y(_125_),
    .A1(_122_),
    .A2(_124_));
 sg13g2_a21o_1 _408_ (.A2(_125_),
    .A1(_117_),
    .B1(_001_),
    .X(_126_));
 sg13g2_nand2b_1 _409_ (.Y(_127_),
    .B(\u_dmtd.shift_reg[70] ),
    .A_N(net228));
 sg13g2_nand2_1 _410_ (.Y(_128_),
    .A(net228),
    .B(\u_dmtd.shift_reg[71] ));
 sg13g2_and3_1 _411_ (.X(_129_),
    .A(net219),
    .B(_127_),
    .C(_128_));
 sg13g2_mux2_1 _412_ (.A0(\u_dmtd.shift_reg[68] ),
    .A1(\u_dmtd.shift_reg[69] ),
    .S(net228),
    .X(_130_));
 sg13g2_o21ai_1 _413_ (.B1(net214),
    .Y(_131_),
    .A1(net219),
    .A2(_130_));
 sg13g2_mux4_1 _414_ (.S0(net228),
    .A0(\u_dmtd.shift_reg[64] ),
    .A1(\u_dmtd.shift_reg[65] ),
    .A2(\u_dmtd.shift_reg[66] ),
    .A3(\u_dmtd.shift_reg[67] ),
    .S1(net219),
    .X(_132_));
 sg13g2_nand2b_1 _415_ (.Y(_133_),
    .B(_132_),
    .A_N(net214));
 sg13g2_o21ai_1 _416_ (.B1(_133_),
    .Y(_134_),
    .A1(_129_),
    .A2(_131_));
 sg13g2_mux4_1 _417_ (.S0(net229),
    .A0(\u_dmtd.shift_reg[72] ),
    .A1(\u_dmtd.shift_reg[73] ),
    .A2(\u_dmtd.shift_reg[74] ),
    .A3(\u_dmtd.shift_reg[75] ),
    .S1(net219),
    .X(_135_));
 sg13g2_nand2b_1 _418_ (.Y(_136_),
    .B(_135_),
    .A_N(net214));
 sg13g2_nand2b_1 _419_ (.Y(_137_),
    .B(\u_dmtd.shift_reg[78] ),
    .A_N(net229));
 sg13g2_nand2_1 _420_ (.Y(_138_),
    .A(net228),
    .B(\u_dmtd.shift_reg[79] ));
 sg13g2_and3_1 _421_ (.X(_139_),
    .A(net219),
    .B(_137_),
    .C(_138_));
 sg13g2_mux2_1 _422_ (.A0(\u_dmtd.shift_reg[76] ),
    .A1(\u_dmtd.shift_reg[77] ),
    .S(net228),
    .X(_140_));
 sg13g2_o21ai_1 _423_ (.B1(net214),
    .Y(_141_),
    .A1(net219),
    .A2(_140_));
 sg13g2_o21ai_1 _424_ (.B1(_136_),
    .Y(_142_),
    .A1(_139_),
    .A2(_141_));
 sg13g2_mux2_1 _425_ (.A0(_134_),
    .A1(_142_),
    .S(net4),
    .X(_143_));
 sg13g2_a21oi_1 _426_ (.A1(_001_),
    .A2(_143_),
    .Y(_144_),
    .B1(net6));
 sg13g2_a22oi_1 _427_ (.Y(_145_),
    .B1(_126_),
    .B2(_144_),
    .A2(_109_),
    .A1(_108_));
 sg13g2_a221oi_1 _428_ (.B2(_074_),
    .C1(net7),
    .B1(_056_),
    .A1(_021_),
    .Y(_146_),
    .A2(_039_));
 sg13g2_a21o_1 _429_ (.A2(_145_),
    .A1(net7),
    .B1(_146_),
    .X(_147_));
 sg13g2_xnor2_1 _430_ (.Y(\u_dmtd.dmtd_out ),
    .A(_004_),
    .B(_147_));
 sg13g2_mux2_1 _431_ (.A0(\u_dmtd.async_reg2[2] ),
    .A1(\u_dmtd.async_reg1[2] ),
    .S(net3),
    .X(\u_dmtd.sync_out2 ));
 sg13g2_dfrbp_1 _432_ (.CLK(net259),
    .RESET_B(net283),
    .D(\u_dmtd.async_reg1[1] ),
    .Q_N(_149_),
    .Q(\u_dmtd.async_reg1[2] ));
 sg13g2_dfrbp_1 _433_ (.CLK(net259),
    .RESET_B(net283),
    .D(\u_dmtd.sync_out2 ),
    .Q_N(_150_),
    .Q(\u_dmtd.shift_reg[0] ));
 sg13g2_dfrbp_1 _434_ (.CLK(net258),
    .RESET_B(net282),
    .D(\u_dmtd.shift_reg[0] ),
    .Q_N(_151_),
    .Q(\u_dmtd.shift_reg[1] ));
 sg13g2_dfrbp_1 _435_ (.CLK(net258),
    .RESET_B(net282),
    .D(\u_dmtd.shift_reg[1] ),
    .Q_N(_152_),
    .Q(\u_dmtd.shift_reg[2] ));
 sg13g2_dfrbp_1 _436_ (.CLK(net258),
    .RESET_B(net282),
    .D(\u_dmtd.shift_reg[2] ),
    .Q_N(_153_),
    .Q(\u_dmtd.shift_reg[3] ));
 sg13g2_dfrbp_1 _437_ (.CLK(net258),
    .RESET_B(net282),
    .D(\u_dmtd.shift_reg[3] ),
    .Q_N(_154_),
    .Q(\u_dmtd.shift_reg[4] ));
 sg13g2_dfrbp_1 _438_ (.CLK(net258),
    .RESET_B(net282),
    .D(\u_dmtd.shift_reg[4] ),
    .Q_N(_155_),
    .Q(\u_dmtd.shift_reg[5] ));
 sg13g2_dfrbp_1 _439_ (.CLK(net258),
    .RESET_B(net282),
    .D(\u_dmtd.shift_reg[5] ),
    .Q_N(_156_),
    .Q(\u_dmtd.shift_reg[6] ));
 sg13g2_dfrbp_1 _440_ (.CLK(net260),
    .RESET_B(net284),
    .D(\u_dmtd.shift_reg[6] ),
    .Q_N(_157_),
    .Q(\u_dmtd.shift_reg[7] ));
 sg13g2_dfrbp_1 _441_ (.CLK(net260),
    .RESET_B(net284),
    .D(\u_dmtd.shift_reg[7] ),
    .Q_N(_158_),
    .Q(\u_dmtd.shift_reg[8] ));
 sg13g2_dfrbp_1 _442_ (.CLK(net257),
    .RESET_B(net281),
    .D(\u_dmtd.shift_reg[8] ),
    .Q_N(_159_),
    .Q(\u_dmtd.shift_reg[9] ));
 sg13g2_dfrbp_1 _443_ (.CLK(net257),
    .RESET_B(net281),
    .D(\u_dmtd.shift_reg[9] ),
    .Q_N(_160_),
    .Q(\u_dmtd.shift_reg[10] ));
 sg13g2_dfrbp_1 _444_ (.CLK(net257),
    .RESET_B(net281),
    .D(\u_dmtd.shift_reg[10] ),
    .Q_N(_161_),
    .Q(\u_dmtd.shift_reg[11] ));
 sg13g2_dfrbp_1 _445_ (.CLK(net257),
    .RESET_B(net281),
    .D(\u_dmtd.shift_reg[11] ),
    .Q_N(_162_),
    .Q(\u_dmtd.shift_reg[12] ));
 sg13g2_dfrbp_1 _446_ (.CLK(net256),
    .RESET_B(net280),
    .D(\u_dmtd.shift_reg[12] ),
    .Q_N(_163_),
    .Q(\u_dmtd.shift_reg[13] ));
 sg13g2_dfrbp_1 _447_ (.CLK(net256),
    .RESET_B(net280),
    .D(\u_dmtd.shift_reg[13] ),
    .Q_N(_164_),
    .Q(\u_dmtd.shift_reg[14] ));
 sg13g2_dfrbp_1 _448_ (.CLK(net257),
    .RESET_B(net281),
    .D(\u_dmtd.shift_reg[14] ),
    .Q_N(_165_),
    .Q(\u_dmtd.shift_reg[15] ));
 sg13g2_dfrbp_1 _449_ (.CLK(net257),
    .RESET_B(net281),
    .D(\u_dmtd.shift_reg[15] ),
    .Q_N(_166_),
    .Q(\u_dmtd.shift_reg[16] ));
 sg13g2_dfrbp_1 _450_ (.CLK(net249),
    .RESET_B(net273),
    .D(\u_dmtd.shift_reg[16] ),
    .Q_N(_167_),
    .Q(\u_dmtd.shift_reg[17] ));
 sg13g2_dfrbp_1 _451_ (.CLK(net249),
    .RESET_B(net273),
    .D(\u_dmtd.shift_reg[17] ),
    .Q_N(_168_),
    .Q(\u_dmtd.shift_reg[18] ));
 sg13g2_dfrbp_1 _452_ (.CLK(net248),
    .RESET_B(net272),
    .D(\u_dmtd.shift_reg[18] ),
    .Q_N(_169_),
    .Q(\u_dmtd.shift_reg[19] ));
 sg13g2_dfrbp_1 _453_ (.CLK(net248),
    .RESET_B(net272),
    .D(\u_dmtd.shift_reg[19] ),
    .Q_N(_170_),
    .Q(\u_dmtd.shift_reg[20] ));
 sg13g2_dfrbp_1 _454_ (.CLK(net248),
    .RESET_B(net272),
    .D(\u_dmtd.shift_reg[20] ),
    .Q_N(_171_),
    .Q(\u_dmtd.shift_reg[21] ));
 sg13g2_dfrbp_1 _455_ (.CLK(net248),
    .RESET_B(net272),
    .D(\u_dmtd.shift_reg[21] ),
    .Q_N(_172_),
    .Q(\u_dmtd.shift_reg[22] ));
 sg13g2_dfrbp_1 _456_ (.CLK(net248),
    .RESET_B(net272),
    .D(\u_dmtd.shift_reg[22] ),
    .Q_N(_173_),
    .Q(\u_dmtd.shift_reg[23] ));
 sg13g2_dfrbp_1 _457_ (.CLK(net243),
    .RESET_B(net267),
    .D(\u_dmtd.shift_reg[23] ),
    .Q_N(_174_),
    .Q(\u_dmtd.shift_reg[24] ));
 sg13g2_dfrbp_1 _458_ (.CLK(net243),
    .RESET_B(net267),
    .D(\u_dmtd.shift_reg[24] ),
    .Q_N(_175_),
    .Q(\u_dmtd.shift_reg[25] ));
 sg13g2_dfrbp_1 _459_ (.CLK(net252),
    .RESET_B(net276),
    .D(\u_dmtd.shift_reg[25] ),
    .Q_N(_176_),
    .Q(\u_dmtd.shift_reg[26] ));
 sg13g2_dfrbp_1 _460_ (.CLK(net252),
    .RESET_B(net276),
    .D(\u_dmtd.shift_reg[26] ),
    .Q_N(_177_),
    .Q(\u_dmtd.shift_reg[27] ));
 sg13g2_dfrbp_1 _461_ (.CLK(net252),
    .RESET_B(net276),
    .D(\u_dmtd.shift_reg[27] ),
    .Q_N(_178_),
    .Q(\u_dmtd.shift_reg[28] ));
 sg13g2_dfrbp_1 _462_ (.CLK(net252),
    .RESET_B(net276),
    .D(\u_dmtd.shift_reg[28] ),
    .Q_N(_179_),
    .Q(\u_dmtd.shift_reg[29] ));
 sg13g2_dfrbp_1 _463_ (.CLK(net252),
    .RESET_B(net276),
    .D(\u_dmtd.shift_reg[29] ),
    .Q_N(_180_),
    .Q(\u_dmtd.shift_reg[30] ));
 sg13g2_dfrbp_1 _464_ (.CLK(net251),
    .RESET_B(net275),
    .D(\u_dmtd.shift_reg[30] ),
    .Q_N(_181_),
    .Q(\u_dmtd.shift_reg[31] ));
 sg13g2_dfrbp_1 _465_ (.CLK(net253),
    .RESET_B(net277),
    .D(\u_dmtd.shift_reg[31] ),
    .Q_N(_182_),
    .Q(\u_dmtd.shift_reg[32] ));
 sg13g2_dfrbp_1 _466_ (.CLK(net253),
    .RESET_B(net277),
    .D(\u_dmtd.shift_reg[32] ),
    .Q_N(_183_),
    .Q(\u_dmtd.shift_reg[33] ));
 sg13g2_dfrbp_1 _467_ (.CLK(net253),
    .RESET_B(net277),
    .D(\u_dmtd.shift_reg[33] ),
    .Q_N(_184_),
    .Q(\u_dmtd.shift_reg[34] ));
 sg13g2_dfrbp_1 _468_ (.CLK(net253),
    .RESET_B(net277),
    .D(\u_dmtd.shift_reg[34] ),
    .Q_N(_185_),
    .Q(\u_dmtd.shift_reg[35] ));
 sg13g2_dfrbp_1 _469_ (.CLK(net253),
    .RESET_B(net277),
    .D(\u_dmtd.shift_reg[35] ),
    .Q_N(_186_),
    .Q(\u_dmtd.shift_reg[36] ));
 sg13g2_dfrbp_1 _470_ (.CLK(net253),
    .RESET_B(net277),
    .D(\u_dmtd.shift_reg[36] ),
    .Q_N(_187_),
    .Q(\u_dmtd.shift_reg[37] ));
 sg13g2_dfrbp_1 _471_ (.CLK(net255),
    .RESET_B(net279),
    .D(\u_dmtd.shift_reg[37] ),
    .Q_N(_188_),
    .Q(\u_dmtd.shift_reg[38] ));
 sg13g2_dfrbp_1 _472_ (.CLK(net253),
    .RESET_B(net277),
    .D(\u_dmtd.shift_reg[38] ),
    .Q_N(_189_),
    .Q(\u_dmtd.shift_reg[39] ));
 sg13g2_dfrbp_1 _473_ (.CLK(net253),
    .RESET_B(net277),
    .D(\u_dmtd.shift_reg[39] ),
    .Q_N(_190_),
    .Q(\u_dmtd.shift_reg[40] ));
 sg13g2_dfrbp_1 _474_ (.CLK(net251),
    .RESET_B(net275),
    .D(\u_dmtd.shift_reg[40] ),
    .Q_N(_191_),
    .Q(\u_dmtd.shift_reg[41] ));
 sg13g2_dfrbp_1 _475_ (.CLK(net251),
    .RESET_B(net275),
    .D(\u_dmtd.shift_reg[41] ),
    .Q_N(_192_),
    .Q(\u_dmtd.shift_reg[42] ));
 sg13g2_dfrbp_1 _476_ (.CLK(net251),
    .RESET_B(net275),
    .D(\u_dmtd.shift_reg[42] ),
    .Q_N(_193_),
    .Q(\u_dmtd.shift_reg[43] ));
 sg13g2_dfrbp_1 _477_ (.CLK(net251),
    .RESET_B(net275),
    .D(\u_dmtd.shift_reg[43] ),
    .Q_N(_194_),
    .Q(\u_dmtd.shift_reg[44] ));
 sg13g2_dfrbp_1 _478_ (.CLK(net251),
    .RESET_B(net275),
    .D(\u_dmtd.shift_reg[44] ),
    .Q_N(_195_),
    .Q(\u_dmtd.shift_reg[45] ));
 sg13g2_dfrbp_1 _479_ (.CLK(net251),
    .RESET_B(net275),
    .D(\u_dmtd.shift_reg[45] ),
    .Q_N(_196_),
    .Q(\u_dmtd.shift_reg[46] ));
 sg13g2_dfrbp_1 _480_ (.CLK(net251),
    .RESET_B(net275),
    .D(\u_dmtd.shift_reg[46] ),
    .Q_N(_197_),
    .Q(\u_dmtd.shift_reg[47] ));
 sg13g2_dfrbp_1 _481_ (.CLK(net242),
    .RESET_B(net266),
    .D(\u_dmtd.shift_reg[47] ),
    .Q_N(_198_),
    .Q(\u_dmtd.shift_reg[48] ));
 sg13g2_dfrbp_1 _482_ (.CLK(net242),
    .RESET_B(net266),
    .D(\u_dmtd.shift_reg[48] ),
    .Q_N(_199_),
    .Q(\u_dmtd.shift_reg[49] ));
 sg13g2_dfrbp_1 _483_ (.CLK(net242),
    .RESET_B(net266),
    .D(\u_dmtd.shift_reg[49] ),
    .Q_N(_200_),
    .Q(\u_dmtd.shift_reg[50] ));
 sg13g2_dfrbp_1 _484_ (.CLK(net242),
    .RESET_B(net266),
    .D(\u_dmtd.shift_reg[50] ),
    .Q_N(_201_),
    .Q(\u_dmtd.shift_reg[51] ));
 sg13g2_dfrbp_1 _485_ (.CLK(net242),
    .RESET_B(net266),
    .D(\u_dmtd.shift_reg[51] ),
    .Q_N(_202_),
    .Q(\u_dmtd.shift_reg[52] ));
 sg13g2_dfrbp_1 _486_ (.CLK(net242),
    .RESET_B(net266),
    .D(\u_dmtd.shift_reg[52] ),
    .Q_N(_203_),
    .Q(\u_dmtd.shift_reg[53] ));
 sg13g2_dfrbp_1 _487_ (.CLK(net242),
    .RESET_B(net266),
    .D(\u_dmtd.shift_reg[53] ),
    .Q_N(_204_),
    .Q(\u_dmtd.shift_reg[54] ));
 sg13g2_dfrbp_1 _488_ (.CLK(net242),
    .RESET_B(net266),
    .D(\u_dmtd.shift_reg[54] ),
    .Q_N(_205_),
    .Q(\u_dmtd.shift_reg[55] ));
 sg13g2_dfrbp_1 _489_ (.CLK(net243),
    .RESET_B(net267),
    .D(\u_dmtd.shift_reg[55] ),
    .Q_N(_206_),
    .Q(\u_dmtd.shift_reg[56] ));
 sg13g2_dfrbp_1 _490_ (.CLK(net243),
    .RESET_B(net267),
    .D(\u_dmtd.shift_reg[56] ),
    .Q_N(_207_),
    .Q(\u_dmtd.shift_reg[57] ));
 sg13g2_dfrbp_1 _491_ (.CLK(net243),
    .RESET_B(net267),
    .D(\u_dmtd.shift_reg[57] ),
    .Q_N(_208_),
    .Q(\u_dmtd.shift_reg[58] ));
 sg13g2_dfrbp_1 _492_ (.CLK(net243),
    .RESET_B(net267),
    .D(\u_dmtd.shift_reg[58] ),
    .Q_N(_209_),
    .Q(\u_dmtd.shift_reg[59] ));
 sg13g2_dfrbp_1 _493_ (.CLK(net241),
    .RESET_B(net265),
    .D(\u_dmtd.shift_reg[59] ),
    .Q_N(_210_),
    .Q(\u_dmtd.shift_reg[60] ));
 sg13g2_dfrbp_1 _494_ (.CLK(net240),
    .RESET_B(net264),
    .D(\u_dmtd.shift_reg[60] ),
    .Q_N(_211_),
    .Q(\u_dmtd.shift_reg[61] ));
 sg13g2_dfrbp_1 _495_ (.CLK(net239),
    .RESET_B(net263),
    .D(\u_dmtd.shift_reg[61] ),
    .Q_N(_212_),
    .Q(\u_dmtd.shift_reg[62] ));
 sg13g2_dfrbp_1 _496_ (.CLK(net241),
    .RESET_B(net265),
    .D(\u_dmtd.shift_reg[62] ),
    .Q_N(_213_),
    .Q(\u_dmtd.shift_reg[63] ));
 sg13g2_dfrbp_1 _497_ (.CLK(net241),
    .RESET_B(net265),
    .D(\u_dmtd.shift_reg[63] ),
    .Q_N(_214_),
    .Q(\u_dmtd.shift_reg[64] ));
 sg13g2_dfrbp_1 _498_ (.CLK(net241),
    .RESET_B(net265),
    .D(\u_dmtd.shift_reg[64] ),
    .Q_N(_215_),
    .Q(\u_dmtd.shift_reg[65] ));
 sg13g2_dfrbp_1 _499_ (.CLK(net239),
    .RESET_B(net263),
    .D(\u_dmtd.shift_reg[65] ),
    .Q_N(_216_),
    .Q(\u_dmtd.shift_reg[66] ));
 sg13g2_dfrbp_1 _500_ (.CLK(net239),
    .RESET_B(net263),
    .D(\u_dmtd.shift_reg[66] ),
    .Q_N(_217_),
    .Q(\u_dmtd.shift_reg[67] ));
 sg13g2_dfrbp_1 _501_ (.CLK(net239),
    .RESET_B(net263),
    .D(\u_dmtd.shift_reg[67] ),
    .Q_N(_218_),
    .Q(\u_dmtd.shift_reg[68] ));
 sg13g2_dfrbp_1 _502_ (.CLK(net239),
    .RESET_B(net263),
    .D(\u_dmtd.shift_reg[68] ),
    .Q_N(_219_),
    .Q(\u_dmtd.shift_reg[69] ));
 sg13g2_dfrbp_1 _503_ (.CLK(net239),
    .RESET_B(net263),
    .D(\u_dmtd.shift_reg[69] ),
    .Q_N(_220_),
    .Q(\u_dmtd.shift_reg[70] ));
 sg13g2_dfrbp_1 _504_ (.CLK(net239),
    .RESET_B(net263),
    .D(\u_dmtd.shift_reg[70] ),
    .Q_N(_221_),
    .Q(\u_dmtd.shift_reg[71] ));
 sg13g2_dfrbp_1 _505_ (.CLK(net239),
    .RESET_B(net263),
    .D(\u_dmtd.shift_reg[71] ),
    .Q_N(_222_),
    .Q(\u_dmtd.shift_reg[72] ));
 sg13g2_dfrbp_1 _506_ (.CLK(net240),
    .RESET_B(net264),
    .D(\u_dmtd.shift_reg[72] ),
    .Q_N(_223_),
    .Q(\u_dmtd.shift_reg[73] ));
 sg13g2_dfrbp_1 _507_ (.CLK(net240),
    .RESET_B(net264),
    .D(\u_dmtd.shift_reg[73] ),
    .Q_N(_224_),
    .Q(\u_dmtd.shift_reg[74] ));
 sg13g2_dfrbp_1 _508_ (.CLK(net240),
    .RESET_B(net264),
    .D(\u_dmtd.shift_reg[74] ),
    .Q_N(_225_),
    .Q(\u_dmtd.shift_reg[75] ));
 sg13g2_dfrbp_1 _509_ (.CLK(net240),
    .RESET_B(net264),
    .D(\u_dmtd.shift_reg[75] ),
    .Q_N(_226_),
    .Q(\u_dmtd.shift_reg[76] ));
 sg13g2_dfrbp_1 _510_ (.CLK(net240),
    .RESET_B(net264),
    .D(\u_dmtd.shift_reg[76] ),
    .Q_N(_227_),
    .Q(\u_dmtd.shift_reg[77] ));
 sg13g2_dfrbp_1 _511_ (.CLK(net240),
    .RESET_B(net264),
    .D(\u_dmtd.shift_reg[77] ),
    .Q_N(_228_),
    .Q(\u_dmtd.shift_reg[78] ));
 sg13g2_dfrbp_1 _512_ (.CLK(net240),
    .RESET_B(net264),
    .D(\u_dmtd.shift_reg[78] ),
    .Q_N(_229_),
    .Q(\u_dmtd.shift_reg[79] ));
 sg13g2_dfrbp_1 _513_ (.CLK(net244),
    .RESET_B(net268),
    .D(\u_dmtd.shift_reg[79] ),
    .Q_N(_230_),
    .Q(\u_dmtd.shift_reg[80] ));
 sg13g2_dfrbp_1 _514_ (.CLK(net244),
    .RESET_B(net268),
    .D(\u_dmtd.shift_reg[80] ),
    .Q_N(_231_),
    .Q(\u_dmtd.shift_reg[81] ));
 sg13g2_dfrbp_1 _515_ (.CLK(net244),
    .RESET_B(net268),
    .D(\u_dmtd.shift_reg[81] ),
    .Q_N(_232_),
    .Q(\u_dmtd.shift_reg[82] ));
 sg13g2_dfrbp_1 _516_ (.CLK(net244),
    .RESET_B(net268),
    .D(\u_dmtd.shift_reg[82] ),
    .Q_N(_233_),
    .Q(\u_dmtd.shift_reg[83] ));
 sg13g2_dfrbp_1 _517_ (.CLK(net244),
    .RESET_B(net268),
    .D(\u_dmtd.shift_reg[83] ),
    .Q_N(_234_),
    .Q(\u_dmtd.shift_reg[84] ));
 sg13g2_dfrbp_1 _518_ (.CLK(net244),
    .RESET_B(net268),
    .D(\u_dmtd.shift_reg[84] ),
    .Q_N(_235_),
    .Q(\u_dmtd.shift_reg[85] ));
 sg13g2_dfrbp_1 _519_ (.CLK(net247),
    .RESET_B(net271),
    .D(\u_dmtd.shift_reg[85] ),
    .Q_N(_236_),
    .Q(\u_dmtd.shift_reg[86] ));
 sg13g2_dfrbp_1 _520_ (.CLK(net244),
    .RESET_B(net268),
    .D(\u_dmtd.shift_reg[86] ),
    .Q_N(_237_),
    .Q(\u_dmtd.shift_reg[87] ));
 sg13g2_dfrbp_1 _521_ (.CLK(net244),
    .RESET_B(net268),
    .D(\u_dmtd.shift_reg[87] ),
    .Q_N(_238_),
    .Q(\u_dmtd.shift_reg[88] ));
 sg13g2_dfrbp_1 _522_ (.CLK(net245),
    .RESET_B(net269),
    .D(\u_dmtd.shift_reg[88] ),
    .Q_N(_239_),
    .Q(\u_dmtd.shift_reg[89] ));
 sg13g2_dfrbp_1 _523_ (.CLK(net245),
    .RESET_B(net269),
    .D(\u_dmtd.shift_reg[89] ),
    .Q_N(_240_),
    .Q(\u_dmtd.shift_reg[90] ));
 sg13g2_dfrbp_1 _524_ (.CLK(net245),
    .RESET_B(net269),
    .D(\u_dmtd.shift_reg[90] ),
    .Q_N(_241_),
    .Q(\u_dmtd.shift_reg[91] ));
 sg13g2_dfrbp_1 _525_ (.CLK(net245),
    .RESET_B(net269),
    .D(\u_dmtd.shift_reg[91] ),
    .Q_N(_242_),
    .Q(\u_dmtd.shift_reg[92] ));
 sg13g2_dfrbp_1 _526_ (.CLK(net245),
    .RESET_B(net269),
    .D(\u_dmtd.shift_reg[92] ),
    .Q_N(_243_),
    .Q(\u_dmtd.shift_reg[93] ));
 sg13g2_dfrbp_1 _527_ (.CLK(net245),
    .RESET_B(net269),
    .D(\u_dmtd.shift_reg[93] ),
    .Q_N(_244_),
    .Q(\u_dmtd.shift_reg[94] ));
 sg13g2_dfrbp_1 _528_ (.CLK(net245),
    .RESET_B(net269),
    .D(\u_dmtd.shift_reg[94] ),
    .Q_N(_245_),
    .Q(\u_dmtd.shift_reg[95] ));
 sg13g2_dfrbp_1 _529_ (.CLK(net245),
    .RESET_B(net269),
    .D(\u_dmtd.shift_reg[95] ),
    .Q_N(_246_),
    .Q(\u_dmtd.shift_reg[96] ));
 sg13g2_dfrbp_1 _530_ (.CLK(net246),
    .RESET_B(net270),
    .D(\u_dmtd.shift_reg[96] ),
    .Q_N(_247_),
    .Q(\u_dmtd.shift_reg[97] ));
 sg13g2_dfrbp_1 _531_ (.CLK(net246),
    .RESET_B(net270),
    .D(\u_dmtd.shift_reg[97] ),
    .Q_N(_248_),
    .Q(\u_dmtd.shift_reg[98] ));
 sg13g2_dfrbp_1 _532_ (.CLK(net246),
    .RESET_B(net270),
    .D(\u_dmtd.shift_reg[98] ),
    .Q_N(_249_),
    .Q(\u_dmtd.shift_reg[99] ));
 sg13g2_dfrbp_1 _533_ (.CLK(net246),
    .RESET_B(net270),
    .D(\u_dmtd.shift_reg[99] ),
    .Q_N(_250_),
    .Q(\u_dmtd.shift_reg[100] ));
 sg13g2_dfrbp_1 _534_ (.CLK(net248),
    .RESET_B(net272),
    .D(\u_dmtd.shift_reg[100] ),
    .Q_N(_251_),
    .Q(\u_dmtd.shift_reg[101] ));
 sg13g2_dfrbp_1 _535_ (.CLK(net249),
    .RESET_B(net273),
    .D(\u_dmtd.shift_reg[101] ),
    .Q_N(_252_),
    .Q(\u_dmtd.shift_reg[102] ));
 sg13g2_dfrbp_1 _536_ (.CLK(net248),
    .RESET_B(net272),
    .D(\u_dmtd.shift_reg[102] ),
    .Q_N(_253_),
    .Q(\u_dmtd.shift_reg[103] ));
 sg13g2_dfrbp_1 _537_ (.CLK(net248),
    .RESET_B(net272),
    .D(\u_dmtd.shift_reg[103] ),
    .Q_N(_254_),
    .Q(\u_dmtd.shift_reg[104] ));
 sg13g2_dfrbp_1 _538_ (.CLK(net256),
    .RESET_B(net280),
    .D(\u_dmtd.shift_reg[104] ),
    .Q_N(_255_),
    .Q(\u_dmtd.shift_reg[105] ));
 sg13g2_dfrbp_1 _539_ (.CLK(net256),
    .RESET_B(net280),
    .D(\u_dmtd.shift_reg[105] ),
    .Q_N(_256_),
    .Q(\u_dmtd.shift_reg[106] ));
 sg13g2_dfrbp_1 _540_ (.CLK(net256),
    .RESET_B(net280),
    .D(\u_dmtd.shift_reg[106] ),
    .Q_N(_257_),
    .Q(\u_dmtd.shift_reg[107] ));
 sg13g2_dfrbp_1 _541_ (.CLK(net256),
    .RESET_B(net280),
    .D(\u_dmtd.shift_reg[107] ),
    .Q_N(_258_),
    .Q(\u_dmtd.shift_reg[108] ));
 sg13g2_dfrbp_1 _542_ (.CLK(net256),
    .RESET_B(net280),
    .D(\u_dmtd.shift_reg[108] ),
    .Q_N(_259_),
    .Q(\u_dmtd.shift_reg[109] ));
 sg13g2_dfrbp_1 _543_ (.CLK(net256),
    .RESET_B(net280),
    .D(\u_dmtd.shift_reg[109] ),
    .Q_N(_260_),
    .Q(\u_dmtd.shift_reg[110] ));
 sg13g2_dfrbp_1 _544_ (.CLK(net261),
    .RESET_B(net285),
    .D(\u_dmtd.shift_reg[110] ),
    .Q_N(_261_),
    .Q(\u_dmtd.shift_reg[111] ));
 sg13g2_dfrbp_1 _545_ (.CLK(net261),
    .RESET_B(net285),
    .D(\u_dmtd.shift_reg[111] ),
    .Q_N(_262_),
    .Q(\u_dmtd.shift_reg[112] ));
 sg13g2_dfrbp_1 _546_ (.CLK(net261),
    .RESET_B(net285),
    .D(\u_dmtd.shift_reg[112] ),
    .Q_N(_263_),
    .Q(\u_dmtd.shift_reg[113] ));
 sg13g2_dfrbp_1 _547_ (.CLK(net261),
    .RESET_B(net285),
    .D(\u_dmtd.shift_reg[113] ),
    .Q_N(_264_),
    .Q(\u_dmtd.shift_reg[114] ));
 sg13g2_dfrbp_1 _548_ (.CLK(net261),
    .RESET_B(net285),
    .D(\u_dmtd.shift_reg[114] ),
    .Q_N(_265_),
    .Q(\u_dmtd.shift_reg[115] ));
 sg13g2_dfrbp_1 _549_ (.CLK(net261),
    .RESET_B(net285),
    .D(\u_dmtd.shift_reg[115] ),
    .Q_N(_266_),
    .Q(\u_dmtd.shift_reg[116] ));
 sg13g2_dfrbp_1 _550_ (.CLK(net261),
    .RESET_B(net285),
    .D(\u_dmtd.shift_reg[116] ),
    .Q_N(_267_),
    .Q(\u_dmtd.shift_reg[117] ));
 sg13g2_dfrbp_1 _551_ (.CLK(net255),
    .RESET_B(net279),
    .D(\u_dmtd.shift_reg[117] ),
    .Q_N(_268_),
    .Q(\u_dmtd.shift_reg[118] ));
 sg13g2_dfrbp_1 _552_ (.CLK(net255),
    .RESET_B(net279),
    .D(\u_dmtd.shift_reg[118] ),
    .Q_N(_269_),
    .Q(\u_dmtd.shift_reg[119] ));
 sg13g2_dfrbp_1 _553_ (.CLK(net254),
    .RESET_B(net278),
    .D(\u_dmtd.shift_reg[119] ),
    .Q_N(_270_),
    .Q(\u_dmtd.shift_reg[120] ));
 sg13g2_dfrbp_1 _554_ (.CLK(net254),
    .RESET_B(net278),
    .D(\u_dmtd.shift_reg[120] ),
    .Q_N(_271_),
    .Q(\u_dmtd.shift_reg[121] ));
 sg13g2_dfrbp_1 _555_ (.CLK(net254),
    .RESET_B(net278),
    .D(\u_dmtd.shift_reg[121] ),
    .Q_N(_272_),
    .Q(\u_dmtd.shift_reg[122] ));
 sg13g2_dfrbp_1 _556_ (.CLK(net254),
    .RESET_B(net278),
    .D(\u_dmtd.shift_reg[122] ),
    .Q_N(_273_),
    .Q(\u_dmtd.shift_reg[123] ));
 sg13g2_dfrbp_1 _557_ (.CLK(net254),
    .RESET_B(net278),
    .D(\u_dmtd.shift_reg[123] ),
    .Q_N(_274_),
    .Q(\u_dmtd.shift_reg[124] ));
 sg13g2_dfrbp_1 _558_ (.CLK(net254),
    .RESET_B(net278),
    .D(\u_dmtd.shift_reg[124] ),
    .Q_N(_275_),
    .Q(\u_dmtd.shift_reg[125] ));
 sg13g2_dfrbp_1 _559_ (.CLK(net254),
    .RESET_B(net278),
    .D(\u_dmtd.shift_reg[125] ),
    .Q_N(_276_),
    .Q(\u_dmtd.shift_reg[126] ));
 sg13g2_dfrbp_1 _560_ (.CLK(net254),
    .RESET_B(net278),
    .D(\u_dmtd.shift_reg[126] ),
    .Q_N(_277_),
    .Q(\u_dmtd.shift_reg[127] ));
 sg13g2_dfrbp_1 _561_ (.CLK(net259),
    .RESET_B(net283),
    .D(net2),
    .Q_N(_278_),
    .Q(\u_dmtd.async_reg2[0] ));
 sg13g2_dfrbp_1 _562_ (.CLK(net259),
    .RESET_B(net283),
    .D(\u_dmtd.async_reg2[0] ),
    .Q_N(_279_),
    .Q(\u_dmtd.async_reg2[1] ));
 sg13g2_dfrbp_1 _563_ (.CLK(net259),
    .RESET_B(net283),
    .D(\u_dmtd.async_reg2[1] ),
    .Q_N(_280_),
    .Q(\u_dmtd.async_reg2[2] ));
 sg13g2_dfrbp_1 _564_ (.CLK(net258),
    .RESET_B(net282),
    .D(net1),
    .Q_N(_281_),
    .Q(\u_dmtd.async_reg1[0] ));
 sg13g2_dfrbp_1 _565_ (.CLK(net258),
    .RESET_B(net282),
    .D(\u_dmtd.async_reg1[0] ),
    .Q_N(_148_),
    .Q(\u_dmtd.async_reg1[1] ));
 sg13g2_tielo tt_um_dmtd_arghunter_9 (.L_LO(net9));
 sg13g2_tielo tt_um_dmtd_arghunter_10 (.L_LO(net10));
 sg13g2_tielo tt_um_dmtd_arghunter_11 (.L_LO(net11));
 sg13g2_tielo tt_um_dmtd_arghunter_12 (.L_LO(net12));
 sg13g2_tielo tt_um_dmtd_arghunter_13 (.L_LO(net13));
 sg13g2_tielo tt_um_dmtd_arghunter_14 (.L_LO(net14));
 sg13g2_tielo tt_um_dmtd_arghunter_15 (.L_LO(net15));
 sg13g2_tielo tt_um_dmtd_arghunter_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dmtd_arghunter_17 (.L_LO(net17));
 sg13g2_tielo tt_um_dmtd_arghunter_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dmtd_arghunter_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dmtd_arghunter_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dmtd_arghunter_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dmtd_arghunter_22 (.L_LO(net22));
 sg13g2_tielo tt_um_dmtd_arghunter_23 (.L_LO(net23));
 sg13g2_tielo tt_um_dmtd_arghunter_24 (.L_LO(net24));
 sg13g2_tielo tt_um_dmtd_arghunter_25 (.L_LO(net25));
 sg13g2_tielo tt_um_dmtd_arghunter_26 (.L_LO(net26));
 sg13g2_tielo tt_um_dmtd_arghunter_27 (.L_LO(net27));
 sg13g2_tielo tt_um_dmtd_arghunter_28 (.L_LO(net28));
 sg13g2_tielo tt_um_dmtd_arghunter_29 (.L_LO(net29));
 sg13g2_tielo tt_um_dmtd_arghunter_30 (.L_LO(net30));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 _589_ (.A(\u_dmtd.dmtd_out ),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout214 (.A(net218),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(net218),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(net218),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(net218),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(uio_in[3]),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(net223),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(net223),
    .X(net220));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(net223));
 sg13g2_buf_1 fanout222 (.A(net223),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(uio_in[2]),
    .X(net223));
 sg13g2_buf_4 fanout224 (.X(net224),
    .A(net227));
 sg13g2_buf_2 fanout225 (.A(net227),
    .X(net225));
 sg13g2_buf_4 fanout226 (.X(net226),
    .A(net227));
 sg13g2_buf_2 fanout227 (.A(uio_in[2]),
    .X(net227));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(net230));
 sg13g2_buf_2 fanout229 (.A(net230),
    .X(net229));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(net238));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(net232));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(net238));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(net234));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(net237));
 sg13g2_buf_4 fanout235 (.X(net235),
    .A(net237));
 sg13g2_buf_2 fanout236 (.A(net237),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(net238),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(uio_in[1]),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(net241),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(net250),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(net250),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(net250),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(net247),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(net247),
    .X(net245));
 sg13g2_buf_1 fanout246 (.A(net247),
    .X(net246));
 sg13g2_buf_1 fanout247 (.A(net249),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(net249),
    .X(net248));
 sg13g2_buf_1 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_1 fanout250 (.A(ui_in[0]),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(net262),
    .X(net251));
 sg13g2_buf_1 fanout252 (.A(net262),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net255),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(net255),
    .X(net254));
 sg13g2_buf_1 fanout255 (.A(net262),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(net262),
    .X(net256));
 sg13g2_buf_1 fanout257 (.A(net262),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net260),
    .X(net258));
 sg13g2_buf_1 fanout259 (.A(net260),
    .X(net259));
 sg13g2_buf_1 fanout260 (.A(net261),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(net262),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(ui_in[0]),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(net265));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(net265));
 sg13g2_buf_2 fanout265 (.A(net274),
    .X(net265));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(net274));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(net274));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(net271));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(net271));
 sg13g2_buf_2 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(net273),
    .X(net271));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(net273));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(rst_n),
    .X(net274));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(net286));
 sg13g2_buf_2 fanout276 (.A(net286),
    .X(net276));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(net279));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(net279));
 sg13g2_buf_2 fanout279 (.A(net286),
    .X(net279));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(net286));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(net286));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(net284));
 sg13g2_buf_2 fanout283 (.A(net284),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(net285),
    .X(net284));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(net286));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[0]),
    .X(net3));
 sg13g2_buf_4 input4 (.X(net4),
    .A(uio_in[4]));
 sg13g2_buf_1 input5 (.A(uio_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[6]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[7]),
    .X(net7));
 sg13g2_tielo tt_um_dmtd_arghunter_8 (.L_LO(net8));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_fill_2 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_4 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_95 ();
 sg13g2_decap_8 FILLER_17_122 ();
 sg13g2_decap_4 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_4 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_decap_8 FILLER_17_220 ();
 sg13g2_decap_4 FILLER_17_227 ();
 sg13g2_fill_2 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_fill_2 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_fill_2 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_124 ();
 sg13g2_fill_2 FILLER_18_131 ();
 sg13g2_decap_8 FILLER_18_185 ();
 sg13g2_decap_4 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_decap_4 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_fill_2 FILLER_18_267 ();
 sg13g2_fill_1 FILLER_18_269 ();
 sg13g2_decap_8 FILLER_18_296 ();
 sg13g2_decap_8 FILLER_18_303 ();
 sg13g2_fill_2 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_fill_2 FILLER_19_128 ();
 sg13g2_decap_8 FILLER_19_187 ();
 sg13g2_decap_8 FILLER_19_194 ();
 sg13g2_fill_2 FILLER_19_201 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_fill_2 FILLER_19_303 ();
 sg13g2_fill_1 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_332 ();
 sg13g2_decap_8 FILLER_19_339 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_4 FILLER_20_84 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_174 ();
 sg13g2_decap_8 FILLER_20_181 ();
 sg13g2_decap_8 FILLER_20_188 ();
 sg13g2_fill_1 FILLER_20_195 ();
 sg13g2_decap_8 FILLER_20_222 ();
 sg13g2_decap_4 FILLER_20_229 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_fill_2 FILLER_20_280 ();
 sg13g2_fill_1 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_304 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_fill_2 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_370 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_4 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_4 FILLER_21_189 ();
 sg13g2_fill_1 FILLER_21_193 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_254 ();
 sg13g2_fill_2 FILLER_21_261 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_290 ();
 sg13g2_decap_4 FILLER_21_297 ();
 sg13g2_fill_1 FILLER_21_301 ();
 sg13g2_fill_2 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_fill_2 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_86 ();
 sg13g2_decap_8 FILLER_22_113 ();
 sg13g2_decap_8 FILLER_22_120 ();
 sg13g2_decap_4 FILLER_22_127 ();
 sg13g2_fill_1 FILLER_22_131 ();
 sg13g2_decap_4 FILLER_22_137 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_decap_8 FILLER_22_148 ();
 sg13g2_fill_1 FILLER_22_155 ();
 sg13g2_fill_2 FILLER_22_166 ();
 sg13g2_fill_2 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_decap_4 FILLER_22_215 ();
 sg13g2_fill_1 FILLER_22_219 ();
 sg13g2_decap_4 FILLER_22_225 ();
 sg13g2_decap_8 FILLER_22_239 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_262 ();
 sg13g2_fill_2 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_4 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_2 FILLER_23_130 ();
 sg13g2_fill_1 FILLER_23_132 ();
 sg13g2_fill_2 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_fill_2 FILLER_23_185 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_246 ();
 sg13g2_decap_4 FILLER_23_253 ();
 sg13g2_fill_2 FILLER_23_257 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_332 ();
 sg13g2_fill_1 FILLER_23_338 ();
 sg13g2_fill_2 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_fill_1 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_367 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_4 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_176 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_301 ();
 sg13g2_fill_2 FILLER_24_316 ();
 sg13g2_decap_4 FILLER_24_323 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_4 FILLER_24_338 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_decap_4 FILLER_24_364 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_84 ();
 sg13g2_decap_4 FILLER_25_124 ();
 sg13g2_decap_8 FILLER_25_164 ();
 sg13g2_decap_4 FILLER_25_171 ();
 sg13g2_decap_8 FILLER_25_180 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_decap_4 FILLER_25_221 ();
 sg13g2_decap_4 FILLER_25_251 ();
 sg13g2_decap_4 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_291 ();
 sg13g2_decap_8 FILLER_25_298 ();
 sg13g2_fill_2 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_375 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_110 ();
 sg13g2_decap_8 FILLER_26_117 ();
 sg13g2_decap_8 FILLER_26_124 ();
 sg13g2_decap_8 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_159 ();
 sg13g2_decap_4 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_170 ();
 sg13g2_decap_4 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_184 ();
 sg13g2_decap_4 FILLER_26_191 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_decap_4 FILLER_26_207 ();
 sg13g2_decap_4 FILLER_26_215 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_255 ();
 sg13g2_decap_8 FILLER_26_262 ();
 sg13g2_decap_4 FILLER_26_269 ();
 sg13g2_fill_2 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_302 ();
 sg13g2_fill_2 FILLER_26_361 ();
 sg13g2_fill_1 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_132 ();
 sg13g2_decap_8 FILLER_27_139 ();
 sg13g2_decap_8 FILLER_27_146 ();
 sg13g2_decap_8 FILLER_27_153 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_fill_1 FILLER_27_162 ();
 sg13g2_fill_1 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_fill_2 FILLER_27_222 ();
 sg13g2_decap_8 FILLER_27_239 ();
 sg13g2_decap_8 FILLER_27_246 ();
 sg13g2_decap_8 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_262 ();
 sg13g2_fill_2 FILLER_27_268 ();
 sg13g2_decap_4 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_decap_4 FILLER_27_367 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_146 ();
 sg13g2_decap_8 FILLER_28_153 ();
 sg13g2_decap_4 FILLER_28_160 ();
 sg13g2_fill_2 FILLER_28_164 ();
 sg13g2_decap_8 FILLER_28_248 ();
 sg13g2_decap_8 FILLER_28_255 ();
 sg13g2_decap_8 FILLER_28_262 ();
 sg13g2_decap_8 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_276 ();
 sg13g2_decap_8 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_313 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_decap_4 FILLER_28_332 ();
 sg13g2_fill_2 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_4 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_4 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_148 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_fill_2 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_decap_8 FILLER_29_299 ();
 sg13g2_decap_8 FILLER_29_306 ();
 sg13g2_fill_2 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_decap_8 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_29_352 ();
 sg13g2_decap_8 FILLER_29_359 ();
 sg13g2_decap_8 FILLER_29_366 ();
 sg13g2_decap_4 FILLER_29_373 ();
 sg13g2_fill_1 FILLER_29_377 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_186 ();
 sg13g2_decap_8 FILLER_30_193 ();
 sg13g2_decap_4 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_204 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_fill_1 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_302 ();
 sg13g2_fill_2 FILLER_30_309 ();
 sg13g2_decap_4 FILLER_30_347 ();
 sg13g2_fill_2 FILLER_30_351 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_4 FILLER_31_105 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_decap_8 FILLER_31_172 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_decap_8 FILLER_31_226 ();
 sg13g2_decap_4 FILLER_31_233 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_333 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_decap_8 FILLER_32_120 ();
 sg13g2_fill_1 FILLER_32_127 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_decap_4 FILLER_32_143 ();
 sg13g2_decap_4 FILLER_32_162 ();
 sg13g2_decap_8 FILLER_32_223 ();
 sg13g2_decap_8 FILLER_32_230 ();
 sg13g2_decap_8 FILLER_32_237 ();
 sg13g2_fill_2 FILLER_32_244 ();
 sg13g2_fill_1 FILLER_32_246 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_decap_8 FILLER_32_332 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_fill_1 FILLER_32_350 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_137 ();
 sg13g2_decap_4 FILLER_33_144 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_decap_4 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_164 ();
 sg13g2_decap_8 FILLER_33_232 ();
 sg13g2_decap_8 FILLER_33_239 ();
 sg13g2_fill_2 FILLER_33_246 ();
 sg13g2_fill_1 FILLER_33_248 ();
 sg13g2_decap_8 FILLER_33_297 ();
 sg13g2_decap_8 FILLER_33_304 ();
 sg13g2_fill_2 FILLER_33_311 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_157 ();
 sg13g2_decap_4 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_216 ();
 sg13g2_decap_4 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_227 ();
 sg13g2_decap_8 FILLER_34_242 ();
 sg13g2_decap_8 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_256 ();
 sg13g2_fill_2 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_285 ();
 sg13g2_decap_8 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_299 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_163 ();
 sg13g2_fill_1 FILLER_35_174 ();
 sg13g2_fill_2 FILLER_35_201 ();
 sg13g2_decap_8 FILLER_35_208 ();
 sg13g2_decap_4 FILLER_35_215 ();
 sg13g2_fill_2 FILLER_35_219 ();
 sg13g2_fill_1 FILLER_35_298 ();
 sg13g2_fill_2 FILLER_35_325 ();
 sg13g2_fill_2 FILLER_35_353 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_130 ();
 sg13g2_fill_2 FILLER_36_142 ();
 sg13g2_decap_4 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_174 ();
 sg13g2_decap_8 FILLER_36_201 ();
 sg13g2_decap_8 FILLER_36_208 ();
 sg13g2_decap_4 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_decap_4 FILLER_36_362 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_4 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_109 ();
 sg13g2_decap_8 FILLER_37_162 ();
 sg13g2_decap_4 FILLER_37_169 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_200 ();
 sg13g2_decap_8 FILLER_37_207 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_decap_8 FILLER_37_221 ();
 sg13g2_fill_2 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_292 ();
 sg13g2_fill_2 FILLER_37_299 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_4 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_fill_2 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_decap_4 FILLER_38_268 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_4 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_377 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net8;
 assign uio_oe[1] = net9;
 assign uio_oe[2] = net10;
 assign uio_oe[3] = net11;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
 assign uio_out[7] = net23;
 assign uo_out[1] = net24;
 assign uo_out[2] = net25;
 assign uo_out[3] = net26;
 assign uo_out[4] = net27;
 assign uo_out[5] = net28;
 assign uo_out[6] = net29;
 assign uo_out[7] = net30;
endmodule

module tt_um_virantha_enigma (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire \enigma.fsm.cnt[0] ;
 wire \enigma.fsm.cnt[1] ;
 wire \enigma.fsm.double_step ;
 wire \enigma.fsm.fsm_state[0] ;
 wire \enigma.fsm.fsm_state[1] ;
 wire \enigma.fsm.fsm_state[2] ;
 wire \enigma.fsm.fsm_state[3] ;
 wire \enigma.fsm.fsm_state[4] ;
 wire \enigma.fsm.ready ;
 wire \enigma.plugboard.$31[0] ;
 wire \enigma.plugboard.bits_0_0.clk ;
 wire \enigma.plugboard.bits_0_0.q ;
 wire \enigma.plugboard.bits_0_1.q ;
 wire \enigma.plugboard.bits_0_2.q ;
 wire \enigma.plugboard.bits_0_3.q ;
 wire \enigma.plugboard.bits_0_4.q ;
 wire \enigma.plugboard.bits_10_0.clk ;
 wire \enigma.plugboard.bits_10_0.q ;
 wire \enigma.plugboard.bits_10_1.q ;
 wire \enigma.plugboard.bits_10_2.q ;
 wire \enigma.plugboard.bits_10_3.q ;
 wire \enigma.plugboard.bits_10_4.q ;
 wire \enigma.plugboard.bits_11_0.clk ;
 wire \enigma.plugboard.bits_11_0.q ;
 wire \enigma.plugboard.bits_11_1.q ;
 wire \enigma.plugboard.bits_11_2.q ;
 wire \enigma.plugboard.bits_11_3.q ;
 wire \enigma.plugboard.bits_11_4.q ;
 wire \enigma.plugboard.bits_12_0.clk ;
 wire \enigma.plugboard.bits_12_0.q ;
 wire \enigma.plugboard.bits_12_1.q ;
 wire \enigma.plugboard.bits_12_2.q ;
 wire \enigma.plugboard.bits_12_3.q ;
 wire \enigma.plugboard.bits_12_4.q ;
 wire \enigma.plugboard.bits_13_0.clk ;
 wire \enigma.plugboard.bits_13_0.q ;
 wire \enigma.plugboard.bits_13_1.q ;
 wire \enigma.plugboard.bits_13_2.q ;
 wire \enigma.plugboard.bits_13_3.q ;
 wire \enigma.plugboard.bits_13_4.q ;
 wire \enigma.plugboard.bits_14_0.clk ;
 wire \enigma.plugboard.bits_14_0.q ;
 wire \enigma.plugboard.bits_14_1.q ;
 wire \enigma.plugboard.bits_14_2.q ;
 wire \enigma.plugboard.bits_14_3.q ;
 wire \enigma.plugboard.bits_14_4.q ;
 wire \enigma.plugboard.bits_15_0.clk ;
 wire \enigma.plugboard.bits_15_0.q ;
 wire \enigma.plugboard.bits_15_1.q ;
 wire \enigma.plugboard.bits_15_2.q ;
 wire \enigma.plugboard.bits_15_3.q ;
 wire \enigma.plugboard.bits_15_4.q ;
 wire \enigma.plugboard.bits_16_0.clk ;
 wire \enigma.plugboard.bits_16_0.q ;
 wire \enigma.plugboard.bits_16_1.q ;
 wire \enigma.plugboard.bits_16_2.q ;
 wire \enigma.plugboard.bits_16_3.q ;
 wire \enigma.plugboard.bits_16_4.q ;
 wire \enigma.plugboard.bits_17_0.clk ;
 wire \enigma.plugboard.bits_17_0.q ;
 wire \enigma.plugboard.bits_17_1.q ;
 wire \enigma.plugboard.bits_17_2.q ;
 wire \enigma.plugboard.bits_17_3.q ;
 wire \enigma.plugboard.bits_17_4.q ;
 wire \enigma.plugboard.bits_18_0.clk ;
 wire \enigma.plugboard.bits_18_0.q ;
 wire \enigma.plugboard.bits_18_1.q ;
 wire \enigma.plugboard.bits_18_2.q ;
 wire \enigma.plugboard.bits_18_3.q ;
 wire \enigma.plugboard.bits_18_4.q ;
 wire \enigma.plugboard.bits_19_0.clk ;
 wire \enigma.plugboard.bits_19_0.q ;
 wire \enigma.plugboard.bits_19_1.q ;
 wire \enigma.plugboard.bits_19_2.q ;
 wire \enigma.plugboard.bits_19_3.q ;
 wire \enigma.plugboard.bits_19_4.q ;
 wire \enigma.plugboard.bits_1_0.clk ;
 wire \enigma.plugboard.bits_1_0.q ;
 wire \enigma.plugboard.bits_1_1.q ;
 wire \enigma.plugboard.bits_1_2.q ;
 wire \enigma.plugboard.bits_1_3.q ;
 wire \enigma.plugboard.bits_1_4.q ;
 wire \enigma.plugboard.bits_20_0.clk ;
 wire \enigma.plugboard.bits_20_0.q ;
 wire \enigma.plugboard.bits_20_1.q ;
 wire \enigma.plugboard.bits_20_2.q ;
 wire \enigma.plugboard.bits_20_3.q ;
 wire \enigma.plugboard.bits_20_4.q ;
 wire \enigma.plugboard.bits_21_0.clk ;
 wire \enigma.plugboard.bits_21_0.q ;
 wire \enigma.plugboard.bits_21_1.q ;
 wire \enigma.plugboard.bits_21_2.q ;
 wire \enigma.plugboard.bits_21_3.q ;
 wire \enigma.plugboard.bits_21_4.q ;
 wire \enigma.plugboard.bits_22_0.clk ;
 wire \enigma.plugboard.bits_22_0.q ;
 wire \enigma.plugboard.bits_22_1.q ;
 wire \enigma.plugboard.bits_22_2.q ;
 wire \enigma.plugboard.bits_22_3.q ;
 wire \enigma.plugboard.bits_22_4.q ;
 wire \enigma.plugboard.bits_23_0.clk ;
 wire \enigma.plugboard.bits_23_0.q ;
 wire \enigma.plugboard.bits_23_1.q ;
 wire \enigma.plugboard.bits_23_2.q ;
 wire \enigma.plugboard.bits_23_3.q ;
 wire \enigma.plugboard.bits_23_4.q ;
 wire \enigma.plugboard.bits_24_0.clk ;
 wire \enigma.plugboard.bits_24_0.q ;
 wire \enigma.plugboard.bits_24_1.q ;
 wire \enigma.plugboard.bits_24_2.q ;
 wire \enigma.plugboard.bits_24_3.q ;
 wire \enigma.plugboard.bits_24_4.q ;
 wire \enigma.plugboard.bits_25_0.clk ;
 wire \enigma.plugboard.bits_25_0.q ;
 wire \enigma.plugboard.bits_25_1.q ;
 wire \enigma.plugboard.bits_25_2.q ;
 wire \enigma.plugboard.bits_25_3.q ;
 wire \enigma.plugboard.bits_25_4.q ;
 wire \enigma.plugboard.bits_2_0.clk ;
 wire \enigma.plugboard.bits_2_0.q ;
 wire \enigma.plugboard.bits_2_1.q ;
 wire \enigma.plugboard.bits_2_2.q ;
 wire \enigma.plugboard.bits_2_3.q ;
 wire \enigma.plugboard.bits_2_4.q ;
 wire \enigma.plugboard.bits_3_0.clk ;
 wire \enigma.plugboard.bits_3_0.q ;
 wire \enigma.plugboard.bits_3_1.q ;
 wire \enigma.plugboard.bits_3_2.q ;
 wire \enigma.plugboard.bits_3_3.q ;
 wire \enigma.plugboard.bits_3_4.q ;
 wire \enigma.plugboard.bits_4_0.clk ;
 wire \enigma.plugboard.bits_4_0.q ;
 wire \enigma.plugboard.bits_4_1.q ;
 wire \enigma.plugboard.bits_4_2.q ;
 wire \enigma.plugboard.bits_4_3.q ;
 wire \enigma.plugboard.bits_4_4.q ;
 wire \enigma.plugboard.bits_5_0.clk ;
 wire \enigma.plugboard.bits_5_0.q ;
 wire \enigma.plugboard.bits_5_1.q ;
 wire \enigma.plugboard.bits_5_2.q ;
 wire \enigma.plugboard.bits_5_3.q ;
 wire \enigma.plugboard.bits_5_4.q ;
 wire \enigma.plugboard.bits_6_0.clk ;
 wire \enigma.plugboard.bits_6_0.q ;
 wire \enigma.plugboard.bits_6_1.q ;
 wire \enigma.plugboard.bits_6_2.q ;
 wire \enigma.plugboard.bits_6_3.q ;
 wire \enigma.plugboard.bits_6_4.q ;
 wire \enigma.plugboard.bits_7_0.clk ;
 wire \enigma.plugboard.bits_7_0.q ;
 wire \enigma.plugboard.bits_7_1.q ;
 wire \enigma.plugboard.bits_7_2.q ;
 wire \enigma.plugboard.bits_7_3.q ;
 wire \enigma.plugboard.bits_7_4.q ;
 wire \enigma.plugboard.bits_8_0.clk ;
 wire \enigma.plugboard.bits_8_0.q ;
 wire \enigma.plugboard.bits_8_1.q ;
 wire \enigma.plugboard.bits_8_2.q ;
 wire \enigma.plugboard.bits_8_3.q ;
 wire \enigma.plugboard.bits_8_4.q ;
 wire \enigma.plugboard.bits_9_0.clk ;
 wire \enigma.plugboard.bits_9_0.q ;
 wire \enigma.plugboard.bits_9_1.q ;
 wire \enigma.plugboard.bits_9_2.q ;
 wire \enigma.plugboard.bits_9_3.q ;
 wire \enigma.plugboard.bits_9_4.q ;
 wire \enigma.plugboard.cnt[0] ;
 wire \enigma.plugboard.cnt[1] ;
 wire \enigma.plugboard.cnt[2] ;
 wire \enigma.plugboard.cnt[3] ;
 wire \enigma.plugboard.cnt[4] ;
 wire \enigma.plugboard.plug_limiter[0] ;
 wire \enigma.plugboard.plug_limiter[1] ;
 wire \enigma.plugboard.plug_limiter[2] ;
 wire \enigma.plugboard.plug_limiter[3] ;
 wire \enigma.plugboard.plug_limiter[4] ;
 wire \enigma.r.$signal$13[0] ;
 wire \enigma.r.$signal$13[1] ;
 wire \enigma.r.$signal$13[2] ;
 wire \enigma.r.$signal$13[3] ;
 wire \enigma.r.$signal$13[4] ;
 wire \enigma.r.$signal$17[0] ;
 wire \enigma.r.$signal$17[1] ;
 wire \enigma.r.$signal$17[2] ;
 wire \enigma.r.$signal$20[0] ;
 wire \enigma.r.$signal$20[1] ;
 wire \enigma.r.$signal$20[2] ;
 wire \enigma.r.$signal$20[3] ;
 wire \enigma.r.$signal$20[4] ;
 wire \enigma.r.$signal$21[0] ;
 wire \enigma.r.$signal$21[1] ;
 wire \enigma.r.$signal$21[2] ;
 wire \enigma.r.$signal$22[0] ;
 wire \enigma.r.$signal$22[1] ;
 wire \enigma.r.$signal$22[2] ;
 wire \enigma.r.$signal$22[3] ;
 wire \enigma.r.$signal$22[4] ;
 wire \enigma.r.$signal$23[0] ;
 wire \enigma.r.$signal$23[1] ;
 wire \enigma.r.$signal$23[2] ;
 wire \enigma.r.cnts_debug0[0] ;
 wire \enigma.r.cnts_debug0[1] ;
 wire \enigma.r.cnts_debug0[2] ;
 wire \enigma.r.cnts_debug0[3] ;
 wire \enigma.r.cnts_debug0[4] ;
 wire \enigma.r.cnts_debug1[0] ;
 wire \enigma.r.cnts_debug1[1] ;
 wire \enigma.r.cnts_debug1[2] ;
 wire \enigma.r.cnts_debug1[3] ;
 wire \enigma.r.cnts_debug1[4] ;
 wire \enigma.r.cnts_debug2[0] ;
 wire \enigma.r.cnts_debug2[1] ;
 wire \enigma.r.cnts_debug2[2] ;
 wire \enigma.r.cnts_debug2[3] ;
 wire \enigma.r.cnts_debug2[4] ;
 wire \enigma.r.dout[0] ;
 wire \enigma.r.dout[1] ;
 wire \enigma.r.dout[2] ;
 wire \enigma.r.dout[3] ;
 wire \enigma.r.dout[4] ;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire clknet_0_clk;
 wire net6;
 wire net7;
 wire net8;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;

 sg13g2_inv_1 _1402_ (.Y(_0638_),
    .A(net556));
 sg13g2_inv_1 _1403_ (.Y(_0639_),
    .A(net559));
 sg13g2_inv_1 _1404_ (.Y(_0640_),
    .A(net560));
 sg13g2_inv_2 _1405_ (.Y(_0641_),
    .A(net567));
 sg13g2_inv_1 _1406_ (.Y(_0642_),
    .A(net570));
 sg13g2_inv_1 _1407_ (.Y(_0643_),
    .A(net134));
 sg13g2_inv_1 _1408_ (.Y(_0644_),
    .A(net108));
 sg13g2_inv_1 _1409_ (.Y(_0645_),
    .A(net589));
 sg13g2_inv_1 _1410_ (.Y(_0646_),
    .A(net130));
 sg13g2_inv_1 _1411_ (.Y(_0647_),
    .A(net136));
 sg13g2_inv_1 _1412_ (.Y(_0648_),
    .A(net597));
 sg13g2_inv_2 _1413_ (.Y(_0649_),
    .A(net135));
 sg13g2_inv_1 _1414_ (.Y(_0650_),
    .A(net603));
 sg13g2_inv_1 _1415_ (.Y(_0651_),
    .A(net141));
 sg13g2_inv_1 _1416_ (.Y(_0652_),
    .A(net606));
 sg13g2_inv_1 _1417_ (.Y(_0653_),
    .A(net83));
 sg13g2_inv_1 _1418_ (.Y(_0654_),
    .A(\enigma.r.cnts_debug0[0] ));
 sg13g2_inv_1 _1419_ (.Y(_0655_),
    .A(\enigma.r.cnts_debug1[4] ));
 sg13g2_inv_1 _1420_ (.Y(_0656_),
    .A(\enigma.r.cnts_debug1[0] ));
 sg13g2_inv_1 _1421_ (.Y(_0657_),
    .A(\enigma.r.cnts_debug2[2] ));
 sg13g2_inv_1 _1422_ (.Y(_0658_),
    .A(\enigma.r.cnts_debug2[1] ));
 sg13g2_inv_1 _1423_ (.Y(_0659_),
    .A(\enigma.r.cnts_debug2[0] ));
 sg13g2_inv_1 _1424_ (.Y(_0660_),
    .A(\enigma.r.$signal$22[2] ));
 sg13g2_inv_1 _1425_ (.Y(_0661_),
    .A(\enigma.r.$signal$22[1] ));
 sg13g2_inv_1 _1426_ (.Y(_0662_),
    .A(\enigma.r.$signal$22[0] ));
 sg13g2_inv_2 _1427_ (.Y(_0663_),
    .A(net582));
 sg13g2_inv_1 _1428_ (.Y(_0664_),
    .A(\enigma.r.dout[4] ));
 sg13g2_inv_1 _1429_ (.Y(_0665_),
    .A(\enigma.r.dout[1] ));
 sg13g2_inv_1 _1430_ (.Y(_0666_),
    .A(net581));
 sg13g2_inv_4 _1431_ (.A(net616),
    .Y(_0667_));
 sg13g2_nor2_2 _1432_ (.A(net573),
    .B(_0643_),
    .Y(_0668_));
 sg13g2_nor2_1 _1433_ (.A(net569),
    .B(net571),
    .Y(_0669_));
 sg13g2_or2_1 _1434_ (.X(_0670_),
    .B(net571),
    .A(net569));
 sg13g2_nor3_2 _1435_ (.A(net570),
    .B(net572),
    .C(net573),
    .Y(_0671_));
 sg13g2_nand2_2 _1436_ (.Y(_0672_),
    .A(net575),
    .B(_0671_));
 sg13g2_nor2_1 _1437_ (.A(net567),
    .B(_0672_),
    .Y(\enigma.fsm.ready ));
 sg13g2_inv_1 _1438_ (.Y(_0673_),
    .A(\enigma.fsm.ready ));
 sg13g2_nand2_2 _1439_ (.Y(_0674_),
    .A(_0640_),
    .B(net564));
 sg13g2_a21oi_1 _1440_ (.A1(_0640_),
    .A2(uio_out[0]),
    .Y(_0675_),
    .B1(net558));
 sg13g2_nor2_1 _1441_ (.A(uio_out[1]),
    .B(uio_out[0]),
    .Y(_0676_));
 sg13g2_or2_1 _1442_ (.X(_0677_),
    .B(net564),
    .A(uio_out[1]));
 sg13g2_o21ai_1 _1443_ (.B1(_0675_),
    .Y(_0678_),
    .A1(_0640_),
    .A2(_0677_));
 sg13g2_and2_2 _1444_ (.A(uio_out[1]),
    .B(net564),
    .X(_0679_));
 sg13g2_o21ai_1 _1445_ (.B1(net560),
    .Y(_0680_),
    .A1(_0676_),
    .A2(_0679_));
 sg13g2_nand2_1 _1446_ (.Y(_0681_),
    .A(_0640_),
    .B(uio_out[1]));
 sg13g2_nor2b_1 _1447_ (.A(uio_out[0]),
    .B_N(uio_out[1]),
    .Y(_0682_));
 sg13g2_o21ai_1 _1448_ (.B1(_0680_),
    .Y(_0683_),
    .A1(uio_out[0]),
    .A2(_0681_));
 sg13g2_xor2_1 _1449_ (.B(_0683_),
    .A(_0678_),
    .X(_0684_));
 sg13g2_o21ai_1 _1450_ (.B1(net559),
    .Y(_0685_),
    .A1(uio_out[1]),
    .A2(_0674_));
 sg13g2_o21ai_1 _1451_ (.B1(_0639_),
    .Y(_0686_),
    .A1(net560),
    .A2(uio_out[0]));
 sg13g2_nand3_1 _1452_ (.B(_0685_),
    .C(_0686_),
    .A(uio_out[4]),
    .Y(_0687_));
 sg13g2_o21ai_1 _1453_ (.B1(_0687_),
    .Y(uo_out[0]),
    .A1(uio_out[4]),
    .A2(_0684_));
 sg13g2_nor2_1 _1454_ (.A(uio_out[2]),
    .B(uio_out[1]),
    .Y(_0688_));
 sg13g2_nor3_1 _1455_ (.A(net560),
    .B(net562),
    .C(uio_out[0]),
    .Y(_0689_));
 sg13g2_nor2_1 _1456_ (.A(_0679_),
    .B(_0689_),
    .Y(_0690_));
 sg13g2_nor3_1 _1457_ (.A(net559),
    .B(_0679_),
    .C(_0689_),
    .Y(_0691_));
 sg13g2_a21oi_1 _1458_ (.A1(net560),
    .A2(_0679_),
    .Y(_0692_),
    .B1(_0685_));
 sg13g2_or3_1 _1459_ (.A(uio_out[4]),
    .B(_0691_),
    .C(_0692_),
    .X(_0693_));
 sg13g2_nand3_1 _1460_ (.B(net558),
    .C(_0688_),
    .A(net556),
    .Y(_0694_));
 sg13g2_nand4_1 _1461_ (.B(_0675_),
    .C(_0680_),
    .A(net556),
    .Y(_0695_),
    .D(_0681_));
 sg13g2_nand3_1 _1462_ (.B(_0694_),
    .C(_0695_),
    .A(_0693_),
    .Y(uo_out[1]));
 sg13g2_nand2b_1 _1463_ (.Y(_0696_),
    .B(net556),
    .A_N(_0689_));
 sg13g2_o21ai_1 _1464_ (.B1(_0696_),
    .Y(_0697_),
    .A1(net556),
    .A2(_0690_));
 sg13g2_nand2_1 _1465_ (.Y(_0698_),
    .A(uio_out[2]),
    .B(_0682_));
 sg13g2_nand2_1 _1466_ (.Y(_0699_),
    .A(_0674_),
    .B(_0698_));
 sg13g2_and4_1 _1467_ (.A(_0638_),
    .B(_0674_),
    .C(_0691_),
    .D(_0698_),
    .X(_0700_));
 sg13g2_o21ai_1 _1468_ (.B1(_0698_),
    .Y(_0701_),
    .A1(net560),
    .A2(_0005_));
 sg13g2_nor2_1 _1469_ (.A(_0638_),
    .B(net558),
    .Y(_0702_));
 sg13g2_a221oi_1 _1470_ (.B2(_0702_),
    .C1(_0700_),
    .B1(_0701_),
    .A1(net559),
    .Y(uo_out[2]),
    .A2(_0697_));
 sg13g2_nor2_1 _1471_ (.A(net556),
    .B(_0675_),
    .Y(_0703_));
 sg13g2_nor2_1 _1472_ (.A(net558),
    .B(_0688_),
    .Y(_0704_));
 sg13g2_nand2b_1 _1473_ (.Y(_0705_),
    .B(net560),
    .A_N(_0005_));
 sg13g2_a22oi_1 _1474_ (.Y(_0706_),
    .B1(_0704_),
    .B2(_0705_),
    .A2(_0703_),
    .A1(_0699_));
 sg13g2_nand2_1 _1475_ (.Y(uo_out[3]),
    .A(_0694_),
    .B(_0706_));
 sg13g2_a21o_1 _1476_ (.A2(_0685_),
    .A1(_0678_),
    .B1(_0003_),
    .X(uo_out[4]));
 sg13g2_a21oi_1 _1477_ (.A1(_0677_),
    .A2(_0704_),
    .Y(_0707_),
    .B1(_0696_));
 sg13g2_nor2_1 _1478_ (.A(net558),
    .B(_0681_),
    .Y(_0708_));
 sg13g2_nor2b_1 _1479_ (.A(net564),
    .B_N(_0004_),
    .Y(_0709_));
 sg13g2_nor3_1 _1480_ (.A(_0639_),
    .B(_0679_),
    .C(_0709_),
    .Y(_0710_));
 sg13g2_or2_1 _1481_ (.X(_0711_),
    .B(_0710_),
    .A(_0708_));
 sg13g2_a21oi_2 _1482_ (.B1(_0707_),
    .Y(uo_out[5]),
    .A2(_0711_),
    .A1(_0638_));
 sg13g2_nand3_1 _1483_ (.B(_0674_),
    .C(_0677_),
    .A(net558),
    .Y(_0712_));
 sg13g2_o21ai_1 _1484_ (.B1(_0712_),
    .Y(_0713_),
    .A1(net558),
    .A2(_0682_));
 sg13g2_a21oi_1 _1485_ (.A1(net556),
    .A2(_0679_),
    .Y(_0714_),
    .B1(_0004_));
 sg13g2_o21ai_1 _1486_ (.B1(_0694_),
    .Y(_0715_),
    .A1(net558),
    .A2(_0714_));
 sg13g2_a21o_1 _1487_ (.A2(_0713_),
    .A1(_0638_),
    .B1(_0715_),
    .X(uo_out[6]));
 sg13g2_nand2_2 _1488_ (.Y(_0716_),
    .A(_0649_),
    .B(\enigma.plugboard.cnt[0] ));
 sg13g2_nand3b_1 _1489_ (.B(net566),
    .C(net574),
    .Y(_0717_),
    .A_N(net575));
 sg13g2_nor2b_2 _1490_ (.A(net570),
    .B_N(net572),
    .Y(_0718_));
 sg13g2_nor2b_2 _1491_ (.A(_0717_),
    .B_N(_0718_),
    .Y(_0719_));
 sg13g2_a21oi_1 _1492_ (.A1(\enigma.plugboard.plug_limiter[2] ),
    .A2(\enigma.plugboard.plug_limiter[1] ),
    .Y(_0720_),
    .B1(\enigma.plugboard.plug_limiter[3] ));
 sg13g2_nand3b_1 _1493_ (.B(_0719_),
    .C(_0720_),
    .Y(_0721_),
    .A_N(\enigma.plugboard.plug_limiter[4] ));
 sg13g2_nor2_2 _1494_ (.A(\enigma.plugboard.cnt[4] ),
    .B(_0721_),
    .Y(_0722_));
 sg13g2_nor2_1 _1495_ (.A(\enigma.plugboard.cnt[3] ),
    .B(_0647_),
    .Y(_0723_));
 sg13g2_nand2_2 _1496_ (.Y(_0724_),
    .A(_0722_),
    .B(_0723_));
 sg13g2_nor2_2 _1497_ (.A(_0716_),
    .B(_0724_),
    .Y(\enigma.plugboard.bits_5_0.clk ));
 sg13g2_nand2_2 _1498_ (.Y(_0725_),
    .A(_0649_),
    .B(_0651_));
 sg13g2_nor2_2 _1499_ (.A(_0724_),
    .B(_0725_),
    .Y(\enigma.plugboard.bits_4_0.clk ));
 sg13g2_nand2_2 _1500_ (.Y(_0726_),
    .A(\enigma.plugboard.cnt[1] ),
    .B(\enigma.plugboard.cnt[0] ));
 sg13g2_nor2_1 _1501_ (.A(\enigma.plugboard.cnt[3] ),
    .B(\enigma.plugboard.cnt[2] ),
    .Y(_0727_));
 sg13g2_nand2_2 _1502_ (.Y(_0728_),
    .A(_0722_),
    .B(_0727_));
 sg13g2_nor2_2 _1503_ (.A(_0726_),
    .B(_0728_),
    .Y(\enigma.plugboard.bits_3_0.clk ));
 sg13g2_nand2_2 _1504_ (.Y(_0729_),
    .A(\enigma.plugboard.cnt[1] ),
    .B(_0651_));
 sg13g2_nor2_2 _1505_ (.A(_0728_),
    .B(_0729_),
    .Y(\enigma.plugboard.bits_2_0.clk ));
 sg13g2_nor2_2 _1506_ (.A(_0716_),
    .B(_0728_),
    .Y(\enigma.plugboard.bits_1_0.clk ));
 sg13g2_nor2_2 _1507_ (.A(_0725_),
    .B(_0728_),
    .Y(\enigma.plugboard.bits_0_0.clk ));
 sg13g2_nor2_1 _1508_ (.A(_0007_),
    .B(_0721_),
    .Y(_0730_));
 sg13g2_or2_1 _1509_ (.X(_0731_),
    .B(_0721_),
    .A(_0007_));
 sg13g2_nand2_1 _1510_ (.Y(_0732_),
    .A(\enigma.plugboard.cnt[3] ),
    .B(_0647_));
 sg13g2_nor3_2 _1511_ (.A(_0716_),
    .B(_0731_),
    .C(_0732_),
    .Y(\enigma.plugboard.bits_25_0.clk ));
 sg13g2_nor3_2 _1512_ (.A(_0725_),
    .B(_0731_),
    .C(_0732_),
    .Y(\enigma.plugboard.bits_24_0.clk ));
 sg13g2_nand2_2 _1513_ (.Y(_0733_),
    .A(_0723_),
    .B(_0730_));
 sg13g2_nor2_2 _1514_ (.A(_0726_),
    .B(_0733_),
    .Y(\enigma.plugboard.bits_23_0.clk ));
 sg13g2_nor2_2 _1515_ (.A(_0729_),
    .B(_0733_),
    .Y(\enigma.plugboard.bits_22_0.clk ));
 sg13g2_nor2_2 _1516_ (.A(_0716_),
    .B(_0733_),
    .Y(\enigma.plugboard.bits_21_0.clk ));
 sg13g2_nor2_2 _1517_ (.A(_0725_),
    .B(_0733_),
    .Y(\enigma.plugboard.bits_20_0.clk ));
 sg13g2_nand2_2 _1518_ (.Y(_0734_),
    .A(_0727_),
    .B(_0730_));
 sg13g2_nor2_2 _1519_ (.A(_0726_),
    .B(_0734_),
    .Y(\enigma.plugboard.bits_19_0.clk ));
 sg13g2_nor2_2 _1520_ (.A(_0729_),
    .B(_0734_),
    .Y(\enigma.plugboard.bits_18_0.clk ));
 sg13g2_nor2_2 _1521_ (.A(_0716_),
    .B(_0734_),
    .Y(\enigma.plugboard.bits_17_0.clk ));
 sg13g2_nor2_2 _1522_ (.A(_0725_),
    .B(_0734_),
    .Y(\enigma.plugboard.bits_16_0.clk ));
 sg13g2_nand3_1 _1523_ (.B(\enigma.plugboard.cnt[2] ),
    .C(_0722_),
    .A(\enigma.plugboard.cnt[3] ),
    .Y(_0735_));
 sg13g2_nor2_2 _1524_ (.A(_0726_),
    .B(_0735_),
    .Y(\enigma.plugboard.bits_15_0.clk ));
 sg13g2_nor2_2 _1525_ (.A(_0729_),
    .B(_0735_),
    .Y(\enigma.plugboard.bits_14_0.clk ));
 sg13g2_nor2_2 _1526_ (.A(_0716_),
    .B(_0735_),
    .Y(\enigma.plugboard.bits_13_0.clk ));
 sg13g2_nor2_2 _1527_ (.A(_0725_),
    .B(_0735_),
    .Y(\enigma.plugboard.bits_12_0.clk ));
 sg13g2_nand3_1 _1528_ (.B(_0647_),
    .C(_0722_),
    .A(\enigma.plugboard.cnt[3] ),
    .Y(_0736_));
 sg13g2_nor2_2 _1529_ (.A(_0726_),
    .B(_0736_),
    .Y(\enigma.plugboard.bits_11_0.clk ));
 sg13g2_nor2_2 _1530_ (.A(_0729_),
    .B(_0736_),
    .Y(\enigma.plugboard.bits_10_0.clk ));
 sg13g2_nor2_2 _1531_ (.A(_0716_),
    .B(_0736_),
    .Y(\enigma.plugboard.bits_9_0.clk ));
 sg13g2_nor2_2 _1532_ (.A(_0725_),
    .B(_0736_),
    .Y(\enigma.plugboard.bits_8_0.clk ));
 sg13g2_nor2_2 _1533_ (.A(_0724_),
    .B(_0726_),
    .Y(\enigma.plugboard.bits_7_0.clk ));
 sg13g2_nor2_2 _1534_ (.A(_0724_),
    .B(_0729_),
    .Y(\enigma.plugboard.bits_6_0.clk ));
 sg13g2_and2_2 _1535_ (.A(net568),
    .B(_0671_),
    .X(_0737_));
 sg13g2_nand2_2 _1536_ (.Y(_0738_),
    .A(net568),
    .B(_0671_));
 sg13g2_nor2_2 _1537_ (.A(net574),
    .B(net575),
    .Y(_0739_));
 sg13g2_nand2_2 _1538_ (.Y(_0740_),
    .A(net570),
    .B(net572));
 sg13g2_nor3_2 _1539_ (.A(net568),
    .B(_0739_),
    .C(_0740_),
    .Y(_0741_));
 sg13g2_or3_2 _1540_ (.A(net568),
    .B(_0739_),
    .C(_0740_),
    .X(_0742_));
 sg13g2_nor2_2 _1541_ (.A(_0737_),
    .B(_0741_),
    .Y(_0743_));
 sg13g2_nand2_2 _1542_ (.Y(_0744_),
    .A(_0738_),
    .B(_0742_));
 sg13g2_and2_1 _1543_ (.A(net573),
    .B(net575),
    .X(_0745_));
 sg13g2_nand3_1 _1544_ (.B(_0669_),
    .C(_0745_),
    .A(_0641_),
    .Y(_0746_));
 sg13g2_nor2_2 _1545_ (.A(_0670_),
    .B(_0717_),
    .Y(_0747_));
 sg13g2_or2_2 _1546_ (.X(_0748_),
    .B(_0717_),
    .A(_0670_));
 sg13g2_nand3_1 _1547_ (.B(_0718_),
    .C(_0739_),
    .A(net565),
    .Y(_0749_));
 sg13g2_nand3_1 _1548_ (.B(_0748_),
    .C(_0749_),
    .A(_0746_),
    .Y(_0750_));
 sg13g2_nand2_1 _1549_ (.Y(_0751_),
    .A(\enigma.fsm.cnt[0] ),
    .B(_0750_));
 sg13g2_inv_1 _1550_ (.Y(_0752_),
    .A(net542));
 sg13g2_nor4_1 _1551_ (.A(net567),
    .B(net573),
    .C(_0643_),
    .D(_0740_),
    .Y(_0753_));
 sg13g2_nand3_1 _1552_ (.B(net573),
    .C(net575),
    .A(net567),
    .Y(_0754_));
 sg13g2_nor2_1 _1553_ (.A(_0670_),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_and4_1 _1554_ (.A(net569),
    .B(net571),
    .C(net565),
    .D(_0739_),
    .X(_0756_));
 sg13g2_nand4_1 _1555_ (.B(net572),
    .C(net566),
    .A(net570),
    .Y(_0757_),
    .D(_0739_));
 sg13g2_nor3_2 _1556_ (.A(_0753_),
    .B(_0755_),
    .C(_0756_),
    .Y(_0758_));
 sg13g2_nand4_1 _1557_ (.B(net571),
    .C(net565),
    .A(net569),
    .Y(_0759_),
    .D(_0745_));
 sg13g2_nor2b_1 _1558_ (.A(net571),
    .B_N(net569),
    .Y(_0760_));
 sg13g2_nor2b_1 _1559_ (.A(_0717_),
    .B_N(_0760_),
    .Y(_0761_));
 sg13g2_nand2_1 _1560_ (.Y(_0762_),
    .A(_0718_),
    .B(_0745_));
 sg13g2_and3_1 _1561_ (.X(_0763_),
    .A(net565),
    .B(_0718_),
    .C(_0745_));
 sg13g2_nor2_1 _1562_ (.A(_0761_),
    .B(_0763_),
    .Y(_0764_));
 sg13g2_and3_1 _1563_ (.X(_0765_),
    .A(_0758_),
    .B(_0759_),
    .C(_0764_));
 sg13g2_nand3_1 _1564_ (.B(_0759_),
    .C(_0764_),
    .A(_0758_),
    .Y(_0766_));
 sg13g2_nand2_1 _1565_ (.Y(_0767_),
    .A(\enigma.fsm.cnt[1] ),
    .B(_0750_));
 sg13g2_or2_1 _1566_ (.X(_0768_),
    .B(_0740_),
    .A(_0717_));
 sg13g2_nand2_1 _1567_ (.Y(_0769_),
    .A(net566),
    .B(_0668_));
 sg13g2_nand3_1 _1568_ (.B(_0668_),
    .C(_0760_),
    .A(net565),
    .Y(_0770_));
 sg13g2_nand3_1 _1569_ (.B(_0745_),
    .C(_0760_),
    .A(net565),
    .Y(_0771_));
 sg13g2_and4_1 _1570_ (.A(_0758_),
    .B(_0768_),
    .C(_0770_),
    .D(_0771_),
    .X(_0772_));
 sg13g2_nand4_1 _1571_ (.B(_0768_),
    .C(_0770_),
    .A(_0758_),
    .Y(_0773_),
    .D(_0771_));
 sg13g2_nand2_1 _1572_ (.Y(_0774_),
    .A(net540),
    .B(net539));
 sg13g2_a22oi_1 _1573_ (.Y(_0775_),
    .B1(net540),
    .B2(net539),
    .A2(net541),
    .A1(net542));
 sg13g2_a221oi_1 _1574_ (.B2(net539),
    .C1(_0659_),
    .B1(net540),
    .A1(net542),
    .Y(_0776_),
    .A2(net541));
 sg13g2_a221oi_1 _1575_ (.B2(net539),
    .C1(_0766_),
    .B1(net540),
    .A1(\enigma.fsm.cnt[0] ),
    .Y(_0777_),
    .A2(_0750_));
 sg13g2_nand3_1 _1576_ (.B(net541),
    .C(_0774_),
    .A(net542),
    .Y(_0778_));
 sg13g2_a221oi_1 _1577_ (.B2(net541),
    .C1(_0773_),
    .B1(_0751_),
    .A1(\enigma.fsm.cnt[1] ),
    .Y(_0779_),
    .A2(_0750_));
 sg13g2_inv_1 _1578_ (.Y(_0780_),
    .A(net521));
 sg13g2_a22oi_1 _1579_ (.Y(_0781_),
    .B1(net521),
    .B2(\enigma.r.cnts_debug0[0] ),
    .A2(net524),
    .A1(\enigma.r.cnts_debug1[0] ));
 sg13g2_a221oi_1 _1580_ (.B2(\enigma.r.cnts_debug0[0] ),
    .C1(_0776_),
    .B1(net521),
    .A1(\enigma.r.cnts_debug1[0] ),
    .Y(_0782_),
    .A2(net524));
 sg13g2_nand2b_1 _1581_ (.Y(_0783_),
    .B(_0781_),
    .A_N(_0776_));
 sg13g2_a221oi_1 _1582_ (.B2(_0772_),
    .C1(_0662_),
    .B1(_0767_),
    .A1(_0751_),
    .Y(_0784_),
    .A2(_0765_));
 sg13g2_a221oi_1 _1583_ (.B2(\enigma.r.$signal$13[0] ),
    .C1(_0784_),
    .B1(net522),
    .A1(\enigma.r.$signal$20[0] ),
    .Y(_0785_),
    .A2(net524));
 sg13g2_nand2b_1 _1584_ (.Y(_0786_),
    .B(_0782_),
    .A_N(_0785_));
 sg13g2_xor2_1 _1585_ (.B(_0785_),
    .A(_0782_),
    .X(_0787_));
 sg13g2_inv_1 _1586_ (.Y(_0788_),
    .A(_0787_));
 sg13g2_nor2_1 _1587_ (.A(\enigma.r.$signal$23[1] ),
    .B(\enigma.r.$signal$23[0] ),
    .Y(_0789_));
 sg13g2_o21ai_1 _1588_ (.B1(net525),
    .Y(_0790_),
    .A1(_0000_),
    .A2(_0789_));
 sg13g2_inv_2 _1589_ (.Y(_0791_),
    .A(_0790_));
 sg13g2_and2_1 _1590_ (.A(_0000_),
    .B(_0789_),
    .X(_0792_));
 sg13g2_nor3_2 _1591_ (.A(_0009_),
    .B(_0010_),
    .C(_0769_),
    .Y(_0793_));
 sg13g2_nor2_1 _1592_ (.A(net572),
    .B(net575),
    .Y(_0794_));
 sg13g2_nor4_2 _1593_ (.A(net567),
    .B(_0642_),
    .C(_0668_),
    .Y(_0795_),
    .D(_0794_));
 sg13g2_nor2_2 _1594_ (.A(_0793_),
    .B(_0795_),
    .Y(_0796_));
 sg13g2_o21ai_1 _1595_ (.B1(net569),
    .Y(_0797_),
    .A1(net571),
    .A2(net573));
 sg13g2_a21oi_1 _1596_ (.A1(_0762_),
    .A2(_0797_),
    .Y(_0798_),
    .B1(net568));
 sg13g2_nor2_1 _1597_ (.A(_0737_),
    .B(_0798_),
    .Y(_0799_));
 sg13g2_o21ai_1 _1598_ (.B1(_0665_),
    .Y(_0800_),
    .A1(_0737_),
    .A2(_0741_));
 sg13g2_nand3_1 _1599_ (.B(_0738_),
    .C(_0742_),
    .A(_0650_),
    .Y(_0801_));
 sg13g2_nand3_1 _1600_ (.B(_0738_),
    .C(_0742_),
    .A(net602),
    .Y(_0802_));
 sg13g2_o21ai_1 _1601_ (.B1(\enigma.r.dout[1] ),
    .Y(_0803_),
    .A1(_0737_),
    .A2(_0741_));
 sg13g2_nand3_1 _1602_ (.B(_0802_),
    .C(_0803_),
    .A(_0799_),
    .Y(_0804_));
 sg13g2_a21o_1 _1603_ (.A2(_0742_),
    .A1(_0738_),
    .B1(net585),
    .X(_0805_));
 sg13g2_nand3_1 _1604_ (.B(_0738_),
    .C(_0742_),
    .A(_0652_),
    .Y(_0806_));
 sg13g2_nand3_1 _1605_ (.B(_0738_),
    .C(_0742_),
    .A(net606),
    .Y(_0807_));
 sg13g2_o21ai_1 _1606_ (.B1(net585),
    .Y(_0808_),
    .A1(_0737_),
    .A2(_0741_));
 sg13g2_nand4_1 _1607_ (.B(_0803_),
    .C(_0805_),
    .A(_0802_),
    .Y(_0809_),
    .D(_0806_));
 sg13g2_nand3_1 _1608_ (.B(_0738_),
    .C(_0742_),
    .A(net592),
    .Y(_0810_));
 sg13g2_o21ai_1 _1609_ (.B1(net581),
    .Y(_0811_),
    .A1(_0737_),
    .A2(_0741_));
 sg13g2_nand2_1 _1610_ (.Y(_0812_),
    .A(_0810_),
    .B(_0811_));
 sg13g2_and2_1 _1611_ (.A(_0810_),
    .B(_0811_),
    .X(_0813_));
 sg13g2_mux2_1 _1612_ (.A0(net588),
    .A1(net580),
    .S(_0744_),
    .X(_0814_));
 sg13g2_mux2_1 _1613_ (.A0(_0645_),
    .A1(_0664_),
    .S(_0744_),
    .X(_0815_));
 sg13g2_mux2_1 _1614_ (.A0(net598),
    .A1(\enigma.r.dout[2] ),
    .S(_0744_),
    .X(_0816_));
 sg13g2_mux2_1 _1615_ (.A0(_0648_),
    .A1(_0663_),
    .S(_0744_),
    .X(_0817_));
 sg13g2_nor4_2 _1616_ (.A(_0809_),
    .B(net537),
    .C(net530),
    .Y(_0818_),
    .D(net529));
 sg13g2_nand4_1 _1617_ (.B(_0801_),
    .C(_0807_),
    .A(_0800_),
    .Y(_0819_),
    .D(_0808_));
 sg13g2_nor4_2 _1618_ (.A(net536),
    .B(net533),
    .C(net526),
    .Y(_0820_),
    .D(_0819_));
 sg13g2_nand2_1 _1619_ (.Y(_0821_),
    .A(\enigma.plugboard.bits_6_1.q ),
    .B(_0820_));
 sg13g2_nor4_2 _1620_ (.A(net537),
    .B(net530),
    .C(net527),
    .Y(_0822_),
    .D(_0819_));
 sg13g2_nor4_2 _1621_ (.A(net536),
    .B(net533),
    .C(net528),
    .Y(_0823_),
    .D(_0819_));
 sg13g2_nand4_1 _1622_ (.B(_0803_),
    .C(_0807_),
    .A(_0802_),
    .Y(_0824_),
    .D(_0808_));
 sg13g2_nor4_2 _1623_ (.A(net536),
    .B(net533),
    .C(net528),
    .Y(_0825_),
    .D(_0824_));
 sg13g2_nor4_2 _1624_ (.A(net534),
    .B(net533),
    .C(net526),
    .Y(_0826_),
    .D(_0824_));
 sg13g2_nor4_2 _1625_ (.A(net534),
    .B(net532),
    .C(net528),
    .Y(_0827_),
    .D(_0819_));
 sg13g2_a22oi_1 _1626_ (.Y(_0828_),
    .B1(_0807_),
    .B2(_0808_),
    .A2(_0803_),
    .A1(_0802_));
 sg13g2_and4_2 _1627_ (.A(net536),
    .B(net530),
    .C(net528),
    .D(_0828_),
    .X(_0829_));
 sg13g2_nor4_2 _1628_ (.A(_0809_),
    .B(net536),
    .C(net532),
    .Y(_0830_),
    .D(net526));
 sg13g2_nor4_2 _1629_ (.A(net537),
    .B(net531),
    .C(net529),
    .Y(_0831_),
    .D(_0819_));
 sg13g2_nor4_2 _1630_ (.A(net535),
    .B(net533),
    .C(net529),
    .Y(_0832_),
    .D(_0824_));
 sg13g2_and4_2 _1631_ (.A(net535),
    .B(net532),
    .C(net527),
    .D(_0828_),
    .X(_0833_));
 sg13g2_nor4_2 _1632_ (.A(_0809_),
    .B(net536),
    .C(net533),
    .Y(_0834_),
    .D(net528));
 sg13g2_and4_2 _1633_ (.A(net535),
    .B(net532),
    .C(net529),
    .D(_0828_),
    .X(_0835_));
 sg13g2_and4_2 _1634_ (.A(net534),
    .B(net530),
    .C(net528),
    .D(_0828_),
    .X(_0836_));
 sg13g2_nor4_2 _1635_ (.A(net535),
    .B(net531),
    .C(net529),
    .Y(_0837_),
    .D(_0824_));
 sg13g2_nor4_2 _1636_ (.A(net534),
    .B(net532),
    .C(net526),
    .Y(_0838_),
    .D(_0819_));
 sg13g2_and4_2 _1637_ (.A(net534),
    .B(net530),
    .C(net526),
    .D(_0828_),
    .X(_0839_));
 sg13g2_nor4_2 _1638_ (.A(_0809_),
    .B(net534),
    .C(net532),
    .Y(_0840_),
    .D(net526));
 sg13g2_nor4_2 _1639_ (.A(_0809_),
    .B(net535),
    .C(net531),
    .Y(_0841_),
    .D(net529));
 sg13g2_nor4_2 _1640_ (.A(net536),
    .B(net530),
    .C(net526),
    .Y(_0842_),
    .D(_0824_));
 sg13g2_nor4_2 _1641_ (.A(_0809_),
    .B(net534),
    .C(net532),
    .Y(_0843_),
    .D(net528));
 sg13g2_nor4_2 _1642_ (.A(net537),
    .B(net532),
    .C(net527),
    .Y(_0844_),
    .D(_0824_));
 sg13g2_and4_2 _1643_ (.A(net536),
    .B(net530),
    .C(net526),
    .D(_0828_),
    .X(_0845_));
 sg13g2_nor4_2 _1644_ (.A(_0809_),
    .B(net537),
    .C(net531),
    .Y(_0846_),
    .D(net527));
 sg13g2_nor4_2 _1645_ (.A(net537),
    .B(net530),
    .C(net528),
    .Y(_0847_),
    .D(_0824_));
 sg13g2_a22oi_1 _1646_ (.Y(_0848_),
    .B1(_0829_),
    .B2(\enigma.plugboard.bits_15_1.q ),
    .A2(_0822_),
    .A1(\enigma.plugboard.bits_22_1.q ));
 sg13g2_a22oi_1 _1647_ (.Y(_0849_),
    .B1(_0846_),
    .B2(\enigma.plugboard.bits_21_1.q ),
    .A2(_0823_),
    .A1(\enigma.plugboard.bits_2_1.q ));
 sg13g2_a22oi_1 _1648_ (.Y(_0850_),
    .B1(_0845_),
    .B2(\enigma.plugboard.bits_11_1.q ),
    .A2(_0840_),
    .A1(\enigma.plugboard.bits_13_1.q ));
 sg13g2_a22oi_1 _1649_ (.Y(_0851_),
    .B1(_0837_),
    .B2(\enigma.plugboard.bits_24_1.q ),
    .A2(_0831_),
    .A1(\enigma.plugboard.bits_18_1.q ));
 sg13g2_a22oi_1 _1650_ (.Y(_0852_),
    .B1(_0844_),
    .B2(\enigma.plugboard.bits_4_1.q ),
    .A2(_0835_),
    .A1(\enigma.plugboard.bits_23_1.q ));
 sg13g2_nand3_1 _1651_ (.B(_0849_),
    .C(_0852_),
    .A(_0848_),
    .Y(_0853_));
 sg13g2_a221oi_1 _1652_ (.B2(\enigma.plugboard.bits_8_1.q ),
    .C1(_0853_),
    .B1(_0832_),
    .A1(\enigma.plugboard.bits_17_1.q ),
    .Y(_0854_),
    .A2(_0818_));
 sg13g2_a21oi_1 _1653_ (.A1(\enigma.plugboard.bits_14_1.q ),
    .A2(_0838_),
    .Y(_0855_),
    .B1(net538));
 sg13g2_a22oi_1 _1654_ (.Y(_0856_),
    .B1(_0833_),
    .B2(\enigma.plugboard.bits_19_1.q ),
    .A2(_0826_),
    .A1(\enigma.plugboard.bits_12_1.q ));
 sg13g2_a22oi_1 _1655_ (.Y(_0857_),
    .B1(_0847_),
    .B2(\enigma.plugboard.bits_16_1.q ),
    .A2(_0842_),
    .A1(\enigma.plugboard.bits_20_1.q ));
 sg13g2_nand4_1 _1656_ (.B(_0855_),
    .C(_0856_),
    .A(_0850_),
    .Y(_0858_),
    .D(_0857_));
 sg13g2_a22oi_1 _1657_ (.Y(_0859_),
    .B1(_0839_),
    .B2(\enigma.plugboard.bits_3_1.q ),
    .A2(_0827_),
    .A1(\enigma.plugboard.bits_10_1.q ));
 sg13g2_a22oi_1 _1658_ (.Y(_0860_),
    .B1(_0836_),
    .B2(\enigma.plugboard.bits_7_1.q ),
    .A2(_0830_),
    .A1(\enigma.plugboard.bits_5_1.q ));
 sg13g2_a22oi_1 _1659_ (.Y(_0861_),
    .B1(_0841_),
    .B2(\enigma.plugboard.bits_25_1.q ),
    .A2(_0834_),
    .A1(\enigma.plugboard.bits_1_1.q ));
 sg13g2_a22oi_1 _1660_ (.Y(_0862_),
    .B1(_0843_),
    .B2(\enigma.plugboard.bits_9_1.q ),
    .A2(_0825_),
    .A1(\enigma.plugboard.bits_0_1.q ));
 sg13g2_nand4_1 _1661_ (.B(_0860_),
    .C(_0861_),
    .A(_0859_),
    .Y(_0863_),
    .D(_0862_));
 sg13g2_nor2_1 _1662_ (.A(_0858_),
    .B(_0863_),
    .Y(_0864_));
 sg13g2_nand4_1 _1663_ (.B(_0851_),
    .C(_0854_),
    .A(_0821_),
    .Y(_0865_),
    .D(_0864_));
 sg13g2_and2_1 _1664_ (.A(_0804_),
    .B(_0865_),
    .X(_0866_));
 sg13g2_nor2_1 _1665_ (.A(net584),
    .B(net583),
    .Y(_0867_));
 sg13g2_a21oi_1 _1666_ (.A1(net585),
    .A2(net583),
    .Y(_0868_),
    .B1(net582));
 sg13g2_nand2_2 _1667_ (.Y(_0869_),
    .A(_0663_),
    .B(net584));
 sg13g2_o21ai_1 _1668_ (.B1(net581),
    .Y(_0870_),
    .A1(net583),
    .A2(_0869_));
 sg13g2_nor2_1 _1669_ (.A(_0663_),
    .B(net583),
    .Y(_0871_));
 sg13g2_nor3_1 _1670_ (.A(\enigma.r.dout[3] ),
    .B(_0867_),
    .C(_0868_),
    .Y(_0872_));
 sg13g2_nor2_1 _1671_ (.A(\enigma.r.dout[4] ),
    .B(_0665_),
    .Y(_0873_));
 sg13g2_a22oi_1 _1672_ (.Y(_0874_),
    .B1(_0869_),
    .B2(_0873_),
    .A2(_0666_),
    .A1(_0664_));
 sg13g2_o21ai_1 _1673_ (.B1(_0870_),
    .Y(_0875_),
    .A1(\enigma.r.dout[3] ),
    .A2(_0871_));
 sg13g2_o21ai_1 _1674_ (.B1(_0793_),
    .Y(_0876_),
    .A1(_0872_),
    .A2(_0874_));
 sg13g2_a21oi_1 _1675_ (.A1(net580),
    .A2(_0875_),
    .Y(_0877_),
    .B1(_0876_));
 sg13g2_a221oi_1 _1676_ (.B2(_0866_),
    .C1(_0877_),
    .B1(_0796_),
    .A1(net583),
    .Y(_0878_),
    .A2(_0795_));
 sg13g2_inv_1 _1677_ (.Y(_0879_),
    .A(_0878_));
 sg13g2_a221oi_1 _1678_ (.B2(net539),
    .C1(_0658_),
    .B1(net540),
    .A1(net542),
    .Y(_0880_),
    .A2(net541));
 sg13g2_a221oi_1 _1679_ (.B2(\enigma.r.cnts_debug0[1] ),
    .C1(_0880_),
    .B1(net521),
    .A1(\enigma.r.cnts_debug1[1] ),
    .Y(_0881_),
    .A2(net523));
 sg13g2_a221oi_1 _1680_ (.B2(net539),
    .C1(_0661_),
    .B1(net540),
    .A1(net542),
    .Y(_0882_),
    .A2(net541));
 sg13g2_a221oi_1 _1681_ (.B2(\enigma.r.$signal$13[1] ),
    .C1(_0882_),
    .B1(net521),
    .A1(\enigma.r.$signal$20[1] ),
    .Y(_0883_),
    .A2(net523));
 sg13g2_nand2b_1 _1682_ (.Y(_0884_),
    .B(_0883_),
    .A_N(_0881_));
 sg13g2_nand2b_1 _1683_ (.Y(_0885_),
    .B(_0881_),
    .A_N(_0883_));
 sg13g2_xor2_1 _1684_ (.B(_0883_),
    .A(_0881_),
    .X(_0886_));
 sg13g2_nand2_1 _1685_ (.Y(_0887_),
    .A(_0786_),
    .B(_0886_));
 sg13g2_xnor2_1 _1686_ (.Y(_0888_),
    .A(_0786_),
    .B(_0886_));
 sg13g2_a22oi_1 _1687_ (.Y(_0889_),
    .B1(net522),
    .B2(\enigma.r.cnts_debug0[4] ),
    .A2(net525),
    .A1(\enigma.r.cnts_debug2[4] ));
 sg13g2_o21ai_1 _1688_ (.B1(_0889_),
    .Y(_0890_),
    .A1(_0655_),
    .A2(_0778_));
 sg13g2_nand2_1 _1689_ (.Y(_0891_),
    .A(\enigma.r.$signal$22[4] ),
    .B(net525));
 sg13g2_a22oi_1 _1690_ (.Y(_0892_),
    .B1(net521),
    .B2(\enigma.r.$signal$13[4] ),
    .A2(net524),
    .A1(\enigma.r.$signal$20[4] ));
 sg13g2_and3_1 _1691_ (.X(_0893_),
    .A(_0890_),
    .B(_0891_),
    .C(_0892_));
 sg13g2_nand3_1 _1692_ (.B(_0891_),
    .C(_0892_),
    .A(_0890_),
    .Y(_0894_));
 sg13g2_a21oi_1 _1693_ (.A1(_0891_),
    .A2(_0892_),
    .Y(_0895_),
    .B1(_0890_));
 sg13g2_and2_1 _1694_ (.A(\enigma.r.$signal$13[3] ),
    .B(net521),
    .X(_0896_));
 sg13g2_a221oi_1 _1695_ (.B2(\enigma.r.$signal$20[3] ),
    .C1(_0896_),
    .B1(net523),
    .A1(\enigma.r.$signal$22[3] ),
    .Y(_0897_),
    .A2(net525));
 sg13g2_nand2_1 _1696_ (.Y(_0898_),
    .A(\enigma.r.cnts_debug1[3] ),
    .B(net523));
 sg13g2_a22oi_1 _1697_ (.Y(_0899_),
    .B1(net522),
    .B2(\enigma.r.cnts_debug0[3] ),
    .A2(_0775_),
    .A1(\enigma.r.cnts_debug2[3] ));
 sg13g2_and2_1 _1698_ (.A(_0898_),
    .B(_0899_),
    .X(_0900_));
 sg13g2_nand2_2 _1699_ (.Y(_0901_),
    .A(_0898_),
    .B(_0899_));
 sg13g2_nor2_2 _1700_ (.A(_0897_),
    .B(_0901_),
    .Y(_0902_));
 sg13g2_a221oi_1 _1701_ (.B2(net539),
    .C1(_0657_),
    .B1(net540),
    .A1(net542),
    .Y(_0903_),
    .A2(net541));
 sg13g2_a221oi_1 _1702_ (.B2(\enigma.r.cnts_debug0[2] ),
    .C1(_0903_),
    .B1(net522),
    .A1(\enigma.r.cnts_debug1[2] ),
    .Y(_0904_),
    .A2(net523));
 sg13g2_a221oi_1 _1703_ (.B2(net539),
    .C1(_0660_),
    .B1(net540),
    .A1(net542),
    .Y(_0905_),
    .A2(net541));
 sg13g2_a221oi_1 _1704_ (.B2(\enigma.r.$signal$13[2] ),
    .C1(_0905_),
    .B1(net521),
    .A1(\enigma.r.$signal$20[2] ),
    .Y(_0906_),
    .A2(net523));
 sg13g2_nor2b_1 _1705_ (.A(_0904_),
    .B_N(_0906_),
    .Y(_0907_));
 sg13g2_xnor2_1 _1706_ (.Y(_0908_),
    .A(_0904_),
    .B(_0906_));
 sg13g2_nand2b_1 _1707_ (.Y(_0909_),
    .B(_0884_),
    .A_N(_0786_));
 sg13g2_and2_1 _1708_ (.A(_0885_),
    .B(_0908_),
    .X(_0910_));
 sg13g2_nand2_1 _1709_ (.Y(_0911_),
    .A(_0885_),
    .B(_0908_));
 sg13g2_nand2_1 _1710_ (.Y(_0912_),
    .A(_0909_),
    .B(_0910_));
 sg13g2_a221oi_1 _1711_ (.B2(_0910_),
    .C1(_0907_),
    .B1(_0909_),
    .A1(_0897_),
    .Y(_0913_),
    .A2(_0901_));
 sg13g2_nor2_1 _1712_ (.A(_0902_),
    .B(_0913_),
    .Y(_0914_));
 sg13g2_nor3_1 _1713_ (.A(_0895_),
    .B(_0902_),
    .C(_0913_),
    .Y(_0915_));
 sg13g2_or3_1 _1714_ (.A(_0895_),
    .B(_0902_),
    .C(_0913_),
    .X(_0916_));
 sg13g2_nor2_2 _1715_ (.A(_0893_),
    .B(_0915_),
    .Y(_0917_));
 sg13g2_a21oi_2 _1716_ (.B1(_0888_),
    .Y(_0918_),
    .A2(_0916_),
    .A1(_0894_));
 sg13g2_and3_1 _1717_ (.X(_0919_),
    .A(_0888_),
    .B(_0894_),
    .C(_0916_));
 sg13g2_or2_2 _1718_ (.X(_0920_),
    .B(_0919_),
    .A(_0918_));
 sg13g2_nor3_1 _1719_ (.A(net513),
    .B(_0918_),
    .C(_0919_),
    .Y(_0921_));
 sg13g2_nand3_1 _1720_ (.B(_0807_),
    .C(_0808_),
    .A(_0799_),
    .Y(_0922_));
 sg13g2_nand2_1 _1721_ (.Y(_0923_),
    .A(\enigma.plugboard.bits_24_0.q ),
    .B(_0837_));
 sg13g2_a22oi_1 _1722_ (.Y(_0924_),
    .B1(_0838_),
    .B2(\enigma.plugboard.bits_14_0.q ),
    .A2(_0832_),
    .A1(\enigma.plugboard.bits_8_0.q ));
 sg13g2_a22oi_1 _1723_ (.Y(_0925_),
    .B1(_0835_),
    .B2(\enigma.plugboard.bits_23_0.q ),
    .A2(_0831_),
    .A1(\enigma.plugboard.bits_18_0.q ));
 sg13g2_a22oi_1 _1724_ (.Y(_0926_),
    .B1(_0829_),
    .B2(\enigma.plugboard.bits_15_0.q ),
    .A2(_0825_),
    .A1(\enigma.plugboard.bits_0_0.q ));
 sg13g2_a22oi_1 _1725_ (.Y(_0927_),
    .B1(_0846_),
    .B2(\enigma.plugboard.bits_21_0.q ),
    .A2(_0843_),
    .A1(\enigma.plugboard.bits_9_0.q ));
 sg13g2_a22oi_1 _1726_ (.Y(_0928_),
    .B1(_0842_),
    .B2(\enigma.plugboard.bits_20_0.q ),
    .A2(_0839_),
    .A1(\enigma.plugboard.bits_3_0.q ));
 sg13g2_nand3_1 _1727_ (.B(_0926_),
    .C(_0928_),
    .A(_0925_),
    .Y(_0929_));
 sg13g2_a221oi_1 _1728_ (.B2(\enigma.plugboard.bits_1_0.q ),
    .C1(_0929_),
    .B1(_0834_),
    .A1(\enigma.plugboard.bits_12_0.q ),
    .Y(_0930_),
    .A2(_0826_));
 sg13g2_a21oi_1 _1729_ (.A1(\enigma.plugboard.bits_11_0.q ),
    .A2(_0845_),
    .Y(_0931_),
    .B1(net538));
 sg13g2_a22oi_1 _1730_ (.Y(_0932_),
    .B1(_0840_),
    .B2(\enigma.plugboard.bits_13_0.q ),
    .A2(_0833_),
    .A1(\enigma.plugboard.bits_19_0.q ));
 sg13g2_a22oi_1 _1731_ (.Y(_0933_),
    .B1(_0841_),
    .B2(\enigma.plugboard.bits_25_0.q ),
    .A2(_0823_),
    .A1(\enigma.plugboard.bits_2_0.q ));
 sg13g2_nand4_1 _1732_ (.B(_0931_),
    .C(_0932_),
    .A(_0924_),
    .Y(_0934_),
    .D(_0933_));
 sg13g2_a22oi_1 _1733_ (.Y(_0935_),
    .B1(_0836_),
    .B2(\enigma.plugboard.bits_7_0.q ),
    .A2(_0818_),
    .A1(\enigma.plugboard.bits_17_0.q ));
 sg13g2_a22oi_1 _1734_ (.Y(_0936_),
    .B1(_0847_),
    .B2(\enigma.plugboard.bits_16_0.q ),
    .A2(_0830_),
    .A1(\enigma.plugboard.bits_5_0.q ));
 sg13g2_a22oi_1 _1735_ (.Y(_0937_),
    .B1(_0827_),
    .B2(\enigma.plugboard.bits_10_0.q ),
    .A2(_0820_),
    .A1(\enigma.plugboard.bits_6_0.q ));
 sg13g2_a22oi_1 _1736_ (.Y(_0938_),
    .B1(_0844_),
    .B2(\enigma.plugboard.bits_4_0.q ),
    .A2(_0822_),
    .A1(\enigma.plugboard.bits_22_0.q ));
 sg13g2_nand4_1 _1737_ (.B(_0936_),
    .C(_0937_),
    .A(_0935_),
    .Y(_0939_),
    .D(_0938_));
 sg13g2_nor2_1 _1738_ (.A(_0934_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_nand4_1 _1739_ (.B(_0927_),
    .C(_0930_),
    .A(_0923_),
    .Y(_0941_),
    .D(_0940_));
 sg13g2_and2_1 _1740_ (.A(_0922_),
    .B(_0941_),
    .X(_0942_));
 sg13g2_and2_1 _1741_ (.A(net582),
    .B(_0012_),
    .X(_0943_));
 sg13g2_a21oi_1 _1742_ (.A1(_0663_),
    .A2(_0867_),
    .Y(_0944_),
    .B1(_0943_));
 sg13g2_nand2_1 _1743_ (.Y(_0945_),
    .A(_0870_),
    .B(_0944_));
 sg13g2_nand2_1 _1744_ (.Y(_0946_),
    .A(_0663_),
    .B(_0011_));
 sg13g2_nor2_1 _1745_ (.A(net581),
    .B(_0943_),
    .Y(_0947_));
 sg13g2_a221oi_1 _1746_ (.B2(_0947_),
    .C1(net580),
    .B1(_0946_),
    .A1(net581),
    .Y(_0948_),
    .A2(_0868_));
 sg13g2_a21oi_1 _1747_ (.A1(net580),
    .A2(_0945_),
    .Y(_0949_),
    .B1(_0948_));
 sg13g2_and2_1 _1748_ (.A(net584),
    .B(_0795_),
    .X(_0950_));
 sg13g2_a221oi_1 _1749_ (.B2(_0793_),
    .C1(_0950_),
    .B1(_0949_),
    .A1(_0796_),
    .Y(_0951_),
    .A2(_0942_));
 sg13g2_nor2_1 _1750_ (.A(_0788_),
    .B(net512),
    .Y(_0952_));
 sg13g2_o21ai_1 _1751_ (.B1(net513),
    .Y(_0953_),
    .A1(_0918_),
    .A2(_0919_));
 sg13g2_nor2b_1 _1752_ (.A(_0921_),
    .B_N(_0953_),
    .Y(_0954_));
 sg13g2_a21oi_1 _1753_ (.A1(_0952_),
    .A2(_0953_),
    .Y(_0955_),
    .B1(_0921_));
 sg13g2_a21o_1 _1754_ (.A2(_0953_),
    .A1(_0952_),
    .B1(_0921_),
    .X(_0956_));
 sg13g2_nand2_1 _1755_ (.Y(_0957_),
    .A(\enigma.plugboard.bits_4_2.q ),
    .B(_0844_));
 sg13g2_a22oi_1 _1756_ (.Y(_0958_),
    .B1(_0839_),
    .B2(\enigma.plugboard.bits_3_2.q ),
    .A2(_0820_),
    .A1(\enigma.plugboard.bits_6_2.q ));
 sg13g2_a22oi_1 _1757_ (.Y(_0959_),
    .B1(_0833_),
    .B2(\enigma.plugboard.bits_19_2.q ),
    .A2(_0831_),
    .A1(\enigma.plugboard.bits_18_2.q ));
 sg13g2_a22oi_1 _1758_ (.Y(_0960_),
    .B1(_0846_),
    .B2(\enigma.plugboard.bits_21_2.q ),
    .A2(_0837_),
    .A1(\enigma.plugboard.bits_24_2.q ));
 sg13g2_a22oi_1 _1759_ (.Y(_0961_),
    .B1(_0843_),
    .B2(\enigma.plugboard.bits_9_2.q ),
    .A2(_0830_),
    .A1(\enigma.plugboard.bits_5_2.q ));
 sg13g2_a22oi_1 _1760_ (.Y(_0962_),
    .B1(_0841_),
    .B2(\enigma.plugboard.bits_25_2.q ),
    .A2(_0832_),
    .A1(\enigma.plugboard.bits_8_2.q ));
 sg13g2_nand2_1 _1761_ (.Y(_0963_),
    .A(_0957_),
    .B(_0962_));
 sg13g2_a22oi_1 _1762_ (.Y(_0964_),
    .B1(_0834_),
    .B2(\enigma.plugboard.bits_1_2.q ),
    .A2(_0823_),
    .A1(\enigma.plugboard.bits_2_2.q ));
 sg13g2_nand4_1 _1763_ (.B(_0960_),
    .C(_0961_),
    .A(_0959_),
    .Y(_0965_),
    .D(_0964_));
 sg13g2_nor2_1 _1764_ (.A(_0963_),
    .B(_0965_),
    .Y(_0966_));
 sg13g2_a21oi_1 _1765_ (.A1(\enigma.plugboard.bits_0_2.q ),
    .A2(_0825_),
    .Y(_0967_),
    .B1(net538));
 sg13g2_a22oi_1 _1766_ (.Y(_0968_),
    .B1(_0840_),
    .B2(\enigma.plugboard.bits_13_2.q ),
    .A2(_0836_),
    .A1(\enigma.plugboard.bits_7_2.q ));
 sg13g2_a22oi_1 _1767_ (.Y(_0969_),
    .B1(_0835_),
    .B2(\enigma.plugboard.bits_23_2.q ),
    .A2(_0822_),
    .A1(\enigma.plugboard.bits_22_2.q ));
 sg13g2_nand4_1 _1768_ (.B(_0967_),
    .C(_0968_),
    .A(_0958_),
    .Y(_0970_),
    .D(_0969_));
 sg13g2_a22oi_1 _1769_ (.Y(_0971_),
    .B1(_0829_),
    .B2(\enigma.plugboard.bits_15_2.q ),
    .A2(_0818_),
    .A1(\enigma.plugboard.bits_17_2.q ));
 sg13g2_a22oi_1 _1770_ (.Y(_0972_),
    .B1(_0845_),
    .B2(\enigma.plugboard.bits_11_2.q ),
    .A2(_0842_),
    .A1(\enigma.plugboard.bits_20_2.q ));
 sg13g2_a22oi_1 _1771_ (.Y(_0973_),
    .B1(_0827_),
    .B2(\enigma.plugboard.bits_10_2.q ),
    .A2(_0826_),
    .A1(\enigma.plugboard.bits_12_2.q ));
 sg13g2_a22oi_1 _1772_ (.Y(_0974_),
    .B1(_0847_),
    .B2(\enigma.plugboard.bits_16_2.q ),
    .A2(_0838_),
    .A1(\enigma.plugboard.bits_14_2.q ));
 sg13g2_nand4_1 _1773_ (.B(_0972_),
    .C(_0973_),
    .A(_0971_),
    .Y(_0975_),
    .D(_0974_));
 sg13g2_nor2_2 _1774_ (.A(_0970_),
    .B(_0975_),
    .Y(_0976_));
 sg13g2_a22oi_1 _1775_ (.Y(_0977_),
    .B1(_0966_),
    .B2(_0976_),
    .A2(net527),
    .A1(net538));
 sg13g2_nand2_1 _1776_ (.Y(_0978_),
    .A(_0796_),
    .B(_0977_));
 sg13g2_nand2_1 _1777_ (.Y(_0979_),
    .A(_0663_),
    .B(net583));
 sg13g2_a221oi_1 _1778_ (.B2(_0979_),
    .C1(net580),
    .B1(_0666_),
    .A1(net582),
    .Y(_0980_),
    .A2(net584));
 sg13g2_xnor2_1 _1779_ (.Y(_0981_),
    .A(net584),
    .B(net583));
 sg13g2_nor2b_1 _1780_ (.A(net581),
    .B_N(net580),
    .Y(_0982_));
 sg13g2_nand2_1 _1781_ (.Y(_0983_),
    .A(_0869_),
    .B(_0982_));
 sg13g2_a21oi_1 _1782_ (.A1(net582),
    .A2(_0981_),
    .Y(_0984_),
    .B1(_0983_));
 sg13g2_o21ai_1 _1783_ (.B1(_0793_),
    .Y(_0985_),
    .A1(_0980_),
    .A2(_0984_));
 sg13g2_nand2_1 _1784_ (.Y(_0986_),
    .A(net582),
    .B(_0795_));
 sg13g2_and3_2 _1785_ (.X(_0987_),
    .A(_0978_),
    .B(_0985_),
    .C(_0986_));
 sg13g2_nand3_1 _1786_ (.B(_0985_),
    .C(_0986_),
    .A(_0978_),
    .Y(_0988_));
 sg13g2_a21o_1 _1787_ (.A2(_0909_),
    .A1(_0885_),
    .B1(_0908_),
    .X(_0989_));
 sg13g2_nand2_1 _1788_ (.Y(_0990_),
    .A(_0912_),
    .B(_0989_));
 sg13g2_nor2_1 _1789_ (.A(_0885_),
    .B(_0908_),
    .Y(_0991_));
 sg13g2_or2_1 _1790_ (.X(_0992_),
    .B(_0991_),
    .A(_0910_));
 sg13g2_xnor2_1 _1791_ (.Y(_0993_),
    .A(_0887_),
    .B(_0992_));
 sg13g2_o21ai_1 _1792_ (.B1(_0990_),
    .Y(_0994_),
    .A1(_0893_),
    .A2(_0915_));
 sg13g2_nand3_1 _1793_ (.B(_0916_),
    .C(_0993_),
    .A(_0894_),
    .Y(_0995_));
 sg13g2_and2_1 _1794_ (.A(_0994_),
    .B(_0995_),
    .X(_0996_));
 sg13g2_nand3_1 _1795_ (.B(_0994_),
    .C(_0995_),
    .A(_0988_),
    .Y(_0997_));
 sg13g2_nor2_1 _1796_ (.A(_0988_),
    .B(_0996_),
    .Y(_0998_));
 sg13g2_xnor2_1 _1797_ (.Y(_0999_),
    .A(_0987_),
    .B(_0996_));
 sg13g2_xnor2_1 _1798_ (.Y(_1000_),
    .A(_0955_),
    .B(_0999_));
 sg13g2_xnor2_1 _1799_ (.Y(_1001_),
    .A(_0956_),
    .B(_0999_));
 sg13g2_xnor2_1 _1800_ (.Y(_1002_),
    .A(_0952_),
    .B(_0954_));
 sg13g2_inv_1 _1801_ (.Y(_1003_),
    .A(_1002_));
 sg13g2_nand2_2 _1802_ (.Y(_1004_),
    .A(_1001_),
    .B(_1002_));
 sg13g2_nand2_1 _1803_ (.Y(_1005_),
    .A(\enigma.plugboard.bits_22_3.q ),
    .B(_0822_));
 sg13g2_a22oi_1 _1804_ (.Y(_1006_),
    .B1(_0842_),
    .B2(\enigma.plugboard.bits_20_3.q ),
    .A2(_0839_),
    .A1(\enigma.plugboard.bits_3_3.q ));
 sg13g2_a22oi_1 _1805_ (.Y(_1007_),
    .B1(_0845_),
    .B2(\enigma.plugboard.bits_11_3.q ),
    .A2(_0825_),
    .A1(\enigma.plugboard.bits_0_3.q ));
 sg13g2_a22oi_1 _1806_ (.Y(_1008_),
    .B1(_0846_),
    .B2(\enigma.plugboard.bits_21_3.q ),
    .A2(_0826_),
    .A1(\enigma.plugboard.bits_12_3.q ));
 sg13g2_a22oi_1 _1807_ (.Y(_1009_),
    .B1(_0838_),
    .B2(\enigma.plugboard.bits_14_3.q ),
    .A2(_0823_),
    .A1(\enigma.plugboard.bits_2_3.q ));
 sg13g2_a22oi_1 _1808_ (.Y(_1010_),
    .B1(_0841_),
    .B2(\enigma.plugboard.bits_25_3.q ),
    .A2(_0818_),
    .A1(\enigma.plugboard.bits_17_3.q ));
 sg13g2_a22oi_1 _1809_ (.Y(_1011_),
    .B1(_0834_),
    .B2(\enigma.plugboard.bits_1_3.q ),
    .A2(_0820_),
    .A1(\enigma.plugboard.bits_6_3.q ));
 sg13g2_nand4_1 _1810_ (.B(_1008_),
    .C(_1009_),
    .A(_1007_),
    .Y(_1012_),
    .D(_1011_));
 sg13g2_nand3b_1 _1811_ (.B(_1005_),
    .C(_1010_),
    .Y(_1013_),
    .A_N(_1012_));
 sg13g2_a21oi_1 _1812_ (.A1(\enigma.plugboard.bits_24_3.q ),
    .A2(_0837_),
    .Y(_1014_),
    .B1(net538));
 sg13g2_a22oi_1 _1813_ (.Y(_1015_),
    .B1(_0847_),
    .B2(\enigma.plugboard.bits_16_3.q ),
    .A2(_0844_),
    .A1(\enigma.plugboard.bits_4_3.q ));
 sg13g2_a22oi_1 _1814_ (.Y(_1016_),
    .B1(_0835_),
    .B2(\enigma.plugboard.bits_23_3.q ),
    .A2(_0833_),
    .A1(\enigma.plugboard.bits_19_3.q ));
 sg13g2_nand4_1 _1815_ (.B(_1014_),
    .C(_1015_),
    .A(_1006_),
    .Y(_1017_),
    .D(_1016_));
 sg13g2_a22oi_1 _1816_ (.Y(_1018_),
    .B1(_0840_),
    .B2(\enigma.plugboard.bits_13_3.q ),
    .A2(_0827_),
    .A1(\enigma.plugboard.bits_10_3.q ));
 sg13g2_a22oi_1 _1817_ (.Y(_1019_),
    .B1(_0843_),
    .B2(\enigma.plugboard.bits_9_3.q ),
    .A2(_0829_),
    .A1(\enigma.plugboard.bits_15_3.q ));
 sg13g2_a22oi_1 _1818_ (.Y(_1020_),
    .B1(_0832_),
    .B2(\enigma.plugboard.bits_8_3.q ),
    .A2(_0831_),
    .A1(\enigma.plugboard.bits_18_3.q ));
 sg13g2_a22oi_1 _1819_ (.Y(_1021_),
    .B1(_0836_),
    .B2(\enigma.plugboard.bits_7_3.q ),
    .A2(_0830_),
    .A1(\enigma.plugboard.bits_5_3.q ));
 sg13g2_nand4_1 _1820_ (.B(_1019_),
    .C(_1020_),
    .A(_1018_),
    .Y(_1022_),
    .D(_1021_));
 sg13g2_nor3_2 _1821_ (.A(_1013_),
    .B(_1017_),
    .C(_1022_),
    .Y(_1023_));
 sg13g2_a21oi_2 _1822_ (.B1(_1023_),
    .Y(_1024_),
    .A2(net534),
    .A1(net538));
 sg13g2_nand2_1 _1823_ (.Y(_1025_),
    .A(_0796_),
    .B(_1024_));
 sg13g2_nand3_1 _1824_ (.B(net583),
    .C(_0982_),
    .A(net584),
    .Y(_1026_));
 sg13g2_nor2_1 _1825_ (.A(net584),
    .B(_0871_),
    .Y(_1027_));
 sg13g2_a22oi_1 _1826_ (.Y(_1028_),
    .B1(_0979_),
    .B2(_1027_),
    .A2(_0869_),
    .A1(net581));
 sg13g2_o21ai_1 _1827_ (.B1(_1026_),
    .Y(_1029_),
    .A1(net580),
    .A2(_1028_));
 sg13g2_nand2_1 _1828_ (.Y(_1030_),
    .A(_0793_),
    .B(_1029_));
 sg13g2_nand2_1 _1829_ (.Y(_1031_),
    .A(net581),
    .B(_0795_));
 sg13g2_and3_2 _1830_ (.X(_1032_),
    .A(_1025_),
    .B(_1030_),
    .C(_1031_));
 sg13g2_nand3_1 _1831_ (.B(_1030_),
    .C(_1031_),
    .A(_1025_),
    .Y(_1033_));
 sg13g2_xnor2_1 _1832_ (.Y(_1034_),
    .A(_0897_),
    .B(_0900_));
 sg13g2_nor2b_1 _1833_ (.A(_1034_),
    .B_N(_0907_),
    .Y(_1035_));
 sg13g2_xnor2_1 _1834_ (.Y(_1036_),
    .A(_0907_),
    .B(_1034_));
 sg13g2_mux2_1 _1835_ (.A0(_1034_),
    .A1(_1036_),
    .S(_0912_),
    .X(_1037_));
 sg13g2_nor2b_1 _1836_ (.A(_0917_),
    .B_N(_1037_),
    .Y(_1038_));
 sg13g2_o21ai_1 _1837_ (.B1(_0911_),
    .Y(_1039_),
    .A1(_0887_),
    .A2(_0991_));
 sg13g2_xnor2_1 _1838_ (.Y(_1040_),
    .A(_1036_),
    .B(_1039_));
 sg13g2_a21oi_2 _1839_ (.B1(_1038_),
    .Y(_1041_),
    .A2(_1040_),
    .A1(_0917_));
 sg13g2_mux2_1 _1840_ (.A0(_1037_),
    .A1(_1040_),
    .S(_0917_),
    .X(_1042_));
 sg13g2_nand2_1 _1841_ (.Y(_1043_),
    .A(_1032_),
    .B(_1042_));
 sg13g2_inv_1 _1842_ (.Y(_1044_),
    .A(_1043_));
 sg13g2_xnor2_1 _1843_ (.Y(_1045_),
    .A(_1033_),
    .B(_1041_));
 sg13g2_o21ai_1 _1844_ (.B1(_0997_),
    .Y(_1046_),
    .A1(_0955_),
    .A2(_0998_));
 sg13g2_xnor2_1 _1845_ (.Y(_1047_),
    .A(_1045_),
    .B(_1046_));
 sg13g2_xor2_1 _1846_ (.B(_1046_),
    .A(_1045_),
    .X(_1048_));
 sg13g2_and2_1 _1847_ (.A(_1004_),
    .B(_1047_),
    .X(_1049_));
 sg13g2_nand2_1 _1848_ (.Y(_1050_),
    .A(_1004_),
    .B(_1047_));
 sg13g2_nand2_1 _1849_ (.Y(_1051_),
    .A(\enigma.plugboard.bits_7_4.q ),
    .B(_0836_));
 sg13g2_a22oi_1 _1850_ (.Y(_1052_),
    .B1(_0834_),
    .B2(\enigma.plugboard.bits_1_4.q ),
    .A2(_0825_),
    .A1(\enigma.plugboard.bits_0_4.q ));
 sg13g2_a22oi_1 _1851_ (.Y(_1053_),
    .B1(_0845_),
    .B2(\enigma.plugboard.bits_11_4.q ),
    .A2(_0844_),
    .A1(\enigma.plugboard.bits_4_4.q ));
 sg13g2_a22oi_1 _1852_ (.Y(_1054_),
    .B1(_0839_),
    .B2(\enigma.plugboard.bits_3_4.q ),
    .A2(_0827_),
    .A1(\enigma.plugboard.bits_10_4.q ));
 sg13g2_a22oi_1 _1853_ (.Y(_1055_),
    .B1(_0846_),
    .B2(\enigma.plugboard.bits_21_4.q ),
    .A2(_0835_),
    .A1(\enigma.plugboard.bits_23_4.q ));
 sg13g2_a22oi_1 _1854_ (.Y(_1056_),
    .B1(_0838_),
    .B2(\enigma.plugboard.bits_14_4.q ),
    .A2(_0820_),
    .A1(\enigma.plugboard.bits_6_4.q ));
 sg13g2_a22oi_1 _1855_ (.Y(_1057_),
    .B1(_0843_),
    .B2(\enigma.plugboard.bits_9_4.q ),
    .A2(_0830_),
    .A1(\enigma.plugboard.bits_5_4.q ));
 sg13g2_a22oi_1 _1856_ (.Y(_1058_),
    .B1(_0837_),
    .B2(\enigma.plugboard.bits_24_4.q ),
    .A2(_0832_),
    .A1(\enigma.plugboard.bits_8_4.q ));
 sg13g2_nand3_1 _1857_ (.B(_1056_),
    .C(_1057_),
    .A(_1055_),
    .Y(_1059_));
 sg13g2_a221oi_1 _1858_ (.B2(\enigma.plugboard.bits_16_4.q ),
    .C1(_1059_),
    .B1(_0847_),
    .A1(\enigma.plugboard.bits_13_4.q ),
    .Y(_1060_),
    .A2(_0840_));
 sg13g2_nand3_1 _1859_ (.B(_1058_),
    .C(_1060_),
    .A(_1051_),
    .Y(_1061_));
 sg13g2_a21oi_1 _1860_ (.A1(\enigma.plugboard.bits_22_4.q ),
    .A2(_0822_),
    .Y(_1062_),
    .B1(net538));
 sg13g2_a22oi_1 _1861_ (.Y(_1063_),
    .B1(_0833_),
    .B2(\enigma.plugboard.bits_19_4.q ),
    .A2(_0831_),
    .A1(\enigma.plugboard.bits_18_4.q ));
 sg13g2_nand4_1 _1862_ (.B(_1053_),
    .C(_1062_),
    .A(_1052_),
    .Y(_1064_),
    .D(_1063_));
 sg13g2_a22oi_1 _1863_ (.Y(_1065_),
    .B1(_0842_),
    .B2(\enigma.plugboard.bits_20_4.q ),
    .A2(_0841_),
    .A1(\enigma.plugboard.bits_25_4.q ));
 sg13g2_a22oi_1 _1864_ (.Y(_1066_),
    .B1(_0829_),
    .B2(\enigma.plugboard.bits_15_4.q ),
    .A2(_0818_),
    .A1(\enigma.plugboard.bits_17_4.q ));
 sg13g2_a22oi_1 _1865_ (.Y(_1067_),
    .B1(_0826_),
    .B2(\enigma.plugboard.bits_12_4.q ),
    .A2(_0823_),
    .A1(\enigma.plugboard.bits_2_4.q ));
 sg13g2_nand4_1 _1866_ (.B(_1065_),
    .C(_1066_),
    .A(_1054_),
    .Y(_1068_),
    .D(_1067_));
 sg13g2_nor3_2 _1867_ (.A(_1061_),
    .B(_1064_),
    .C(_1068_),
    .Y(_1069_));
 sg13g2_a21oi_2 _1868_ (.B1(_1069_),
    .Y(_1070_),
    .A2(net531),
    .A1(net538));
 sg13g2_o21ai_1 _1869_ (.B1(_0873_),
    .Y(_1071_),
    .A1(net582),
    .A2(net584));
 sg13g2_a21o_1 _1870_ (.A2(_0981_),
    .A1(net582),
    .B1(_0868_),
    .X(_1072_));
 sg13g2_nand3_1 _1871_ (.B(_0870_),
    .C(_1071_),
    .A(_0793_),
    .Y(_1073_));
 sg13g2_a21oi_1 _1872_ (.A1(_0982_),
    .A2(_1072_),
    .Y(_1074_),
    .B1(_1073_));
 sg13g2_a221oi_1 _1873_ (.B2(_1070_),
    .C1(_1074_),
    .B1(_0796_),
    .A1(net580),
    .Y(_1075_),
    .A2(_0795_));
 sg13g2_inv_1 _1874_ (.Y(_1076_),
    .A(_1075_));
 sg13g2_a21oi_1 _1875_ (.A1(_1036_),
    .A2(_1039_),
    .Y(_1077_),
    .B1(_1035_));
 sg13g2_nor2_1 _1876_ (.A(_0893_),
    .B(_0895_),
    .Y(_1078_));
 sg13g2_xnor2_1 _1877_ (.Y(_1079_),
    .A(_0902_),
    .B(_1078_));
 sg13g2_nor2_1 _1878_ (.A(_1077_),
    .B(_1079_),
    .Y(_1080_));
 sg13g2_nand2_1 _1879_ (.Y(_1081_),
    .A(_1077_),
    .B(_1079_));
 sg13g2_nor2b_1 _1880_ (.A(_1080_),
    .B_N(_0917_),
    .Y(_1082_));
 sg13g2_a22oi_1 _1881_ (.Y(_1083_),
    .B1(_1081_),
    .B2(_1082_),
    .A2(_0914_),
    .A1(_0893_));
 sg13g2_inv_1 _1882_ (.Y(_1084_),
    .A(_1083_));
 sg13g2_nor2_1 _1883_ (.A(_1075_),
    .B(_1083_),
    .Y(_1085_));
 sg13g2_xnor2_1 _1884_ (.Y(_1086_),
    .A(_1075_),
    .B(_1083_));
 sg13g2_o21ai_1 _1885_ (.B1(_0997_),
    .Y(_1087_),
    .A1(_1032_),
    .A2(_1042_));
 sg13g2_a21oi_1 _1886_ (.A1(_0956_),
    .A2(_0999_),
    .Y(_1088_),
    .B1(_1087_));
 sg13g2_or3_2 _1887_ (.A(_1044_),
    .B(_1086_),
    .C(_1088_),
    .X(_1089_));
 sg13g2_o21ai_1 _1888_ (.B1(_1086_),
    .Y(_1090_),
    .A1(_1044_),
    .A2(_1088_));
 sg13g2_and2_1 _1889_ (.A(_1089_),
    .B(_1090_),
    .X(_1091_));
 sg13g2_and4_2 _1890_ (.A(_1004_),
    .B(_1047_),
    .C(_1089_),
    .D(_1090_),
    .X(_1092_));
 sg13g2_nand4_1 _1891_ (.B(_1047_),
    .C(_1089_),
    .A(_1004_),
    .Y(_1093_),
    .D(_1090_));
 sg13g2_nor2b_2 _1892_ (.A(_1085_),
    .B_N(_1089_),
    .Y(_1094_));
 sg13g2_nand2b_2 _1893_ (.Y(_1095_),
    .B(_1089_),
    .A_N(_1085_));
 sg13g2_a21oi_1 _1894_ (.A1(_1093_),
    .A2(_1094_),
    .Y(_1096_),
    .B1(_1050_));
 sg13g2_o21ai_1 _1895_ (.B1(_1049_),
    .Y(_1097_),
    .A1(_1092_),
    .A2(_1095_));
 sg13g2_a21oi_1 _1896_ (.A1(_1049_),
    .A2(_1095_),
    .Y(_1098_),
    .B1(_1091_));
 sg13g2_nand2b_1 _1897_ (.Y(_1099_),
    .B(_1097_),
    .A_N(_1091_));
 sg13g2_nor2_1 _1898_ (.A(_1092_),
    .B(_1098_),
    .Y(_1100_));
 sg13g2_or2_1 _1899_ (.X(_1101_),
    .B(_1098_),
    .A(_1092_));
 sg13g2_o21ai_1 _1900_ (.B1(_1004_),
    .Y(_1102_),
    .A1(_1092_),
    .A2(_1095_));
 sg13g2_nand2_1 _1901_ (.Y(_1103_),
    .A(_1048_),
    .B(_1102_));
 sg13g2_a21oi_1 _1902_ (.A1(_1048_),
    .A2(_1102_),
    .Y(_1104_),
    .B1(_1096_));
 sg13g2_a21o_1 _1903_ (.A2(_1102_),
    .A1(_1048_),
    .B1(_1096_),
    .X(_1105_));
 sg13g2_xnor2_1 _1904_ (.Y(_1106_),
    .A(_0787_),
    .B(net512));
 sg13g2_xnor2_1 _1905_ (.Y(_1107_),
    .A(_0788_),
    .B(net512));
 sg13g2_a21oi_2 _1906_ (.B1(_1003_),
    .Y(_1108_),
    .A2(_1094_),
    .A1(_1093_));
 sg13g2_o21ai_1 _1907_ (.B1(_1002_),
    .Y(_1109_),
    .A1(_1092_),
    .A2(_1095_));
 sg13g2_nor3_2 _1908_ (.A(_1002_),
    .B(_1092_),
    .C(_1095_),
    .Y(_1110_));
 sg13g2_nand3_1 _1909_ (.B(_1093_),
    .C(_1094_),
    .A(_1003_),
    .Y(_1111_));
 sg13g2_nor2_2 _1910_ (.A(_1108_),
    .B(_1110_),
    .Y(_1112_));
 sg13g2_nand2_2 _1911_ (.Y(_1113_),
    .A(_1109_),
    .B(_1111_));
 sg13g2_nor3_1 _1912_ (.A(_1000_),
    .B(_1108_),
    .C(_1110_),
    .Y(_1114_));
 sg13g2_nand2_1 _1913_ (.Y(_1115_),
    .A(_1001_),
    .B(_1112_));
 sg13g2_nor3_2 _1914_ (.A(net505),
    .B(_1108_),
    .C(_1110_),
    .Y(_1116_));
 sg13g2_nand3_1 _1915_ (.B(_1109_),
    .C(_1111_),
    .A(net508),
    .Y(_1117_));
 sg13g2_nand4_1 _1916_ (.B(net508),
    .C(_1109_),
    .A(_1001_),
    .Y(_1118_),
    .D(_1111_));
 sg13g2_a21oi_2 _1917_ (.B1(net496),
    .Y(_1119_),
    .A2(_1118_),
    .A1(net492));
 sg13g2_xnor2_1 _1918_ (.Y(_1120_),
    .A(_1000_),
    .B(_1108_));
 sg13g2_xnor2_1 _1919_ (.Y(_1121_),
    .A(_1001_),
    .B(_1108_));
 sg13g2_a21oi_2 _1920_ (.B1(net509),
    .Y(_1122_),
    .A2(_1111_),
    .A1(_1109_));
 sg13g2_o21ai_1 _1921_ (.B1(net505),
    .Y(_1123_),
    .A1(_1108_),
    .A2(_1110_));
 sg13g2_nor2_1 _1922_ (.A(net476),
    .B(_1122_),
    .Y(_1124_));
 sg13g2_nand2_1 _1923_ (.Y(_1125_),
    .A(net481),
    .B(_1123_));
 sg13g2_nand2_2 _1924_ (.Y(_1126_),
    .A(net505),
    .B(net474));
 sg13g2_a21oi_2 _1925_ (.B1(net494),
    .Y(_1127_),
    .A2(net473),
    .A1(net507));
 sg13g2_a221oi_1 _1926_ (.B2(_1127_),
    .C1(net498),
    .B1(_1125_),
    .A1(net491),
    .Y(_1128_),
    .A2(_1118_));
 sg13g2_a21oi_1 _1927_ (.A1(_1109_),
    .A2(_1111_),
    .Y(_1129_),
    .B1(net505));
 sg13g2_o21ai_1 _1928_ (.B1(net509),
    .Y(_1130_),
    .A1(_1108_),
    .A2(_1110_));
 sg13g2_nand2_1 _1929_ (.Y(_1131_),
    .A(net494),
    .B(net470));
 sg13g2_nor3_1 _1930_ (.A(net509),
    .B(_1108_),
    .C(_1110_),
    .Y(_1132_));
 sg13g2_nand3_1 _1931_ (.B(_1109_),
    .C(_1111_),
    .A(net505),
    .Y(_1133_));
 sg13g2_nor2_2 _1932_ (.A(_1112_),
    .B(net479),
    .Y(_1134_));
 sg13g2_nand2_1 _1933_ (.Y(_1135_),
    .A(_1113_),
    .B(net476));
 sg13g2_nand2_1 _1934_ (.Y(_1136_),
    .A(net511),
    .B(net473));
 sg13g2_nand2_2 _1935_ (.Y(_1137_),
    .A(net474),
    .B(_1133_));
 sg13g2_nor2_1 _1936_ (.A(net482),
    .B(net471),
    .Y(_1138_));
 sg13g2_nor2_2 _1937_ (.A(net500),
    .B(net494),
    .Y(_1139_));
 sg13g2_a221oi_1 _1938_ (.B2(net494),
    .C1(net502),
    .B1(_1138_),
    .A1(_1131_),
    .Y(_1140_),
    .A2(_1137_));
 sg13g2_or2_1 _1939_ (.X(_1141_),
    .B(_1140_),
    .A(_1128_));
 sg13g2_nand2_1 _1940_ (.Y(_1142_),
    .A(\enigma.r.$signal$23[0] ),
    .B(_0000_));
 sg13g2_nor2_1 _1941_ (.A(\enigma.r.$signal$23[1] ),
    .B(_1142_),
    .Y(_1143_));
 sg13g2_or2_1 _1942_ (.X(_1144_),
    .B(_1142_),
    .A(\enigma.r.$signal$23[1] ));
 sg13g2_nor2_1 _1943_ (.A(net496),
    .B(net493),
    .Y(_1145_));
 sg13g2_nor2_1 _1944_ (.A(net475),
    .B(net472),
    .Y(_1146_));
 sg13g2_nand2_2 _1945_ (.Y(_1147_),
    .A(net479),
    .B(net469));
 sg13g2_mux2_1 _1946_ (.A0(_1112_),
    .A1(net472),
    .S(net480),
    .X(_1148_));
 sg13g2_nand2b_1 _1947_ (.Y(_1149_),
    .B(net466),
    .A_N(_1148_));
 sg13g2_nand2_1 _1948_ (.Y(_1150_),
    .A(net469),
    .B(_1133_));
 sg13g2_nor3_2 _1949_ (.A(net473),
    .B(net471),
    .C(net468),
    .Y(_1151_));
 sg13g2_nand3_1 _1950_ (.B(net470),
    .C(_1133_),
    .A(net480),
    .Y(_1152_));
 sg13g2_a221oi_1 _1951_ (.B2(net477),
    .C1(net504),
    .B1(_1117_),
    .A1(_1097_),
    .Y(_1153_),
    .A2(_1103_));
 sg13g2_o21ai_1 _1952_ (.B1(net470),
    .Y(_1154_),
    .A1(net508),
    .A2(net481));
 sg13g2_a221oi_1 _1953_ (.B2(_1048_),
    .C1(_1096_),
    .B1(_1102_),
    .A1(_1050_),
    .Y(_1155_),
    .A2(_1091_));
 sg13g2_nand2_1 _1954_ (.Y(_1156_),
    .A(net495),
    .B(net494));
 sg13g2_nand4_1 _1955_ (.B(net505),
    .C(_1109_),
    .A(_1001_),
    .Y(_1157_),
    .D(_1111_));
 sg13g2_nor2_2 _1956_ (.A(net495),
    .B(net485),
    .Y(_1158_));
 sg13g2_and3_1 _1957_ (.X(_1159_),
    .A(net503),
    .B(net492),
    .C(_1157_));
 sg13g2_a221oi_1 _1958_ (.B2(net467),
    .C1(_1159_),
    .B1(_1154_),
    .A1(_1152_),
    .Y(_1160_),
    .A2(_1153_));
 sg13g2_and2_2 _1959_ (.A(_1149_),
    .B(_1160_),
    .X(_1161_));
 sg13g2_nand2_1 _1960_ (.Y(_1162_),
    .A(\enigma.r.$signal$23[1] ),
    .B(_0000_));
 sg13g2_nor2_1 _1961_ (.A(\enigma.r.$signal$23[0] ),
    .B(_1162_),
    .Y(_1163_));
 sg13g2_inv_1 _1962_ (.Y(_1164_),
    .A(net551));
 sg13g2_nor2_2 _1963_ (.A(net487),
    .B(net483),
    .Y(_1165_));
 sg13g2_a21oi_1 _1964_ (.A1(net505),
    .A2(net481),
    .Y(_1166_),
    .B1(net502));
 sg13g2_o21ai_1 _1965_ (.B1(net490),
    .Y(_1167_),
    .A1(net510),
    .A2(net478));
 sg13g2_nor2_1 _1966_ (.A(net500),
    .B(net483),
    .Y(_1168_));
 sg13g2_nor2_1 _1967_ (.A(net495),
    .B(net483),
    .Y(_1169_));
 sg13g2_nor3_2 _1968_ (.A(net497),
    .B(net493),
    .C(net483),
    .Y(_1170_));
 sg13g2_nand2_2 _1969_ (.Y(_1171_),
    .A(net473),
    .B(net471));
 sg13g2_o21ai_1 _1970_ (.B1(net475),
    .Y(_1172_),
    .A1(net472),
    .A2(net468));
 sg13g2_a21oi_2 _1971_ (.B1(net480),
    .Y(_1173_),
    .A2(_1133_),
    .A1(net469));
 sg13g2_nor2_1 _1972_ (.A(net490),
    .B(_1116_),
    .Y(_1174_));
 sg13g2_nor2_1 _1973_ (.A(net501),
    .B(_1122_),
    .Y(_1175_));
 sg13g2_o21ai_1 _1974_ (.B1(net485),
    .Y(_1176_),
    .A1(net471),
    .A2(net468));
 sg13g2_nor4_1 _1975_ (.A(net504),
    .B(net491),
    .C(_1116_),
    .D(_1122_),
    .Y(_1177_));
 sg13g2_a221oi_1 _1976_ (.B2(_1172_),
    .C1(_1177_),
    .B1(_1170_),
    .A1(_1165_),
    .Y(_1178_),
    .A2(_1166_));
 sg13g2_nor2_1 _1977_ (.A(_1164_),
    .B(_1178_),
    .Y(_1179_));
 sg13g2_a221oi_1 _1978_ (.B2(_1161_),
    .C1(_1179_),
    .B1(net552),
    .A1(_0792_),
    .Y(_1180_),
    .A2(_1141_));
 sg13g2_nor3_2 _1979_ (.A(\enigma.r.$signal$23[1] ),
    .B(\enigma.r.$signal$23[0] ),
    .C(_0000_),
    .Y(_1181_));
 sg13g2_nand2b_1 _1980_ (.Y(_1182_),
    .B(_0789_),
    .A_N(_0000_));
 sg13g2_o21ai_1 _1981_ (.B1(net486),
    .Y(_1183_),
    .A1(_1112_),
    .A2(net479));
 sg13g2_a221oi_1 _1982_ (.B2(_1113_),
    .C1(net492),
    .B1(net474),
    .A1(net508),
    .Y(_1184_),
    .A2(net483));
 sg13g2_nor3_1 _1983_ (.A(net496),
    .B(_1165_),
    .C(_1184_),
    .Y(_1185_));
 sg13g2_a21oi_2 _1984_ (.B1(net493),
    .Y(_1186_),
    .A2(net468),
    .A1(net474));
 sg13g2_a22oi_1 _1985_ (.Y(_1187_),
    .B1(_1186_),
    .B2(net470),
    .A2(_1148_),
    .A1(net492));
 sg13g2_a21o_2 _1986_ (.A2(_1187_),
    .A1(net496),
    .B1(_1185_),
    .X(_1188_));
 sg13g2_and3_1 _1987_ (.X(_1189_),
    .A(\enigma.r.$signal$23[1] ),
    .B(\enigma.r.$signal$23[0] ),
    .C(_0000_));
 sg13g2_nand3_1 _1988_ (.B(_1109_),
    .C(_1111_),
    .A(_1000_),
    .Y(_1190_));
 sg13g2_a22oi_1 _1989_ (.Y(_1191_),
    .B1(net481),
    .B2(net506),
    .A2(_1112_),
    .A1(_1000_));
 sg13g2_nand2b_1 _1990_ (.Y(_1192_),
    .B(_1127_),
    .A_N(_1191_));
 sg13g2_a21o_2 _1991_ (.A2(_1118_),
    .A1(net503),
    .B1(net465),
    .X(_1193_));
 sg13g2_nor2_1 _1992_ (.A(net473),
    .B(_1123_),
    .Y(_1194_));
 sg13g2_nand2_2 _1993_ (.Y(_1195_),
    .A(net480),
    .B(_1122_));
 sg13g2_a21oi_2 _1994_ (.B1(net487),
    .Y(_1196_),
    .A2(net475),
    .A1(net508));
 sg13g2_a22oi_1 _1995_ (.Y(_1197_),
    .B1(_1196_),
    .B2(_1150_),
    .A2(_1195_),
    .A1(_1186_));
 sg13g2_a22oi_1 _1996_ (.Y(_1198_),
    .B1(_1197_),
    .B2(net499),
    .A2(_1193_),
    .A1(_1192_));
 sg13g2_a22oi_1 _1997_ (.Y(_1199_),
    .B1(net555),
    .B2(_1198_),
    .A2(_1188_),
    .A1(_1181_));
 sg13g2_a21oi_1 _1998_ (.A1(_1180_),
    .A2(_1199_),
    .Y(_1200_),
    .B1(_0790_));
 sg13g2_nand2_1 _1999_ (.Y(_1201_),
    .A(\enigma.r.$signal$21[1] ),
    .B(net579));
 sg13g2_nand2_2 _2000_ (.Y(_1202_),
    .A(_0001_),
    .B(_1201_));
 sg13g2_nor2_2 _2001_ (.A(\enigma.r.$signal$21[1] ),
    .B(net579),
    .Y(_1203_));
 sg13g2_nor2_1 _2002_ (.A(\enigma.r.$signal$21[2] ),
    .B(_1201_),
    .Y(_1204_));
 sg13g2_a21oi_2 _2003_ (.B1(_1204_),
    .Y(_1205_),
    .A2(_1203_),
    .A1(\enigma.r.$signal$21[2] ));
 sg13g2_a21oi_2 _2004_ (.B1(_0778_),
    .Y(_1206_),
    .A2(_1205_),
    .A1(_1202_));
 sg13g2_a21o_2 _2005_ (.A2(_1205_),
    .A1(_1202_),
    .B1(_0778_),
    .X(_1207_));
 sg13g2_nand2_1 _2006_ (.Y(_1208_),
    .A(net579),
    .B(_0001_));
 sg13g2_nor2_2 _2007_ (.A(\enigma.r.$signal$21[1] ),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_nand2_1 _2008_ (.Y(_1210_),
    .A(_1161_),
    .B(net550));
 sg13g2_and2_1 _2009_ (.A(_0001_),
    .B(_1203_),
    .X(_1211_));
 sg13g2_o21ai_1 _2010_ (.B1(_1211_),
    .Y(_1212_),
    .A1(_1128_),
    .A2(_1140_));
 sg13g2_nand2_1 _2011_ (.Y(_1213_),
    .A(\enigma.r.$signal$21[1] ),
    .B(_0001_));
 sg13g2_nor2_1 _2012_ (.A(net579),
    .B(_1213_),
    .Y(_1214_));
 sg13g2_or2_1 _2013_ (.X(_1215_),
    .B(_1213_),
    .A(net579));
 sg13g2_nand2b_1 _2014_ (.Y(_1216_),
    .B(_1214_),
    .A_N(_1178_));
 sg13g2_and3_1 _2015_ (.X(_1217_),
    .A(\enigma.r.$signal$21[1] ),
    .B(net579),
    .C(_0001_));
 sg13g2_nor3_2 _2016_ (.A(\enigma.r.$signal$21[1] ),
    .B(net579),
    .C(_0001_),
    .Y(_1218_));
 sg13g2_nand2b_2 _2017_ (.Y(_1219_),
    .B(_1203_),
    .A_N(_0001_));
 sg13g2_a22oi_1 _2018_ (.Y(_1220_),
    .B1(_1218_),
    .B2(_1188_),
    .A2(net554),
    .A1(_1198_));
 sg13g2_nand4_1 _2019_ (.B(_1212_),
    .C(_1216_),
    .A(_1210_),
    .Y(_1221_),
    .D(_1220_));
 sg13g2_nand2_1 _2020_ (.Y(_1222_),
    .A(\enigma.r.$signal$17[1] ),
    .B(net578));
 sg13g2_nand2_1 _2021_ (.Y(_1223_),
    .A(net576),
    .B(_1222_));
 sg13g2_nor2_2 _2022_ (.A(net577),
    .B(\enigma.r.$signal$17[0] ),
    .Y(_1224_));
 sg13g2_nor2_1 _2023_ (.A(\enigma.r.$signal$17[2] ),
    .B(_1222_),
    .Y(_1225_));
 sg13g2_a21oi_2 _2024_ (.B1(_1225_),
    .Y(_1226_),
    .A2(_1224_),
    .A1(\enigma.r.$signal$17[2] ));
 sg13g2_nand2_1 _2025_ (.Y(_1227_),
    .A(_1223_),
    .B(_1226_));
 sg13g2_and2_2 _2026_ (.A(net522),
    .B(_1227_),
    .X(_1228_));
 sg13g2_nand2_2 _2027_ (.Y(_1229_),
    .A(net522),
    .B(_1227_));
 sg13g2_nand2_1 _2028_ (.Y(_1230_),
    .A(net577),
    .B(net576));
 sg13g2_nor2_2 _2029_ (.A(\enigma.r.$signal$17[0] ),
    .B(_1230_),
    .Y(_1231_));
 sg13g2_or2_1 _2030_ (.X(_1232_),
    .B(_1230_),
    .A(net578));
 sg13g2_nand2b_1 _2031_ (.Y(_1233_),
    .B(_1231_),
    .A_N(_1178_));
 sg13g2_nand2_1 _2032_ (.Y(_1234_),
    .A(net578),
    .B(_0002_));
 sg13g2_nor2_1 _2033_ (.A(net577),
    .B(_1234_),
    .Y(_1235_));
 sg13g2_inv_1 _2034_ (.Y(_1236_),
    .A(net546));
 sg13g2_nand2_1 _2035_ (.Y(_1237_),
    .A(_1161_),
    .B(net546));
 sg13g2_and2_1 _2036_ (.A(net576),
    .B(_1224_),
    .X(_1238_));
 sg13g2_o21ai_1 _2037_ (.B1(_1238_),
    .Y(_1239_),
    .A1(_1128_),
    .A2(_1140_));
 sg13g2_and3_2 _2038_ (.X(_1240_),
    .A(net577),
    .B(net578),
    .C(net576));
 sg13g2_nand3_1 _2039_ (.B(net578),
    .C(net576),
    .A(net577),
    .Y(_1241_));
 sg13g2_nor3_2 _2040_ (.A(net577),
    .B(net578),
    .C(net576),
    .Y(_1242_));
 sg13g2_nand2b_2 _2041_ (.Y(_1243_),
    .B(_1224_),
    .A_N(net576));
 sg13g2_a22oi_1 _2042_ (.Y(_1244_),
    .B1(_1242_),
    .B2(_1188_),
    .A2(_1240_),
    .A1(_1198_));
 sg13g2_nand4_1 _2043_ (.B(_1237_),
    .C(_1239_),
    .A(_1233_),
    .Y(_1245_),
    .D(_1244_));
 sg13g2_a221oi_1 _2044_ (.B2(_1245_),
    .C1(_1200_),
    .B1(_1228_),
    .A1(_1206_),
    .Y(_1246_),
    .A2(_1221_));
 sg13g2_nand2_1 _2045_ (.Y(_1247_),
    .A(_0787_),
    .B(_1246_));
 sg13g2_xnor2_1 _2046_ (.Y(_1248_),
    .A(_0787_),
    .B(_1246_));
 sg13g2_nand3_1 _2047_ (.B(net484),
    .C(net507),
    .A(net495),
    .Y(_1249_));
 sg13g2_nand3_1 _2048_ (.B(_1139_),
    .C(_1147_),
    .A(_1136_),
    .Y(_1250_));
 sg13g2_o21ai_1 _2049_ (.B1(net467),
    .Y(_1251_),
    .A1(net479),
    .A2(net471));
 sg13g2_nand2_1 _2050_ (.Y(_1252_),
    .A(_1117_),
    .B(net480));
 sg13g2_a21oi_1 _2051_ (.A1(net469),
    .A2(_1133_),
    .Y(_1253_),
    .B1(net473));
 sg13g2_o21ai_1 _2052_ (.B1(net479),
    .Y(_1254_),
    .A1(net471),
    .A2(net468));
 sg13g2_o21ai_1 _2053_ (.B1(_1119_),
    .Y(_1255_),
    .A1(_1183_),
    .A2(_1253_));
 sg13g2_nand3_1 _2054_ (.B(_1251_),
    .C(_1255_),
    .A(_1250_),
    .Y(_1256_));
 sg13g2_nand2_1 _2055_ (.Y(_1257_),
    .A(net484),
    .B(net511));
 sg13g2_nor3_1 _2056_ (.A(net502),
    .B(net491),
    .C(net506),
    .Y(_1258_));
 sg13g2_a21oi_2 _2057_ (.B1(net500),
    .Y(_1259_),
    .A2(_1257_),
    .A1(_1134_));
 sg13g2_nand2b_1 _2058_ (.Y(_1260_),
    .B(_1119_),
    .A_N(_1154_));
 sg13g2_o21ai_1 _2059_ (.B1(net487),
    .Y(_1261_),
    .A1(net480),
    .A2(net472));
 sg13g2_a21oi_1 _2060_ (.A1(net481),
    .A2(net472),
    .Y(_1262_),
    .B1(_1261_));
 sg13g2_o21ai_1 _2061_ (.B1(net496),
    .Y(_1263_),
    .A1(net487),
    .A2(net474));
 sg13g2_o21ai_1 _2062_ (.B1(_1260_),
    .Y(_1264_),
    .A1(_1262_),
    .A2(_1263_));
 sg13g2_nor2_1 _2063_ (.A(net482),
    .B(_1122_),
    .Y(_1265_));
 sg13g2_nand2_1 _2064_ (.Y(_1266_),
    .A(net489),
    .B(net477));
 sg13g2_a21oi_1 _2065_ (.A1(net473),
    .A2(_1123_),
    .Y(_1267_),
    .B1(net490));
 sg13g2_o21ai_1 _2066_ (.B1(net489),
    .Y(_1268_),
    .A1(net482),
    .A2(_1122_));
 sg13g2_a21oi_1 _2067_ (.A1(_1147_),
    .A2(_1267_),
    .Y(_1269_),
    .B1(net499));
 sg13g2_a21oi_2 _2068_ (.B1(_1269_),
    .Y(_1270_),
    .A2(_1268_),
    .A1(_1167_));
 sg13g2_nor3_1 _2069_ (.A(net504),
    .B(net493),
    .C(_1132_),
    .Y(_1271_));
 sg13g2_o21ai_1 _2070_ (.B1(net509),
    .Y(_1272_),
    .A1(_1113_),
    .A2(net476));
 sg13g2_a221oi_1 _2071_ (.B2(net476),
    .C1(net488),
    .B1(_1117_),
    .A1(_1093_),
    .Y(_1273_),
    .A2(_1099_));
 sg13g2_nand2_2 _2072_ (.Y(_1274_),
    .A(_1116_),
    .B(net474));
 sg13g2_a221oi_1 _2073_ (.B2(_1170_),
    .C1(_1273_),
    .B1(_1274_),
    .A1(_1271_),
    .Y(_1275_),
    .A2(_1272_));
 sg13g2_nand2b_1 _2074_ (.Y(_1276_),
    .B(_1209_),
    .A_N(_1275_));
 sg13g2_a22oi_1 _2075_ (.Y(_1277_),
    .B1(_1270_),
    .B2(_1218_),
    .A2(_1259_),
    .A1(net548));
 sg13g2_a22oi_1 _2076_ (.Y(_1278_),
    .B1(_1264_),
    .B2(net554),
    .A2(_1256_),
    .A1(_1211_));
 sg13g2_nand3_1 _2077_ (.B(_1277_),
    .C(_1278_),
    .A(_1276_),
    .Y(_1279_));
 sg13g2_nor2_1 _2078_ (.A(_1236_),
    .B(_1275_),
    .Y(_1280_));
 sg13g2_a22oi_1 _2079_ (.Y(_1281_),
    .B1(_1264_),
    .B2(_1240_),
    .A2(_1259_),
    .A1(net547));
 sg13g2_a221oi_1 _2080_ (.B2(_1242_),
    .C1(_1280_),
    .B1(_1270_),
    .A1(_1238_),
    .Y(_0080_),
    .A2(_1256_));
 sg13g2_a21oi_1 _2081_ (.A1(_1281_),
    .A2(_0080_),
    .Y(_0081_),
    .B1(_1229_));
 sg13g2_a22oi_1 _2082_ (.Y(_0082_),
    .B1(_1264_),
    .B2(_1189_),
    .A2(_1259_),
    .A1(net551));
 sg13g2_nand2b_1 _2083_ (.Y(_0083_),
    .B(net552),
    .A_N(_1275_));
 sg13g2_a22oi_1 _2084_ (.Y(_0084_),
    .B1(_1270_),
    .B2(_1181_),
    .A2(_1256_),
    .A1(_0792_));
 sg13g2_nand3_1 _2085_ (.B(_0083_),
    .C(_0084_),
    .A(_0082_),
    .Y(_0085_));
 sg13g2_a221oi_1 _2086_ (.B2(_0791_),
    .C1(_0081_),
    .B1(_0085_),
    .A1(_1206_),
    .Y(_0086_),
    .A2(_1279_));
 sg13g2_nor2_1 _2087_ (.A(_0787_),
    .B(_0086_),
    .Y(_0087_));
 sg13g2_and2_2 _2088_ (.A(_0787_),
    .B(_0086_),
    .X(_0088_));
 sg13g2_nor3_1 _2089_ (.A(_0744_),
    .B(_0087_),
    .C(_0088_),
    .Y(_0089_));
 sg13g2_o21ai_1 _2090_ (.B1(net611),
    .Y(_0090_),
    .A1(_0743_),
    .A2(_1248_));
 sg13g2_nor2_1 _2091_ (.A(_0089_),
    .B(_0090_),
    .Y(_0013_));
 sg13g2_nor2_1 _2092_ (.A(net493),
    .B(_1113_),
    .Y(_0091_));
 sg13g2_o21ai_1 _2093_ (.B1(_1166_),
    .Y(_0092_),
    .A1(_1137_),
    .A2(_0091_));
 sg13g2_a21oi_2 _2094_ (.B1(net497),
    .Y(_0093_),
    .A2(_1157_),
    .A1(net493));
 sg13g2_a21o_2 _2095_ (.A2(_1157_),
    .A1(net492),
    .B1(net496),
    .X(_0094_));
 sg13g2_nor2_1 _2096_ (.A(net476),
    .B(net468),
    .Y(_0095_));
 sg13g2_a221oi_1 _2097_ (.B2(net472),
    .C1(_0095_),
    .B1(net476),
    .A1(_1097_),
    .Y(_0096_),
    .A2(_1103_));
 sg13g2_o21ai_1 _2098_ (.B1(_0092_),
    .Y(_0097_),
    .A1(_0094_),
    .A2(_0096_));
 sg13g2_a221oi_1 _2099_ (.B2(_0093_),
    .C1(_1258_),
    .B1(_1266_),
    .A1(net467),
    .Y(_0098_),
    .A2(_1265_));
 sg13g2_nor2b_1 _2100_ (.A(_0098_),
    .B_N(net545),
    .Y(_0099_));
 sg13g2_a21oi_1 _2101_ (.A1(_1242_),
    .A2(_0097_),
    .Y(_0100_),
    .B1(_0099_));
 sg13g2_nor2_1 _2102_ (.A(net506),
    .B(net477),
    .Y(_0101_));
 sg13g2_nand2_2 _2103_ (.Y(_0102_),
    .A(net508),
    .B(net481));
 sg13g2_mux2_1 _2104_ (.A0(net488),
    .A1(net509),
    .S(net482),
    .X(_0103_));
 sg13g2_a21oi_1 _2105_ (.A1(_1112_),
    .A2(_0103_),
    .Y(_0104_),
    .B1(net497));
 sg13g2_nor2_2 _2106_ (.A(net490),
    .B(net483),
    .Y(_0105_));
 sg13g2_a221oi_1 _2107_ (.B2(_1126_),
    .C1(net502),
    .B1(_0105_),
    .A1(_1135_),
    .Y(_0106_),
    .A2(_1165_));
 sg13g2_nor2_1 _2108_ (.A(_0104_),
    .B(_0106_),
    .Y(_0107_));
 sg13g2_a21oi_1 _2109_ (.A1(_1195_),
    .A2(_1267_),
    .Y(_0108_),
    .B1(_0094_));
 sg13g2_a21oi_1 _2110_ (.A1(net510),
    .A2(net482),
    .Y(_0109_),
    .B1(net502));
 sg13g2_a21o_1 _2111_ (.A2(_0109_),
    .A1(_1131_),
    .B1(_0108_),
    .X(_0110_));
 sg13g2_and4_1 _2112_ (.A(net498),
    .B(net489),
    .C(net506),
    .D(_1190_),
    .X(_0111_));
 sg13g2_a221oi_1 _2113_ (.B2(net476),
    .C1(net488),
    .B1(net508),
    .A1(_1093_),
    .Y(_0112_),
    .A2(_1099_));
 sg13g2_a221oi_1 _2114_ (.B2(_0112_),
    .C1(_0111_),
    .B1(_1195_),
    .A1(_1123_),
    .Y(_0113_),
    .A2(_1170_));
 sg13g2_nor2_1 _2115_ (.A(_1241_),
    .B(_0113_),
    .Y(_0114_));
 sg13g2_a221oi_1 _2116_ (.B2(net547),
    .C1(_0114_),
    .B1(_0110_),
    .A1(net546),
    .Y(_0115_),
    .A2(_0107_));
 sg13g2_a21oi_1 _2117_ (.A1(_0100_),
    .A2(_0115_),
    .Y(_0116_),
    .B1(_1229_));
 sg13g2_nor2b_1 _2118_ (.A(_0113_),
    .B_N(_1217_),
    .Y(_0117_));
 sg13g2_a21oi_1 _2119_ (.A1(_1218_),
    .A2(_0097_),
    .Y(_0118_),
    .B1(_0117_));
 sg13g2_nor2b_1 _2120_ (.A(_0098_),
    .B_N(net549),
    .Y(_0119_));
 sg13g2_a221oi_1 _2121_ (.B2(net548),
    .C1(_0119_),
    .B1(_0110_),
    .A1(net550),
    .Y(_0120_),
    .A2(_0107_));
 sg13g2_a21oi_1 _2122_ (.A1(_0118_),
    .A2(_0120_),
    .Y(_0121_),
    .B1(_1207_));
 sg13g2_a22oi_1 _2123_ (.Y(_0122_),
    .B1(_0110_),
    .B2(net551),
    .A2(_0097_),
    .A1(_1181_));
 sg13g2_nor2b_1 _2124_ (.A(_0113_),
    .B_N(net555),
    .Y(_0123_));
 sg13g2_nor2b_1 _2125_ (.A(_0098_),
    .B_N(net553),
    .Y(_0124_));
 sg13g2_nor3_1 _2126_ (.A(_1144_),
    .B(_0104_),
    .C(_0106_),
    .Y(_0125_));
 sg13g2_nor3_1 _2127_ (.A(_0123_),
    .B(_0124_),
    .C(_0125_),
    .Y(_0126_));
 sg13g2_a21oi_1 _2128_ (.A1(_0122_),
    .A2(_0126_),
    .Y(_0127_),
    .B1(_0790_));
 sg13g2_nor3_1 _2129_ (.A(_0116_),
    .B(_0121_),
    .C(_0127_),
    .Y(_0128_));
 sg13g2_nor2b_2 _2130_ (.A(_0128_),
    .B_N(_0920_),
    .Y(_0129_));
 sg13g2_nor4_2 _2131_ (.A(_0920_),
    .B(_0116_),
    .C(_0121_),
    .Y(_0130_),
    .D(_0127_));
 sg13g2_o21ai_1 _2132_ (.B1(_1247_),
    .Y(_0131_),
    .A1(_0129_),
    .A2(_0130_));
 sg13g2_or3_1 _2133_ (.A(_1247_),
    .B(_0129_),
    .C(_0130_),
    .X(_0132_));
 sg13g2_and2_1 _2134_ (.A(_0131_),
    .B(_0132_),
    .X(_0133_));
 sg13g2_a221oi_1 _2135_ (.B2(_1171_),
    .C1(net500),
    .B1(_1165_),
    .A1(net485),
    .Y(_0134_),
    .A2(_1147_));
 sg13g2_nor2_1 _2136_ (.A(_1151_),
    .B(_1173_),
    .Y(_0135_));
 sg13g2_o21ai_1 _2137_ (.B1(net465),
    .Y(_0136_),
    .A1(_1151_),
    .A2(_1173_));
 sg13g2_nand2b_2 _2138_ (.Y(_0137_),
    .B(_0136_),
    .A_N(_0134_));
 sg13g2_nor2_1 _2139_ (.A(net489),
    .B(_1133_),
    .Y(_0138_));
 sg13g2_nand2_1 _2140_ (.Y(_0139_),
    .A(net492),
    .B(_1137_));
 sg13g2_a21oi_1 _2141_ (.A1(_1261_),
    .A2(_0139_),
    .Y(_0140_),
    .B1(net503));
 sg13g2_nor3_1 _2142_ (.A(net495),
    .B(net484),
    .C(net483),
    .Y(_0141_));
 sg13g2_nand2_1 _2143_ (.Y(_0142_),
    .A(net503),
    .B(_1165_));
 sg13g2_nand3_1 _2144_ (.B(_1157_),
    .C(_1274_),
    .A(net465),
    .Y(_0143_));
 sg13g2_nand2_1 _2145_ (.Y(_0144_),
    .A(_0142_),
    .B(_0143_));
 sg13g2_nor2_2 _2146_ (.A(_0140_),
    .B(_0144_),
    .Y(_0145_));
 sg13g2_a21o_2 _2147_ (.A2(net475),
    .A1(_1113_),
    .B1(net483),
    .X(_0146_));
 sg13g2_nor3_2 _2148_ (.A(net501),
    .B(net494),
    .C(_0146_),
    .Y(_0147_));
 sg13g2_nor4_1 _2149_ (.A(net511),
    .B(_1158_),
    .C(_1232_),
    .D(_0147_),
    .Y(_0148_));
 sg13g2_a221oi_1 _2150_ (.B2(net546),
    .C1(_0148_),
    .B1(_0145_),
    .A1(net545),
    .Y(_0149_),
    .A2(_0137_));
 sg13g2_nand2b_1 _2151_ (.Y(_0150_),
    .B(_0102_),
    .A_N(_0146_));
 sg13g2_a221oi_1 _2152_ (.B2(_1155_),
    .C1(_1269_),
    .B1(_0150_),
    .A1(_1177_),
    .Y(_0151_),
    .A2(_0102_));
 sg13g2_nand3_1 _2153_ (.B(net465),
    .C(_0146_),
    .A(net507),
    .Y(_0152_));
 sg13g2_nand3_1 _2154_ (.B(_1126_),
    .C(_1152_),
    .A(net490),
    .Y(_0153_));
 sg13g2_a21oi_1 _2155_ (.A1(net484),
    .A2(_1191_),
    .Y(_0154_),
    .B1(net501));
 sg13g2_nand2_1 _2156_ (.Y(_0155_),
    .A(_0153_),
    .B(_0154_));
 sg13g2_nand2_2 _2157_ (.Y(_0156_),
    .A(_0152_),
    .B(_0155_));
 sg13g2_a22oi_1 _2158_ (.Y(_0157_),
    .B1(_0156_),
    .B2(_1242_),
    .A2(_0151_),
    .A1(_1240_));
 sg13g2_a21oi_1 _2159_ (.A1(_0149_),
    .A2(_0157_),
    .Y(_0158_),
    .B1(_1229_));
 sg13g2_nor4_1 _2160_ (.A(net511),
    .B(_1158_),
    .C(_1215_),
    .D(_0147_),
    .Y(_0159_));
 sg13g2_a221oi_1 _2161_ (.B2(net550),
    .C1(_0159_),
    .B1(_0145_),
    .A1(net549),
    .Y(_0160_),
    .A2(_0137_));
 sg13g2_a22oi_1 _2162_ (.Y(_0161_),
    .B1(_0156_),
    .B2(_1218_),
    .A2(_0151_),
    .A1(net554));
 sg13g2_a21oi_1 _2163_ (.A1(_0160_),
    .A2(_0161_),
    .Y(_0162_),
    .B1(_1207_));
 sg13g2_nor4_1 _2164_ (.A(net511),
    .B(_1158_),
    .C(_1164_),
    .D(_0147_),
    .Y(_0163_));
 sg13g2_a221oi_1 _2165_ (.B2(net552),
    .C1(_0163_),
    .B1(_0145_),
    .A1(net553),
    .Y(_0164_),
    .A2(_0137_));
 sg13g2_a22oi_1 _2166_ (.Y(_0165_),
    .B1(_0156_),
    .B2(_1181_),
    .A2(_0151_),
    .A1(net555));
 sg13g2_a21oi_1 _2167_ (.A1(_0164_),
    .A2(_0165_),
    .Y(_0166_),
    .B1(_0790_));
 sg13g2_nor3_1 _2168_ (.A(_0158_),
    .B(_0162_),
    .C(_0166_),
    .Y(_0167_));
 sg13g2_and2_1 _2169_ (.A(_1084_),
    .B(_0167_),
    .X(_0168_));
 sg13g2_o21ai_1 _2170_ (.B1(net489),
    .Y(_0169_),
    .A1(_0101_),
    .A2(_0146_));
 sg13g2_nand3b_1 _2171_ (.B(net491),
    .C(_1152_),
    .Y(_0170_),
    .A_N(_1265_));
 sg13g2_a21oi_1 _2172_ (.A1(_0169_),
    .A2(_0170_),
    .Y(_0171_),
    .B1(net502));
 sg13g2_nand2_2 _2173_ (.Y(_0172_),
    .A(net475),
    .B(_1122_));
 sg13g2_a21oi_2 _2174_ (.B1(_0094_),
    .Y(_0173_),
    .A2(_0172_),
    .A1(_0105_));
 sg13g2_o21ai_1 _2175_ (.B1(net545),
    .Y(_0174_),
    .A1(_0171_),
    .A2(_0173_));
 sg13g2_a21oi_2 _2176_ (.B1(net503),
    .Y(_0175_),
    .A2(_1174_),
    .A1(_1126_));
 sg13g2_a21oi_2 _2177_ (.B1(net487),
    .Y(_0176_),
    .A2(net470),
    .A1(net475));
 sg13g2_o21ai_1 _2178_ (.B1(_1157_),
    .Y(_0177_),
    .A1(_0138_),
    .A2(_0176_));
 sg13g2_a21oi_2 _2179_ (.B1(net493),
    .Y(_0178_),
    .A2(net481),
    .A1(_1117_));
 sg13g2_mux2_1 _2180_ (.A0(_1116_),
    .A1(net471),
    .S(net474),
    .X(_0179_));
 sg13g2_nand2_1 _2181_ (.Y(_0180_),
    .A(net486),
    .B(_0179_));
 sg13g2_a22oi_1 _2182_ (.Y(_0181_),
    .B1(_0180_),
    .B2(_1193_),
    .A2(_0177_),
    .A1(_0175_));
 sg13g2_a221oi_1 _2183_ (.B2(_1193_),
    .C1(_1241_),
    .B1(_0180_),
    .A1(_0175_),
    .Y(_0182_),
    .A2(_0177_));
 sg13g2_and2_1 _2184_ (.A(net507),
    .B(net467),
    .X(_0183_));
 sg13g2_a221oi_1 _2185_ (.B2(_0183_),
    .C1(_0141_),
    .B1(_0146_),
    .A1(_1186_),
    .Y(_0184_),
    .A2(_1195_));
 sg13g2_and2_1 _2186_ (.A(net547),
    .B(_0184_),
    .X(_0185_));
 sg13g2_a21oi_1 _2187_ (.A1(_1152_),
    .A2(_1172_),
    .Y(_0186_),
    .B1(_1156_));
 sg13g2_a221oi_1 _2188_ (.B2(net479),
    .C1(net495),
    .B1(net468),
    .A1(net484),
    .Y(_0187_),
    .A2(net471));
 sg13g2_a21o_1 _2189_ (.A2(_1139_),
    .A1(net479),
    .B1(_0187_),
    .X(_0188_));
 sg13g2_nor2_1 _2190_ (.A(_0186_),
    .B(_0188_),
    .Y(_0189_));
 sg13g2_nor3_1 _2191_ (.A(_1243_),
    .B(_0186_),
    .C(_0188_),
    .Y(_0190_));
 sg13g2_o21ai_1 _2192_ (.B1(_0093_),
    .Y(_0191_),
    .A1(_1261_),
    .A2(_0095_));
 sg13g2_o21ai_1 _2193_ (.B1(_1133_),
    .Y(_0192_),
    .A1(net479),
    .A2(net469));
 sg13g2_a221oi_1 _2194_ (.B2(net474),
    .C1(net492),
    .B1(_1117_),
    .A1(_1001_),
    .Y(_0193_),
    .A2(_1112_));
 sg13g2_o21ai_1 _2195_ (.B1(_0105_),
    .Y(_0194_),
    .A1(_1116_),
    .A2(net480));
 sg13g2_a22oi_1 _2196_ (.Y(_0195_),
    .B1(_0193_),
    .B2(_0109_),
    .A2(_0192_),
    .A1(net467));
 sg13g2_nand2_1 _2197_ (.Y(_0196_),
    .A(_0191_),
    .B(_0195_));
 sg13g2_a21oi_1 _2198_ (.A1(_0191_),
    .A2(_0195_),
    .Y(_0197_),
    .B1(_1236_));
 sg13g2_nor4_1 _2199_ (.A(_0182_),
    .B(_0185_),
    .C(_0190_),
    .D(_0197_),
    .Y(_0198_));
 sg13g2_a21oi_1 _2200_ (.A1(_0174_),
    .A2(_0198_),
    .Y(_0199_),
    .B1(_1229_));
 sg13g2_o21ai_1 _2201_ (.B1(net549),
    .Y(_0200_),
    .A1(_0171_),
    .A2(_0173_));
 sg13g2_a22oi_1 _2202_ (.Y(_0201_),
    .B1(_0196_),
    .B2(net550),
    .A2(_0184_),
    .A1(net548));
 sg13g2_a22oi_1 _2203_ (.Y(_0202_),
    .B1(_0189_),
    .B2(_1218_),
    .A2(_0181_),
    .A1(net554));
 sg13g2_nand3_1 _2204_ (.B(_0201_),
    .C(_0202_),
    .A(_0200_),
    .Y(_0203_));
 sg13g2_o21ai_1 _2205_ (.B1(net553),
    .Y(_0204_),
    .A1(_0171_),
    .A2(_0173_));
 sg13g2_nand2_1 _2206_ (.Y(_0205_),
    .A(net555),
    .B(_0181_));
 sg13g2_nand2_1 _2207_ (.Y(_0206_),
    .A(net552),
    .B(_0196_));
 sg13g2_a22oi_1 _2208_ (.Y(_0207_),
    .B1(_0189_),
    .B2(_1181_),
    .A2(_0184_),
    .A1(_1163_));
 sg13g2_nand4_1 _2209_ (.B(_0205_),
    .C(_0206_),
    .A(_0204_),
    .Y(_0208_),
    .D(_0207_));
 sg13g2_a221oi_1 _2210_ (.B2(_0791_),
    .C1(_0199_),
    .B1(_0208_),
    .A1(_1206_),
    .Y(_0209_),
    .A2(_0203_));
 sg13g2_nand2_1 _2211_ (.Y(_0210_),
    .A(net514),
    .B(_0209_));
 sg13g2_nand3_1 _2212_ (.B(_1147_),
    .C(_1190_),
    .A(net486),
    .Y(_0211_));
 sg13g2_a221oi_1 _2213_ (.B2(net476),
    .C1(net488),
    .B1(net505),
    .A1(_1093_),
    .Y(_0212_),
    .A2(_1099_));
 sg13g2_a21oi_1 _2214_ (.A1(_1136_),
    .A2(_1147_),
    .Y(_0213_),
    .B1(_1156_));
 sg13g2_a221oi_1 _2215_ (.B2(net500),
    .C1(_0213_),
    .B1(_0211_),
    .A1(_1139_),
    .Y(_0214_),
    .A2(_0135_));
 sg13g2_a22oi_1 _2216_ (.Y(_0215_),
    .B1(_0179_),
    .B2(_1139_),
    .A2(_1253_),
    .A1(net467));
 sg13g2_o21ai_1 _2217_ (.B1(_0215_),
    .Y(_0216_),
    .A1(_0094_),
    .A2(_0193_));
 sg13g2_a22oi_1 _2218_ (.Y(_0217_),
    .B1(_0216_),
    .B2(_1240_),
    .A2(_0214_),
    .A1(net546));
 sg13g2_nand3_1 _2219_ (.B(_1171_),
    .C(_1195_),
    .A(_1139_),
    .Y(_0218_));
 sg13g2_nand3_1 _2220_ (.B(net467),
    .C(_0172_),
    .A(_1117_),
    .Y(_0219_));
 sg13g2_nand2_1 _2221_ (.Y(_0220_),
    .A(net466),
    .B(_0192_));
 sg13g2_o21ai_1 _2222_ (.B1(net466),
    .Y(_0221_),
    .A1(_1146_),
    .A2(_1173_));
 sg13g2_and4_2 _2223_ (.A(_0142_),
    .B(_0218_),
    .C(_0219_),
    .D(_0221_),
    .X(_0222_));
 sg13g2_a22oi_1 _2224_ (.Y(_0223_),
    .B1(net473),
    .B2(net507),
    .A2(_1112_),
    .A1(net485));
 sg13g2_nand2_1 _2225_ (.Y(_0224_),
    .A(_1168_),
    .B(_0223_));
 sg13g2_o21ai_1 _2226_ (.B1(net465),
    .Y(_0225_),
    .A1(_1173_),
    .A2(_1194_));
 sg13g2_a21oi_1 _2227_ (.A1(_0224_),
    .A2(_0225_),
    .Y(_0226_),
    .B1(_1243_));
 sg13g2_or3_1 _2228_ (.A(_1186_),
    .B(_0138_),
    .C(_0176_),
    .X(_0227_));
 sg13g2_a22oi_1 _2229_ (.Y(_0228_),
    .B1(_0227_),
    .B2(net495),
    .A2(_1257_),
    .A1(_1169_));
 sg13g2_a221oi_1 _2230_ (.B2(net547),
    .C1(_0226_),
    .B1(_0228_),
    .A1(net545),
    .Y(_0229_),
    .A2(_0222_));
 sg13g2_a21oi_1 _2231_ (.A1(_0217_),
    .A2(_0229_),
    .Y(_0230_),
    .B1(_1229_));
 sg13g2_a21oi_1 _2232_ (.A1(_0224_),
    .A2(_0225_),
    .Y(_0231_),
    .B1(_1219_));
 sg13g2_a22oi_1 _2233_ (.Y(_0232_),
    .B1(_0222_),
    .B2(net549),
    .A2(_0214_),
    .A1(net550));
 sg13g2_a221oi_1 _2234_ (.B2(net548),
    .C1(_0231_),
    .B1(_0228_),
    .A1(net554),
    .Y(_0233_),
    .A2(_0216_));
 sg13g2_a21oi_1 _2235_ (.A1(_0232_),
    .A2(_0233_),
    .Y(_0234_),
    .B1(_1207_));
 sg13g2_a22oi_1 _2236_ (.Y(_0235_),
    .B1(_0216_),
    .B2(net555),
    .A2(_0214_),
    .A1(net552));
 sg13g2_a21oi_1 _2237_ (.A1(_0224_),
    .A2(_0225_),
    .Y(_0236_),
    .B1(_1182_));
 sg13g2_a221oi_1 _2238_ (.B2(net551),
    .C1(_0236_),
    .B1(_0228_),
    .A1(net553),
    .Y(_0237_),
    .A2(_0222_));
 sg13g2_a21oi_1 _2239_ (.A1(_0235_),
    .A2(_0237_),
    .Y(_0238_),
    .B1(_0790_));
 sg13g2_nor3_2 _2240_ (.A(_0230_),
    .B(_0234_),
    .C(_0238_),
    .Y(_0239_));
 sg13g2_nand2_1 _2241_ (.Y(_0240_),
    .A(_1041_),
    .B(_0239_));
 sg13g2_nor2_1 _2242_ (.A(_1041_),
    .B(_0239_),
    .Y(_0241_));
 sg13g2_xnor2_1 _2243_ (.Y(_0242_),
    .A(_1041_),
    .B(_0239_));
 sg13g2_nor2_1 _2244_ (.A(net514),
    .B(_0209_),
    .Y(_0243_));
 sg13g2_nor2_1 _2245_ (.A(_0242_),
    .B(_0243_),
    .Y(_0244_));
 sg13g2_inv_1 _2246_ (.Y(_0245_),
    .A(_0244_));
 sg13g2_xor2_1 _2247_ (.B(_0209_),
    .A(net514),
    .X(_0246_));
 sg13g2_nor2b_1 _2248_ (.A(_0242_),
    .B_N(_0246_),
    .Y(_0247_));
 sg13g2_nor3_1 _2249_ (.A(_0787_),
    .B(_1246_),
    .C(_0130_),
    .Y(_0248_));
 sg13g2_nor2_1 _2250_ (.A(_0129_),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_a21oi_1 _2251_ (.A1(_0210_),
    .A2(_0240_),
    .Y(_0250_),
    .B1(_0241_));
 sg13g2_a21o_1 _2252_ (.A2(_0249_),
    .A1(_0247_),
    .B1(_0250_),
    .X(_0251_));
 sg13g2_nor2_1 _2253_ (.A(_1084_),
    .B(_0167_),
    .Y(_0252_));
 sg13g2_nor3_1 _2254_ (.A(_1248_),
    .B(_0129_),
    .C(_0130_),
    .Y(_0253_));
 sg13g2_a21oi_1 _2255_ (.A1(_0247_),
    .A2(_0253_),
    .Y(_0254_),
    .B1(_0252_));
 sg13g2_a21oi_2 _2256_ (.B1(_0168_),
    .Y(_0255_),
    .A2(_0254_),
    .A1(_0251_));
 sg13g2_a21oi_1 _2257_ (.A1(_0133_),
    .A2(_0255_),
    .Y(_0256_),
    .B1(_0743_));
 sg13g2_o21ai_1 _2258_ (.B1(_0256_),
    .Y(_0257_),
    .A1(_0133_),
    .A2(_0255_));
 sg13g2_a21oi_1 _2259_ (.A1(_1127_),
    .A2(_0146_),
    .Y(_0258_),
    .B1(_0094_));
 sg13g2_nand2_1 _2260_ (.Y(_0259_),
    .A(_1152_),
    .B(_1186_));
 sg13g2_a21oi_1 _2261_ (.A1(net494),
    .A2(_1137_),
    .Y(_0260_),
    .B1(net501));
 sg13g2_a21o_1 _2262_ (.A2(_0260_),
    .A1(_0259_),
    .B1(_0258_),
    .X(_0261_));
 sg13g2_mux4_1 _2263_ (.S0(net487),
    .A0(_1115_),
    .A1(_1117_),
    .A2(net468),
    .A3(_1126_),
    .S1(net496),
    .X(_0262_));
 sg13g2_nor2_1 _2264_ (.A(_1219_),
    .B(_0262_),
    .Y(_0263_));
 sg13g2_nand3_1 _2265_ (.B(net469),
    .C(_1190_),
    .A(net490),
    .Y(_0264_));
 sg13g2_nor2_1 _2266_ (.A(_0094_),
    .B(_0178_),
    .Y(_0265_));
 sg13g2_a21o_1 _2267_ (.A2(_0264_),
    .A1(_0175_),
    .B1(_0265_),
    .X(_0266_));
 sg13g2_a221oi_1 _2268_ (.B2(net549),
    .C1(_0263_),
    .B1(_0266_),
    .A1(net554),
    .Y(_0267_),
    .A2(_0261_));
 sg13g2_nand2_1 _2269_ (.Y(_0268_),
    .A(net484),
    .B(_1134_));
 sg13g2_o21ai_1 _2270_ (.B1(_1249_),
    .Y(_0269_),
    .A1(_1151_),
    .A2(_1156_));
 sg13g2_o21ai_1 _2271_ (.B1(net484),
    .Y(_0270_),
    .A1(_1151_),
    .A2(_1173_));
 sg13g2_a22oi_1 _2272_ (.Y(_0271_),
    .B1(_0270_),
    .B2(_1193_),
    .A2(_0269_),
    .A1(_0268_));
 sg13g2_nand3_1 _2273_ (.B(_1118_),
    .C(_0172_),
    .A(net490),
    .Y(_0272_));
 sg13g2_a21oi_1 _2274_ (.A1(_1137_),
    .A2(_0105_),
    .Y(_0273_),
    .B1(net503));
 sg13g2_nand2_1 _2275_ (.Y(_0274_),
    .A(_1137_),
    .B(_1252_));
 sg13g2_a221oi_1 _2276_ (.B2(net465),
    .C1(_1159_),
    .B1(_0274_),
    .A1(_0272_),
    .Y(_0275_),
    .A2(_0273_));
 sg13g2_a22oi_1 _2277_ (.Y(_0276_),
    .B1(_0275_),
    .B2(net550),
    .A2(_0271_),
    .A1(net548));
 sg13g2_a21oi_1 _2278_ (.A1(_0267_),
    .A2(_0276_),
    .Y(_0277_),
    .B1(_1207_));
 sg13g2_nor2_1 _2279_ (.A(_1182_),
    .B(_0262_),
    .Y(_0278_));
 sg13g2_a221oi_1 _2280_ (.B2(net553),
    .C1(_0278_),
    .B1(_0266_),
    .A1(net555),
    .Y(_0279_),
    .A2(_0261_));
 sg13g2_a22oi_1 _2281_ (.Y(_0280_),
    .B1(_0275_),
    .B2(net552),
    .A2(_0271_),
    .A1(net551));
 sg13g2_a21oi_1 _2282_ (.A1(_0279_),
    .A2(_0280_),
    .Y(_0281_),
    .B1(_0790_));
 sg13g2_nor2_1 _2283_ (.A(_1243_),
    .B(_0262_),
    .Y(_0282_));
 sg13g2_a221oi_1 _2284_ (.B2(net545),
    .C1(_0282_),
    .B1(_0266_),
    .A1(_1240_),
    .Y(_0283_),
    .A2(_0261_));
 sg13g2_a22oi_1 _2285_ (.Y(_0284_),
    .B1(_0275_),
    .B2(net546),
    .A2(_0271_),
    .A1(net547));
 sg13g2_a21oi_1 _2286_ (.A1(_0283_),
    .A2(_0284_),
    .Y(_0285_),
    .B1(_1229_));
 sg13g2_nor3_2 _2287_ (.A(_0277_),
    .B(_0281_),
    .C(_0285_),
    .Y(_0286_));
 sg13g2_nor2b_1 _2288_ (.A(_0920_),
    .B_N(_0286_),
    .Y(_0287_));
 sg13g2_nand2b_1 _2289_ (.Y(_0288_),
    .B(_0286_),
    .A_N(_0920_));
 sg13g2_nor2b_1 _2290_ (.A(_0286_),
    .B_N(_0920_),
    .Y(_0289_));
 sg13g2_xnor2_1 _2291_ (.Y(_0290_),
    .A(_0920_),
    .B(_0286_));
 sg13g2_nor2_1 _2292_ (.A(_0088_),
    .B(_0290_),
    .Y(_0291_));
 sg13g2_xnor2_1 _2293_ (.Y(_0292_),
    .A(_0088_),
    .B(_0290_));
 sg13g2_nand2_1 _2294_ (.Y(_0293_),
    .A(_1137_),
    .B(_0178_));
 sg13g2_a21oi_1 _2295_ (.A1(_0102_),
    .A2(_0176_),
    .Y(_0294_),
    .B1(net502));
 sg13g2_a22oi_1 _2296_ (.Y(_0295_),
    .B1(_0294_),
    .B2(_0169_),
    .A2(_0293_),
    .A1(net502));
 sg13g2_nor2_1 _2297_ (.A(_1184_),
    .B(_0094_),
    .Y(_0296_));
 sg13g2_or2_1 _2298_ (.X(_0297_),
    .B(_0296_),
    .A(_0112_));
 sg13g2_nand2_1 _2299_ (.Y(_0298_),
    .A(net548),
    .B(_0297_));
 sg13g2_nand3_1 _2300_ (.B(_1126_),
    .C(_0102_),
    .A(net487),
    .Y(_0299_));
 sg13g2_a21oi_1 _2301_ (.A1(net508),
    .A2(net480),
    .Y(_0300_),
    .B1(_1113_));
 sg13g2_o21ai_1 _2302_ (.B1(net496),
    .Y(_0301_),
    .A1(net487),
    .A2(_0300_));
 sg13g2_a21oi_2 _2303_ (.B1(_1153_),
    .Y(_0302_),
    .A2(_0301_),
    .A1(_0299_));
 sg13g2_o21ai_1 _2304_ (.B1(net467),
    .Y(_0303_),
    .A1(_1173_),
    .A2(_1194_));
 sg13g2_o21ai_1 _2305_ (.B1(_0303_),
    .Y(_0304_),
    .A1(net499),
    .A2(_1262_));
 sg13g2_a21oi_2 _2306_ (.B1(_0304_),
    .Y(_0305_),
    .A2(_1171_),
    .A1(_1139_));
 sg13g2_a22oi_1 _2307_ (.Y(_0306_),
    .B1(_1165_),
    .B2(net511),
    .A2(_1134_),
    .A1(net484));
 sg13g2_nor2b_2 _2308_ (.A(_1159_),
    .B_N(_1249_),
    .Y(_0307_));
 sg13g2_o21ai_1 _2309_ (.B1(_0307_),
    .Y(_0308_),
    .A1(net500),
    .A2(_0306_));
 sg13g2_a21oi_2 _2310_ (.B1(_0308_),
    .Y(_0309_),
    .A2(_1195_),
    .A1(net465));
 sg13g2_a22oi_1 _2311_ (.Y(_0310_),
    .B1(_0305_),
    .B2(net549),
    .A2(_0295_),
    .A1(_1218_));
 sg13g2_a22oi_1 _2312_ (.Y(_0311_),
    .B1(_0309_),
    .B2(net554),
    .A2(_0302_),
    .A1(net550));
 sg13g2_nand3_1 _2313_ (.B(_0310_),
    .C(_0311_),
    .A(_0298_),
    .Y(_0312_));
 sg13g2_a22oi_1 _2314_ (.Y(_0313_),
    .B1(_0309_),
    .B2(net555),
    .A2(_0302_),
    .A1(net552));
 sg13g2_nand2_1 _2315_ (.Y(_0314_),
    .A(net551),
    .B(_0297_));
 sg13g2_a22oi_1 _2316_ (.Y(_0315_),
    .B1(_0305_),
    .B2(net553),
    .A2(_0295_),
    .A1(_1181_));
 sg13g2_nand3_1 _2317_ (.B(_0314_),
    .C(_0315_),
    .A(_0313_),
    .Y(_0316_));
 sg13g2_nand2_1 _2318_ (.Y(_0317_),
    .A(_0791_),
    .B(_0316_));
 sg13g2_nand2_1 _2319_ (.Y(_0318_),
    .A(net545),
    .B(_0305_));
 sg13g2_a22oi_1 _2320_ (.Y(_0319_),
    .B1(_0302_),
    .B2(net546),
    .A2(_0295_),
    .A1(_1242_));
 sg13g2_a22oi_1 _2321_ (.Y(_0320_),
    .B1(_0309_),
    .B2(_1240_),
    .A2(_0297_),
    .A1(net547));
 sg13g2_nand3_1 _2322_ (.B(_0319_),
    .C(_0320_),
    .A(_0318_),
    .Y(_0321_));
 sg13g2_a22oi_1 _2323_ (.Y(_0322_),
    .B1(_0321_),
    .B2(_1228_),
    .A2(_0312_),
    .A1(_1206_));
 sg13g2_nand3_1 _2324_ (.B(_0317_),
    .C(_0322_),
    .A(_1084_),
    .Y(_0323_));
 sg13g2_a21o_1 _2325_ (.A2(_0259_),
    .A1(_0153_),
    .B1(net500),
    .X(_0324_));
 sg13g2_o21ai_1 _2326_ (.B1(_1193_),
    .Y(_0325_),
    .A1(_1257_),
    .A2(_0146_));
 sg13g2_nand3_1 _2327_ (.B(_0324_),
    .C(_0325_),
    .A(net553),
    .Y(_0326_));
 sg13g2_o21ai_1 _2328_ (.B1(_1252_),
    .Y(_0327_),
    .A1(_1127_),
    .A2(_1196_));
 sg13g2_a22oi_1 _2329_ (.Y(_0328_),
    .B1(_0327_),
    .B2(net498),
    .A2(_0194_),
    .A1(_1193_));
 sg13g2_nand2_1 _2330_ (.Y(_0329_),
    .A(_1181_),
    .B(_0328_));
 sg13g2_o21ai_1 _2331_ (.B1(_1119_),
    .Y(_0330_),
    .A1(net492),
    .A2(_0300_));
 sg13g2_nand2_1 _2332_ (.Y(_0331_),
    .A(net498),
    .B(_1268_));
 sg13g2_o21ai_1 _2333_ (.B1(_0330_),
    .Y(_0332_),
    .A1(_0176_),
    .A2(_0331_));
 sg13g2_a22oi_1 _2334_ (.Y(_0333_),
    .B1(_0146_),
    .B2(net465),
    .A2(_1183_),
    .A1(_1175_));
 sg13g2_and3_1 _2335_ (.X(_0334_),
    .A(net552),
    .B(_0307_),
    .C(_0333_));
 sg13g2_a22oi_1 _2336_ (.Y(_0335_),
    .B1(_0176_),
    .B2(_1152_),
    .A2(_0105_),
    .A1(net469));
 sg13g2_o21ai_1 _2337_ (.B1(_0220_),
    .Y(_0336_),
    .A1(net503),
    .A2(_0335_));
 sg13g2_a221oi_1 _2338_ (.B2(net555),
    .C1(_0334_),
    .B1(_0336_),
    .A1(net551),
    .Y(_0337_),
    .A2(_0332_));
 sg13g2_nand3_1 _2339_ (.B(_0329_),
    .C(_0337_),
    .A(_0326_),
    .Y(_0338_));
 sg13g2_nand3_1 _2340_ (.B(_0324_),
    .C(_0325_),
    .A(net549),
    .Y(_0339_));
 sg13g2_nand2_1 _2341_ (.Y(_0340_),
    .A(_1218_),
    .B(_0328_));
 sg13g2_nand3_1 _2342_ (.B(_0307_),
    .C(_0333_),
    .A(net550),
    .Y(_0341_));
 sg13g2_nand2_1 _2343_ (.Y(_0342_),
    .A(net548),
    .B(_0332_));
 sg13g2_nand2_1 _2344_ (.Y(_0343_),
    .A(net554),
    .B(_0336_));
 sg13g2_nand3_1 _2345_ (.B(_0341_),
    .C(_0342_),
    .A(_0340_),
    .Y(_0344_));
 sg13g2_nand2_1 _2346_ (.Y(_0345_),
    .A(_0339_),
    .B(_0343_));
 sg13g2_o21ai_1 _2347_ (.B1(_1206_),
    .Y(_0346_),
    .A1(_0344_),
    .A2(_0345_));
 sg13g2_nand3_1 _2348_ (.B(_0324_),
    .C(_0325_),
    .A(net545),
    .Y(_0347_));
 sg13g2_nand2_1 _2349_ (.Y(_0348_),
    .A(_1242_),
    .B(_0328_));
 sg13g2_nand3_1 _2350_ (.B(_0307_),
    .C(_0333_),
    .A(net546),
    .Y(_0349_));
 sg13g2_a22oi_1 _2351_ (.Y(_0350_),
    .B1(_0336_),
    .B2(_1240_),
    .A2(_0332_),
    .A1(net547));
 sg13g2_nand4_1 _2352_ (.B(_0348_),
    .C(_0349_),
    .A(_0347_),
    .Y(_0351_),
    .D(_0350_));
 sg13g2_a22oi_1 _2353_ (.Y(_0352_),
    .B1(_0351_),
    .B2(_1228_),
    .A2(_0338_),
    .A1(_0791_));
 sg13g2_nand3_1 _2354_ (.B(_0346_),
    .C(_0352_),
    .A(_1041_),
    .Y(_0353_));
 sg13g2_a21o_2 _2355_ (.A2(_0352_),
    .A1(_0346_),
    .B1(_1041_),
    .X(_0354_));
 sg13g2_nand2_2 _2356_ (.Y(_0355_),
    .A(_0353_),
    .B(_0354_));
 sg13g2_a22oi_1 _2357_ (.Y(_0356_),
    .B1(_1274_),
    .B2(_0178_),
    .A2(_1196_),
    .A1(_1191_));
 sg13g2_a22oi_1 _2358_ (.Y(_0357_),
    .B1(_0356_),
    .B2(net497),
    .A2(net466),
    .A1(_1124_));
 sg13g2_nor2b_1 _2359_ (.A(_0357_),
    .B_N(net549),
    .Y(_0358_));
 sg13g2_a21oi_2 _2360_ (.B1(_0094_),
    .Y(_0359_),
    .A2(_0105_),
    .A1(net469));
 sg13g2_a21o_1 _2361_ (.A2(net475),
    .A1(net489),
    .B1(_1114_),
    .X(_0360_));
 sg13g2_a221oi_1 _2362_ (.B2(_1133_),
    .C1(net503),
    .B1(_0360_),
    .A1(net490),
    .Y(_0361_),
    .A2(_1150_));
 sg13g2_o21ai_1 _2363_ (.B1(_1217_),
    .Y(_0362_),
    .A1(_0359_),
    .A2(_0361_));
 sg13g2_a22oi_1 _2364_ (.Y(_0363_),
    .B1(_0223_),
    .B2(_1168_),
    .A2(_1176_),
    .A1(_1119_));
 sg13g2_nand2b_1 _2365_ (.Y(_0364_),
    .B(net548),
    .A_N(_0363_));
 sg13g2_nand3b_1 _2366_ (.B(_1127_),
    .C(net500),
    .Y(_0365_),
    .A_N(_1191_));
 sg13g2_a221oi_1 _2367_ (.B2(_0212_),
    .C1(_0141_),
    .B1(_1254_),
    .A1(_1139_),
    .Y(_0366_),
    .A2(_1171_));
 sg13g2_nand3_1 _2368_ (.B(_0365_),
    .C(_0366_),
    .A(_1209_),
    .Y(_0367_));
 sg13g2_a21o_1 _2369_ (.A2(_1254_),
    .A1(_1186_),
    .B1(net495),
    .X(_0368_));
 sg13g2_a21oi_2 _2370_ (.B1(_1271_),
    .Y(_0369_),
    .A2(_1196_),
    .A1(_1113_));
 sg13g2_nand3_1 _2371_ (.B(_0368_),
    .C(_0369_),
    .A(_1218_),
    .Y(_0370_));
 sg13g2_nand4_1 _2372_ (.B(_0364_),
    .C(_0367_),
    .A(_0362_),
    .Y(_0371_),
    .D(_0370_));
 sg13g2_o21ai_1 _2373_ (.B1(_1206_),
    .Y(_0372_),
    .A1(_0358_),
    .A2(_0371_));
 sg13g2_nor2b_1 _2374_ (.A(_0357_),
    .B_N(net553),
    .Y(_0373_));
 sg13g2_nand3_1 _2375_ (.B(_0365_),
    .C(_0366_),
    .A(_1143_),
    .Y(_0374_));
 sg13g2_nand2b_1 _2376_ (.Y(_0375_),
    .B(net551),
    .A_N(_0363_));
 sg13g2_nand3_1 _2377_ (.B(_0368_),
    .C(_0369_),
    .A(_1181_),
    .Y(_0376_));
 sg13g2_o21ai_1 _2378_ (.B1(_1189_),
    .Y(_0377_),
    .A1(_0359_),
    .A2(_0361_));
 sg13g2_nand4_1 _2379_ (.B(_0375_),
    .C(_0376_),
    .A(_0374_),
    .Y(_0378_),
    .D(_0377_));
 sg13g2_o21ai_1 _2380_ (.B1(_0791_),
    .Y(_0379_),
    .A1(_0373_),
    .A2(_0378_));
 sg13g2_nor2b_1 _2381_ (.A(_0357_),
    .B_N(net545),
    .Y(_0380_));
 sg13g2_o21ai_1 _2382_ (.B1(_1240_),
    .Y(_0381_),
    .A1(_0359_),
    .A2(_0361_));
 sg13g2_nand3_1 _2383_ (.B(_0365_),
    .C(_0366_),
    .A(_1235_),
    .Y(_0382_));
 sg13g2_nand2b_1 _2384_ (.Y(_0383_),
    .B(_1231_),
    .A_N(_0363_));
 sg13g2_nand3_1 _2385_ (.B(_0368_),
    .C(_0369_),
    .A(_1242_),
    .Y(_0384_));
 sg13g2_nand4_1 _2386_ (.B(_0382_),
    .C(_0383_),
    .A(_0381_),
    .Y(_0385_),
    .D(_0384_));
 sg13g2_o21ai_1 _2387_ (.B1(_1228_),
    .Y(_0386_),
    .A1(_0380_),
    .A2(_0385_));
 sg13g2_and3_2 _2388_ (.X(_0387_),
    .A(_0372_),
    .B(_0379_),
    .C(_0386_));
 sg13g2_nand2_1 _2389_ (.Y(_0388_),
    .A(net514),
    .B(_0387_));
 sg13g2_nor2_1 _2390_ (.A(net514),
    .B(_0387_),
    .Y(_0389_));
 sg13g2_or2_1 _2391_ (.X(_0390_),
    .B(_0387_),
    .A(net514));
 sg13g2_xor2_1 _2392_ (.B(_0387_),
    .A(net514),
    .X(_0391_));
 sg13g2_xnor2_1 _2393_ (.Y(_0392_),
    .A(net514),
    .B(_0387_));
 sg13g2_nor2_1 _2394_ (.A(_0355_),
    .B(_0389_),
    .Y(_0393_));
 sg13g2_and3_1 _2395_ (.X(_0394_),
    .A(_0353_),
    .B(_0354_),
    .C(_0391_));
 sg13g2_nand3_1 _2396_ (.B(_0354_),
    .C(_0391_),
    .A(_0353_),
    .Y(_0395_));
 sg13g2_a21oi_1 _2397_ (.A1(_0087_),
    .A2(_0288_),
    .Y(_0396_),
    .B1(_0289_));
 sg13g2_nand2_1 _2398_ (.Y(_0397_),
    .A(_0353_),
    .B(_0388_));
 sg13g2_a22oi_1 _2399_ (.Y(_0398_),
    .B1(_0397_),
    .B2(_0354_),
    .A2(_0396_),
    .A1(_0394_));
 sg13g2_a21o_1 _2400_ (.A2(_0322_),
    .A1(_0317_),
    .B1(_1084_),
    .X(_0399_));
 sg13g2_or4_1 _2401_ (.A(_0087_),
    .B(_0088_),
    .C(_0287_),
    .D(_0289_),
    .X(_0400_));
 sg13g2_o21ai_1 _2402_ (.B1(_0399_),
    .Y(_0401_),
    .A1(_0395_),
    .A2(_0400_));
 sg13g2_nand2_1 _2403_ (.Y(_0402_),
    .A(_0323_),
    .B(_0399_));
 sg13g2_o21ai_1 _2404_ (.B1(_0323_),
    .Y(_0403_),
    .A1(_0398_),
    .A2(_0401_));
 sg13g2_a21oi_1 _2405_ (.A1(_0292_),
    .A2(_0403_),
    .Y(_0404_),
    .B1(_0744_));
 sg13g2_o21ai_1 _2406_ (.B1(_0404_),
    .Y(_0405_),
    .A1(_0292_),
    .A2(_0403_));
 sg13g2_a21oi_1 _2407_ (.A1(_0257_),
    .A2(_0405_),
    .Y(_0014_),
    .B1(_0667_));
 sg13g2_nor2b_1 _2408_ (.A(_0130_),
    .B_N(_0246_),
    .Y(_0406_));
 sg13g2_xnor2_1 _2409_ (.Y(_0407_),
    .A(_0130_),
    .B(_0246_));
 sg13g2_nor2b_1 _2410_ (.A(_0131_),
    .B_N(_0407_),
    .Y(_0408_));
 sg13g2_xor2_1 _2411_ (.B(_0407_),
    .A(_0131_),
    .X(_0409_));
 sg13g2_nor2_1 _2412_ (.A(_0255_),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_a21oi_1 _2413_ (.A1(_0787_),
    .A2(_1246_),
    .Y(_0411_),
    .B1(_0130_));
 sg13g2_nor2_1 _2414_ (.A(_0129_),
    .B(_0411_),
    .Y(_0412_));
 sg13g2_o21ai_1 _2415_ (.B1(_0246_),
    .Y(_0413_),
    .A1(_0129_),
    .A2(_0411_));
 sg13g2_xnor2_1 _2416_ (.Y(_0414_),
    .A(_0246_),
    .B(_0412_));
 sg13g2_a21o_1 _2417_ (.A2(_0414_),
    .A1(_0255_),
    .B1(_0743_),
    .X(_0415_));
 sg13g2_nor2_1 _2418_ (.A(_0287_),
    .B(_0392_),
    .Y(_0416_));
 sg13g2_nand2_1 _2419_ (.Y(_0417_),
    .A(_0288_),
    .B(_0391_));
 sg13g2_nand2_1 _2420_ (.Y(_0418_),
    .A(_0287_),
    .B(_0392_));
 sg13g2_and2_1 _2421_ (.A(_0417_),
    .B(_0418_),
    .X(_0419_));
 sg13g2_xor2_1 _2422_ (.B(_0419_),
    .A(_0291_),
    .X(_0420_));
 sg13g2_nor2b_1 _2423_ (.A(_0289_),
    .B_N(_0088_),
    .Y(_0421_));
 sg13g2_o21ai_1 _2424_ (.B1(_0392_),
    .Y(_0422_),
    .A1(_0287_),
    .A2(_0421_));
 sg13g2_o21ai_1 _2425_ (.B1(_0422_),
    .Y(_0423_),
    .A1(_0417_),
    .A2(_0421_));
 sg13g2_nor2_1 _2426_ (.A(_0403_),
    .B(_0423_),
    .Y(_0424_));
 sg13g2_a21oi_1 _2427_ (.A1(_0403_),
    .A2(_0420_),
    .Y(_0425_),
    .B1(_0424_));
 sg13g2_o21ai_1 _2428_ (.B1(net615),
    .Y(_0426_),
    .A1(_0410_),
    .A2(_0415_));
 sg13g2_a21oi_1 _2429_ (.A1(_0743_),
    .A2(_0425_),
    .Y(_0015_),
    .B1(_0426_));
 sg13g2_nand2_1 _2430_ (.Y(_0427_),
    .A(_0242_),
    .B(_0243_));
 sg13g2_nand2b_1 _2431_ (.Y(_0428_),
    .B(_0427_),
    .A_N(_0406_));
 sg13g2_nand2_1 _2432_ (.Y(_0429_),
    .A(_0245_),
    .B(_0427_));
 sg13g2_nor2_1 _2433_ (.A(_0406_),
    .B(_0408_),
    .Y(_0430_));
 sg13g2_xor2_1 _2434_ (.B(_0430_),
    .A(_0429_),
    .X(_0431_));
 sg13g2_nand2b_1 _2435_ (.Y(_0432_),
    .B(_0413_),
    .A_N(_0243_));
 sg13g2_xor2_1 _2436_ (.B(_0432_),
    .A(_0242_),
    .X(_0433_));
 sg13g2_a21oi_1 _2437_ (.A1(_0255_),
    .A2(_0433_),
    .Y(_0434_),
    .B1(_0743_));
 sg13g2_o21ai_1 _2438_ (.B1(_0434_),
    .Y(_0435_),
    .A1(_0255_),
    .A2(_0431_));
 sg13g2_o21ai_1 _2439_ (.B1(_0390_),
    .Y(_0436_),
    .A1(_0417_),
    .A2(_0421_));
 sg13g2_xnor2_1 _2440_ (.Y(_0437_),
    .A(_0355_),
    .B(_0436_));
 sg13g2_xnor2_1 _2441_ (.Y(_0438_),
    .A(_0355_),
    .B(_0390_));
 sg13g2_a21oi_1 _2442_ (.A1(_0291_),
    .A2(_0418_),
    .Y(_0439_),
    .B1(_0416_));
 sg13g2_a221oi_1 _2443_ (.B2(_0291_),
    .C1(_0416_),
    .B1(_0418_),
    .A1(_0355_),
    .Y(_0440_),
    .A2(_0389_));
 sg13g2_xnor2_1 _2444_ (.Y(_0441_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_mux2_1 _2445_ (.A0(_0437_),
    .A1(_0441_),
    .S(_0403_),
    .X(_0442_));
 sg13g2_nand2_1 _2446_ (.Y(_0443_),
    .A(_0743_),
    .B(_0442_));
 sg13g2_a21oi_1 _2447_ (.A1(_0435_),
    .A2(_0443_),
    .Y(_0016_),
    .B1(_0667_));
 sg13g2_o21ai_1 _2448_ (.B1(_0245_),
    .Y(_0444_),
    .A1(_0408_),
    .A2(_0428_));
 sg13g2_nor2_1 _2449_ (.A(_0168_),
    .B(_0252_),
    .Y(_0445_));
 sg13g2_xnor2_1 _2450_ (.Y(_0446_),
    .A(_0240_),
    .B(_0445_));
 sg13g2_xnor2_1 _2451_ (.Y(_0447_),
    .A(_0444_),
    .B(_0446_));
 sg13g2_nand2b_1 _2452_ (.Y(_0448_),
    .B(_0447_),
    .A_N(_0255_));
 sg13g2_o21ai_1 _2453_ (.B1(_0240_),
    .Y(_0449_),
    .A1(_0241_),
    .A2(_0432_));
 sg13g2_xnor2_1 _2454_ (.Y(_0450_),
    .A(_0445_),
    .B(_0449_));
 sg13g2_a21oi_1 _2455_ (.A1(_0255_),
    .A2(_0450_),
    .Y(_0451_),
    .B1(_0743_));
 sg13g2_nor2_1 _2456_ (.A(_0393_),
    .B(_0440_),
    .Y(_0452_));
 sg13g2_xnor2_1 _2457_ (.Y(_0453_),
    .A(_0353_),
    .B(_0402_));
 sg13g2_xnor2_1 _2458_ (.Y(_0454_),
    .A(_0452_),
    .B(_0453_));
 sg13g2_nand2_1 _2459_ (.Y(_0455_),
    .A(_0353_),
    .B(_0436_));
 sg13g2_a21oi_1 _2460_ (.A1(_0354_),
    .A2(_0455_),
    .Y(_0456_),
    .B1(_0399_));
 sg13g2_a21oi_1 _2461_ (.A1(_0403_),
    .A2(_0454_),
    .Y(_0457_),
    .B1(_0456_));
 sg13g2_a221oi_1 _2462_ (.B2(_0743_),
    .C1(_0667_),
    .B1(_0457_),
    .A1(_0448_),
    .Y(_0017_),
    .A2(_0451_));
 sg13g2_nand3_1 _2463_ (.B(_0642_),
    .C(_0739_),
    .A(_0641_),
    .Y(_0458_));
 sg13g2_nor2_2 _2464_ (.A(_0009_),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_and2_1 _2465_ (.A(net525),
    .B(_0459_),
    .X(_0460_));
 sg13g2_nand2_1 _2466_ (.Y(_0461_),
    .A(net525),
    .B(_0459_));
 sg13g2_o21ai_1 _2467_ (.B1(net610),
    .Y(_0462_),
    .A1(net140),
    .A2(_0460_));
 sg13g2_a21oi_1 _2468_ (.A1(net512),
    .A2(_0460_),
    .Y(_0018_),
    .B1(_0462_));
 sg13g2_a21oi_1 _2469_ (.A1(net138),
    .A2(_0461_),
    .Y(_0463_),
    .B1(_0667_));
 sg13g2_o21ai_1 _2470_ (.B1(_0463_),
    .Y(_0019_),
    .A1(net513),
    .A2(_0461_));
 sg13g2_o21ai_1 _2471_ (.B1(net610),
    .Y(_0464_),
    .A1(net95),
    .A2(_0460_));
 sg13g2_a21oi_1 _2472_ (.A1(_0987_),
    .A2(_0460_),
    .Y(_0020_),
    .B1(_0464_));
 sg13g2_nor2b_1 _2473_ (.A(_0746_),
    .B_N(net525),
    .Y(_0465_));
 sg13g2_o21ai_1 _2474_ (.B1(net613),
    .Y(_0466_),
    .A1(net117),
    .A2(net520));
 sg13g2_a21oi_1 _2475_ (.A1(_0951_),
    .A2(net520),
    .Y(_0021_),
    .B1(_0466_));
 sg13g2_o21ai_1 _2476_ (.B1(net613),
    .Y(_0467_),
    .A1(net106),
    .A2(net520));
 sg13g2_a21oi_1 _2477_ (.A1(net513),
    .A2(net520),
    .Y(_0022_),
    .B1(_0467_));
 sg13g2_o21ai_1 _2478_ (.B1(net613),
    .Y(_0468_),
    .A1(net103),
    .A2(net520));
 sg13g2_a21oi_1 _2479_ (.A1(_0987_),
    .A2(net520),
    .Y(_0023_),
    .B1(_0468_));
 sg13g2_o21ai_1 _2480_ (.B1(net614),
    .Y(_0469_),
    .A1(net113),
    .A2(_0465_));
 sg13g2_a21oi_1 _2481_ (.A1(_1032_),
    .A2(_0465_),
    .Y(_0024_),
    .B1(_0469_));
 sg13g2_o21ai_1 _2482_ (.B1(net615),
    .Y(_0470_),
    .A1(net96),
    .A2(net520));
 sg13g2_a21oi_1 _2483_ (.A1(_1075_),
    .A2(net520),
    .Y(_0025_),
    .B1(_0470_));
 sg13g2_nand3_1 _2484_ (.B(_0009_),
    .C(_0668_),
    .A(net569),
    .Y(_0471_));
 sg13g2_nand2_1 _2485_ (.Y(_0472_),
    .A(_0762_),
    .B(_0471_));
 sg13g2_nor2_1 _2486_ (.A(net571),
    .B(_0754_),
    .Y(_0473_));
 sg13g2_a221oi_1 _2487_ (.B2(_0010_),
    .C1(_0747_),
    .B1(_0473_),
    .A1(_0641_),
    .Y(_0474_),
    .A2(_0472_));
 sg13g2_nor2b_1 _2488_ (.A(_0474_),
    .B_N(net525),
    .Y(_0475_));
 sg13g2_nor2_1 _2489_ (.A(_0748_),
    .B(_0951_),
    .Y(_0476_));
 sg13g2_a21oi_2 _2490_ (.B1(_0476_),
    .Y(_0477_),
    .A2(_0782_),
    .A1(_0748_));
 sg13g2_o21ai_1 _2491_ (.B1(net612),
    .Y(_0478_),
    .A1(net101),
    .A2(_0475_));
 sg13g2_a21oi_1 _2492_ (.A1(_0475_),
    .A2(_0477_),
    .Y(_0026_),
    .B1(_0478_));
 sg13g2_and4_1 _2493_ (.A(_0881_),
    .B(_0890_),
    .C(_0901_),
    .D(_0904_),
    .X(_0479_));
 sg13g2_a21oi_2 _2494_ (.B1(_0747_),
    .Y(_0480_),
    .A2(_0479_),
    .A1(_0783_));
 sg13g2_xor2_1 _2495_ (.B(_0881_),
    .A(_0782_),
    .X(_0481_));
 sg13g2_a22oi_1 _2496_ (.Y(_0482_),
    .B1(_0480_),
    .B2(_0481_),
    .A2(_0879_),
    .A1(_0747_));
 sg13g2_o21ai_1 _2497_ (.B1(net612),
    .Y(_0483_),
    .A1(net97),
    .A2(net519));
 sg13g2_a21oi_1 _2498_ (.A1(net519),
    .A2(_0482_),
    .Y(_0027_),
    .B1(_0483_));
 sg13g2_nor3_2 _2499_ (.A(_0782_),
    .B(_0881_),
    .C(_0904_),
    .Y(_0484_));
 sg13g2_o21ai_1 _2500_ (.B1(_0904_),
    .Y(_0485_),
    .A1(_0782_),
    .A2(_0881_));
 sg13g2_nor2b_1 _2501_ (.A(_0484_),
    .B_N(_0485_),
    .Y(_0486_));
 sg13g2_a22oi_1 _2502_ (.Y(_0487_),
    .B1(_0480_),
    .B2(_0486_),
    .A2(_0988_),
    .A1(_0747_));
 sg13g2_o21ai_1 _2503_ (.B1(net612),
    .Y(_0488_),
    .A1(net98),
    .A2(net519));
 sg13g2_a21oi_1 _2504_ (.A1(net519),
    .A2(_0487_),
    .Y(_0028_),
    .B1(_0488_));
 sg13g2_nand2_1 _2505_ (.Y(_0489_),
    .A(_0901_),
    .B(_0484_));
 sg13g2_xnor2_1 _2506_ (.Y(_0490_),
    .A(_0900_),
    .B(_0484_));
 sg13g2_a22oi_1 _2507_ (.Y(_0491_),
    .B1(_0480_),
    .B2(_0490_),
    .A2(_1033_),
    .A1(_0747_));
 sg13g2_o21ai_1 _2508_ (.B1(net609),
    .Y(_0492_),
    .A1(net100),
    .A2(net519));
 sg13g2_a21oi_1 _2509_ (.A1(net519),
    .A2(_0491_),
    .Y(_0029_),
    .B1(_0492_));
 sg13g2_xnor2_1 _2510_ (.Y(_0493_),
    .A(_0890_),
    .B(_0489_));
 sg13g2_a22oi_1 _2511_ (.Y(_0494_),
    .B1(_0480_),
    .B2(_0493_),
    .A2(_1076_),
    .A1(_0747_));
 sg13g2_o21ai_1 _2512_ (.B1(net609),
    .Y(_0495_),
    .A1(net115),
    .A2(net519));
 sg13g2_a21oi_1 _2513_ (.A1(net519),
    .A2(_0494_),
    .Y(_0030_),
    .B1(_0495_));
 sg13g2_and2_1 _2514_ (.A(net523),
    .B(_0459_),
    .X(_0496_));
 sg13g2_nand2_1 _2515_ (.Y(_0497_),
    .A(net523),
    .B(_0459_));
 sg13g2_a21oi_1 _2516_ (.A1(net579),
    .A2(_0497_),
    .Y(_0498_),
    .B1(_0667_));
 sg13g2_o21ai_1 _2517_ (.B1(_0498_),
    .Y(_0031_),
    .A1(net512),
    .A2(_0497_));
 sg13g2_o21ai_1 _2518_ (.B1(net610),
    .Y(_0499_),
    .A1(net143),
    .A2(_0496_));
 sg13g2_a21oi_1 _2519_ (.A1(net513),
    .A2(_0496_),
    .Y(_0032_),
    .B1(_0499_));
 sg13g2_o21ai_1 _2520_ (.B1(net610),
    .Y(_0500_),
    .A1(net128),
    .A2(_0496_));
 sg13g2_a21oi_1 _2521_ (.A1(_0987_),
    .A2(_0496_),
    .Y(_0033_),
    .B1(_0500_));
 sg13g2_nor2_1 _2522_ (.A(_0746_),
    .B(_0778_),
    .Y(_0501_));
 sg13g2_o21ai_1 _2523_ (.B1(net613),
    .Y(_0502_),
    .A1(net111),
    .A2(net518));
 sg13g2_a21oi_1 _2524_ (.A1(net512),
    .A2(net518),
    .Y(_0034_),
    .B1(_0502_));
 sg13g2_o21ai_1 _2525_ (.B1(net612),
    .Y(_0503_),
    .A1(net102),
    .A2(net518));
 sg13g2_a21oi_1 _2526_ (.A1(net513),
    .A2(net518),
    .Y(_0035_),
    .B1(_0503_));
 sg13g2_o21ai_1 _2527_ (.B1(net613),
    .Y(_0504_),
    .A1(net104),
    .A2(net518));
 sg13g2_a21oi_1 _2528_ (.A1(_0987_),
    .A2(net518),
    .Y(_0036_),
    .B1(_0504_));
 sg13g2_o21ai_1 _2529_ (.B1(net614),
    .Y(_0505_),
    .A1(net99),
    .A2(_0501_));
 sg13g2_a21oi_1 _2530_ (.A1(_1032_),
    .A2(_0501_),
    .Y(_0037_),
    .B1(_0505_));
 sg13g2_o21ai_1 _2531_ (.B1(net612),
    .Y(_0506_),
    .A1(net107),
    .A2(net518));
 sg13g2_a21oi_1 _2532_ (.A1(_1075_),
    .A2(net518),
    .Y(_0038_),
    .B1(_0506_));
 sg13g2_nor2_1 _2533_ (.A(_0778_),
    .B(_0474_),
    .Y(_0507_));
 sg13g2_o21ai_1 _2534_ (.B1(net612),
    .Y(_0508_),
    .A1(net133),
    .A2(net517));
 sg13g2_a21oi_1 _2535_ (.A1(_0477_),
    .A2(net517),
    .Y(_0039_),
    .B1(_0508_));
 sg13g2_o21ai_1 _2536_ (.B1(net609),
    .Y(_0509_),
    .A1(net124),
    .A2(net517));
 sg13g2_a21oi_1 _2537_ (.A1(_0482_),
    .A2(net517),
    .Y(_0040_),
    .B1(_0509_));
 sg13g2_o21ai_1 _2538_ (.B1(net611),
    .Y(_0510_),
    .A1(net121),
    .A2(_0507_));
 sg13g2_a21oi_1 _2539_ (.A1(_0487_),
    .A2(_0507_),
    .Y(_0041_),
    .B1(_0510_));
 sg13g2_o21ai_1 _2540_ (.B1(net611),
    .Y(_0511_),
    .A1(net120),
    .A2(net517));
 sg13g2_a21oi_1 _2541_ (.A1(_0491_),
    .A2(net517),
    .Y(_0042_),
    .B1(_0511_));
 sg13g2_o21ai_1 _2542_ (.B1(net609),
    .Y(_0512_),
    .A1(net110),
    .A2(net517));
 sg13g2_a21oi_1 _2543_ (.A1(_0494_),
    .A2(net517),
    .Y(_0043_),
    .B1(_0512_));
 sg13g2_and2_2 _2544_ (.A(net522),
    .B(_0459_),
    .X(_0513_));
 sg13g2_o21ai_1 _2545_ (.B1(net610),
    .Y(_0514_),
    .A1(net578),
    .A2(_0513_));
 sg13g2_a21oi_1 _2546_ (.A1(net512),
    .A2(_0513_),
    .Y(_0044_),
    .B1(_0514_));
 sg13g2_o21ai_1 _2547_ (.B1(net610),
    .Y(_0515_),
    .A1(net577),
    .A2(_0513_));
 sg13g2_a21oi_1 _2548_ (.A1(net513),
    .A2(_0513_),
    .Y(_0045_),
    .B1(_0515_));
 sg13g2_o21ai_1 _2549_ (.B1(net610),
    .Y(_0516_),
    .A1(net132),
    .A2(_0513_));
 sg13g2_a21oi_1 _2550_ (.A1(_0987_),
    .A2(_0513_),
    .Y(_0046_),
    .B1(_0516_));
 sg13g2_nor2_1 _2551_ (.A(_0746_),
    .B(_0780_),
    .Y(_0517_));
 sg13g2_o21ai_1 _2552_ (.B1(net613),
    .Y(_0518_),
    .A1(net114),
    .A2(net516));
 sg13g2_a21oi_1 _2553_ (.A1(net512),
    .A2(net516),
    .Y(_0047_),
    .B1(_0518_));
 sg13g2_o21ai_1 _2554_ (.B1(net612),
    .Y(_0519_),
    .A1(net118),
    .A2(net516));
 sg13g2_a21oi_1 _2555_ (.A1(net513),
    .A2(net516),
    .Y(_0048_),
    .B1(_0519_));
 sg13g2_o21ai_1 _2556_ (.B1(net613),
    .Y(_0520_),
    .A1(net112),
    .A2(net516));
 sg13g2_a21oi_1 _2557_ (.A1(_0987_),
    .A2(net516),
    .Y(_0049_),
    .B1(_0520_));
 sg13g2_o21ai_1 _2558_ (.B1(net614),
    .Y(_0521_),
    .A1(net116),
    .A2(_0517_));
 sg13g2_a21oi_1 _2559_ (.A1(_1032_),
    .A2(_0517_),
    .Y(_0050_),
    .B1(_0521_));
 sg13g2_o21ai_1 _2560_ (.B1(net613),
    .Y(_0522_),
    .A1(net105),
    .A2(net516));
 sg13g2_a21oi_1 _2561_ (.A1(_1075_),
    .A2(net516),
    .Y(_0051_),
    .B1(_0522_));
 sg13g2_nor2_1 _2562_ (.A(_0780_),
    .B(_0474_),
    .Y(_0523_));
 sg13g2_o21ai_1 _2563_ (.B1(net612),
    .Y(_0524_),
    .A1(net129),
    .A2(_0523_));
 sg13g2_a21oi_1 _2564_ (.A1(_0477_),
    .A2(_0523_),
    .Y(_0052_),
    .B1(_0524_));
 sg13g2_o21ai_1 _2565_ (.B1(net609),
    .Y(_0525_),
    .A1(net126),
    .A2(net515));
 sg13g2_a21oi_1 _2566_ (.A1(_0482_),
    .A2(net515),
    .Y(_0053_),
    .B1(_0525_));
 sg13g2_o21ai_1 _2567_ (.B1(net609),
    .Y(_0526_),
    .A1(net125),
    .A2(net515));
 sg13g2_a21oi_1 _2568_ (.A1(_0487_),
    .A2(net515),
    .Y(_0054_),
    .B1(_0526_));
 sg13g2_o21ai_1 _2569_ (.B1(net609),
    .Y(_0527_),
    .A1(net123),
    .A2(net515));
 sg13g2_a21oi_1 _2570_ (.A1(_0491_),
    .A2(net515),
    .Y(_0055_),
    .B1(_0527_));
 sg13g2_o21ai_1 _2571_ (.B1(net609),
    .Y(_0528_),
    .A1(net122),
    .A2(net515));
 sg13g2_a21oi_1 _2572_ (.A1(_0494_),
    .A2(net515),
    .Y(_0056_),
    .B1(_0528_));
 sg13g2_nand2_1 _2573_ (.Y(_0529_),
    .A(_0647_),
    .B(net597));
 sg13g2_nand2_1 _2574_ (.Y(_0530_),
    .A(\enigma.plugboard.cnt[0] ),
    .B(_0652_));
 sg13g2_xor2_1 _2575_ (.B(net593),
    .A(\enigma.plugboard.cnt[3] ),
    .X(_0531_));
 sg13g2_a221oi_1 _2576_ (.B2(net606),
    .C1(_0531_),
    .B1(_0651_),
    .A1(\enigma.plugboard.cnt[4] ),
    .Y(_0532_),
    .A2(_0645_));
 sg13g2_a22oi_1 _2577_ (.Y(_0533_),
    .B1(_0649_),
    .B2(net602),
    .A2(_0648_),
    .A1(\enigma.plugboard.cnt[2] ));
 sg13g2_a22oi_1 _2578_ (.Y(_0534_),
    .B1(\enigma.plugboard.cnt[1] ),
    .B2(_0650_),
    .A2(net589),
    .A1(_0644_));
 sg13g2_and4_1 _2579_ (.A(_0530_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .X(_0535_));
 sg13g2_a21oi_1 _2580_ (.A1(_0529_),
    .A2(_0535_),
    .Y(_0536_),
    .B1(_0721_));
 sg13g2_o21ai_1 _2581_ (.B1(net617),
    .Y(_0537_),
    .A1(\enigma.plugboard.plug_limiter[0] ),
    .A2(_0536_));
 sg13g2_a21oi_1 _2582_ (.A1(_0653_),
    .A2(_0536_),
    .Y(_0057_),
    .B1(_0537_));
 sg13g2_and2_1 _2583_ (.A(\enigma.plugboard.plug_limiter[0] ),
    .B(_0536_),
    .X(_0538_));
 sg13g2_o21ai_1 _2584_ (.B1(net617),
    .Y(_0539_),
    .A1(net91),
    .A2(_0538_));
 sg13g2_a21oi_1 _2585_ (.A1(net91),
    .A2(_0538_),
    .Y(_0058_),
    .B1(_0539_));
 sg13g2_a21oi_1 _2586_ (.A1(\enigma.plugboard.plug_limiter[1] ),
    .A2(_0538_),
    .Y(_0540_),
    .B1(net87));
 sg13g2_nor2_1 _2587_ (.A(_0667_),
    .B(net88),
    .Y(_0059_));
 sg13g2_and2_1 _2588_ (.A(net85),
    .B(net617),
    .X(_0060_));
 sg13g2_and2_1 _2589_ (.A(net86),
    .B(net617),
    .X(_0061_));
 sg13g2_nand3_1 _2590_ (.B(_0668_),
    .C(_0718_),
    .A(net566),
    .Y(_0541_));
 sg13g2_o21ai_1 _2591_ (.B1(net616),
    .Y(_0542_),
    .A1(net606),
    .A2(net543));
 sg13g2_a21oi_1 _2592_ (.A1(_0651_),
    .A2(net543),
    .Y(_0062_),
    .B1(_0542_));
 sg13g2_o21ai_1 _2593_ (.B1(net616),
    .Y(_0543_),
    .A1(net603),
    .A2(net543));
 sg13g2_a21oi_1 _2594_ (.A1(_0649_),
    .A2(net543),
    .Y(_0063_),
    .B1(_0543_));
 sg13g2_o21ai_1 _2595_ (.B1(net617),
    .Y(_0544_),
    .A1(net597),
    .A2(net543));
 sg13g2_a21oi_1 _2596_ (.A1(_0647_),
    .A2(net543),
    .Y(_0064_),
    .B1(_0544_));
 sg13g2_o21ai_1 _2597_ (.B1(net616),
    .Y(_0545_),
    .A1(net593),
    .A2(net543));
 sg13g2_a21oi_1 _2598_ (.A1(_0646_),
    .A2(net544),
    .Y(_0065_),
    .B1(_0545_));
 sg13g2_o21ai_1 _2599_ (.B1(net616),
    .Y(_0546_),
    .A1(net589),
    .A2(net543));
 sg13g2_a21oi_1 _2600_ (.A1(_0644_),
    .A2(net544),
    .Y(_0066_),
    .B1(_0546_));
 sg13g2_nor2_1 _2601_ (.A(_1223_),
    .B(_1224_),
    .Y(_0547_));
 sg13g2_a21oi_1 _2602_ (.A1(\enigma.r.$signal$17[2] ),
    .A2(net577),
    .Y(_0548_),
    .B1(net578));
 sg13g2_o21ai_1 _2603_ (.B1(_0548_),
    .Y(_0549_),
    .A1(\enigma.r.$signal$17[2] ),
    .A2(net576));
 sg13g2_xnor2_1 _2604_ (.Y(_0550_),
    .A(\enigma.r.cnts_debug0[2] ),
    .B(_0547_));
 sg13g2_o21ai_1 _2605_ (.B1(_0550_),
    .Y(_0551_),
    .A1(\enigma.r.cnts_debug0[4] ),
    .A2(_0549_));
 sg13g2_nand2_1 _2606_ (.Y(_0552_),
    .A(\enigma.r.cnts_debug0[0] ),
    .B(_1232_));
 sg13g2_a21oi_1 _2607_ (.A1(_1226_),
    .A2(_0552_),
    .Y(_0553_),
    .B1(\enigma.r.cnts_debug0[3] ));
 sg13g2_o21ai_1 _2608_ (.B1(\enigma.r.cnts_debug0[3] ),
    .Y(_0554_),
    .A1(_0654_),
    .A2(_1226_));
 sg13g2_a221oi_1 _2609_ (.B2(\enigma.r.cnts_debug0[4] ),
    .C1(\enigma.r.cnts_debug0[1] ),
    .B1(_0549_),
    .A1(_0654_),
    .Y(_0555_),
    .A2(net547));
 sg13g2_nand2_1 _2610_ (.Y(_0556_),
    .A(_0554_),
    .B(_0555_));
 sg13g2_or3_2 _2611_ (.A(_0551_),
    .B(_0553_),
    .C(_0556_),
    .X(_0557_));
 sg13g2_nand2_1 _2612_ (.Y(_0558_),
    .A(net89),
    .B(_0557_));
 sg13g2_nand3_1 _2613_ (.B(_0739_),
    .C(_0760_),
    .A(net565),
    .Y(_0559_));
 sg13g2_o21ai_1 _2614_ (.B1(_0458_),
    .Y(_0560_),
    .A1(_0641_),
    .A2(_0672_));
 sg13g2_nand3_1 _2615_ (.B(_0748_),
    .C(_0559_),
    .A(_0746_),
    .Y(_0561_));
 sg13g2_or2_1 _2616_ (.X(_0562_),
    .B(_0561_),
    .A(_0560_));
 sg13g2_nand4_1 _2617_ (.B(net573),
    .C(_0643_),
    .A(net567),
    .Y(_0563_),
    .D(_0669_));
 sg13g2_nor2_1 _2618_ (.A(net89),
    .B(_0563_),
    .Y(_0564_));
 sg13g2_nor4_2 _2619_ (.A(net573),
    .B(net575),
    .C(net565),
    .Y(_0565_),
    .D(_0670_));
 sg13g2_inv_1 _2620_ (.Y(_0566_),
    .A(_0565_));
 sg13g2_o21ai_1 _2621_ (.B1(_0757_),
    .Y(_0567_),
    .A1(_0642_),
    .A2(_0717_));
 sg13g2_nor4_1 _2622_ (.A(_0562_),
    .B(_0564_),
    .C(_0565_),
    .D(_0567_),
    .Y(_0568_));
 sg13g2_a21oi_1 _2623_ (.A1(_0717_),
    .A2(_0769_),
    .Y(_0569_),
    .B1(_0740_));
 sg13g2_nand3_1 _2624_ (.B(_0718_),
    .C(_0739_),
    .A(net567),
    .Y(_0570_));
 sg13g2_nor2b_1 _2625_ (.A(_0755_),
    .B_N(_0570_),
    .Y(_0571_));
 sg13g2_nand2b_1 _2626_ (.Y(_0572_),
    .B(_0571_),
    .A_N(_0569_));
 sg13g2_nand2_1 _2627_ (.Y(_0573_),
    .A(_0757_),
    .B(_0771_));
 sg13g2_nor3_1 _2628_ (.A(_0719_),
    .B(_0572_),
    .C(_0573_),
    .Y(_0574_));
 sg13g2_nand3_1 _2629_ (.B(net544),
    .C(_0574_),
    .A(_0764_),
    .Y(_0575_));
 sg13g2_nand2_1 _2630_ (.Y(_0576_),
    .A(_0759_),
    .B(_0770_));
 sg13g2_nand4_1 _2631_ (.B(_0770_),
    .C(_0563_),
    .A(_0759_),
    .Y(_0577_),
    .D(_0566_));
 sg13g2_nor3_2 _2632_ (.A(_0562_),
    .B(_0575_),
    .C(_0577_),
    .Y(_0578_));
 sg13g2_nor2_1 _2633_ (.A(net2),
    .B(net4),
    .Y(_0579_));
 sg13g2_nand2b_1 _2634_ (.Y(_0580_),
    .B(net4),
    .A_N(net3));
 sg13g2_nor2b_1 _2635_ (.A(_0579_),
    .B_N(_0580_),
    .Y(_0581_));
 sg13g2_a21oi_1 _2636_ (.A1(_0671_),
    .A2(_0581_),
    .Y(_0582_),
    .B1(_0643_));
 sg13g2_a22oi_1 _2637_ (.Y(_0583_),
    .B1(_0578_),
    .B2(_0582_),
    .A2(_0558_),
    .A1(_0763_));
 sg13g2_a21oi_1 _2638_ (.A1(_0568_),
    .A2(_0583_),
    .Y(_0067_),
    .B1(_0667_));
 sg13g2_nand2_1 _2639_ (.Y(_0584_),
    .A(\enigma.r.cnts_debug1[0] ),
    .B(_1215_));
 sg13g2_a21oi_1 _2640_ (.A1(_1205_),
    .A2(_0584_),
    .Y(_0585_),
    .B1(\enigma.r.cnts_debug1[3] ));
 sg13g2_o21ai_1 _2641_ (.B1(\enigma.r.cnts_debug1[3] ),
    .Y(_0586_),
    .A1(_0656_),
    .A2(_1205_));
 sg13g2_nor2b_1 _2642_ (.A(_0585_),
    .B_N(_0586_),
    .Y(_0587_));
 sg13g2_a21oi_1 _2643_ (.A1(\enigma.r.$signal$21[2] ),
    .A2(\enigma.r.$signal$21[1] ),
    .Y(_0588_),
    .B1(\enigma.r.$signal$21[0] ));
 sg13g2_o21ai_1 _2644_ (.B1(_0588_),
    .Y(_0589_),
    .A1(\enigma.r.$signal$21[2] ),
    .A2(_0001_));
 sg13g2_xnor2_1 _2645_ (.Y(_0590_),
    .A(_0655_),
    .B(_0589_));
 sg13g2_o21ai_1 _2646_ (.B1(\enigma.r.cnts_debug1[2] ),
    .Y(_0591_),
    .A1(_1202_),
    .A2(_1203_));
 sg13g2_nor3_1 _2647_ (.A(\enigma.r.cnts_debug1[2] ),
    .B(_1202_),
    .C(_1203_),
    .Y(_0592_));
 sg13g2_nor2_1 _2648_ (.A(\enigma.r.cnts_debug1[0] ),
    .B(_1215_),
    .Y(_0593_));
 sg13g2_nor3_1 _2649_ (.A(\enigma.r.cnts_debug1[1] ),
    .B(_0592_),
    .C(_0593_),
    .Y(_0594_));
 sg13g2_nand4_1 _2650_ (.B(_0590_),
    .C(_0591_),
    .A(_0587_),
    .Y(_0595_),
    .D(_0594_));
 sg13g2_nor2_1 _2651_ (.A(\enigma.fsm.double_step ),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_nand2b_1 _2652_ (.Y(_0597_),
    .B(_0770_),
    .A_N(_0572_));
 sg13g2_nand3b_1 _2653_ (.B(_0763_),
    .C(_0557_),
    .Y(_0598_),
    .A_N(\enigma.fsm.double_step ));
 sg13g2_o21ai_1 _2654_ (.B1(_0598_),
    .Y(_0599_),
    .A1(_0563_),
    .A2(_0596_));
 sg13g2_nor4_1 _2655_ (.A(_0761_),
    .B(_0578_),
    .C(_0597_),
    .D(_0599_),
    .Y(_0600_));
 sg13g2_nand2_1 _2656_ (.Y(_0601_),
    .A(_0672_),
    .B(_0578_));
 sg13g2_nor2_1 _2657_ (.A(net3),
    .B(net4),
    .Y(_0602_));
 sg13g2_xor2_1 _2658_ (.B(_0602_),
    .A(net2),
    .X(_0603_));
 sg13g2_o21ai_1 _2659_ (.B1(_0578_),
    .Y(_0604_),
    .A1(_0672_),
    .A2(_0603_));
 sg13g2_o21ai_1 _2660_ (.B1(net615),
    .Y(_0605_),
    .A1(net574),
    .A2(_0604_));
 sg13g2_nor2_1 _2661_ (.A(_0600_),
    .B(_0605_),
    .Y(_0068_));
 sg13g2_nor2_1 _2662_ (.A(_0563_),
    .B(_0595_),
    .Y(_0606_));
 sg13g2_nand2_1 _2663_ (.Y(_0607_),
    .A(net89),
    .B(_0606_));
 sg13g2_nor3_1 _2664_ (.A(_0569_),
    .B(_0573_),
    .C(_0578_),
    .Y(_0608_));
 sg13g2_nor2_1 _2665_ (.A(net4),
    .B(_0672_),
    .Y(_0609_));
 sg13g2_o21ai_1 _2666_ (.B1(net615),
    .Y(_0610_),
    .A1(net572),
    .A2(_0601_));
 sg13g2_a221oi_1 _2667_ (.B2(_0578_),
    .C1(_0610_),
    .B1(_0609_),
    .A1(_0607_),
    .Y(_0069_),
    .A2(_0608_));
 sg13g2_nor2_1 _2668_ (.A(net137),
    .B(_0563_),
    .Y(_0611_));
 sg13g2_a221oi_1 _2669_ (.B2(_0611_),
    .C1(_0575_),
    .B1(_0595_),
    .A1(net569),
    .Y(_0612_),
    .A2(_0578_));
 sg13g2_nor2_1 _2670_ (.A(_0667_),
    .B(_0612_),
    .Y(_0070_));
 sg13g2_nor4_1 _2671_ (.A(_0564_),
    .B(_0565_),
    .C(_0576_),
    .D(_0606_),
    .Y(_0613_));
 sg13g2_o21ai_1 _2672_ (.B1(net615),
    .Y(_0614_),
    .A1(net567),
    .A2(_0601_));
 sg13g2_a21oi_1 _2673_ (.A1(_0601_),
    .A2(_0613_),
    .Y(_0071_),
    .B1(_0614_));
 sg13g2_o21ai_1 _2674_ (.B1(net137),
    .Y(_0615_),
    .A1(net571),
    .A2(_0458_));
 sg13g2_o21ai_1 _2675_ (.B1(_0570_),
    .Y(_0616_),
    .A1(_0755_),
    .A2(_0615_));
 sg13g2_and2_1 _2676_ (.A(net614),
    .B(_0616_),
    .X(_0072_));
 sg13g2_a22oi_1 _2677_ (.Y(_0617_),
    .B1(_0752_),
    .B2(net127),
    .A2(_0671_),
    .A1(_0641_));
 sg13g2_xnor2_1 _2678_ (.Y(_0618_),
    .A(net2),
    .B(net4));
 sg13g2_a221oi_1 _2679_ (.B2(net3),
    .C1(_0673_),
    .B1(_0618_),
    .A1(net2),
    .Y(_0619_),
    .A2(_0602_));
 sg13g2_nor2_1 _2680_ (.A(_0617_),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_a21oi_1 _2681_ (.A1(net575),
    .A2(_0620_),
    .Y(_0621_),
    .B1(net93));
 sg13g2_nand2_1 _2682_ (.Y(_0622_),
    .A(net93),
    .B(_0620_));
 sg13g2_nand2_1 _2683_ (.Y(_0623_),
    .A(net614),
    .B(_0622_));
 sg13g2_nor2_1 _2684_ (.A(net94),
    .B(_0623_),
    .Y(_0073_));
 sg13g2_xor2_1 _2685_ (.B(_0622_),
    .A(net127),
    .X(_0624_));
 sg13g2_o21ai_1 _2686_ (.B1(net614),
    .Y(_0625_),
    .A1(\enigma.fsm.ready ),
    .A2(_0617_));
 sg13g2_nor2_1 _2687_ (.A(_0624_),
    .B(_0625_),
    .Y(_0074_));
 sg13g2_or3_2 _2688_ (.A(net2),
    .B(_0566_),
    .C(_0580_),
    .X(_0626_));
 sg13g2_nor2_1 _2689_ (.A(_0942_),
    .B(_0626_),
    .Y(_0627_));
 sg13g2_nor3_2 _2690_ (.A(net2),
    .B(_0566_),
    .C(_0580_),
    .Y(_0628_));
 sg13g2_o21ai_1 _2691_ (.B1(net615),
    .Y(_0629_),
    .A1(uio_out[0]),
    .A2(_0628_));
 sg13g2_nor2_1 _2692_ (.A(_0627_),
    .B(_0629_),
    .Y(_0075_));
 sg13g2_nor2_1 _2693_ (.A(_0866_),
    .B(_0626_),
    .Y(_0630_));
 sg13g2_o21ai_1 _2694_ (.B1(net616),
    .Y(_0631_),
    .A1(net119),
    .A2(_0628_));
 sg13g2_nor2_1 _2695_ (.A(_0630_),
    .B(_0631_),
    .Y(_0076_));
 sg13g2_nor2_1 _2696_ (.A(_0977_),
    .B(_0626_),
    .Y(_0632_));
 sg13g2_o21ai_1 _2697_ (.B1(net615),
    .Y(_0633_),
    .A1(net560),
    .A2(_0628_));
 sg13g2_nor2_1 _2698_ (.A(_0632_),
    .B(_0633_),
    .Y(_0077_));
 sg13g2_nor2_1 _2699_ (.A(_1024_),
    .B(_0626_),
    .Y(_0634_));
 sg13g2_o21ai_1 _2700_ (.B1(net616),
    .Y(_0635_),
    .A1(net559),
    .A2(_0628_));
 sg13g2_nor2_1 _2701_ (.A(_0634_),
    .B(_0635_),
    .Y(_0078_));
 sg13g2_nor2_1 _2702_ (.A(_1070_),
    .B(_0626_),
    .Y(_0636_));
 sg13g2_o21ai_1 _2703_ (.B1(net616),
    .Y(_0637_),
    .A1(net556),
    .A2(_0628_));
 sg13g2_nor2_1 _2704_ (.A(_0636_),
    .B(_0637_),
    .Y(_0079_));
 sg13g2_dfrbp_1 _2705_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net14),
    .D(_0013_),
    .Q_N(_0011_),
    .Q(\enigma.r.dout[0] ));
 sg13g2_dfrbp_1 _2706_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net12),
    .D(_0014_),
    .Q_N(_0012_),
    .Q(\enigma.r.dout[1] ));
 sg13g2_dfrbp_1 _2707_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net11),
    .D(_0015_),
    .Q_N(_1334_),
    .Q(\enigma.r.dout[2] ));
 sg13g2_dfrbp_1 _2708_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net10),
    .D(_0016_),
    .Q_N(_1333_),
    .Q(\enigma.r.dout[3] ));
 sg13g2_dfrbp_1 _2709_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net9),
    .D(_0017_),
    .Q_N(_1332_),
    .Q(\enigma.r.dout[4] ));
 sg13g2_dfrbp_1 _2710_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net8),
    .D(_0018_),
    .Q_N(_1331_),
    .Q(\enigma.r.$signal$23[0] ));
 sg13g2_dfrbp_1 _2711_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net73),
    .D(net139),
    .Q_N(_1330_),
    .Q(\enigma.r.$signal$23[1] ));
 sg13g2_dfrbp_1 _2712_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net71),
    .D(_0020_),
    .Q_N(_0000_),
    .Q(\enigma.r.$signal$23[2] ));
 sg13g2_dfrbp_1 _2713_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net69),
    .D(_0021_),
    .Q_N(_1329_),
    .Q(\enigma.r.$signal$22[0] ));
 sg13g2_dfrbp_1 _2714_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net67),
    .D(_0022_),
    .Q_N(_1328_),
    .Q(\enigma.r.$signal$22[1] ));
 sg13g2_dfrbp_1 _2715_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net65),
    .D(_0023_),
    .Q_N(_1327_),
    .Q(\enigma.r.$signal$22[2] ));
 sg13g2_dfrbp_1 _2716_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net63),
    .D(_0024_),
    .Q_N(_1326_),
    .Q(\enigma.r.$signal$22[3] ));
 sg13g2_dfrbp_1 _2717_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net61),
    .D(_0025_),
    .Q_N(_1325_),
    .Q(\enigma.r.$signal$22[4] ));
 sg13g2_dfrbp_1 _2718_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net59),
    .D(_0026_),
    .Q_N(_1324_),
    .Q(\enigma.r.cnts_debug2[0] ));
 sg13g2_dfrbp_1 _2719_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net57),
    .D(_0027_),
    .Q_N(_1323_),
    .Q(\enigma.r.cnts_debug2[1] ));
 sg13g2_dfrbp_1 _2720_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net55),
    .D(_0028_),
    .Q_N(_1322_),
    .Q(\enigma.r.cnts_debug2[2] ));
 sg13g2_dfrbp_1 _2721_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net53),
    .D(_0029_),
    .Q_N(_1321_),
    .Q(\enigma.r.cnts_debug2[3] ));
 sg13g2_dfrbp_1 _2722_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net51),
    .D(_0030_),
    .Q_N(_1320_),
    .Q(\enigma.r.cnts_debug2[4] ));
 sg13g2_dfrbp_1 _2723_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net49),
    .D(net148),
    .Q_N(_1319_),
    .Q(\enigma.r.$signal$21[0] ));
 sg13g2_dfrbp_1 _2724_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net47),
    .D(_0032_),
    .Q_N(_1318_),
    .Q(\enigma.r.$signal$21[1] ));
 sg13g2_dfrbp_1 _2725_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net45),
    .D(_0033_),
    .Q_N(_0001_),
    .Q(\enigma.r.$signal$21[2] ));
 sg13g2_dfrbp_1 _2726_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net43),
    .D(_0034_),
    .Q_N(_1317_),
    .Q(\enigma.r.$signal$20[0] ));
 sg13g2_dfrbp_1 _2727_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net41),
    .D(_0035_),
    .Q_N(_1316_),
    .Q(\enigma.r.$signal$20[1] ));
 sg13g2_dfrbp_1 _2728_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net39),
    .D(_0036_),
    .Q_N(_1315_),
    .Q(\enigma.r.$signal$20[2] ));
 sg13g2_dfrbp_1 _2729_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net37),
    .D(_0037_),
    .Q_N(_1314_),
    .Q(\enigma.r.$signal$20[3] ));
 sg13g2_dfrbp_1 _2730_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net35),
    .D(_0038_),
    .Q_N(_1313_),
    .Q(\enigma.r.$signal$20[4] ));
 sg13g2_dfrbp_1 _2731_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net33),
    .D(_0039_),
    .Q_N(_1312_),
    .Q(\enigma.r.cnts_debug1[0] ));
 sg13g2_dfrbp_1 _2732_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net31),
    .D(_0040_),
    .Q_N(_1311_),
    .Q(\enigma.r.cnts_debug1[1] ));
 sg13g2_dfrbp_1 _2733_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net29),
    .D(_0041_),
    .Q_N(_1310_),
    .Q(\enigma.r.cnts_debug1[2] ));
 sg13g2_dfrbp_1 _2734_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net27),
    .D(_0042_),
    .Q_N(_1309_),
    .Q(\enigma.r.cnts_debug1[3] ));
 sg13g2_dfrbp_1 _2735_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net25),
    .D(_0043_),
    .Q_N(_1308_),
    .Q(\enigma.r.cnts_debug1[4] ));
 sg13g2_dfrbp_1 _2736_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net23),
    .D(_0044_),
    .Q_N(_1307_),
    .Q(\enigma.r.$signal$17[0] ));
 sg13g2_dfrbp_1 _2737_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net21),
    .D(_0045_),
    .Q_N(_1306_),
    .Q(\enigma.r.$signal$17[1] ));
 sg13g2_dfrbp_1 _2738_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net19),
    .D(_0046_),
    .Q_N(_0002_),
    .Q(\enigma.r.$signal$17[2] ));
 sg13g2_dfrbp_1 _2739_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net17),
    .D(_0047_),
    .Q_N(_1305_),
    .Q(\enigma.r.$signal$13[0] ));
 sg13g2_dfrbp_1 _2740_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net15),
    .D(_0048_),
    .Q_N(_1304_),
    .Q(\enigma.r.$signal$13[1] ));
 sg13g2_dfrbp_1 _2741_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net13),
    .D(_0049_),
    .Q_N(_1303_),
    .Q(\enigma.r.$signal$13[2] ));
 sg13g2_dfrbp_1 _2742_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net72),
    .D(_0050_),
    .Q_N(_1302_),
    .Q(\enigma.r.$signal$13[3] ));
 sg13g2_dfrbp_1 _2743_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net68),
    .D(_0051_),
    .Q_N(_1301_),
    .Q(\enigma.r.$signal$13[4] ));
 sg13g2_dfrbp_1 _2744_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net64),
    .D(_0052_),
    .Q_N(_1300_),
    .Q(\enigma.r.cnts_debug0[0] ));
 sg13g2_dfrbp_1 _2745_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net60),
    .D(_0053_),
    .Q_N(_1299_),
    .Q(\enigma.r.cnts_debug0[1] ));
 sg13g2_dfrbp_1 _2746_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net56),
    .D(_0054_),
    .Q_N(_1298_),
    .Q(\enigma.r.cnts_debug0[2] ));
 sg13g2_dfrbp_1 _2747_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net52),
    .D(_0055_),
    .Q_N(_1297_),
    .Q(\enigma.r.cnts_debug0[3] ));
 sg13g2_dfrbp_1 _2748_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net48),
    .D(_0056_),
    .Q_N(_1296_),
    .Q(\enigma.r.cnts_debug0[4] ));
 sg13g2_dlhq_1 _2749_ (.D(net605),
    .GATE(\enigma.plugboard.bits_0_0.clk ),
    .Q(\enigma.plugboard.bits_0_0.q ));
 sg13g2_dlhq_1 _2750_ (.D(net600),
    .GATE(\enigma.plugboard.bits_0_0.clk ),
    .Q(\enigma.plugboard.bits_0_1.q ));
 sg13g2_dlhq_1 _2751_ (.D(net596),
    .GATE(\enigma.plugboard.bits_0_0.clk ),
    .Q(\enigma.plugboard.bits_0_2.q ));
 sg13g2_dlhq_1 _2752_ (.D(net590),
    .GATE(\enigma.plugboard.bits_0_0.clk ),
    .Q(\enigma.plugboard.bits_0_3.q ));
 sg13g2_dlhq_1 _2753_ (.D(net587),
    .GATE(\enigma.plugboard.bits_0_0.clk ),
    .Q(\enigma.plugboard.bits_0_4.q ));
 sg13g2_dlhq_1 _2754_ (.D(net604),
    .GATE(\enigma.plugboard.bits_10_0.clk ),
    .Q(\enigma.plugboard.bits_10_0.q ));
 sg13g2_dlhq_1 _2755_ (.D(net599),
    .GATE(\enigma.plugboard.bits_10_0.clk ),
    .Q(\enigma.plugboard.bits_10_1.q ));
 sg13g2_dlhq_1 _2756_ (.D(net1),
    .GATE(\enigma.plugboard.bits_10_0.clk ),
    .Q(\enigma.plugboard.bits_10_2.q ));
 sg13g2_dlhq_1 _2757_ (.D(net590),
    .GATE(\enigma.plugboard.bits_10_0.clk ),
    .Q(\enigma.plugboard.bits_10_3.q ));
 sg13g2_dlhq_1 _2758_ (.D(net587),
    .GATE(\enigma.plugboard.bits_10_0.clk ),
    .Q(\enigma.plugboard.bits_10_4.q ));
 sg13g2_dlhq_1 _2759_ (.D(net604),
    .GATE(\enigma.plugboard.bits_11_0.clk ),
    .Q(\enigma.plugboard.bits_11_0.q ));
 sg13g2_dlhq_1 _2760_ (.D(net600),
    .GATE(\enigma.plugboard.bits_11_0.clk ),
    .Q(\enigma.plugboard.bits_11_1.q ));
 sg13g2_dlhq_1 _2761_ (.D(net596),
    .GATE(\enigma.plugboard.bits_11_0.clk ),
    .Q(\enigma.plugboard.bits_11_2.q ));
 sg13g2_dlhq_1 _2762_ (.D(net591),
    .GATE(\enigma.plugboard.bits_11_0.clk ),
    .Q(\enigma.plugboard.bits_11_3.q ));
 sg13g2_dlhq_1 _2763_ (.D(net588),
    .GATE(\enigma.plugboard.bits_11_0.clk ),
    .Q(\enigma.plugboard.bits_11_4.q ));
 sg13g2_dlhq_1 _2764_ (.D(net605),
    .GATE(\enigma.plugboard.bits_12_0.clk ),
    .Q(\enigma.plugboard.bits_12_0.q ));
 sg13g2_dlhq_1 _2765_ (.D(net599),
    .GATE(\enigma.plugboard.bits_12_0.clk ),
    .Q(\enigma.plugboard.bits_12_1.q ));
 sg13g2_dlhq_1 _2766_ (.D(net596),
    .GATE(\enigma.plugboard.bits_12_0.clk ),
    .Q(\enigma.plugboard.bits_12_2.q ));
 sg13g2_dlhq_1 _2767_ (.D(net592),
    .GATE(\enigma.plugboard.bits_12_0.clk ),
    .Q(\enigma.plugboard.bits_12_3.q ));
 sg13g2_dlhq_1 _2768_ (.D(net588),
    .GATE(\enigma.plugboard.bits_12_0.clk ),
    .Q(\enigma.plugboard.bits_12_4.q ));
 sg13g2_dlhq_1 _2769_ (.D(net604),
    .GATE(\enigma.plugboard.bits_13_0.clk ),
    .Q(\enigma.plugboard.bits_13_0.q ));
 sg13g2_dlhq_1 _2770_ (.D(net600),
    .GATE(\enigma.plugboard.bits_13_0.clk ),
    .Q(\enigma.plugboard.bits_13_1.q ));
 sg13g2_dlhq_1 _2771_ (.D(net595),
    .GATE(\enigma.plugboard.bits_13_0.clk ),
    .Q(\enigma.plugboard.bits_13_2.q ));
 sg13g2_dlhq_1 _2772_ (.D(net590),
    .GATE(\enigma.plugboard.bits_13_0.clk ),
    .Q(\enigma.plugboard.bits_13_3.q ));
 sg13g2_dlhq_1 _2773_ (.D(net586),
    .GATE(\enigma.plugboard.bits_13_0.clk ),
    .Q(\enigma.plugboard.bits_13_4.q ));
 sg13g2_dlhq_1 _2774_ (.D(net608),
    .GATE(\enigma.plugboard.bits_14_0.clk ),
    .Q(\enigma.plugboard.bits_14_0.q ));
 sg13g2_dlhq_1 _2775_ (.D(net599),
    .GATE(\enigma.plugboard.bits_14_0.clk ),
    .Q(\enigma.plugboard.bits_14_1.q ));
 sg13g2_dlhq_1 _2776_ (.D(net595),
    .GATE(\enigma.plugboard.bits_14_0.clk ),
    .Q(\enigma.plugboard.bits_14_2.q ));
 sg13g2_dlhq_1 _2777_ (.D(net591),
    .GATE(\enigma.plugboard.bits_14_0.clk ),
    .Q(\enigma.plugboard.bits_14_3.q ));
 sg13g2_dlhq_1 _2778_ (.D(net586),
    .GATE(\enigma.plugboard.bits_14_0.clk ),
    .Q(\enigma.plugboard.bits_14_4.q ));
 sg13g2_dlhq_1 _2779_ (.D(net605),
    .GATE(\enigma.plugboard.bits_15_0.clk ),
    .Q(\enigma.plugboard.bits_15_0.q ));
 sg13g2_dlhq_1 _2780_ (.D(net601),
    .GATE(\enigma.plugboard.bits_15_0.clk ),
    .Q(\enigma.plugboard.bits_15_1.q ));
 sg13g2_dlhq_1 _2781_ (.D(net595),
    .GATE(\enigma.plugboard.bits_15_0.clk ),
    .Q(\enigma.plugboard.bits_15_2.q ));
 sg13g2_dlhq_1 _2782_ (.D(net590),
    .GATE(\enigma.plugboard.bits_15_0.clk ),
    .Q(\enigma.plugboard.bits_15_3.q ));
 sg13g2_dlhq_1 _2783_ (.D(net586),
    .GATE(\enigma.plugboard.bits_15_0.clk ),
    .Q(\enigma.plugboard.bits_15_4.q ));
 sg13g2_dlhq_1 _2784_ (.D(net604),
    .GATE(\enigma.plugboard.bits_16_0.clk ),
    .Q(\enigma.plugboard.bits_16_0.q ));
 sg13g2_dlhq_1 _2785_ (.D(net599),
    .GATE(\enigma.plugboard.bits_16_0.clk ),
    .Q(\enigma.plugboard.bits_16_1.q ));
 sg13g2_dlhq_1 _2786_ (.D(net596),
    .GATE(\enigma.plugboard.bits_16_0.clk ),
    .Q(\enigma.plugboard.bits_16_2.q ));
 sg13g2_dlhq_1 _2787_ (.D(net593),
    .GATE(\enigma.plugboard.bits_16_0.clk ),
    .Q(\enigma.plugboard.bits_16_3.q ));
 sg13g2_dlhq_1 _2788_ (.D(net586),
    .GATE(\enigma.plugboard.bits_16_0.clk ),
    .Q(\enigma.plugboard.bits_16_4.q ));
 sg13g2_dlhq_1 _2789_ (.D(net605),
    .GATE(\enigma.plugboard.bits_17_0.clk ),
    .Q(\enigma.plugboard.bits_17_0.q ));
 sg13g2_dlhq_1 _2790_ (.D(net602),
    .GATE(\enigma.plugboard.bits_17_0.clk ),
    .Q(\enigma.plugboard.bits_17_1.q ));
 sg13g2_dlhq_1 _2791_ (.D(net595),
    .GATE(\enigma.plugboard.bits_17_0.clk ),
    .Q(\enigma.plugboard.bits_17_2.q ));
 sg13g2_dlhq_1 _2792_ (.D(net592),
    .GATE(\enigma.plugboard.bits_17_0.clk ),
    .Q(\enigma.plugboard.bits_17_3.q ));
 sg13g2_dlhq_1 _2793_ (.D(net586),
    .GATE(\enigma.plugboard.bits_17_0.clk ),
    .Q(\enigma.plugboard.bits_17_4.q ));
 sg13g2_dlhq_1 _2794_ (.D(net607),
    .GATE(\enigma.plugboard.bits_18_0.clk ),
    .Q(\enigma.plugboard.bits_18_0.q ));
 sg13g2_dlhq_1 _2795_ (.D(net602),
    .GATE(\enigma.plugboard.bits_18_0.clk ),
    .Q(\enigma.plugboard.bits_18_1.q ));
 sg13g2_dlhq_1 _2796_ (.D(net598),
    .GATE(\enigma.plugboard.bits_18_0.clk ),
    .Q(\enigma.plugboard.bits_18_2.q ));
 sg13g2_dlhq_1 _2797_ (.D(net593),
    .GATE(\enigma.plugboard.bits_18_0.clk ),
    .Q(\enigma.plugboard.bits_18_3.q ));
 sg13g2_dlhq_1 _2798_ (.D(net589),
    .GATE(\enigma.plugboard.bits_18_0.clk ),
    .Q(\enigma.plugboard.bits_18_4.q ));
 sg13g2_dlhq_1 _2799_ (.D(net607),
    .GATE(\enigma.plugboard.bits_19_0.clk ),
    .Q(\enigma.plugboard.bits_19_0.q ));
 sg13g2_dlhq_1 _2800_ (.D(net601),
    .GATE(\enigma.plugboard.bits_19_0.clk ),
    .Q(\enigma.plugboard.bits_19_1.q ));
 sg13g2_dlhq_1 _2801_ (.D(net597),
    .GATE(\enigma.plugboard.bits_19_0.clk ),
    .Q(\enigma.plugboard.bits_19_2.q ));
 sg13g2_dlhq_1 _2802_ (.D(net593),
    .GATE(\enigma.plugboard.bits_19_0.clk ),
    .Q(\enigma.plugboard.bits_19_3.q ));
 sg13g2_dlhq_1 _2803_ (.D(net589),
    .GATE(\enigma.plugboard.bits_19_0.clk ),
    .Q(\enigma.plugboard.bits_19_4.q ));
 sg13g2_dlhq_1 _2804_ (.D(net605),
    .GATE(\enigma.plugboard.bits_1_0.clk ),
    .Q(\enigma.plugboard.bits_1_0.q ));
 sg13g2_dlhq_1 _2805_ (.D(net600),
    .GATE(\enigma.plugboard.bits_1_0.clk ),
    .Q(\enigma.plugboard.bits_1_1.q ));
 sg13g2_dlhq_1 _2806_ (.D(net596),
    .GATE(\enigma.plugboard.bits_1_0.clk ),
    .Q(\enigma.plugboard.bits_1_2.q ));
 sg13g2_dlhq_1 _2807_ (.D(net591),
    .GATE(\enigma.plugboard.bits_1_0.clk ),
    .Q(\enigma.plugboard.bits_1_3.q ));
 sg13g2_dlhq_1 _2808_ (.D(net587),
    .GATE(\enigma.plugboard.bits_1_0.clk ),
    .Q(\enigma.plugboard.bits_1_4.q ));
 sg13g2_dlhq_1 _2809_ (.D(net605),
    .GATE(\enigma.plugboard.bits_20_0.clk ),
    .Q(\enigma.plugboard.bits_20_0.q ));
 sg13g2_dlhq_1 _2810_ (.D(net599),
    .GATE(\enigma.plugboard.bits_20_0.clk ),
    .Q(\enigma.plugboard.bits_20_1.q ));
 sg13g2_dlhq_1 _2811_ (.D(net596),
    .GATE(\enigma.plugboard.bits_20_0.clk ),
    .Q(\enigma.plugboard.bits_20_2.q ));
 sg13g2_dlhq_1 _2812_ (.D(net591),
    .GATE(\enigma.plugboard.bits_20_0.clk ),
    .Q(\enigma.plugboard.bits_20_3.q ));
 sg13g2_dlhq_1 _2813_ (.D(net587),
    .GATE(\enigma.plugboard.bits_20_0.clk ),
    .Q(\enigma.plugboard.bits_20_4.q ));
 sg13g2_dlhq_1 _2814_ (.D(net606),
    .GATE(\enigma.plugboard.bits_21_0.clk ),
    .Q(\enigma.plugboard.bits_21_0.q ));
 sg13g2_dlhq_1 _2815_ (.D(net602),
    .GATE(\enigma.plugboard.bits_21_0.clk ),
    .Q(\enigma.plugboard.bits_21_1.q ));
 sg13g2_dlhq_1 _2816_ (.D(net598),
    .GATE(\enigma.plugboard.bits_21_0.clk ),
    .Q(\enigma.plugboard.bits_21_2.q ));
 sg13g2_dlhq_1 _2817_ (.D(net592),
    .GATE(\enigma.plugboard.bits_21_0.clk ),
    .Q(\enigma.plugboard.bits_21_3.q ));
 sg13g2_dlhq_1 _2818_ (.D(net588),
    .GATE(\enigma.plugboard.bits_21_0.clk ),
    .Q(\enigma.plugboard.bits_21_4.q ));
 sg13g2_dlhq_1 _2819_ (.D(net607),
    .GATE(\enigma.plugboard.bits_22_0.clk ),
    .Q(\enigma.plugboard.bits_22_0.q ));
 sg13g2_dlhq_1 _2820_ (.D(net601),
    .GATE(\enigma.plugboard.bits_22_0.clk ),
    .Q(\enigma.plugboard.bits_22_1.q ));
 sg13g2_dlhq_1 _2821_ (.D(net598),
    .GATE(\enigma.plugboard.bits_22_0.clk ),
    .Q(\enigma.plugboard.bits_22_2.q ));
 sg13g2_dlhq_1 _2822_ (.D(net592),
    .GATE(\enigma.plugboard.bits_22_0.clk ),
    .Q(\enigma.plugboard.bits_22_3.q ));
 sg13g2_dlhq_1 _2823_ (.D(net588),
    .GATE(\enigma.plugboard.bits_22_0.clk ),
    .Q(\enigma.plugboard.bits_22_4.q ));
 sg13g2_dlhq_1 _2824_ (.D(net607),
    .GATE(\enigma.plugboard.bits_23_0.clk ),
    .Q(\enigma.plugboard.bits_23_0.q ));
 sg13g2_dlhq_1 _2825_ (.D(net602),
    .GATE(\enigma.plugboard.bits_23_0.clk ),
    .Q(\enigma.plugboard.bits_23_1.q ));
 sg13g2_dlhq_1 _2826_ (.D(net597),
    .GATE(\enigma.plugboard.bits_23_0.clk ),
    .Q(\enigma.plugboard.bits_23_2.q ));
 sg13g2_dlhq_1 _2827_ (.D(net593),
    .GATE(\enigma.plugboard.bits_23_0.clk ),
    .Q(\enigma.plugboard.bits_23_3.q ));
 sg13g2_dlhq_1 _2828_ (.D(net588),
    .GATE(\enigma.plugboard.bits_23_0.clk ),
    .Q(\enigma.plugboard.bits_23_4.q ));
 sg13g2_dlhq_1 _2829_ (.D(net606),
    .GATE(\enigma.plugboard.bits_24_0.clk ),
    .Q(\enigma.plugboard.bits_24_0.q ));
 sg13g2_dlhq_1 _2830_ (.D(net603),
    .GATE(\enigma.plugboard.bits_24_0.clk ),
    .Q(\enigma.plugboard.bits_24_1.q ));
 sg13g2_dlhq_1 _2831_ (.D(net597),
    .GATE(\enigma.plugboard.bits_24_0.clk ),
    .Q(\enigma.plugboard.bits_24_2.q ));
 sg13g2_dlhq_1 _2832_ (.D(net594),
    .GATE(\enigma.plugboard.bits_24_0.clk ),
    .Q(\enigma.plugboard.bits_24_3.q ));
 sg13g2_dlhq_1 _2833_ (.D(net589),
    .GATE(\enigma.plugboard.bits_24_0.clk ),
    .Q(\enigma.plugboard.bits_24_4.q ));
 sg13g2_dlhq_1 _2834_ (.D(net606),
    .GATE(\enigma.plugboard.bits_25_0.clk ),
    .Q(\enigma.plugboard.bits_25_0.q ));
 sg13g2_dlhq_1 _2835_ (.D(net601),
    .GATE(\enigma.plugboard.bits_25_0.clk ),
    .Q(\enigma.plugboard.bits_25_1.q ));
 sg13g2_dlhq_1 _2836_ (.D(net597),
    .GATE(\enigma.plugboard.bits_25_0.clk ),
    .Q(\enigma.plugboard.bits_25_2.q ));
 sg13g2_dlhq_1 _2837_ (.D(net592),
    .GATE(\enigma.plugboard.bits_25_0.clk ),
    .Q(\enigma.plugboard.bits_25_3.q ));
 sg13g2_dlhq_1 _2838_ (.D(net587),
    .GATE(\enigma.plugboard.bits_25_0.clk ),
    .Q(\enigma.plugboard.bits_25_4.q ));
 sg13g2_dlhq_1 _2839_ (.D(net606),
    .GATE(\enigma.plugboard.bits_2_0.clk ),
    .Q(\enigma.plugboard.bits_2_0.q ));
 sg13g2_dlhq_1 _2840_ (.D(net601),
    .GATE(\enigma.plugboard.bits_2_0.clk ),
    .Q(\enigma.plugboard.bits_2_1.q ));
 sg13g2_dlhq_1 _2841_ (.D(net598),
    .GATE(\enigma.plugboard.bits_2_0.clk ),
    .Q(\enigma.plugboard.bits_2_2.q ));
 sg13g2_dlhq_1 _2842_ (.D(net592),
    .GATE(\enigma.plugboard.bits_2_0.clk ),
    .Q(\enigma.plugboard.bits_2_3.q ));
 sg13g2_dlhq_1 _2843_ (.D(net588),
    .GATE(\enigma.plugboard.bits_2_0.clk ),
    .Q(\enigma.plugboard.bits_2_4.q ));
 sg13g2_dlhq_1 _2844_ (.D(net604),
    .GATE(\enigma.plugboard.bits_3_0.clk ),
    .Q(\enigma.plugboard.bits_3_0.q ));
 sg13g2_dlhq_1 _2845_ (.D(net599),
    .GATE(\enigma.plugboard.bits_3_0.clk ),
    .Q(\enigma.plugboard.bits_3_1.q ));
 sg13g2_dlhq_1 _2846_ (.D(net596),
    .GATE(\enigma.plugboard.bits_3_0.clk ),
    .Q(\enigma.plugboard.bits_3_2.q ));
 sg13g2_dlhq_1 _2847_ (.D(net591),
    .GATE(\enigma.plugboard.bits_3_0.clk ),
    .Q(\enigma.plugboard.bits_3_3.q ));
 sg13g2_dlhq_1 _2848_ (.D(net587),
    .GATE(\enigma.plugboard.bits_3_0.clk ),
    .Q(\enigma.plugboard.bits_3_4.q ));
 sg13g2_dlhq_1 _2849_ (.D(net607),
    .GATE(\enigma.plugboard.bits_4_0.clk ),
    .Q(\enigma.plugboard.bits_4_0.q ));
 sg13g2_dlhq_1 _2850_ (.D(net602),
    .GATE(\enigma.plugboard.bits_4_0.clk ),
    .Q(\enigma.plugboard.bits_4_1.q ));
 sg13g2_dlhq_1 _2851_ (.D(net598),
    .GATE(\enigma.plugboard.bits_4_0.clk ),
    .Q(\enigma.plugboard.bits_4_2.q ));
 sg13g2_dlhq_1 _2852_ (.D(net592),
    .GATE(\enigma.plugboard.bits_4_0.clk ),
    .Q(\enigma.plugboard.bits_4_3.q ));
 sg13g2_dlhq_1 _2853_ (.D(net588),
    .GATE(\enigma.plugboard.bits_4_0.clk ),
    .Q(\enigma.plugboard.bits_4_4.q ));
 sg13g2_dlhq_1 _2854_ (.D(net604),
    .GATE(\enigma.plugboard.bits_5_0.clk ),
    .Q(\enigma.plugboard.bits_5_0.q ));
 sg13g2_dlhq_1 _2855_ (.D(net599),
    .GATE(\enigma.plugboard.bits_5_0.clk ),
    .Q(\enigma.plugboard.bits_5_1.q ));
 sg13g2_dlhq_1 _2856_ (.D(net595),
    .GATE(\enigma.plugboard.bits_5_0.clk ),
    .Q(\enigma.plugboard.bits_5_2.q ));
 sg13g2_dlhq_1 _2857_ (.D(net590),
    .GATE(\enigma.plugboard.bits_5_0.clk ),
    .Q(\enigma.plugboard.bits_5_3.q ));
 sg13g2_dlhq_1 _2858_ (.D(net587),
    .GATE(\enigma.plugboard.bits_5_0.clk ),
    .Q(\enigma.plugboard.bits_5_4.q ));
 sg13g2_dlhq_1 _2859_ (.D(net604),
    .GATE(\enigma.plugboard.bits_6_0.clk ),
    .Q(\enigma.plugboard.bits_6_0.q ));
 sg13g2_dlhq_1 _2860_ (.D(net600),
    .GATE(\enigma.plugboard.bits_6_0.clk ),
    .Q(\enigma.plugboard.bits_6_1.q ));
 sg13g2_dlhq_1 _2861_ (.D(net595),
    .GATE(\enigma.plugboard.bits_6_0.clk ),
    .Q(\enigma.plugboard.bits_6_2.q ));
 sg13g2_dlhq_1 _2862_ (.D(net590),
    .GATE(\enigma.plugboard.bits_6_0.clk ),
    .Q(\enigma.plugboard.bits_6_3.q ));
 sg13g2_dlhq_1 _2863_ (.D(net586),
    .GATE(\enigma.plugboard.bits_6_0.clk ),
    .Q(\enigma.plugboard.bits_6_4.q ));
 sg13g2_dlhq_1 _2864_ (.D(net604),
    .GATE(\enigma.plugboard.bits_7_0.clk ),
    .Q(\enigma.plugboard.bits_7_0.q ));
 sg13g2_dlhq_1 _2865_ (.D(net599),
    .GATE(\enigma.plugboard.bits_7_0.clk ),
    .Q(\enigma.plugboard.bits_7_1.q ));
 sg13g2_dlhq_1 _2866_ (.D(net595),
    .GATE(\enigma.plugboard.bits_7_0.clk ),
    .Q(\enigma.plugboard.bits_7_2.q ));
 sg13g2_dlhq_1 _2867_ (.D(net590),
    .GATE(\enigma.plugboard.bits_7_0.clk ),
    .Q(\enigma.plugboard.bits_7_3.q ));
 sg13g2_dlhq_1 _2868_ (.D(net586),
    .GATE(\enigma.plugboard.bits_7_0.clk ),
    .Q(\enigma.plugboard.bits_7_4.q ));
 sg13g2_dlhq_1 _2869_ (.D(net607),
    .GATE(\enigma.plugboard.bits_8_0.clk ),
    .Q(\enigma.plugboard.bits_8_0.q ));
 sg13g2_dlhq_1 _2870_ (.D(net602),
    .GATE(\enigma.plugboard.bits_8_0.clk ),
    .Q(\enigma.plugboard.bits_8_1.q ));
 sg13g2_dlhq_1 _2871_ (.D(net597),
    .GATE(\enigma.plugboard.bits_8_0.clk ),
    .Q(\enigma.plugboard.bits_8_2.q ));
 sg13g2_dlhq_1 _2872_ (.D(net593),
    .GATE(\enigma.plugboard.bits_8_0.clk ),
    .Q(\enigma.plugboard.bits_8_3.q ));
 sg13g2_dlhq_1 _2873_ (.D(net589),
    .GATE(\enigma.plugboard.bits_8_0.clk ),
    .Q(\enigma.plugboard.bits_8_4.q ));
 sg13g2_dlhq_1 _2874_ (.D(net605),
    .GATE(\enigma.plugboard.bits_9_0.clk ),
    .Q(\enigma.plugboard.bits_9_0.q ));
 sg13g2_dlhq_1 _2875_ (.D(net600),
    .GATE(\enigma.plugboard.bits_9_0.clk ),
    .Q(\enigma.plugboard.bits_9_1.q ));
 sg13g2_dlhq_1 _2876_ (.D(net595),
    .GATE(\enigma.plugboard.bits_9_0.clk ),
    .Q(\enigma.plugboard.bits_9_2.q ));
 sg13g2_dlhq_1 _2877_ (.D(net590),
    .GATE(\enigma.plugboard.bits_9_0.clk ),
    .Q(\enigma.plugboard.bits_9_3.q ));
 sg13g2_dlhq_1 _2878_ (.D(net586),
    .GATE(\enigma.plugboard.bits_9_0.clk ),
    .Q(\enigma.plugboard.bits_9_4.q ));
 sg13g2_dfrbp_1 _2879_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net44),
    .D(net84),
    .Q_N(\enigma.plugboard.$31[0] ),
    .Q(\enigma.plugboard.plug_limiter[0] ));
 sg13g2_dfrbp_1 _2880_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net40),
    .D(net92),
    .Q_N(_1295_),
    .Q(\enigma.plugboard.plug_limiter[1] ));
 sg13g2_dfrbp_1 _2881_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net36),
    .D(_0059_),
    .Q_N(_1294_),
    .Q(\enigma.plugboard.plug_limiter[2] ));
 sg13g2_dfrbp_1 _2882_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net32),
    .D(_0060_),
    .Q_N(_1293_),
    .Q(\enigma.plugboard.plug_limiter[3] ));
 sg13g2_dfrbp_1 _2883_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net28),
    .D(_0061_),
    .Q_N(_1292_),
    .Q(\enigma.plugboard.plug_limiter[4] ));
 sg13g2_dfrbp_1 _2884_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net24),
    .D(_0062_),
    .Q_N(_1291_),
    .Q(\enigma.plugboard.cnt[0] ));
 sg13g2_dfrbp_1 _2885_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net20),
    .D(_0063_),
    .Q_N(_1290_),
    .Q(\enigma.plugboard.cnt[1] ));
 sg13g2_dfrbp_1 _2886_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net16),
    .D(_0064_),
    .Q_N(_1289_),
    .Q(\enigma.plugboard.cnt[2] ));
 sg13g2_dfrbp_1 _2887_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net74),
    .D(net131),
    .Q_N(_1288_),
    .Q(\enigma.plugboard.cnt[3] ));
 sg13g2_dfrbp_1 _2888_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net66),
    .D(net109),
    .Q_N(_0007_),
    .Q(\enigma.plugboard.cnt[4] ));
 sg13g2_dfrbp_1 _2889_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net58),
    .D(_0067_),
    .Q_N(_1287_),
    .Q(\enigma.fsm.fsm_state[0] ));
 sg13g2_dfrbp_1 _2890_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net50),
    .D(net145),
    .Q_N(_1286_),
    .Q(\enigma.fsm.fsm_state[1] ));
 sg13g2_dfrbp_1 _2891_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net42),
    .D(net90),
    .Q_N(_0009_),
    .Q(\enigma.fsm.fsm_state[2] ));
 sg13g2_dfrbp_1 _2892_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net34),
    .D(_0070_),
    .Q_N(_0010_),
    .Q(\enigma.fsm.fsm_state[3] ));
 sg13g2_dfrbp_1 _2893_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net26),
    .D(_0071_),
    .Q_N(_0008_),
    .Q(\enigma.fsm.fsm_state[4] ));
 sg13g2_dfrbp_1 _2894_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net18),
    .D(_0072_),
    .Q_N(_0006_),
    .Q(\enigma.fsm.double_step ));
 sg13g2_dfrbp_1 _2895_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net70),
    .D(_0073_),
    .Q_N(_1285_),
    .Q(\enigma.fsm.cnt[0] ));
 sg13g2_dfrbp_1 _2896_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net54),
    .D(_0074_),
    .Q_N(_1284_),
    .Q(\enigma.fsm.cnt[1] ));
 sg13g2_dfrbp_1 _2897_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net38),
    .D(_0075_),
    .Q_N(_0005_),
    .Q(net563));
 sg13g2_dfrbp_1 _2898_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net22),
    .D(_0076_),
    .Q_N(_1283_),
    .Q(net562));
 sg13g2_dfrbp_1 _2899_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net62),
    .D(_0077_),
    .Q_N(_0004_),
    .Q(net561));
 sg13g2_dfrbp_1 _2900_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net30),
    .D(_0078_),
    .Q_N(_1282_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _2901_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net46),
    .D(_0079_),
    .Q_N(_0003_),
    .Q(net557));
 sg13g2_tiehi _2709__9 (.L_HI(net9));
 sg13g2_tiehi _2708__10 (.L_HI(net10));
 sg13g2_tiehi _2707__11 (.L_HI(net11));
 sg13g2_tiehi _2706__12 (.L_HI(net12));
 sg13g2_tiehi _2741__13 (.L_HI(net13));
 sg13g2_tiehi _2705__14 (.L_HI(net14));
 sg13g2_tiehi _2740__15 (.L_HI(net15));
 sg13g2_tiehi _2886__16 (.L_HI(net16));
 sg13g2_tiehi _2739__17 (.L_HI(net17));
 sg13g2_tiehi _2894__18 (.L_HI(net18));
 sg13g2_tiehi _2738__19 (.L_HI(net19));
 sg13g2_tiehi _2885__20 (.L_HI(net20));
 sg13g2_tiehi _2737__21 (.L_HI(net21));
 sg13g2_tiehi _2898__22 (.L_HI(net22));
 sg13g2_tiehi _2736__23 (.L_HI(net23));
 sg13g2_tiehi _2884__24 (.L_HI(net24));
 sg13g2_tiehi _2735__25 (.L_HI(net25));
 sg13g2_tiehi _2893__26 (.L_HI(net26));
 sg13g2_tiehi _2734__27 (.L_HI(net27));
 sg13g2_tiehi _2883__28 (.L_HI(net28));
 sg13g2_tiehi _2733__29 (.L_HI(net29));
 sg13g2_tiehi _2900__30 (.L_HI(net30));
 sg13g2_tiehi _2732__31 (.L_HI(net31));
 sg13g2_tiehi _2882__32 (.L_HI(net32));
 sg13g2_tiehi _2731__33 (.L_HI(net33));
 sg13g2_tiehi _2892__34 (.L_HI(net34));
 sg13g2_tiehi _2730__35 (.L_HI(net35));
 sg13g2_tiehi _2881__36 (.L_HI(net36));
 sg13g2_tiehi _2729__37 (.L_HI(net37));
 sg13g2_tiehi _2897__38 (.L_HI(net38));
 sg13g2_tiehi _2728__39 (.L_HI(net39));
 sg13g2_tiehi _2880__40 (.L_HI(net40));
 sg13g2_tiehi _2727__41 (.L_HI(net41));
 sg13g2_tiehi _2891__42 (.L_HI(net42));
 sg13g2_tiehi _2726__43 (.L_HI(net43));
 sg13g2_tiehi _2879__44 (.L_HI(net44));
 sg13g2_tiehi _2725__45 (.L_HI(net45));
 sg13g2_tiehi _2901__46 (.L_HI(net46));
 sg13g2_tiehi _2724__47 (.L_HI(net47));
 sg13g2_tiehi _2748__48 (.L_HI(net48));
 sg13g2_tiehi _2723__49 (.L_HI(net49));
 sg13g2_tiehi _2890__50 (.L_HI(net50));
 sg13g2_tiehi _2722__51 (.L_HI(net51));
 sg13g2_tiehi _2747__52 (.L_HI(net52));
 sg13g2_tiehi _2721__53 (.L_HI(net53));
 sg13g2_tiehi _2896__54 (.L_HI(net54));
 sg13g2_tiehi _2720__55 (.L_HI(net55));
 sg13g2_tiehi _2746__56 (.L_HI(net56));
 sg13g2_tiehi _2719__57 (.L_HI(net57));
 sg13g2_tiehi _2889__58 (.L_HI(net58));
 sg13g2_tiehi _2718__59 (.L_HI(net59));
 sg13g2_tiehi _2745__60 (.L_HI(net60));
 sg13g2_tiehi _2717__61 (.L_HI(net61));
 sg13g2_tiehi _2899__62 (.L_HI(net62));
 sg13g2_tiehi _2716__63 (.L_HI(net63));
 sg13g2_tiehi _2744__64 (.L_HI(net64));
 sg13g2_tiehi _2715__65 (.L_HI(net65));
 sg13g2_tiehi _2888__66 (.L_HI(net66));
 sg13g2_tiehi _2714__67 (.L_HI(net67));
 sg13g2_tiehi _2743__68 (.L_HI(net68));
 sg13g2_tiehi _2713__69 (.L_HI(net69));
 sg13g2_tiehi _2895__70 (.L_HI(net70));
 sg13g2_tiehi _2712__71 (.L_HI(net71));
 sg13g2_tiehi _2742__72 (.L_HI(net72));
 sg13g2_tiehi _2711__73 (.L_HI(net73));
 sg13g2_tiehi _2887__74 (.L_HI(net74));
 sg13g2_tiehi tt_um_virantha_enigma_75 (.L_HI(net75));
 sg13g2_tiehi tt_um_virantha_enigma_76 (.L_HI(net76));
 sg13g2_tiehi tt_um_virantha_enigma_77 (.L_HI(net77));
 sg13g2_tiehi tt_um_virantha_enigma_78 (.L_HI(net78));
 sg13g2_tiehi tt_um_virantha_enigma_79 (.L_HI(net79));
 sg13g2_tiehi tt_um_virantha_enigma_80 (.L_HI(net80));
 sg13g2_tiehi tt_um_virantha_enigma_81 (.L_HI(net81));
 sg13g2_tiehi tt_um_virantha_enigma_82 (.L_HI(net82));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_virantha_enigma_6 (.L_LO(net6));
 sg13g2_tielo tt_um_virantha_enigma_7 (.L_LO(net7));
 sg13g2_tiehi _2710__8 (.L_HI(net8));
 sg13g2_buf_1 _2980_ (.A(\enigma.fsm.ready ),
    .X(uio_out[5]));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(_1145_));
 sg13g2_buf_2 fanout466 (.A(_1145_),
    .X(net466));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(_1155_));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(_1132_));
 sg13g2_buf_2 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_1130_),
    .X(net470));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(_1129_));
 sg13g2_buf_2 fanout472 (.A(_1129_),
    .X(net472));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(net478));
 sg13g2_buf_4 fanout474 (.X(net474),
    .A(net475));
 sg13g2_buf_4 fanout475 (.X(net475),
    .A(net478));
 sg13g2_buf_2 fanout476 (.A(net477),
    .X(net476));
 sg13g2_buf_1 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_1121_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(net482),
    .X(net479));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(net481));
 sg13g2_buf_4 fanout481 (.X(net481),
    .A(net482));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(_1120_));
 sg13g2_buf_4 fanout483 (.X(net483),
    .A(_1114_));
 sg13g2_buf_2 fanout484 (.A(net485),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_1105_),
    .X(net486));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(net489));
 sg13g2_buf_1 fanout488 (.A(net489),
    .X(net488));
 sg13g2_buf_4 fanout489 (.X(net489),
    .A(_1105_));
 sg13g2_buf_2 fanout490 (.A(_1104_),
    .X(net490));
 sg13g2_buf_1 fanout491 (.A(_1104_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(net493),
    .X(net492));
 sg13g2_buf_4 fanout493 (.X(net493),
    .A(net494));
 sg13g2_buf_4 fanout494 (.X(net494),
    .A(_1104_));
 sg13g2_buf_2 fanout495 (.A(net499),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(net498),
    .X(net496));
 sg13g2_buf_1 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(net499),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_1101_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_1100_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(net504),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_1100_),
    .X(net503));
 sg13g2_buf_1 fanout504 (.A(_1100_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(net506),
    .X(net505));
 sg13g2_buf_1 fanout506 (.A(net507),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_1107_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net510),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_1 fanout510 (.A(net511),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_1106_),
    .X(net511));
 sg13g2_buf_4 fanout512 (.X(net512),
    .A(_0951_));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(_0878_));
 sg13g2_buf_2 fanout514 (.A(_0996_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_0523_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_0517_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_0507_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_0501_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_0475_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_0465_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(net522),
    .X(net521));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(_0779_));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(_0777_));
 sg13g2_buf_1 fanout524 (.A(_0777_),
    .X(net524));
 sg13g2_buf_4 fanout525 (.X(net525),
    .A(_0775_));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(_0817_));
 sg13g2_buf_2 fanout527 (.A(_0817_),
    .X(net527));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(_0816_));
 sg13g2_buf_2 fanout529 (.A(_0816_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(net531),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_0815_),
    .X(net531));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(net533));
 sg13g2_buf_4 fanout533 (.X(net533),
    .A(_0814_));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(_0813_));
 sg13g2_buf_2 fanout535 (.A(_0813_),
    .X(net535));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(_0812_));
 sg13g2_buf_2 fanout537 (.A(_0812_),
    .X(net537));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(_0799_));
 sg13g2_buf_2 fanout539 (.A(_0772_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_0767_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_0765_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_0751_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(net544),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_0541_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_1238_),
    .X(net545));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(_1235_));
 sg13g2_buf_4 fanout547 (.X(net547),
    .A(_1231_));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(_1214_));
 sg13g2_buf_2 fanout549 (.A(_1211_),
    .X(net549));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(_1209_));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(_1163_));
 sg13g2_buf_2 fanout552 (.A(_1143_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_0792_),
    .X(net553));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(_1217_));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(_1189_));
 sg13g2_buf_2 fanout556 (.A(uio_out[4]),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(net557),
    .X(uio_out[4]));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(uio_out[3]),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(uio_out[2]),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net561),
    .X(uio_out[2]));
 sg13g2_buf_2 fanout562 (.A(net562),
    .X(uio_out[1]));
 sg13g2_buf_4 fanout563 (.X(uio_out[0]),
    .A(net142));
 sg13g2_buf_1 fanout564 (.A(net563),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_0008_),
    .X(net565));
 sg13g2_buf_1 fanout566 (.A(_0008_),
    .X(net566));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(net146));
 sg13g2_buf_2 fanout568 (.A(\enigma.fsm.fsm_state[4] ),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(\enigma.fsm.fsm_state[3] ),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(\enigma.fsm.fsm_state[3] ),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(\enigma.fsm.fsm_state[2] ),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(\enigma.fsm.fsm_state[2] ),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_1 fanout574 (.A(net144),
    .X(net574));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(\enigma.fsm.fsm_state[0] ));
 sg13g2_buf_2 fanout576 (.A(_0002_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net149),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net150),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net147),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(\enigma.r.dout[4] ),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(\enigma.r.dout[3] ),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(\enigma.r.dout[2] ),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(\enigma.r.dout[1] ),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_1 fanout585 (.A(\enigma.r.dout[0] ),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(ui_in[4]),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(ui_in[4]),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(ui_in[4]),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(net594),
    .X(net590));
 sg13g2_buf_1 fanout591 (.A(net594),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(ui_in[3]),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(net596),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(net1),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(net598),
    .X(net597));
 sg13g2_buf_4 fanout598 (.X(net598),
    .A(net1));
 sg13g2_buf_2 fanout599 (.A(net600),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(net601),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(net603),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(ui_in[1]),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(net608),
    .X(net605));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(net608));
 sg13g2_buf_2 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_1 fanout608 (.A(ui_in[0]),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(net610),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(net611),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(net618),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(net614),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_4 fanout615 (.X(net615),
    .A(net618));
 sg13g2_buf_2 fanout616 (.A(net618),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(rst_n),
    .X(net618));
 sg13g2_buf_2 input1 (.A(ui_in[2]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[5]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[6]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[7]),
    .X(net4));
 sg13g2_tielo tt_um_virantha_enigma_5 (.L_LO(net5));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\enigma.plugboard.$31[0] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0057_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold3 (.A(\enigma.plugboard.plug_limiter[3] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold4 (.A(\enigma.plugboard.plug_limiter[4] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold5 (.A(\enigma.plugboard.plug_limiter[2] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0540_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0006_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0069_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold9 (.A(\enigma.plugboard.plug_limiter[1] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0058_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold11 (.A(\enigma.fsm.cnt[0] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0621_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold13 (.A(\enigma.r.$signal$23[2] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold14 (.A(\enigma.r.$signal$22[4] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold15 (.A(\enigma.r.cnts_debug2[1] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold16 (.A(\enigma.r.cnts_debug2[2] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold17 (.A(\enigma.r.$signal$20[3] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold18 (.A(\enigma.r.cnts_debug2[3] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold19 (.A(\enigma.r.cnts_debug2[0] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold20 (.A(\enigma.r.$signal$20[1] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold21 (.A(\enigma.r.$signal$22[2] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold22 (.A(\enigma.r.$signal$20[2] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold23 (.A(\enigma.r.$signal$13[4] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold24 (.A(\enigma.r.$signal$22[1] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold25 (.A(\enigma.r.$signal$20[4] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold26 (.A(\enigma.plugboard.cnt[4] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0066_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold28 (.A(\enigma.r.cnts_debug1[4] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold29 (.A(\enigma.r.$signal$20[0] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold30 (.A(\enigma.r.$signal$13[2] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold31 (.A(\enigma.r.$signal$22[3] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold32 (.A(\enigma.r.$signal$13[0] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold33 (.A(\enigma.r.cnts_debug2[4] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold34 (.A(\enigma.r.$signal$13[3] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold35 (.A(\enigma.r.$signal$22[0] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold36 (.A(\enigma.r.$signal$13[1] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold37 (.A(net562),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold38 (.A(\enigma.r.cnts_debug1[3] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold39 (.A(\enigma.r.cnts_debug1[2] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold40 (.A(\enigma.r.cnts_debug0[4] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold41 (.A(\enigma.r.cnts_debug0[3] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold42 (.A(\enigma.r.cnts_debug1[1] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold43 (.A(\enigma.r.cnts_debug0[2] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold44 (.A(\enigma.r.cnts_debug0[1] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold45 (.A(\enigma.fsm.cnt[1] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold46 (.A(\enigma.r.$signal$21[2] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold47 (.A(\enigma.r.cnts_debug0[0] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold48 (.A(\enigma.plugboard.cnt[3] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0065_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold50 (.A(\enigma.r.$signal$17[2] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold51 (.A(\enigma.r.cnts_debug1[0] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold52 (.A(\enigma.fsm.fsm_state[0] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold53 (.A(\enigma.plugboard.cnt[1] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold54 (.A(\enigma.plugboard.cnt[2] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold55 (.A(\enigma.fsm.double_step ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold56 (.A(\enigma.r.$signal$23[1] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0019_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold58 (.A(\enigma.r.$signal$23[0] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold59 (.A(\enigma.plugboard.cnt[0] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold60 (.A(net563),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold61 (.A(\enigma.r.$signal$21[1] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold62 (.A(\enigma.fsm.fsm_state[1] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0068_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold64 (.A(\enigma.fsm.fsm_state[4] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold65 (.A(\enigma.r.$signal$21[0] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0031_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold67 (.A(\enigma.r.$signal$17[1] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold68 (.A(\enigma.r.$signal$17[0] ),
    .X(net150));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_fill_1 FILLER_0_49 ();
 sg13g2_decap_4 FILLER_0_59 ();
 sg13g2_fill_2 FILLER_0_63 ();
 sg13g2_decap_4 FILLER_0_87 ();
 sg13g2_fill_1 FILLER_0_91 ();
 sg13g2_fill_2 FILLER_0_96 ();
 sg13g2_decap_4 FILLER_0_126 ();
 sg13g2_fill_1 FILLER_0_135 ();
 sg13g2_decap_4 FILLER_0_147 ();
 sg13g2_fill_2 FILLER_0_151 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_fill_1 FILLER_0_175 ();
 sg13g2_fill_1 FILLER_0_193 ();
 sg13g2_fill_1 FILLER_0_202 ();
 sg13g2_fill_1 FILLER_0_208 ();
 sg13g2_fill_2 FILLER_0_234 ();
 sg13g2_fill_1 FILLER_0_236 ();
 sg13g2_fill_2 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_fill_2 FILLER_0_270 ();
 sg13g2_fill_1 FILLER_0_272 ();
 sg13g2_decap_8 FILLER_0_307 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_4 FILLER_0_321 ();
 sg13g2_fill_2 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_361 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_4 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_fill_1 FILLER_1_32 ();
 sg13g2_fill_1 FILLER_1_73 ();
 sg13g2_fill_1 FILLER_1_108 ();
 sg13g2_fill_2 FILLER_1_127 ();
 sg13g2_fill_2 FILLER_1_142 ();
 sg13g2_fill_1 FILLER_1_144 ();
 sg13g2_fill_2 FILLER_1_171 ();
 sg13g2_fill_1 FILLER_1_195 ();
 sg13g2_fill_2 FILLER_1_206 ();
 sg13g2_fill_2 FILLER_1_218 ();
 sg13g2_fill_1 FILLER_1_225 ();
 sg13g2_fill_1 FILLER_1_244 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_fill_2 FILLER_1_273 ();
 sg13g2_decap_4 FILLER_1_292 ();
 sg13g2_fill_1 FILLER_1_296 ();
 sg13g2_decap_4 FILLER_1_314 ();
 sg13g2_fill_1 FILLER_1_318 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_fill_2 FILLER_1_343 ();
 sg13g2_fill_1 FILLER_1_345 ();
 sg13g2_decap_4 FILLER_1_363 ();
 sg13g2_fill_2 FILLER_1_367 ();
 sg13g2_fill_2 FILLER_1_386 ();
 sg13g2_fill_1 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_21 ();
 sg13g2_fill_1 FILLER_2_23 ();
 sg13g2_decap_4 FILLER_2_40 ();
 sg13g2_fill_1 FILLER_2_82 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_fill_2 FILLER_2_95 ();
 sg13g2_fill_2 FILLER_2_115 ();
 sg13g2_fill_1 FILLER_2_117 ();
 sg13g2_decap_4 FILLER_2_148 ();
 sg13g2_fill_2 FILLER_2_152 ();
 sg13g2_fill_2 FILLER_2_161 ();
 sg13g2_fill_1 FILLER_2_163 ();
 sg13g2_decap_4 FILLER_2_176 ();
 sg13g2_decap_4 FILLER_2_185 ();
 sg13g2_fill_2 FILLER_2_189 ();
 sg13g2_decap_4 FILLER_2_212 ();
 sg13g2_decap_4 FILLER_2_236 ();
 sg13g2_fill_2 FILLER_2_240 ();
 sg13g2_fill_1 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_fill_1 FILLER_2_272 ();
 sg13g2_fill_1 FILLER_2_290 ();
 sg13g2_decap_8 FILLER_2_341 ();
 sg13g2_fill_1 FILLER_2_348 ();
 sg13g2_fill_1 FILLER_2_389 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_fill_2 FILLER_3_41 ();
 sg13g2_fill_1 FILLER_3_43 ();
 sg13g2_fill_2 FILLER_3_73 ();
 sg13g2_fill_1 FILLER_3_75 ();
 sg13g2_fill_2 FILLER_3_82 ();
 sg13g2_fill_1 FILLER_3_84 ();
 sg13g2_decap_4 FILLER_3_98 ();
 sg13g2_fill_1 FILLER_3_107 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_fill_2 FILLER_3_123 ();
 sg13g2_fill_1 FILLER_3_125 ();
 sg13g2_fill_2 FILLER_3_130 ();
 sg13g2_fill_2 FILLER_3_147 ();
 sg13g2_fill_2 FILLER_3_153 ();
 sg13g2_fill_1 FILLER_3_155 ();
 sg13g2_fill_2 FILLER_3_165 ();
 sg13g2_decap_4 FILLER_3_194 ();
 sg13g2_decap_4 FILLER_3_209 ();
 sg13g2_fill_2 FILLER_3_213 ();
 sg13g2_fill_1 FILLER_3_220 ();
 sg13g2_decap_4 FILLER_3_231 ();
 sg13g2_fill_1 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_257 ();
 sg13g2_decap_4 FILLER_3_264 ();
 sg13g2_fill_1 FILLER_3_268 ();
 sg13g2_decap_4 FILLER_3_314 ();
 sg13g2_fill_2 FILLER_3_340 ();
 sg13g2_fill_1 FILLER_3_342 ();
 sg13g2_decap_8 FILLER_3_372 ();
 sg13g2_decap_4 FILLER_3_379 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_4 FILLER_4_7 ();
 sg13g2_decap_4 FILLER_4_15 ();
 sg13g2_fill_2 FILLER_4_19 ();
 sg13g2_fill_1 FILLER_4_43 ();
 sg13g2_fill_2 FILLER_4_54 ();
 sg13g2_fill_1 FILLER_4_56 ();
 sg13g2_decap_4 FILLER_4_72 ();
 sg13g2_fill_2 FILLER_4_88 ();
 sg13g2_decap_4 FILLER_4_95 ();
 sg13g2_fill_2 FILLER_4_99 ();
 sg13g2_decap_8 FILLER_4_152 ();
 sg13g2_fill_2 FILLER_4_173 ();
 sg13g2_fill_1 FILLER_4_203 ();
 sg13g2_fill_2 FILLER_4_218 ();
 sg13g2_fill_1 FILLER_4_220 ();
 sg13g2_fill_2 FILLER_4_239 ();
 sg13g2_decap_8 FILLER_4_269 ();
 sg13g2_fill_1 FILLER_4_276 ();
 sg13g2_decap_4 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_327 ();
 sg13g2_fill_2 FILLER_4_336 ();
 sg13g2_fill_2 FILLER_4_344 ();
 sg13g2_fill_1 FILLER_4_346 ();
 sg13g2_fill_1 FILLER_4_370 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_fill_2 FILLER_5_26 ();
 sg13g2_fill_1 FILLER_5_28 ();
 sg13g2_fill_2 FILLER_5_55 ();
 sg13g2_fill_1 FILLER_5_57 ();
 sg13g2_fill_1 FILLER_5_68 ();
 sg13g2_fill_2 FILLER_5_100 ();
 sg13g2_fill_1 FILLER_5_102 ();
 sg13g2_fill_1 FILLER_5_110 ();
 sg13g2_fill_1 FILLER_5_121 ();
 sg13g2_decap_8 FILLER_5_127 ();
 sg13g2_fill_1 FILLER_5_134 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_fill_1 FILLER_5_153 ();
 sg13g2_fill_2 FILLER_5_171 ();
 sg13g2_fill_1 FILLER_5_173 ();
 sg13g2_decap_8 FILLER_5_190 ();
 sg13g2_fill_2 FILLER_5_197 ();
 sg13g2_decap_4 FILLER_5_209 ();
 sg13g2_fill_2 FILLER_5_213 ();
 sg13g2_decap_8 FILLER_5_268 ();
 sg13g2_decap_8 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_282 ();
 sg13g2_decap_8 FILLER_5_289 ();
 sg13g2_fill_2 FILLER_5_318 ();
 sg13g2_decap_4 FILLER_5_354 ();
 sg13g2_fill_1 FILLER_5_358 ();
 sg13g2_decap_4 FILLER_5_382 ();
 sg13g2_fill_2 FILLER_6_19 ();
 sg13g2_fill_2 FILLER_6_29 ();
 sg13g2_fill_2 FILLER_6_40 ();
 sg13g2_fill_1 FILLER_6_42 ();
 sg13g2_fill_2 FILLER_6_53 ();
 sg13g2_fill_1 FILLER_6_55 ();
 sg13g2_decap_4 FILLER_6_78 ();
 sg13g2_fill_1 FILLER_6_82 ();
 sg13g2_decap_4 FILLER_6_89 ();
 sg13g2_fill_1 FILLER_6_93 ();
 sg13g2_fill_2 FILLER_6_121 ();
 sg13g2_fill_2 FILLER_6_138 ();
 sg13g2_fill_2 FILLER_6_151 ();
 sg13g2_fill_1 FILLER_6_153 ();
 sg13g2_decap_4 FILLER_6_170 ();
 sg13g2_fill_2 FILLER_6_174 ();
 sg13g2_fill_1 FILLER_6_184 ();
 sg13g2_fill_1 FILLER_6_194 ();
 sg13g2_decap_4 FILLER_6_214 ();
 sg13g2_fill_2 FILLER_6_232 ();
 sg13g2_fill_1 FILLER_6_234 ();
 sg13g2_decap_4 FILLER_6_252 ();
 sg13g2_decap_4 FILLER_6_264 ();
 sg13g2_fill_2 FILLER_6_268 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_fill_2 FILLER_6_350 ();
 sg13g2_fill_1 FILLER_6_352 ();
 sg13g2_fill_1 FILLER_6_382 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_fill_2 FILLER_7_38 ();
 sg13g2_fill_2 FILLER_7_55 ();
 sg13g2_fill_1 FILLER_7_57 ();
 sg13g2_decap_4 FILLER_7_73 ();
 sg13g2_fill_1 FILLER_7_77 ();
 sg13g2_fill_2 FILLER_7_102 ();
 sg13g2_decap_8 FILLER_7_138 ();
 sg13g2_fill_1 FILLER_7_145 ();
 sg13g2_fill_1 FILLER_7_171 ();
 sg13g2_fill_2 FILLER_7_188 ();
 sg13g2_decap_8 FILLER_7_216 ();
 sg13g2_fill_2 FILLER_7_223 ();
 sg13g2_decap_8 FILLER_7_233 ();
 sg13g2_fill_2 FILLER_7_240 ();
 sg13g2_decap_4 FILLER_7_271 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_decap_8 FILLER_7_293 ();
 sg13g2_fill_2 FILLER_7_300 ();
 sg13g2_decap_4 FILLER_7_320 ();
 sg13g2_fill_2 FILLER_7_324 ();
 sg13g2_decap_4 FILLER_7_343 ();
 sg13g2_fill_1 FILLER_7_347 ();
 sg13g2_decap_4 FILLER_7_353 ();
 sg13g2_decap_4 FILLER_7_380 ();
 sg13g2_fill_1 FILLER_7_384 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_35 ();
 sg13g2_fill_1 FILLER_8_37 ();
 sg13g2_fill_2 FILLER_8_55 ();
 sg13g2_fill_1 FILLER_8_57 ();
 sg13g2_fill_2 FILLER_8_69 ();
 sg13g2_decap_8 FILLER_8_101 ();
 sg13g2_fill_1 FILLER_8_108 ();
 sg13g2_decap_8 FILLER_8_132 ();
 sg13g2_decap_8 FILLER_8_139 ();
 sg13g2_decap_4 FILLER_8_146 ();
 sg13g2_fill_2 FILLER_8_160 ();
 sg13g2_decap_4 FILLER_8_179 ();
 sg13g2_fill_1 FILLER_8_183 ();
 sg13g2_fill_1 FILLER_8_197 ();
 sg13g2_fill_2 FILLER_8_208 ();
 sg13g2_fill_2 FILLER_8_231 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_decap_4 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_298 ();
 sg13g2_fill_1 FILLER_8_300 ();
 sg13g2_decap_4 FILLER_8_323 ();
 sg13g2_fill_2 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_fill_2 FILLER_8_381 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_32 ();
 sg13g2_fill_2 FILLER_9_58 ();
 sg13g2_fill_2 FILLER_9_90 ();
 sg13g2_fill_1 FILLER_9_100 ();
 sg13g2_fill_1 FILLER_9_119 ();
 sg13g2_fill_2 FILLER_9_142 ();
 sg13g2_fill_1 FILLER_9_144 ();
 sg13g2_decap_4 FILLER_9_183 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_215 ();
 sg13g2_fill_2 FILLER_9_237 ();
 sg13g2_decap_4 FILLER_9_244 ();
 sg13g2_decap_8 FILLER_9_264 ();
 sg13g2_decap_4 FILLER_9_271 ();
 sg13g2_fill_2 FILLER_9_275 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_303 ();
 sg13g2_fill_1 FILLER_9_310 ();
 sg13g2_fill_2 FILLER_9_319 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_fill_2 FILLER_9_352 ();
 sg13g2_fill_1 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_360 ();
 sg13g2_decap_8 FILLER_9_367 ();
 sg13g2_fill_2 FILLER_9_374 ();
 sg13g2_decap_4 FILLER_9_382 ();
 sg13g2_fill_2 FILLER_9_386 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_fill_2 FILLER_10_46 ();
 sg13g2_decap_4 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_fill_2 FILLER_10_77 ();
 sg13g2_decap_4 FILLER_10_95 ();
 sg13g2_fill_2 FILLER_10_99 ();
 sg13g2_fill_2 FILLER_10_106 ();
 sg13g2_fill_1 FILLER_10_108 ();
 sg13g2_fill_1 FILLER_10_132 ();
 sg13g2_fill_2 FILLER_10_142 ();
 sg13g2_fill_1 FILLER_10_144 ();
 sg13g2_decap_4 FILLER_10_165 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_decap_8 FILLER_10_187 ();
 sg13g2_fill_1 FILLER_10_194 ();
 sg13g2_fill_2 FILLER_10_208 ();
 sg13g2_fill_1 FILLER_10_219 ();
 sg13g2_fill_1 FILLER_10_230 ();
 sg13g2_fill_2 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_243 ();
 sg13g2_fill_1 FILLER_10_339 ();
 sg13g2_fill_2 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_37 ();
 sg13g2_fill_2 FILLER_11_54 ();
 sg13g2_fill_2 FILLER_11_95 ();
 sg13g2_decap_4 FILLER_11_116 ();
 sg13g2_fill_1 FILLER_11_141 ();
 sg13g2_fill_2 FILLER_11_186 ();
 sg13g2_fill_2 FILLER_11_209 ();
 sg13g2_fill_1 FILLER_11_211 ();
 sg13g2_fill_2 FILLER_11_216 ();
 sg13g2_fill_2 FILLER_11_239 ();
 sg13g2_fill_1 FILLER_11_241 ();
 sg13g2_decap_4 FILLER_11_250 ();
 sg13g2_decap_8 FILLER_11_271 ();
 sg13g2_decap_4 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_fill_1 FILLER_11_329 ();
 sg13g2_fill_2 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_75 ();
 sg13g2_decap_8 FILLER_12_83 ();
 sg13g2_decap_8 FILLER_12_90 ();
 sg13g2_fill_2 FILLER_12_97 ();
 sg13g2_fill_1 FILLER_12_99 ();
 sg13g2_decap_4 FILLER_12_116 ();
 sg13g2_fill_2 FILLER_12_120 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_decap_8 FILLER_12_144 ();
 sg13g2_fill_1 FILLER_12_151 ();
 sg13g2_fill_2 FILLER_12_166 ();
 sg13g2_fill_2 FILLER_12_181 ();
 sg13g2_decap_8 FILLER_12_191 ();
 sg13g2_fill_1 FILLER_12_207 ();
 sg13g2_fill_2 FILLER_12_218 ();
 sg13g2_fill_1 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_fill_1 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_299 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_fill_1 FILLER_12_329 ();
 sg13g2_decap_4 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_fill_1 FILLER_12_352 ();
 sg13g2_decap_4 FILLER_12_359 ();
 sg13g2_fill_1 FILLER_12_386 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_2 FILLER_13_31 ();
 sg13g2_fill_2 FILLER_13_43 ();
 sg13g2_fill_2 FILLER_13_87 ();
 sg13g2_fill_2 FILLER_13_116 ();
 sg13g2_fill_1 FILLER_13_118 ();
 sg13g2_decap_4 FILLER_13_145 ();
 sg13g2_fill_1 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_186 ();
 sg13g2_fill_1 FILLER_13_199 ();
 sg13g2_fill_2 FILLER_13_208 ();
 sg13g2_fill_1 FILLER_13_210 ();
 sg13g2_fill_1 FILLER_13_233 ();
 sg13g2_decap_8 FILLER_13_243 ();
 sg13g2_decap_4 FILLER_13_292 ();
 sg13g2_fill_1 FILLER_13_296 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_fill_2 FILLER_13_354 ();
 sg13g2_decap_4 FILLER_13_385 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_11 ();
 sg13g2_fill_2 FILLER_14_37 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_1 FILLER_14_46 ();
 sg13g2_fill_2 FILLER_14_73 ();
 sg13g2_fill_2 FILLER_14_84 ();
 sg13g2_decap_4 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_103 ();
 sg13g2_decap_4 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_120 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_4 FILLER_14_147 ();
 sg13g2_fill_1 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_159 ();
 sg13g2_decap_4 FILLER_14_166 ();
 sg13g2_fill_1 FILLER_14_180 ();
 sg13g2_decap_4 FILLER_14_194 ();
 sg13g2_fill_1 FILLER_14_198 ();
 sg13g2_fill_1 FILLER_14_207 ();
 sg13g2_fill_1 FILLER_14_213 ();
 sg13g2_decap_4 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_232 ();
 sg13g2_fill_2 FILLER_14_238 ();
 sg13g2_decap_4 FILLER_14_257 ();
 sg13g2_decap_4 FILLER_14_301 ();
 sg13g2_decap_4 FILLER_14_328 ();
 sg13g2_fill_2 FILLER_14_332 ();
 sg13g2_decap_4 FILLER_14_346 ();
 sg13g2_fill_1 FILLER_14_350 ();
 sg13g2_fill_2 FILLER_14_363 ();
 sg13g2_fill_1 FILLER_14_365 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_2 FILLER_15_26 ();
 sg13g2_fill_1 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_53 ();
 sg13g2_fill_1 FILLER_15_55 ();
 sg13g2_fill_2 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_111 ();
 sg13g2_fill_2 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_177 ();
 sg13g2_fill_1 FILLER_15_179 ();
 sg13g2_fill_2 FILLER_15_187 ();
 sg13g2_decap_8 FILLER_15_205 ();
 sg13g2_decap_4 FILLER_15_228 ();
 sg13g2_fill_2 FILLER_15_232 ();
 sg13g2_fill_2 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_fill_1 FILLER_15_357 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_fill_1 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_25 ();
 sg13g2_fill_2 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_88 ();
 sg13g2_fill_2 FILLER_16_97 ();
 sg13g2_fill_1 FILLER_16_132 ();
 sg13g2_fill_2 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_153 ();
 sg13g2_decap_4 FILLER_16_172 ();
 sg13g2_fill_2 FILLER_16_176 ();
 sg13g2_decap_4 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_202 ();
 sg13g2_fill_2 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_decap_4 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_fill_2 FILLER_16_298 ();
 sg13g2_fill_1 FILLER_16_300 ();
 sg13g2_decap_4 FILLER_16_307 ();
 sg13g2_fill_1 FILLER_16_311 ();
 sg13g2_decap_4 FILLER_16_324 ();
 sg13g2_fill_1 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_fill_2 FILLER_16_351 ();
 sg13g2_fill_2 FILLER_16_361 ();
 sg13g2_fill_2 FILLER_16_391 ();
 sg13g2_fill_1 FILLER_16_393 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_2 FILLER_17_47 ();
 sg13g2_fill_2 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_86 ();
 sg13g2_fill_2 FILLER_17_96 ();
 sg13g2_decap_4 FILLER_17_105 ();
 sg13g2_fill_1 FILLER_17_109 ();
 sg13g2_fill_2 FILLER_17_115 ();
 sg13g2_fill_1 FILLER_17_117 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_fill_1 FILLER_17_134 ();
 sg13g2_fill_2 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_155 ();
 sg13g2_decap_8 FILLER_17_160 ();
 sg13g2_fill_1 FILLER_17_167 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_decap_4 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_248 ();
 sg13g2_fill_1 FILLER_17_255 ();
 sg13g2_fill_1 FILLER_17_262 ();
 sg13g2_fill_1 FILLER_17_275 ();
 sg13g2_fill_1 FILLER_17_288 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_fill_2 FILLER_17_328 ();
 sg13g2_decap_4 FILLER_17_347 ();
 sg13g2_fill_1 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_4 FILLER_17_381 ();
 sg13g2_fill_1 FILLER_17_390 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_32 ();
 sg13g2_fill_2 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_45 ();
 sg13g2_fill_2 FILLER_18_51 ();
 sg13g2_fill_1 FILLER_18_53 ();
 sg13g2_fill_2 FILLER_18_62 ();
 sg13g2_fill_1 FILLER_18_69 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_153 ();
 sg13g2_fill_1 FILLER_18_155 ();
 sg13g2_fill_2 FILLER_18_174 ();
 sg13g2_fill_2 FILLER_18_188 ();
 sg13g2_decap_8 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_226 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_251 ();
 sg13g2_fill_1 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_4 FILLER_18_284 ();
 sg13g2_fill_2 FILLER_18_288 ();
 sg13g2_fill_2 FILLER_18_302 ();
 sg13g2_fill_1 FILLER_18_304 ();
 sg13g2_decap_4 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_330 ();
 sg13g2_fill_2 FILLER_18_371 ();
 sg13g2_fill_1 FILLER_18_373 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_1 FILLER_19_26 ();
 sg13g2_fill_2 FILLER_19_67 ();
 sg13g2_fill_1 FILLER_19_100 ();
 sg13g2_fill_1 FILLER_19_106 ();
 sg13g2_fill_2 FILLER_19_138 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_156 ();
 sg13g2_decap_4 FILLER_19_195 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_decap_4 FILLER_19_205 ();
 sg13g2_fill_1 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_236 ();
 sg13g2_decap_8 FILLER_19_243 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_decap_8 FILLER_19_272 ();
 sg13g2_decap_4 FILLER_19_302 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_334 ();
 sg13g2_decap_4 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_350 ();
 sg13g2_fill_2 FILLER_19_362 ();
 sg13g2_fill_2 FILLER_19_373 ();
 sg13g2_fill_1 FILLER_19_375 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_decap_8 FILLER_20_29 ();
 sg13g2_decap_8 FILLER_20_79 ();
 sg13g2_fill_1 FILLER_20_86 ();
 sg13g2_decap_4 FILLER_20_100 ();
 sg13g2_fill_1 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_139 ();
 sg13g2_fill_2 FILLER_20_146 ();
 sg13g2_fill_1 FILLER_20_148 ();
 sg13g2_fill_1 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_176 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_decap_8 FILLER_20_205 ();
 sg13g2_fill_2 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_219 ();
 sg13g2_decap_4 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_fill_2 FILLER_20_311 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_fill_2 FILLER_20_326 ();
 sg13g2_fill_1 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_fill_1 FILLER_20_348 ();
 sg13g2_decap_4 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_25 ();
 sg13g2_fill_1 FILLER_21_27 ();
 sg13g2_fill_1 FILLER_21_41 ();
 sg13g2_fill_1 FILLER_21_47 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_fill_1 FILLER_21_68 ();
 sg13g2_fill_2 FILLER_21_74 ();
 sg13g2_fill_1 FILLER_21_76 ();
 sg13g2_decap_4 FILLER_21_86 ();
 sg13g2_decap_4 FILLER_21_106 ();
 sg13g2_fill_1 FILLER_21_114 ();
 sg13g2_fill_1 FILLER_21_118 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_fill_2 FILLER_21_145 ();
 sg13g2_decap_8 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_4 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_decap_4 FILLER_21_251 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_269 ();
 sg13g2_fill_2 FILLER_21_287 ();
 sg13g2_fill_1 FILLER_21_289 ();
 sg13g2_fill_2 FILLER_21_302 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_fill_1 FILLER_21_358 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_1 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_70 ();
 sg13g2_fill_2 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_96 ();
 sg13g2_decap_8 FILLER_22_103 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_131 ();
 sg13g2_decap_4 FILLER_22_145 ();
 sg13g2_fill_2 FILLER_22_159 ();
 sg13g2_fill_2 FILLER_22_187 ();
 sg13g2_fill_2 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_220 ();
 sg13g2_fill_1 FILLER_22_222 ();
 sg13g2_fill_2 FILLER_22_232 ();
 sg13g2_fill_1 FILLER_22_234 ();
 sg13g2_fill_2 FILLER_22_251 ();
 sg13g2_fill_1 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_275 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_302 ();
 sg13g2_fill_2 FILLER_22_332 ();
 sg13g2_decap_4 FILLER_22_357 ();
 sg13g2_decap_4 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_1 FILLER_23_26 ();
 sg13g2_fill_2 FILLER_23_71 ();
 sg13g2_fill_1 FILLER_23_73 ();
 sg13g2_fill_2 FILLER_23_114 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_122 ();
 sg13g2_fill_2 FILLER_23_134 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_fill_2 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_162 ();
 sg13g2_fill_1 FILLER_23_169 ();
 sg13g2_decap_4 FILLER_23_200 ();
 sg13g2_decap_4 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_decap_4 FILLER_23_244 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_decap_4 FILLER_23_263 ();
 sg13g2_fill_2 FILLER_23_291 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_decap_4 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_314 ();
 sg13g2_fill_2 FILLER_23_327 ();
 sg13g2_fill_1 FILLER_23_329 ();
 sg13g2_fill_2 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_fill_1 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_44 ();
 sg13g2_fill_1 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_110 ();
 sg13g2_fill_1 FILLER_24_129 ();
 sg13g2_decap_8 FILLER_24_143 ();
 sg13g2_decap_4 FILLER_24_167 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_fill_2 FILLER_24_178 ();
 sg13g2_decap_4 FILLER_24_214 ();
 sg13g2_fill_2 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_243 ();
 sg13g2_fill_2 FILLER_24_247 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_fill_2 FILLER_24_340 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_48 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_fill_1 FILLER_25_116 ();
 sg13g2_decap_4 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_fill_1 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_253 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_288 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_315 ();
 sg13g2_fill_2 FILLER_25_333 ();
 sg13g2_fill_1 FILLER_25_362 ();
 sg13g2_fill_1 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_386 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_4 FILLER_26_96 ();
 sg13g2_fill_2 FILLER_26_100 ();
 sg13g2_fill_1 FILLER_26_144 ();
 sg13g2_fill_2 FILLER_26_157 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_182 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_244 ();
 sg13g2_fill_2 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_275 ();
 sg13g2_decap_4 FILLER_26_311 ();
 sg13g2_decap_8 FILLER_26_321 ();
 sg13g2_fill_1 FILLER_26_328 ();
 sg13g2_decap_4 FILLER_26_352 ();
 sg13g2_fill_1 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_15 ();
 sg13g2_fill_2 FILLER_27_31 ();
 sg13g2_fill_1 FILLER_27_53 ();
 sg13g2_fill_2 FILLER_27_64 ();
 sg13g2_fill_2 FILLER_27_71 ();
 sg13g2_fill_2 FILLER_27_95 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_146 ();
 sg13g2_fill_2 FILLER_27_157 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_decap_4 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_decap_4 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_287 ();
 sg13g2_decap_4 FILLER_27_352 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_28_26 ();
 sg13g2_fill_2 FILLER_28_101 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_114 ();
 sg13g2_fill_2 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_135 ();
 sg13g2_fill_2 FILLER_28_178 ();
 sg13g2_fill_1 FILLER_28_180 ();
 sg13g2_decap_4 FILLER_28_189 ();
 sg13g2_fill_1 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_247 ();
 sg13g2_fill_2 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_decap_4 FILLER_28_297 ();
 sg13g2_decap_8 FILLER_28_309 ();
 sg13g2_decap_8 FILLER_28_316 ();
 sg13g2_decap_8 FILLER_28_323 ();
 sg13g2_decap_4 FILLER_28_330 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_fill_1 FILLER_28_338 ();
 sg13g2_decap_4 FILLER_28_345 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_fill_2 FILLER_29_146 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_232 ();
 sg13g2_decap_4 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_243 ();
 sg13g2_decap_4 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_37 ();
 sg13g2_fill_1 FILLER_30_60 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_fill_1 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_111 ();
 sg13g2_fill_2 FILLER_30_128 ();
 sg13g2_fill_1 FILLER_30_130 ();
 sg13g2_fill_1 FILLER_30_145 ();
 sg13g2_fill_1 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_185 ();
 sg13g2_fill_1 FILLER_30_190 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_248 ();
 sg13g2_fill_1 FILLER_30_255 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_2 FILLER_30_275 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_fill_2 FILLER_30_380 ();
 sg13g2_fill_2 FILLER_31_26 ();
 sg13g2_fill_2 FILLER_31_87 ();
 sg13g2_fill_2 FILLER_31_99 ();
 sg13g2_fill_2 FILLER_31_138 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_fill_1 FILLER_31_148 ();
 sg13g2_fill_1 FILLER_31_178 ();
 sg13g2_fill_2 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_decap_4 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_326 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_32_68 ();
 sg13g2_fill_1 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_84 ();
 sg13g2_fill_1 FILLER_32_101 ();
 sg13g2_fill_2 FILLER_32_130 ();
 sg13g2_fill_2 FILLER_32_153 ();
 sg13g2_fill_2 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_fill_2 FILLER_32_183 ();
 sg13g2_fill_1 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_decap_8 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_decap_4 FILLER_32_232 ();
 sg13g2_fill_2 FILLER_32_252 ();
 sg13g2_fill_1 FILLER_32_262 ();
 sg13g2_fill_1 FILLER_32_281 ();
 sg13g2_fill_2 FILLER_32_286 ();
 sg13g2_fill_1 FILLER_32_305 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_fill_2 FILLER_32_317 ();
 sg13g2_fill_2 FILLER_32_398 ();
 sg13g2_fill_2 FILLER_33_26 ();
 sg13g2_fill_1 FILLER_33_62 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_173 ();
 sg13g2_fill_2 FILLER_33_181 ();
 sg13g2_fill_1 FILLER_33_183 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_202 ();
 sg13g2_decap_4 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_41 ();
 sg13g2_fill_2 FILLER_34_60 ();
 sg13g2_fill_2 FILLER_34_67 ();
 sg13g2_fill_1 FILLER_34_69 ();
 sg13g2_fill_2 FILLER_34_75 ();
 sg13g2_fill_2 FILLER_34_82 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_239 ();
 sg13g2_decap_4 FILLER_34_246 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_decap_8 FILLER_34_264 ();
 sg13g2_decap_4 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_fill_2 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_34_314 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_35_102 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_223 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_fill_2 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_319 ();
 sg13g2_fill_2 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_fill_2 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_fill_1 FILLER_36_118 ();
 sg13g2_fill_1 FILLER_36_205 ();
 sg13g2_fill_1 FILLER_36_212 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_241 ();
 sg13g2_decap_4 FILLER_36_272 ();
 sg13g2_fill_1 FILLER_36_320 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_373 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_30 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_fill_2 FILLER_37_166 ();
 sg13g2_fill_1 FILLER_37_188 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_1 FILLER_37_217 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_decap_4 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_271 ();
 sg13g2_fill_2 FILLER_37_282 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_fill_2 FILLER_37_336 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_fill_1 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_61 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_fill_2 FILLER_38_282 ();
 sg13g2_fill_1 FILLER_38_284 ();
 sg13g2_fill_2 FILLER_38_332 ();
 sg13g2_fill_2 FILLER_38_359 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net75;
 assign uio_oe[1] = net76;
 assign uio_oe[2] = net77;
 assign uio_oe[3] = net78;
 assign uio_oe[4] = net79;
 assign uio_oe[5] = net80;
 assign uio_oe[6] = net81;
 assign uio_oe[7] = net82;
 assign uio_out[6] = net5;
 assign uio_out[7] = net6;
 assign uo_out[7] = net7;
endmodule

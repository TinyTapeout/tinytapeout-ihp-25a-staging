module tt_um_rebeccargb_styler (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire clknet_0_clk;
 wire \bitmapIn[0] ;
 wire \bitmapIn[10] ;
 wire \bitmapIn[11] ;
 wire \bitmapIn[12] ;
 wire \bitmapIn[13] ;
 wire \bitmapIn[14] ;
 wire \bitmapIn[15] ;
 wire \bitmapIn[1] ;
 wire \bitmapIn[2] ;
 wire \bitmapIn[3] ;
 wire \bitmapIn[4] ;
 wire \bitmapIn[5] ;
 wire \bitmapIn[6] ;
 wire \bitmapIn[7] ;
 wire \bitmapIn[8] ;
 wire \bitmapIn[9] ;
 wire \ctrl[0] ;
 wire \ctrl[1] ;
 wire \ctrl[2] ;
 wire \ctrl[3] ;
 wire \ctrl[4] ;
 wire \ctrl[5] ;
 wire \ctrl[6] ;
 wire \ctrl[7] ;
 wire \s.alternate ;
 wire \s.blink ;
 wire \s.bold ;
 wire \s.dottedOverline ;
 wire \s.dottedStrikethru ;
 wire \s.dottedUnderline ;
 wire \s.doubleOverline ;
 wire \s.doubleStrikethru ;
 wire \s.doubleUnderline ;
 wire \s.faint ;
 wire \s.hidden ;
 wire \s.inv.xPostMirror ;
 wire \s.inverse ;
 wire \s.italic ;
 wire \s.lg.overline ;
 wire \s.lg.s0[0] ;
 wire \s.lg.s0[1] ;
 wire \s.lg.s0[2] ;
 wire \s.lg.s0[3] ;
 wire \s.lg.strikethru ;
 wire \s.lg.underline ;
 wire \s.lg.yPostMirror ;
 wire \s.lg.yPreMirror ;
 wire \s.lg.yoffset ;
 wire \s.lg.yscale ;
 wire \s.reverseItalic ;
 wire \s.sty.xPreMirror ;
 wire \s.sty.xoffset ;
 wire \s.sty.xscale ;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;

 sg13g2_inv_1 _0730_ (.Y(_0059_),
    .A(net85));
 sg13g2_inv_1 _0731_ (.Y(_0060_),
    .A(net16));
 sg13g2_inv_1 _0732_ (.Y(_0061_),
    .A(net89));
 sg13g2_inv_1 _0733_ (.Y(_0062_),
    .A(net15));
 sg13g2_inv_1 _0734_ (.Y(_0063_),
    .A(net84));
 sg13g2_inv_1 _0735_ (.Y(_0064_),
    .A(net14));
 sg13g2_inv_1 _0736_ (.Y(_0065_),
    .A(net78));
 sg13g2_inv_1 _0737_ (.Y(_0066_),
    .A(net13));
 sg13g2_inv_1 _0738_ (.Y(_0067_),
    .A(net91));
 sg13g2_inv_1 _0739_ (.Y(_0068_),
    .A(net12));
 sg13g2_inv_1 _0740_ (.Y(_0069_),
    .A(net87));
 sg13g2_inv_1 _0741_ (.Y(_0070_),
    .A(net11));
 sg13g2_inv_1 _0742_ (.Y(_0071_),
    .A(net93));
 sg13g2_inv_1 _0743_ (.Y(_0072_),
    .A(net10));
 sg13g2_inv_1 _0744_ (.Y(_0073_),
    .A(net95));
 sg13g2_inv_1 _0745_ (.Y(_0074_),
    .A(net9));
 sg13g2_inv_1 _0746_ (.Y(_0075_),
    .A(net90));
 sg13g2_inv_1 _0747_ (.Y(_0076_),
    .A(net94));
 sg13g2_inv_1 _0748_ (.Y(_0077_),
    .A(net81));
 sg13g2_inv_1 _0749_ (.Y(_0078_),
    .A(net77));
 sg13g2_inv_1 _0750_ (.Y(_0079_),
    .A(net111));
 sg13g2_inv_1 _0751_ (.Y(_0080_),
    .A(net108));
 sg13g2_inv_1 _0752_ (.Y(_0081_),
    .A(net80));
 sg13g2_inv_1 _0753_ (.Y(_0082_),
    .A(net79));
 sg13g2_inv_1 _0754_ (.Y(_0083_),
    .A(net118));
 sg13g2_inv_1 _0755_ (.Y(_0084_),
    .A(net72));
 sg13g2_inv_1 _0756_ (.Y(_0085_),
    .A(net272));
 sg13g2_inv_2 _0757_ (.Y(_0086_),
    .A(net275));
 sg13g2_inv_1 _0758_ (.Y(_0087_),
    .A(net116));
 sg13g2_inv_1 _0759_ (.Y(_0088_),
    .A(net115));
 sg13g2_inv_1 _0760_ (.Y(_0089_),
    .A(net278));
 sg13g2_inv_1 _0761_ (.Y(_0090_),
    .A(net280));
 sg13g2_inv_1 _0762_ (.Y(_0091_),
    .A(net86));
 sg13g2_inv_1 _0763_ (.Y(_0092_),
    .A(net96));
 sg13g2_inv_1 _0764_ (.Y(_0093_),
    .A(net74));
 sg13g2_inv_1 _0765_ (.Y(_0094_),
    .A(net83));
 sg13g2_inv_1 _0766_ (.Y(_0095_),
    .A(net73));
 sg13g2_inv_1 _0767_ (.Y(_0096_),
    .A(net75));
 sg13g2_inv_1 _0768_ (.Y(_0097_),
    .A(net71));
 sg13g2_inv_1 _0769_ (.Y(_0098_),
    .A(net70));
 sg13g2_inv_1 _0770_ (.Y(_0099_),
    .A(\ctrl[4] ));
 sg13g2_inv_1 _0771_ (.Y(_0100_),
    .A(net105));
 sg13g2_inv_1 _0772_ (.Y(_0101_),
    .A(net107));
 sg13g2_inv_1 _0773_ (.Y(_0102_),
    .A(net101));
 sg13g2_inv_1 _0774_ (.Y(_0103_),
    .A(net97));
 sg13g2_inv_1 _0775_ (.Y(_0104_),
    .A(net88));
 sg13g2_inv_1 _0776_ (.Y(_0105_),
    .A(net3));
 sg13g2_inv_1 _0777_ (.Y(_0106_),
    .A(net5));
 sg13g2_inv_2 _0778_ (.Y(uio_oe[7]),
    .A(net7));
 sg13g2_nand2_1 _0779_ (.Y(_0107_),
    .A(_0102_),
    .B(_0103_));
 sg13g2_nand4_1 _0780_ (.B(\s.lg.s0[3] ),
    .C(\s.lg.s0[2] ),
    .A(\ctrl[0] ),
    .Y(_0108_),
    .D(_0107_));
 sg13g2_nand3_1 _0781_ (.B(_0100_),
    .C(_0101_),
    .A(\ctrl[1] ),
    .Y(_0109_));
 sg13g2_a21oi_1 _0782_ (.A1(\s.lg.s0[1] ),
    .A2(\s.lg.s0[0] ),
    .Y(_0110_),
    .B1(_0109_));
 sg13g2_o21ai_1 _0783_ (.B1(_0108_),
    .Y(_0111_),
    .A1(\ctrl[1] ),
    .A2(\ctrl[0] ));
 sg13g2_nor2_1 _0784_ (.A(\ctrl[7] ),
    .B(net5),
    .Y(_0112_));
 sg13g2_a21oi_1 _0785_ (.A1(\ctrl[7] ),
    .A2(net4),
    .Y(_0113_),
    .B1(_0112_));
 sg13g2_nand2_1 _0786_ (.Y(_0114_),
    .A(\ctrl[3] ),
    .B(net6));
 sg13g2_a21oi_1 _0787_ (.A1(\ctrl[2] ),
    .A2(_0113_),
    .Y(_0115_),
    .B1(_0114_));
 sg13g2_o21ai_1 _0788_ (.B1(_0115_),
    .Y(_0116_),
    .A1(_0110_),
    .A2(_0111_));
 sg13g2_a21oi_1 _0789_ (.A1(\ctrl[5] ),
    .A2(_0106_),
    .Y(_0117_),
    .B1(_0077_));
 sg13g2_xnor2_1 _0790_ (.Y(_0118_),
    .A(_0076_),
    .B(_0117_));
 sg13g2_xnor2_1 _0791_ (.Y(_0119_),
    .A(_0116_),
    .B(_0118_));
 sg13g2_nand3_1 _0792_ (.B(\ctrl[5] ),
    .C(net5),
    .A(\s.blink ),
    .Y(_0120_));
 sg13g2_and2_1 _0793_ (.A(_0075_),
    .B(_0120_),
    .X(_0121_));
 sg13g2_nand2_1 _0794_ (.Y(_0122_),
    .A(_0075_),
    .B(_0120_));
 sg13g2_xnor2_1 _0795_ (.Y(_0123_),
    .A(\s.lg.yPostMirror ),
    .B(\s.lg.s0[1] ));
 sg13g2_xnor2_1 _0796_ (.Y(_0124_),
    .A(\s.lg.yPostMirror ),
    .B(\s.lg.s0[2] ));
 sg13g2_xor2_1 _0797_ (.B(\s.lg.s0[2] ),
    .A(\s.lg.yPostMirror ),
    .X(_0125_));
 sg13g2_mux2_2 _0798_ (.A0(_0123_),
    .A1(_0124_),
    .S(\s.lg.yscale ),
    .X(_0126_));
 sg13g2_xnor2_1 _0799_ (.Y(_0127_),
    .A(\s.lg.yPostMirror ),
    .B(\s.lg.s0[0] ));
 sg13g2_mux2_2 _0800_ (.A0(_0123_),
    .A1(_0127_),
    .S(_0087_),
    .X(_0128_));
 sg13g2_xnor2_1 _0801_ (.Y(_0129_),
    .A(\s.lg.yPostMirror ),
    .B(\s.lg.s0[3] ));
 sg13g2_xor2_1 _0802_ (.B(\s.lg.s0[3] ),
    .A(\s.lg.yPostMirror ),
    .X(_0130_));
 sg13g2_and3_2 _0803_ (.X(_0131_),
    .A(\s.lg.yoffset ),
    .B(_0001_),
    .C(_0130_));
 sg13g2_nand3_1 _0804_ (.B(_0001_),
    .C(_0130_),
    .A(\s.lg.yoffset ),
    .Y(_0132_));
 sg13g2_a21oi_2 _0805_ (.B1(\s.lg.yoffset ),
    .Y(_0133_),
    .A2(_0130_),
    .A1(_0001_));
 sg13g2_a21o_2 _0806_ (.A2(_0130_),
    .A1(_0001_),
    .B1(\s.lg.yoffset ),
    .X(_0134_));
 sg13g2_nand3_1 _0807_ (.B(_0001_),
    .C(_0130_),
    .A(_0088_),
    .Y(_0135_));
 sg13g2_a21o_1 _0808_ (.A2(_0130_),
    .A1(_0001_),
    .B1(_0088_),
    .X(_0136_));
 sg13g2_nor2_2 _0809_ (.A(_0131_),
    .B(_0133_),
    .Y(_0137_));
 sg13g2_nand2_1 _0810_ (.Y(_0138_),
    .A(_0132_),
    .B(_0134_));
 sg13g2_nor2_1 _0811_ (.A(\s.dottedStrikethru ),
    .B(\s.lg.strikethru ),
    .Y(_0139_));
 sg13g2_nor3_1 _0812_ (.A(_0126_),
    .B(_0128_),
    .C(_0139_),
    .Y(_0140_));
 sg13g2_nand2_1 _0813_ (.Y(_0141_),
    .A(\s.doubleStrikethru ),
    .B(_0067_));
 sg13g2_nor2b_1 _0814_ (.A(_0128_),
    .B_N(_0126_),
    .Y(_0142_));
 sg13g2_a22oi_1 _0815_ (.Y(_0143_),
    .B1(_0142_),
    .B2(\s.doubleStrikethru ),
    .A2(_0140_),
    .A1(net237));
 sg13g2_nand2_1 _0816_ (.Y(_0144_),
    .A(_0126_),
    .B(_0128_));
 sg13g2_a21o_1 _0817_ (.A2(_0144_),
    .A1(_0067_),
    .B1(net237),
    .X(_0145_));
 sg13g2_mux2_1 _0818_ (.A0(_0124_),
    .A1(_0129_),
    .S(\s.lg.yscale ),
    .X(_0146_));
 sg13g2_mux2_1 _0819_ (.A0(_0125_),
    .A1(_0130_),
    .S(\s.lg.yscale ),
    .X(_0147_));
 sg13g2_nor2b_1 _0820_ (.A(_0126_),
    .B_N(_0128_),
    .Y(_0148_));
 sg13g2_nand2b_1 _0821_ (.Y(_0149_),
    .B(_0128_),
    .A_N(_0126_));
 sg13g2_o21ai_1 _0822_ (.B1(net250),
    .Y(_0150_),
    .A1(_0141_),
    .A2(_0148_));
 sg13g2_a21oi_1 _0823_ (.A1(net256),
    .A2(net255),
    .Y(_0151_),
    .B1(net253));
 sg13g2_nand2b_1 _0824_ (.Y(_0152_),
    .B(\ctrl[4] ),
    .A_N(net233));
 sg13g2_a21oi_2 _0825_ (.B1(net250),
    .Y(_0153_),
    .A2(_0134_),
    .A1(_0132_));
 sg13g2_nand3_1 _0826_ (.B(net255),
    .C(net252),
    .A(net256),
    .Y(_0154_));
 sg13g2_a221oi_1 _0827_ (.B2(_0150_),
    .C1(_0152_),
    .B1(_0145_),
    .A1(_0141_),
    .Y(_0155_),
    .A2(_0143_));
 sg13g2_nand2_1 _0828_ (.Y(_0156_),
    .A(\s.dottedStrikethru ),
    .B(_0155_));
 sg13g2_nand2_1 _0829_ (.Y(_0157_),
    .A(_0061_),
    .B(_0128_));
 sg13g2_nand3_1 _0830_ (.B(_0149_),
    .C(_0157_),
    .A(\s.doubleOverline ),
    .Y(_0158_));
 sg13g2_nor2_1 _0831_ (.A(\s.lg.overline ),
    .B(\s.dottedOverline ),
    .Y(_0159_));
 sg13g2_o21ai_1 _0832_ (.B1(_0059_),
    .Y(_0160_),
    .A1(_0144_),
    .A2(_0159_));
 sg13g2_and4_1 _0833_ (.A(\ctrl[4] ),
    .B(_0153_),
    .C(_0158_),
    .D(_0160_),
    .X(_0161_));
 sg13g2_a21oi_1 _0834_ (.A1(\s.dottedOverline ),
    .A2(_0161_),
    .Y(_0162_),
    .B1(\s.faint ));
 sg13g2_a21oi_1 _0835_ (.A1(\s.lg.underline ),
    .A2(_0126_),
    .Y(_0163_),
    .B1(_0128_));
 sg13g2_nand2_1 _0836_ (.Y(_0164_),
    .A(_0069_),
    .B(_0073_));
 sg13g2_a21oi_1 _0837_ (.A1(_0142_),
    .A2(_0164_),
    .Y(_0165_),
    .B1(\s.doubleUnderline ));
 sg13g2_o21ai_1 _0838_ (.B1(net233),
    .Y(_0166_),
    .A1(_0071_),
    .A2(_0163_));
 sg13g2_nor3_1 _0839_ (.A(_0099_),
    .B(_0165_),
    .C(_0166_),
    .Y(_0167_));
 sg13g2_nand2_1 _0840_ (.Y(_0168_),
    .A(\s.dottedUnderline ),
    .B(_0167_));
 sg13g2_and3_1 _0841_ (.X(_0169_),
    .A(_0156_),
    .B(_0162_),
    .C(_0168_));
 sg13g2_nand3_1 _0842_ (.B(_0162_),
    .C(_0168_),
    .A(_0156_),
    .Y(_0170_));
 sg13g2_nor2b_1 _0843_ (.A(\ctrl[7] ),
    .B_N(net4),
    .Y(_0171_));
 sg13g2_xnor2_1 _0844_ (.Y(_0172_),
    .A(_0127_),
    .B(_0171_));
 sg13g2_xor2_1 _0845_ (.B(_0171_),
    .A(_0127_),
    .X(_0173_));
 sg13g2_a21oi_2 _0846_ (.B1(_0122_),
    .Y(_0174_),
    .A2(_0173_),
    .A1(_0170_));
 sg13g2_o21ai_1 _0847_ (.B1(_0121_),
    .Y(_0175_),
    .A1(_0169_),
    .A2(_0172_));
 sg13g2_nor2b_2 _0848_ (.A(\s.italic ),
    .B_N(\s.reverseItalic ),
    .Y(_0176_));
 sg13g2_nand2_1 _0849_ (.Y(_0177_),
    .A(\s.reverseItalic ),
    .B(_0080_));
 sg13g2_a21oi_1 _0850_ (.A1(_0135_),
    .A2(_0136_),
    .Y(_0178_),
    .B1(net246));
 sg13g2_nand3_1 _0851_ (.B(_0134_),
    .C(_0176_),
    .A(_0132_),
    .Y(_0179_));
 sg13g2_nor2b_2 _0852_ (.A(\s.reverseItalic ),
    .B_N(\s.italic ),
    .Y(_0180_));
 sg13g2_nand2_2 _0853_ (.Y(_0181_),
    .A(_0079_),
    .B(\s.italic ));
 sg13g2_nor2_2 _0854_ (.A(_0176_),
    .B(_0180_),
    .Y(_0182_));
 sg13g2_nand2_2 _0855_ (.Y(_0183_),
    .A(net246),
    .B(_0181_));
 sg13g2_nor2_1 _0856_ (.A(\bitmapIn[9] ),
    .B(net273),
    .Y(_0184_));
 sg13g2_a21oi_2 _0857_ (.B1(_0184_),
    .Y(_0185_),
    .A2(_0092_),
    .A1(net274));
 sg13g2_nor2_1 _0858_ (.A(_0183_),
    .B(_0185_),
    .Y(_0186_));
 sg13g2_nor2_1 _0859_ (.A(\bitmapIn[8] ),
    .B(net273),
    .Y(_0187_));
 sg13g2_a21oi_2 _0860_ (.B1(_0187_),
    .Y(_0188_),
    .A2(_0091_),
    .A1(net273));
 sg13g2_nand2_1 _0861_ (.Y(_0189_),
    .A(\bitmapIn[8] ),
    .B(net273));
 sg13g2_o21ai_1 _0862_ (.B1(_0189_),
    .Y(_0190_),
    .A1(net273),
    .A2(_0091_));
 sg13g2_inv_1 _0863_ (.Y(_0191_),
    .A(net245));
 sg13g2_a21o_1 _0864_ (.A2(net245),
    .A1(net251),
    .B1(net247),
    .X(_0192_));
 sg13g2_a21oi_1 _0865_ (.A1(net249),
    .A2(_0188_),
    .Y(_0193_),
    .B1(_0192_));
 sg13g2_o21ai_1 _0866_ (.B1(net228),
    .Y(_0194_),
    .A1(_0186_),
    .A2(_0193_));
 sg13g2_nor2_2 _0867_ (.A(_0153_),
    .B(_0181_),
    .Y(_0195_));
 sg13g2_nand2_2 _0868_ (.Y(_0196_),
    .A(_0154_),
    .B(_0180_));
 sg13g2_nor2_1 _0869_ (.A(\bitmapIn[10] ),
    .B(net276),
    .Y(_0197_));
 sg13g2_a21oi_2 _0870_ (.B1(_0197_),
    .Y(_0198_),
    .A2(_0093_),
    .A1(net273));
 sg13g2_and3_1 _0871_ (.X(_0199_),
    .A(net256),
    .B(net255),
    .C(_0198_));
 sg13g2_and2_1 _0872_ (.A(net251),
    .B(_0185_),
    .X(_0200_));
 sg13g2_a221oi_1 _0873_ (.B2(net234),
    .C1(_0200_),
    .B1(_0198_),
    .A1(net230),
    .Y(_0201_),
    .A2(_0188_));
 sg13g2_nor2_2 _0874_ (.A(_0154_),
    .B(_0181_),
    .Y(_0202_));
 sg13g2_nand4_1 _0875_ (.B(net255),
    .C(net254),
    .A(net256),
    .Y(_0203_),
    .D(_0180_));
 sg13g2_nor2_1 _0876_ (.A(\bitmapIn[11] ),
    .B(net276),
    .Y(_0204_));
 sg13g2_a21oi_2 _0877_ (.B1(_0204_),
    .Y(_0205_),
    .A2(_0094_),
    .A1(net276));
 sg13g2_nor2_1 _0878_ (.A(_0203_),
    .B(_0205_),
    .Y(_0206_));
 sg13g2_nand2_1 _0879_ (.Y(_0207_),
    .A(net230),
    .B(_0198_));
 sg13g2_nor2_1 _0880_ (.A(net228),
    .B(_0200_),
    .Y(_0208_));
 sg13g2_a221oi_1 _0881_ (.B2(_0208_),
    .C1(_0206_),
    .B1(_0207_),
    .A1(_0195_),
    .Y(_0209_),
    .A2(_0201_));
 sg13g2_and2_1 _0882_ (.A(_0194_),
    .B(_0209_),
    .X(_0210_));
 sg13g2_nand2b_1 _0883_ (.Y(_0211_),
    .B(_0182_),
    .A_N(_0188_));
 sg13g2_nand4_1 _0884_ (.B(_0136_),
    .C(net248),
    .A(net256),
    .Y(_0212_),
    .D(_0190_));
 sg13g2_nand2_1 _0885_ (.Y(_0213_),
    .A(\bitmapIn[9] ),
    .B(net273));
 sg13g2_o21ai_1 _0886_ (.B1(_0213_),
    .Y(_0214_),
    .A1(net273),
    .A2(_0092_));
 sg13g2_inv_1 _0887_ (.Y(_0215_),
    .A(_0214_));
 sg13g2_a21oi_1 _0888_ (.A1(net253),
    .A2(_0214_),
    .Y(_0216_),
    .B1(net246));
 sg13g2_o21ai_1 _0889_ (.B1(_0212_),
    .Y(_0217_),
    .A1(_0178_),
    .A2(_0216_));
 sg13g2_and2_1 _0890_ (.A(net252),
    .B(_0188_),
    .X(_0218_));
 sg13g2_a21o_1 _0891_ (.A2(_0185_),
    .A1(net233),
    .B1(_0218_),
    .X(_0219_));
 sg13g2_a22oi_1 _0892_ (.Y(_0220_),
    .B1(_0219_),
    .B2(net229),
    .A2(_0217_),
    .A1(_0211_));
 sg13g2_nor2_1 _0893_ (.A(_0198_),
    .B(_0203_),
    .Y(_0221_));
 sg13g2_and2_1 _0894_ (.A(net230),
    .B(net245),
    .X(_0222_));
 sg13g2_and3_1 _0895_ (.X(_0223_),
    .A(net256),
    .B(net255),
    .C(_0185_));
 sg13g2_nor4_1 _0896_ (.A(_0196_),
    .B(_0218_),
    .C(_0222_),
    .D(_0223_),
    .Y(_0224_));
 sg13g2_nor3_2 _0897_ (.A(_0220_),
    .B(_0221_),
    .C(_0224_),
    .Y(_0225_));
 sg13g2_and2_1 _0898_ (.A(net270),
    .B(\ctrl[6] ),
    .X(_0226_));
 sg13g2_nand2_1 _0899_ (.Y(_0227_),
    .A(net270),
    .B(\ctrl[6] ));
 sg13g2_a22oi_1 _0900_ (.Y(_0228_),
    .B1(net245),
    .B2(net253),
    .A2(_0188_),
    .A1(net232));
 sg13g2_nand2b_1 _0901_ (.Y(_0229_),
    .B(net229),
    .A_N(_0228_));
 sg13g2_nand4_1 _0902_ (.B(net255),
    .C(net248),
    .A(net256),
    .Y(_0230_),
    .D(_0214_));
 sg13g2_mux2_2 _0903_ (.A0(\bitmapIn[5] ),
    .A1(\bitmapIn[10] ),
    .S(net274),
    .X(_0231_));
 sg13g2_inv_1 _0904_ (.Y(_0232_),
    .A(_0231_));
 sg13g2_nor2_1 _0905_ (.A(net249),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_nand2_1 _0906_ (.Y(_0234_),
    .A(net253),
    .B(_0231_));
 sg13g2_a21oi_1 _0907_ (.A1(net253),
    .A2(_0231_),
    .Y(_0235_),
    .B1(net246));
 sg13g2_o21ai_1 _0908_ (.B1(_0230_),
    .Y(_0236_),
    .A1(net229),
    .A2(_0235_));
 sg13g2_o21ai_1 _0909_ (.B1(_0236_),
    .Y(_0237_),
    .A1(_0183_),
    .A2(net245));
 sg13g2_nand4_1 _0910_ (.B(_0134_),
    .C(net248),
    .A(_0132_),
    .Y(_0238_),
    .D(_0214_));
 sg13g2_a221oi_1 _0911_ (.B2(net253),
    .C1(_0196_),
    .B1(net245),
    .A1(net236),
    .Y(_0239_),
    .A2(_0188_));
 sg13g2_nor2_1 _0912_ (.A(_0185_),
    .B(_0203_),
    .Y(_0240_));
 sg13g2_a221oi_1 _0913_ (.B2(_0239_),
    .C1(_0240_),
    .B1(_0238_),
    .A1(_0229_),
    .Y(_0241_),
    .A2(_0237_));
 sg13g2_a221oi_1 _0914_ (.B2(_0241_),
    .C1(_0225_),
    .B1(net261),
    .A1(net268),
    .Y(_0242_),
    .A2(_0210_));
 sg13g2_nor2_1 _0915_ (.A(net275),
    .B(_0004_),
    .Y(_0243_));
 sg13g2_nand2b_1 _0916_ (.Y(_0244_),
    .B(net275),
    .A_N(_0005_));
 sg13g2_nor2b_1 _0917_ (.A(_0243_),
    .B_N(_0244_),
    .Y(_0245_));
 sg13g2_nand2b_1 _0918_ (.Y(_0246_),
    .B(_0244_),
    .A_N(_0243_));
 sg13g2_and2_1 _0919_ (.A(net277),
    .B(_0003_),
    .X(_0247_));
 sg13g2_a21oi_2 _0920_ (.B1(_0247_),
    .Y(_0248_),
    .A2(_0002_),
    .A1(_0086_));
 sg13g2_mux2_1 _0921_ (.A0(_0248_),
    .A1(_0246_),
    .S(net232),
    .X(_0249_));
 sg13g2_or2_1 _0922_ (.X(_0250_),
    .B(_0248_),
    .A(_0180_));
 sg13g2_a22oi_1 _0923_ (.Y(_0251_),
    .B1(_0250_),
    .B2(_0177_),
    .A2(_0249_),
    .A1(net229));
 sg13g2_mux2_1 _0924_ (.A0(_0246_),
    .A1(_0248_),
    .S(net254),
    .X(_0252_));
 sg13g2_nor2_1 _0925_ (.A(net232),
    .B(_0153_),
    .Y(_0253_));
 sg13g2_nand2_1 _0926_ (.Y(_0254_),
    .A(\bitmapIn[13] ),
    .B(net276));
 sg13g2_o21ai_1 _0927_ (.B1(_0254_),
    .Y(_0255_),
    .A1(net277),
    .A2(_0096_));
 sg13g2_and2_1 _0928_ (.A(net254),
    .B(_0255_),
    .X(_0256_));
 sg13g2_a221oi_1 _0929_ (.B2(net236),
    .C1(_0181_),
    .B1(_0256_),
    .A1(_0252_),
    .Y(_0257_),
    .A2(_0253_));
 sg13g2_nor2_1 _0930_ (.A(_0251_),
    .B(_0257_),
    .Y(_0258_));
 sg13g2_and2_1 _0931_ (.A(net248),
    .B(_0255_),
    .X(_0259_));
 sg13g2_nor4_1 _0932_ (.A(_0131_),
    .B(_0133_),
    .C(net250),
    .D(_0245_),
    .Y(_0260_));
 sg13g2_a221oi_1 _0933_ (.B2(net232),
    .C1(_0260_),
    .B1(_0255_),
    .A1(net236),
    .Y(_0261_),
    .A2(_0248_));
 sg13g2_o21ai_1 _0934_ (.B1(_0176_),
    .Y(_0262_),
    .A1(_0153_),
    .A2(_0261_));
 sg13g2_nand2_1 _0935_ (.Y(_0263_),
    .A(net232),
    .B(_0248_));
 sg13g2_nor2_1 _0936_ (.A(net275),
    .B(\bitmapIn[3] ),
    .Y(_0264_));
 sg13g2_nand2b_1 _0937_ (.Y(_0265_),
    .B(net274),
    .A_N(\bitmapIn[12] ));
 sg13g2_nor2b_2 _0938_ (.A(_0264_),
    .B_N(_0265_),
    .Y(_0266_));
 sg13g2_nand2b_1 _0939_ (.Y(_0267_),
    .B(_0265_),
    .A_N(_0264_));
 sg13g2_nor2_1 _0940_ (.A(net248),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_o21ai_1 _0941_ (.B1(net236),
    .Y(_0269_),
    .A1(_0259_),
    .A2(_0268_));
 sg13g2_nor2_1 _0942_ (.A(_0181_),
    .B(_0260_),
    .Y(_0270_));
 sg13g2_nand3_1 _0943_ (.B(_0269_),
    .C(_0270_),
    .A(_0263_),
    .Y(_0271_));
 sg13g2_nand2_1 _0944_ (.Y(_0272_),
    .A(_0182_),
    .B(_0245_));
 sg13g2_and3_2 _0945_ (.X(_0273_),
    .A(_0262_),
    .B(_0271_),
    .C(_0272_));
 sg13g2_a21oi_1 _0946_ (.A1(net270),
    .A2(_0273_),
    .Y(_0274_),
    .B1(_0258_));
 sg13g2_mux2_1 _0947_ (.A0(_0242_),
    .A1(_0274_),
    .S(net280),
    .X(_0275_));
 sg13g2_nand2b_1 _0948_ (.Y(_0276_),
    .B(net265),
    .A_N(_0275_));
 sg13g2_nor3_2 _0949_ (.A(_0155_),
    .B(_0161_),
    .C(_0167_),
    .Y(_0277_));
 sg13g2_inv_1 _0950_ (.Y(_0278_),
    .A(_0277_));
 sg13g2_nor2_1 _0951_ (.A(net275),
    .B(_0005_),
    .Y(_0279_));
 sg13g2_nand2b_1 _0952_ (.Y(_0280_),
    .B(net275),
    .A_N(_0004_));
 sg13g2_nor2b_2 _0953_ (.A(_0279_),
    .B_N(_0280_),
    .Y(_0281_));
 sg13g2_nand2b_2 _0954_ (.Y(_0282_),
    .B(_0280_),
    .A_N(_0279_));
 sg13g2_a21oi_1 _0955_ (.A1(_0132_),
    .A2(_0134_),
    .Y(_0283_),
    .B1(_0281_));
 sg13g2_or2_1 _0956_ (.X(_0284_),
    .B(net275),
    .A(\bitmapIn[12] ));
 sg13g2_o21ai_1 _0957_ (.B1(_0284_),
    .Y(_0285_),
    .A1(_0086_),
    .A2(\bitmapIn[3] ));
 sg13g2_nor4_2 _0958_ (.A(_0131_),
    .B(_0133_),
    .C(net253),
    .Y(_0286_),
    .D(_0285_));
 sg13g2_o21ai_1 _0959_ (.B1(_0154_),
    .Y(_0287_),
    .A1(_0283_),
    .A2(_0286_));
 sg13g2_mux2_2 _0960_ (.A0(\bitmapIn[13] ),
    .A1(\bitmapIn[2] ),
    .S(net276),
    .X(_0288_));
 sg13g2_inv_1 _0961_ (.Y(_0289_),
    .A(_0288_));
 sg13g2_nor2_1 _0962_ (.A(net249),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_and2_1 _0963_ (.A(net277),
    .B(_0002_),
    .X(_0291_));
 sg13g2_a21oi_2 _0964_ (.B1(_0291_),
    .Y(_0292_),
    .A2(_0003_),
    .A1(_0086_));
 sg13g2_a221oi_1 _0965_ (.B2(_0153_),
    .C1(_0181_),
    .B1(_0292_),
    .A1(_0137_),
    .Y(_0293_),
    .A2(_0290_));
 sg13g2_nor2_1 _0966_ (.A(_0183_),
    .B(_0288_),
    .Y(_0294_));
 sg13g2_a21oi_1 _0967_ (.A1(_0132_),
    .A2(_0134_),
    .Y(_0295_),
    .B1(_0285_));
 sg13g2_o21ai_1 _0968_ (.B1(_0154_),
    .Y(_0296_),
    .A1(_0290_),
    .A2(_0295_));
 sg13g2_and2_1 _0969_ (.A(net252),
    .B(_0205_),
    .X(_0297_));
 sg13g2_a221oi_1 _0970_ (.B2(net235),
    .C1(net247),
    .B1(_0297_),
    .A1(net231),
    .Y(_0298_),
    .A2(_0282_));
 sg13g2_a221oi_1 _0971_ (.B2(_0298_),
    .C1(_0294_),
    .B1(_0296_),
    .A1(_0287_),
    .Y(_0299_),
    .A2(_0293_));
 sg13g2_nand2_1 _0972_ (.Y(_0300_),
    .A(_0182_),
    .B(_0285_));
 sg13g2_and2_1 _0973_ (.A(net251),
    .B(_0198_),
    .X(_0301_));
 sg13g2_mux2_1 _0974_ (.A0(_0198_),
    .A1(_0205_),
    .S(net249),
    .X(_0302_));
 sg13g2_o21ai_1 _0975_ (.B1(_0300_),
    .Y(_0303_),
    .A1(net247),
    .A2(_0302_));
 sg13g2_nand2_1 _0976_ (.Y(_0304_),
    .A(net228),
    .B(_0303_));
 sg13g2_nor2_1 _0977_ (.A(net249),
    .B(_0285_),
    .Y(_0305_));
 sg13g2_a221oi_1 _0978_ (.B2(net235),
    .C1(_0305_),
    .B1(_0288_),
    .A1(net231),
    .Y(_0306_),
    .A2(_0205_));
 sg13g2_nor2_1 _0979_ (.A(_0203_),
    .B(_0282_),
    .Y(_0307_));
 sg13g2_nand2_1 _0980_ (.Y(_0308_),
    .A(net231),
    .B(_0288_));
 sg13g2_nor2_1 _0981_ (.A(net228),
    .B(_0305_),
    .Y(_0309_));
 sg13g2_a221oi_1 _0982_ (.B2(_0309_),
    .C1(_0307_),
    .B1(_0308_),
    .A1(_0195_),
    .Y(_0310_),
    .A2(_0306_));
 sg13g2_and2_1 _0983_ (.A(_0304_),
    .B(_0310_),
    .X(_0311_));
 sg13g2_o21ai_1 _0984_ (.B1(net229),
    .Y(_0312_),
    .A1(_0286_),
    .A2(_0297_));
 sg13g2_nor2_1 _0985_ (.A(_0183_),
    .B(_0205_),
    .Y(_0313_));
 sg13g2_a221oi_1 _0986_ (.B2(net234),
    .C1(net247),
    .B1(_0200_),
    .A1(net249),
    .Y(_0314_),
    .A2(_0199_));
 sg13g2_o21ai_1 _0987_ (.B1(_0312_),
    .Y(_0315_),
    .A1(_0313_),
    .A2(_0314_));
 sg13g2_nor4_1 _0988_ (.A(_0153_),
    .B(_0181_),
    .C(_0295_),
    .D(_0297_),
    .Y(_0316_));
 sg13g2_a22oi_1 _0989_ (.Y(_0317_),
    .B1(_0316_),
    .B2(_0207_),
    .A2(_0289_),
    .A1(_0202_));
 sg13g2_and2_1 _0990_ (.A(_0315_),
    .B(_0317_),
    .X(_0318_));
 sg13g2_nand2_1 _0991_ (.Y(_0319_),
    .A(_0315_),
    .B(_0317_));
 sg13g2_a22oi_1 _0992_ (.Y(_0320_),
    .B1(_0304_),
    .B2(_0310_),
    .A2(_0299_),
    .A1(net269));
 sg13g2_o21ai_1 _0993_ (.B1(_0320_),
    .Y(_0321_),
    .A1(_0227_),
    .A2(_0319_));
 sg13g2_nand2_1 _0994_ (.Y(_0322_),
    .A(\bitmapIn[11] ),
    .B(net276));
 sg13g2_o21ai_1 _0995_ (.B1(_0322_),
    .Y(_0323_),
    .A1(net276),
    .A2(_0094_));
 sg13g2_and3_1 _0996_ (.X(_0324_),
    .A(_0135_),
    .B(net255),
    .C(_0323_));
 sg13g2_a221oi_1 _0997_ (.B2(net230),
    .C1(net228),
    .B1(_0323_),
    .A1(net251),
    .Y(_0325_),
    .A2(_0266_));
 sg13g2_a221oi_1 _0998_ (.B2(net236),
    .C1(_0268_),
    .B1(_0323_),
    .A1(net233),
    .Y(_0326_),
    .A2(_0255_));
 sg13g2_nand2_1 _0999_ (.Y(_0327_),
    .A(_0182_),
    .B(_0267_));
 sg13g2_o21ai_1 _1000_ (.B1(_0176_),
    .Y(_0328_),
    .A1(net248),
    .A2(_0245_));
 sg13g2_o21ai_1 _1001_ (.B1(_0327_),
    .Y(_0329_),
    .A1(_0259_),
    .A2(_0328_));
 sg13g2_a21oi_1 _1002_ (.A1(_0202_),
    .A2(_0232_),
    .Y(_0330_),
    .B1(_0325_));
 sg13g2_a22oi_1 _1003_ (.Y(_0331_),
    .B1(_0329_),
    .B2(net228),
    .A2(_0326_),
    .A1(_0195_));
 sg13g2_and2_1 _1004_ (.A(_0330_),
    .B(_0331_),
    .X(_0332_));
 sg13g2_nand3_1 _1005_ (.B(_0330_),
    .C(_0331_),
    .A(net261),
    .Y(_0333_));
 sg13g2_nand2_1 _1006_ (.Y(_0334_),
    .A(net251),
    .B(_0323_));
 sg13g2_mux2_1 _1007_ (.A0(_0231_),
    .A1(_0323_),
    .S(net251),
    .X(_0335_));
 sg13g2_nand2_1 _1008_ (.Y(_0336_),
    .A(net229),
    .B(_0335_));
 sg13g2_nor2_1 _1009_ (.A(_0183_),
    .B(_0323_),
    .Y(_0337_));
 sg13g2_a21oi_1 _1010_ (.A1(_0132_),
    .A2(_0134_),
    .Y(_0338_),
    .B1(_0267_));
 sg13g2_a221oi_1 _1011_ (.B2(net248),
    .C1(net246),
    .B1(_0338_),
    .A1(net237),
    .Y(_0339_),
    .A2(_0256_));
 sg13g2_o21ai_1 _1012_ (.B1(_0336_),
    .Y(_0340_),
    .A1(_0337_),
    .A2(_0339_));
 sg13g2_nor4_1 _1013_ (.A(_0131_),
    .B(_0133_),
    .C(net253),
    .D(_0267_),
    .Y(_0341_));
 sg13g2_nand2_1 _1014_ (.Y(_0342_),
    .A(net231),
    .B(_0266_));
 sg13g2_nand3_1 _1015_ (.B(net255),
    .C(_0231_),
    .A(net256),
    .Y(_0343_));
 sg13g2_and4_1 _1016_ (.A(_0154_),
    .B(_0180_),
    .C(_0334_),
    .D(_0343_),
    .X(_0344_));
 sg13g2_a22oi_1 _1017_ (.Y(_0345_),
    .B1(_0342_),
    .B2(_0344_),
    .A2(_0215_),
    .A1(_0202_));
 sg13g2_and2_1 _1018_ (.A(_0340_),
    .B(_0345_),
    .X(_0346_));
 sg13g2_nand2_1 _1019_ (.Y(_0347_),
    .A(_0340_),
    .B(_0345_));
 sg13g2_a21o_1 _1020_ (.A2(_0238_),
    .A1(_0234_),
    .B1(_0179_),
    .X(_0348_));
 sg13g2_nor2_1 _1021_ (.A(_0183_),
    .B(_0231_),
    .Y(_0349_));
 sg13g2_a221oi_1 _1022_ (.B2(net248),
    .C1(net246),
    .B1(_0324_),
    .A1(net237),
    .Y(_0350_),
    .A2(_0268_));
 sg13g2_o21ai_1 _1023_ (.B1(_0348_),
    .Y(_0351_),
    .A1(_0349_),
    .A2(_0350_));
 sg13g2_a221oi_1 _1024_ (.B2(net230),
    .C1(_0233_),
    .B1(_0323_),
    .A1(net234),
    .Y(_0352_),
    .A2(_0214_));
 sg13g2_a22oi_1 _1025_ (.Y(_0353_),
    .B1(_0352_),
    .B2(_0195_),
    .A2(_0202_),
    .A1(_0191_));
 sg13g2_and2_1 _1026_ (.A(_0351_),
    .B(_0353_),
    .X(_0354_));
 sg13g2_nand3_1 _1027_ (.B(_0351_),
    .C(_0353_),
    .A(net268),
    .Y(_0355_));
 sg13g2_nand3_1 _1028_ (.B(_0347_),
    .C(_0355_),
    .A(_0333_),
    .Y(_0356_));
 sg13g2_mux2_1 _1029_ (.A0(_0321_),
    .A1(_0356_),
    .S(net281),
    .X(_0357_));
 sg13g2_a21oi_1 _1030_ (.A1(net279),
    .A2(_0357_),
    .Y(_0358_),
    .B1(_0278_));
 sg13g2_a21oi_1 _1031_ (.A1(_0276_),
    .A2(_0358_),
    .Y(_0359_),
    .B1(_0175_));
 sg13g2_xnor2_1 _1032_ (.Y(_0360_),
    .A(_0119_),
    .B(_0359_));
 sg13g2_and2_2 _1033_ (.A(net1),
    .B(net2),
    .X(_0361_));
 sg13g2_nand2_2 _1034_ (.Y(_0362_),
    .A(net1),
    .B(net2));
 sg13g2_a21oi_2 _1035_ (.B1(_0122_),
    .Y(_0363_),
    .A2(_0172_),
    .A1(_0170_));
 sg13g2_o21ai_1 _1036_ (.B1(_0121_),
    .Y(_0364_),
    .A1(_0169_),
    .A2(_0173_));
 sg13g2_nand3_1 _1037_ (.B(_0304_),
    .C(_0310_),
    .A(net269),
    .Y(_0365_));
 sg13g2_nand2_1 _1038_ (.Y(_0366_),
    .A(net229),
    .B(_0302_));
 sg13g2_nor2_1 _1039_ (.A(_0183_),
    .B(_0198_),
    .Y(_0367_));
 sg13g2_a221oi_1 _1040_ (.B2(net249),
    .C1(net247),
    .B1(_0223_),
    .A1(net234),
    .Y(_0368_),
    .A2(_0218_));
 sg13g2_o21ai_1 _1041_ (.B1(_0366_),
    .Y(_0369_),
    .A1(_0367_),
    .A2(_0368_));
 sg13g2_a221oi_1 _1042_ (.B2(net234),
    .C1(_0301_),
    .B1(_0205_),
    .A1(net230),
    .Y(_0370_),
    .A2(_0185_));
 sg13g2_a22oi_1 _1043_ (.Y(_0371_),
    .B1(_0370_),
    .B2(_0195_),
    .A2(_0285_),
    .A1(_0202_));
 sg13g2_and2_1 _1044_ (.A(_0369_),
    .B(_0371_),
    .X(_0372_));
 sg13g2_nand3_1 _1045_ (.B(_0369_),
    .C(_0371_),
    .A(net261),
    .Y(_0373_));
 sg13g2_nand3_1 _1046_ (.B(_0365_),
    .C(_0373_),
    .A(_0319_),
    .Y(_0374_));
 sg13g2_o21ai_1 _1047_ (.B1(net229),
    .Y(_0375_),
    .A1(_0256_),
    .A2(_0341_));
 sg13g2_a21oi_1 _1048_ (.A1(_0132_),
    .A2(_0134_),
    .Y(_0376_),
    .B1(net246));
 sg13g2_a221oi_1 _1049_ (.B2(_0252_),
    .C1(_0180_),
    .B1(_0376_),
    .A1(net246),
    .Y(_0377_),
    .A2(_0255_));
 sg13g2_nor2_1 _1050_ (.A(_0203_),
    .B(_0323_),
    .Y(_0378_));
 sg13g2_a221oi_1 _1051_ (.B2(net236),
    .C1(_0256_),
    .B1(_0266_),
    .A1(net232),
    .Y(_0379_),
    .A2(_0246_));
 sg13g2_a221oi_1 _1052_ (.B2(_0195_),
    .C1(_0378_),
    .B1(_0379_),
    .A1(_0375_),
    .Y(_0380_),
    .A2(_0377_));
 sg13g2_nand2_1 _1053_ (.Y(_0381_),
    .A(net261),
    .B(_0380_));
 sg13g2_nand3_1 _1054_ (.B(_0340_),
    .C(_0345_),
    .A(net268),
    .Y(_0382_));
 sg13g2_nand3b_1 _1055_ (.B(_0381_),
    .C(_0382_),
    .Y(_0383_),
    .A_N(_0332_));
 sg13g2_mux2_1 _1056_ (.A0(_0374_),
    .A1(_0383_),
    .S(net280),
    .X(_0384_));
 sg13g2_a21oi_1 _1057_ (.A1(net279),
    .A2(_0384_),
    .Y(_0385_),
    .B1(_0278_));
 sg13g2_mux2_1 _1058_ (.A0(_0292_),
    .A1(_0282_),
    .S(net233),
    .X(_0386_));
 sg13g2_nand3_1 _1059_ (.B(_0180_),
    .C(_0386_),
    .A(_0137_),
    .Y(_0387_));
 sg13g2_a21o_1 _1060_ (.A2(_0292_),
    .A1(net252),
    .B1(_0283_),
    .X(_0388_));
 sg13g2_nand3_1 _1061_ (.B(_0176_),
    .C(_0388_),
    .A(_0154_),
    .Y(_0389_));
 sg13g2_nand2_1 _1062_ (.Y(_0390_),
    .A(_0182_),
    .B(_0292_));
 sg13g2_nand2_1 _1063_ (.Y(_0391_),
    .A(_0290_),
    .B(_0376_));
 sg13g2_nand4_1 _1064_ (.B(_0389_),
    .C(_0390_),
    .A(_0387_),
    .Y(_0392_),
    .D(_0391_));
 sg13g2_nor4_2 _1065_ (.A(_0131_),
    .B(_0133_),
    .C(net250),
    .Y(_0393_),
    .D(_0281_));
 sg13g2_a21oi_1 _1066_ (.A1(net235),
    .A2(_0292_),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_a21oi_1 _1067_ (.A1(_0308_),
    .A2(_0394_),
    .Y(_0395_),
    .B1(_0196_));
 sg13g2_a221oi_1 _1068_ (.B2(net233),
    .C1(_0393_),
    .B1(_0292_),
    .A1(net235),
    .Y(_0396_),
    .A2(_0288_));
 sg13g2_a21oi_1 _1069_ (.A1(net234),
    .A2(_0305_),
    .Y(_0397_),
    .B1(net247));
 sg13g2_o21ai_1 _1070_ (.B1(_0397_),
    .Y(_0398_),
    .A1(_0153_),
    .A2(_0396_));
 sg13g2_o21ai_1 _1071_ (.B1(net247),
    .Y(_0399_),
    .A1(_0180_),
    .A2(_0281_));
 sg13g2_a21o_1 _1072_ (.A2(_0399_),
    .A1(_0398_),
    .B1(_0395_),
    .X(_0400_));
 sg13g2_a21oi_1 _1073_ (.A1(net262),
    .A2(_0400_),
    .Y(_0401_),
    .B1(_0392_));
 sg13g2_nand2_1 _1074_ (.Y(_0402_),
    .A(net281),
    .B(_0401_));
 sg13g2_a22oi_1 _1075_ (.Y(_0403_),
    .B1(_0214_),
    .B2(net251),
    .A2(net245),
    .A1(net234));
 sg13g2_a221oi_1 _1076_ (.B2(net230),
    .C1(_0181_),
    .B1(_0231_),
    .A1(net234),
    .Y(_0404_),
    .A2(_0218_));
 sg13g2_o21ai_1 _1077_ (.B1(_0404_),
    .Y(_0405_),
    .A1(_0153_),
    .A2(_0403_));
 sg13g2_nand2b_1 _1078_ (.Y(_0406_),
    .B(_0182_),
    .A_N(_0214_));
 sg13g2_o21ai_1 _1079_ (.B1(_0406_),
    .Y(_0407_),
    .A1(net247),
    .A2(_0335_));
 sg13g2_a221oi_1 _1080_ (.B2(net251),
    .C1(net228),
    .B1(_0214_),
    .A1(net230),
    .Y(_0408_),
    .A2(net245));
 sg13g2_a21oi_1 _1081_ (.A1(net228),
    .A2(_0407_),
    .Y(_0409_),
    .B1(_0408_));
 sg13g2_and2_1 _1082_ (.A(_0405_),
    .B(_0409_),
    .X(_0410_));
 sg13g2_a221oi_1 _1083_ (.B2(_0410_),
    .C1(_0241_),
    .B1(net261),
    .A1(net268),
    .Y(_0411_),
    .A2(_0225_));
 sg13g2_a21oi_1 _1084_ (.A1(net263),
    .A2(_0411_),
    .Y(_0412_),
    .B1(net278));
 sg13g2_nand2_1 _1085_ (.Y(_0413_),
    .A(_0402_),
    .B(_0412_));
 sg13g2_a21oi_1 _1086_ (.A1(_0385_),
    .A2(_0413_),
    .Y(_0414_),
    .B1(_0364_));
 sg13g2_xnor2_1 _1087_ (.Y(_0415_),
    .A(net227),
    .B(_0414_));
 sg13g2_nand2_1 _1088_ (.Y(_0416_),
    .A(\s.inv.xPostMirror ),
    .B(_0415_));
 sg13g2_a21oi_1 _1089_ (.A1(_0085_),
    .A2(_0360_),
    .Y(_0417_),
    .B1(_0362_));
 sg13g2_o21ai_1 _1090_ (.B1(_0277_),
    .Y(_0418_),
    .A1(net265),
    .A2(_0275_));
 sg13g2_a21o_1 _1091_ (.A2(_0274_),
    .A1(net263),
    .B1(net278),
    .X(_0419_));
 sg13g2_a21oi_1 _1092_ (.A1(net281),
    .A2(_0242_),
    .Y(_0420_),
    .B1(_0419_));
 sg13g2_o21ai_1 _1093_ (.B1(_0174_),
    .Y(_0421_),
    .A1(_0418_),
    .A2(_0420_));
 sg13g2_xor2_1 _1094_ (.B(_0421_),
    .A(net227),
    .X(_0422_));
 sg13g2_nor2b_1 _1095_ (.A(net1),
    .B_N(net2),
    .Y(_0423_));
 sg13g2_nand2b_2 _1096_ (.Y(_0424_),
    .B(net2),
    .A_N(net1));
 sg13g2_mux2_1 _1097_ (.A0(_0401_),
    .A1(_0411_),
    .S(net281),
    .X(_0425_));
 sg13g2_a21oi_1 _1098_ (.A1(_0277_),
    .A2(_0425_),
    .Y(_0426_),
    .B1(_0364_));
 sg13g2_xor2_1 _1099_ (.B(_0426_),
    .A(net227),
    .X(_0427_));
 sg13g2_nor2_1 _1100_ (.A(net267),
    .B(_0427_),
    .Y(_0428_));
 sg13g2_a21oi_1 _1101_ (.A1(net267),
    .A2(_0422_),
    .Y(_0429_),
    .B1(_0428_));
 sg13g2_nor2_1 _1102_ (.A(net1),
    .B(net2),
    .Y(_0430_));
 sg13g2_xor2_1 _1103_ (.B(_0128_),
    .A(_0000_),
    .X(_0431_));
 sg13g2_nor2b_1 _1104_ (.A(net2),
    .B_N(net1),
    .Y(_0432_));
 sg13g2_a22oi_1 _1105_ (.Y(_0433_),
    .B1(net283),
    .B2(\ctrl[0] ),
    .A2(_0431_),
    .A1(net286));
 sg13g2_nand2_1 _1106_ (.Y(_0434_),
    .A(net288),
    .B(_0433_));
 sg13g2_a221oi_1 _1107_ (.B2(_0429_),
    .C1(_0434_),
    .B1(net287),
    .A1(_0416_),
    .Y(_0435_),
    .A2(_0417_));
 sg13g2_nor2_1 _1108_ (.A(_0073_),
    .B(_0424_),
    .Y(_0436_));
 sg13g2_a21oi_1 _1109_ (.A1(\s.sty.xoffset ),
    .A2(net285),
    .Y(_0437_),
    .B1(net288));
 sg13g2_a221oi_1 _1110_ (.B2(\s.bold ),
    .C1(_0436_),
    .B1(net282),
    .A1(\s.dottedOverline ),
    .Y(_0438_),
    .A2(_0361_));
 sg13g2_a21oi_2 _1111_ (.B1(_0435_),
    .Y(uio_out[0]),
    .A2(_0438_),
    .A1(_0437_));
 sg13g2_a221oi_1 _1112_ (.B2(net269),
    .C1(_0210_),
    .B1(_0372_),
    .A1(_0225_),
    .Y(_0439_),
    .A2(net262));
 sg13g2_and2_1 _1113_ (.A(net268),
    .B(_0380_),
    .X(_0440_));
 sg13g2_nor3_1 _1114_ (.A(_0227_),
    .B(_0251_),
    .C(_0257_),
    .Y(_0441_));
 sg13g2_nor4_1 _1115_ (.A(net263),
    .B(_0273_),
    .C(_0440_),
    .D(_0441_),
    .Y(_0442_));
 sg13g2_a21oi_1 _1116_ (.A1(net263),
    .A2(_0439_),
    .Y(_0443_),
    .B1(_0442_));
 sg13g2_nand2_1 _1117_ (.Y(_0444_),
    .A(net264),
    .B(_0443_));
 sg13g2_a21oi_1 _1118_ (.A1(_0358_),
    .A2(_0444_),
    .Y(_0445_),
    .B1(_0364_));
 sg13g2_xnor2_1 _1119_ (.Y(_0446_),
    .A(net226),
    .B(_0445_));
 sg13g2_nor4_1 _1120_ (.A(net281),
    .B(_0273_),
    .C(_0440_),
    .D(_0441_),
    .Y(_0447_));
 sg13g2_a21oi_1 _1121_ (.A1(net281),
    .A2(_0439_),
    .Y(_0448_),
    .B1(_0447_));
 sg13g2_and2_1 _1122_ (.A(net264),
    .B(_0448_),
    .X(_0449_));
 sg13g2_o21ai_1 _1123_ (.B1(_0363_),
    .Y(_0450_),
    .A1(_0418_),
    .A2(_0449_));
 sg13g2_xor2_1 _1124_ (.B(_0450_),
    .A(net227),
    .X(_0451_));
 sg13g2_xor2_1 _1125_ (.B(_0126_),
    .A(_0000_),
    .X(_0452_));
 sg13g2_a21o_1 _1126_ (.A2(net284),
    .A1(\ctrl[1] ),
    .B1(net3),
    .X(_0453_));
 sg13g2_a221oi_1 _1127_ (.B2(net261),
    .C1(_0410_),
    .B1(_0354_),
    .A1(net268),
    .Y(_0454_),
    .A2(_0241_));
 sg13g2_nand2_1 _1128_ (.Y(_0455_),
    .A(_0090_),
    .B(_0454_));
 sg13g2_a221oi_1 _1129_ (.B2(net270),
    .C1(_0400_),
    .B1(_0392_),
    .A1(net262),
    .Y(_0456_),
    .A2(_0299_));
 sg13g2_a21oi_1 _1130_ (.A1(net280),
    .A2(_0456_),
    .Y(_0457_),
    .B1(net278));
 sg13g2_nand2_1 _1131_ (.Y(_0458_),
    .A(_0455_),
    .B(_0457_));
 sg13g2_a21oi_1 _1132_ (.A1(_0385_),
    .A2(_0458_),
    .Y(_0459_),
    .B1(_0175_));
 sg13g2_xnor2_1 _1133_ (.Y(_0460_),
    .A(net226),
    .B(_0459_));
 sg13g2_mux2_1 _1134_ (.A0(_0454_),
    .A1(_0456_),
    .S(_0090_),
    .X(_0461_));
 sg13g2_mux2_1 _1135_ (.A0(_0425_),
    .A1(_0461_),
    .S(net265),
    .X(_0462_));
 sg13g2_a21oi_1 _1136_ (.A1(_0277_),
    .A2(_0462_),
    .Y(_0463_),
    .B1(_0175_));
 sg13g2_xnor2_1 _1137_ (.Y(_0464_),
    .A(net227),
    .B(_0463_));
 sg13g2_nand2_1 _1138_ (.Y(_0465_),
    .A(net267),
    .B(_0451_));
 sg13g2_a21oi_1 _1139_ (.A1(\s.inv.xPostMirror ),
    .A2(_0464_),
    .Y(_0466_),
    .B1(_0424_));
 sg13g2_nand2_1 _1140_ (.Y(_0467_),
    .A(net266),
    .B(_0446_));
 sg13g2_a21oi_1 _1141_ (.A1(net272),
    .A2(_0460_),
    .Y(_0468_),
    .B1(_0362_));
 sg13g2_nand2_1 _1142_ (.Y(_0469_),
    .A(_0467_),
    .B(_0468_));
 sg13g2_a221oi_1 _1143_ (.B2(_0466_),
    .C1(_0453_),
    .B1(_0465_),
    .A1(net285),
    .Y(_0470_),
    .A2(_0452_));
 sg13g2_a21oi_1 _1144_ (.A1(\s.faint ),
    .A2(net282),
    .Y(_0471_),
    .B1(net288));
 sg13g2_a22oi_1 _1145_ (.Y(_0472_),
    .B1(net285),
    .B2(net278),
    .A2(net287),
    .A1(\s.doubleUnderline ));
 sg13g2_a22oi_1 _1146_ (.Y(uio_out[1]),
    .B1(_0471_),
    .B2(_0472_),
    .A2(_0470_),
    .A1(_0469_));
 sg13g2_a21oi_1 _1147_ (.A1(net279),
    .A2(_0443_),
    .Y(_0473_),
    .B1(_0278_));
 sg13g2_a221oi_1 _1148_ (.B2(net269),
    .C1(_0372_),
    .B1(_0318_),
    .A1(_0210_),
    .Y(_0474_),
    .A2(net261));
 sg13g2_nand2_1 _1149_ (.Y(_0475_),
    .A(net280),
    .B(_0474_));
 sg13g2_a221oi_1 _1150_ (.B2(net268),
    .C1(_0380_),
    .B1(_0332_),
    .A1(net262),
    .Y(_0476_),
    .A2(_0273_));
 sg13g2_a21oi_1 _1151_ (.A1(net263),
    .A2(_0476_),
    .Y(_0477_),
    .B1(net278));
 sg13g2_nand2_1 _1152_ (.Y(_0478_),
    .A(_0475_),
    .B(_0477_));
 sg13g2_a21oi_1 _1153_ (.A1(_0473_),
    .A2(_0478_),
    .Y(_0479_),
    .B1(_0175_));
 sg13g2_xnor2_1 _1154_ (.Y(_0480_),
    .A(net226),
    .B(_0479_));
 sg13g2_nand2_1 _1155_ (.Y(_0481_),
    .A(net266),
    .B(_0480_));
 sg13g2_a221oi_1 _1156_ (.B2(net270),
    .C1(_0299_),
    .B1(_0400_),
    .A1(net262),
    .Y(_0482_),
    .A2(_0311_));
 sg13g2_a221oi_1 _1157_ (.B2(net268),
    .C1(_0354_),
    .B1(_0410_),
    .A1(net261),
    .Y(_0483_),
    .A2(_0346_));
 sg13g2_mux2_1 _1158_ (.A0(_0482_),
    .A1(_0483_),
    .S(net281),
    .X(_0484_));
 sg13g2_nor2_1 _1159_ (.A(net279),
    .B(_0484_),
    .Y(_0485_));
 sg13g2_o21ai_1 _1160_ (.B1(_0277_),
    .Y(_0486_),
    .A1(net265),
    .A2(_0461_));
 sg13g2_o21ai_1 _1161_ (.B1(_0363_),
    .Y(_0487_),
    .A1(_0485_),
    .A2(_0486_));
 sg13g2_xor2_1 _1162_ (.B(_0487_),
    .A(net227),
    .X(_0488_));
 sg13g2_a21oi_1 _1163_ (.A1(net271),
    .A2(_0488_),
    .Y(_0489_),
    .B1(_0424_));
 sg13g2_o21ai_1 _1164_ (.B1(_0277_),
    .Y(_0490_),
    .A1(net264),
    .A2(_0484_));
 sg13g2_mux2_1 _1165_ (.A0(_0474_),
    .A1(_0476_),
    .S(net280),
    .X(_0491_));
 sg13g2_nor2_1 _1166_ (.A(net278),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_o21ai_1 _1167_ (.B1(_0174_),
    .Y(_0493_),
    .A1(_0490_),
    .A2(_0492_));
 sg13g2_xor2_1 _1168_ (.B(_0493_),
    .A(net226),
    .X(_0494_));
 sg13g2_nand2_1 _1169_ (.Y(_0495_),
    .A(net266),
    .B(_0494_));
 sg13g2_o21ai_1 _1170_ (.B1(_0277_),
    .Y(_0496_),
    .A1(net264),
    .A2(_0491_));
 sg13g2_a21o_1 _1171_ (.A2(_0482_),
    .A1(net280),
    .B1(net278),
    .X(_0497_));
 sg13g2_a21oi_1 _1172_ (.A1(net263),
    .A2(_0483_),
    .Y(_0498_),
    .B1(_0497_));
 sg13g2_o21ai_1 _1173_ (.B1(_0363_),
    .Y(_0499_),
    .A1(_0496_),
    .A2(_0498_));
 sg13g2_xor2_1 _1174_ (.B(_0499_),
    .A(net226),
    .X(_0500_));
 sg13g2_a21oi_1 _1175_ (.A1(net271),
    .A2(_0500_),
    .Y(_0501_),
    .B1(_0362_));
 sg13g2_xnor2_1 _1176_ (.Y(_0502_),
    .A(_0000_),
    .B(net250));
 sg13g2_a22oi_1 _1177_ (.Y(_0503_),
    .B1(_0502_),
    .B2(net286),
    .A2(net283),
    .A1(\ctrl[2] ));
 sg13g2_nand2_1 _1178_ (.Y(_0504_),
    .A(net289),
    .B(_0503_));
 sg13g2_a221oi_1 _1179_ (.B2(_0501_),
    .C1(_0504_),
    .B1(_0495_),
    .A1(_0481_),
    .Y(_0505_),
    .A2(_0489_));
 sg13g2_a22oi_1 _1180_ (.Y(_0506_),
    .B1(net284),
    .B2(\s.italic ),
    .A2(net286),
    .A1(\s.lg.yoffset ));
 sg13g2_a21oi_1 _1181_ (.A1(\s.dottedUnderline ),
    .A2(net287),
    .Y(_0507_),
    .B1(net289));
 sg13g2_a21oi_2 _1182_ (.B1(_0505_),
    .Y(uio_out[2]),
    .A2(_0507_),
    .A1(_0506_));
 sg13g2_mux2_1 _1183_ (.A0(_0374_),
    .A1(_0383_),
    .S(net263),
    .X(_0508_));
 sg13g2_nand2_1 _1184_ (.Y(_0509_),
    .A(net264),
    .B(_0508_));
 sg13g2_a21oi_1 _1185_ (.A1(_0473_),
    .A2(_0509_),
    .Y(_0510_),
    .B1(_0364_));
 sg13g2_xnor2_1 _1186_ (.Y(_0511_),
    .A(net226),
    .B(_0510_));
 sg13g2_nand2_1 _1187_ (.Y(_0512_),
    .A(net266),
    .B(_0511_));
 sg13g2_and2_1 _1188_ (.A(net265),
    .B(_0357_),
    .X(_0513_));
 sg13g2_o21ai_1 _1189_ (.B1(_0174_),
    .Y(_0514_),
    .A1(_0486_),
    .A2(_0513_));
 sg13g2_xor2_1 _1190_ (.B(_0514_),
    .A(net227),
    .X(_0515_));
 sg13g2_a21oi_1 _1191_ (.A1(\s.inv.xPostMirror ),
    .A2(_0515_),
    .Y(_0516_),
    .B1(_0424_));
 sg13g2_and2_1 _1192_ (.A(net264),
    .B(_0384_),
    .X(_0517_));
 sg13g2_o21ai_1 _1193_ (.B1(_0363_),
    .Y(_0518_),
    .A1(_0490_),
    .A2(_0517_));
 sg13g2_xor2_1 _1194_ (.B(_0518_),
    .A(net226),
    .X(_0519_));
 sg13g2_nand2_1 _1195_ (.Y(_0520_),
    .A(net266),
    .B(_0519_));
 sg13g2_nor2_1 _1196_ (.A(_0090_),
    .B(_0321_),
    .Y(_0521_));
 sg13g2_o21ai_1 _1197_ (.B1(net264),
    .Y(_0522_),
    .A1(net280),
    .A2(_0356_));
 sg13g2_nor2_1 _1198_ (.A(_0521_),
    .B(_0522_),
    .Y(_0523_));
 sg13g2_o21ai_1 _1199_ (.B1(_0174_),
    .Y(_0524_),
    .A1(_0496_),
    .A2(_0523_));
 sg13g2_xor2_1 _1200_ (.B(_0524_),
    .A(net226),
    .X(_0525_));
 sg13g2_a21oi_1 _1201_ (.A1(net271),
    .A2(_0525_),
    .Y(_0526_),
    .B1(_0362_));
 sg13g2_xnor2_1 _1202_ (.Y(_0527_),
    .A(_0000_),
    .B(_0137_));
 sg13g2_a22oi_1 _1203_ (.Y(_0528_),
    .B1(_0527_),
    .B2(net286),
    .A2(net283),
    .A1(\ctrl[3] ));
 sg13g2_nand2_1 _1204_ (.Y(_0529_),
    .A(net289),
    .B(_0528_));
 sg13g2_a221oi_1 _1205_ (.B2(_0526_),
    .C1(_0529_),
    .B1(_0520_),
    .A1(_0512_),
    .Y(_0530_),
    .A2(_0516_));
 sg13g2_a21oi_1 _1206_ (.A1(\s.lg.yscale ),
    .A2(net285),
    .Y(_0531_),
    .B1(net289));
 sg13g2_a22oi_1 _1207_ (.Y(_0532_),
    .B1(net284),
    .B2(\s.reverseItalic ),
    .A2(_0423_),
    .A1(\s.lg.strikethru ));
 sg13g2_a21oi_2 _1208_ (.B1(_0530_),
    .Y(uio_out[3]),
    .A2(_0532_),
    .A1(_0531_));
 sg13g2_nand2_1 _1209_ (.Y(_0533_),
    .A(net271),
    .B(_0511_));
 sg13g2_a21oi_1 _1210_ (.A1(_0085_),
    .A2(_0515_),
    .Y(_0534_),
    .B1(_0362_));
 sg13g2_nand2_1 _1211_ (.Y(_0535_),
    .A(net271),
    .B(_0519_));
 sg13g2_a21oi_1 _1212_ (.A1(net266),
    .A2(_0525_),
    .Y(_0536_),
    .B1(_0424_));
 sg13g2_nand2_1 _1213_ (.Y(_0537_),
    .A(_0535_),
    .B(_0536_));
 sg13g2_a221oi_1 _1214_ (.B2(_0534_),
    .C1(net3),
    .B1(_0533_),
    .A1(\ctrl[4] ),
    .Y(_0538_),
    .A2(net282));
 sg13g2_a21oi_1 _1215_ (.A1(\s.blink ),
    .A2(net282),
    .Y(_0539_),
    .B1(net288));
 sg13g2_a22oi_1 _1216_ (.Y(_0540_),
    .B1(net286),
    .B2(net277),
    .A2(_0423_),
    .A1(\s.doubleStrikethru ));
 sg13g2_a22oi_1 _1217_ (.Y(uio_out[4]),
    .B1(_0539_),
    .B2(_0540_),
    .A2(_0538_),
    .A1(_0537_));
 sg13g2_nand2_1 _1218_ (.Y(_0541_),
    .A(net271),
    .B(_0480_));
 sg13g2_a21oi_1 _1219_ (.A1(net267),
    .A2(_0488_),
    .Y(_0542_),
    .B1(_0362_));
 sg13g2_nand2_1 _1220_ (.Y(_0543_),
    .A(net271),
    .B(_0494_));
 sg13g2_a21oi_1 _1221_ (.A1(net266),
    .A2(_0500_),
    .Y(_0544_),
    .B1(_0424_));
 sg13g2_nand2_1 _1222_ (.Y(_0545_),
    .A(_0543_),
    .B(_0544_));
 sg13g2_a221oi_1 _1223_ (.B2(_0542_),
    .C1(net3),
    .B1(_0541_),
    .A1(\ctrl[5] ),
    .Y(_0546_),
    .A2(net282));
 sg13g2_a21oi_1 _1224_ (.A1(net272),
    .A2(net285),
    .Y(_0547_),
    .B1(net288));
 sg13g2_a22oi_1 _1225_ (.Y(_0548_),
    .B1(net283),
    .B2(\s.alternate ),
    .A2(net287),
    .A1(\s.dottedStrikethru ));
 sg13g2_a22oi_1 _1226_ (.Y(uio_out[5]),
    .B1(_0547_),
    .B2(_0548_),
    .A2(_0546_),
    .A1(_0545_));
 sg13g2_nand2_1 _1227_ (.Y(_0549_),
    .A(net267),
    .B(_0464_));
 sg13g2_a21oi_1 _1228_ (.A1(net272),
    .A2(_0451_),
    .Y(_0550_),
    .B1(_0362_));
 sg13g2_nand2_1 _1229_ (.Y(_0551_),
    .A(net271),
    .B(_0446_));
 sg13g2_a21oi_1 _1230_ (.A1(net266),
    .A2(_0460_),
    .Y(_0552_),
    .B1(_0424_));
 sg13g2_nand2_1 _1231_ (.Y(_0553_),
    .A(_0551_),
    .B(_0552_));
 sg13g2_a221oi_1 _1232_ (.B2(_0550_),
    .C1(net3),
    .B1(_0549_),
    .A1(\ctrl[6] ),
    .Y(_0554_),
    .A2(net282));
 sg13g2_a21oi_1 _1233_ (.A1(\s.lg.overline ),
    .A2(net287),
    .Y(_0555_),
    .B1(net288));
 sg13g2_a22oi_1 _1234_ (.Y(_0556_),
    .B1(net283),
    .B2(\s.inverse ),
    .A2(net286),
    .A1(\s.lg.yPreMirror ));
 sg13g2_a22oi_1 _1235_ (.Y(uio_out[6]),
    .B1(_0555_),
    .B2(_0556_),
    .A2(_0554_),
    .A1(_0553_));
 sg13g2_nand2_1 _1236_ (.Y(_0557_),
    .A(net267),
    .B(_0415_));
 sg13g2_a21oi_1 _1237_ (.A1(net272),
    .A2(_0360_),
    .Y(_0558_),
    .B1(_0424_));
 sg13g2_nand2_1 _1238_ (.Y(_0559_),
    .A(_0557_),
    .B(_0558_));
 sg13g2_o21ai_1 _1239_ (.B1(_0361_),
    .Y(_0560_),
    .A1(net272),
    .A2(_0427_));
 sg13g2_a21oi_1 _1240_ (.A1(net272),
    .A2(_0422_),
    .Y(_0561_),
    .B1(_0560_));
 sg13g2_a21oi_1 _1241_ (.A1(\ctrl[7] ),
    .A2(net283),
    .Y(_0562_),
    .B1(net3));
 sg13g2_nor2b_1 _1242_ (.A(_0561_),
    .B_N(_0562_),
    .Y(_0563_));
 sg13g2_a22oi_1 _1243_ (.Y(_0564_),
    .B1(net282),
    .B2(\s.hidden ),
    .A2(net287),
    .A1(\s.doubleOverline ));
 sg13g2_a21oi_1 _1244_ (.A1(\s.lg.yPostMirror ),
    .A2(net285),
    .Y(_0565_),
    .B1(net288));
 sg13g2_a22oi_1 _1245_ (.Y(uio_out[7]),
    .B1(_0564_),
    .B2(_0565_),
    .A2(_0563_),
    .A1(_0559_));
 sg13g2_nor2_2 _1246_ (.A(net8),
    .B(net288),
    .Y(_0566_));
 sg13g2_nand2_1 _1247_ (.Y(_0567_),
    .A(_0361_),
    .B(_0566_));
 sg13g2_o21ai_1 _1248_ (.B1(net291),
    .Y(_0568_),
    .A1(net9),
    .A2(_0567_));
 sg13g2_a21oi_1 _1249_ (.A1(_0104_),
    .A2(_0567_),
    .Y(_0006_),
    .B1(_0568_));
 sg13g2_nor2_2 _1250_ (.A(net8),
    .B(net3),
    .Y(_0569_));
 sg13g2_nand2_2 _1251_ (.Y(_0570_),
    .A(net285),
    .B(_0569_));
 sg13g2_o21ai_1 _1252_ (.B1(net296),
    .Y(_0571_),
    .A1(net9),
    .A2(_0570_));
 sg13g2_a21oi_1 _1253_ (.A1(_0103_),
    .A2(_0570_),
    .Y(_0007_),
    .B1(_0571_));
 sg13g2_o21ai_1 _1254_ (.B1(net296),
    .Y(_0572_),
    .A1(net10),
    .A2(_0570_));
 sg13g2_a21oi_1 _1255_ (.A1(_0102_),
    .A2(_0570_),
    .Y(_0008_),
    .B1(_0572_));
 sg13g2_o21ai_1 _1256_ (.B1(net298),
    .Y(_0573_),
    .A1(net11),
    .A2(_0570_));
 sg13g2_a21oi_1 _1257_ (.A1(_0101_),
    .A2(_0570_),
    .Y(_0009_),
    .B1(_0573_));
 sg13g2_o21ai_1 _1258_ (.B1(net298),
    .Y(_0574_),
    .A1(net12),
    .A2(_0570_));
 sg13g2_a21oi_1 _1259_ (.A1(_0100_),
    .A2(_0570_),
    .Y(_0010_),
    .B1(_0574_));
 sg13g2_and2_2 _1260_ (.A(net283),
    .B(_0569_),
    .X(_0575_));
 sg13g2_nand2_2 _1261_ (.Y(_0576_),
    .A(net283),
    .B(_0569_));
 sg13g2_o21ai_1 _1262_ (.B1(net296),
    .Y(_0577_),
    .A1(net110),
    .A2(_0575_));
 sg13g2_a21oi_1 _1263_ (.A1(_0074_),
    .A2(_0575_),
    .Y(_0011_),
    .B1(_0577_));
 sg13g2_o21ai_1 _1264_ (.B1(net296),
    .Y(_0578_),
    .A1(net114),
    .A2(_0575_));
 sg13g2_a21oi_1 _1265_ (.A1(_0072_),
    .A2(_0575_),
    .Y(_0012_),
    .B1(_0578_));
 sg13g2_o21ai_1 _1266_ (.B1(net296),
    .Y(_0579_),
    .A1(_0070_),
    .A2(_0576_));
 sg13g2_a21o_1 _1267_ (.A2(_0576_),
    .A1(net99),
    .B1(_0579_),
    .X(_0013_));
 sg13g2_o21ai_1 _1268_ (.B1(net296),
    .Y(_0580_),
    .A1(_0068_),
    .A2(_0576_));
 sg13g2_a21o_1 _1269_ (.A2(_0576_),
    .A1(net92),
    .B1(_0580_),
    .X(_0014_));
 sg13g2_o21ai_1 _1270_ (.B1(net293),
    .Y(_0581_),
    .A1(_0066_),
    .A2(_0576_));
 sg13g2_a21o_1 _1271_ (.A2(_0576_),
    .A1(net113),
    .B1(_0581_),
    .X(_0015_));
 sg13g2_o21ai_1 _1272_ (.B1(net296),
    .Y(_0582_),
    .A1(_0064_),
    .A2(_0576_));
 sg13g2_a21o_1 _1273_ (.A2(_0576_),
    .A1(net109),
    .B1(_0582_),
    .X(_0016_));
 sg13g2_o21ai_1 _1274_ (.B1(net293),
    .Y(_0583_),
    .A1(net117),
    .A2(_0575_));
 sg13g2_a21oi_1 _1275_ (.A1(_0062_),
    .A2(_0575_),
    .Y(_0017_),
    .B1(_0583_));
 sg13g2_o21ai_1 _1276_ (.B1(net296),
    .Y(_0584_),
    .A1(net112),
    .A2(_0575_));
 sg13g2_a21oi_1 _1277_ (.A1(_0060_),
    .A2(_0575_),
    .Y(_0018_),
    .B1(_0584_));
 sg13g2_nand2_1 _1278_ (.Y(_0585_),
    .A(net287),
    .B(_0569_));
 sg13g2_o21ai_1 _1279_ (.B1(net293),
    .Y(_0586_),
    .A1(net9),
    .A2(net260));
 sg13g2_a21oi_1 _1280_ (.A1(_0098_),
    .A2(net260),
    .Y(_0019_),
    .B1(_0586_));
 sg13g2_o21ai_1 _1281_ (.B1(net293),
    .Y(_0587_),
    .A1(net10),
    .A2(net260));
 sg13g2_a21oi_1 _1282_ (.A1(_0097_),
    .A2(net260),
    .Y(_0020_),
    .B1(_0587_));
 sg13g2_o21ai_1 _1283_ (.B1(net295),
    .Y(_0588_),
    .A1(net11),
    .A2(net260));
 sg13g2_a21oi_1 _1284_ (.A1(_0096_),
    .A2(net260),
    .Y(_0021_),
    .B1(_0588_));
 sg13g2_o21ai_1 _1285_ (.B1(net293),
    .Y(_0589_),
    .A1(net12),
    .A2(net260));
 sg13g2_a21oi_1 _1286_ (.A1(_0095_),
    .A2(net259),
    .Y(_0022_),
    .B1(_0589_));
 sg13g2_o21ai_1 _1287_ (.B1(net294),
    .Y(_0590_),
    .A1(net13),
    .A2(net259));
 sg13g2_a21oi_1 _1288_ (.A1(_0094_),
    .A2(net259),
    .Y(_0023_),
    .B1(_0590_));
 sg13g2_o21ai_1 _1289_ (.B1(net294),
    .Y(_0591_),
    .A1(net14),
    .A2(net259));
 sg13g2_a21oi_1 _1290_ (.A1(_0093_),
    .A2(net259),
    .Y(_0024_),
    .B1(_0591_));
 sg13g2_o21ai_1 _1291_ (.B1(net294),
    .Y(_0592_),
    .A1(net15),
    .A2(net259));
 sg13g2_a21oi_1 _1292_ (.A1(_0092_),
    .A2(net259),
    .Y(_0025_),
    .B1(_0592_));
 sg13g2_o21ai_1 _1293_ (.B1(net293),
    .Y(_0593_),
    .A1(net16),
    .A2(net260));
 sg13g2_a21oi_1 _1294_ (.A1(_0091_),
    .A2(net259),
    .Y(_0026_),
    .B1(_0593_));
 sg13g2_nand2_1 _1295_ (.Y(_0594_),
    .A(net285),
    .B(_0566_));
 sg13g2_o21ai_1 _1296_ (.B1(net292),
    .Y(_0595_),
    .A1(net9),
    .A2(net244));
 sg13g2_a21oi_1 _1297_ (.A1(net263),
    .A2(net244),
    .Y(_0027_),
    .B1(_0595_));
 sg13g2_o21ai_1 _1298_ (.B1(net292),
    .Y(_0596_),
    .A1(net10),
    .A2(net244));
 sg13g2_a21oi_1 _1299_ (.A1(net264),
    .A2(net244),
    .Y(_0028_),
    .B1(_0596_));
 sg13g2_o21ai_1 _1300_ (.B1(net295),
    .Y(_0597_),
    .A1(net11),
    .A2(net242));
 sg13g2_a21oi_1 _1301_ (.A1(_0088_),
    .A2(net242),
    .Y(_0029_),
    .B1(_0597_));
 sg13g2_o21ai_1 _1302_ (.B1(net297),
    .Y(_0598_),
    .A1(net12),
    .A2(net242));
 sg13g2_a21oi_1 _1303_ (.A1(_0087_),
    .A2(net242),
    .Y(_0030_),
    .B1(_0598_));
 sg13g2_o21ai_1 _1304_ (.B1(net295),
    .Y(_0599_),
    .A1(net13),
    .A2(net242));
 sg13g2_a21oi_1 _1305_ (.A1(_0086_),
    .A2(net242),
    .Y(_0031_),
    .B1(_0599_));
 sg13g2_o21ai_1 _1306_ (.B1(net291),
    .Y(_0600_),
    .A1(net14),
    .A2(net243));
 sg13g2_a21oi_1 _1307_ (.A1(net267),
    .A2(net244),
    .Y(_0032_),
    .B1(_0600_));
 sg13g2_o21ai_1 _1308_ (.B1(net297),
    .Y(_0601_),
    .A1(net15),
    .A2(net243));
 sg13g2_a21oi_1 _1309_ (.A1(_0084_),
    .A2(net243),
    .Y(_0033_),
    .B1(_0601_));
 sg13g2_o21ai_1 _1310_ (.B1(net297),
    .Y(_0602_),
    .A1(net16),
    .A2(net242));
 sg13g2_a21oi_1 _1311_ (.A1(_0083_),
    .A2(net242),
    .Y(_0034_),
    .B1(_0602_));
 sg13g2_nand2_1 _1312_ (.Y(_0603_),
    .A(net282),
    .B(_0566_));
 sg13g2_o21ai_1 _1313_ (.B1(net292),
    .Y(_0604_),
    .A1(net9),
    .A2(net241));
 sg13g2_a21oi_1 _1314_ (.A1(_0082_),
    .A2(net241),
    .Y(_0035_),
    .B1(_0604_));
 sg13g2_o21ai_1 _1315_ (.B1(net291),
    .Y(_0605_),
    .A1(net10),
    .A2(net241));
 sg13g2_a21oi_1 _1316_ (.A1(_0081_),
    .A2(net241),
    .Y(_0036_),
    .B1(_0605_));
 sg13g2_o21ai_1 _1317_ (.B1(net292),
    .Y(_0606_),
    .A1(net11),
    .A2(net240));
 sg13g2_a21oi_1 _1318_ (.A1(_0080_),
    .A2(net240),
    .Y(_0037_),
    .B1(_0606_));
 sg13g2_o21ai_1 _1319_ (.B1(net292),
    .Y(_0607_),
    .A1(net12),
    .A2(net240));
 sg13g2_a21oi_1 _1320_ (.A1(_0079_),
    .A2(net240),
    .Y(_0038_),
    .B1(_0607_));
 sg13g2_o21ai_1 _1321_ (.B1(net297),
    .Y(_0608_),
    .A1(net13),
    .A2(_0603_));
 sg13g2_a21oi_1 _1322_ (.A1(_0078_),
    .A2(net241),
    .Y(_0039_),
    .B1(_0608_));
 sg13g2_o21ai_1 _1323_ (.B1(net297),
    .Y(_0609_),
    .A1(net14),
    .A2(net240));
 sg13g2_a21oi_1 _1324_ (.A1(_0077_),
    .A2(net240),
    .Y(_0040_),
    .B1(_0609_));
 sg13g2_o21ai_1 _1325_ (.B1(net297),
    .Y(_0610_),
    .A1(net15),
    .A2(net240));
 sg13g2_a21oi_1 _1326_ (.A1(_0076_),
    .A2(net240),
    .Y(_0041_),
    .B1(_0610_));
 sg13g2_o21ai_1 _1327_ (.B1(net290),
    .Y(_0611_),
    .A1(net16),
    .A2(net241));
 sg13g2_a21oi_1 _1328_ (.A1(_0075_),
    .A2(net241),
    .Y(_0042_),
    .B1(_0611_));
 sg13g2_and2_1 _1329_ (.A(_0361_),
    .B(_0569_),
    .X(_0612_));
 sg13g2_o21ai_1 _1330_ (.B1(net294),
    .Y(_0613_),
    .A1(net106),
    .A2(net257));
 sg13g2_a21oi_1 _1331_ (.A1(_0074_),
    .A2(net257),
    .Y(_0043_),
    .B1(_0613_));
 sg13g2_o21ai_1 _1332_ (.B1(net294),
    .Y(_0614_),
    .A1(net102),
    .A2(net257));
 sg13g2_a21oi_1 _1333_ (.A1(_0072_),
    .A2(net257),
    .Y(_0044_),
    .B1(_0614_));
 sg13g2_o21ai_1 _1334_ (.B1(net294),
    .Y(_0615_),
    .A1(net104),
    .A2(net257));
 sg13g2_a21oi_1 _1335_ (.A1(_0070_),
    .A2(net257),
    .Y(_0045_),
    .B1(_0615_));
 sg13g2_o21ai_1 _1336_ (.B1(net294),
    .Y(_0616_),
    .A1(net103),
    .A2(net257));
 sg13g2_a21oi_1 _1337_ (.A1(_0068_),
    .A2(_0612_),
    .Y(_0046_),
    .B1(_0616_));
 sg13g2_o21ai_1 _1338_ (.B1(net294),
    .Y(_0617_),
    .A1(net100),
    .A2(net258));
 sg13g2_a21oi_1 _1339_ (.A1(_0066_),
    .A2(net257),
    .Y(_0047_),
    .B1(_0617_));
 sg13g2_o21ai_1 _1340_ (.B1(net293),
    .Y(_0618_),
    .A1(net98),
    .A2(net258));
 sg13g2_a21oi_1 _1341_ (.A1(_0064_),
    .A2(net258),
    .Y(_0048_),
    .B1(_0618_));
 sg13g2_o21ai_1 _1342_ (.B1(net295),
    .Y(_0619_),
    .A1(net76),
    .A2(net258));
 sg13g2_a21oi_1 _1343_ (.A1(_0062_),
    .A2(net258),
    .Y(_0049_),
    .B1(_0619_));
 sg13g2_o21ai_1 _1344_ (.B1(net293),
    .Y(_0620_),
    .A1(net82),
    .A2(net258));
 sg13g2_a21oi_1 _1345_ (.A1(_0060_),
    .A2(net258),
    .Y(_0050_),
    .B1(_0620_));
 sg13g2_nand2_1 _1346_ (.Y(_0621_),
    .A(net287),
    .B(_0566_));
 sg13g2_o21ai_1 _1347_ (.B1(net290),
    .Y(_0622_),
    .A1(net9),
    .A2(net238));
 sg13g2_a21oi_1 _1348_ (.A1(_0073_),
    .A2(net238),
    .Y(_0051_),
    .B1(_0622_));
 sg13g2_o21ai_1 _1349_ (.B1(net290),
    .Y(_0623_),
    .A1(net10),
    .A2(net238));
 sg13g2_a21oi_1 _1350_ (.A1(_0071_),
    .A2(net238),
    .Y(_0052_),
    .B1(_0623_));
 sg13g2_o21ai_1 _1351_ (.B1(net290),
    .Y(_0624_),
    .A1(net11),
    .A2(net238));
 sg13g2_a21oi_1 _1352_ (.A1(_0069_),
    .A2(net238),
    .Y(_0053_),
    .B1(_0624_));
 sg13g2_o21ai_1 _1353_ (.B1(net290),
    .Y(_0625_),
    .A1(net12),
    .A2(net239));
 sg13g2_a21oi_1 _1354_ (.A1(_0067_),
    .A2(net239),
    .Y(_0054_),
    .B1(_0625_));
 sg13g2_o21ai_1 _1355_ (.B1(net297),
    .Y(_0626_),
    .A1(net13),
    .A2(net239));
 sg13g2_a21oi_1 _1356_ (.A1(_0065_),
    .A2(net239),
    .Y(_0055_),
    .B1(_0626_));
 sg13g2_o21ai_1 _1357_ (.B1(net290),
    .Y(_0627_),
    .A1(net14),
    .A2(net239));
 sg13g2_a21oi_1 _1358_ (.A1(_0063_),
    .A2(net239),
    .Y(_0056_),
    .B1(_0627_));
 sg13g2_o21ai_1 _1359_ (.B1(net290),
    .Y(_0628_),
    .A1(net15),
    .A2(net239));
 sg13g2_a21oi_1 _1360_ (.A1(_0061_),
    .A2(net239),
    .Y(_0057_),
    .B1(_0628_));
 sg13g2_o21ai_1 _1361_ (.B1(net290),
    .Y(_0629_),
    .A1(net16),
    .A2(net238));
 sg13g2_a21oi_1 _1362_ (.A1(_0059_),
    .A2(net238),
    .Y(_0058_),
    .B1(_0629_));
 sg13g2_dfrbp_1 _1363_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net66),
    .D(_0006_),
    .Q_N(_0676_),
    .Q(\s.dottedOverline ));
 sg13g2_dfrbp_1 _1364_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net54),
    .D(_0007_),
    .Q_N(_0675_),
    .Q(\s.lg.s0[0] ));
 sg13g2_dfrbp_1 _1365_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net52),
    .D(_0008_),
    .Q_N(_0674_),
    .Q(\s.lg.s0[1] ));
 sg13g2_dfrbp_1 _1366_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net50),
    .D(_0009_),
    .Q_N(_0673_),
    .Q(\s.lg.s0[2] ));
 sg13g2_dfrbp_1 _1367_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net48),
    .D(_0010_),
    .Q_N(_0672_),
    .Q(\s.lg.s0[3] ));
 sg13g2_dfrbp_1 _1368_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net46),
    .D(_0011_),
    .Q_N(_0671_),
    .Q(\ctrl[0] ));
 sg13g2_dfrbp_1 _1369_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net44),
    .D(_0012_),
    .Q_N(_0670_),
    .Q(\ctrl[1] ));
 sg13g2_dfrbp_1 _1370_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net42),
    .D(_0013_),
    .Q_N(_0669_),
    .Q(\ctrl[2] ));
 sg13g2_dfrbp_1 _1371_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net40),
    .D(_0014_),
    .Q_N(_0668_),
    .Q(\ctrl[3] ));
 sg13g2_dfrbp_1 _1372_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net38),
    .D(_0015_),
    .Q_N(_0667_),
    .Q(\ctrl[4] ));
 sg13g2_dfrbp_1 _1373_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net36),
    .D(_0016_),
    .Q_N(_0666_),
    .Q(\ctrl[5] ));
 sg13g2_dfrbp_1 _1374_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net34),
    .D(_0017_),
    .Q_N(_0665_),
    .Q(\ctrl[6] ));
 sg13g2_dfrbp_1 _1375_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net32),
    .D(_0018_),
    .Q_N(_0664_),
    .Q(\ctrl[7] ));
 sg13g2_dfrbp_1 _1376_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net30),
    .D(_0019_),
    .Q_N(_0002_),
    .Q(\bitmapIn[0] ));
 sg13g2_dfrbp_1 _1377_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net28),
    .D(_0020_),
    .Q_N(_0004_),
    .Q(\bitmapIn[1] ));
 sg13g2_dfrbp_1 _1378_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net26),
    .D(_0021_),
    .Q_N(_0663_),
    .Q(\bitmapIn[2] ));
 sg13g2_dfrbp_1 _1379_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net24),
    .D(_0022_),
    .Q_N(_0662_),
    .Q(\bitmapIn[3] ));
 sg13g2_dfrbp_1 _1380_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net22),
    .D(_0023_),
    .Q_N(_0661_),
    .Q(\bitmapIn[4] ));
 sg13g2_dfrbp_1 _1381_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net20),
    .D(_0024_),
    .Q_N(_0660_),
    .Q(\bitmapIn[5] ));
 sg13g2_dfrbp_1 _1382_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net18),
    .D(_0025_),
    .Q_N(_0659_),
    .Q(\bitmapIn[6] ));
 sg13g2_dfrbp_1 _1383_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net69),
    .D(_0026_),
    .Q_N(_0658_),
    .Q(\bitmapIn[7] ));
 sg13g2_dfrbp_1 _1384_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net67),
    .D(_0027_),
    .Q_N(_0657_),
    .Q(\s.sty.xoffset ));
 sg13g2_dfrbp_1 _1385_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net65),
    .D(_0028_),
    .Q_N(_0656_),
    .Q(\s.sty.xscale ));
 sg13g2_dfrbp_1 _1386_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net63),
    .D(_0029_),
    .Q_N(_0655_),
    .Q(\s.lg.yoffset ));
 sg13g2_dfrbp_1 _1387_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net61),
    .D(_0030_),
    .Q_N(_0001_),
    .Q(\s.lg.yscale ));
 sg13g2_dfrbp_1 _1388_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net59),
    .D(_0031_),
    .Q_N(_0654_),
    .Q(\s.sty.xPreMirror ));
 sg13g2_dfrbp_1 _1389_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net57),
    .D(_0032_),
    .Q_N(_0653_),
    .Q(\s.inv.xPostMirror ));
 sg13g2_dfrbp_1 _1390_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net55),
    .D(_0033_),
    .Q_N(_0000_),
    .Q(\s.lg.yPreMirror ));
 sg13g2_dfrbp_1 _1391_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net51),
    .D(_0034_),
    .Q_N(_0652_),
    .Q(\s.lg.yPostMirror ));
 sg13g2_dfrbp_1 _1392_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net47),
    .D(_0035_),
    .Q_N(_0651_),
    .Q(\s.bold ));
 sg13g2_dfrbp_1 _1393_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net43),
    .D(_0036_),
    .Q_N(_0650_),
    .Q(\s.faint ));
 sg13g2_dfrbp_1 _1394_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net39),
    .D(_0037_),
    .Q_N(_0649_),
    .Q(\s.italic ));
 sg13g2_dfrbp_1 _1395_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net35),
    .D(_0038_),
    .Q_N(_0648_),
    .Q(\s.reverseItalic ));
 sg13g2_dfrbp_1 _1396_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net31),
    .D(_0039_),
    .Q_N(_0647_),
    .Q(\s.blink ));
 sg13g2_dfrbp_1 _1397_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net27),
    .D(_0040_),
    .Q_N(_0646_),
    .Q(\s.alternate ));
 sg13g2_dfrbp_1 _1398_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net23),
    .D(_0041_),
    .Q_N(_0645_),
    .Q(\s.inverse ));
 sg13g2_dfrbp_1 _1399_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net19),
    .D(_0042_),
    .Q_N(_0644_),
    .Q(\s.hidden ));
 sg13g2_dfrbp_1 _1400_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net68),
    .D(_0043_),
    .Q_N(_0643_),
    .Q(\bitmapIn[8] ));
 sg13g2_dfrbp_1 _1401_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net64),
    .D(_0044_),
    .Q_N(_0642_),
    .Q(\bitmapIn[9] ));
 sg13g2_dfrbp_1 _1402_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net60),
    .D(_0045_),
    .Q_N(_0641_),
    .Q(\bitmapIn[10] ));
 sg13g2_dfrbp_1 _1403_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net56),
    .D(_0046_),
    .Q_N(_0640_),
    .Q(\bitmapIn[11] ));
 sg13g2_dfrbp_1 _1404_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net49),
    .D(_0047_),
    .Q_N(_0639_),
    .Q(\bitmapIn[12] ));
 sg13g2_dfrbp_1 _1405_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net41),
    .D(_0048_),
    .Q_N(_0638_),
    .Q(\bitmapIn[13] ));
 sg13g2_dfrbp_1 _1406_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net33),
    .D(_0049_),
    .Q_N(_0005_),
    .Q(\bitmapIn[14] ));
 sg13g2_dfrbp_1 _1407_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net25),
    .D(_0050_),
    .Q_N(_0003_),
    .Q(\bitmapIn[15] ));
 sg13g2_dfrbp_1 _1408_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net17),
    .D(_0051_),
    .Q_N(_0637_),
    .Q(\s.lg.underline ));
 sg13g2_dfrbp_1 _1409_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net62),
    .D(_0052_),
    .Q_N(_0636_),
    .Q(\s.doubleUnderline ));
 sg13g2_dfrbp_1 _1410_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net53),
    .D(_0053_),
    .Q_N(_0635_),
    .Q(\s.dottedUnderline ));
 sg13g2_dfrbp_1 _1411_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net37),
    .D(_0054_),
    .Q_N(_0634_),
    .Q(\s.lg.strikethru ));
 sg13g2_dfrbp_1 _1412_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net21),
    .D(_0055_),
    .Q_N(_0633_),
    .Q(\s.doubleStrikethru ));
 sg13g2_dfrbp_1 _1413_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net58),
    .D(_0056_),
    .Q_N(_0632_),
    .Q(\s.dottedStrikethru ));
 sg13g2_dfrbp_1 _1414_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net29),
    .D(_0057_),
    .Q_N(_0631_),
    .Q(\s.lg.overline ));
 sg13g2_dfrbp_1 _1415_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net45),
    .D(_0058_),
    .Q_N(_0630_),
    .Q(\s.doubleOverline ));
 sg13g2_tiehi _1382__18 (.L_HI(net18));
 sg13g2_tiehi _1399__19 (.L_HI(net19));
 sg13g2_tiehi _1381__20 (.L_HI(net20));
 sg13g2_tiehi _1412__21 (.L_HI(net21));
 sg13g2_tiehi _1380__22 (.L_HI(net22));
 sg13g2_tiehi _1398__23 (.L_HI(net23));
 sg13g2_tiehi _1379__24 (.L_HI(net24));
 sg13g2_tiehi _1407__25 (.L_HI(net25));
 sg13g2_tiehi _1378__26 (.L_HI(net26));
 sg13g2_tiehi _1397__27 (.L_HI(net27));
 sg13g2_tiehi _1377__28 (.L_HI(net28));
 sg13g2_tiehi _1414__29 (.L_HI(net29));
 sg13g2_tiehi _1376__30 (.L_HI(net30));
 sg13g2_tiehi _1396__31 (.L_HI(net31));
 sg13g2_tiehi _1375__32 (.L_HI(net32));
 sg13g2_tiehi _1406__33 (.L_HI(net33));
 sg13g2_tiehi _1374__34 (.L_HI(net34));
 sg13g2_tiehi _1395__35 (.L_HI(net35));
 sg13g2_tiehi _1373__36 (.L_HI(net36));
 sg13g2_tiehi _1411__37 (.L_HI(net37));
 sg13g2_tiehi _1372__38 (.L_HI(net38));
 sg13g2_tiehi _1394__39 (.L_HI(net39));
 sg13g2_tiehi _1371__40 (.L_HI(net40));
 sg13g2_tiehi _1405__41 (.L_HI(net41));
 sg13g2_tiehi _1370__42 (.L_HI(net42));
 sg13g2_tiehi _1393__43 (.L_HI(net43));
 sg13g2_tiehi _1369__44 (.L_HI(net44));
 sg13g2_tiehi _1415__45 (.L_HI(net45));
 sg13g2_tiehi _1368__46 (.L_HI(net46));
 sg13g2_tiehi _1392__47 (.L_HI(net47));
 sg13g2_tiehi _1367__48 (.L_HI(net48));
 sg13g2_tiehi _1404__49 (.L_HI(net49));
 sg13g2_tiehi _1366__50 (.L_HI(net50));
 sg13g2_tiehi _1391__51 (.L_HI(net51));
 sg13g2_tiehi _1365__52 (.L_HI(net52));
 sg13g2_tiehi _1410__53 (.L_HI(net53));
 sg13g2_tiehi _1364__54 (.L_HI(net54));
 sg13g2_tiehi _1390__55 (.L_HI(net55));
 sg13g2_tiehi _1403__56 (.L_HI(net56));
 sg13g2_tiehi _1389__57 (.L_HI(net57));
 sg13g2_tiehi _1413__58 (.L_HI(net58));
 sg13g2_tiehi _1388__59 (.L_HI(net59));
 sg13g2_tiehi _1402__60 (.L_HI(net60));
 sg13g2_tiehi _1387__61 (.L_HI(net61));
 sg13g2_tiehi _1409__62 (.L_HI(net62));
 sg13g2_tiehi _1386__63 (.L_HI(net63));
 sg13g2_tiehi _1401__64 (.L_HI(net64));
 sg13g2_tiehi _1385__65 (.L_HI(net65));
 sg13g2_tiehi _1363__66 (.L_HI(net66));
 sg13g2_tiehi _1384__67 (.L_HI(net67));
 sg13g2_tiehi _1400__68 (.L_HI(net68));
 sg13g2_tiehi _1383__69 (.L_HI(net69));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _1469_ (.A(uio_oe[7]),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1470_ (.A(uio_oe[7]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1471_ (.A(uio_oe[7]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1472_ (.A(uio_oe[7]),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1473_ (.A(uio_oe[7]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1474_ (.A(uio_oe[7]),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1475_ (.A(uio_oe[7]),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1476_ (.A(uio_out[0]),
    .X(uo_out[0]));
 sg13g2_buf_1 _1477_ (.A(uio_out[1]),
    .X(uo_out[1]));
 sg13g2_buf_1 _1478_ (.A(uio_out[2]),
    .X(uo_out[2]));
 sg13g2_buf_1 _1479_ (.A(uio_out[3]),
    .X(uo_out[3]));
 sg13g2_buf_1 _1480_ (.A(uio_out[4]),
    .X(uo_out[4]));
 sg13g2_buf_1 _1481_ (.A(uio_out[5]),
    .X(uo_out[5]));
 sg13g2_buf_1 _1482_ (.A(uio_out[6]),
    .X(uo_out[6]));
 sg13g2_buf_1 _1483_ (.A(uio_out[7]),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout226 (.X(net226),
    .A(net227));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(_0119_));
 sg13g2_buf_2 fanout228 (.A(_0179_),
    .X(net228));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(_0178_));
 sg13g2_buf_2 fanout230 (.A(net232),
    .X(net230));
 sg13g2_buf_1 fanout231 (.A(net232),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(net233),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_0151_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(net236),
    .X(net234));
 sg13g2_buf_1 fanout235 (.A(net236),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(net237),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_0138_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_0621_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_0621_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_0603_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(net243),
    .X(net242));
 sg13g2_buf_1 fanout243 (.A(net244),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_0594_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_0190_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_0177_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_0177_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(net249),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(_0147_));
 sg13g2_buf_2 fanout251 (.A(net252),
    .X(net251));
 sg13g2_buf_1 fanout252 (.A(net254),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net254),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_0146_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_0136_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_0135_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(net258),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_0612_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_0585_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_0585_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(net262),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_0226_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_0090_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_0089_),
    .X(net264));
 sg13g2_buf_1 fanout265 (.A(_0089_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(net267),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_0085_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(net269),
    .X(net268));
 sg13g2_buf_1 fanout269 (.A(net270),
    .X(net269));
 sg13g2_buf_1 fanout270 (.A(\s.bold ),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(net272),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(\s.inv.xPostMirror ),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_buf_1 fanout274 (.A(net275),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(net276),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(net277),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(\s.sty.xPreMirror ),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(\s.sty.xscale ),
    .X(net278));
 sg13g2_buf_1 fanout279 (.A(\s.sty.xscale ),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(\s.sty.xoffset ),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(net284),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(net284),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_0432_),
    .X(net284));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_0430_));
 sg13g2_buf_2 fanout286 (.A(_0430_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_0423_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_0105_),
    .X(net288));
 sg13g2_buf_1 fanout289 (.A(_0105_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net291),
    .X(net290));
 sg13g2_buf_1 fanout291 (.A(net292),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(rst_n),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net295),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(net295),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(net298),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(net297),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(net298),
    .X(net297));
 sg13g2_buf_1 fanout298 (.A(rst_n),
    .X(net298));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[2]));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_4 input9 (.X(net9),
    .A(uio_in[0]));
 sg13g2_buf_4 input10 (.X(net10),
    .A(uio_in[1]));
 sg13g2_buf_4 input11 (.X(net11),
    .A(uio_in[2]));
 sg13g2_buf_2 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_2 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_2 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_2 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tiehi _1408__17 (.L_HI(net17));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\bitmapIn[0] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold2 (.A(\bitmapIn[1] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold3 (.A(\s.lg.yPreMirror ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold4 (.A(\bitmapIn[3] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold5 (.A(\bitmapIn[5] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold6 (.A(\bitmapIn[2] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold7 (.A(\bitmapIn[14] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold8 (.A(\s.blink ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold9 (.A(\s.doubleStrikethru ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold10 (.A(\s.bold ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold11 (.A(\s.faint ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold12 (.A(\s.alternate ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold13 (.A(\bitmapIn[15] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold14 (.A(\bitmapIn[4] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold15 (.A(\s.dottedStrikethru ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold16 (.A(\s.doubleOverline ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold17 (.A(\bitmapIn[7] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold18 (.A(\s.dottedUnderline ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold19 (.A(\s.dottedOverline ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold20 (.A(\s.lg.overline ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold21 (.A(\s.hidden ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold22 (.A(\s.lg.strikethru ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold23 (.A(\ctrl[3] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold24 (.A(\s.doubleUnderline ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold25 (.A(\s.inverse ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold26 (.A(\s.lg.underline ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold27 (.A(\bitmapIn[6] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold28 (.A(\s.lg.s0[0] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold29 (.A(\bitmapIn[13] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold30 (.A(\ctrl[2] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold31 (.A(\bitmapIn[12] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold32 (.A(\s.lg.s0[1] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold33 (.A(\bitmapIn[9] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold34 (.A(\bitmapIn[11] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold35 (.A(\bitmapIn[10] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold36 (.A(\s.lg.s0[3] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold37 (.A(\bitmapIn[8] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold38 (.A(\s.lg.s0[2] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold39 (.A(\s.italic ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold40 (.A(\ctrl[5] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold41 (.A(\ctrl[0] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold42 (.A(\s.reverseItalic ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold43 (.A(\ctrl[7] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold44 (.A(\ctrl[4] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold45 (.A(\ctrl[1] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold46 (.A(\s.lg.yoffset ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold47 (.A(\s.lg.yscale ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold48 (.A(\ctrl[6] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold49 (.A(\s.lg.yPostMirror ),
    .X(net118));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_4 FILLER_14_196 ();
 sg13g2_fill_1 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_8 FILLER_14_213 ();
 sg13g2_decap_8 FILLER_14_220 ();
 sg13g2_decap_8 FILLER_14_227 ();
 sg13g2_decap_8 FILLER_14_234 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_decap_8 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_255 ();
 sg13g2_decap_8 FILLER_14_262 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_decap_8 FILLER_14_276 ();
 sg13g2_decap_8 FILLER_14_283 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_decap_8 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_decap_4 FILLER_15_173 ();
 sg13g2_decap_4 FILLER_15_188 ();
 sg13g2_decap_4 FILLER_15_235 ();
 sg13g2_fill_2 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_262 ();
 sg13g2_fill_1 FILLER_15_278 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_fill_2 FILLER_15_308 ();
 sg13g2_fill_1 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_344 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_fill_2 FILLER_15_358 ();
 sg13g2_fill_1 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_fill_2 FILLER_16_175 ();
 sg13g2_decap_4 FILLER_16_193 ();
 sg13g2_decap_4 FILLER_16_219 ();
 sg13g2_decap_4 FILLER_16_234 ();
 sg13g2_decap_4 FILLER_16_260 ();
 sg13g2_decap_4 FILLER_16_270 ();
 sg13g2_fill_2 FILLER_16_282 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_321 ();
 sg13g2_fill_1 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_179 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_decap_4 FILLER_17_200 ();
 sg13g2_fill_1 FILLER_17_204 ();
 sg13g2_decap_4 FILLER_17_209 ();
 sg13g2_fill_2 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_fill_2 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_264 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_296 ();
 sg13g2_fill_2 FILLER_17_303 ();
 sg13g2_fill_1 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_327 ();
 sg13g2_fill_2 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_fill_2 FILLER_17_373 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_fill_2 FILLER_18_112 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_139 ();
 sg13g2_fill_2 FILLER_18_146 ();
 sg13g2_fill_2 FILLER_18_177 ();
 sg13g2_fill_1 FILLER_18_217 ();
 sg13g2_decap_4 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_241 ();
 sg13g2_fill_1 FILLER_18_253 ();
 sg13g2_decap_4 FILLER_18_270 ();
 sg13g2_fill_1 FILLER_18_274 ();
 sg13g2_fill_1 FILLER_18_280 ();
 sg13g2_decap_4 FILLER_18_298 ();
 sg13g2_fill_2 FILLER_18_302 ();
 sg13g2_fill_2 FILLER_18_317 ();
 sg13g2_fill_1 FILLER_18_330 ();
 sg13g2_decap_4 FILLER_18_362 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_136 ();
 sg13g2_fill_1 FILLER_19_138 ();
 sg13g2_fill_1 FILLER_19_155 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_4 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_208 ();
 sg13g2_fill_1 FILLER_19_214 ();
 sg13g2_decap_4 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_decap_4 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_248 ();
 sg13g2_decap_4 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_fill_2 FILLER_19_312 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_fill_1 FILLER_19_329 ();
 sg13g2_fill_2 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_353 ();
 sg13g2_fill_1 FILLER_19_355 ();
 sg13g2_decap_4 FILLER_19_370 ();
 sg13g2_decap_4 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_4 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_1 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_134 ();
 sg13g2_decap_8 FILLER_20_141 ();
 sg13g2_fill_2 FILLER_20_158 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_fill_2 FILLER_20_202 ();
 sg13g2_fill_1 FILLER_20_204 ();
 sg13g2_fill_1 FILLER_20_208 ();
 sg13g2_decap_8 FILLER_20_213 ();
 sg13g2_fill_2 FILLER_20_220 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_decap_4 FILLER_20_237 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_254 ();
 sg13g2_decap_8 FILLER_20_260 ();
 sg13g2_decap_4 FILLER_20_267 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_295 ();
 sg13g2_decap_4 FILLER_20_302 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_fill_1 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_391 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_103 ();
 sg13g2_fill_2 FILLER_21_115 ();
 sg13g2_fill_1 FILLER_21_129 ();
 sg13g2_fill_2 FILLER_21_151 ();
 sg13g2_fill_1 FILLER_21_153 ();
 sg13g2_fill_2 FILLER_21_164 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_180 ();
 sg13g2_fill_2 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_254 ();
 sg13g2_fill_2 FILLER_21_264 ();
 sg13g2_decap_8 FILLER_21_304 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_decap_4 FILLER_21_318 ();
 sg13g2_fill_2 FILLER_21_331 ();
 sg13g2_fill_1 FILLER_21_333 ();
 sg13g2_decap_4 FILLER_21_339 ();
 sg13g2_fill_1 FILLER_21_343 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_fill_1 FILLER_21_358 ();
 sg13g2_fill_2 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_370 ();
 sg13g2_fill_2 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_91 ();
 sg13g2_fill_2 FILLER_22_103 ();
 sg13g2_fill_1 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_4 FILLER_22_123 ();
 sg13g2_fill_2 FILLER_22_127 ();
 sg13g2_decap_8 FILLER_22_135 ();
 sg13g2_decap_8 FILLER_22_142 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_decap_4 FILLER_22_187 ();
 sg13g2_fill_2 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_fill_1 FILLER_22_262 ();
 sg13g2_decap_4 FILLER_22_285 ();
 sg13g2_fill_1 FILLER_22_289 ();
 sg13g2_decap_4 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_304 ();
 sg13g2_decap_4 FILLER_22_328 ();
 sg13g2_decap_4 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_345 ();
 sg13g2_fill_2 FILLER_22_352 ();
 sg13g2_fill_1 FILLER_22_354 ();
 sg13g2_fill_1 FILLER_22_363 ();
 sg13g2_fill_2 FILLER_22_369 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_fill_1 FILLER_23_97 ();
 sg13g2_decap_8 FILLER_23_111 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_fill_2 FILLER_23_185 ();
 sg13g2_decap_4 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_216 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_decap_8 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_decap_4 FILLER_23_285 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_4 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_312 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_decap_4 FILLER_23_367 ();
 sg13g2_fill_1 FILLER_23_371 ();
 sg13g2_decap_4 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_4 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_fill_2 FILLER_24_219 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_258 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_268 ();
 sg13g2_decap_4 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_315 ();
 sg13g2_decap_4 FILLER_24_321 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_379 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_81 ();
 sg13g2_decap_4 FILLER_25_88 ();
 sg13g2_fill_1 FILLER_25_92 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_decap_4 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_124 ();
 sg13g2_decap_8 FILLER_25_150 ();
 sg13g2_fill_2 FILLER_25_157 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_222 ();
 sg13g2_decap_4 FILLER_25_227 ();
 sg13g2_fill_1 FILLER_25_231 ();
 sg13g2_fill_1 FILLER_25_245 ();
 sg13g2_fill_1 FILLER_25_251 ();
 sg13g2_decap_8 FILLER_25_272 ();
 sg13g2_fill_2 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_302 ();
 sg13g2_fill_1 FILLER_25_337 ();
 sg13g2_decap_4 FILLER_25_351 ();
 sg13g2_decap_4 FILLER_25_367 ();
 sg13g2_fill_2 FILLER_25_371 ();
 sg13g2_fill_1 FILLER_25_378 ();
 sg13g2_fill_2 FILLER_25_389 ();
 sg13g2_fill_1 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_65 ();
 sg13g2_decap_4 FILLER_26_106 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_fill_2 FILLER_26_134 ();
 sg13g2_decap_8 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_226 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_260 ();
 sg13g2_fill_2 FILLER_26_341 ();
 sg13g2_fill_2 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_decap_4 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_fill_2 FILLER_27_104 ();
 sg13g2_decap_8 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_decap_4 FILLER_27_156 ();
 sg13g2_fill_1 FILLER_27_160 ();
 sg13g2_fill_2 FILLER_27_176 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_fill_2 FILLER_27_220 ();
 sg13g2_decap_4 FILLER_27_236 ();
 sg13g2_decap_4 FILLER_27_260 ();
 sg13g2_decap_4 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_281 ();
 sg13g2_fill_2 FILLER_27_288 ();
 sg13g2_fill_1 FILLER_27_290 ();
 sg13g2_fill_1 FILLER_27_337 ();
 sg13g2_decap_4 FILLER_27_342 ();
 sg13g2_fill_1 FILLER_27_368 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_4 FILLER_28_70 ();
 sg13g2_fill_1 FILLER_28_74 ();
 sg13g2_decap_8 FILLER_28_79 ();
 sg13g2_decap_4 FILLER_28_86 ();
 sg13g2_fill_1 FILLER_28_120 ();
 sg13g2_fill_2 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_158 ();
 sg13g2_fill_2 FILLER_28_165 ();
 sg13g2_fill_1 FILLER_28_167 ();
 sg13g2_fill_1 FILLER_28_197 ();
 sg13g2_fill_2 FILLER_28_250 ();
 sg13g2_decap_4 FILLER_28_283 ();
 sg13g2_fill_1 FILLER_28_291 ();
 sg13g2_decap_4 FILLER_28_323 ();
 sg13g2_fill_2 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_4 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_81 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_fill_1 FILLER_29_99 ();
 sg13g2_decap_4 FILLER_29_110 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_decap_4 FILLER_29_120 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_decap_8 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_137 ();
 sg13g2_fill_2 FILLER_29_144 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_decap_8 FILLER_29_173 ();
 sg13g2_decap_4 FILLER_29_180 ();
 sg13g2_fill_2 FILLER_29_184 ();
 sg13g2_decap_8 FILLER_29_191 ();
 sg13g2_decap_4 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_202 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_234 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_307 ();
 sg13g2_fill_1 FILLER_29_314 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_4 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_105 ();
 sg13g2_fill_2 FILLER_30_117 ();
 sg13g2_fill_1 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_157 ();
 sg13g2_decap_4 FILLER_30_163 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_decap_4 FILLER_30_212 ();
 sg13g2_fill_1 FILLER_30_216 ();
 sg13g2_decap_8 FILLER_30_233 ();
 sg13g2_decap_8 FILLER_30_240 ();
 sg13g2_fill_1 FILLER_30_247 ();
 sg13g2_fill_1 FILLER_30_272 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_79 ();
 sg13g2_fill_2 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_100 ();
 sg13g2_fill_2 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_fill_2 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_153 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_fill_1 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_209 ();
 sg13g2_decap_4 FILLER_31_216 ();
 sg13g2_decap_4 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_decap_4 FILLER_31_279 ();
 sg13g2_fill_2 FILLER_31_283 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_325 ();
 sg13g2_fill_1 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_384 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_84 ();
 sg13g2_decap_4 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_124 ();
 sg13g2_decap_4 FILLER_32_141 ();
 sg13g2_fill_1 FILLER_32_145 ();
 sg13g2_decap_8 FILLER_32_160 ();
 sg13g2_fill_2 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_decap_4 FILLER_32_183 ();
 sg13g2_fill_2 FILLER_32_187 ();
 sg13g2_decap_4 FILLER_32_234 ();
 sg13g2_fill_2 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_283 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_decap_8 FILLER_32_303 ();
 sg13g2_fill_2 FILLER_32_310 ();
 sg13g2_fill_2 FILLER_32_372 ();
 sg13g2_fill_1 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_100 ();
 sg13g2_decap_4 FILLER_33_109 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_decap_8 FILLER_33_122 ();
 sg13g2_fill_2 FILLER_33_129 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_decap_4 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_decap_4 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_decap_4 FILLER_33_181 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_fill_2 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_4 FILLER_33_249 ();
 sg13g2_fill_2 FILLER_33_253 ();
 sg13g2_fill_2 FILLER_33_260 ();
 sg13g2_fill_1 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_291 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_decap_4 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_341 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_110 ();
 sg13g2_fill_1 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_decap_4 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_193 ();
 sg13g2_decap_4 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_fill_2 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_4 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_121 ();
 sg13g2_fill_1 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_160 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_fill_1 FILLER_35_182 ();
 sg13g2_fill_2 FILLER_35_188 ();
 sg13g2_fill_2 FILLER_35_203 ();
 sg13g2_fill_2 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_319 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_fill_2 FILLER_35_388 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_4 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_135 ();
 sg13g2_decap_8 FILLER_36_142 ();
 sg13g2_fill_2 FILLER_36_149 ();
 sg13g2_fill_2 FILLER_36_160 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_decap_4 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_fill_2 FILLER_36_256 ();
 sg13g2_fill_1 FILLER_36_258 ();
 sg13g2_fill_1 FILLER_36_269 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_111 ();
 sg13g2_fill_2 FILLER_37_118 ();
 sg13g2_decap_8 FILLER_37_124 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_decap_4 FILLER_37_169 ();
 sg13g2_decap_4 FILLER_37_185 ();
 sg13g2_fill_2 FILLER_37_189 ();
 sg13g2_decap_4 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_200 ();
 sg13g2_fill_2 FILLER_37_238 ();
 sg13g2_fill_2 FILLER_37_247 ();
 sg13g2_fill_1 FILLER_37_249 ();
 sg13g2_fill_1 FILLER_37_295 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_115 ();
 sg13g2_decap_8 FILLER_38_122 ();
 sg13g2_decap_8 FILLER_38_129 ();
 sg13g2_decap_8 FILLER_38_136 ();
 sg13g2_decap_4 FILLER_38_143 ();
 sg13g2_fill_2 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_153 ();
 sg13g2_fill_2 FILLER_38_160 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_decap_4 FILLER_38_223 ();
 sg13g2_fill_2 FILLER_38_227 ();
 sg13g2_fill_1 FILLER_38_380 ();
 sg13g2_fill_2 FILLER_38_407 ();
endmodule

module tt_um_wokwi_411379488132926465 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net693;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net156;
 wire net187;
 wire net199;
 wire net218;
 wire net406;
 wire net412;
 wire net521;
 wire net526;
 wire net527;
 wire net553;
 wire net586;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire \flop1/_0_ ;
 wire \flop1/_1_ ;
 wire net641;
 wire net642;
 wire \flop10/_0_ ;
 wire \flop10/_1_ ;
 wire net643;
 wire net644;
 wire \flop11/_0_ ;
 wire \flop11/_1_ ;
 wire net645;
 wire net646;
 wire \flop12/_0_ ;
 wire \flop12/_1_ ;
 wire net647;
 wire net648;
 wire \flop13/_0_ ;
 wire \flop13/_1_ ;
 wire net649;
 wire net650;
 wire \flop14/_0_ ;
 wire \flop14/_1_ ;
 wire net651;
 wire net652;
 wire \flop15/_0_ ;
 wire \flop15/_1_ ;
 wire net653;
 wire net654;
 wire \flop16/_0_ ;
 wire \flop16/_1_ ;
 wire net655;
 wire net656;
 wire \flop17/_0_ ;
 wire \flop17/_1_ ;
 wire net657;
 wire net658;
 wire \flop18/_0_ ;
 wire \flop18/_1_ ;
 wire net659;
 wire net660;
 wire \flop19/_0_ ;
 wire \flop19/_1_ ;
 wire net661;
 wire net662;
 wire \flop2/_0_ ;
 wire \flop2/_1_ ;
 wire net663;
 wire net664;
 wire \flop20/_0_ ;
 wire \flop20/_1_ ;
 wire net665;
 wire net666;
 wire \flop21/_0_ ;
 wire \flop21/_1_ ;
 wire net667;
 wire net668;
 wire \flop22/_0_ ;
 wire \flop22/_1_ ;
 wire net669;
 wire net670;
 wire \flop23/_0_ ;
 wire \flop23/_1_ ;
 wire net671;
 wire net672;
 wire \flop24/_0_ ;
 wire \flop24/_1_ ;
 wire net673;
 wire net674;
 wire \flop25/_0_ ;
 wire \flop25/_1_ ;
 wire net675;
 wire net676;
 wire \flop26/_0_ ;
 wire \flop26/_1_ ;
 wire net677;
 wire net678;
 wire \flop26/notq ;
 wire \flop3/_0_ ;
 wire \flop3/_1_ ;
 wire net679;
 wire net680;
 wire \flop4/_0_ ;
 wire \flop4/_1_ ;
 wire net681;
 wire net682;
 wire \flop5/_0_ ;
 wire \flop5/_1_ ;
 wire net683;
 wire net684;
 wire \flop6/_0_ ;
 wire \flop6/_1_ ;
 wire net685;
 wire net686;
 wire \flop7/_0_ ;
 wire \flop7/_1_ ;
 wire net687;
 wire net688;
 wire \flop8/_0_ ;
 wire \flop8/_1_ ;
 wire net689;
 wire net690;
 wire \flop9/_0_ ;
 wire \flop9/_1_ ;
 wire net691;
 wire net692;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;

 sg13g2_tiehi \not9/_0__101  (.L_HI(net693));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tielo \flop10/_4__6  (.L_LO(net6));
 sg13g2_tielo \flop11/_4__7  (.L_LO(net7));
 sg13g2_tielo \flop15/_4__8  (.L_LO(net8));
 sg13g2_tielo \flop16/_4__9  (.L_LO(net9));
 sg13g2_tielo \flop17/_4__10  (.L_LO(net17));
 sg13g2_tielo \flop18/_4__11  (.L_LO(net18));
 sg13g2_tielo \flop19/_4__12  (.L_LO(net19));
 sg13g2_tielo \flop2/_4__13  (.L_LO(net20));
 sg13g2_tielo \flop20/_4__14  (.L_LO(net156));
 sg13g2_tielo \flop21/_4__15  (.L_LO(net187));
 sg13g2_tielo \flop22/_4__16  (.L_LO(net199));
 sg13g2_tielo \flop23/_4__17  (.L_LO(net218));
 sg13g2_tielo \flop24/_4__18  (.L_LO(net406));
 sg13g2_tielo \flop25/_4__19  (.L_LO(net412));
 sg13g2_tielo \flop26/_4__20  (.L_LO(net521));
 sg13g2_tielo \flop3/_4__21  (.L_LO(net526));
 sg13g2_tielo \flop4/_4__22  (.L_LO(net527));
 sg13g2_tielo \flop5/_4__23  (.L_LO(net553));
 sg13g2_tielo \flop6/_4__24  (.L_LO(net586));
 sg13g2_tielo \flop7/_4__25  (.L_LO(net617));
 sg13g2_tielo \flop8/_4__26  (.L_LO(net618));
 sg13g2_tielo \flop9/_4__27  (.L_LO(net619));
 sg13g2_tielo \mux60/_0__28  (.L_LO(net620));
 sg13g2_tielo \mux69/_0__29  (.L_LO(net621));
 sg13g2_tielo \not130/_0__30  (.L_LO(net622));
 sg13g2_tielo tt_um_wokwi_411379488132926465_31 (.L_LO(net623));
 sg13g2_tielo tt_um_wokwi_411379488132926465_32 (.L_LO(net624));
 sg13g2_tielo tt_um_wokwi_411379488132926465_33 (.L_LO(net625));
 sg13g2_tielo tt_um_wokwi_411379488132926465_34 (.L_LO(net626));
 sg13g2_tielo tt_um_wokwi_411379488132926465_35 (.L_LO(net627));
 sg13g2_tielo tt_um_wokwi_411379488132926465_36 (.L_LO(net628));
 sg13g2_tielo tt_um_wokwi_411379488132926465_37 (.L_LO(net629));
 sg13g2_tielo tt_um_wokwi_411379488132926465_38 (.L_LO(net630));
 sg13g2_tielo tt_um_wokwi_411379488132926465_39 (.L_LO(net631));
 sg13g2_tielo tt_um_wokwi_411379488132926465_40 (.L_LO(net632));
 sg13g2_tielo tt_um_wokwi_411379488132926465_41 (.L_LO(net633));
 sg13g2_tielo tt_um_wokwi_411379488132926465_42 (.L_LO(net634));
 sg13g2_tielo tt_um_wokwi_411379488132926465_43 (.L_LO(net635));
 sg13g2_tielo tt_um_wokwi_411379488132926465_44 (.L_LO(net636));
 sg13g2_tielo tt_um_wokwi_411379488132926465_45 (.L_LO(net637));
 sg13g2_tielo tt_um_wokwi_411379488132926465_46 (.L_LO(net638));
 sg13g2_tielo tt_um_wokwi_411379488132926465_47 (.L_LO(net639));
 sg13g2_tielo \flop1/dffsr_48  (.L_LO(net640));
 sg13g2_buf_1 _73_ (.A(net10),
    .X(uo_out[0]));
 sg13g2_buf_1 _74_ (.A(net11),
    .X(uo_out[1]));
 sg13g2_buf_1 _75_ (.A(net12),
    .X(uo_out[2]));
 sg13g2_buf_1 _76_ (.A(net13),
    .X(uo_out[3]));
 sg13g2_buf_1 _77_ (.A(net14),
    .X(uo_out[4]));
 sg13g2_buf_1 _78_ (.A(net15),
    .X(uo_out[5]));
 sg13g2_buf_1 _79_ (.A(net16),
    .X(uo_out[6]));
 sg13g2_and2_1 \and1/_0_  (.A(net2),
    .B(net749),
    .X(net136));
 sg13g2_and2_1 \and10/_0_  (.A(net725),
    .B(net159),
    .X(net163));
 sg13g2_and2_1 \and100/_0_  (.A(net388),
    .B(net389),
    .X(net387));
 sg13g2_and2_1 \and101/_0_  (.A(net390),
    .B(net718),
    .X(net391));
 sg13g2_and2_1 \and102/_0_  (.A(net395),
    .B(net718),
    .X(net394));
 sg13g2_and2_1 \and103/_0_  (.A(net397),
    .B(net396),
    .X(net393));
 sg13g2_and2_1 \and104/_0_  (.A(net718),
    .B(net398),
    .X(net399));
 sg13g2_and2_1 \and105/_0_  (.A(net402),
    .B(net718),
    .X(net400));
 sg13g2_and2_1 \and106/_0_  (.A(net721),
    .B(net404),
    .X(net403));
 sg13g2_and2_1 \and107/_0_  (.A(net419),
    .B(net416),
    .X(net423));
 sg13g2_and2_1 \and108/_0_  (.A(net422),
    .B(net416),
    .X(net426));
 sg13g2_and2_1 \and109/_0_  (.A(net420),
    .B(net418),
    .X(net427));
 sg13g2_and2_1 \and11/_0_  (.A(net158),
    .B(net161),
    .X(net164));
 sg13g2_and2_1 \and110/_0_  (.A(net422),
    .B(net418),
    .X(net428));
 sg13g2_and2_1 \and111/_0_  (.A(net421),
    .B(net416),
    .X(net429));
 sg13g2_and2_1 \and112/_0_  (.A(net419),
    .B(net418),
    .X(net430));
 sg13g2_and2_1 \and113/_0_  (.A(net422),
    .B(net421),
    .X(net431));
 sg13g2_and2_1 \and114/_0_  (.A(net429),
    .B(net419),
    .X(net432));
 sg13g2_and2_1 \and115/_0_  (.A(net422),
    .B(net420),
    .X(net424));
 sg13g2_and2_1 \and116/_0_  (.A(net446),
    .B(net448),
    .X(net450));
 sg13g2_and2_1 \and117/_0_  (.A(net447),
    .B(net720),
    .X(net451));
 sg13g2_and2_1 \and118/_0_  (.A(net444),
    .B(net448),
    .X(net454));
 sg13g2_and2_1 \and119/_0_  (.A(net445),
    .B(net720),
    .X(net456));
 sg13g2_and2_1 \and12/_0_  (.A(net158),
    .B(net159),
    .X(net165));
 sg13g2_and2_1 \and120/_0_  (.A(net447),
    .B(net444),
    .X(net460));
 sg13g2_and2_1 \and121/_0_  (.A(net444),
    .B(net720),
    .X(net461));
 sg13g2_and2_1 \and122/_0_  (.A(net447),
    .B(net449),
    .X(net463));
 sg13g2_and2_1 \and123/_0_  (.A(net446),
    .B(net448),
    .X(net464));
 sg13g2_and2_1 \and124/_0_  (.A(net445),
    .B(net464),
    .X(net465));
 sg13g2_and2_1 \and125/_0_  (.A(net444),
    .B(net720),
    .X(net468));
 sg13g2_and2_1 \and126/_0_  (.A(net447),
    .B(net720),
    .X(net469));
 sg13g2_and2_1 \and127/_0_  (.A(net445),
    .B(net446),
    .X(net471));
 sg13g2_and2_1 \and128/_0_  (.A(net446),
    .B(net720),
    .X(net472));
 sg13g2_and2_1 \and129/_0_  (.A(net445),
    .B(net720),
    .X(net474));
 sg13g2_and2_1 \and13/_0_  (.A(net158),
    .B(net160),
    .X(net166));
 sg13g2_and2_1 \and130/_0_  (.A(net445),
    .B(net446),
    .X(net476));
 sg13g2_and2_1 \and131/_0_  (.A(net446),
    .B(net720),
    .X(net477));
 sg13g2_and2_1 \and132/_0_  (.A(net444),
    .B(net447),
    .X(net479));
 sg13g2_and2_1 \and133/_0_  (.A(net489),
    .B(net487),
    .X(net490));
 sg13g2_and2_1 \and134/_0_  (.A(net488),
    .B(net486),
    .X(net491));
 sg13g2_and2_1 \and135/_0_  (.A(net484),
    .B(net487),
    .X(net492));
 sg13g2_and2_1 \and136/_0_  (.A(net485),
    .B(net493),
    .X(net494));
 sg13g2_and2_1 \and137/_0_  (.A(net488),
    .B(net486),
    .X(net493));
 sg13g2_and2_1 \and138/_0_  (.A(net489),
    .B(net484),
    .X(net495));
 sg13g2_and2_1 \and139/_0_  (.A(net489),
    .B(net485),
    .X(net496));
 sg13g2_and2_1 \and14/_0_  (.A(net158),
    .B(net162),
    .X(net167));
 sg13g2_and2_1 \and140/_0_  (.A(net488),
    .B(net484),
    .X(net497));
 sg13g2_and2_1 \and141/_0_  (.A(net489),
    .B(net486),
    .X(net498));
 sg13g2_and2_1 \and142/_0_  (.A(net485),
    .B(net486),
    .X(net499));
 sg13g2_and2_1 \and143/_0_  (.A(net557),
    .B(net529),
    .X(net558));
 sg13g2_and2_1 \and144/_0_  (.A(net560),
    .B(net559),
    .X(net561));
 sg13g2_and2_1 \and145/_0_  (.A(net562),
    .B(net537),
    .X(net563));
 sg13g2_and2_1 \and146/_0_  (.A(net565),
    .B(net564),
    .X(net566));
 sg13g2_and2_1 \and147/_0_  (.A(net561),
    .B(net558),
    .X(net567));
 sg13g2_and2_1 \and148/_0_  (.A(net566),
    .B(net563),
    .X(net568));
 sg13g2_and2_1 \and149/_0_  (.A(net568),
    .B(net567),
    .X(net544));
 sg13g2_and2_1 \and15/_0_  (.A(net725),
    .B(net161),
    .X(net168));
 sg13g2_and2_1 \and150/_0_  (.A(net571),
    .B(net570),
    .X(net572));
 sg13g2_and2_1 \and151/_0_  (.A(net539),
    .B(net537),
    .X(net573));
 sg13g2_and2_1 \and152/_0_  (.A(net531),
    .B(net574),
    .X(net575));
 sg13g2_and2_1 \and153/_0_  (.A(net543),
    .B(net569),
    .X(net576));
 sg13g2_and2_1 \and154/_0_  (.A(net572),
    .B(net575),
    .X(net577));
 sg13g2_and2_1 \and155/_0_  (.A(net578),
    .B(net577),
    .X(net546));
 sg13g2_and2_1 \and156/_0_  (.A(net576),
    .B(net573),
    .X(net578));
 sg13g2_and2_1 \and157/_0_  (.A(net531),
    .B(net529),
    .X(net579));
 sg13g2_and2_1 \and158/_0_  (.A(net535),
    .B(net533),
    .X(net580));
 sg13g2_and2_1 \and159/_0_  (.A(net539),
    .B(net537),
    .X(net581));
 sg13g2_and2_1 \and16/_0_  (.A(net162),
    .B(net159),
    .X(net169));
 sg13g2_and2_1 \and160/_0_  (.A(net582),
    .B(net541),
    .X(net583));
 sg13g2_and2_1 \and161/_0_  (.A(net580),
    .B(net579),
    .X(net584));
 sg13g2_and2_1 \and162/_0_  (.A(net583),
    .B(net581),
    .X(net585));
 sg13g2_and2_1 \and163/_0_  (.A(net585),
    .B(net584),
    .X(net549));
 sg13g2_and2_1 \and164/_0_  (.A(net535),
    .B(net529),
    .X(net587));
 sg13g2_and2_1 \and165/_0_  (.A(net589),
    .B(net588),
    .X(net590));
 sg13g2_and2_1 \and166/_0_  (.A(net592),
    .B(net591),
    .X(net593));
 sg13g2_and2_1 \and167/_0_  (.A(net594),
    .B(net541),
    .X(net595));
 sg13g2_and2_1 \and168/_0_  (.A(net593),
    .B(net595),
    .X(net596));
 sg13g2_and2_1 \and169/_0_  (.A(net590),
    .B(net587),
    .X(net597));
 sg13g2_and2_1 \and17/_0_  (.A(net161),
    .B(net160),
    .X(net170));
 sg13g2_and2_1 \and170/_0_  (.A(net597),
    .B(net596),
    .X(net550));
 sg13g2_and2_1 \and171/_0_  (.A(net533),
    .B(net529),
    .X(net598));
 sg13g2_and2_1 \and172/_0_  (.A(net600),
    .B(net599),
    .X(net601));
 sg13g2_and2_1 \and173/_0_  (.A(net541),
    .B(net537),
    .X(net602));
 sg13g2_and2_1 \and174/_0_  (.A(net604),
    .B(net603),
    .X(net605));
 sg13g2_and2_1 \and175/_0_  (.A(net601),
    .B(net598),
    .X(net606));
 sg13g2_and2_1 \and176/_0_  (.A(net605),
    .B(net602),
    .X(net607));
 sg13g2_and2_1 \and177/_0_  (.A(net607),
    .B(net606),
    .X(net552));
 sg13g2_and2_1 \and178/_0_  (.A(net532),
    .B(net530),
    .X(net608));
 sg13g2_and2_1 \and179/_0_  (.A(net536),
    .B(net534),
    .X(net609));
 sg13g2_and2_1 \and18/_0_  (.A(net162),
    .B(net159),
    .X(net171));
 sg13g2_and2_1 \and180/_0_  (.A(net540),
    .B(net538),
    .X(net610));
 sg13g2_and2_1 \and181/_0_  (.A(net543),
    .B(net542),
    .X(net611));
 sg13g2_and2_1 \and182/_0_  (.A(net609),
    .B(net608),
    .X(net612));
 sg13g2_and2_1 \and183/_0_  (.A(net611),
    .B(net610),
    .X(net613));
 sg13g2_and2_1 \and184/_0_  (.A(net613),
    .B(net612),
    .X(net614));
 sg13g2_and2_1 \and19/_0_  (.A(net181),
    .B(net158),
    .X(net95));
 sg13g2_and2_1 \and2/_0_  (.A(net135),
    .B(net749),
    .X(net139));
 sg13g2_and2_1 \and20/_0_  (.A(net725),
    .B(net171),
    .X(net180));
 sg13g2_and2_1 \and21/_0_  (.A(net157),
    .B(net191),
    .X(net196));
 sg13g2_and2_1 \and22/_0_  (.A(net195),
    .B(net174),
    .X(net197));
 sg13g2_and2_1 \and23/_0_  (.A(net197),
    .B(net196),
    .X(net198));
 sg13g2_and2_1 \and24/_0_  (.A(net692),
    .B(net189),
    .X(net200));
 sg13g2_and2_1 \and25/_0_  (.A(net157),
    .B(net203),
    .X(net201));
 sg13g2_and2_1 \and26/_0_  (.A(net202),
    .B(net204),
    .X(net186));
 sg13g2_and2_1 \and27/_0_  (.A(net725),
    .B(net191),
    .X(net205));
 sg13g2_and2_1 \and28/_0_  (.A(net161),
    .B(net206),
    .X(net207));
 sg13g2_and2_1 \and29/_0_  (.A(net211),
    .B(net195),
    .X(net209));
 sg13g2_and2_1 \and3/_0_  (.A(net133),
    .B(net740),
    .X(net140));
 sg13g2_and2_1 \and30/_0_  (.A(net159),
    .B(net212),
    .X(net210));
 sg13g2_and2_1 \and31/_0_  (.A(net161),
    .B(net725),
    .X(net211));
 sg13g2_and2_1 \and32/_0_  (.A(net216),
    .B(net193),
    .X(net213));
 sg13g2_and2_1 \and33/_0_  (.A(net174),
    .B(net217),
    .X(net214));
 sg13g2_and2_1 \and34/_0_  (.A(net211),
    .B(net159),
    .X(net216));
 sg13g2_and2_1 \and35/_0_  (.A(net204),
    .B(net215),
    .X(net192));
 sg13g2_and2_1 \and36/_0_  (.A(net204),
    .B(net208),
    .X(net190));
 sg13g2_and2_1 \and37/_0_  (.A(net220),
    .B(net219),
    .X(net221));
 sg13g2_and2_1 \and38/_0_  (.A(net739),
    .B(net757),
    .X(net222));
 sg13g2_and2_1 \and39/_0_  (.A(net225),
    .B(net224),
    .X(net226));
 sg13g2_and2_1 \and4/_0_  (.A(net135),
    .B(net740),
    .X(net141));
 sg13g2_and2_1 \and40/_0_  (.A(net735),
    .B(net745),
    .X(net227));
 sg13g2_and2_1 \and41/_0_  (.A(net233),
    .B(net232),
    .X(net234));
 sg13g2_and2_1 \and42/_0_  (.A(net748),
    .B(net232),
    .X(net235));
 sg13g2_and2_1 \and43/_0_  (.A(net739),
    .B(net236),
    .X(net237));
 sg13g2_and2_1 \and44/_0_  (.A(net238),
    .B(net747),
    .X(net239));
 sg13g2_and2_1 \and45/_0_  (.A(net242),
    .B(net753),
    .X(net236));
 sg13g2_and2_1 \and46/_0_  (.A(net244),
    .B(net243),
    .X(net245));
 sg13g2_and2_1 \and47/_0_  (.A(net246),
    .B(net744),
    .X(net247));
 sg13g2_and2_1 \and48/_0_  (.A(net249),
    .B(net248),
    .X(net250));
 sg13g2_and2_1 \and49/_0_  (.A(net251),
    .B(net755),
    .X(net252));
 sg13g2_and2_1 \and5/_0_  (.A(net134),
    .B(net749),
    .X(net142));
 sg13g2_and2_1 \and50/_0_  (.A(net253),
    .B(net755),
    .X(net254));
 sg13g2_and2_1 \and51/_0_  (.A(net743),
    .B(net256),
    .X(net257));
 sg13g2_and2_1 \and52/_0_  (.A(net258),
    .B(net752),
    .X(net259));
 sg13g2_and2_1 \and53/_0_  (.A(net260),
    .B(net744),
    .X(net261));
 sg13g2_and2_1 \and54/_0_  (.A(net264),
    .B(net263),
    .X(net265));
 sg13g2_and2_1 \and55/_0_  (.A(net740),
    .B(net757),
    .X(net267));
 sg13g2_and2_1 \and56/_0_  (.A(net735),
    .B(net745),
    .X(net269));
 sg13g2_and2_1 \and57/_0_  (.A(net273),
    .B(net272),
    .X(net271));
 sg13g2_and2_1 \and58/_0_  (.A(net283),
    .B(net282),
    .X(net276));
 sg13g2_and2_1 \and59/_0_  (.A(net747),
    .B(net284),
    .X(net277));
 sg13g2_and2_1 \and6/_0_  (.A(net2),
    .B(net740),
    .X(net143));
 sg13g2_and2_1 \and60/_0_  (.A(net287),
    .B(net757),
    .X(net280));
 sg13g2_and2_1 \and61/_0_  (.A(net288),
    .B(net747),
    .X(net279));
 sg13g2_and2_1 \and62/_0_  (.A(net738),
    .B(net285),
    .X(net287));
 sg13g2_and2_1 \and63/_0_  (.A(net291),
    .B(net286),
    .X(net289));
 sg13g2_and2_1 \and64/_0_  (.A(net292),
    .B(net745),
    .X(net290));
 sg13g2_and2_1 \and65/_0_  (.A(net298),
    .B(net297),
    .X(net295));
 sg13g2_and2_1 \and66/_0_  (.A(net299),
    .B(net755),
    .X(net296));
 sg13g2_and2_1 \and67/_0_  (.A(net300),
    .B(net755),
    .X(net294));
 sg13g2_and2_1 \and68/_0_  (.A(net305),
    .B(net752),
    .X(net302));
 sg13g2_and2_1 \and69/_0_  (.A(net306),
    .B(net744),
    .X(net304));
 sg13g2_and2_1 \and7/_0_  (.A(net135),
    .B(net134),
    .X(net144));
 sg13g2_and2_1 \and70/_0_  (.A(net743),
    .B(net307),
    .X(net303));
 sg13g2_and2_1 \and71/_0_  (.A(net308),
    .B(net751),
    .X(net309));
 sg13g2_and2_1 \and72/_0_  (.A(net313),
    .B(net752),
    .X(net312));
 sg13g2_and2_1 \and73/_0_  (.A(net315),
    .B(net314),
    .X(net311));
 sg13g2_and2_1 \and74/_0_  (.A(net751),
    .B(net316),
    .X(net317));
 sg13g2_and2_1 \and75/_0_  (.A(net320),
    .B(net751),
    .X(net318));
 sg13g2_and2_1 \and76/_0_  (.A(net743),
    .B(net322),
    .X(net321));
 sg13g2_and2_1 \and77/_0_  (.A(net746),
    .B(net323),
    .X(net324));
 sg13g2_and2_1 \and78/_0_  (.A(net326),
    .B(net327),
    .X(net325));
 sg13g2_and2_1 \and79/_0_  (.A(net330),
    .B(net331),
    .X(net332));
 sg13g2_and2_1 \and8/_0_  (.A(net142),
    .B(net2),
    .X(net145));
 sg13g2_and2_1 \and80/_0_  (.A(net747),
    .B(net335),
    .X(net333));
 sg13g2_and2_1 \and81/_0_  (.A(net748),
    .B(net336),
    .X(net337));
 sg13g2_and2_1 \and82/_0_  (.A(net738),
    .B(net753),
    .X(net338));
 sg13g2_and2_1 \and83/_0_  (.A(net339),
    .B(net338),
    .X(net340));
 sg13g2_and2_1 \and84/_0_  (.A(net347),
    .B(net345),
    .X(net342));
 sg13g2_and2_1 \and85/_0_  (.A(net747),
    .B(net346),
    .X(net343));
 sg13g2_and2_1 \and86/_0_  (.A(net738),
    .B(net754),
    .X(net348));
 sg13g2_and2_1 \and87/_0_  (.A(net351),
    .B(net350),
    .X(net352));
 sg13g2_and2_1 \and88/_0_  (.A(net735),
    .B(net746),
    .X(net354));
 sg13g2_and2_1 \and89/_0_  (.A(net359),
    .B(net361),
    .X(net355));
 sg13g2_and2_1 \and9/_0_  (.A(net135),
    .B(net133),
    .X(net137));
 sg13g2_and2_1 \and90/_0_  (.A(net722),
    .B(net362),
    .X(net356));
 sg13g2_and2_1 \and91/_0_  (.A(net724),
    .B(net719),
    .X(net364));
 sg13g2_and2_1 \and92/_0_  (.A(net367),
    .B(net366),
    .X(net368));
 sg13g2_and2_1 \and93/_0_  (.A(net723),
    .B(net721),
    .X(net370));
 sg13g2_and2_1 \and94/_0_  (.A(net373),
    .B(net374),
    .X(net375));
 sg13g2_and2_1 \and95/_0_  (.A(net722),
    .B(net378),
    .X(net376));
 sg13g2_and2_1 \and96/_0_  (.A(net722),
    .B(net379),
    .X(net380));
 sg13g2_and2_1 \and97/_0_  (.A(net724),
    .B(net719),
    .X(net381));
 sg13g2_and2_1 \and98/_0_  (.A(net382),
    .B(net381),
    .X(net383));
 sg13g2_and2_1 \and99/_0_  (.A(net721),
    .B(net385),
    .X(net386));
 sg13g2_inv_1 \flop1/_4_  (.Y(\flop1/_1_ ),
    .A(net5));
 sg13g2_inv_1 \flop1/_5_  (.Y(\flop1/_0_ ),
    .A(net188));
 sg13g2_tielo \flop1/dffsr_49  (.L_LO(net641));
 sg13g2_tielo \flop10/dffsr_50  (.L_LO(net642));
 sg13g2_sdfbbp_1 \flop1/dffsr  (.Q(net157),
    .Q_N(net189),
    .RESET_B(\flop1/_0_ ),
    .SET_B(\flop1/_1_ ),
    .D(net186),
    .SCE(net641),
    .SCD(net640),
    .CLK(net757));
 sg13g2_inv_1 \flop10/_4_  (.Y(\flop10/_1_ ),
    .A(net6));
 sg13g2_inv_1 \flop10/_5_  (.Y(\flop10/_0_ ),
    .A(net413));
 sg13g2_tielo \flop10/dffsr_51  (.L_LO(net643));
 sg13g2_tielo \flop11/dffsr_52  (.L_LO(net644));
 sg13g2_sdfbbp_1 \flop10/dffsr  (.Q(net418),
    .Q_N(net415),
    .RESET_B(\flop10/_0_ ),
    .SET_B(\flop10/_1_ ),
    .D(net415),
    .SCE(net643),
    .SCD(net642),
    .CLK(net417));
 sg13g2_inv_1 \flop11/_4_  (.Y(\flop11/_1_ ),
    .A(net7));
 sg13g2_inv_1 \flop11/_5_  (.Y(\flop11/_0_ ),
    .A(net413));
 sg13g2_tielo \flop11/dffsr_53  (.L_LO(net645));
 sg13g2_tielo \flop12/dffsr_54  (.L_LO(net646));
 sg13g2_sdfbbp_1 \flop11/dffsr  (.Q(net419),
    .Q_N(net417),
    .RESET_B(\flop11/_0_ ),
    .SET_B(\flop11/_1_ ),
    .D(net417),
    .SCE(net645),
    .SCD(net644),
    .CLK(net751));
 sg13g2_inv_1 \flop12/_4_  (.Y(\flop12/_1_ ),
    .A(net751));
 sg13g2_inv_1 \flop12/_5_  (.Y(\flop12/_0_ ),
    .A(net443));
 sg13g2_tielo \flop12/dffsr_55  (.L_LO(net647));
 sg13g2_tielo \flop13/dffsr_56  (.L_LO(net648));
 sg13g2_sdfbbp_1 \flop12/dffsr  (.Q(net448),
    .Q_N(net481),
    .RESET_B(\flop12/_0_ ),
    .SET_B(\flop12/_1_ ),
    .D(net481),
    .SCE(net647),
    .SCD(net646),
    .CLK(net743));
 sg13g2_inv_1 \flop13/_4_  (.Y(\flop13/_1_ ),
    .A(net751));
 sg13g2_inv_1 \flop13/_5_  (.Y(\flop13/_0_ ),
    .A(net443));
 sg13g2_tielo \flop13/dffsr_57  (.L_LO(net649));
 sg13g2_tielo \flop14/dffsr_58  (.L_LO(net650));
 sg13g2_sdfbbp_1 \flop13/dffsr  (.Q(net446),
    .Q_N(net482),
    .RESET_B(\flop13/_0_ ),
    .SET_B(\flop13/_1_ ),
    .D(net482),
    .SCE(net649),
    .SCD(net648),
    .CLK(net483));
 sg13g2_inv_1 \flop14/_4_  (.Y(\flop14/_1_ ),
    .A(net751));
 sg13g2_inv_1 \flop14/_5_  (.Y(\flop14/_0_ ),
    .A(net443));
 sg13g2_tielo \flop14/dffsr_59  (.L_LO(net651));
 sg13g2_tielo \flop15/dffsr_60  (.L_LO(net652));
 sg13g2_sdfbbp_1 \flop14/dffsr  (.Q(net444),
    .Q_N(net483),
    .RESET_B(\flop14/_0_ ),
    .SET_B(\flop14/_1_ ),
    .D(net483),
    .SCE(net651),
    .SCD(net650),
    .CLK(net481));
 sg13g2_inv_1 \flop15/_4_  (.Y(\flop15/_1_ ),
    .A(net8));
 sg13g2_inv_1 \flop15/_5_  (.Y(\flop15/_0_ ),
    .A(net520));
 sg13g2_tielo \flop15/dffsr_61  (.L_LO(net653));
 sg13g2_tielo \flop16/dffsr_62  (.L_LO(net654));
 sg13g2_sdfbbp_1 \flop15/dffsr  (.Q(net484),
    .Q_N(net522),
    .RESET_B(\flop15/_0_ ),
    .SET_B(\flop15/_1_ ),
    .D(net522),
    .SCE(net653),
    .SCD(net652),
    .CLK(net523));
 sg13g2_inv_1 \flop16/_4_  (.Y(\flop16/_1_ ),
    .A(net9));
 sg13g2_inv_1 \flop16/_5_  (.Y(\flop16/_0_ ),
    .A(net520));
 sg13g2_tielo \flop16/dffsr_63  (.L_LO(net655));
 sg13g2_tielo \flop17/dffsr_64  (.L_LO(net656));
 sg13g2_sdfbbp_1 \flop16/dffsr  (.Q(net486),
    .Q_N(net524),
    .RESET_B(\flop16/_0_ ),
    .SET_B(\flop16/_1_ ),
    .D(net524),
    .SCE(net655),
    .SCD(net654),
    .CLK(net522));
 sg13g2_inv_1 \flop17/_4_  (.Y(\flop17/_1_ ),
    .A(net17));
 sg13g2_inv_1 \flop17/_5_  (.Y(\flop17/_0_ ),
    .A(net520));
 sg13g2_tielo \flop17/dffsr_65  (.L_LO(net657));
 sg13g2_tielo \flop18/dffsr_66  (.L_LO(net658));
 sg13g2_sdfbbp_1 \flop17/dffsr  (.Q(net488),
    .Q_N(net523),
    .RESET_B(\flop17/_0_ ),
    .SET_B(\flop17/_1_ ),
    .D(net523),
    .SCE(net657),
    .SCD(net656),
    .CLK(net752));
 sg13g2_inv_1 \flop18/_4_  (.Y(\flop18/_1_ ),
    .A(net18));
 sg13g2_inv_1 \flop18/_5_  (.Y(\flop18/_0_ ),
    .A(net520));
 sg13g2_tielo \flop18/dffsr_67  (.L_LO(net659));
 sg13g2_tielo \flop19/dffsr_68  (.L_LO(net660));
 sg13g2_sdfbbp_1 \flop18/dffsr  (.Q(net515),
    .Q_N(net525),
    .RESET_B(\flop18/_0_ ),
    .SET_B(\flop18/_1_ ),
    .D(net525),
    .SCE(net659),
    .SCD(net658),
    .CLK(net524));
 sg13g2_inv_1 \flop19/_4_  (.Y(\flop19/_1_ ),
    .A(net19));
 sg13g2_inv_1 \flop19/_5_  (.Y(\flop19/_0_ ),
    .A(net528));
 sg13g2_tielo \flop19/dffsr_69  (.L_LO(net661));
 sg13g2_tielo \flop2/dffsr_70  (.L_LO(net662));
 sg13g2_sdfbbp_1 \flop19/dffsr  (.Q(net529),
    .Q_N(net530),
    .RESET_B(\flop19/_0_ ),
    .SET_B(\flop19/_1_ ),
    .D(net752),
    .SCE(net661),
    .SCD(net660),
    .CLK(net742));
 sg13g2_inv_1 \flop2/_4_  (.Y(\flop2/_1_ ),
    .A(net20));
 sg13g2_inv_1 \flop2/_5_  (.Y(\flop2/_0_ ),
    .A(net188));
 sg13g2_tielo \flop2/dffsr_71  (.L_LO(net663));
 sg13g2_tielo \flop20/dffsr_72  (.L_LO(net664));
 sg13g2_sdfbbp_1 \flop2/dffsr  (.Q(net161),
    .Q_N(net191),
    .RESET_B(\flop2/_0_ ),
    .SET_B(\flop2/_1_ ),
    .D(net190),
    .SCE(net663),
    .SCD(net662),
    .CLK(net757));
 sg13g2_inv_1 \flop20/_4_  (.Y(\flop20/_1_ ),
    .A(net156));
 sg13g2_inv_1 \flop20/_5_  (.Y(\flop20/_0_ ),
    .A(net528));
 sg13g2_tielo \flop20/dffsr_73  (.L_LO(net665));
 sg13g2_tielo \flop21/dffsr_74  (.L_LO(net666));
 sg13g2_sdfbbp_1 \flop20/dffsr  (.Q(net531),
    .Q_N(net532),
    .RESET_B(\flop20/_0_ ),
    .SET_B(\flop20/_1_ ),
    .D(net529),
    .SCE(net665),
    .SCD(net664),
    .CLK(net742));
 sg13g2_inv_1 \flop21/_4_  (.Y(\flop21/_1_ ),
    .A(net187));
 sg13g2_inv_1 \flop21/_5_  (.Y(\flop21/_0_ ),
    .A(net528));
 sg13g2_tielo \flop21/dffsr_75  (.L_LO(net667));
 sg13g2_tielo \flop22/dffsr_76  (.L_LO(net668));
 sg13g2_sdfbbp_1 \flop21/dffsr  (.Q(net533),
    .Q_N(net534),
    .RESET_B(\flop21/_0_ ),
    .SET_B(\flop21/_1_ ),
    .D(net531),
    .SCE(net667),
    .SCD(net666),
    .CLK(net742));
 sg13g2_inv_1 \flop22/_4_  (.Y(\flop22/_1_ ),
    .A(net199));
 sg13g2_inv_1 \flop22/_5_  (.Y(\flop22/_0_ ),
    .A(net528));
 sg13g2_tielo \flop22/dffsr_77  (.L_LO(net669));
 sg13g2_tielo \flop23/dffsr_78  (.L_LO(net670));
 sg13g2_sdfbbp_1 \flop22/dffsr  (.Q(net535),
    .Q_N(net536),
    .RESET_B(\flop22/_0_ ),
    .SET_B(\flop22/_1_ ),
    .D(net533),
    .SCE(net669),
    .SCD(net668),
    .CLK(net742));
 sg13g2_inv_1 \flop23/_4_  (.Y(\flop23/_1_ ),
    .A(net218));
 sg13g2_inv_1 \flop23/_5_  (.Y(\flop23/_0_ ),
    .A(net528));
 sg13g2_tielo \flop23/dffsr_79  (.L_LO(net671));
 sg13g2_tielo \flop24/dffsr_80  (.L_LO(net672));
 sg13g2_sdfbbp_1 \flop23/dffsr  (.Q(net537),
    .Q_N(net538),
    .RESET_B(\flop23/_0_ ),
    .SET_B(\flop23/_1_ ),
    .D(net535),
    .SCE(net671),
    .SCD(net670),
    .CLK(net742));
 sg13g2_inv_1 \flop24/_4_  (.Y(\flop24/_1_ ),
    .A(net406));
 sg13g2_inv_1 \flop24/_5_  (.Y(\flop24/_0_ ),
    .A(net528));
 sg13g2_tielo \flop24/dffsr_81  (.L_LO(net673));
 sg13g2_tielo \flop25/dffsr_82  (.L_LO(net674));
 sg13g2_sdfbbp_1 \flop24/dffsr  (.Q(net539),
    .Q_N(net540),
    .RESET_B(\flop24/_0_ ),
    .SET_B(\flop24/_1_ ),
    .D(net537),
    .SCE(net673),
    .SCD(net672),
    .CLK(net742));
 sg13g2_inv_1 \flop25/_4_  (.Y(\flop25/_1_ ),
    .A(net412));
 sg13g2_inv_1 \flop25/_5_  (.Y(\flop25/_0_ ),
    .A(net528));
 sg13g2_tielo \flop25/dffsr_83  (.L_LO(net675));
 sg13g2_tielo \flop26/dffsr_84  (.L_LO(net676));
 sg13g2_sdfbbp_1 \flop25/dffsr  (.Q(net541),
    .Q_N(net542),
    .RESET_B(\flop25/_0_ ),
    .SET_B(\flop25/_1_ ),
    .D(net539),
    .SCE(net675),
    .SCD(net674),
    .CLK(net742));
 sg13g2_inv_1 \flop26/_4_  (.Y(\flop26/_1_ ),
    .A(net521));
 sg13g2_inv_1 \flop26/_5_  (.Y(\flop26/_0_ ),
    .A(net528));
 sg13g2_tielo \flop26/dffsr_85  (.L_LO(net677));
 sg13g2_tielo \flop3/dffsr_86  (.L_LO(net678));
 sg13g2_sdfbbp_1 \flop26/dffsr  (.Q(net543),
    .Q_N(\flop26/notq ),
    .RESET_B(\flop26/_0_ ),
    .SET_B(\flop26/_1_ ),
    .D(net541),
    .SCE(net677),
    .SCD(net676),
    .CLK(net742));
 sg13g2_inv_1 \flop3/_4_  (.Y(\flop3/_1_ ),
    .A(net526));
 sg13g2_inv_1 \flop3/_5_  (.Y(\flop3/_0_ ),
    .A(net188));
 sg13g2_tielo \flop3/dffsr_87  (.L_LO(net679));
 sg13g2_tielo \flop4/dffsr_88  (.L_LO(net680));
 sg13g2_sdfbbp_1 \flop3/dffsr  (.Q(net174),
    .Q_N(net193),
    .RESET_B(\flop3/_0_ ),
    .SET_B(\flop3/_1_ ),
    .D(net192),
    .SCE(net679),
    .SCD(net678),
    .CLK(net758));
 sg13g2_inv_1 \flop4/_4_  (.Y(\flop4/_1_ ),
    .A(net527));
 sg13g2_inv_1 \flop4/_5_  (.Y(\flop4/_0_ ),
    .A(net188));
 sg13g2_tielo \flop4/dffsr_89  (.L_LO(net681));
 sg13g2_tielo \flop5/dffsr_90  (.L_LO(net682));
 sg13g2_sdfbbp_1 \flop4/dffsr  (.Q(net159),
    .Q_N(net195),
    .RESET_B(\flop4/_0_ ),
    .SET_B(\flop4/_1_ ),
    .D(net194),
    .SCE(net681),
    .SCD(net680),
    .CLK(net757));
 sg13g2_inv_1 \flop5/_4_  (.Y(\flop5/_1_ ),
    .A(net553));
 sg13g2_inv_1 \flop5/_5_  (.Y(\flop5/_0_ ),
    .A(net407));
 sg13g2_tielo \flop5/dffsr_91  (.L_LO(net683));
 sg13g2_tielo \flop6/dffsr_92  (.L_LO(net684));
 sg13g2_sdfbbp_1 \flop5/dffsr  (.Q(net358),
    .Q_N(net405),
    .RESET_B(\flop5/_0_ ),
    .SET_B(\flop5/_1_ ),
    .D(net405),
    .SCE(net683),
    .SCD(net682),
    .CLK(net754));
 sg13g2_inv_1 \flop6/_4_  (.Y(\flop6/_1_ ),
    .A(net586));
 sg13g2_inv_1 \flop6/_5_  (.Y(\flop6/_0_ ),
    .A(net407));
 sg13g2_tielo \flop6/dffsr_93  (.L_LO(net685));
 sg13g2_tielo \flop7/dffsr_94  (.L_LO(net686));
 sg13g2_sdfbbp_1 \flop6/dffsr  (.Q(net363),
    .Q_N(net408),
    .RESET_B(\flop6/_0_ ),
    .SET_B(\flop6/_1_ ),
    .D(net408),
    .SCE(net685),
    .SCD(net684),
    .CLK(net405));
 sg13g2_inv_1 \flop7/_4_  (.Y(\flop7/_1_ ),
    .A(net617));
 sg13g2_inv_1 \flop7/_5_  (.Y(\flop7/_0_ ),
    .A(net407));
 sg13g2_tielo \flop7/dffsr_95  (.L_LO(net687));
 sg13g2_tielo \flop8/dffsr_96  (.L_LO(net688));
 sg13g2_sdfbbp_1 \flop7/dffsr  (.Q(net360),
    .Q_N(net409),
    .RESET_B(\flop7/_0_ ),
    .SET_B(\flop7/_1_ ),
    .D(net409),
    .SCE(net687),
    .SCD(net686),
    .CLK(net408));
 sg13g2_inv_1 \flop8/_4_  (.Y(\flop8/_1_ ),
    .A(net618));
 sg13g2_inv_1 \flop8/_5_  (.Y(\flop8/_0_ ),
    .A(net413));
 sg13g2_tielo \flop8/dffsr_97  (.L_LO(net689));
 sg13g2_tielo \flop9/dffsr_98  (.L_LO(net690));
 sg13g2_sdfbbp_1 \flop8/dffsr  (.Q(net414),
    .Q_N(net410),
    .RESET_B(\flop8/_0_ ),
    .SET_B(\flop8/_1_ ),
    .D(net410),
    .SCE(net689),
    .SCD(net688),
    .CLK(net411));
 sg13g2_inv_1 \flop9/_4_  (.Y(\flop9/_1_ ),
    .A(net619));
 sg13g2_inv_1 \flop9/_5_  (.Y(\flop9/_0_ ),
    .A(net413));
 sg13g2_tielo \flop9/dffsr_99  (.L_LO(net691));
 sg13g2_tiehi \and24/_0__100  (.L_HI(net692));
 sg13g2_sdfbbp_1 \flop9/dffsr  (.Q(net416),
    .Q_N(net411),
    .RESET_B(\flop9/_0_ ),
    .SET_B(\flop9/_1_ ),
    .D(net411),
    .SCE(net691),
    .SCD(net690),
    .CLK(net415));
 sg13g2_mux2_1 \mux1/_0_  (.A0(net21),
    .A1(net22),
    .S(net732),
    .X(net23));
 sg13g2_mux2_1 \mux10/_0_  (.A0(net40),
    .A1(net41),
    .S(net732),
    .X(net42));
 sg13g2_mux2_1 \mux11/_0_  (.A0(net43),
    .A1(net44),
    .S(net733),
    .X(net45));
 sg13g2_mux2_1 \mux12/_0_  (.A0(net46),
    .A1(net47),
    .S(net733),
    .X(net48));
 sg13g2_mux2_1 \mux13/_0_  (.A0(net42),
    .A1(net39),
    .S(net728),
    .X(net49));
 sg13g2_mux2_1 \mux14/_0_  (.A0(net48),
    .A1(net45),
    .S(net729),
    .X(net50));
 sg13g2_mux2_1 \mux15/_0_  (.A0(net50),
    .A1(net49),
    .S(net3),
    .X(net51));
 sg13g2_mux2_1 \mux16/_0_  (.A0(net51),
    .A1(net52),
    .S(net4),
    .X(net11));
 sg13g2_mux2_1 \mux17/_0_  (.A0(net53),
    .A1(net54),
    .S(net731),
    .X(net55));
 sg13g2_mux2_1 \mux18/_0_  (.A0(net56),
    .A1(net57),
    .S(net732),
    .X(net58));
 sg13g2_mux2_1 \mux19/_0_  (.A0(net59),
    .A1(net60),
    .S(net733),
    .X(net61));
 sg13g2_mux2_1 \mux2/_0_  (.A0(net24),
    .A1(net25),
    .S(net734),
    .X(net26));
 sg13g2_mux2_1 \mux20/_0_  (.A0(net62),
    .A1(net63),
    .S(net734),
    .X(net64));
 sg13g2_mux2_1 \mux21/_0_  (.A0(net58),
    .A1(net55),
    .S(net726),
    .X(net65));
 sg13g2_mux2_1 \mux22/_0_  (.A0(net64),
    .A1(net61),
    .S(net729),
    .X(net66));
 sg13g2_mux2_1 \mux23/_0_  (.A0(net66),
    .A1(net65),
    .S(net3),
    .X(net67));
 sg13g2_mux2_1 \mux24/_0_  (.A0(net67),
    .A1(net68),
    .S(net4),
    .X(net12));
 sg13g2_mux2_1 \mux25/_0_  (.A0(net69),
    .A1(net70),
    .S(net732),
    .X(net71));
 sg13g2_mux2_1 \mux26/_0_  (.A0(net72),
    .A1(net73),
    .S(net732),
    .X(net74));
 sg13g2_mux2_1 \mux27/_0_  (.A0(net75),
    .A1(net76),
    .S(net732),
    .X(net77));
 sg13g2_mux2_1 \mux28/_0_  (.A0(net78),
    .A1(net79),
    .S(net734),
    .X(net80));
 sg13g2_mux2_1 \mux29/_0_  (.A0(net74),
    .A1(net71),
    .S(net728),
    .X(net81));
 sg13g2_mux2_1 \mux3/_0_  (.A0(net27),
    .A1(net28),
    .S(net732),
    .X(net29));
 sg13g2_mux2_1 \mux30/_0_  (.A0(net80),
    .A1(net77),
    .S(net728),
    .X(net82));
 sg13g2_mux2_1 \mux31/_0_  (.A0(net82),
    .A1(net81),
    .S(net3),
    .X(net83));
 sg13g2_mux2_1 \mux32/_0_  (.A0(net83),
    .A1(net84),
    .S(net4),
    .X(net13));
 sg13g2_mux2_1 \mux33/_0_  (.A0(net85),
    .A1(net86),
    .S(net730),
    .X(net87));
 sg13g2_mux2_1 \mux34/_0_  (.A0(net88),
    .A1(net89),
    .S(net732),
    .X(net90));
 sg13g2_mux2_1 \mux35/_0_  (.A0(net91),
    .A1(net92),
    .S(net733),
    .X(net93));
 sg13g2_mux2_1 \mux36/_0_  (.A0(net94),
    .A1(net95),
    .S(net733),
    .X(net96));
 sg13g2_mux2_1 \mux37/_0_  (.A0(net90),
    .A1(net87),
    .S(net728),
    .X(net97));
 sg13g2_mux2_1 \mux38/_0_  (.A0(net96),
    .A1(net93),
    .S(net728),
    .X(net98));
 sg13g2_mux2_1 \mux39/_0_  (.A0(net98),
    .A1(net97),
    .S(net3),
    .X(net99));
 sg13g2_mux2_1 \mux4/_0_  (.A0(net30),
    .A1(net31),
    .S(net734),
    .X(net32));
 sg13g2_mux2_1 \mux40/_0_  (.A0(net99),
    .A1(net100),
    .S(net4),
    .X(net14));
 sg13g2_mux2_1 \mux41/_0_  (.A0(net101),
    .A1(net102),
    .S(net730),
    .X(net103));
 sg13g2_mux2_1 \mux42/_0_  (.A0(net104),
    .A1(net105),
    .S(net730),
    .X(net106));
 sg13g2_mux2_1 \mux43/_0_  (.A0(net107),
    .A1(net108),
    .S(net733),
    .X(net109));
 sg13g2_mux2_1 \mux44/_0_  (.A0(net110),
    .A1(net111),
    .S(net733),
    .X(net112));
 sg13g2_mux2_1 \mux45/_0_  (.A0(net106),
    .A1(net103),
    .S(net726),
    .X(net113));
 sg13g2_mux2_1 \mux46/_0_  (.A0(net112),
    .A1(net109),
    .S(net728),
    .X(net114));
 sg13g2_mux2_1 \mux47/_0_  (.A0(net114),
    .A1(net113),
    .S(net3),
    .X(net115));
 sg13g2_mux2_1 \mux48/_0_  (.A0(net115),
    .A1(net116),
    .S(net4),
    .X(net15));
 sg13g2_mux2_1 \mux49/_0_  (.A0(net117),
    .A1(net118),
    .S(net730),
    .X(net119));
 sg13g2_mux2_1 \mux5/_0_  (.A0(net26),
    .A1(net23),
    .S(net728),
    .X(net33));
 sg13g2_mux2_1 \mux50/_0_  (.A0(net120),
    .A1(net121),
    .S(net730),
    .X(net122));
 sg13g2_mux2_1 \mux51/_0_  (.A0(net123),
    .A1(net124),
    .S(net731),
    .X(net125));
 sg13g2_mux2_1 \mux52/_0_  (.A0(net126),
    .A1(net127),
    .S(net733),
    .X(net128));
 sg13g2_mux2_1 \mux53/_0_  (.A0(net122),
    .A1(net119),
    .S(net726),
    .X(net129));
 sg13g2_mux2_1 \mux54/_0_  (.A0(net128),
    .A1(net125),
    .S(net726),
    .X(net130));
 sg13g2_mux2_1 \mux55/_0_  (.A0(net130),
    .A1(net129),
    .S(net3),
    .X(net131));
 sg13g2_mux2_1 \mux56/_0_  (.A0(net131),
    .A1(net132),
    .S(net4),
    .X(net16));
 sg13g2_mux2_1 \mux57/_0_  (.A0(net502),
    .A1(net544),
    .S(net731),
    .X(net545));
 sg13g2_mux2_1 \mux58/_0_  (.A0(net546),
    .A1(net547),
    .S(net731),
    .X(net548));
 sg13g2_mux2_1 \mux59/_0_  (.A0(net549),
    .A1(net550),
    .S(net730),
    .X(net551));
 sg13g2_mux2_1 \mux6/_0_  (.A0(net32),
    .A1(net29),
    .S(net728),
    .X(net34));
 sg13g2_mux2_1 \mux60/_0_  (.A0(net552),
    .A1(net620),
    .S(net730),
    .X(net554));
 sg13g2_mux2_1 \mux61/_0_  (.A0(net545),
    .A1(net548),
    .S(net726),
    .X(net555));
 sg13g2_mux2_1 \mux62/_0_  (.A0(net551),
    .A1(net554),
    .S(net726),
    .X(net556));
 sg13g2_mux2_1 \mux63/_0_  (.A0(net555),
    .A1(net556),
    .S(net3),
    .X(net36));
 sg13g2_mux2_1 \mux64/_0_  (.A0(net514),
    .A1(net615),
    .S(net727),
    .X(net52));
 sg13g2_mux2_1 \mux65/_0_  (.A0(net511),
    .A1(net616),
    .S(net727),
    .X(net68));
 sg13g2_mux2_1 \mux66/_0_  (.A0(net517),
    .A1(net547),
    .S(net727),
    .X(net84));
 sg13g2_mux2_1 \mux67/_0_  (.A0(net509),
    .A1(net547),
    .S(net727),
    .X(net100));
 sg13g2_mux2_1 \mux68/_0_  (.A0(net505),
    .A1(net547),
    .S(net726),
    .X(net116));
 sg13g2_mux2_1 \mux69/_0_  (.A0(net508),
    .A1(net621),
    .S(net726),
    .X(net132));
 sg13g2_mux2_1 \mux7/_0_  (.A0(net34),
    .A1(net33),
    .S(net3),
    .X(net35));
 sg13g2_mux2_1 \mux8/_0_  (.A0(net35),
    .A1(net36),
    .S(net4),
    .X(net10));
 sg13g2_mux2_1 \mux9/_0_  (.A0(net37),
    .A1(net38),
    .S(net730),
    .X(net39));
 sg13g2_nand2_2 \nand1/_0_  (.Y(net547),
    .A(net613),
    .B(net612));
 sg13g2_inv_1 \not1/_0_  (.Y(net133),
    .A(net749));
 sg13g2_inv_1 \not10/_0_  (.Y(net204),
    .A(net198));
 sg13g2_inv_1 \not100/_0_  (.Y(net413),
    .A(net1));
 sg13g2_inv_1 \not101/_0_  (.Y(net420),
    .A(net416));
 sg13g2_inv_1 \not102/_0_  (.Y(net421),
    .A(net418));
 sg13g2_inv_1 \not103/_0_  (.Y(net422),
    .A(net419));
 sg13g2_inv_1 \not104/_0_  (.Y(net443),
    .A(net1));
 sg13g2_inv_1 \not105/_0_  (.Y(net445),
    .A(net444));
 sg13g2_inv_1 \not106/_0_  (.Y(net447),
    .A(net446));
 sg13g2_inv_1 \not107/_0_  (.Y(net449),
    .A(net448));
 sg13g2_inv_1 \not108/_0_  (.Y(net22),
    .A(net453));
 sg13g2_inv_1 \not109/_0_  (.Y(net38),
    .A(net457));
 sg13g2_inv_1 \not11/_0_  (.Y(net206),
    .A(net725));
 sg13g2_inv_1 \not110/_0_  (.Y(net70),
    .A(net467));
 sg13g2_inv_1 \not111/_0_  (.Y(net54),
    .A(net459));
 sg13g2_inv_1 \not112/_0_  (.Y(net118),
    .A(net480));
 sg13g2_inv_1 \not113/_0_  (.Y(net102),
    .A(net475));
 sg13g2_inv_1 \not114/_0_  (.Y(net86),
    .A(net470));
 sg13g2_inv_1 \not115/_0_  (.Y(net485),
    .A(net484));
 sg13g2_inv_1 \not116/_0_  (.Y(net487),
    .A(net486));
 sg13g2_inv_1 \not117/_0_  (.Y(net489),
    .A(net488));
 sg13g2_inv_1 \not118/_0_  (.Y(net520),
    .A(net1));
 sg13g2_inv_2 \not119/_0_  (.Y(net528),
    .A(net1));
 sg13g2_inv_1 \not12/_0_  (.Y(net212),
    .A(net211));
 sg13g2_inv_1 \not120/_0_  (.Y(net557),
    .A(net531));
 sg13g2_inv_1 \not121/_0_  (.Y(net559),
    .A(net533));
 sg13g2_inv_1 \not122/_0_  (.Y(net560),
    .A(net535));
 sg13g2_inv_1 \not123/_0_  (.Y(net562),
    .A(net539));
 sg13g2_inv_1 \not124/_0_  (.Y(net564),
    .A(net541));
 sg13g2_inv_1 \not125/_0_  (.Y(net565),
    .A(net543));
 sg13g2_inv_1 \not126/_0_  (.Y(net569),
    .A(net541));
 sg13g2_inv_1 \not127/_0_  (.Y(net570),
    .A(net533));
 sg13g2_inv_1 \not128/_0_  (.Y(net574),
    .A(net529));
 sg13g2_inv_1 \not129/_0_  (.Y(net571),
    .A(net535));
 sg13g2_inv_1 \not13/_0_  (.Y(net217),
    .A(net216));
 sg13g2_inv_1 \not130/_0_  (.Y(net582),
    .A(net622));
 sg13g2_inv_1 \not131/_0_  (.Y(net588),
    .A(net531));
 sg13g2_inv_1 \not132/_0_  (.Y(net589),
    .A(net533));
 sg13g2_inv_1 \not133/_0_  (.Y(net591),
    .A(net537));
 sg13g2_inv_1 \not134/_0_  (.Y(net592),
    .A(net539));
 sg13g2_inv_1 \not135/_0_  (.Y(net594),
    .A(net543));
 sg13g2_inv_1 \not136/_0_  (.Y(net604),
    .A(net543));
 sg13g2_inv_1 \not137/_0_  (.Y(net603),
    .A(net539));
 sg13g2_inv_1 \not138/_0_  (.Y(net599),
    .A(net531));
 sg13g2_inv_1 \not139/_0_  (.Y(net600),
    .A(net535));
 sg13g2_inv_1 \not14/_0_  (.Y(net219),
    .A(net757));
 sg13g2_inv_1 \not15/_0_  (.Y(net220),
    .A(net739));
 sg13g2_inv_1 \not16/_0_  (.Y(net224),
    .A(net745));
 sg13g2_inv_1 \not17/_0_  (.Y(net225),
    .A(net735));
 sg13g2_inv_1 \not18/_0_  (.Y(net229),
    .A(net755));
 sg13g2_inv_1 \not19/_0_  (.Y(net230),
    .A(net745));
 sg13g2_inv_1 \not2/_0_  (.Y(net134),
    .A(net740));
 sg13g2_inv_1 \not20/_0_  (.Y(net232),
    .A(net753));
 sg13g2_inv_1 \not21/_0_  (.Y(net233),
    .A(net738));
 sg13g2_inv_1 \not22/_0_  (.Y(net242),
    .A(net747));
 sg13g2_inv_1 \not23/_0_  (.Y(net238),
    .A(net739));
 sg13g2_inv_1 \not24/_0_  (.Y(net243),
    .A(net756));
 sg13g2_inv_1 \not25/_0_  (.Y(net244),
    .A(net737));
 sg13g2_inv_1 \not26/_0_  (.Y(net246),
    .A(net737));
 sg13g2_inv_1 \not27/_0_  (.Y(net248),
    .A(net744));
 sg13g2_inv_1 \not28/_0_  (.Y(net249),
    .A(net736));
 sg13g2_inv_1 \not29/_0_  (.Y(net251),
    .A(net744));
 sg13g2_inv_1 \not3/_0_  (.Y(net135),
    .A(net2));
 sg13g2_inv_1 \not30/_0_  (.Y(net253),
    .A(net736));
 sg13g2_inv_1 \not31/_0_  (.Y(net256),
    .A(net752));
 sg13g2_inv_1 \not32/_0_  (.Y(net258),
    .A(net743));
 sg13g2_inv_1 \not33/_0_  (.Y(net260),
    .A(net736));
 sg13g2_inv_1 \not34/_0_  (.Y(net263),
    .A(net757));
 sg13g2_inv_1 \not35/_0_  (.Y(net264),
    .A(net740));
 sg13g2_inv_1 \not36/_0_  (.Y(net273),
    .A(net737));
 sg13g2_inv_1 \not37/_0_  (.Y(net272),
    .A(net745));
 sg13g2_inv_1 \not38/_0_  (.Y(net270),
    .A(net755));
 sg13g2_inv_1 \not39/_0_  (.Y(net275),
    .A(net745));
 sg13g2_inv_1 \not4/_0_  (.Y(net158),
    .A(net725));
 sg13g2_inv_1 \not40/_0_  (.Y(net284),
    .A(net753));
 sg13g2_inv_1 \not41/_0_  (.Y(net283),
    .A(net738));
 sg13g2_inv_1 \not42/_0_  (.Y(net282),
    .A(net753));
 sg13g2_inv_1 \not43/_0_  (.Y(net285),
    .A(net747));
 sg13g2_inv_1 \not44/_0_  (.Y(net286),
    .A(net755));
 sg13g2_inv_1 \not45/_0_  (.Y(net292),
    .A(net737));
 sg13g2_inv_1 \not46/_0_  (.Y(net291),
    .A(net737));
 sg13g2_inv_1 \not47/_0_  (.Y(net300),
    .A(net736));
 sg13g2_inv_1 \not48/_0_  (.Y(net297),
    .A(net744));
 sg13g2_inv_1 \not49/_0_  (.Y(net299),
    .A(net744));
 sg13g2_inv_1 \not5/_0_  (.Y(net160),
    .A(net159));
 sg13g2_inv_1 \not50/_0_  (.Y(net298),
    .A(net736));
 sg13g2_inv_1 \not51/_0_  (.Y(net307),
    .A(net752));
 sg13g2_inv_1 \not52/_0_  (.Y(net305),
    .A(net743));
 sg13g2_inv_1 \not53/_0_  (.Y(net306),
    .A(net737));
 sg13g2_inv_1 \not54/_0_  (.Y(net288),
    .A(net739));
 sg13g2_inv_1 \not55/_0_  (.Y(net308),
    .A(net744));
 sg13g2_inv_1 \not56/_0_  (.Y(net313),
    .A(net736));
 sg13g2_inv_1 \not57/_0_  (.Y(net315),
    .A(net736));
 sg13g2_inv_1 \not58/_0_  (.Y(net314),
    .A(net746));
 sg13g2_inv_1 \not59/_0_  (.Y(net316),
    .A(net743));
 sg13g2_inv_1 \not6/_0_  (.Y(net162),
    .A(net161));
 sg13g2_inv_1 \not60/_0_  (.Y(net320),
    .A(net736));
 sg13g2_inv_1 \not61/_0_  (.Y(net322),
    .A(net751));
 sg13g2_inv_1 \not62/_0_  (.Y(net323),
    .A(net735));
 sg13g2_inv_1 \not63/_0_  (.Y(net326),
    .A(net735));
 sg13g2_inv_1 \not64/_0_  (.Y(net327),
    .A(net754));
 sg13g2_inv_1 \not65/_0_  (.Y(net329),
    .A(net746));
 sg13g2_inv_1 \not66/_0_  (.Y(net330),
    .A(net738));
 sg13g2_inv_1 \not67/_0_  (.Y(net331),
    .A(net753));
 sg13g2_inv_1 \not68/_0_  (.Y(net335),
    .A(net753));
 sg13g2_inv_1 \not69/_0_  (.Y(net336),
    .A(net738));
 sg13g2_inv_1 \not7/_0_  (.Y(net181),
    .A(net169));
 sg13g2_inv_1 \not70/_0_  (.Y(net339),
    .A(net747));
 sg13g2_inv_1 \not71/_0_  (.Y(net345),
    .A(net754));
 sg13g2_inv_1 \not72/_0_  (.Y(net346),
    .A(net753));
 sg13g2_inv_1 \not73/_0_  (.Y(net347),
    .A(net738));
 sg13g2_inv_1 \not74/_0_  (.Y(net349),
    .A(net755));
 sg13g2_inv_1 \not75/_0_  (.Y(net350),
    .A(net748));
 sg13g2_inv_1 \not76/_0_  (.Y(net351),
    .A(net735));
 sg13g2_inv_1 \not77/_0_  (.Y(net359),
    .A(net724));
 sg13g2_inv_1 \not78/_0_  (.Y(net361),
    .A(net719));
 sg13g2_inv_1 \not79/_0_  (.Y(net362),
    .A(net719));
 sg13g2_inv_1 \not8/_0_  (.Y(net188),
    .A(net1));
 sg13g2_inv_1 \not80/_0_  (.Y(net365),
    .A(net718));
 sg13g2_inv_1 \not81/_0_  (.Y(net366),
    .A(net721));
 sg13g2_inv_1 \not82/_0_  (.Y(net367),
    .A(net723));
 sg13g2_inv_1 \not83/_0_  (.Y(net372),
    .A(net721));
 sg13g2_inv_1 \not84/_0_  (.Y(net373),
    .A(net724));
 sg13g2_inv_1 \not85/_0_  (.Y(net374),
    .A(net719));
 sg13g2_inv_1 \not86/_0_  (.Y(net378),
    .A(net719));
 sg13g2_inv_1 \not87/_0_  (.Y(net379),
    .A(net724));
 sg13g2_inv_1 \not88/_0_  (.Y(net382),
    .A(net722));
 sg13g2_inv_1 \not89/_0_  (.Y(net385),
    .A(net723));
 sg13g2_inv_1 \not9/_0_  (.Y(net203),
    .A(net693));
 sg13g2_inv_1 \not90/_0_  (.Y(net388),
    .A(net723));
 sg13g2_inv_1 \not91/_0_  (.Y(net389),
    .A(net718));
 sg13g2_inv_1 \not92/_0_  (.Y(net390),
    .A(net721));
 sg13g2_inv_1 \not93/_0_  (.Y(net395),
    .A(net723));
 sg13g2_inv_1 \not94/_0_  (.Y(net397),
    .A(net723));
 sg13g2_inv_1 \not95/_0_  (.Y(net396),
    .A(net721));
 sg13g2_inv_1 \not96/_0_  (.Y(net398),
    .A(net721));
 sg13g2_inv_1 \not97/_0_  (.Y(net402),
    .A(net723));
 sg13g2_inv_1 \not98/_0_  (.Y(net404),
    .A(net718));
 sg13g2_inv_1 \not99/_0_  (.Y(net407),
    .A(net1));
 sg13g2_or2_1 \or1/_0_  (.X(net138),
    .B(net136),
    .A(net137));
 sg13g2_or2_1 \or10/_0_  (.X(net151),
    .B(net149),
    .A(net150));
 sg13g2_or2_1 \or100/_0_  (.X(net37),
    .B(net434),
    .A(net420));
 sg13g2_or2_1 \or101/_0_  (.X(net435),
    .B(net416),
    .A(net421));
 sg13g2_or2_1 \or102/_0_  (.X(net53),
    .B(net435),
    .A(net419));
 sg13g2_or2_1 \or103/_0_  (.X(net436),
    .B(net428),
    .A(net427));
 sg13g2_or2_1 \or104/_0_  (.X(net437),
    .B(net414),
    .A(net424));
 sg13g2_or2_1 \or105/_0_  (.X(net438),
    .B(net436),
    .A(net437));
 sg13g2_or2_1 \or106/_0_  (.X(net69),
    .B(net438),
    .A(net432));
 sg13g2_or2_1 \or107/_0_  (.X(net85),
    .B(net428),
    .A(net424));
 sg13g2_or2_1 \or108/_0_  (.X(net439),
    .B(net429),
    .A(net426));
 sg13g2_or2_1 \or109/_0_  (.X(net440),
    .B(net431),
    .A(net414));
 sg13g2_or2_1 \or11/_0_  (.X(net110),
    .B(net151),
    .A(net145));
 sg13g2_or2_1 \or110/_0_  (.X(net101),
    .B(net439),
    .A(net440));
 sg13g2_or2_1 \or111/_0_  (.X(net441),
    .B(net428),
    .A(net429));
 sg13g2_or2_1 \or112/_0_  (.X(net442),
    .B(net414),
    .A(net427));
 sg13g2_or2_1 \or113/_0_  (.X(net117),
    .B(net441),
    .A(net442));
 sg13g2_or2_1 \or114/_0_  (.X(net452),
    .B(net450),
    .A(net444));
 sg13g2_or2_1 \or115/_0_  (.X(net453),
    .B(net452),
    .A(net451));
 sg13g2_or2_1 \or116/_0_  (.X(net455),
    .B(net447),
    .A(net454));
 sg13g2_or2_1 \or117/_0_  (.X(net457),
    .B(net455),
    .A(net456));
 sg13g2_or2_1 \or118/_0_  (.X(net458),
    .B(net448),
    .A(net446));
 sg13g2_or2_1 \or119/_0_  (.X(net459),
    .B(net458),
    .A(net445));
 sg13g2_or2_1 \or12/_0_  (.X(net94),
    .B(net141),
    .A(net137));
 sg13g2_or2_1 \or120/_0_  (.X(net462),
    .B(net460),
    .A(net461));
 sg13g2_or2_1 \or121/_0_  (.X(net466),
    .B(net463),
    .A(net465));
 sg13g2_or2_1 \or122/_0_  (.X(net467),
    .B(net462),
    .A(net466));
 sg13g2_or2_1 \or123/_0_  (.X(net470),
    .B(net468),
    .A(net469));
 sg13g2_or2_1 \or124/_0_  (.X(net473),
    .B(net471),
    .A(net472));
 sg13g2_or2_1 \or125/_0_  (.X(net475),
    .B(net473),
    .A(net474));
 sg13g2_or2_1 \or126/_0_  (.X(net478),
    .B(net476),
    .A(net477));
 sg13g2_or2_1 \or127/_0_  (.X(net480),
    .B(net478),
    .A(net479));
 sg13g2_or2_1 \or128/_0_  (.X(net502),
    .B(net500),
    .A(net501));
 sg13g2_or2_1 \or129/_0_  (.X(net505),
    .B(net503),
    .A(net504));
 sg13g2_or2_1 \or13/_0_  (.X(net152),
    .B(net142),
    .A(net139));
 sg13g2_or2_1 \or130/_0_  (.X(net508),
    .B(net506),
    .A(net507));
 sg13g2_or2_1 \or131/_0_  (.X(net509),
    .B(net490),
    .A(net495));
 sg13g2_or2_1 \or132/_0_  (.X(net511),
    .B(net510),
    .A(net496));
 sg13g2_or2_1 \or133/_0_  (.X(net514),
    .B(net512),
    .A(net513));
 sg13g2_or2_1 \or134/_0_  (.X(net503),
    .B(net496),
    .A(net499));
 sg13g2_or2_1 \or135/_0_  (.X(net504),
    .B(net515),
    .A(net498));
 sg13g2_or2_1 \or136/_0_  (.X(net517),
    .B(net516),
    .A(net492));
 sg13g2_or2_1 \or137/_0_  (.X(net516),
    .B(net518),
    .A(net519));
 sg13g2_or2_1 \or138/_0_  (.X(net519),
    .B(net495),
    .A(net494));
 sg13g2_or2_1 \or139/_0_  (.X(net518),
    .B(net515),
    .A(net490));
 sg13g2_or2_1 \or14/_0_  (.X(net153),
    .B(net144),
    .A(net758));
 sg13g2_or2_1 \or140/_0_  (.X(net510),
    .B(net486),
    .A(net488));
 sg13g2_or2_1 \or141/_0_  (.X(net513),
    .B(net497),
    .A(net496));
 sg13g2_or2_1 \or142/_0_  (.X(net512),
    .B(net515),
    .A(net487));
 sg13g2_or2_1 \or143/_0_  (.X(net501),
    .B(net491),
    .A(net484));
 sg13g2_or2_1 \or144/_0_  (.X(net500),
    .B(net515),
    .A(net490));
 sg13g2_or2_1 \or145/_0_  (.X(net506),
    .B(net515),
    .A(net499));
 sg13g2_or2_1 \or146/_0_  (.X(net507),
    .B(net498),
    .A(net492));
 sg13g2_or2_1 \or147/_0_  (.X(net615),
    .B(net614),
    .A(net547));
 sg13g2_or2_1 \or148/_0_  (.X(net616),
    .B(net614),
    .A(net547));
 sg13g2_or2_1 \or15/_0_  (.X(net62),
    .B(net152),
    .A(net153));
 sg13g2_or2_1 \or16/_0_  (.X(net154),
    .B(net141),
    .A(net142));
 sg13g2_or2_1 \or17/_0_  (.X(net155),
    .B(net758),
    .A(net140));
 sg13g2_or2_1 \or18/_0_  (.X(net78),
    .B(net154),
    .A(net155));
 sg13g2_or2_1 \or19/_0_  (.X(net31),
    .B(net172),
    .A(net173));
 sg13g2_or2_1 \or2/_0_  (.X(net146),
    .B(net756),
    .A(net740));
 sg13g2_or2_1 \or20/_0_  (.X(net173),
    .B(net163),
    .A(net161));
 sg13g2_or2_1 \or21/_0_  (.X(net172),
    .B(net174),
    .A(net166));
 sg13g2_or2_1 \or22/_0_  (.X(net47),
    .B(net175),
    .A(net176));
 sg13g2_or2_1 \or23/_0_  (.X(net176),
    .B(net168),
    .A(net167));
 sg13g2_or2_1 \or24/_0_  (.X(net175),
    .B(net160),
    .A(net174));
 sg13g2_or2_1 \or25/_0_  (.X(net177),
    .B(net164),
    .A(net170));
 sg13g2_or2_1 \or26/_0_  (.X(net63),
    .B(net178),
    .A(net725));
 sg13g2_or2_1 \or27/_0_  (.X(net178),
    .B(net159),
    .A(net167));
 sg13g2_or2_1 \or28/_0_  (.X(net79),
    .B(net177),
    .A(net179));
 sg13g2_or2_1 \or29/_0_  (.X(net179),
    .B(net166),
    .A(net180));
 sg13g2_or2_1 \or3/_0_  (.X(net46),
    .B(net138),
    .A(net146));
 sg13g2_or2_1 \or30/_0_  (.X(net111),
    .B(net182),
    .A(net183));
 sg13g2_or2_1 \or31/_0_  (.X(net183),
    .B(net167),
    .A(net169));
 sg13g2_or2_1 \or32/_0_  (.X(net182),
    .B(net174),
    .A(net165));
 sg13g2_or2_1 \or33/_0_  (.X(net127),
    .B(net184),
    .A(net185));
 sg13g2_or2_1 \or34/_0_  (.X(net185),
    .B(net170),
    .A(net169));
 sg13g2_or2_1 \or35/_0_  (.X(net184),
    .B(net174),
    .A(net164));
 sg13g2_or2_1 \or36/_0_  (.X(net202),
    .B(net200),
    .A(net201));
 sg13g2_or2_1 \or37/_0_  (.X(net208),
    .B(net205),
    .A(net207));
 sg13g2_or2_1 \or38/_0_  (.X(net194),
    .B(net209),
    .A(net210));
 sg13g2_or2_1 \or39/_0_  (.X(net215),
    .B(net213),
    .A(net214));
 sg13g2_or2_1 \or4/_0_  (.X(net147),
    .B(net143),
    .A(net144));
 sg13g2_or2_1 \or40/_0_  (.X(net223),
    .B(net221),
    .A(net222));
 sg13g2_or2_1 \or41/_0_  (.X(net27),
    .B(net223),
    .A(net749));
 sg13g2_or2_1 \or42/_0_  (.X(net228),
    .B(net226),
    .A(net227));
 sg13g2_or2_1 \or43/_0_  (.X(net43),
    .B(net228),
    .A(net229));
 sg13g2_or2_1 \or44/_0_  (.X(net231),
    .B(net230),
    .A(net741));
 sg13g2_or2_1 \or45/_0_  (.X(net59),
    .B(net231),
    .A(net756));
 sg13g2_or2_1 \or46/_0_  (.X(net240),
    .B(net234),
    .A(net235));
 sg13g2_or2_1 \or47/_0_  (.X(net75),
    .B(net240),
    .A(net241));
 sg13g2_or2_1 \or48/_0_  (.X(net241),
    .B(net237),
    .A(net239));
 sg13g2_or2_1 \or49/_0_  (.X(net91),
    .B(net245),
    .A(net247));
 sg13g2_or2_1 \or5/_0_  (.X(net30),
    .B(net147),
    .A(net133));
 sg13g2_or2_1 \or50/_0_  (.X(net255),
    .B(net250),
    .A(net252));
 sg13g2_or2_1 \or51/_0_  (.X(net107),
    .B(net255),
    .A(net254));
 sg13g2_or2_1 \or52/_0_  (.X(net262),
    .B(net257),
    .A(net259));
 sg13g2_or2_1 \or53/_0_  (.X(net123),
    .B(net262),
    .A(net261));
 sg13g2_or2_1 \or54/_0_  (.X(net266),
    .B(net749),
    .A(net265));
 sg13g2_or2_1 \or55/_0_  (.X(net28),
    .B(net266),
    .A(net267));
 sg13g2_or2_1 \or56/_0_  (.X(net44),
    .B(net268),
    .A(net269));
 sg13g2_or2_1 \or57/_0_  (.X(net268),
    .B(net270),
    .A(net271));
 sg13g2_or2_1 \or58/_0_  (.X(net60),
    .B(net274),
    .A(net275));
 sg13g2_or2_1 \or59/_0_  (.X(net274),
    .B(net756),
    .A(net741));
 sg13g2_or2_1 \or6/_0_  (.X(net148),
    .B(net749),
    .A(net134));
 sg13g2_or2_1 \or60/_0_  (.X(net278),
    .B(net276),
    .A(net277));
 sg13g2_or2_1 \or61/_0_  (.X(net281),
    .B(net279),
    .A(net280));
 sg13g2_or2_1 \or62/_0_  (.X(net76),
    .B(net278),
    .A(net281));
 sg13g2_or2_1 \or63/_0_  (.X(net92),
    .B(net289),
    .A(net290));
 sg13g2_or2_1 \or64/_0_  (.X(net108),
    .B(net293),
    .A(net294));
 sg13g2_or2_1 \or65/_0_  (.X(net293),
    .B(net295),
    .A(net296));
 sg13g2_or2_1 \or66/_0_  (.X(net124),
    .B(net301),
    .A(net302));
 sg13g2_or2_1 \or67/_0_  (.X(net301),
    .B(net303),
    .A(net304));
 sg13g2_or2_1 \or68/_0_  (.X(net104),
    .B(net310),
    .A(net311));
 sg13g2_or2_1 \or69/_0_  (.X(net310),
    .B(net309),
    .A(net312));
 sg13g2_or2_1 \or7/_0_  (.X(net126),
    .B(net148),
    .A(net2));
 sg13g2_or2_1 \or70/_0_  (.X(net319),
    .B(net317),
    .A(net318));
 sg13g2_or2_1 \or71/_0_  (.X(net120),
    .B(net319),
    .A(net321));
 sg13g2_or2_1 \or72/_0_  (.X(net88),
    .B(net324),
    .A(net325));
 sg13g2_or2_1 \or73/_0_  (.X(net328),
    .B(net754),
    .A(net735));
 sg13g2_or2_1 \or74/_0_  (.X(net56),
    .B(net328),
    .A(net329));
 sg13g2_or2_1 \or75/_0_  (.X(net334),
    .B(net332),
    .A(net333));
 sg13g2_or2_1 \or76/_0_  (.X(net341),
    .B(net337),
    .A(net340));
 sg13g2_or2_1 \or77/_0_  (.X(net72),
    .B(net334),
    .A(net341));
 sg13g2_or2_1 \or78/_0_  (.X(net344),
    .B(net342),
    .A(net343));
 sg13g2_or2_1 \or79/_0_  (.X(net24),
    .B(net344),
    .A(net348));
 sg13g2_or2_1 \or8/_0_  (.X(net149),
    .B(net141),
    .A(net140));
 sg13g2_or2_1 \or80/_0_  (.X(net40),
    .B(net353),
    .A(net354));
 sg13g2_or2_1 \or81/_0_  (.X(net353),
    .B(net349),
    .A(net352));
 sg13g2_or2_1 \or82/_0_  (.X(net357),
    .B(net355),
    .A(net356));
 sg13g2_or2_1 \or83/_0_  (.X(net25),
    .B(net357),
    .A(net364));
 sg13g2_or2_1 \or84/_0_  (.X(net41),
    .B(net369),
    .A(net370));
 sg13g2_or2_1 \or85/_0_  (.X(net369),
    .B(net365),
    .A(net368));
 sg13g2_or2_1 \or86/_0_  (.X(net371),
    .B(net718),
    .A(net723));
 sg13g2_or2_1 \or87/_0_  (.X(net57),
    .B(net371),
    .A(net372));
 sg13g2_or2_1 \or88/_0_  (.X(net377),
    .B(net375),
    .A(net376));
 sg13g2_or2_1 \or89/_0_  (.X(net384),
    .B(net380),
    .A(net383));
 sg13g2_or2_1 \or9/_0_  (.X(net150),
    .B(net756),
    .A(net137));
 sg13g2_or2_1 \or90/_0_  (.X(net73),
    .B(net377),
    .A(net384));
 sg13g2_or2_1 \or91/_0_  (.X(net89),
    .B(net386),
    .A(net387));
 sg13g2_or2_1 \or92/_0_  (.X(net105),
    .B(net392),
    .A(net393));
 sg13g2_or2_1 \or93/_0_  (.X(net392),
    .B(net391),
    .A(net394));
 sg13g2_or2_1 \or94/_0_  (.X(net401),
    .B(net399),
    .A(net400));
 sg13g2_or2_1 \or95/_0_  (.X(net121),
    .B(net401),
    .A(net403));
 sg13g2_or2_1 \or96/_0_  (.X(net425),
    .B(net423),
    .A(net424));
 sg13g2_or2_1 \or97/_0_  (.X(net433),
    .B(net414),
    .A(net418));
 sg13g2_or2_1 \or98/_0_  (.X(net21),
    .B(net425),
    .A(net433));
 sg13g2_or2_1 \or99/_0_  (.X(net434),
    .B(net430),
    .A(net431));
 sg13g2_buf_2 fanout126 (.A(net360),
    .X(net718));
 sg13g2_buf_1 fanout127 (.A(net360),
    .X(net719));
 sg13g2_buf_2 fanout128 (.A(net449),
    .X(net720));
 sg13g2_buf_2 fanout129 (.A(net363),
    .X(net721));
 sg13g2_buf_1 fanout130 (.A(net363),
    .X(net722));
 sg13g2_buf_2 fanout131 (.A(net358),
    .X(net723));
 sg13g2_buf_1 fanout132 (.A(net358),
    .X(net724));
 sg13g2_buf_2 fanout133 (.A(net157),
    .X(net725));
 sg13g2_buf_4 fanout134 (.X(net726),
    .A(net729));
 sg13g2_buf_2 fanout135 (.A(net729),
    .X(net727));
 sg13g2_buf_4 fanout136 (.X(net728),
    .A(net729));
 sg13g2_buf_2 fanout137 (.A(ui_in[5]),
    .X(net729));
 sg13g2_buf_4 fanout138 (.X(net730),
    .A(net731));
 sg13g2_buf_2 fanout139 (.A(ui_in[4]),
    .X(net731));
 sg13g2_buf_4 fanout140 (.X(net732),
    .A(net734));
 sg13g2_buf_4 fanout141 (.X(net733),
    .A(net734));
 sg13g2_buf_2 fanout142 (.A(ui_in[4]),
    .X(net734));
 sg13g2_buf_2 fanout143 (.A(net737),
    .X(net735));
 sg13g2_buf_2 fanout144 (.A(net737),
    .X(net736));
 sg13g2_buf_2 fanout145 (.A(net741),
    .X(net737));
 sg13g2_buf_2 fanout146 (.A(net739),
    .X(net738));
 sg13g2_buf_1 fanout147 (.A(net740),
    .X(net739));
 sg13g2_buf_2 fanout148 (.A(net741),
    .X(net740));
 sg13g2_buf_1 fanout149 (.A(ui_in[2]),
    .X(net741));
 sg13g2_buf_4 fanout150 (.X(net742),
    .A(net750));
 sg13g2_buf_2 fanout151 (.A(net750),
    .X(net743));
 sg13g2_buf_2 fanout152 (.A(net745),
    .X(net744));
 sg13g2_buf_2 fanout153 (.A(net746),
    .X(net745));
 sg13g2_buf_2 fanout154 (.A(net750),
    .X(net746));
 sg13g2_buf_2 fanout155 (.A(net748),
    .X(net747));
 sg13g2_buf_1 fanout156 (.A(net749),
    .X(net748));
 sg13g2_buf_2 fanout157 (.A(net750),
    .X(net749));
 sg13g2_buf_2 fanout158 (.A(ui_in[1]),
    .X(net750));
 sg13g2_buf_2 fanout159 (.A(net759),
    .X(net751));
 sg13g2_buf_2 fanout160 (.A(net759),
    .X(net752));
 sg13g2_buf_2 fanout161 (.A(net754),
    .X(net753));
 sg13g2_buf_2 fanout162 (.A(net759),
    .X(net754));
 sg13g2_buf_2 fanout163 (.A(net758),
    .X(net755));
 sg13g2_buf_1 fanout164 (.A(net758),
    .X(net756));
 sg13g2_buf_2 fanout165 (.A(net758),
    .X(net757));
 sg13g2_buf_2 fanout166 (.A(net759),
    .X(net758));
 sg13g2_buf_2 fanout167 (.A(ui_in[0]),
    .X(net759));
 sg13g2_buf_4 input1 (.X(net1),
    .A(rst_n));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[6]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[7]));
 sg13g2_tielo \flop1/_4__5  (.L_LO(net5));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_4 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_144 ();
 sg13g2_fill_1 FILLER_17_151 ();
 sg13g2_decap_8 FILLER_17_159 ();
 sg13g2_decap_8 FILLER_17_166 ();
 sg13g2_fill_1 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_fill_2 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_fill_2 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_127 ();
 sg13g2_decap_8 FILLER_18_167 ();
 sg13g2_decap_4 FILLER_18_186 ();
 sg13g2_fill_1 FILLER_18_190 ();
 sg13g2_fill_2 FILLER_18_197 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_109 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_decap_4 FILLER_19_127 ();
 sg13g2_fill_2 FILLER_19_131 ();
 sg13g2_decap_8 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_150 ();
 sg13g2_fill_1 FILLER_19_152 ();
 sg13g2_decap_8 FILLER_19_156 ();
 sg13g2_decap_4 FILLER_19_163 ();
 sg13g2_fill_2 FILLER_19_167 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_220 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_233 ();
 sg13g2_decap_8 FILLER_19_240 ();
 sg13g2_decap_8 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_254 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_decap_4 FILLER_19_282 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_decap_4 FILLER_20_154 ();
 sg13g2_fill_1 FILLER_20_193 ();
 sg13g2_decap_4 FILLER_20_200 ();
 sg13g2_fill_1 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_4 FILLER_20_264 ();
 sg13g2_fill_2 FILLER_20_268 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_112 ();
 sg13g2_fill_1 FILLER_21_114 ();
 sg13g2_decap_8 FILLER_21_123 ();
 sg13g2_fill_2 FILLER_21_130 ();
 sg13g2_fill_1 FILLER_21_132 ();
 sg13g2_fill_2 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_142 ();
 sg13g2_decap_8 FILLER_21_146 ();
 sg13g2_decap_4 FILLER_21_153 ();
 sg13g2_fill_2 FILLER_21_157 ();
 sg13g2_fill_2 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_177 ();
 sg13g2_decap_4 FILLER_21_184 ();
 sg13g2_fill_2 FILLER_21_188 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_207 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_decap_8 FILLER_21_215 ();
 sg13g2_decap_8 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_234 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_decap_8 FILLER_21_263 ();
 sg13g2_fill_2 FILLER_21_270 ();
 sg13g2_fill_2 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_282 ();
 sg13g2_fill_2 FILLER_21_290 ();
 sg13g2_fill_1 FILLER_21_292 ();
 sg13g2_decap_4 FILLER_21_296 ();
 sg13g2_fill_2 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_4 FILLER_22_73 ();
 sg13g2_fill_1 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_4 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_149 ();
 sg13g2_fill_1 FILLER_22_155 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_172 ();
 sg13g2_fill_1 FILLER_22_183 ();
 sg13g2_decap_4 FILLER_22_209 ();
 sg13g2_fill_2 FILLER_22_213 ();
 sg13g2_decap_8 FILLER_22_225 ();
 sg13g2_decap_8 FILLER_22_232 ();
 sg13g2_decap_4 FILLER_22_239 ();
 sg13g2_fill_1 FILLER_22_243 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_fill_1 FILLER_22_261 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_fill_2 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_318 ();
 sg13g2_decap_8 FILLER_22_325 ();
 sg13g2_decap_8 FILLER_22_332 ();
 sg13g2_decap_8 FILLER_22_339 ();
 sg13g2_decap_8 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_353 ();
 sg13g2_decap_8 FILLER_22_360 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_4 FILLER_23_45 ();
 sg13g2_fill_2 FILLER_23_49 ();
 sg13g2_fill_2 FILLER_23_86 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_151 ();
 sg13g2_fill_2 FILLER_23_163 ();
 sg13g2_decap_8 FILLER_23_180 ();
 sg13g2_fill_2 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_201 ();
 sg13g2_decap_4 FILLER_23_207 ();
 sg13g2_fill_2 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_254 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_4 FILLER_23_301 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_decap_4 FILLER_23_320 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_decap_8 FILLER_23_344 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_4 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_25 ();
 sg13g2_decap_4 FILLER_24_66 ();
 sg13g2_fill_1 FILLER_24_70 ();
 sg13g2_decap_4 FILLER_24_75 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_131 ();
 sg13g2_decap_8 FILLER_24_138 ();
 sg13g2_fill_2 FILLER_24_145 ();
 sg13g2_decap_4 FILLER_24_162 ();
 sg13g2_decap_8 FILLER_24_181 ();
 sg13g2_decap_8 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_195 ();
 sg13g2_decap_4 FILLER_24_207 ();
 sg13g2_fill_2 FILLER_24_232 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_fill_2 FILLER_24_265 ();
 sg13g2_fill_2 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_274 ();
 sg13g2_fill_2 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_decap_4 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_fill_2 FILLER_24_313 ();
 sg13g2_fill_2 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_24_358 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_28 ();
 sg13g2_decap_4 FILLER_25_38 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_47 ();
 sg13g2_fill_2 FILLER_25_51 ();
 sg13g2_fill_2 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_62 ();
 sg13g2_decap_8 FILLER_25_68 ();
 sg13g2_fill_2 FILLER_25_78 ();
 sg13g2_fill_1 FILLER_25_91 ();
 sg13g2_decap_4 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_137 ();
 sg13g2_fill_1 FILLER_25_171 ();
 sg13g2_decap_4 FILLER_25_177 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_205 ();
 sg13g2_fill_2 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_fill_1 FILLER_25_234 ();
 sg13g2_fill_2 FILLER_25_252 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_fill_2 FILLER_25_279 ();
 sg13g2_decap_4 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_decap_4 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_89 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_fill_2 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_125 ();
 sg13g2_fill_2 FILLER_26_136 ();
 sg13g2_fill_1 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_169 ();
 sg13g2_decap_4 FILLER_26_176 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_fill_2 FILLER_26_186 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_decap_4 FILLER_26_211 ();
 sg13g2_decap_8 FILLER_26_225 ();
 sg13g2_decap_8 FILLER_26_232 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_260 ();
 sg13g2_fill_1 FILLER_26_262 ();
 sg13g2_decap_8 FILLER_26_269 ();
 sg13g2_decap_8 FILLER_26_276 ();
 sg13g2_fill_1 FILLER_26_283 ();
 sg13g2_fill_1 FILLER_26_287 ();
 sg13g2_decap_4 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_decap_4 FILLER_26_321 ();
 sg13g2_fill_1 FILLER_26_325 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_decap_4 FILLER_27_42 ();
 sg13g2_fill_1 FILLER_27_57 ();
 sg13g2_decap_8 FILLER_27_61 ();
 sg13g2_fill_2 FILLER_27_71 ();
 sg13g2_decap_4 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_decap_4 FILLER_27_88 ();
 sg13g2_fill_1 FILLER_27_92 ();
 sg13g2_fill_2 FILLER_27_96 ();
 sg13g2_fill_1 FILLER_27_111 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_138 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_204 ();
 sg13g2_fill_1 FILLER_27_211 ();
 sg13g2_decap_8 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_293 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_336 ();
 sg13g2_fill_1 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_8 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_64 ();
 sg13g2_fill_1 FILLER_28_97 ();
 sg13g2_fill_2 FILLER_28_108 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_146 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_165 ();
 sg13g2_decap_4 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_186 ();
 sg13g2_decap_4 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_fill_1 FILLER_28_211 ();
 sg13g2_decap_4 FILLER_28_230 ();
 sg13g2_fill_2 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_fill_2 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_285 ();
 sg13g2_decap_4 FILLER_28_292 ();
 sg13g2_decap_8 FILLER_28_309 ();
 sg13g2_decap_4 FILLER_28_329 ();
 sg13g2_fill_1 FILLER_28_333 ();
 sg13g2_fill_2 FILLER_28_339 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_decap_8 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_365 ();
 sg13g2_decap_8 FILLER_28_372 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_67 ();
 sg13g2_decap_8 FILLER_29_72 ();
 sg13g2_decap_8 FILLER_29_79 ();
 sg13g2_decap_8 FILLER_29_89 ();
 sg13g2_decap_8 FILLER_29_96 ();
 sg13g2_decap_4 FILLER_29_103 ();
 sg13g2_fill_1 FILLER_29_110 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_decap_8 FILLER_29_124 ();
 sg13g2_decap_4 FILLER_29_131 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_decap_4 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_163 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_fill_2 FILLER_29_183 ();
 sg13g2_fill_1 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_191 ();
 sg13g2_fill_1 FILLER_29_201 ();
 sg13g2_decap_8 FILLER_29_223 ();
 sg13g2_decap_8 FILLER_29_243 ();
 sg13g2_fill_2 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_332 ();
 sg13g2_decap_8 FILLER_29_360 ();
 sg13g2_decap_8 FILLER_29_367 ();
 sg13g2_decap_8 FILLER_29_374 ();
 sg13g2_decap_8 FILLER_29_381 ();
 sg13g2_decap_8 FILLER_29_388 ();
 sg13g2_decap_8 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_28 ();
 sg13g2_decap_4 FILLER_30_38 ();
 sg13g2_fill_2 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_132 ();
 sg13g2_decap_4 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_144 ();
 sg13g2_fill_2 FILLER_30_155 ();
 sg13g2_fill_1 FILLER_30_157 ();
 sg13g2_fill_2 FILLER_30_168 ();
 sg13g2_decap_4 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_204 ();
 sg13g2_decap_4 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_249 ();
 sg13g2_decap_4 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_277 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_decap_4 FILLER_30_302 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_decap_4 FILLER_30_333 ();
 sg13g2_fill_2 FILLER_30_340 ();
 sg13g2_fill_1 FILLER_30_342 ();
 sg13g2_fill_2 FILLER_30_348 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_4 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_fill_2 FILLER_31_74 ();
 sg13g2_fill_1 FILLER_31_76 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_99 ();
 sg13g2_fill_2 FILLER_31_106 ();
 sg13g2_fill_1 FILLER_31_112 ();
 sg13g2_fill_1 FILLER_31_116 ();
 sg13g2_decap_8 FILLER_31_122 ();
 sg13g2_decap_4 FILLER_31_129 ();
 sg13g2_fill_2 FILLER_31_133 ();
 sg13g2_fill_2 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_decap_4 FILLER_31_175 ();
 sg13g2_decap_4 FILLER_31_182 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_decap_4 FILLER_31_203 ();
 sg13g2_decap_4 FILLER_31_226 ();
 sg13g2_fill_2 FILLER_31_230 ();
 sg13g2_fill_1 FILLER_31_237 ();
 sg13g2_decap_8 FILLER_31_256 ();
 sg13g2_fill_1 FILLER_31_263 ();
 sg13g2_decap_4 FILLER_31_277 ();
 sg13g2_decap_4 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_320 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_decap_8 FILLER_31_341 ();
 sg13g2_fill_2 FILLER_31_348 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_fill_2 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_84 ();
 sg13g2_decap_4 FILLER_32_124 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_148 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_211 ();
 sg13g2_decap_8 FILLER_32_216 ();
 sg13g2_decap_4 FILLER_32_223 ();
 sg13g2_decap_4 FILLER_32_258 ();
 sg13g2_fill_1 FILLER_32_262 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_fill_2 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_282 ();
 sg13g2_decap_8 FILLER_32_293 ();
 sg13g2_fill_1 FILLER_32_300 ();
 sg13g2_decap_8 FILLER_32_324 ();
 sg13g2_fill_1 FILLER_32_331 ();
 sg13g2_fill_2 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_decap_4 FILLER_32_353 ();
 sg13g2_fill_1 FILLER_32_357 ();
 sg13g2_decap_4 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_373 ();
 sg13g2_fill_2 FILLER_32_379 ();
 sg13g2_fill_2 FILLER_32_384 ();
 sg13g2_fill_1 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_96 ();
 sg13g2_fill_2 FILLER_33_103 ();
 sg13g2_decap_4 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_116 ();
 sg13g2_fill_2 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_150 ();
 sg13g2_decap_8 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_decap_8 FILLER_33_171 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_decap_8 FILLER_33_191 ();
 sg13g2_fill_2 FILLER_33_198 ();
 sg13g2_decap_4 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_242 ();
 sg13g2_decap_4 FILLER_33_252 ();
 sg13g2_decap_4 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_decap_4 FILLER_33_292 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_308 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_321 ();
 sg13g2_fill_2 FILLER_33_328 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_fill_2 FILLER_33_342 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_356 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_4 FILLER_33_368 ();
 sg13g2_fill_1 FILLER_33_372 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_fill_1 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_383 ();
 sg13g2_fill_1 FILLER_33_390 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_86 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_4 FILLER_34_98 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_decap_4 FILLER_34_108 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_123 ();
 sg13g2_fill_1 FILLER_34_132 ();
 sg13g2_fill_1 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_180 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_decap_4 FILLER_34_197 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_211 ();
 sg13g2_fill_2 FILLER_34_215 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_decap_4 FILLER_34_241 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_decap_8 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_fill_2 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_4 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_148 ();
 sg13g2_decap_8 FILLER_35_155 ();
 sg13g2_decap_8 FILLER_35_162 ();
 sg13g2_decap_4 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_186 ();
 sg13g2_fill_1 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_221 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_decap_8 FILLER_35_249 ();
 sg13g2_decap_4 FILLER_35_256 ();
 sg13g2_decap_4 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_272 ();
 sg13g2_fill_1 FILLER_35_296 ();
 sg13g2_decap_8 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_314 ();
 sg13g2_fill_2 FILLER_35_323 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_decap_8 FILLER_35_339 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_fill_1 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_362 ();
 sg13g2_fill_2 FILLER_35_376 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_fill_2 FILLER_35_388 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_4 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_92 ();
 sg13g2_decap_4 FILLER_36_99 ();
 sg13g2_decap_4 FILLER_36_109 ();
 sg13g2_fill_1 FILLER_36_113 ();
 sg13g2_decap_8 FILLER_36_117 ();
 sg13g2_decap_8 FILLER_36_124 ();
 sg13g2_decap_4 FILLER_36_174 ();
 sg13g2_decap_4 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_196 ();
 sg13g2_fill_1 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_decap_4 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_237 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_fill_2 FILLER_36_276 ();
 sg13g2_fill_1 FILLER_36_278 ();
 sg13g2_decap_4 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_fill_2 FILLER_36_347 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_4 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_2 FILLER_37_132 ();
 sg13g2_fill_1 FILLER_37_147 ();
 sg13g2_fill_2 FILLER_37_153 ();
 sg13g2_fill_1 FILLER_37_155 ();
 sg13g2_decap_4 FILLER_37_161 ();
 sg13g2_fill_2 FILLER_37_175 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_227 ();
 sg13g2_fill_1 FILLER_37_239 ();
 sg13g2_fill_2 FILLER_37_279 ();
 sg13g2_fill_1 FILLER_37_281 ();
 sg13g2_fill_2 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_decap_4 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_337 ();
 sg13g2_decap_4 FILLER_37_344 ();
 sg13g2_fill_2 FILLER_37_348 ();
 sg13g2_fill_1 FILLER_37_354 ();
 sg13g2_decap_4 FILLER_37_363 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_fill_1 FILLER_37_388 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_fill_2 FILLER_38_174 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_195 ();
 sg13g2_decap_4 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_219 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_decap_8 FILLER_38_230 ();
 sg13g2_fill_2 FILLER_38_237 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_4 FILLER_38_273 ();
 sg13g2_fill_1 FILLER_38_277 ();
 sg13g2_fill_2 FILLER_38_283 ();
 sg13g2_fill_1 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_4 FILLER_38_308 ();
 sg13g2_decap_4 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_342 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net623;
 assign uio_oe[1] = net624;
 assign uio_oe[2] = net625;
 assign uio_oe[3] = net626;
 assign uio_oe[4] = net627;
 assign uio_oe[5] = net628;
 assign uio_oe[6] = net629;
 assign uio_oe[7] = net630;
 assign uio_out[0] = net631;
 assign uio_out[1] = net632;
 assign uio_out[2] = net633;
 assign uio_out[3] = net634;
 assign uio_out[4] = net635;
 assign uio_out[5] = net636;
 assign uio_out[6] = net637;
 assign uio_out[7] = net638;
 assign uo_out[7] = net639;
endmodule

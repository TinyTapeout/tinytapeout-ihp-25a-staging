module tt_um_nvious_graphics (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \gradient_sky.x[0] ;
 wire \gradient_sky.x[1] ;
 wire \gradient_sky.y[0] ;
 wire \gradient_sky.y[1] ;
 wire \gradient_sky.y[2] ;
 wire \gradient_sky.y[3] ;
 wire \gradient_sky.y[4] ;
 wire \gradient_sky.y[5] ;
 wire \gradient_sky.y[6] ;
 wire hsync;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \hx0[0] ;
 wire \hy0[0] ;
 wire show;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;

 sg13g2_inv_2 _1595_ (.Y(_0392_),
    .A(net610));
 sg13g2_inv_2 _1596_ (.Y(_0403_),
    .A(net686));
 sg13g2_inv_2 _1597_ (.Y(_0414_),
    .A(net612));
 sg13g2_inv_2 _1598_ (.Y(_0425_),
    .A(net607));
 sg13g2_inv_2 _1599_ (.Y(_0436_),
    .A(net603));
 sg13g2_inv_4 _1600_ (.A(net581),
    .Y(_0447_));
 sg13g2_inv_4 _1601_ (.A(net571),
    .Y(_0458_));
 sg13g2_inv_1 _1602_ (.Y(_0469_),
    .A(net585));
 sg13g2_inv_2 _1603_ (.Y(_0480_),
    .A(net591));
 sg13g2_inv_4 _1604_ (.A(net568),
    .Y(_0491_));
 sg13g2_inv_4 _1605_ (.A(net562),
    .Y(_0502_));
 sg13g2_inv_4 _1606_ (.A(net617),
    .Y(_0513_));
 sg13g2_inv_1 _1607_ (.Y(_0524_),
    .A(net660));
 sg13g2_inv_1 _1608_ (.Y(_0535_),
    .A(net678));
 sg13g2_inv_2 _1609_ (.Y(_0546_),
    .A(net679));
 sg13g2_inv_4 _1610_ (.A(net631),
    .Y(_0557_));
 sg13g2_inv_1 _1611_ (.Y(_0568_),
    .A(net640));
 sg13g2_inv_2 _1612_ (.Y(_0577_),
    .A(net647));
 sg13g2_inv_1 _1613_ (.Y(_0588_),
    .A(net655));
 sg13g2_inv_2 _1614_ (.Y(_0597_),
    .A(net615));
 sg13g2_inv_4 _1615_ (.A(_0028_),
    .Y(_0605_));
 sg13g2_inv_1 _1616_ (.Y(_0614_),
    .A(net569));
 sg13g2_inv_4 _1617_ (.A(net564),
    .Y(_0622_));
 sg13g2_inv_4 _1618_ (.A(net635),
    .Y(_0629_));
 sg13g2_inv_2 _1619_ (.Y(_0639_),
    .A(net643));
 sg13g2_inv_1 _1620_ (.Y(_0648_),
    .A(net587));
 sg13g2_inv_2 _1621_ (.Y(_0656_),
    .A(net669));
 sg13g2_inv_2 _1622_ (.Y(_0666_),
    .A(net593));
 sg13g2_inv_2 _1623_ (.Y(_0675_),
    .A(net600));
 sg13g2_inv_4 _1624_ (.A(net606),
    .Y(_0680_));
 sg13g2_inv_2 _1625_ (.Y(_0683_),
    .A(\counter[6] ));
 sg13g2_inv_1 _1626_ (.Y(_0688_),
    .A(net531));
 sg13g2_inv_1 _1627_ (.Y(_0697_),
    .A(\counter[4] ));
 sg13g2_inv_1 _1628_ (.Y(_0698_),
    .A(\counter[2] ));
 sg13g2_nor2_2 _1629_ (.A(_0458_),
    .B(_0491_),
    .Y(_0699_));
 sg13g2_nand2_2 _1630_ (.Y(_0700_),
    .A(net579),
    .B(net574));
 sg13g2_nand2_1 _1631_ (.Y(_0701_),
    .A(net579),
    .B(_0699_));
 sg13g2_inv_1 _1632_ (.Y(_0702_),
    .A(_0701_));
 sg13g2_nand2_1 _1633_ (.Y(_0703_),
    .A(net567),
    .B(_0502_));
 sg13g2_nor2_2 _1634_ (.A(net552),
    .B(net588),
    .Y(_0704_));
 sg13g2_nand4_1 _1635_ (.B(net597),
    .C(net554),
    .A(net608),
    .Y(_0705_),
    .D(_0704_));
 sg13g2_nor3_1 _1636_ (.A(net562),
    .B(_0701_),
    .C(_0705_),
    .Y(_0011_));
 sg13g2_nand2_2 _1637_ (.Y(_0706_),
    .A(net617),
    .B(net626));
 sg13g2_nor2_2 _1638_ (.A(_0513_),
    .B(_0557_),
    .Y(_0707_));
 sg13g2_nor2_2 _1639_ (.A(net637),
    .B(net655),
    .Y(_0708_));
 sg13g2_nor2_1 _1640_ (.A(net639),
    .B(net647),
    .Y(_0709_));
 sg13g2_nand2_1 _1641_ (.Y(_0710_),
    .A(net545),
    .B(_0577_));
 sg13g2_o21ai_1 _1642_ (.B1(_0707_),
    .Y(_0711_),
    .A1(net656),
    .A2(_0710_));
 sg13g2_nor2_2 _1643_ (.A(_0577_),
    .B(net543),
    .Y(_0712_));
 sg13g2_nand2_2 _1644_ (.Y(_0713_),
    .A(net645),
    .B(net652));
 sg13g2_nand2_1 _1645_ (.Y(_0714_),
    .A(net632),
    .B(net641));
 sg13g2_or2_2 _1646_ (.X(_0715_),
    .B(_0714_),
    .A(_0713_));
 sg13g2_nor2_1 _1647_ (.A(_0513_),
    .B(net626),
    .Y(_0716_));
 sg13g2_a21oi_1 _1648_ (.A1(_0715_),
    .A2(_0716_),
    .Y(_0717_),
    .B1(net615));
 sg13g2_a21oi_2 _1649_ (.B1(_0717_),
    .Y(_0010_),
    .A2(_0711_),
    .A1(_0706_));
 sg13g2_nor2_1 _1650_ (.A(net627),
    .B(net632),
    .Y(_0718_));
 sg13g2_a21oi_1 _1651_ (.A1(net586),
    .A2(_0702_),
    .Y(_0719_),
    .B1(net560));
 sg13g2_o21ai_1 _1652_ (.B1(_0719_),
    .Y(_0720_),
    .A1(net616),
    .A2(_0718_));
 sg13g2_and2_2 _1653_ (.A(net624),
    .B(net639),
    .X(_0721_));
 sg13g2_nor2_1 _1654_ (.A(net617),
    .B(net630),
    .Y(_0722_));
 sg13g2_nor2_1 _1655_ (.A(_0707_),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_nand2_1 _1656_ (.Y(_0724_),
    .A(_0721_),
    .B(_0723_));
 sg13g2_nor2_1 _1657_ (.A(net630),
    .B(net647),
    .Y(_0725_));
 sg13g2_nor2_2 _1658_ (.A(net626),
    .B(net641),
    .Y(_0726_));
 sg13g2_nor3_1 _1659_ (.A(_0721_),
    .B(_0725_),
    .C(_0726_),
    .Y(_0727_));
 sg13g2_xnor2_1 _1660_ (.Y(_0728_),
    .A(net630),
    .B(net647));
 sg13g2_nand2b_1 _1661_ (.Y(_0729_),
    .B(_0728_),
    .A_N(_0708_));
 sg13g2_xnor2_1 _1662_ (.Y(_0730_),
    .A(_0708_),
    .B(_0728_));
 sg13g2_nand2_1 _1663_ (.Y(_0731_),
    .A(net546),
    .B(net655));
 sg13g2_nor2_1 _1664_ (.A(net545),
    .B(net655),
    .Y(_0732_));
 sg13g2_xnor2_1 _1665_ (.Y(_0733_),
    .A(net637),
    .B(net655));
 sg13g2_nand2_1 _1666_ (.Y(_0734_),
    .A(net666),
    .B(net647));
 sg13g2_nor2_1 _1667_ (.A(net666),
    .B(net644),
    .Y(_0735_));
 sg13g2_xor2_1 _1668_ (.B(net645),
    .A(net666),
    .X(_0736_));
 sg13g2_nor2_2 _1669_ (.A(net677),
    .B(net655),
    .Y(_0737_));
 sg13g2_o21ai_1 _1670_ (.B1(_0734_),
    .Y(_0738_),
    .A1(_0735_),
    .A2(_0737_));
 sg13g2_nand3_1 _1671_ (.B(_0733_),
    .C(_0738_),
    .A(_0730_),
    .Y(_0739_));
 sg13g2_o21ai_1 _1672_ (.B1(_0725_),
    .Y(_0740_),
    .A1(_0721_),
    .A2(_0726_));
 sg13g2_nand2b_1 _1673_ (.Y(_0741_),
    .B(_0740_),
    .A_N(_0727_));
 sg13g2_a21oi_1 _1674_ (.A1(_0729_),
    .A2(_0739_),
    .Y(_0742_),
    .B1(_0741_));
 sg13g2_xor2_1 _1675_ (.B(_0723_),
    .A(_0721_),
    .X(_0743_));
 sg13g2_o21ai_1 _1676_ (.B1(_0743_),
    .Y(_0744_),
    .A1(_0727_),
    .A2(_0742_));
 sg13g2_nand2_1 _1677_ (.Y(_0745_),
    .A(_0724_),
    .B(_0744_));
 sg13g2_xnor2_1 _1678_ (.Y(_0746_),
    .A(net620),
    .B(_0707_));
 sg13g2_nand2_1 _1679_ (.Y(_0747_),
    .A(_0745_),
    .B(_0746_));
 sg13g2_nand3_1 _1680_ (.B(_0622_),
    .C(_0747_),
    .A(_0513_),
    .Y(_0748_));
 sg13g2_nand3b_1 _1681_ (.B(_0745_),
    .C(net563),
    .Y(_0749_),
    .A_N(net620));
 sg13g2_nand3_1 _1682_ (.B(_0739_),
    .C(_0741_),
    .A(_0729_),
    .Y(_0750_));
 sg13g2_nor2b_1 _1683_ (.A(_0742_),
    .B_N(_0750_),
    .Y(_0751_));
 sg13g2_xnor2_1 _1684_ (.Y(_0752_),
    .A(_0038_),
    .B(_0751_));
 sg13g2_a21o_1 _1685_ (.A2(_0738_),
    .A1(_0733_),
    .B1(_0730_),
    .X(_0753_));
 sg13g2_and2_1 _1686_ (.A(_0739_),
    .B(_0753_),
    .X(_0754_));
 sg13g2_xnor2_1 _1687_ (.Y(_0755_),
    .A(net593),
    .B(_0754_));
 sg13g2_xor2_1 _1688_ (.B(_0738_),
    .A(_0733_),
    .X(_0756_));
 sg13g2_and2_1 _1689_ (.A(net601),
    .B(_0756_),
    .X(_0757_));
 sg13g2_xnor2_1 _1690_ (.Y(_0758_),
    .A(_0736_),
    .B(_0737_));
 sg13g2_nand2_2 _1691_ (.Y(_0759_),
    .A(net677),
    .B(net655));
 sg13g2_nand2b_2 _1692_ (.Y(_0760_),
    .B(_0759_),
    .A_N(_0737_));
 sg13g2_o21ai_1 _1693_ (.B1(_0502_),
    .Y(_0761_),
    .A1(net556),
    .A2(_0760_));
 sg13g2_a21oi_2 _1694_ (.B1(_0761_),
    .Y(_0762_),
    .A2(_0760_),
    .A1(_0414_));
 sg13g2_o21ai_1 _1695_ (.B1(_0762_),
    .Y(_0763_),
    .A1(net606),
    .A2(_0758_));
 sg13g2_a221oi_1 _1696_ (.B2(_0758_),
    .C1(_0763_),
    .B1(net606),
    .A1(net619),
    .Y(_0764_),
    .A2(net566));
 sg13g2_o21ai_1 _1697_ (.B1(_0764_),
    .Y(_0765_),
    .A1(net601),
    .A2(_0756_));
 sg13g2_nor4_1 _1698_ (.A(_0752_),
    .B(_0755_),
    .C(_0757_),
    .D(_0765_),
    .Y(_0766_));
 sg13g2_or3_1 _1699_ (.A(_0727_),
    .B(_0742_),
    .C(_0743_),
    .X(_0767_));
 sg13g2_and2_1 _1700_ (.A(_0744_),
    .B(_0767_),
    .X(_0768_));
 sg13g2_xor2_1 _1701_ (.B(_0768_),
    .A(net582),
    .X(_0769_));
 sg13g2_nand4_1 _1702_ (.B(_0749_),
    .C(_0766_),
    .A(_0748_),
    .Y(_0770_),
    .D(_0769_));
 sg13g2_nand2_2 _1703_ (.Y(_0771_),
    .A(net625),
    .B(net631));
 sg13g2_o21ai_1 _1704_ (.B1(_0747_),
    .Y(_0772_),
    .A1(_0513_),
    .A2(_0771_));
 sg13g2_xor2_1 _1705_ (.B(net569),
    .A(net615),
    .X(_0773_));
 sg13g2_xor2_1 _1706_ (.B(_0746_),
    .A(_0745_),
    .X(_0774_));
 sg13g2_xnor2_1 _1707_ (.Y(_0775_),
    .A(_0772_),
    .B(_0773_));
 sg13g2_xnor2_1 _1708_ (.Y(_0776_),
    .A(net576),
    .B(_0774_));
 sg13g2_nor3_1 _1709_ (.A(_0770_),
    .B(_0775_),
    .C(_0776_),
    .Y(_0777_));
 sg13g2_nand2_1 _1710_ (.Y(_0778_),
    .A(_0557_),
    .B(net639));
 sg13g2_o21ai_1 _1711_ (.B1(_0778_),
    .Y(_0779_),
    .A1(net639),
    .A2(_0728_));
 sg13g2_xor2_1 _1712_ (.B(_0779_),
    .A(net575),
    .X(_0780_));
 sg13g2_xnor2_1 _1713_ (.Y(_0781_),
    .A(net619),
    .B(net566));
 sg13g2_nor3_2 _1714_ (.A(net630),
    .B(net639),
    .C(net647),
    .Y(_0782_));
 sg13g2_xor2_1 _1715_ (.B(net620),
    .A(net569),
    .X(_0783_));
 sg13g2_a221oi_1 _1716_ (.B2(net624),
    .C1(_0783_),
    .B1(_0781_),
    .A1(net546),
    .Y(_0784_),
    .A2(_0725_));
 sg13g2_nand3_1 _1717_ (.B(_0782_),
    .C(_0783_),
    .A(_0781_),
    .Y(_0785_));
 sg13g2_nand2b_1 _1718_ (.Y(_0786_),
    .B(_0785_),
    .A_N(_0784_));
 sg13g2_xor2_1 _1719_ (.B(net656),
    .A(net598),
    .X(_0787_));
 sg13g2_xnor2_1 _1720_ (.Y(_0788_),
    .A(net589),
    .B(net649));
 sg13g2_xnor2_1 _1721_ (.Y(_0789_),
    .A(net613),
    .B(net684));
 sg13g2_xor2_1 _1722_ (.B(net682),
    .A(net613),
    .X(_0790_));
 sg13g2_xor2_1 _1723_ (.B(net667),
    .A(net604),
    .X(_0791_));
 sg13g2_nand4_1 _1724_ (.B(_0788_),
    .C(_0790_),
    .A(_0787_),
    .Y(_0792_),
    .D(_0791_));
 sg13g2_a21oi_1 _1725_ (.A1(net624),
    .A2(net615),
    .Y(_0793_),
    .B1(_0781_));
 sg13g2_xnor2_1 _1726_ (.Y(_0794_),
    .A(net608),
    .B(net676));
 sg13g2_nor4_1 _1727_ (.A(net562),
    .B(_0792_),
    .C(_0793_),
    .D(_0794_),
    .Y(_0795_));
 sg13g2_nand3_1 _1728_ (.B(_0786_),
    .C(_0795_),
    .A(_0780_),
    .Y(_0796_));
 sg13g2_a21oi_1 _1729_ (.A1(net639),
    .A2(net647),
    .Y(_0797_),
    .B1(net630));
 sg13g2_or2_1 _1730_ (.X(_0798_),
    .B(_0797_),
    .A(_0706_));
 sg13g2_xnor2_1 _1731_ (.Y(_0799_),
    .A(net561),
    .B(_0798_));
 sg13g2_nor2_1 _1732_ (.A(net546),
    .B(_0728_),
    .Y(_0800_));
 sg13g2_a21oi_1 _1733_ (.A1(net630),
    .A2(net546),
    .Y(_0801_),
    .B1(_0800_));
 sg13g2_nor2_2 _1734_ (.A(net617),
    .B(net626),
    .Y(_0802_));
 sg13g2_nand2_2 _1735_ (.Y(_0803_),
    .A(net639),
    .B(net647));
 sg13g2_a21oi_1 _1736_ (.A1(_0722_),
    .A2(_0803_),
    .Y(_0804_),
    .B1(_0802_));
 sg13g2_a21oi_1 _1737_ (.A1(_0798_),
    .A2(_0804_),
    .Y(_0805_),
    .B1(net563));
 sg13g2_a21o_1 _1738_ (.A2(_0801_),
    .A1(net575),
    .B1(_0805_),
    .X(_0806_));
 sg13g2_nand2_1 _1739_ (.Y(_0807_),
    .A(net628),
    .B(_0803_));
 sg13g2_xnor2_1 _1740_ (.Y(_0808_),
    .A(net624),
    .B(net570));
 sg13g2_xnor2_1 _1741_ (.Y(_0809_),
    .A(_0807_),
    .B(_0808_));
 sg13g2_nor3_1 _1742_ (.A(_0787_),
    .B(_0788_),
    .C(_0791_),
    .Y(_0810_));
 sg13g2_nand4_1 _1743_ (.B(_0794_),
    .C(_0809_),
    .A(_0789_),
    .Y(_0811_),
    .D(_0810_));
 sg13g2_nand3_1 _1744_ (.B(_0798_),
    .C(_0804_),
    .A(net563),
    .Y(_0812_));
 sg13g2_o21ai_1 _1745_ (.B1(_0812_),
    .Y(_0813_),
    .A1(net575),
    .A2(_0801_));
 sg13g2_or4_1 _1746_ (.A(_0799_),
    .B(_0806_),
    .C(_0811_),
    .D(_0813_),
    .X(_0814_));
 sg13g2_nor2b_1 _1747_ (.A(_0709_),
    .B_N(_0803_),
    .Y(_0815_));
 sg13g2_xnor2_1 _1748_ (.Y(_0816_),
    .A(net582),
    .B(_0815_));
 sg13g2_a21oi_1 _1749_ (.A1(_0796_),
    .A2(_0814_),
    .Y(_0817_),
    .B1(_0816_));
 sg13g2_nor2_2 _1750_ (.A(net685),
    .B(net680),
    .Y(_0818_));
 sg13g2_or2_2 _1751_ (.X(_0819_),
    .B(net680),
    .A(net686));
 sg13g2_nor3_2 _1752_ (.A(net688),
    .B(net676),
    .C(net682),
    .Y(_0820_));
 sg13g2_nor2_2 _1753_ (.A(net667),
    .B(net654),
    .Y(_0821_));
 sg13g2_nor3_2 _1754_ (.A(net667),
    .B(net649),
    .C(net656),
    .Y(_0822_));
 sg13g2_nor4_2 _1755_ (.A(net689),
    .B(net666),
    .C(net676),
    .Y(_0823_),
    .D(net682));
 sg13g2_nand2_2 _1756_ (.Y(_0824_),
    .A(net550),
    .B(_0820_));
 sg13g2_nor2_1 _1757_ (.A(net645),
    .B(net655),
    .Y(_0825_));
 sg13g2_or2_2 _1758_ (.X(_0826_),
    .B(net656),
    .A(net648));
 sg13g2_nand4_1 _1759_ (.B(_0722_),
    .C(_0823_),
    .A(_0721_),
    .Y(_0827_),
    .D(net539));
 sg13g2_nor2b_2 _1760_ (.A(net653),
    .B_N(net645),
    .Y(_0828_));
 sg13g2_nand2b_2 _1761_ (.Y(_0829_),
    .B(net645),
    .A_N(net653));
 sg13g2_nor2b_2 _1762_ (.A(net644),
    .B_N(net652),
    .Y(_0830_));
 sg13g2_nand2b_2 _1763_ (.Y(_0831_),
    .B(net653),
    .A_N(net645));
 sg13g2_nand2_2 _1764_ (.Y(_0832_),
    .A(_0829_),
    .B(_0831_));
 sg13g2_xnor2_1 _1765_ (.Y(_0833_),
    .A(net582),
    .B(_0832_));
 sg13g2_xnor2_1 _1766_ (.Y(_0834_),
    .A(net565),
    .B(net621));
 sg13g2_xor2_1 _1767_ (.B(net620),
    .A(net563),
    .X(_0835_));
 sg13g2_o21ai_1 _1768_ (.B1(net628),
    .Y(_0836_),
    .A1(_0778_),
    .A2(net538));
 sg13g2_o21ai_1 _1769_ (.B1(_0833_),
    .Y(_0837_),
    .A1(_0835_),
    .A2(_0836_));
 sg13g2_nand2_2 _1770_ (.Y(_0838_),
    .A(net640),
    .B(_0826_));
 sg13g2_a22oi_1 _1771_ (.Y(_0839_),
    .B1(_0826_),
    .B2(net639),
    .A2(_0709_),
    .A1(net544));
 sg13g2_xnor2_1 _1772_ (.Y(_0840_),
    .A(net630),
    .B(net569));
 sg13g2_xnor2_1 _1773_ (.Y(_0841_),
    .A(_0838_),
    .B(_0840_));
 sg13g2_o21ai_1 _1774_ (.B1(_0841_),
    .Y(_0842_),
    .A1(net575),
    .A2(_0839_));
 sg13g2_or2_1 _1775_ (.X(_0843_),
    .B(_0842_),
    .A(_0837_));
 sg13g2_xor2_1 _1776_ (.B(_0028_),
    .A(net616),
    .X(_0844_));
 sg13g2_nor2_1 _1777_ (.A(net625),
    .B(net537),
    .Y(_0845_));
 sg13g2_o21ai_1 _1778_ (.B1(_0835_),
    .Y(_0846_),
    .A1(_0836_),
    .A2(_0845_));
 sg13g2_nand2_2 _1779_ (.Y(_0847_),
    .A(net608),
    .B(net682));
 sg13g2_nand2_1 _1780_ (.Y(_0848_),
    .A(_0425_),
    .B(_0546_));
 sg13g2_nand2_2 _1781_ (.Y(_0849_),
    .A(_0847_),
    .B(_0848_));
 sg13g2_nor2_1 _1782_ (.A(net689),
    .B(net613),
    .Y(_0850_));
 sg13g2_nand2_1 _1783_ (.Y(_0851_),
    .A(_0403_),
    .B(_0414_));
 sg13g2_xnor2_1 _1784_ (.Y(_0852_),
    .A(net689),
    .B(net613));
 sg13g2_xor2_1 _1785_ (.B(net656),
    .A(net589),
    .X(_0853_));
 sg13g2_nand2b_1 _1786_ (.Y(_0854_),
    .B(net667),
    .A_N(net598));
 sg13g2_nand2b_1 _1787_ (.Y(_0855_),
    .B(net598),
    .A_N(net667));
 sg13g2_and2_1 _1788_ (.A(_0854_),
    .B(_0855_),
    .X(_0856_));
 sg13g2_xnor2_1 _1789_ (.Y(_0857_),
    .A(net604),
    .B(net678));
 sg13g2_and2_1 _1790_ (.A(net526),
    .B(_0857_),
    .X(_0858_));
 sg13g2_nand4_1 _1791_ (.B(_0852_),
    .C(_0853_),
    .A(_0849_),
    .Y(_0859_),
    .D(_0858_));
 sg13g2_nand2_1 _1792_ (.Y(_0860_),
    .A(_0716_),
    .B(_0835_));
 sg13g2_a221oi_1 _1793_ (.B2(_0860_),
    .C1(_0859_),
    .B1(net537),
    .A1(net575),
    .Y(_0861_),
    .A2(_0839_));
 sg13g2_nand2_1 _1794_ (.Y(_0862_),
    .A(_0846_),
    .B(_0861_));
 sg13g2_o21ai_1 _1795_ (.B1(_0827_),
    .Y(_0863_),
    .A1(_0843_),
    .A2(_0862_));
 sg13g2_nor3_2 _1796_ (.A(net631),
    .B(net640),
    .C(_0712_),
    .Y(_0864_));
 sg13g2_nor2b_1 _1797_ (.A(net625),
    .B_N(_0864_),
    .Y(_0865_));
 sg13g2_nor3_1 _1798_ (.A(net617),
    .B(net537),
    .C(_0865_),
    .Y(_0866_));
 sg13g2_a21oi_1 _1799_ (.A1(net537),
    .A2(_0865_),
    .Y(_0867_),
    .B1(_0866_));
 sg13g2_xnor2_1 _1800_ (.Y(_0868_),
    .A(net634),
    .B(_0713_));
 sg13g2_xor2_1 _1801_ (.B(_0868_),
    .A(net576),
    .X(_0869_));
 sg13g2_xnor2_1 _1802_ (.Y(_0870_),
    .A(net625),
    .B(_0864_));
 sg13g2_xnor2_1 _1803_ (.Y(_0871_),
    .A(net563),
    .B(_0870_));
 sg13g2_a21oi_1 _1804_ (.A1(net634),
    .A2(_0713_),
    .Y(_0872_),
    .B1(_0840_));
 sg13g2_nand3_1 _1805_ (.B(_0713_),
    .C(_0840_),
    .A(net634),
    .Y(_0873_));
 sg13g2_nor3_1 _1806_ (.A(_0853_),
    .B(_0856_),
    .C(_0872_),
    .Y(_0874_));
 sg13g2_nor3_2 _1807_ (.A(_0849_),
    .B(_0852_),
    .C(_0857_),
    .Y(_0875_));
 sg13g2_nand4_1 _1808_ (.B(_0873_),
    .C(_0874_),
    .A(_0833_),
    .Y(_0876_),
    .D(_0875_));
 sg13g2_nor4_1 _1809_ (.A(_0867_),
    .B(_0869_),
    .C(_0871_),
    .D(_0876_),
    .Y(_0877_));
 sg13g2_nor4_2 _1810_ (.A(_0777_),
    .B(_0817_),
    .C(_0863_),
    .Y(_0878_),
    .D(_0877_));
 sg13g2_nor2_1 _1811_ (.A(net634),
    .B(net539),
    .Y(_0879_));
 sg13g2_xnor2_1 _1812_ (.Y(_0880_),
    .A(net628),
    .B(_0879_));
 sg13g2_nand2_1 _1813_ (.Y(_0881_),
    .A(net615),
    .B(_0880_));
 sg13g2_and2_1 _1814_ (.A(net628),
    .B(_0832_),
    .X(_0882_));
 sg13g2_xor2_1 _1815_ (.B(_0832_),
    .A(net628),
    .X(_0883_));
 sg13g2_a21oi_1 _1816_ (.A1(_0734_),
    .A2(_0759_),
    .Y(_0884_),
    .B1(_0735_));
 sg13g2_o21ai_1 _1817_ (.B1(_0731_),
    .Y(_0885_),
    .A1(_0732_),
    .A2(_0884_));
 sg13g2_a21oi_1 _1818_ (.A1(_0883_),
    .A2(_0885_),
    .Y(_0886_),
    .B1(_0882_));
 sg13g2_xnor2_1 _1819_ (.Y(_0887_),
    .A(net620),
    .B(_0839_));
 sg13g2_nor2b_1 _1820_ (.A(_0886_),
    .B_N(_0887_),
    .Y(_0888_));
 sg13g2_nor2_1 _1821_ (.A(net624),
    .B(_0839_),
    .Y(_0889_));
 sg13g2_nor2_1 _1822_ (.A(_0888_),
    .B(_0889_),
    .Y(_0890_));
 sg13g2_xnor2_1 _1823_ (.Y(_0891_),
    .A(_0597_),
    .B(_0880_));
 sg13g2_o21ai_1 _1824_ (.B1(_0891_),
    .Y(_0892_),
    .A1(_0888_),
    .A2(_0889_));
 sg13g2_nand2_2 _1825_ (.Y(_0893_),
    .A(_0881_),
    .B(_0892_));
 sg13g2_nand2_1 _1826_ (.Y(_0894_),
    .A(_0557_),
    .B(_0838_));
 sg13g2_xor2_1 _1827_ (.B(_0894_),
    .A(net625),
    .X(_0895_));
 sg13g2_inv_1 _1828_ (.Y(_0896_),
    .A(_0895_));
 sg13g2_a21oi_1 _1829_ (.A1(_0557_),
    .A2(_0838_),
    .Y(_0897_),
    .B1(net620));
 sg13g2_xnor2_1 _1830_ (.Y(_0898_),
    .A(net615),
    .B(_0897_));
 sg13g2_nor3_1 _1831_ (.A(_0893_),
    .B(_0896_),
    .C(_0898_),
    .Y(_0899_));
 sg13g2_o21ai_1 _1832_ (.B1(_0898_),
    .Y(_0900_),
    .A1(_0893_),
    .A2(_0896_));
 sg13g2_nor2b_1 _1833_ (.A(_0899_),
    .B_N(_0900_),
    .Y(_0901_));
 sg13g2_xnor2_1 _1834_ (.Y(_0902_),
    .A(net569),
    .B(_0901_));
 sg13g2_a21oi_1 _1835_ (.A1(net625),
    .A2(_0894_),
    .Y(_0903_),
    .B1(net617));
 sg13g2_nor2b_1 _1836_ (.A(_0899_),
    .B_N(_0903_),
    .Y(_0904_));
 sg13g2_xnor2_1 _1837_ (.Y(_0905_),
    .A(_0622_),
    .B(_0904_));
 sg13g2_xnor2_1 _1838_ (.Y(_0906_),
    .A(_0893_),
    .B(_0895_));
 sg13g2_nor2b_1 _1839_ (.A(net576),
    .B_N(_0906_),
    .Y(_0907_));
 sg13g2_xnor2_1 _1840_ (.Y(_0908_),
    .A(_0890_),
    .B(_0891_));
 sg13g2_nand2_1 _1841_ (.Y(_0909_),
    .A(net582),
    .B(_0908_));
 sg13g2_or2_1 _1842_ (.X(_0910_),
    .B(_0908_),
    .A(net582));
 sg13g2_xnor2_1 _1843_ (.Y(_0911_),
    .A(_0886_),
    .B(_0887_));
 sg13g2_nor2_1 _1844_ (.A(_0038_),
    .B(_0911_),
    .Y(_0912_));
 sg13g2_xor2_1 _1845_ (.B(_0885_),
    .A(_0883_),
    .X(_0913_));
 sg13g2_nor2_1 _1846_ (.A(net593),
    .B(_0913_),
    .Y(_0914_));
 sg13g2_xnor2_1 _1847_ (.Y(_0915_),
    .A(_0733_),
    .B(_0884_));
 sg13g2_xor2_1 _1848_ (.B(_0759_),
    .A(_0736_),
    .X(_0916_));
 sg13g2_xnor2_1 _1849_ (.Y(_0917_),
    .A(_0680_),
    .B(_0916_));
 sg13g2_nand2_1 _1850_ (.Y(_0918_),
    .A(_0762_),
    .B(_0917_));
 sg13g2_nor3_1 _1851_ (.A(_0912_),
    .B(_0914_),
    .C(_0918_),
    .Y(_0919_));
 sg13g2_xnor2_1 _1852_ (.Y(_0920_),
    .A(net601),
    .B(_0915_));
 sg13g2_a221oi_1 _1853_ (.B2(net593),
    .C1(_0920_),
    .B1(_0913_),
    .A1(_0038_),
    .Y(_0921_),
    .A2(_0911_));
 sg13g2_nand4_1 _1854_ (.B(_0910_),
    .C(_0919_),
    .A(_0909_),
    .Y(_0922_),
    .D(_0921_));
 sg13g2_nor2b_1 _1855_ (.A(_0903_),
    .B_N(_0899_),
    .Y(_0923_));
 sg13g2_nor2b_1 _1856_ (.A(_0906_),
    .B_N(net576),
    .Y(_0924_));
 sg13g2_nor4_1 _1857_ (.A(_0907_),
    .B(_0922_),
    .C(_0923_),
    .D(_0924_),
    .Y(_0925_));
 sg13g2_nand3_1 _1858_ (.B(_0905_),
    .C(_0925_),
    .A(_0902_),
    .Y(_0926_));
 sg13g2_nor2_2 _1859_ (.A(net568),
    .B(net560),
    .Y(_0927_));
 sg13g2_nor2_2 _1860_ (.A(net552),
    .B(_0480_),
    .Y(_0928_));
 sg13g2_nand2_2 _1861_ (.Y(_0929_),
    .A(net585),
    .B(net588));
 sg13g2_nor2_2 _1862_ (.A(net611),
    .B(net607),
    .Y(_0930_));
 sg13g2_nor4_2 _1863_ (.A(net614),
    .B(net608),
    .C(net596),
    .Y(_0931_),
    .D(net603));
 sg13g2_nor2_2 _1864_ (.A(net581),
    .B(net571),
    .Y(_0932_));
 sg13g2_o21ai_1 _1865_ (.B1(_0932_),
    .Y(_0933_),
    .A1(_0929_),
    .A2(_0931_));
 sg13g2_nand2_1 _1866_ (.Y(_0934_),
    .A(net567),
    .B(_0933_));
 sg13g2_a22oi_1 _1867_ (.Y(_0935_),
    .B1(_0934_),
    .B2(_0502_),
    .A2(_0926_),
    .A1(_0878_));
 sg13g2_nor2_1 _1868_ (.A(_0447_),
    .B(net571),
    .Y(_0936_));
 sg13g2_nand2_2 _1869_ (.Y(_0937_),
    .A(net614),
    .B(net609));
 sg13g2_inv_1 _1870_ (.Y(_0938_),
    .A(_0937_));
 sg13g2_nand3_1 _1871_ (.B(net607),
    .C(net603),
    .A(net611),
    .Y(_0939_));
 sg13g2_nand2_2 _1872_ (.Y(_0940_),
    .A(net595),
    .B(net603));
 sg13g2_or2_1 _1873_ (.X(_0941_),
    .B(_0940_),
    .A(_0937_));
 sg13g2_a21oi_1 _1874_ (.A1(_0704_),
    .A2(net524),
    .Y(_0942_),
    .B1(net584));
 sg13g2_nor2b_1 _1875_ (.A(_0942_),
    .B_N(_0936_),
    .Y(_0943_));
 sg13g2_or2_2 _1876_ (.X(_0944_),
    .B(net532),
    .A(\counter[4] ));
 sg13g2_or2_2 _1877_ (.X(_0945_),
    .B(\counter[1] ),
    .A(net533));
 sg13g2_o21ai_1 _1878_ (.B1(net530),
    .Y(_0946_),
    .A1(_0944_),
    .A2(_0945_));
 sg13g2_xnor2_1 _1879_ (.Y(_0947_),
    .A(_0683_),
    .B(_0946_));
 sg13g2_o21ai_1 _1880_ (.B1(_0022_),
    .Y(_0948_),
    .A1(\counter[6] ),
    .A2(_0946_));
 sg13g2_o21ai_1 _1881_ (.B1(_0948_),
    .Y(_0949_),
    .A1(net581),
    .A2(net570));
 sg13g2_nor2_2 _1882_ (.A(net530),
    .B(\counter[4] ),
    .Y(_0950_));
 sg13g2_nand2b_1 _1883_ (.Y(_0951_),
    .B(_0950_),
    .A_N(net532));
 sg13g2_o21ai_1 _1884_ (.B1(_0946_),
    .Y(_0952_),
    .A1(_0945_),
    .A2(_0951_));
 sg13g2_xnor2_1 _1885_ (.Y(_0953_),
    .A(net542),
    .B(_0952_));
 sg13g2_nor2_1 _1886_ (.A(\counter[3] ),
    .B(net533),
    .Y(_0954_));
 sg13g2_nor2_1 _1887_ (.A(\counter[3] ),
    .B(_0945_),
    .Y(_0955_));
 sg13g2_xor2_1 _1888_ (.B(_0025_),
    .A(net602),
    .X(_0956_));
 sg13g2_xor2_1 _1889_ (.B(_0024_),
    .A(net592),
    .X(_0957_));
 sg13g2_xnor2_1 _1890_ (.Y(_0958_),
    .A(net611),
    .B(\counter[1] ));
 sg13g2_nand2_1 _1891_ (.Y(_0959_),
    .A(net533),
    .B(\counter[1] ));
 sg13g2_a21oi_1 _1892_ (.A1(_0945_),
    .A2(_0959_),
    .Y(_0960_),
    .B1(_0680_));
 sg13g2_nand2_1 _1893_ (.Y(_0961_),
    .A(net606),
    .B(_0945_));
 sg13g2_and2_1 _1894_ (.A(_0959_),
    .B(_0961_),
    .X(_0962_));
 sg13g2_nor2b_1 _1895_ (.A(_0956_),
    .B_N(_0962_),
    .Y(_0963_));
 sg13g2_xnor2_1 _1896_ (.Y(_0964_),
    .A(_0955_),
    .B(_0957_));
 sg13g2_a21oi_1 _1897_ (.A1(net581),
    .A2(net570),
    .Y(_0965_),
    .B1(_0948_));
 sg13g2_xor2_1 _1898_ (.B(_0022_),
    .A(net592),
    .X(_0966_));
 sg13g2_xnor2_1 _1899_ (.Y(_0967_),
    .A(_0951_),
    .B(_0966_));
 sg13g2_nand2_1 _1900_ (.Y(_0968_),
    .A(_0683_),
    .B(_0688_));
 sg13g2_nor2_1 _1901_ (.A(_0944_),
    .B(_0968_),
    .Y(_0969_));
 sg13g2_nor2_1 _1902_ (.A(net585),
    .B(net591),
    .Y(_0970_));
 sg13g2_or2_2 _1903_ (.X(_0971_),
    .B(net588),
    .A(net585));
 sg13g2_and3_1 _1904_ (.X(_0972_),
    .A(_0928_),
    .B(_0932_),
    .C(net524));
 sg13g2_nand2_1 _1905_ (.Y(_0973_),
    .A(\counter[4] ),
    .B(net532));
 sg13g2_nand3_1 _1906_ (.B(_0944_),
    .C(_0973_),
    .A(_0680_),
    .Y(_0974_));
 sg13g2_nor2_2 _1907_ (.A(net578),
    .B(net536),
    .Y(_0975_));
 sg13g2_a21oi_1 _1908_ (.A1(_0944_),
    .A2(_0973_),
    .Y(_0976_),
    .B1(_0680_));
 sg13g2_xor2_1 _1909_ (.B(_0023_),
    .A(net602),
    .X(_0977_));
 sg13g2_xor2_1 _1910_ (.B(net532),
    .A(net611),
    .X(_0978_));
 sg13g2_nand2_1 _1911_ (.Y(_0979_),
    .A(net578),
    .B(net536));
 sg13g2_nor3_1 _1912_ (.A(_0932_),
    .B(_0969_),
    .C(_0971_),
    .Y(_0980_));
 sg13g2_a21oi_1 _1913_ (.A1(_0928_),
    .A2(_0969_),
    .Y(_0981_),
    .B1(_0980_));
 sg13g2_xnor2_1 _1914_ (.Y(_0982_),
    .A(net571),
    .B(_0975_));
 sg13g2_nand3_1 _1915_ (.B(_0978_),
    .C(_0982_),
    .A(_0974_),
    .Y(_0983_));
 sg13g2_nor2b_2 _1916_ (.A(_0975_),
    .B_N(_0979_),
    .Y(_0984_));
 sg13g2_nand2b_2 _1917_ (.Y(_0985_),
    .B(_0979_),
    .A_N(_0975_));
 sg13g2_or4_1 _1918_ (.A(_0967_),
    .B(_0972_),
    .C(_0976_),
    .D(_0985_),
    .X(_0986_));
 sg13g2_xnor2_1 _1919_ (.Y(_0987_),
    .A(_0944_),
    .B(_0977_));
 sg13g2_nor4_1 _1920_ (.A(_0981_),
    .B(_0983_),
    .C(_0986_),
    .D(_0987_),
    .Y(_0988_));
 sg13g2_xor2_1 _1921_ (.B(net533),
    .A(net532),
    .X(_0989_));
 sg13g2_nor2_1 _1922_ (.A(net533),
    .B(_0944_),
    .Y(_0990_));
 sg13g2_xor2_1 _1923_ (.B(_0023_),
    .A(net592),
    .X(_0991_));
 sg13g2_xor2_1 _1924_ (.B(_0024_),
    .A(net602),
    .X(_0992_));
 sg13g2_o21ai_1 _1925_ (.B1(_0936_),
    .Y(_0993_),
    .A1(net556),
    .A2(_0698_));
 sg13g2_a21oi_1 _1926_ (.A1(_0950_),
    .A2(_0954_),
    .Y(_0994_),
    .B1(_0683_));
 sg13g2_a21oi_1 _1927_ (.A1(_0698_),
    .A2(_0969_),
    .Y(_0995_),
    .B1(_0994_));
 sg13g2_xnor2_1 _1928_ (.Y(_0996_),
    .A(net587),
    .B(_0995_));
 sg13g2_xnor2_1 _1929_ (.Y(_0997_),
    .A(net552),
    .B(_0994_));
 sg13g2_xnor2_1 _1930_ (.Y(_0998_),
    .A(net606),
    .B(_0989_));
 sg13g2_xnor2_1 _1931_ (.Y(_0999_),
    .A(_0990_),
    .B(_0991_));
 sg13g2_a22oi_1 _1932_ (.Y(_1000_),
    .B1(_0968_),
    .B2(net601),
    .A2(_0937_),
    .A1(_0436_));
 sg13g2_xor2_1 _1933_ (.B(net530),
    .A(\counter[6] ),
    .X(_1001_));
 sg13g2_o21ai_1 _1934_ (.B1(_1000_),
    .Y(_1002_),
    .A1(net614),
    .A2(net530));
 sg13g2_o21ai_1 _1935_ (.B1(_0688_),
    .Y(_1003_),
    .A1(net601),
    .A2(\counter[6] ));
 sg13g2_a21oi_1 _1936_ (.A1(net614),
    .A2(_1003_),
    .Y(_1004_),
    .B1(_1002_));
 sg13g2_xnor2_1 _1937_ (.Y(_1005_),
    .A(net606),
    .B(_1001_));
 sg13g2_nand2_1 _1938_ (.Y(_1006_),
    .A(net613),
    .B(\counter[6] ));
 sg13g2_a21oi_1 _1939_ (.A1(net608),
    .A2(_0683_),
    .Y(_1007_),
    .B1(net603));
 sg13g2_a22oi_1 _1940_ (.Y(_1008_),
    .B1(_1006_),
    .B2(_1007_),
    .A2(_1005_),
    .A1(_1004_));
 sg13g2_xnor2_1 _1941_ (.Y(_1009_),
    .A(net601),
    .B(_0022_));
 sg13g2_nand2_1 _1942_ (.Y(_1010_),
    .A(_0950_),
    .B(_1009_));
 sg13g2_a21oi_1 _1943_ (.A1(_0683_),
    .A2(_0950_),
    .Y(_1011_),
    .B1(net541));
 sg13g2_nand2b_2 _1944_ (.Y(_1012_),
    .B(_0939_),
    .A_N(net596));
 sg13g2_xor2_1 _1945_ (.B(\counter[4] ),
    .A(net530),
    .X(_1013_));
 sg13g2_xnor2_1 _1946_ (.Y(_1014_),
    .A(_0680_),
    .B(_1013_));
 sg13g2_o21ai_1 _1947_ (.B1(net614),
    .Y(_1015_),
    .A1(net592),
    .A2(_0968_));
 sg13g2_and2_1 _1948_ (.A(_0697_),
    .B(_1015_),
    .X(_1016_));
 sg13g2_nand2_1 _1949_ (.Y(_1017_),
    .A(net613),
    .B(\counter[4] ));
 sg13g2_a21oi_1 _1950_ (.A1(_1009_),
    .A2(_1017_),
    .Y(_1018_),
    .B1(_0950_));
 sg13g2_nor4_1 _1951_ (.A(_1011_),
    .B(_1014_),
    .C(_1016_),
    .D(_1018_),
    .Y(_1019_));
 sg13g2_nand3_1 _1952_ (.B(_1012_),
    .C(_1019_),
    .A(_1010_),
    .Y(_1020_));
 sg13g2_o21ai_1 _1953_ (.B1(_1020_),
    .Y(_1021_),
    .A1(net596),
    .A2(_1008_));
 sg13g2_nand3_1 _1954_ (.B(_0932_),
    .C(_1021_),
    .A(_0928_),
    .Y(_1022_));
 sg13g2_a221oi_1 _1955_ (.B2(_0970_),
    .C1(_0993_),
    .B1(net524),
    .A1(net556),
    .Y(_1023_),
    .A2(_0698_));
 sg13g2_xnor2_1 _1956_ (.Y(_1024_),
    .A(_0954_),
    .B(_0992_));
 sg13g2_nand4_1 _1957_ (.B(_0999_),
    .C(_1023_),
    .A(_0998_),
    .Y(_1025_),
    .D(_1024_));
 sg13g2_nor3_1 _1958_ (.A(_0996_),
    .B(_0997_),
    .C(_1025_),
    .Y(_1026_));
 sg13g2_nor4_1 _1959_ (.A(_0932_),
    .B(_0960_),
    .C(_0963_),
    .D(_0965_),
    .Y(_1027_));
 sg13g2_a21oi_1 _1960_ (.A1(_0945_),
    .A2(_0956_),
    .Y(_1028_),
    .B1(_0958_));
 sg13g2_nand4_1 _1961_ (.B(_0964_),
    .C(_1027_),
    .A(_0949_),
    .Y(_1029_),
    .D(_1028_));
 sg13g2_xnor2_1 _1962_ (.Y(_1030_),
    .A(net584),
    .B(_0947_));
 sg13g2_nor4_1 _1963_ (.A(_0943_),
    .B(_0953_),
    .C(_1029_),
    .D(_1030_),
    .Y(_1031_));
 sg13g2_nor3_1 _1964_ (.A(_0988_),
    .B(_1026_),
    .C(_1031_),
    .Y(_1032_));
 sg13g2_a21oi_1 _1965_ (.A1(_1022_),
    .A2(_1032_),
    .Y(_1033_),
    .B1(_0703_));
 sg13g2_nor2_2 _1966_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .Y(_1034_));
 sg13g2_nand2_2 _1967_ (.Y(_1035_),
    .A(_0698_),
    .B(_1034_));
 sg13g2_o21ai_1 _1968_ (.B1(\counter[4] ),
    .Y(_1036_),
    .A1(\counter[3] ),
    .A2(_1035_));
 sg13g2_o21ai_1 _1969_ (.B1(_0023_),
    .Y(_1037_),
    .A1(net531),
    .A2(_1036_));
 sg13g2_nand2b_1 _1970_ (.Y(_1038_),
    .B(_0683_),
    .A_N(_1037_));
 sg13g2_nand2_1 _1971_ (.Y(_1039_),
    .A(net578),
    .B(_1038_));
 sg13g2_nand2_1 _1972_ (.Y(_1040_),
    .A(\counter[6] ),
    .B(_1037_));
 sg13g2_nand2_1 _1973_ (.Y(_1041_),
    .A(net570),
    .B(_1040_));
 sg13g2_o21ai_1 _1974_ (.B1(_1041_),
    .Y(_1042_),
    .A1(net570),
    .A2(_1039_));
 sg13g2_o21ai_1 _1975_ (.B1(net571),
    .Y(_1043_),
    .A1(net581),
    .A2(_0942_));
 sg13g2_nor2b_1 _1976_ (.A(_0703_),
    .B_N(_1043_),
    .Y(_1044_));
 sg13g2_o21ai_1 _1977_ (.B1(_1036_),
    .Y(_1045_),
    .A1(_0944_),
    .A2(_1035_));
 sg13g2_xnor2_1 _1978_ (.Y(_1046_),
    .A(net587),
    .B(_1045_));
 sg13g2_xor2_1 _1979_ (.B(_0025_),
    .A(net592),
    .X(_1047_));
 sg13g2_xnor2_1 _1980_ (.Y(_1048_),
    .A(_1035_),
    .B(_1047_));
 sg13g2_xnor2_1 _1981_ (.Y(_1049_),
    .A(net601),
    .B(_0027_));
 sg13g2_a21oi_1 _1982_ (.A1(_1034_),
    .A2(_1049_),
    .Y(_1050_),
    .B1(_1048_));
 sg13g2_and2_1 _1983_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .X(_1051_));
 sg13g2_nor2_1 _1984_ (.A(_1034_),
    .B(_1051_),
    .Y(_1052_));
 sg13g2_xnor2_1 _1985_ (.Y(_1053_),
    .A(net605),
    .B(_1052_));
 sg13g2_nor2_1 _1986_ (.A(_1034_),
    .B(_1049_),
    .Y(_1054_));
 sg13g2_xnor2_1 _1987_ (.Y(_1055_),
    .A(net611),
    .B(\counter[0] ));
 sg13g2_nor2_2 _1988_ (.A(net568),
    .B(_0605_),
    .Y(_1056_));
 sg13g2_nor4_1 _1989_ (.A(_0927_),
    .B(_1054_),
    .C(_1055_),
    .D(_1056_),
    .Y(_1057_));
 sg13g2_nand4_1 _1990_ (.B(_1050_),
    .C(_1053_),
    .A(_1046_),
    .Y(_1058_),
    .D(_1057_));
 sg13g2_a21o_1 _1991_ (.A2(_1040_),
    .A1(_1038_),
    .B1(net578),
    .X(_1059_));
 sg13g2_xnor2_1 _1992_ (.Y(_1060_),
    .A(net530),
    .B(_1036_));
 sg13g2_xnor2_1 _1993_ (.Y(_1061_),
    .A(net584),
    .B(_1060_));
 sg13g2_a21oi_1 _1994_ (.A1(_0688_),
    .A2(_1036_),
    .Y(_1062_),
    .B1(_0683_));
 sg13g2_nor2_1 _1995_ (.A(_0028_),
    .B(_1062_),
    .Y(_1063_));
 sg13g2_a21oi_1 _1996_ (.A1(net567),
    .A2(_1062_),
    .Y(_1064_),
    .B1(_1063_));
 sg13g2_nand3_1 _1997_ (.B(_1061_),
    .C(_1064_),
    .A(_1059_),
    .Y(_1065_));
 sg13g2_nor4_1 _1998_ (.A(_1042_),
    .B(_1044_),
    .C(_1058_),
    .D(_1065_),
    .Y(_1066_));
 sg13g2_or3_2 _1999_ (.A(_0935_),
    .B(_1033_),
    .C(_1066_),
    .X(_1067_));
 sg13g2_inv_1 _2000_ (.Y(_1068_),
    .A(_1067_));
 sg13g2_or2_2 _2001_ (.X(_1069_),
    .B(_0929_),
    .A(_0700_));
 sg13g2_xnor2_1 _2002_ (.Y(_1070_),
    .A(_0491_),
    .B(_1069_));
 sg13g2_xnor2_1 _2003_ (.Y(_1071_),
    .A(net567),
    .B(_1069_));
 sg13g2_nand2_1 _2004_ (.Y(_1072_),
    .A(net566),
    .B(_1069_));
 sg13g2_and2_1 _2005_ (.A(_0605_),
    .B(_1072_),
    .X(_1073_));
 sg13g2_nor2_1 _2006_ (.A(_0605_),
    .B(_1072_),
    .Y(_1074_));
 sg13g2_xnor2_1 _2007_ (.Y(_1075_),
    .A(net570),
    .B(_0975_));
 sg13g2_nor4_2 _2008_ (.A(_1070_),
    .B(_1073_),
    .C(_1074_),
    .Y(_1076_),
    .D(_1075_));
 sg13g2_nand2_1 _2009_ (.Y(_1077_),
    .A(_0985_),
    .B(_1076_));
 sg13g2_xor2_1 _2010_ (.B(net641),
    .A(net633),
    .X(_1078_));
 sg13g2_nand2_1 _2011_ (.Y(_1079_),
    .A(net616),
    .B(_0771_));
 sg13g2_nor3_2 _2012_ (.A(_0726_),
    .B(_1078_),
    .C(_1079_),
    .Y(_1080_));
 sg13g2_and2_2 _2013_ (.A(net667),
    .B(net656),
    .X(_1081_));
 sg13g2_nand2_2 _2014_ (.Y(_1082_),
    .A(net666),
    .B(net657));
 sg13g2_nor2_1 _2015_ (.A(net674),
    .B(net683),
    .Y(_1083_));
 sg13g2_o21ai_1 _2016_ (.B1(net654),
    .Y(_1084_),
    .A1(net664),
    .A2(net675));
 sg13g2_a21oi_1 _2017_ (.A1(net550),
    .A2(_1083_),
    .Y(_1085_),
    .B1(net543));
 sg13g2_nor2_2 _2018_ (.A(net646),
    .B(_1085_),
    .Y(_1086_));
 sg13g2_nand2_1 _2019_ (.Y(_1087_),
    .A(net638),
    .B(_1086_));
 sg13g2_nand2_1 _2020_ (.Y(_1088_),
    .A(_0985_),
    .B(_1087_));
 sg13g2_nor2_2 _2021_ (.A(_0928_),
    .B(_0970_),
    .Y(_1089_));
 sg13g2_nand2_2 _2022_ (.Y(_1090_),
    .A(net536),
    .B(_0971_));
 sg13g2_o21ai_1 _2023_ (.B1(net676),
    .Y(_1091_),
    .A1(net688),
    .A2(net683));
 sg13g2_nand2_1 _2024_ (.Y(_1092_),
    .A(_0821_),
    .B(_1091_));
 sg13g2_and2_2 _2025_ (.A(net661),
    .B(net672),
    .X(_1093_));
 sg13g2_nand2b_1 _2026_ (.Y(_1094_),
    .B(net650),
    .A_N(_1093_));
 sg13g2_a22oi_1 _2027_ (.Y(_1095_),
    .B1(_1094_),
    .B2(net646),
    .A2(_1092_),
    .A1(_1086_));
 sg13g2_nand2_2 _2028_ (.Y(_1096_),
    .A(net638),
    .B(_1095_));
 sg13g2_xnor2_1 _2029_ (.Y(_1097_),
    .A(_1090_),
    .B(_1096_));
 sg13g2_and2_1 _2030_ (.A(net685),
    .B(net679),
    .X(_1098_));
 sg13g2_nand2_1 _2031_ (.Y(_1099_),
    .A(net686),
    .B(net680));
 sg13g2_nor2_2 _2032_ (.A(_0656_),
    .B(net534),
    .Y(_1100_));
 sg13g2_nand2_2 _2033_ (.Y(_1101_),
    .A(net671),
    .B(_1099_));
 sg13g2_nand2_1 _2034_ (.Y(_1102_),
    .A(net545),
    .B(net659));
 sg13g2_nand4_1 _2035_ (.B(net659),
    .C(_0708_),
    .A(net643),
    .Y(_1103_),
    .D(_1100_));
 sg13g2_o21ai_1 _2036_ (.B1(net660),
    .Y(_1104_),
    .A1(net672),
    .A2(net680));
 sg13g2_inv_1 _2037_ (.Y(_1105_),
    .A(_1104_));
 sg13g2_nor2_1 _2038_ (.A(net652),
    .B(_1105_),
    .Y(_1106_));
 sg13g2_nand2b_1 _2039_ (.Y(_1107_),
    .B(_0021_),
    .A_N(net674));
 sg13g2_nand3_1 _2040_ (.B(_1091_),
    .C(_1107_),
    .A(net550),
    .Y(_1108_));
 sg13g2_nand2_1 _2041_ (.Y(_1109_),
    .A(_0819_),
    .B(_1093_));
 sg13g2_a221oi_1 _2042_ (.B2(_1085_),
    .C1(net644),
    .B1(_1109_),
    .A1(_1106_),
    .Y(_1110_),
    .A2(_1108_));
 sg13g2_nor2_1 _2043_ (.A(net652),
    .B(_1093_),
    .Y(_1111_));
 sg13g2_o21ai_1 _2044_ (.B1(net637),
    .Y(_1112_),
    .A1(_0829_),
    .A2(_1093_));
 sg13g2_nor2_1 _2045_ (.A(_0577_),
    .B(_0821_),
    .Y(_1113_));
 sg13g2_o21ai_1 _2046_ (.B1(_1103_),
    .Y(_1114_),
    .A1(_1110_),
    .A2(_1112_));
 sg13g2_xnor2_1 _2047_ (.Y(_1115_),
    .A(_0480_),
    .B(_1114_));
 sg13g2_nor2_1 _2048_ (.A(_1097_),
    .B(_1115_),
    .Y(_1116_));
 sg13g2_nand2_1 _2049_ (.Y(_1117_),
    .A(_0036_),
    .B(_1082_));
 sg13g2_nor2_1 _2050_ (.A(net637),
    .B(_1117_),
    .Y(_1118_));
 sg13g2_a22oi_1 _2051_ (.Y(_1119_),
    .B1(_0821_),
    .B2(_1100_),
    .A2(net654),
    .A1(net675));
 sg13g2_nor2b_1 _2052_ (.A(_1104_),
    .B_N(_1091_),
    .Y(_1120_));
 sg13g2_nand2_1 _2053_ (.Y(_1121_),
    .A(net548),
    .B(\hx0[0] ));
 sg13g2_xor2_1 _2054_ (.B(net682),
    .A(net689),
    .X(_1122_));
 sg13g2_xnor2_1 _2055_ (.Y(_1123_),
    .A(net685),
    .B(net679));
 sg13g2_nand2_1 _2056_ (.Y(_1124_),
    .A(net673),
    .B(_1122_));
 sg13g2_a21oi_1 _2057_ (.A1(_1121_),
    .A2(_1124_),
    .Y(_1125_),
    .B1(net663));
 sg13g2_o21ai_1 _2058_ (.B1(net538),
    .Y(_1126_),
    .A1(_1120_),
    .A2(_1125_));
 sg13g2_nand2b_2 _2059_ (.Y(_1127_),
    .B(net661),
    .A_N(net671));
 sg13g2_nor2_1 _2060_ (.A(net540),
    .B(_1127_),
    .Y(_1128_));
 sg13g2_nand2_1 _2061_ (.Y(_1129_),
    .A(net674),
    .B(net683));
 sg13g2_and3_2 _2062_ (.X(_1130_),
    .A(net689),
    .B(net677),
    .C(net682));
 sg13g2_nor2_2 _2063_ (.A(net666),
    .B(_1130_),
    .Y(_1131_));
 sg13g2_inv_1 _2064_ (.Y(_1132_),
    .A(_1131_));
 sg13g2_nor2b_1 _2065_ (.A(net672),
    .B_N(net681),
    .Y(_1133_));
 sg13g2_nor3_1 _2066_ (.A(net665),
    .B(_1083_),
    .C(_1130_),
    .Y(_1134_));
 sg13g2_o21ai_1 _2067_ (.B1(_0830_),
    .Y(_1135_),
    .A1(_1128_),
    .A2(_1134_));
 sg13g2_nand3_1 _2068_ (.B(net527),
    .C(_1129_),
    .A(net659),
    .Y(_1136_));
 sg13g2_nor2b_2 _2069_ (.A(net673),
    .B_N(net663),
    .Y(_1137_));
 sg13g2_nor2b_2 _2070_ (.A(net662),
    .B_N(net674),
    .Y(_1138_));
 sg13g2_nand2_1 _2071_ (.Y(_1139_),
    .A(net549),
    .B(net676));
 sg13g2_nor2_2 _2072_ (.A(_1137_),
    .B(_1138_),
    .Y(_1140_));
 sg13g2_nand2_1 _2073_ (.Y(_1141_),
    .A(_0828_),
    .B(_1140_));
 sg13g2_nand4_1 _2074_ (.B(_1135_),
    .C(_1136_),
    .A(_1126_),
    .Y(_1142_),
    .D(_1141_));
 sg13g2_a22oi_1 _2075_ (.Y(_1143_),
    .B1(_1142_),
    .B2(net638),
    .A2(_1119_),
    .A1(_1118_));
 sg13g2_nand2b_1 _2076_ (.Y(_1144_),
    .B(_1143_),
    .A_N(net594));
 sg13g2_nor2_1 _2077_ (.A(net541),
    .B(_1143_),
    .Y(_1145_));
 sg13g2_xnor2_1 _2078_ (.Y(_1146_),
    .A(net592),
    .B(_1143_));
 sg13g2_nor2b_2 _2079_ (.A(net686),
    .B_N(net672),
    .Y(_1147_));
 sg13g2_nand2b_2 _2080_ (.Y(_1148_),
    .B(net676),
    .A_N(net688));
 sg13g2_a21o_1 _2081_ (.A2(net683),
    .A1(net688),
    .B1(net673),
    .X(_1149_));
 sg13g2_o21ai_1 _2082_ (.B1(_1148_),
    .Y(_1150_),
    .A1(net674),
    .A2(_1123_));
 sg13g2_a21oi_1 _2083_ (.A1(net672),
    .A2(_1122_),
    .Y(_1151_),
    .B1(_1133_));
 sg13g2_nand2_1 _2084_ (.Y(_1152_),
    .A(net663),
    .B(_1151_));
 sg13g2_a21oi_1 _2085_ (.A1(net549),
    .A2(_1150_),
    .Y(_1153_),
    .B1(_0826_));
 sg13g2_a21oi_1 _2086_ (.A1(net673),
    .A2(net683),
    .Y(_1154_),
    .B1(net662));
 sg13g2_a21o_1 _2087_ (.A2(net683),
    .A1(net676),
    .B1(net664),
    .X(_1155_));
 sg13g2_nand2_1 _2088_ (.Y(_1156_),
    .A(_1127_),
    .B(_1155_));
 sg13g2_nand3_1 _2089_ (.B(_0824_),
    .C(_1156_),
    .A(net653),
    .Y(_1157_));
 sg13g2_nor2_1 _2090_ (.A(_0577_),
    .B(_0737_),
    .Y(_1158_));
 sg13g2_nand3b_1 _2091_ (.B(net652),
    .C(net665),
    .Y(_1159_),
    .A_N(net644));
 sg13g2_a21oi_1 _2092_ (.A1(_1091_),
    .A2(_1107_),
    .Y(_1160_),
    .B1(_1159_));
 sg13g2_nor2_1 _2093_ (.A(_0546_),
    .B(_0831_),
    .Y(_1161_));
 sg13g2_nand2b_2 _2094_ (.Y(_1162_),
    .B(net686),
    .A_N(net660));
 sg13g2_nor2_1 _2095_ (.A(net664),
    .B(net675),
    .Y(_1163_));
 sg13g2_nor4_1 _2096_ (.A(net660),
    .B(_0546_),
    .C(_0831_),
    .D(_1147_),
    .Y(_1164_));
 sg13g2_or2_1 _2097_ (.X(_1165_),
    .B(_1164_),
    .A(_1160_));
 sg13g2_a221oi_1 _2098_ (.B2(_1158_),
    .C1(_1165_),
    .B1(_1157_),
    .A1(_1152_),
    .Y(_1166_),
    .A2(_1153_));
 sg13g2_nor2_1 _2099_ (.A(net545),
    .B(_1166_),
    .Y(_1167_));
 sg13g2_nand2_1 _2100_ (.Y(_1168_),
    .A(net644),
    .B(net650));
 sg13g2_nor4_1 _2101_ (.A(net675),
    .B(_0819_),
    .C(_1102_),
    .D(_1168_),
    .Y(_1169_));
 sg13g2_o21ai_1 _2102_ (.B1(_1106_),
    .Y(_1170_),
    .A1(net664),
    .A2(_1101_));
 sg13g2_a21oi_1 _2103_ (.A1(_1084_),
    .A2(_1170_),
    .Y(_1171_),
    .B1(_0710_));
 sg13g2_nor3_2 _2104_ (.A(_1167_),
    .B(_1169_),
    .C(_1171_),
    .Y(_1172_));
 sg13g2_nor2b_2 _2105_ (.A(net680),
    .B_N(net686),
    .Y(_1173_));
 sg13g2_nand2b_2 _2106_ (.Y(_1174_),
    .B(net685),
    .A_N(net679));
 sg13g2_nor2b_2 _2107_ (.A(net685),
    .B_N(net679),
    .Y(_1175_));
 sg13g2_nand2b_2 _2108_ (.Y(_1176_),
    .B(net681),
    .A_N(net687));
 sg13g2_nand3_1 _2109_ (.B(_1174_),
    .C(_1176_),
    .A(net675),
    .Y(_1177_));
 sg13g2_nor2_1 _2110_ (.A(net660),
    .B(_0831_),
    .Y(_1178_));
 sg13g2_nand2_1 _2111_ (.Y(_1179_),
    .A(net549),
    .B(_0830_));
 sg13g2_a21oi_1 _2112_ (.A1(_1121_),
    .A2(_1177_),
    .Y(_1180_),
    .B1(_1179_));
 sg13g2_o21ai_1 _2113_ (.B1(_0828_),
    .Y(_1181_),
    .A1(_0021_),
    .A2(_1138_));
 sg13g2_a21oi_1 _2114_ (.A1(_0819_),
    .A2(_1138_),
    .Y(_1182_),
    .B1(_1181_));
 sg13g2_mux2_1 _2115_ (.A0(_1174_),
    .A1(_1176_),
    .S(net548),
    .X(_1183_));
 sg13g2_nor2_1 _2116_ (.A(_1159_),
    .B(_1183_),
    .Y(_1184_));
 sg13g2_nand2b_1 _2117_ (.Y(_1185_),
    .B(net688),
    .A_N(net676));
 sg13g2_nand2_1 _2118_ (.Y(_1186_),
    .A(net662),
    .B(_1148_));
 sg13g2_nand3_1 _2119_ (.B(_1148_),
    .C(_1185_),
    .A(net662),
    .Y(_1187_));
 sg13g2_o21ai_1 _2120_ (.B1(net549),
    .Y(_1188_),
    .A1(_0820_),
    .A2(_1130_));
 sg13g2_a21oi_1 _2121_ (.A1(_1187_),
    .A2(_1188_),
    .Y(_1189_),
    .B1(_0826_));
 sg13g2_nand2b_1 _2122_ (.Y(_1190_),
    .B(net687),
    .A_N(net670));
 sg13g2_nand3b_1 _2123_ (.B(net679),
    .C(net685),
    .Y(_1191_),
    .A_N(net669));
 sg13g2_o21ai_1 _2124_ (.B1(net669),
    .Y(_1192_),
    .A1(net685),
    .A2(net679));
 sg13g2_and3_1 _2125_ (.X(_1193_),
    .A(net663),
    .B(_1191_),
    .C(_1192_));
 sg13g2_nand2_1 _2126_ (.Y(_1194_),
    .A(_1129_),
    .B(_1149_));
 sg13g2_a221oi_1 _2127_ (.B2(_1149_),
    .C1(net662),
    .B1(_1129_),
    .A1(net548),
    .Y(_1195_),
    .A2(net540));
 sg13g2_o21ai_1 _2128_ (.B1(net527),
    .Y(_1196_),
    .A1(_1193_),
    .A2(_1195_));
 sg13g2_nor4_1 _2129_ (.A(_1180_),
    .B(_1182_),
    .C(_1184_),
    .D(_1189_),
    .Y(_1197_));
 sg13g2_and2_1 _2130_ (.A(net636),
    .B(_1196_),
    .X(_1198_));
 sg13g2_nand3b_1 _2131_ (.B(net681),
    .C(net687),
    .Y(_1199_),
    .A_N(net672));
 sg13g2_nand2_1 _2132_ (.Y(_1200_),
    .A(net673),
    .B(_0021_));
 sg13g2_a21o_1 _2133_ (.A2(_1200_),
    .A1(_1199_),
    .B1(net663),
    .X(_1201_));
 sg13g2_nand4_1 _2134_ (.B(net666),
    .C(net677),
    .A(net688),
    .Y(_1202_),
    .D(net682));
 sg13g2_o21ai_1 _2135_ (.B1(_1201_),
    .Y(_1203_),
    .A1(_1104_),
    .A2(_1130_));
 sg13g2_nand2b_1 _2136_ (.Y(_1204_),
    .B(_0830_),
    .A_N(_1163_));
 sg13g2_nand2_1 _2137_ (.Y(_1205_),
    .A(net670),
    .B(net540));
 sg13g2_nor2_1 _2138_ (.A(net661),
    .B(_1205_),
    .Y(_1206_));
 sg13g2_nand3_1 _2139_ (.B(net670),
    .C(net540),
    .A(net551),
    .Y(_1207_));
 sg13g2_nand2b_1 _2140_ (.Y(_1208_),
    .B(_1207_),
    .A_N(_1168_));
 sg13g2_a21o_1 _2141_ (.A2(_1208_),
    .A1(_1204_),
    .B1(_1105_),
    .X(_1209_));
 sg13g2_a21oi_1 _2142_ (.A1(net538),
    .A2(_1203_),
    .Y(_1210_),
    .B1(net636));
 sg13g2_a22oi_1 _2143_ (.Y(_1211_),
    .B1(_1209_),
    .B2(_1210_),
    .A2(_1198_),
    .A1(_1197_));
 sg13g2_nor2_1 _2144_ (.A(net607),
    .B(_1211_),
    .Y(_1212_));
 sg13g2_or2_1 _2145_ (.X(_1213_),
    .B(_1211_),
    .A(net605));
 sg13g2_nand2_1 _2146_ (.Y(_1214_),
    .A(net605),
    .B(_1211_));
 sg13g2_xnor2_1 _2147_ (.Y(_1215_),
    .A(net605),
    .B(_1211_));
 sg13g2_o21ai_1 _2148_ (.B1(_1200_),
    .Y(_1216_),
    .A1(net673),
    .A2(net540));
 sg13g2_and3_1 _2149_ (.X(_1217_),
    .A(net551),
    .B(_1199_),
    .C(_1216_));
 sg13g2_a22oi_1 _2150_ (.Y(_1218_),
    .B1(_1137_),
    .B2(_0021_),
    .A2(_1122_),
    .A1(_1093_));
 sg13g2_inv_1 _2151_ (.Y(_1219_),
    .A(_1218_));
 sg13g2_o21ai_1 _2152_ (.B1(net538),
    .Y(_1220_),
    .A1(_1217_),
    .A2(_1219_));
 sg13g2_or2_1 _2153_ (.X(_1221_),
    .B(net669),
    .A(net685));
 sg13g2_o21ai_1 _2154_ (.B1(_1192_),
    .Y(_1222_),
    .A1(net679),
    .A2(_1221_));
 sg13g2_nand2_2 _2155_ (.Y(_1223_),
    .A(net551),
    .B(_1222_));
 sg13g2_nand3_1 _2156_ (.B(_1106_),
    .C(_1223_),
    .A(net644),
    .Y(_1224_));
 sg13g2_nor2_1 _2157_ (.A(net637),
    .B(_1160_),
    .Y(_1225_));
 sg13g2_nand3_1 _2158_ (.B(net658),
    .C(net540),
    .A(net671),
    .Y(_1226_));
 sg13g2_o21ai_1 _2159_ (.B1(_1099_),
    .Y(_1227_),
    .A1(net672),
    .A2(net540));
 sg13g2_a21oi_1 _2160_ (.A1(net548),
    .A2(_0819_),
    .Y(_1228_),
    .B1(net534));
 sg13g2_a22oi_1 _2161_ (.Y(_1229_),
    .B1(_1227_),
    .B2(_1178_),
    .A2(_1226_),
    .A1(net527));
 sg13g2_and4_1 _2162_ (.A(_1220_),
    .B(_1224_),
    .C(_1225_),
    .D(_1229_),
    .X(_1230_));
 sg13g2_nand3_1 _2163_ (.B(_1148_),
    .C(_1185_),
    .A(net549),
    .Y(_1231_));
 sg13g2_mux2_1 _2164_ (.A0(_1122_),
    .A1(_1174_),
    .S(net548),
    .X(_1232_));
 sg13g2_nand2_1 _2165_ (.Y(_1233_),
    .A(net662),
    .B(_1232_));
 sg13g2_a21oi_1 _2166_ (.A1(_1231_),
    .A2(_1233_),
    .Y(_1234_),
    .B1(_0713_));
 sg13g2_mux2_1 _2167_ (.A0(_1123_),
    .A1(_1175_),
    .S(net672),
    .X(_1235_));
 sg13g2_nor2_1 _2168_ (.A(net683),
    .B(_1139_),
    .Y(_1236_));
 sg13g2_o21ai_1 _2169_ (.B1(_0830_),
    .Y(_1237_),
    .A1(net683),
    .A2(_1139_));
 sg13g2_o21ai_1 _2170_ (.B1(_0403_),
    .Y(_1238_),
    .A1(net548),
    .A2(net681));
 sg13g2_a21oi_1 _2171_ (.A1(net663),
    .A2(_1192_),
    .Y(_1239_),
    .B1(_0826_));
 sg13g2_o21ai_1 _2172_ (.B1(_1239_),
    .Y(_1240_),
    .A1(net662),
    .A2(_1238_));
 sg13g2_a22oi_1 _2173_ (.Y(_1241_),
    .B1(_1237_),
    .B2(_1240_),
    .A2(_1235_),
    .A1(_1081_));
 sg13g2_o21ai_1 _2174_ (.B1(_0828_),
    .Y(_1242_),
    .A1(net688),
    .A2(_1138_));
 sg13g2_o21ai_1 _2175_ (.B1(net636),
    .Y(_1243_),
    .A1(_1236_),
    .A2(_1242_));
 sg13g2_nor3_2 _2176_ (.A(_1234_),
    .B(_1241_),
    .C(_1243_),
    .Y(_1244_));
 sg13g2_nor2_1 _2177_ (.A(_1230_),
    .B(_1244_),
    .Y(_1245_));
 sg13g2_o21ai_1 _2178_ (.B1(_0392_),
    .Y(_1246_),
    .A1(_1230_),
    .A2(_1244_));
 sg13g2_a21o_1 _2179_ (.A2(_1246_),
    .A1(_1215_),
    .B1(_1212_),
    .X(_1247_));
 sg13g2_xnor2_1 _2180_ (.Y(_1248_),
    .A(net603),
    .B(_1172_));
 sg13g2_a22oi_1 _2181_ (.Y(_1249_),
    .B1(_1247_),
    .B2(_1248_),
    .A2(_1172_),
    .A1(net600));
 sg13g2_o21ai_1 _2182_ (.B1(_1144_),
    .Y(_1250_),
    .A1(_1146_),
    .A2(_1249_));
 sg13g2_o21ai_1 _2183_ (.B1(net588),
    .Y(_1251_),
    .A1(net585),
    .A2(_1096_));
 sg13g2_nor2_1 _2184_ (.A(_1114_),
    .B(_1251_),
    .Y(_1252_));
 sg13g2_a221oi_1 _2185_ (.B2(_1250_),
    .C1(_1252_),
    .B1(_1116_),
    .A1(_1090_),
    .Y(_1253_),
    .A2(_1096_));
 sg13g2_nand3_1 _2186_ (.B(_0984_),
    .C(_1086_),
    .A(net638),
    .Y(_1254_));
 sg13g2_xnor2_1 _2187_ (.Y(_1255_),
    .A(net612),
    .B(_1245_));
 sg13g2_nand4_1 _2188_ (.B(_1215_),
    .C(_1248_),
    .A(_1116_),
    .Y(_1256_),
    .D(_1255_));
 sg13g2_o21ai_1 _2189_ (.B1(_1254_),
    .Y(_1257_),
    .A1(_1146_),
    .A2(_1256_));
 sg13g2_o21ai_1 _2190_ (.B1(_1088_),
    .Y(_1258_),
    .A1(_1253_),
    .A2(_1257_));
 sg13g2_nand3b_1 _2191_ (.B(net681),
    .C(net675),
    .Y(_1259_),
    .A_N(net659));
 sg13g2_a21oi_1 _2192_ (.A1(net650),
    .A2(_1259_),
    .Y(_1260_),
    .B1(_0629_));
 sg13g2_nand2_2 _2193_ (.Y(_1261_),
    .A(_0639_),
    .B(_1260_));
 sg13g2_inv_1 _2194_ (.Y(_1262_),
    .A(_1261_));
 sg13g2_nand2_1 _2195_ (.Y(_1263_),
    .A(_0985_),
    .B(_1261_));
 sg13g2_nand3_1 _2196_ (.B(_1155_),
    .C(_1194_),
    .A(net652),
    .Y(_1264_));
 sg13g2_and2_1 _2197_ (.A(net543),
    .B(_1259_),
    .X(_1265_));
 sg13g2_o21ai_1 _2198_ (.B1(_1265_),
    .Y(_1266_),
    .A1(net664),
    .A2(_1101_));
 sg13g2_nand3_1 _2199_ (.B(_1264_),
    .C(_1266_),
    .A(net644),
    .Y(_1267_));
 sg13g2_nor3_1 _2200_ (.A(net646),
    .B(net650),
    .C(_1163_),
    .Y(_1268_));
 sg13g2_nor2_1 _2201_ (.A(net636),
    .B(_1268_),
    .Y(_1269_));
 sg13g2_nor2_1 _2202_ (.A(net650),
    .B(_0803_),
    .Y(_1270_));
 sg13g2_a22oi_1 _2203_ (.Y(_1271_),
    .B1(_1270_),
    .B2(_1128_),
    .A2(_1269_),
    .A1(_1267_));
 sg13g2_nor3_1 _2204_ (.A(net543),
    .B(net659),
    .C(_1100_),
    .Y(_1272_));
 sg13g2_o21ai_1 _2205_ (.B1(net646),
    .Y(_1273_),
    .A1(_1265_),
    .A2(_1272_));
 sg13g2_a21oi_2 _2206_ (.B1(_0629_),
    .Y(_1274_),
    .A2(_1273_),
    .A1(_1204_));
 sg13g2_nor2_1 _2207_ (.A(_1090_),
    .B(_1274_),
    .Y(_1275_));
 sg13g2_xnor2_1 _2208_ (.Y(_1276_),
    .A(_1089_),
    .B(_1274_));
 sg13g2_xnor2_1 _2209_ (.Y(_1277_),
    .A(net588),
    .B(_1271_));
 sg13g2_nor2_1 _2210_ (.A(_1276_),
    .B(_1277_),
    .Y(_1278_));
 sg13g2_nor2_1 _2211_ (.A(_1082_),
    .B(_1091_),
    .Y(_1279_));
 sg13g2_nor4_1 _2212_ (.A(net545),
    .B(net643),
    .C(_1111_),
    .D(_1279_),
    .Y(_1280_));
 sg13g2_mux2_1 _2213_ (.A0(_1100_),
    .A1(_1216_),
    .S(net663),
    .X(_1281_));
 sg13g2_nor2_1 _2214_ (.A(net673),
    .B(_1122_),
    .Y(_1282_));
 sg13g2_o21ai_1 _2215_ (.B1(_1201_),
    .Y(_1283_),
    .A1(_1186_),
    .A2(_1282_));
 sg13g2_mux4_1 _2216_ (.S0(net652),
    .A0(_1105_),
    .A1(_1140_),
    .A2(_1281_),
    .A3(_1283_),
    .S1(net644),
    .X(_1284_));
 sg13g2_a21oi_2 _2217_ (.B1(_1280_),
    .Y(_1285_),
    .A2(_1284_),
    .A1(net545));
 sg13g2_nor2b_1 _2218_ (.A(net594),
    .B_N(_1285_),
    .Y(_1286_));
 sg13g2_and2_1 _2219_ (.A(net541),
    .B(_1285_),
    .X(_1287_));
 sg13g2_nand2b_1 _2220_ (.Y(_1288_),
    .B(net592),
    .A_N(_1285_));
 sg13g2_nor2b_1 _2221_ (.A(_1287_),
    .B_N(_1288_),
    .Y(_1289_));
 sg13g2_inv_1 _2222_ (.Y(_1290_),
    .A(_1289_));
 sg13g2_a21oi_1 _2223_ (.A1(_1121_),
    .A2(_1177_),
    .Y(_1291_),
    .B1(net551));
 sg13g2_o21ai_1 _2224_ (.B1(net527),
    .Y(_1292_),
    .A1(_1217_),
    .A2(_1291_));
 sg13g2_a221oi_1 _2225_ (.B2(_0021_),
    .C1(_1138_),
    .B1(_1137_),
    .A1(net673),
    .Y(_1293_),
    .A2(net535));
 sg13g2_inv_1 _2226_ (.Y(_1294_),
    .A(_1293_));
 sg13g2_nor2_2 _2227_ (.A(net549),
    .B(_0820_),
    .Y(_1295_));
 sg13g2_nand2b_2 _2228_ (.Y(_1296_),
    .B(net668),
    .A_N(_0820_));
 sg13g2_a221oi_1 _2229_ (.B2(_1295_),
    .C1(_0829_),
    .B1(_1200_),
    .A1(_1149_),
    .Y(_1297_),
    .A2(_1154_));
 sg13g2_a221oi_1 _2230_ (.B2(net538),
    .C1(_1297_),
    .B1(_1294_),
    .A1(_0040_),
    .Y(_1298_),
    .A2(_0830_));
 sg13g2_a21oi_1 _2231_ (.A1(_1292_),
    .A2(_1298_),
    .Y(_1299_),
    .B1(net636));
 sg13g2_a21oi_1 _2232_ (.A1(net652),
    .A2(_1155_),
    .Y(_1300_),
    .B1(_1111_));
 sg13g2_nor3_1 _2233_ (.A(_0803_),
    .B(_1279_),
    .C(_1300_),
    .Y(_1301_));
 sg13g2_nor3_1 _2234_ (.A(net545),
    .B(_1159_),
    .C(_1191_),
    .Y(_1302_));
 sg13g2_nor2_1 _2235_ (.A(net551),
    .B(_1191_),
    .Y(_1303_));
 sg13g2_nor3_2 _2236_ (.A(_1299_),
    .B(_1301_),
    .C(_1302_),
    .Y(_1304_));
 sg13g2_nand2_1 _2237_ (.Y(_1305_),
    .A(net600),
    .B(_1304_));
 sg13g2_xnor2_1 _2238_ (.Y(_1306_),
    .A(net554),
    .B(_1304_));
 sg13g2_o21ai_1 _2239_ (.B1(net666),
    .Y(_1307_),
    .A1(_0820_),
    .A2(_1130_));
 sg13g2_nand2_1 _2240_ (.Y(_1308_),
    .A(_1231_),
    .B(_1307_));
 sg13g2_nand2_1 _2241_ (.Y(_1309_),
    .A(_0403_),
    .B(_1137_));
 sg13g2_o21ai_1 _2242_ (.B1(_1218_),
    .Y(_1310_),
    .A1(net663),
    .A2(_1228_));
 sg13g2_nand2_1 _2243_ (.Y(_1311_),
    .A(net664),
    .B(_1150_));
 sg13g2_a21oi_1 _2244_ (.A1(net551),
    .A2(_1183_),
    .Y(_1312_),
    .B1(_0829_));
 sg13g2_a22oi_1 _2245_ (.Y(_1313_),
    .B1(_1310_),
    .B2(net538),
    .A2(_1308_),
    .A1(net527));
 sg13g2_a221oi_1 _2246_ (.B2(_1312_),
    .C1(net636),
    .B1(_1311_),
    .A1(_1161_),
    .Y(_1314_),
    .A2(_1309_));
 sg13g2_a21oi_1 _2247_ (.A1(net549),
    .A2(_1216_),
    .Y(_1315_),
    .B1(_1120_));
 sg13g2_nand2b_1 _2248_ (.Y(_1316_),
    .B(net527),
    .A_N(_1315_));
 sg13g2_nor2_1 _2249_ (.A(_0831_),
    .B(_1154_),
    .Y(_1317_));
 sg13g2_nand2b_1 _2250_ (.Y(_1318_),
    .B(_1317_),
    .A_N(_1303_));
 sg13g2_nand3_1 _2251_ (.B(_1127_),
    .C(_1155_),
    .A(_0828_),
    .Y(_1319_));
 sg13g2_and3_1 _2252_ (.X(_1320_),
    .A(net636),
    .B(_1318_),
    .C(_1319_));
 sg13g2_a22oi_1 _2253_ (.Y(_1321_),
    .B1(_1316_),
    .B2(_1320_),
    .A2(_1314_),
    .A1(_1313_));
 sg13g2_nor2_1 _2254_ (.A(net607),
    .B(_1321_),
    .Y(_1322_));
 sg13g2_o21ai_1 _2255_ (.B1(net527),
    .Y(_1323_),
    .A1(_1151_),
    .A2(_1162_));
 sg13g2_a21o_1 _2256_ (.A2(_1162_),
    .A1(_1151_),
    .B1(_1323_),
    .X(_1324_));
 sg13g2_a21oi_1 _2257_ (.A1(net661),
    .A2(_1227_),
    .Y(_1325_),
    .B1(_0829_));
 sg13g2_xnor2_1 _2258_ (.Y(_1326_),
    .A(net669),
    .B(net534));
 sg13g2_nand2_1 _2259_ (.Y(_1327_),
    .A(_1101_),
    .B(_1191_));
 sg13g2_nand2_1 _2260_ (.Y(_1328_),
    .A(net660),
    .B(_1326_));
 sg13g2_o21ai_1 _2261_ (.B1(net636),
    .Y(_1329_),
    .A1(_0826_),
    .A2(_1303_));
 sg13g2_a221oi_1 _2262_ (.B2(_1317_),
    .C1(_1329_),
    .B1(_1328_),
    .A1(_1201_),
    .Y(_1330_),
    .A2(_1325_));
 sg13g2_o21ai_1 _2263_ (.B1(_1187_),
    .Y(_1331_),
    .A1(net662),
    .A2(_1235_));
 sg13g2_a21oi_1 _2264_ (.A1(net660),
    .A2(_1133_),
    .Y(_1332_),
    .B1(_0829_));
 sg13g2_o21ai_1 _2265_ (.B1(_1332_),
    .Y(_1333_),
    .A1(net660),
    .A2(_1232_));
 sg13g2_o21ai_1 _2266_ (.B1(_1162_),
    .Y(_1334_),
    .A1(_1104_),
    .A2(_1147_));
 sg13g2_o21ai_1 _2267_ (.B1(net545),
    .Y(_1335_),
    .A1(_0831_),
    .A2(_1334_));
 sg13g2_nand2_1 _2268_ (.Y(_1336_),
    .A(\hx0[0] ),
    .B(_1093_));
 sg13g2_mux2_1 _2269_ (.A0(net534),
    .A1(_1173_),
    .S(net548),
    .X(_1337_));
 sg13g2_o21ai_1 _2270_ (.B1(_1336_),
    .Y(_1338_),
    .A1(_1140_),
    .A2(_1337_));
 sg13g2_a221oi_1 _2271_ (.B2(net527),
    .C1(_1335_),
    .B1(_1338_),
    .A1(net538),
    .Y(_1339_),
    .A2(_1331_));
 sg13g2_a22oi_1 _2272_ (.Y(_1340_),
    .B1(_1333_),
    .B2(_1339_),
    .A2(_1330_),
    .A1(_1324_));
 sg13g2_nand2b_1 _2273_ (.Y(_1341_),
    .B(net612),
    .A_N(_1340_));
 sg13g2_nand2_1 _2274_ (.Y(_1342_),
    .A(net607),
    .B(_1321_));
 sg13g2_a21oi_1 _2275_ (.A1(_1341_),
    .A2(_1342_),
    .Y(_1343_),
    .B1(_1322_));
 sg13g2_o21ai_1 _2276_ (.B1(_1305_),
    .Y(_1344_),
    .A1(_1306_),
    .A2(_1343_));
 sg13g2_a21o_1 _2277_ (.A2(_1344_),
    .A1(_1290_),
    .B1(_1286_),
    .X(_1345_));
 sg13g2_nand3b_1 _2278_ (.B(_1271_),
    .C(net588),
    .Y(_1346_),
    .A_N(_1276_));
 sg13g2_o21ai_1 _2279_ (.B1(_1346_),
    .Y(_1347_),
    .A1(_1089_),
    .A2(_1274_));
 sg13g2_a21oi_1 _2280_ (.A1(_1278_),
    .A2(_1345_),
    .Y(_1348_),
    .B1(_1347_));
 sg13g2_nand2b_1 _2281_ (.Y(_1349_),
    .B(net610),
    .A_N(_1340_));
 sg13g2_xnor2_1 _2282_ (.Y(_1350_),
    .A(_0392_),
    .B(_1340_));
 sg13g2_nand4_1 _2283_ (.B(_1290_),
    .C(_1342_),
    .A(_1278_),
    .Y(_1351_),
    .D(_1350_));
 sg13g2_nor3_1 _2284_ (.A(_1306_),
    .B(_1322_),
    .C(_1351_),
    .Y(_1352_));
 sg13g2_o21ai_1 _2285_ (.B1(_1263_),
    .Y(_1353_),
    .A1(_1348_),
    .A2(_1352_));
 sg13g2_nand3_1 _2286_ (.B(net616),
    .C(_1078_),
    .A(\hvsync_gen.hpos[8] ),
    .Y(_1354_));
 sg13g2_a21oi_1 _2287_ (.A1(_0984_),
    .A2(_1262_),
    .Y(_1355_),
    .B1(_1354_));
 sg13g2_a22oi_1 _2288_ (.Y(_1356_),
    .B1(_1353_),
    .B2(_1355_),
    .A2(_1258_),
    .A1(_1080_));
 sg13g2_a21oi_1 _2289_ (.A1(net552),
    .A2(_1274_),
    .Y(_1357_),
    .B1(net588));
 sg13g2_a21oi_1 _2290_ (.A1(_1271_),
    .A2(_1357_),
    .Y(_1358_),
    .B1(_1275_));
 sg13g2_nor2_1 _2291_ (.A(net605),
    .B(_1321_),
    .Y(_1359_));
 sg13g2_nand2_1 _2292_ (.Y(_1360_),
    .A(net605),
    .B(_1321_));
 sg13g2_a21o_1 _2293_ (.A2(_1360_),
    .A1(_1349_),
    .B1(_1359_),
    .X(_1361_));
 sg13g2_a221oi_1 _2294_ (.B2(_1361_),
    .C1(_1287_),
    .B1(_1306_),
    .A1(_0675_),
    .Y(_1362_),
    .A2(_1304_));
 sg13g2_xnor2_1 _2295_ (.Y(_1363_),
    .A(net542),
    .B(_1271_));
 sg13g2_nand3_1 _2296_ (.B(_1288_),
    .C(_1363_),
    .A(_1276_),
    .Y(_1364_));
 sg13g2_o21ai_1 _2297_ (.B1(_1358_),
    .Y(_1365_),
    .A1(_1362_),
    .A2(_1364_));
 sg13g2_nand3_1 _2298_ (.B(_1360_),
    .C(_1363_),
    .A(_1276_),
    .Y(_1366_));
 sg13g2_nor2_1 _2299_ (.A(_1359_),
    .B(_1366_),
    .Y(_1367_));
 sg13g2_xnor2_1 _2300_ (.Y(_1368_),
    .A(net556),
    .B(_1340_));
 sg13g2_nand4_1 _2301_ (.B(_1306_),
    .C(_1367_),
    .A(_1289_),
    .Y(_1369_),
    .D(_1368_));
 sg13g2_a22oi_1 _2302_ (.Y(_1370_),
    .B1(_1365_),
    .B2(_1369_),
    .A2(_1261_),
    .A1(_0984_));
 sg13g2_nor2_1 _2303_ (.A(_0984_),
    .B(_1261_),
    .Y(_1371_));
 sg13g2_nor3_1 _2304_ (.A(_1354_),
    .B(_1370_),
    .C(_1371_),
    .Y(_1372_));
 sg13g2_nand2_1 _2305_ (.Y(_1373_),
    .A(_0984_),
    .B(_1087_));
 sg13g2_a22oi_1 _2306_ (.Y(_1374_),
    .B1(_1172_),
    .B2(_0675_),
    .A2(_1143_),
    .A1(net541));
 sg13g2_o21ai_1 _2307_ (.B1(_1214_),
    .Y(_1375_),
    .A1(_0392_),
    .A2(_1245_));
 sg13g2_a21o_1 _2308_ (.A2(_1375_),
    .A1(_1213_),
    .B1(_1248_),
    .X(_1376_));
 sg13g2_xnor2_1 _2309_ (.Y(_1377_),
    .A(net587),
    .B(_1114_));
 sg13g2_nand2_1 _2310_ (.Y(_1378_),
    .A(_1097_),
    .B(_1377_));
 sg13g2_or2_1 _2311_ (.X(_1379_),
    .B(_1378_),
    .A(_1145_));
 sg13g2_a21oi_1 _2312_ (.A1(_1374_),
    .A2(_1376_),
    .Y(_1380_),
    .B1(_1379_));
 sg13g2_nand2_1 _2313_ (.Y(_1381_),
    .A(_0480_),
    .B(_1097_));
 sg13g2_nand2_1 _2314_ (.Y(_1382_),
    .A(_1089_),
    .B(_1096_));
 sg13g2_o21ai_1 _2315_ (.B1(_1382_),
    .Y(_1383_),
    .A1(_1114_),
    .A2(_1381_));
 sg13g2_nor2_1 _2316_ (.A(_1215_),
    .B(_1378_),
    .Y(_1384_));
 sg13g2_nor2_1 _2317_ (.A(_1248_),
    .B(_1255_),
    .Y(_1385_));
 sg13g2_nand3_1 _2318_ (.B(_1384_),
    .C(_1385_),
    .A(_1146_),
    .Y(_1386_));
 sg13g2_o21ai_1 _2319_ (.B1(_1386_),
    .Y(_1387_),
    .A1(_1380_),
    .A2(_1383_));
 sg13g2_o21ai_1 _2320_ (.B1(_1080_),
    .Y(_1388_),
    .A1(_0984_),
    .A2(_1087_));
 sg13g2_a21oi_1 _2321_ (.A1(_1373_),
    .A2(_1387_),
    .Y(_1389_),
    .B1(_1388_));
 sg13g2_xnor2_1 _2322_ (.Y(_1390_),
    .A(_0502_),
    .B(_1072_));
 sg13g2_nor3_1 _2323_ (.A(_0982_),
    .B(_1071_),
    .C(_1390_),
    .Y(_1391_));
 sg13g2_o21ai_1 _2324_ (.B1(_1391_),
    .Y(_1392_),
    .A1(_1372_),
    .A2(_1389_));
 sg13g2_o21ai_1 _2325_ (.B1(_1392_),
    .Y(_1393_),
    .A1(_1077_),
    .A2(_1356_));
 sg13g2_inv_1 _2326_ (.Y(_1394_),
    .A(_1393_));
 sg13g2_nor2_2 _2327_ (.A(_1067_),
    .B(_1393_),
    .Y(_1395_));
 sg13g2_o21ai_1 _2328_ (.B1(net646),
    .Y(_1396_),
    .A1(net654),
    .A2(_1295_));
 sg13g2_nor2_1 _2329_ (.A(net546),
    .B(_1396_),
    .Y(_1397_));
 sg13g2_xnor2_1 _2330_ (.Y(_1398_),
    .A(net546),
    .B(_1396_));
 sg13g2_xor2_1 _2331_ (.B(_1398_),
    .A(net577),
    .X(_1399_));
 sg13g2_nand3_1 _2332_ (.B(net544),
    .C(_1296_),
    .A(_0577_),
    .Y(_1400_));
 sg13g2_nand2_1 _2333_ (.Y(_1401_),
    .A(_1396_),
    .B(_1400_));
 sg13g2_xnor2_1 _2334_ (.Y(_1402_),
    .A(net543),
    .B(_1295_));
 sg13g2_nand2_1 _2335_ (.Y(_1403_),
    .A(net589),
    .B(_1402_));
 sg13g2_nor2_1 _2336_ (.A(_0425_),
    .B(_1123_),
    .Y(_1404_));
 sg13g2_xnor2_1 _2337_ (.Y(_1405_),
    .A(net555),
    .B(_1122_));
 sg13g2_a21oi_1 _2338_ (.A1(_0851_),
    .A2(_1405_),
    .Y(_1406_),
    .B1(_1404_));
 sg13g2_xnor2_1 _2339_ (.Y(_1407_),
    .A(_0675_),
    .B(_1222_));
 sg13g2_nor2_1 _2340_ (.A(_1406_),
    .B(_1407_),
    .Y(_1408_));
 sg13g2_nand2_1 _2341_ (.Y(_1409_),
    .A(_0824_),
    .B(_1296_));
 sg13g2_a221oi_1 _2342_ (.B2(net598),
    .C1(_1408_),
    .B1(_1409_),
    .A1(net604),
    .Y(_1410_),
    .A2(_1222_));
 sg13g2_or2_1 _2343_ (.X(_1411_),
    .B(_1402_),
    .A(net589));
 sg13g2_o21ai_1 _2344_ (.B1(_1411_),
    .Y(_1412_),
    .A1(net598),
    .A2(_1409_));
 sg13g2_o21ai_1 _2345_ (.B1(_1403_),
    .Y(_1413_),
    .A1(_1410_),
    .A2(_1412_));
 sg13g2_xnor2_1 _2346_ (.Y(_1414_),
    .A(net584),
    .B(_1401_));
 sg13g2_a22oi_1 _2347_ (.Y(_1415_),
    .B1(_1413_),
    .B2(_1414_),
    .A2(_1401_),
    .A1(net586));
 sg13g2_nor2_1 _2348_ (.A(_1399_),
    .B(_1415_),
    .Y(_1416_));
 sg13g2_xor2_1 _2349_ (.B(_1397_),
    .A(net629),
    .X(_1417_));
 sg13g2_a221oi_1 _2350_ (.B2(net572),
    .C1(_1416_),
    .B1(_1417_),
    .A1(net580),
    .Y(_1418_),
    .A2(_1398_));
 sg13g2_nor2_1 _2351_ (.A(net627),
    .B(_1397_),
    .Y(_1419_));
 sg13g2_nor3_2 _2352_ (.A(net547),
    .B(_0771_),
    .C(_1396_),
    .Y(_1420_));
 sg13g2_nor3_1 _2353_ (.A(_0718_),
    .B(_1419_),
    .C(_1420_),
    .Y(_1421_));
 sg13g2_xnor2_1 _2354_ (.Y(_1422_),
    .A(_0622_),
    .B(_1421_));
 sg13g2_o21ai_1 _2355_ (.B1(_1422_),
    .Y(_1423_),
    .A1(net573),
    .A2(_1417_));
 sg13g2_xnor2_1 _2356_ (.Y(_1424_),
    .A(_0597_),
    .B(_1420_));
 sg13g2_nor2_1 _2357_ (.A(_0491_),
    .B(_1421_),
    .Y(_1425_));
 sg13g2_a21oi_1 _2358_ (.A1(net560),
    .A2(_1424_),
    .Y(_1426_),
    .B1(_1425_));
 sg13g2_o21ai_1 _2359_ (.B1(_1426_),
    .Y(_1427_),
    .A1(_1418_),
    .A2(_1423_));
 sg13g2_nor2_1 _2360_ (.A(net560),
    .B(_1424_),
    .Y(_1428_));
 sg13g2_a21oi_1 _2361_ (.A1(net618),
    .A2(_1420_),
    .Y(_1429_),
    .B1(_1428_));
 sg13g2_nor2_2 _2362_ (.A(net597),
    .B(net590),
    .Y(_1430_));
 sg13g2_xor2_1 _2363_ (.B(_1430_),
    .A(net583),
    .X(_1431_));
 sg13g2_and2_1 _2364_ (.A(net598),
    .B(net667),
    .X(_1432_));
 sg13g2_nor2b_1 _2365_ (.A(net608),
    .B_N(net684),
    .Y(_1433_));
 sg13g2_nand2_1 _2366_ (.Y(_1434_),
    .A(_0403_),
    .B(net613));
 sg13g2_nand2b_1 _2367_ (.Y(_1435_),
    .B(net608),
    .A_N(net682));
 sg13g2_a21oi_1 _2368_ (.A1(_1434_),
    .A2(_1435_),
    .Y(_1436_),
    .B1(_1433_));
 sg13g2_nor3_1 _2369_ (.A(net604),
    .B(net548),
    .C(net526),
    .Y(_1437_));
 sg13g2_nand2b_1 _2370_ (.Y(_1438_),
    .B(_0857_),
    .A_N(net526));
 sg13g2_nor2_1 _2371_ (.A(_1436_),
    .B(_1438_),
    .Y(_1439_));
 sg13g2_nor3_2 _2372_ (.A(_1432_),
    .B(_1437_),
    .C(_1439_),
    .Y(_1440_));
 sg13g2_nand2_2 _2373_ (.Y(_1441_),
    .A(net597),
    .B(net589));
 sg13g2_nor2b_2 _2374_ (.A(_1430_),
    .B_N(_1441_),
    .Y(_1442_));
 sg13g2_nand2b_2 _2375_ (.Y(_1443_),
    .B(_1441_),
    .A_N(_1430_));
 sg13g2_nand2_1 _2376_ (.Y(_1444_),
    .A(net657),
    .B(_1442_));
 sg13g2_a22oi_1 _2377_ (.Y(_1445_),
    .B1(_1443_),
    .B2(net544),
    .A2(_1431_),
    .A1(_0639_));
 sg13g2_o21ai_1 _2378_ (.B1(_1445_),
    .Y(_1446_),
    .A1(_0639_),
    .A2(_1431_));
 sg13g2_a21oi_1 _2379_ (.A1(_1440_),
    .A2(_1444_),
    .Y(_1447_),
    .B1(_1446_));
 sg13g2_a21oi_1 _2380_ (.A1(net648),
    .A2(_1431_),
    .Y(_1448_),
    .B1(_1447_));
 sg13g2_nor2_2 _2381_ (.A(net597),
    .B(_0971_),
    .Y(_1449_));
 sg13g2_nand2_2 _2382_ (.Y(_1450_),
    .A(net552),
    .B(_1430_));
 sg13g2_nand2_1 _2383_ (.Y(_1451_),
    .A(net579),
    .B(_1450_));
 sg13g2_xnor2_1 _2384_ (.Y(_1452_),
    .A(net580),
    .B(_1449_));
 sg13g2_xnor2_1 _2385_ (.Y(_1453_),
    .A(net635),
    .B(_1452_));
 sg13g2_nor2_1 _2386_ (.A(net546),
    .B(_1452_),
    .Y(_1454_));
 sg13g2_xnor2_1 _2387_ (.Y(_1455_),
    .A(_0614_),
    .B(_1451_));
 sg13g2_a21oi_1 _2388_ (.A1(net632),
    .A2(_1455_),
    .Y(_1456_),
    .B1(_1454_));
 sg13g2_o21ai_1 _2389_ (.B1(_1456_),
    .Y(_1457_),
    .A1(_1448_),
    .A2(_1453_));
 sg13g2_a21oi_1 _2390_ (.A1(net580),
    .A2(_1450_),
    .Y(_1458_),
    .B1(net573));
 sg13g2_nor2_1 _2391_ (.A(_0491_),
    .B(_1458_),
    .Y(_1459_));
 sg13g2_xnor2_1 _2392_ (.Y(_1460_),
    .A(net568),
    .B(_1458_));
 sg13g2_xor2_1 _2393_ (.B(_1460_),
    .A(net621),
    .X(_1461_));
 sg13g2_o21ai_1 _2394_ (.B1(_1461_),
    .Y(_1462_),
    .A1(net633),
    .A2(_1455_));
 sg13g2_nand2b_1 _2395_ (.Y(_1463_),
    .B(_1457_),
    .A_N(_1462_));
 sg13g2_nor2b_1 _2396_ (.A(_1460_),
    .B_N(net627),
    .Y(_1464_));
 sg13g2_xnor2_1 _2397_ (.Y(_1465_),
    .A(net560),
    .B(_1459_));
 sg13g2_a21oi_1 _2398_ (.A1(net618),
    .A2(_1465_),
    .Y(_1466_),
    .B1(_1464_));
 sg13g2_nor2_1 _2399_ (.A(net618),
    .B(_1465_),
    .Y(_1467_));
 sg13g2_a221oi_1 _2400_ (.B2(_1466_),
    .C1(_1467_),
    .B1(_1463_),
    .A1(_0605_),
    .Y(_1468_),
    .A2(_1459_));
 sg13g2_a21oi_1 _2401_ (.A1(_1427_),
    .A2(_1429_),
    .Y(_1469_),
    .B1(_1468_));
 sg13g2_a21oi_2 _2402_ (.B1(net648),
    .Y(_1470_),
    .A2(_1132_),
    .A1(net656));
 sg13g2_nand2_1 _2403_ (.Y(_1471_),
    .A(net634),
    .B(_1470_));
 sg13g2_xnor2_1 _2404_ (.Y(_1472_),
    .A(net629),
    .B(_1471_));
 sg13g2_nor2_1 _2405_ (.A(net572),
    .B(_1472_),
    .Y(_1473_));
 sg13g2_nor2_1 _2406_ (.A(net650),
    .B(_1131_),
    .Y(_1474_));
 sg13g2_xnor2_1 _2407_ (.Y(_1475_),
    .A(_0036_),
    .B(_1474_));
 sg13g2_nor2_1 _2408_ (.A(net553),
    .B(_1475_),
    .Y(_1476_));
 sg13g2_nand2b_1 _2409_ (.Y(_1477_),
    .B(_1475_),
    .A_N(net582));
 sg13g2_nand2b_1 _2410_ (.Y(_1478_),
    .B(net582),
    .A_N(_1475_));
 sg13g2_xnor2_1 _2411_ (.Y(_1479_),
    .A(net549),
    .B(_1191_));
 sg13g2_or2_1 _2412_ (.X(_1480_),
    .B(_1479_),
    .A(_0666_));
 sg13g2_nor2b_1 _2413_ (.A(net613),
    .B_N(net689),
    .Y(_1481_));
 sg13g2_nand2_1 _2414_ (.Y(_1482_),
    .A(net688),
    .B(_0414_));
 sg13g2_a21oi_1 _2415_ (.A1(_1405_),
    .A2(_1482_),
    .Y(_1483_),
    .B1(_1404_));
 sg13g2_xnor2_1 _2416_ (.Y(_1484_),
    .A(_0535_),
    .B(net534));
 sg13g2_xnor2_1 _2417_ (.Y(_1485_),
    .A(_0675_),
    .B(_1484_));
 sg13g2_a22oi_1 _2418_ (.Y(_1486_),
    .B1(_1484_),
    .B2(net604),
    .A2(_1479_),
    .A1(net541));
 sg13g2_o21ai_1 _2419_ (.B1(_1486_),
    .Y(_1487_),
    .A1(_1483_),
    .A2(_1485_));
 sg13g2_nand3_1 _2420_ (.B(_1480_),
    .C(_1487_),
    .A(_0648_),
    .Y(_1488_));
 sg13g2_xnor2_1 _2421_ (.Y(_1489_),
    .A(net544),
    .B(_1131_));
 sg13g2_a21oi_2 _2422_ (.B1(net542),
    .Y(_1490_),
    .A2(_1487_),
    .A1(_1480_));
 sg13g2_a221oi_1 _2423_ (.B2(_1489_),
    .C1(_1490_),
    .B1(_1488_),
    .A1(_1477_),
    .Y(_1491_),
    .A2(_1478_));
 sg13g2_xnor2_1 _2424_ (.Y(_1492_),
    .A(net634),
    .B(_1470_));
 sg13g2_xnor2_1 _2425_ (.Y(_1493_),
    .A(net576),
    .B(_1492_));
 sg13g2_o21ai_1 _2426_ (.B1(_1493_),
    .Y(_1494_),
    .A1(_1476_),
    .A2(_1491_));
 sg13g2_a21o_1 _2427_ (.A2(_1470_),
    .A1(net546),
    .B1(_0557_),
    .X(_1495_));
 sg13g2_nand2_1 _2428_ (.Y(_1496_),
    .A(net623),
    .B(_1495_));
 sg13g2_xor2_1 _2429_ (.B(_1495_),
    .A(net623),
    .X(_1497_));
 sg13g2_nor2_1 _2430_ (.A(net564),
    .B(_1497_),
    .Y(_1498_));
 sg13g2_a22oi_1 _2431_ (.Y(_1499_),
    .B1(_1492_),
    .B2(net580),
    .A2(_1472_),
    .A1(net572));
 sg13g2_a21oi_1 _2432_ (.A1(_1494_),
    .A2(_1499_),
    .Y(_1500_),
    .B1(_1473_));
 sg13g2_xnor2_1 _2433_ (.Y(_1501_),
    .A(net537),
    .B(_1496_));
 sg13g2_a21oi_1 _2434_ (.A1(net564),
    .A2(_1497_),
    .Y(_1502_),
    .B1(_1501_));
 sg13g2_o21ai_1 _2435_ (.B1(_1502_),
    .Y(_1503_),
    .A1(_1498_),
    .A2(_1500_));
 sg13g2_nand2b_1 _2436_ (.Y(_1504_),
    .B(net641),
    .A_N(_0822_));
 sg13g2_nor2_1 _2437_ (.A(net629),
    .B(_1504_),
    .Y(_1505_));
 sg13g2_xnor2_1 _2438_ (.Y(_1506_),
    .A(net625),
    .B(_1505_));
 sg13g2_or2_1 _2439_ (.X(_1507_),
    .B(_1504_),
    .A(_0771_));
 sg13g2_xnor2_1 _2440_ (.Y(_1508_),
    .A(net537),
    .B(_1507_));
 sg13g2_a21oi_1 _2441_ (.A1(net564),
    .A2(_1506_),
    .Y(_1509_),
    .B1(_1508_));
 sg13g2_xnor2_1 _2442_ (.Y(_1510_),
    .A(net632),
    .B(_1504_));
 sg13g2_nor2_1 _2443_ (.A(net563),
    .B(_1506_),
    .Y(_1511_));
 sg13g2_a21oi_1 _2444_ (.A1(net572),
    .A2(_1510_),
    .Y(_1512_),
    .B1(_1511_));
 sg13g2_nor2_1 _2445_ (.A(net572),
    .B(_1510_),
    .Y(_1513_));
 sg13g2_xnor2_1 _2446_ (.Y(_1514_),
    .A(_0629_),
    .B(_0822_));
 sg13g2_xnor2_1 _2447_ (.Y(_1515_),
    .A(net575),
    .B(_1514_));
 sg13g2_nor2_1 _2448_ (.A(_0821_),
    .B(_1081_),
    .Y(_1516_));
 sg13g2_nor3_2 _2449_ (.A(net587),
    .B(_0821_),
    .C(_1081_),
    .Y(_1517_));
 sg13g2_nor2_1 _2450_ (.A(net542),
    .B(_1516_),
    .Y(_1518_));
 sg13g2_nor2_1 _2451_ (.A(_1517_),
    .B(_1518_),
    .Y(_1519_));
 sg13g2_nor2_1 _2452_ (.A(_0822_),
    .B(_1113_),
    .Y(_1520_));
 sg13g2_xnor2_1 _2453_ (.Y(_1521_),
    .A(net583),
    .B(_1520_));
 sg13g2_nor2_1 _2454_ (.A(_1519_),
    .B(_1521_),
    .Y(_1522_));
 sg13g2_a21oi_1 _2455_ (.A1(_0847_),
    .A2(_0850_),
    .Y(_1523_),
    .B1(_0857_));
 sg13g2_nand3_1 _2456_ (.B(net526),
    .C(_1523_),
    .A(_0848_),
    .Y(_1524_));
 sg13g2_nand3_1 _2457_ (.B(net678),
    .C(net526),
    .A(net603),
    .Y(_1525_));
 sg13g2_nand3_1 _2458_ (.B(_1524_),
    .C(_1525_),
    .A(_0855_),
    .Y(_1526_));
 sg13g2_nor3_1 _2459_ (.A(net587),
    .B(_1516_),
    .C(_1521_),
    .Y(_1527_));
 sg13g2_nor2_1 _2460_ (.A(net553),
    .B(_1520_),
    .Y(_1528_));
 sg13g2_a21oi_1 _2461_ (.A1(_1522_),
    .A2(_1526_),
    .Y(_1529_),
    .B1(_1528_));
 sg13g2_nand2b_1 _2462_ (.Y(_1530_),
    .B(_1529_),
    .A_N(_1527_));
 sg13g2_a22oi_1 _2463_ (.Y(_1531_),
    .B1(_1515_),
    .B2(_1530_),
    .A2(_1514_),
    .A1(net580));
 sg13g2_o21ai_1 _2464_ (.B1(_1512_),
    .Y(_0082_),
    .A1(_1513_),
    .A2(_1531_));
 sg13g2_a21o_1 _2465_ (.A2(_0082_),
    .A1(_1509_),
    .B1(net561),
    .X(_0083_));
 sg13g2_nand2_2 _2466_ (.Y(_0084_),
    .A(net526),
    .B(_0875_));
 sg13g2_nor2_1 _2467_ (.A(_1513_),
    .B(_0084_),
    .Y(_0085_));
 sg13g2_and2_1 _2468_ (.A(_1515_),
    .B(_1522_),
    .X(_0086_));
 sg13g2_nand4_1 _2469_ (.B(_1512_),
    .C(_0085_),
    .A(_1509_),
    .Y(_0087_),
    .D(_0086_));
 sg13g2_nand2_1 _2470_ (.Y(_0088_),
    .A(net561),
    .B(_1496_));
 sg13g2_nand4_1 _2471_ (.B(_1507_),
    .C(_0087_),
    .A(net615),
    .Y(_0089_),
    .D(_0088_));
 sg13g2_nand3b_1 _2472_ (.B(_0083_),
    .C(_1503_),
    .Y(_0090_),
    .A_N(_0089_));
 sg13g2_o21ai_1 _2473_ (.B1(_0932_),
    .Y(_0091_),
    .A1(net555),
    .A2(net554));
 sg13g2_o21ai_1 _2474_ (.B1(net567),
    .Y(_0092_),
    .A1(_1450_),
    .A2(_0091_));
 sg13g2_a21oi_2 _2475_ (.B1(net586),
    .Y(_0093_),
    .A2(net590),
    .A1(net596));
 sg13g2_o21ai_1 _2476_ (.B1(_1056_),
    .Y(_0094_),
    .A1(_0700_),
    .A2(_0093_));
 sg13g2_mux2_1 _2477_ (.A0(_0018_),
    .A1(net7),
    .S(net529),
    .X(_0095_));
 sg13g2_nand4_1 _2478_ (.B(_0092_),
    .C(_0094_),
    .A(_0502_),
    .Y(_0096_),
    .D(_0095_));
 sg13g2_nor2_1 _2479_ (.A(_0090_),
    .B(_0096_),
    .Y(_0097_));
 sg13g2_nor2_1 _2480_ (.A(_0829_),
    .B(_1295_),
    .Y(_0098_));
 sg13g2_nor3_2 _2481_ (.A(net547),
    .B(net643),
    .C(_0098_),
    .Y(_0099_));
 sg13g2_nor2_2 _2482_ (.A(net631),
    .B(_0099_),
    .Y(_0100_));
 sg13g2_nor2_1 _2483_ (.A(net621),
    .B(_0100_),
    .Y(_0101_));
 sg13g2_xnor2_1 _2484_ (.Y(_0102_),
    .A(net618),
    .B(_0101_));
 sg13g2_nand2b_1 _2485_ (.Y(_0103_),
    .B(net561),
    .A_N(_0102_));
 sg13g2_xor2_1 _2486_ (.B(_0100_),
    .A(net627),
    .X(_0104_));
 sg13g2_nor2_1 _2487_ (.A(net564),
    .B(_0104_),
    .Y(_0105_));
 sg13g2_nor2_1 _2488_ (.A(net635),
    .B(_1396_),
    .Y(_0106_));
 sg13g2_xnor2_1 _2489_ (.Y(_0107_),
    .A(net629),
    .B(_0106_));
 sg13g2_nand2b_1 _2490_ (.Y(_0108_),
    .B(net572),
    .A_N(_0107_));
 sg13g2_o21ai_1 _2491_ (.B1(net650),
    .Y(_0109_),
    .A1(net550),
    .A2(_0820_));
 sg13g2_xnor2_1 _2492_ (.Y(_0110_),
    .A(net651),
    .B(_1296_));
 sg13g2_nand2_1 _2493_ (.Y(_0111_),
    .A(net542),
    .B(_0110_));
 sg13g2_a22oi_1 _2494_ (.Y(_0112_),
    .B1(_1481_),
    .B2(_0847_),
    .A2(_1122_),
    .A1(net555));
 sg13g2_xnor2_1 _2495_ (.Y(_0113_),
    .A(net659),
    .B(_1205_));
 sg13g2_nor2_1 _2496_ (.A(_0436_),
    .B(_1222_),
    .Y(_0114_));
 sg13g2_a221oi_1 _2497_ (.B2(net598),
    .C1(_0114_),
    .B1(_0113_),
    .A1(_1407_),
    .Y(_0115_),
    .A2(_0112_));
 sg13g2_nor2_1 _2498_ (.A(net598),
    .B(_0113_),
    .Y(_0116_));
 sg13g2_o21ai_1 _2499_ (.B1(_0111_),
    .Y(_0117_),
    .A1(_0115_),
    .A2(_0116_));
 sg13g2_xnor2_1 _2500_ (.Y(_0118_),
    .A(_0639_),
    .B(_0109_));
 sg13g2_xnor2_1 _2501_ (.Y(_0119_),
    .A(net583),
    .B(_0118_));
 sg13g2_nor2_1 _2502_ (.A(net542),
    .B(_0110_),
    .Y(_0120_));
 sg13g2_nor2_1 _2503_ (.A(_0119_),
    .B(_0120_),
    .Y(_0121_));
 sg13g2_nand2b_1 _2504_ (.Y(_0122_),
    .B(net586),
    .A_N(_0118_));
 sg13g2_o21ai_1 _2505_ (.B1(_0122_),
    .Y(_0123_),
    .A1(_0447_),
    .A2(_1398_));
 sg13g2_a21oi_2 _2506_ (.B1(_0123_),
    .Y(_0124_),
    .A2(_0121_),
    .A1(_0117_));
 sg13g2_nor3_1 _2507_ (.A(net580),
    .B(net577),
    .C(_1398_),
    .Y(_0125_));
 sg13g2_a21o_1 _2508_ (.A2(_1398_),
    .A1(net577),
    .B1(_0125_),
    .X(_0126_));
 sg13g2_o21ai_1 _2509_ (.B1(_0108_),
    .Y(_0127_),
    .A1(_0124_),
    .A2(_0126_));
 sg13g2_a22oi_1 _2510_ (.Y(_0128_),
    .B1(_0107_),
    .B2(_0458_),
    .A2(_0104_),
    .A1(net565));
 sg13g2_a21oi_1 _2511_ (.A1(_0127_),
    .A2(_0128_),
    .Y(_0129_),
    .B1(_0105_));
 sg13g2_xnor2_1 _2512_ (.Y(_0130_),
    .A(_0028_),
    .B(_0102_));
 sg13g2_o21ai_1 _2513_ (.B1(_0103_),
    .Y(_0131_),
    .A1(_0129_),
    .A2(_0130_));
 sg13g2_o21ai_1 _2514_ (.B1(_0131_),
    .Y(_0132_),
    .A1(_0706_),
    .A2(_0100_));
 sg13g2_nand2_2 _2515_ (.Y(_0133_),
    .A(_0709_),
    .B(_1082_));
 sg13g2_nand2_1 _2516_ (.Y(_0134_),
    .A(net631),
    .B(_0133_));
 sg13g2_a21oi_1 _2517_ (.A1(net630),
    .A2(_0133_),
    .Y(_0135_),
    .B1(net624));
 sg13g2_xnor2_1 _2518_ (.Y(_0136_),
    .A(net617),
    .B(_0135_));
 sg13g2_xor2_1 _2519_ (.B(_0134_),
    .A(net620),
    .X(_0137_));
 sg13g2_xnor2_1 _2520_ (.Y(_0138_),
    .A(_0605_),
    .B(_0136_));
 sg13g2_a21oi_1 _2521_ (.A1(net563),
    .A2(_0137_),
    .Y(_0139_),
    .B1(_0138_));
 sg13g2_xnor2_1 _2522_ (.Y(_0140_),
    .A(net628),
    .B(_0133_));
 sg13g2_nor2_1 _2523_ (.A(net563),
    .B(_0137_),
    .Y(_0141_));
 sg13g2_a21oi_1 _2524_ (.A1(net573),
    .A2(_0140_),
    .Y(_0142_),
    .B1(_0141_));
 sg13g2_nor2_1 _2525_ (.A(net573),
    .B(_0140_),
    .Y(_0143_));
 sg13g2_xnor2_1 _2526_ (.Y(_0144_),
    .A(net547),
    .B(_1117_));
 sg13g2_nor2_1 _2527_ (.A(_0447_),
    .B(_0144_),
    .Y(_0145_));
 sg13g2_xor2_1 _2528_ (.B(_0144_),
    .A(net575),
    .X(_0146_));
 sg13g2_xnor2_1 _2529_ (.Y(_0147_),
    .A(net643),
    .B(_1081_));
 sg13g2_xnor2_1 _2530_ (.Y(_0148_),
    .A(net582),
    .B(_0147_));
 sg13g2_nor2_1 _2531_ (.A(_1518_),
    .B(_0148_),
    .Y(_0149_));
 sg13g2_o21ai_1 _2532_ (.B1(_0149_),
    .Y(_0150_),
    .A1(_1517_),
    .A2(_1526_));
 sg13g2_o21ai_1 _2533_ (.B1(_0150_),
    .Y(_0151_),
    .A1(net553),
    .A2(_0147_));
 sg13g2_a21oi_1 _2534_ (.A1(_0146_),
    .A2(_0151_),
    .Y(_0152_),
    .B1(_0145_));
 sg13g2_o21ai_1 _2535_ (.B1(_0142_),
    .Y(_0153_),
    .A1(_0143_),
    .A2(_0152_));
 sg13g2_a22oi_1 _2536_ (.Y(_0154_),
    .B1(_0139_),
    .B2(_0153_),
    .A2(_0136_),
    .A1(net561));
 sg13g2_nand3_1 _2537_ (.B(_0875_),
    .C(_1519_),
    .A(net526),
    .Y(_0155_));
 sg13g2_nor3_1 _2538_ (.A(_0143_),
    .B(_0148_),
    .C(_0155_),
    .Y(_0156_));
 sg13g2_nand4_1 _2539_ (.B(_0142_),
    .C(_0146_),
    .A(_0139_),
    .Y(_0157_),
    .D(_0156_));
 sg13g2_o21ai_1 _2540_ (.B1(_0157_),
    .Y(_0158_),
    .A1(net615),
    .A2(_0135_));
 sg13g2_nor2_1 _2541_ (.A(_0154_),
    .B(_0158_),
    .Y(_0159_));
 sg13g2_nand2_2 _2542_ (.Y(_0160_),
    .A(_0132_),
    .B(_0159_));
 sg13g2_or4_1 _2543_ (.A(net618),
    .B(net641),
    .C(_0771_),
    .D(net538),
    .X(_0161_));
 sg13g2_nand2b_1 _2544_ (.Y(_0162_),
    .B(net529),
    .A_N(net3));
 sg13g2_o21ai_1 _2545_ (.B1(_0162_),
    .Y(_0163_),
    .A1(net528),
    .A2(_0014_));
 sg13g2_nor3_1 _2546_ (.A(_0160_),
    .B(_0161_),
    .C(_0163_),
    .Y(_0164_));
 sg13g2_o21ai_1 _2547_ (.B1(_1469_),
    .Y(_0165_),
    .A1(_0097_),
    .A2(_0164_));
 sg13g2_nor3_1 _2548_ (.A(_0771_),
    .B(_0803_),
    .C(_0821_),
    .Y(_0166_));
 sg13g2_nor2_1 _2549_ (.A(_0597_),
    .B(_0166_),
    .Y(_0167_));
 sg13g2_nand2_1 _2550_ (.Y(_0168_),
    .A(net561),
    .B(_0167_));
 sg13g2_nor3_2 _2551_ (.A(net628),
    .B(_0803_),
    .C(_0821_),
    .Y(_0169_));
 sg13g2_o21ai_1 _2552_ (.B1(net628),
    .Y(_0170_),
    .A1(_0803_),
    .A2(_0821_));
 sg13g2_nor2b_1 _2553_ (.A(_0169_),
    .B_N(_0170_),
    .Y(_0171_));
 sg13g2_xnor2_1 _2554_ (.Y(_0172_),
    .A(_0834_),
    .B(_0169_));
 sg13g2_a21oi_1 _2555_ (.A1(_0458_),
    .A2(_0171_),
    .Y(_0173_),
    .B1(_0172_));
 sg13g2_xnor2_1 _2556_ (.Y(_0174_),
    .A(_0629_),
    .B(_1113_));
 sg13g2_xnor2_1 _2557_ (.Y(_0175_),
    .A(net575),
    .B(_0174_));
 sg13g2_o21ai_1 _2558_ (.B1(_1435_),
    .Y(_0176_),
    .A1(_1433_),
    .A2(_1481_));
 sg13g2_nor2b_1 _2559_ (.A(_1438_),
    .B_N(_0176_),
    .Y(_0177_));
 sg13g2_nor3_1 _2560_ (.A(net554),
    .B(net678),
    .C(net526),
    .Y(_0178_));
 sg13g2_nor4_1 _2561_ (.A(_1432_),
    .B(_1517_),
    .C(_0177_),
    .D(_0178_),
    .Y(_0179_));
 sg13g2_nor3_1 _2562_ (.A(_1518_),
    .B(_1521_),
    .C(_0179_),
    .Y(_0180_));
 sg13g2_o21ai_1 _2563_ (.B1(_0175_),
    .Y(_0181_),
    .A1(_1528_),
    .A2(_0180_));
 sg13g2_nand2b_1 _2564_ (.Y(_0182_),
    .B(net572),
    .A_N(_0171_));
 sg13g2_nand2_1 _2565_ (.Y(_0183_),
    .A(net579),
    .B(_0174_));
 sg13g2_nand3_1 _2566_ (.B(_0182_),
    .C(_0183_),
    .A(_0181_),
    .Y(_0184_));
 sg13g2_xor2_1 _2567_ (.B(_0169_),
    .A(net621),
    .X(_0185_));
 sg13g2_a22oi_1 _2568_ (.Y(_0186_),
    .B1(_0185_),
    .B2(net568),
    .A2(_0184_),
    .A1(_0173_));
 sg13g2_nand3b_1 _2569_ (.B(_0852_),
    .C(_0849_),
    .Y(_0187_),
    .A_N(_1438_));
 sg13g2_nor4_1 _2570_ (.A(_1517_),
    .B(_1518_),
    .C(_1521_),
    .D(_0187_),
    .Y(_0188_));
 sg13g2_and4_1 _2571_ (.A(_0173_),
    .B(_0175_),
    .C(_0182_),
    .D(_0188_),
    .X(_0189_));
 sg13g2_o21ai_1 _2572_ (.B1(_0168_),
    .Y(_0190_),
    .A1(_0186_),
    .A2(_0189_));
 sg13g2_nor2_2 _2573_ (.A(net552),
    .B(_1430_),
    .Y(_0191_));
 sg13g2_o21ai_1 _2574_ (.B1(net586),
    .Y(_0192_),
    .A1(net596),
    .A2(net589));
 sg13g2_nand3_1 _2575_ (.B(_0614_),
    .C(_0191_),
    .A(net579),
    .Y(_0193_));
 sg13g2_xnor2_1 _2576_ (.Y(_0194_),
    .A(_0491_),
    .B(_0193_));
 sg13g2_nor3_1 _2577_ (.A(net568),
    .B(_0700_),
    .C(_0192_),
    .Y(_0195_));
 sg13g2_nand2b_2 _2578_ (.Y(_0196_),
    .B(net565),
    .A_N(_0195_));
 sg13g2_xnor2_1 _2579_ (.Y(_0197_),
    .A(_0844_),
    .B(_0196_));
 sg13g2_a21o_1 _2580_ (.A2(_0194_),
    .A1(net622),
    .B1(_0197_),
    .X(_0198_));
 sg13g2_o21ai_1 _2581_ (.B1(_0030_),
    .Y(_0199_),
    .A1(_0447_),
    .A2(_0192_));
 sg13g2_and2_1 _2582_ (.A(_0193_),
    .B(_0199_),
    .X(_0200_));
 sg13g2_nand2_1 _2583_ (.Y(_0201_),
    .A(_0557_),
    .B(_0200_));
 sg13g2_nand2b_1 _2584_ (.Y(_0202_),
    .B(net632),
    .A_N(_0200_));
 sg13g2_xnor2_1 _2585_ (.Y(_0203_),
    .A(net577),
    .B(_0192_));
 sg13g2_xnor2_1 _2586_ (.Y(_0204_),
    .A(net634),
    .B(_0203_));
 sg13g2_nand3_1 _2587_ (.B(_0202_),
    .C(_0204_),
    .A(_0201_),
    .Y(_0205_));
 sg13g2_nor2_2 _2588_ (.A(_1449_),
    .B(_0191_),
    .Y(_0206_));
 sg13g2_inv_1 _2589_ (.Y(_0207_),
    .A(_0206_));
 sg13g2_xnor2_1 _2590_ (.Y(_0208_),
    .A(net643),
    .B(_0206_));
 sg13g2_xnor2_1 _2591_ (.Y(_0209_),
    .A(net544),
    .B(_1442_));
 sg13g2_nand2b_1 _2592_ (.Y(_0210_),
    .B(_0209_),
    .A_N(_0208_));
 sg13g2_nor2_1 _2593_ (.A(_0205_),
    .B(_0210_),
    .Y(_0211_));
 sg13g2_nor2b_1 _2594_ (.A(_1440_),
    .B_N(_0211_),
    .Y(_0212_));
 sg13g2_and3_1 _2595_ (.X(_0213_),
    .A(net642),
    .B(_0201_),
    .C(_0203_));
 sg13g2_nor2_1 _2596_ (.A(net621),
    .B(_0194_),
    .Y(_0214_));
 sg13g2_o21ai_1 _2597_ (.B1(_0202_),
    .Y(_0215_),
    .A1(net621),
    .A2(_0194_));
 sg13g2_nor2_1 _2598_ (.A(_1444_),
    .B(_0208_),
    .Y(_0216_));
 sg13g2_a21oi_1 _2599_ (.A1(net648),
    .A2(_0207_),
    .Y(_0217_),
    .B1(_0216_));
 sg13g2_nor2_1 _2600_ (.A(_0205_),
    .B(_0217_),
    .Y(_0218_));
 sg13g2_nor4_1 _2601_ (.A(_0212_),
    .B(_0213_),
    .C(_0215_),
    .D(_0218_),
    .Y(_0219_));
 sg13g2_a21oi_1 _2602_ (.A1(_0605_),
    .A2(_0196_),
    .Y(_0220_),
    .B1(_0513_));
 sg13g2_o21ai_1 _2603_ (.B1(_0220_),
    .Y(_0221_),
    .A1(_0605_),
    .A2(_0196_));
 sg13g2_o21ai_1 _2604_ (.B1(_0221_),
    .Y(_0222_),
    .A1(_0198_),
    .A2(_0219_));
 sg13g2_nor3_1 _2605_ (.A(_0187_),
    .B(_0198_),
    .C(_0214_),
    .Y(_0223_));
 sg13g2_a21oi_1 _2606_ (.A1(_0167_),
    .A2(_0196_),
    .Y(_0224_),
    .B1(net560));
 sg13g2_a221oi_1 _2607_ (.B2(_0223_),
    .C1(_0224_),
    .B1(_0211_),
    .A1(_0597_),
    .Y(_0225_),
    .A2(_0166_));
 sg13g2_nand3_1 _2608_ (.B(_0222_),
    .C(_0225_),
    .A(_0190_),
    .Y(_0226_));
 sg13g2_mux2_1 _2609_ (.A0(_0015_),
    .A1(net4),
    .S(net529),
    .X(_0227_));
 sg13g2_nand2_1 _2610_ (.Y(_0228_),
    .A(_0719_),
    .B(_0227_));
 sg13g2_nand3_1 _2611_ (.B(net554),
    .C(_0930_),
    .A(net596),
    .Y(_0229_));
 sg13g2_and2_1 _2612_ (.A(net541),
    .B(_0229_),
    .X(_0230_));
 sg13g2_nor2b_1 _2613_ (.A(_0701_),
    .B_N(_0230_),
    .Y(_0231_));
 sg13g2_o21ai_1 _2614_ (.B1(_0699_),
    .Y(_0232_),
    .A1(net579),
    .A2(_0191_));
 sg13g2_nor2_1 _2615_ (.A(net585),
    .B(_0480_),
    .Y(_0233_));
 sg13g2_nand2_1 _2616_ (.Y(_0234_),
    .A(net552),
    .B(net590));
 sg13g2_nor4_2 _2617_ (.A(_0700_),
    .B(_0703_),
    .C(_0229_),
    .Y(_0235_),
    .D(_0234_));
 sg13g2_nand2b_1 _2618_ (.Y(_0236_),
    .B(net528),
    .A_N(net2));
 sg13g2_o21ai_1 _2619_ (.B1(_0236_),
    .Y(_0237_),
    .A1(net528),
    .A2(_0013_));
 sg13g2_nor3_1 _2620_ (.A(_0090_),
    .B(_0161_),
    .C(_0237_),
    .Y(_0238_));
 sg13g2_and2_1 _2621_ (.A(_0928_),
    .B(_0230_),
    .X(_0239_));
 sg13g2_nand2b_1 _2622_ (.Y(_0240_),
    .B(net528),
    .A_N(net1));
 sg13g2_or4_1 _2623_ (.A(net581),
    .B(net574),
    .C(net536),
    .D(_0229_),
    .X(_0241_));
 sg13g2_o21ai_1 _2624_ (.B1(_0240_),
    .Y(_0242_),
    .A1(_0012_),
    .A2(net528));
 sg13g2_a21oi_1 _2625_ (.A1(_1056_),
    .A2(_1449_),
    .Y(_0243_),
    .B1(_0242_));
 sg13g2_nand4_1 _2626_ (.B(_0932_),
    .C(_0241_),
    .A(_0927_),
    .Y(_0244_),
    .D(_0243_));
 sg13g2_nand2_2 _2627_ (.Y(_0245_),
    .A(net539),
    .B(_1131_));
 sg13g2_nand2b_1 _2628_ (.Y(_0246_),
    .B(_0245_),
    .A_N(_0714_));
 sg13g2_a21o_1 _2629_ (.A2(_0245_),
    .A1(net641),
    .B1(net632),
    .X(_0247_));
 sg13g2_and2_1 _2630_ (.A(_0246_),
    .B(_0247_),
    .X(_0248_));
 sg13g2_xnor2_1 _2631_ (.Y(_0249_),
    .A(net635),
    .B(_0245_));
 sg13g2_nand2_1 _2632_ (.Y(_0250_),
    .A(net580),
    .B(_0249_));
 sg13g2_nand2_1 _2633_ (.Y(_0251_),
    .A(net650),
    .B(_1131_));
 sg13g2_xnor2_1 _2634_ (.Y(_0252_),
    .A(_0577_),
    .B(_0251_));
 sg13g2_inv_1 _2635_ (.Y(_0253_),
    .A(_0252_));
 sg13g2_nand3b_1 _2636_ (.B(_1488_),
    .C(_0251_),
    .Y(_0254_),
    .A_N(_1474_));
 sg13g2_xnor2_1 _2637_ (.Y(_0255_),
    .A(net583),
    .B(_0252_));
 sg13g2_nor2_1 _2638_ (.A(_1490_),
    .B(_0255_),
    .Y(_0256_));
 sg13g2_a22oi_1 _2639_ (.Y(_0257_),
    .B1(_0254_),
    .B2(_0256_),
    .A2(_0253_),
    .A1(net586));
 sg13g2_xor2_1 _2640_ (.B(_0249_),
    .A(net576),
    .X(_0258_));
 sg13g2_o21ai_1 _2641_ (.B1(_0250_),
    .Y(_0259_),
    .A1(_0257_),
    .A2(_0258_));
 sg13g2_o21ai_1 _2642_ (.B1(_0259_),
    .Y(_0260_),
    .A1(net572),
    .A2(_0248_));
 sg13g2_xor2_1 _2643_ (.B(_0246_),
    .A(net627),
    .X(_0261_));
 sg13g2_nor2_1 _2644_ (.A(net565),
    .B(_0261_),
    .Y(_0262_));
 sg13g2_a21oi_1 _2645_ (.A1(net573),
    .A2(_0248_),
    .Y(_0263_),
    .B1(_0262_));
 sg13g2_nor2_1 _2646_ (.A(net621),
    .B(_0246_),
    .Y(_0264_));
 sg13g2_xnor2_1 _2647_ (.Y(_0265_),
    .A(net537),
    .B(_0264_));
 sg13g2_a22oi_1 _2648_ (.Y(_0266_),
    .B1(_0263_),
    .B2(_0260_),
    .A2(_0261_),
    .A1(net565));
 sg13g2_and3_2 _2649_ (.X(_0267_),
    .A(net596),
    .B(net586),
    .C(net589));
 sg13g2_nand2_1 _2650_ (.Y(_0268_),
    .A(net580),
    .B(_0267_));
 sg13g2_nor2_1 _2651_ (.A(net569),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_xnor2_1 _2652_ (.Y(_0270_),
    .A(net566),
    .B(_0269_));
 sg13g2_nor2b_1 _2653_ (.A(_0700_),
    .B_N(_0267_),
    .Y(_0271_));
 sg13g2_nor2_1 _2654_ (.A(net568),
    .B(_0271_),
    .Y(_0272_));
 sg13g2_xnor2_1 _2655_ (.Y(_0273_),
    .A(net537),
    .B(_0272_));
 sg13g2_a21o_1 _2656_ (.A2(_0270_),
    .A1(net621),
    .B1(_0273_),
    .X(_0274_));
 sg13g2_a21oi_1 _2657_ (.A1(_0458_),
    .A2(_0268_),
    .Y(_0275_),
    .B1(_0271_));
 sg13g2_nand2_1 _2658_ (.Y(_0276_),
    .A(net632),
    .B(_0275_));
 sg13g2_o21ai_1 _2659_ (.B1(_0276_),
    .Y(_0277_),
    .A1(net622),
    .A2(_0270_));
 sg13g2_or2_1 _2660_ (.X(_0278_),
    .B(_0275_),
    .A(net632));
 sg13g2_nand3_1 _2661_ (.B(_1524_),
    .C(_1525_),
    .A(_0854_),
    .Y(_0279_));
 sg13g2_nor2_1 _2662_ (.A(net583),
    .B(_1441_),
    .Y(_0280_));
 sg13g2_xnor2_1 _2663_ (.Y(_0281_),
    .A(_0447_),
    .B(_0280_));
 sg13g2_xnor2_1 _2664_ (.Y(_0282_),
    .A(_0629_),
    .B(_0281_));
 sg13g2_nor2_2 _2665_ (.A(_0093_),
    .B(_0267_),
    .Y(_0283_));
 sg13g2_xnor2_1 _2666_ (.Y(_0284_),
    .A(net643),
    .B(_0283_));
 sg13g2_nand2_1 _2667_ (.Y(_0285_),
    .A(_0209_),
    .B(_0284_));
 sg13g2_inv_1 _2668_ (.Y(_0286_),
    .A(_0285_));
 sg13g2_nand2_1 _2669_ (.Y(_0287_),
    .A(net641),
    .B(_0281_));
 sg13g2_a221oi_1 _2670_ (.B2(_0279_),
    .C1(_0216_),
    .B1(_0286_),
    .A1(net648),
    .Y(_0288_),
    .A2(_0283_));
 sg13g2_o21ai_1 _2671_ (.B1(_0287_),
    .Y(_0289_),
    .A1(_0282_),
    .A2(_0288_));
 sg13g2_a21oi_1 _2672_ (.A1(_0278_),
    .A2(_0289_),
    .Y(_0290_),
    .B1(_0277_));
 sg13g2_o21ai_1 _2673_ (.B1(_0513_),
    .Y(_0291_),
    .A1(_0274_),
    .A2(_0290_));
 sg13g2_o21ai_1 _2674_ (.B1(net560),
    .Y(_0292_),
    .A1(net616),
    .A2(_0264_));
 sg13g2_a21oi_1 _2675_ (.A1(net616),
    .A2(_0264_),
    .Y(_0293_),
    .B1(_0292_));
 sg13g2_a21oi_1 _2676_ (.A1(_0265_),
    .A2(_0266_),
    .Y(_0294_),
    .B1(_0293_));
 sg13g2_nand2b_1 _2677_ (.Y(_0295_),
    .B(_0286_),
    .A_N(_0084_));
 sg13g2_nand2b_1 _2678_ (.Y(_0296_),
    .B(_0278_),
    .A_N(_0282_));
 sg13g2_nor4_1 _2679_ (.A(_0274_),
    .B(_0277_),
    .C(_0295_),
    .D(_0296_),
    .Y(_0297_));
 sg13g2_nor2_1 _2680_ (.A(_0271_),
    .B(_0297_),
    .Y(_0298_));
 sg13g2_nand3_1 _2681_ (.B(_0291_),
    .C(_0298_),
    .A(_1056_),
    .Y(_0299_));
 sg13g2_nor3_1 _2682_ (.A(_0239_),
    .B(_0244_),
    .C(_0299_),
    .Y(_0300_));
 sg13g2_and2_1 _2683_ (.A(_0294_),
    .B(_0300_),
    .X(_0301_));
 sg13g2_o21ai_1 _2684_ (.B1(net593),
    .Y(_0302_),
    .A1(net596),
    .A2(_0939_));
 sg13g2_nor2_1 _2685_ (.A(net590),
    .B(_0302_),
    .Y(_0303_));
 sg13g2_o21ai_1 _2686_ (.B1(net581),
    .Y(_0304_),
    .A1(_0971_),
    .A2(_0302_));
 sg13g2_o21ai_1 _2687_ (.B1(net570),
    .Y(_0305_),
    .A1(net574),
    .A2(_0304_));
 sg13g2_and2_1 _2688_ (.A(net567),
    .B(_0305_),
    .X(_0306_));
 sg13g2_xnor2_1 _2689_ (.Y(_0307_),
    .A(_0605_),
    .B(_0306_));
 sg13g2_xnor2_1 _2690_ (.Y(_0308_),
    .A(_0491_),
    .B(_0305_));
 sg13g2_nor2b_1 _2691_ (.A(_0308_),
    .B_N(net627),
    .Y(_0309_));
 sg13g2_xnor2_1 _2692_ (.Y(_0310_),
    .A(_0458_),
    .B(_0304_));
 sg13g2_xnor2_1 _2693_ (.Y(_0311_),
    .A(net622),
    .B(_0308_));
 sg13g2_a21oi_1 _2694_ (.A1(_0557_),
    .A2(_0310_),
    .Y(_0312_),
    .B1(_0311_));
 sg13g2_xnor2_1 _2695_ (.Y(_0313_),
    .A(net583),
    .B(_0303_));
 sg13g2_nor2_1 _2696_ (.A(_0577_),
    .B(_0313_),
    .Y(_0314_));
 sg13g2_a21oi_1 _2697_ (.A1(net525),
    .A2(_1012_),
    .Y(_0315_),
    .B1(net668));
 sg13g2_xnor2_1 _2698_ (.Y(_0316_),
    .A(net554),
    .B(_0937_));
 sg13g2_nand2_1 _2699_ (.Y(_0317_),
    .A(_0937_),
    .B(_0176_));
 sg13g2_xnor2_1 _2700_ (.Y(_0318_),
    .A(_0040_),
    .B(_0316_));
 sg13g2_a22oi_1 _2701_ (.Y(_0319_),
    .B1(_0317_),
    .B2(_0318_),
    .A2(_0316_),
    .A1(net678));
 sg13g2_or2_1 _2702_ (.X(_0320_),
    .B(_0319_),
    .A(_0315_));
 sg13g2_and3_1 _2703_ (.X(_0321_),
    .A(net668),
    .B(net525),
    .C(_1012_));
 sg13g2_xnor2_1 _2704_ (.Y(_0322_),
    .A(net542),
    .B(_0302_));
 sg13g2_or2_1 _2705_ (.X(_0323_),
    .B(_0322_),
    .A(net651));
 sg13g2_nor2b_1 _2706_ (.A(_0321_),
    .B_N(_0323_),
    .Y(_0324_));
 sg13g2_nor2_1 _2707_ (.A(_0315_),
    .B(_0321_),
    .Y(_0325_));
 sg13g2_xnor2_1 _2708_ (.Y(_0326_),
    .A(_0036_),
    .B(_0313_));
 sg13g2_nand2_1 _2709_ (.Y(_0327_),
    .A(net651),
    .B(_0322_));
 sg13g2_a21oi_1 _2710_ (.A1(_0320_),
    .A2(_0324_),
    .Y(_0328_),
    .B1(_0326_));
 sg13g2_a21oi_1 _2711_ (.A1(_0327_),
    .A2(_0328_),
    .Y(_0329_),
    .B1(_0314_));
 sg13g2_nand3_1 _2712_ (.B(net553),
    .C(_0303_),
    .A(_0447_),
    .Y(_0330_));
 sg13g2_nand2_1 _2713_ (.Y(_0331_),
    .A(_0304_),
    .B(_0330_));
 sg13g2_xnor2_1 _2714_ (.Y(_0332_),
    .A(_0629_),
    .B(_0331_));
 sg13g2_nor2_1 _2715_ (.A(_0557_),
    .B(_0310_),
    .Y(_0333_));
 sg13g2_a21oi_1 _2716_ (.A1(net638),
    .A2(_0331_),
    .Y(_0334_),
    .B1(_0333_));
 sg13g2_o21ai_1 _2717_ (.B1(_0334_),
    .Y(_0335_),
    .A1(_0329_),
    .A2(_0332_));
 sg13g2_a21oi_1 _2718_ (.A1(_0312_),
    .A2(_0335_),
    .Y(_0336_),
    .B1(_0309_));
 sg13g2_inv_1 _2719_ (.Y(_0337_),
    .A(_0336_));
 sg13g2_nor2_1 _2720_ (.A(net619),
    .B(_0307_),
    .Y(_0338_));
 sg13g2_nand2_1 _2721_ (.Y(_0339_),
    .A(_0849_),
    .B(_1481_));
 sg13g2_o21ai_1 _2722_ (.B1(_0339_),
    .Y(_0340_),
    .A1(_0849_),
    .A2(_1434_));
 sg13g2_and3_1 _2723_ (.X(_0341_),
    .A(_0323_),
    .B(_0327_),
    .C(_0340_));
 sg13g2_nor3_1 _2724_ (.A(_0326_),
    .B(_0332_),
    .C(_0333_),
    .Y(_0342_));
 sg13g2_and4_1 _2725_ (.A(_0318_),
    .B(_0325_),
    .C(_0341_),
    .D(_0342_),
    .X(_0343_));
 sg13g2_a21oi_1 _2726_ (.A1(_0312_),
    .A2(_0343_),
    .Y(_0344_),
    .B1(_0338_));
 sg13g2_a22oi_1 _2727_ (.Y(_0345_),
    .B1(_0337_),
    .B2(_0344_),
    .A2(_0307_),
    .A1(net619));
 sg13g2_xor2_1 _2728_ (.B(_1441_),
    .A(net583),
    .X(_0346_));
 sg13g2_inv_1 _2729_ (.Y(_0347_),
    .A(_0346_));
 sg13g2_nand2_1 _2730_ (.Y(_0348_),
    .A(net657),
    .B(_1443_));
 sg13g2_o21ai_1 _2731_ (.B1(_0348_),
    .Y(_0349_),
    .A1(_1440_),
    .A2(_0209_));
 sg13g2_xnor2_1 _2732_ (.Y(_0350_),
    .A(_0639_),
    .B(_0346_));
 sg13g2_a22oi_1 _2733_ (.Y(_0351_),
    .B1(_0349_),
    .B2(_0350_),
    .A2(_0347_),
    .A1(net648));
 sg13g2_xor2_1 _2734_ (.B(_0280_),
    .A(net577),
    .X(_0352_));
 sg13g2_xnor2_1 _2735_ (.Y(_0353_),
    .A(_0629_),
    .B(_0352_));
 sg13g2_a22oi_1 _2736_ (.Y(_0354_),
    .B1(_0352_),
    .B2(net641),
    .A2(_0275_),
    .A1(net633));
 sg13g2_o21ai_1 _2737_ (.B1(_0354_),
    .Y(_0355_),
    .A1(_0351_),
    .A2(_0353_));
 sg13g2_nand2_1 _2738_ (.Y(_0356_),
    .A(net569),
    .B(_0268_));
 sg13g2_xnor2_1 _2739_ (.Y(_0357_),
    .A(_0834_),
    .B(_0356_));
 sg13g2_nand3_1 _2740_ (.B(_0355_),
    .C(_0357_),
    .A(_0278_),
    .Y(_0358_));
 sg13g2_xnor2_1 _2741_ (.Y(_0359_),
    .A(net565),
    .B(_0356_));
 sg13g2_and3_1 _2742_ (.X(_0360_),
    .A(_0458_),
    .B(_0491_),
    .C(_0268_));
 sg13g2_xnor2_1 _2743_ (.Y(_0361_),
    .A(net560),
    .B(_0360_));
 sg13g2_inv_1 _2744_ (.Y(_0362_),
    .A(_0361_));
 sg13g2_a22oi_1 _2745_ (.Y(_0363_),
    .B1(_0362_),
    .B2(net617),
    .A2(_0359_),
    .A1(net627));
 sg13g2_or2_1 _2746_ (.X(_0364_),
    .B(_0360_),
    .A(_0028_));
 sg13g2_a22oi_1 _2747_ (.Y(_0365_),
    .B1(_0363_),
    .B2(_0358_),
    .A2(_0361_),
    .A1(_0513_));
 sg13g2_a221oi_1 _2748_ (.B2(_0365_),
    .C1(_0345_),
    .B1(_0364_),
    .A1(net561),
    .Y(_0366_),
    .A2(_0306_));
 sg13g2_o21ai_1 _2749_ (.B1(_0366_),
    .Y(_0367_),
    .A1(_0238_),
    .A2(_0301_));
 sg13g2_nor2_1 _2750_ (.A(net651),
    .B(_1202_),
    .Y(_0368_));
 sg13g2_xor2_1 _2751_ (.B(_1202_),
    .A(net651),
    .X(_0369_));
 sg13g2_xnor2_1 _2752_ (.Y(_0370_),
    .A(net651),
    .B(_1202_));
 sg13g2_nor2_1 _2753_ (.A(net669),
    .B(net534),
    .Y(_0371_));
 sg13g2_xnor2_1 _2754_ (.Y(_0372_),
    .A(net658),
    .B(_1191_));
 sg13g2_nor2b_1 _2755_ (.A(_0371_),
    .B_N(_0372_),
    .Y(_0373_));
 sg13g2_nor3_1 _2756_ (.A(net658),
    .B(net534),
    .C(_1147_),
    .Y(_0374_));
 sg13g2_o21ai_1 _2757_ (.B1(_0369_),
    .Y(_0375_),
    .A1(_0373_),
    .A2(_0374_));
 sg13g2_nand2b_1 _2758_ (.Y(_0376_),
    .B(_0370_),
    .A_N(_0372_));
 sg13g2_nor2_1 _2759_ (.A(_1175_),
    .B(_1326_),
    .Y(_0377_));
 sg13g2_nor2_1 _2760_ (.A(_0546_),
    .B(net670),
    .Y(_0378_));
 sg13g2_nand2b_1 _2761_ (.Y(_0379_),
    .B(net680),
    .A_N(net669));
 sg13g2_a21oi_1 _2762_ (.A1(_0403_),
    .A2(_0379_),
    .Y(_0380_),
    .B1(net658));
 sg13g2_o21ai_1 _2763_ (.B1(_0546_),
    .Y(_0381_),
    .A1(net669),
    .A2(net658));
 sg13g2_nand3b_1 _2764_ (.B(_0381_),
    .C(_0369_),
    .Y(_0382_),
    .A_N(_0380_));
 sg13g2_o21ai_1 _2765_ (.B1(_0382_),
    .Y(_0383_),
    .A1(_0376_),
    .A2(_0377_));
 sg13g2_nor2_1 _2766_ (.A(net607),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_xnor2_1 _2767_ (.Y(_0385_),
    .A(net607),
    .B(_0383_));
 sg13g2_o21ai_1 _2768_ (.B1(_1221_),
    .Y(_0386_),
    .A1(_0021_),
    .A2(_1326_));
 sg13g2_nor2_1 _2769_ (.A(_0656_),
    .B(net658),
    .Y(_0387_));
 sg13g2_a22oi_1 _2770_ (.Y(_0388_),
    .B1(_0387_),
    .B2(_1123_),
    .A2(_0386_),
    .A1(_0372_));
 sg13g2_a21oi_1 _2771_ (.A1(_1174_),
    .A2(_1222_),
    .Y(_0389_),
    .B1(_0376_));
 sg13g2_a21oi_2 _2772_ (.B1(_0389_),
    .Y(_0390_),
    .A2(_0388_),
    .A1(_0369_));
 sg13g2_o21ai_1 _2773_ (.B1(_0385_),
    .Y(_0391_),
    .A1(_0392_),
    .A2(_0390_));
 sg13g2_o21ai_1 _2774_ (.B1(_0391_),
    .Y(_0393_),
    .A1(net605),
    .A2(_0383_));
 sg13g2_xnor2_1 _2775_ (.Y(_0394_),
    .A(net554),
    .B(_0375_));
 sg13g2_a22oi_1 _2776_ (.Y(_0395_),
    .B1(_0393_),
    .B2(_0394_),
    .A2(_0375_),
    .A1(_0675_));
 sg13g2_o21ai_1 _2777_ (.B1(_0379_),
    .Y(_0396_),
    .A1(_0656_),
    .A2(net534));
 sg13g2_o21ai_1 _2778_ (.B1(_0369_),
    .Y(_0397_),
    .A1(net658),
    .A2(_0396_));
 sg13g2_nor2_2 _2779_ (.A(_0373_),
    .B(_0397_),
    .Y(_0398_));
 sg13g2_xnor2_1 _2780_ (.Y(_0399_),
    .A(net556),
    .B(_0390_));
 sg13g2_and2_1 _2781_ (.A(_0385_),
    .B(_0394_),
    .X(_0400_));
 sg13g2_a221oi_1 _2782_ (.B2(_0400_),
    .C1(_0395_),
    .B1(_0399_),
    .A1(net594),
    .Y(_0401_),
    .A2(_0398_));
 sg13g2_nor3_2 _2783_ (.A(net658),
    .B(_1327_),
    .C(_0370_),
    .Y(_0402_));
 sg13g2_nand2b_1 _2784_ (.Y(_0404_),
    .B(_1442_),
    .A_N(_0402_));
 sg13g2_o21ai_1 _2785_ (.B1(_0404_),
    .Y(_0405_),
    .A1(net594),
    .A2(_0398_));
 sg13g2_nor2_1 _2786_ (.A(net543),
    .B(_1202_),
    .Y(_0406_));
 sg13g2_nor2_1 _2787_ (.A(_0713_),
    .B(_1202_),
    .Y(_0407_));
 sg13g2_nor2_1 _2788_ (.A(_0715_),
    .B(_1202_),
    .Y(_0408_));
 sg13g2_nor3_1 _2789_ (.A(net620),
    .B(_0715_),
    .C(_1202_),
    .Y(_0409_));
 sg13g2_xnor2_1 _2790_ (.Y(_0410_),
    .A(_0513_),
    .B(_0409_));
 sg13g2_xnor2_1 _2791_ (.Y(_0411_),
    .A(net625),
    .B(_0408_));
 sg13g2_xnor2_1 _2792_ (.Y(_0412_),
    .A(net643),
    .B(_0368_));
 sg13g2_xnor2_1 _2793_ (.Y(_0413_),
    .A(net640),
    .B(_0407_));
 sg13g2_nor2b_1 _2794_ (.A(_0412_),
    .B_N(_0413_),
    .Y(_0415_));
 sg13g2_nor3_1 _2795_ (.A(net634),
    .B(_0713_),
    .C(_1202_),
    .Y(_0416_));
 sg13g2_xnor2_1 _2796_ (.Y(_0417_),
    .A(net631),
    .B(_0416_));
 sg13g2_nand4_1 _2797_ (.B(_0411_),
    .C(_0415_),
    .A(_0410_),
    .Y(_0418_),
    .D(_0417_));
 sg13g2_a21oi_1 _2798_ (.A1(_1443_),
    .A2(_0402_),
    .Y(_0419_),
    .B1(_0418_));
 sg13g2_o21ai_1 _2799_ (.B1(_0419_),
    .Y(_0420_),
    .A1(_0401_),
    .A2(_0405_));
 sg13g2_nor2_1 _2800_ (.A(_1173_),
    .B(_1223_),
    .Y(_0421_));
 sg13g2_nand2_1 _2801_ (.Y(_0422_),
    .A(net543),
    .B(_0823_));
 sg13g2_xnor2_1 _2802_ (.Y(_0423_),
    .A(net654),
    .B(_0823_));
 sg13g2_xnor2_1 _2803_ (.Y(_0424_),
    .A(net543),
    .B(_0823_));
 sg13g2_nand3_1 _2804_ (.B(_1207_),
    .C(_0423_),
    .A(_1127_),
    .Y(_0426_));
 sg13g2_nor2_1 _2805_ (.A(_0421_),
    .B(_0426_),
    .Y(_0427_));
 sg13g2_nor2_1 _2806_ (.A(_1223_),
    .B(_0424_),
    .Y(_0428_));
 sg13g2_o21ai_1 _2807_ (.B1(_1443_),
    .Y(_0429_),
    .A1(_1223_),
    .A2(_0424_));
 sg13g2_nand2_1 _2808_ (.Y(_0430_),
    .A(_1442_),
    .B(_0428_));
 sg13g2_a22oi_1 _2809_ (.Y(_0431_),
    .B1(_0429_),
    .B2(_0430_),
    .A2(_0427_),
    .A1(net594));
 sg13g2_or2_1 _2810_ (.X(_0432_),
    .B(_0427_),
    .A(net594));
 sg13g2_o21ai_1 _2811_ (.B1(net661),
    .Y(_0433_),
    .A1(_0656_),
    .A2(_0819_));
 sg13g2_o21ai_1 _2812_ (.B1(_1190_),
    .Y(_0434_),
    .A1(net686),
    .A2(_0021_));
 sg13g2_a221oi_1 _2813_ (.B2(_0434_),
    .C1(_1206_),
    .B1(_0433_),
    .A1(net661),
    .Y(_0435_),
    .A2(_0656_));
 sg13g2_nand2b_2 _2814_ (.Y(_0437_),
    .B(_0423_),
    .A_N(_0435_));
 sg13g2_xnor2_1 _2815_ (.Y(_0438_),
    .A(net554),
    .B(_0437_));
 sg13g2_nand3_1 _2816_ (.B(_0432_),
    .C(_0438_),
    .A(_0431_),
    .Y(_0439_));
 sg13g2_a21oi_1 _2817_ (.A1(net551),
    .A2(_1190_),
    .Y(_0440_),
    .B1(net680));
 sg13g2_nor3_1 _2818_ (.A(_0546_),
    .B(_0656_),
    .C(_1162_),
    .Y(_0441_));
 sg13g2_o21ai_1 _2819_ (.B1(_0423_),
    .Y(_0442_),
    .A1(_0440_),
    .A2(_0441_));
 sg13g2_nand4_1 _2820_ (.B(_1205_),
    .C(_0379_),
    .A(net551),
    .Y(_0443_),
    .D(_0424_));
 sg13g2_and2_2 _2821_ (.A(_0442_),
    .B(_0443_),
    .X(_0444_));
 sg13g2_xnor2_1 _2822_ (.Y(_0445_),
    .A(net555),
    .B(_0444_));
 sg13g2_nand4_1 _2823_ (.B(_0396_),
    .C(_0424_),
    .A(_1207_),
    .Y(_0446_),
    .D(_0433_));
 sg13g2_a221oi_1 _2824_ (.B2(_1207_),
    .C1(_0378_),
    .B1(_0433_),
    .A1(\hx0[0] ),
    .Y(_0448_),
    .A2(_1222_));
 sg13g2_nand2_1 _2825_ (.Y(_0449_),
    .A(_0656_),
    .B(_1123_));
 sg13g2_o21ai_1 _2826_ (.B1(_0423_),
    .Y(_0450_),
    .A1(net661),
    .A2(_0449_));
 sg13g2_o21ai_1 _2827_ (.B1(_0446_),
    .Y(_0451_),
    .A1(_0448_),
    .A2(_0450_));
 sg13g2_nand2_1 _2828_ (.Y(_0452_),
    .A(net610),
    .B(_0451_));
 sg13g2_a22oi_1 _2829_ (.Y(_0453_),
    .B1(_0445_),
    .B2(_0452_),
    .A2(_0444_),
    .A1(_0680_));
 sg13g2_nor2_1 _2830_ (.A(_1443_),
    .B(_0428_),
    .Y(_0454_));
 sg13g2_nand2_1 _2831_ (.Y(_0455_),
    .A(_0675_),
    .B(_0437_));
 sg13g2_nand2_1 _2832_ (.Y(_0456_),
    .A(_0432_),
    .B(_0455_));
 sg13g2_a21oi_1 _2833_ (.A1(_0431_),
    .A2(_0456_),
    .Y(_0457_),
    .B1(_0454_));
 sg13g2_o21ai_1 _2834_ (.B1(_0457_),
    .Y(_0459_),
    .A1(_0439_),
    .A2(_0453_));
 sg13g2_nand2_1 _2835_ (.Y(_0460_),
    .A(net612),
    .B(_0451_));
 sg13g2_xnor2_1 _2836_ (.Y(_0461_),
    .A(net612),
    .B(_0451_));
 sg13g2_nand3b_1 _2837_ (.B(_0445_),
    .C(_0461_),
    .Y(_0462_),
    .A_N(_0439_));
 sg13g2_a22oi_1 _2838_ (.Y(_0463_),
    .B1(_0422_),
    .B2(net648),
    .A2(net539),
    .A1(_0823_));
 sg13g2_xnor2_1 _2839_ (.Y(_0464_),
    .A(net624),
    .B(_0782_));
 sg13g2_nor4_2 _2840_ (.A(_1514_),
    .B(_0140_),
    .C(_0463_),
    .Y(_0465_),
    .D(_0464_));
 sg13g2_nand2_1 _2841_ (.Y(_0466_),
    .A(_0136_),
    .B(_0465_));
 sg13g2_nand4_1 _2842_ (.B(_0459_),
    .C(_0462_),
    .A(_0136_),
    .Y(_0467_),
    .D(_0465_));
 sg13g2_o21ai_1 _2843_ (.B1(_0614_),
    .Y(_0468_),
    .A1(net579),
    .A2(_0267_));
 sg13g2_xnor2_1 _2844_ (.Y(_0470_),
    .A(_0622_),
    .B(_0468_));
 sg13g2_o21ai_1 _2845_ (.B1(_0699_),
    .Y(_0471_),
    .A1(net579),
    .A2(_0267_));
 sg13g2_xnor2_1 _2846_ (.Y(_0472_),
    .A(_0028_),
    .B(_0471_));
 sg13g2_nor2b_1 _2847_ (.A(_0281_),
    .B_N(_0283_),
    .Y(_0473_));
 sg13g2_nand4_1 _2848_ (.B(_0470_),
    .C(_0472_),
    .A(_1455_),
    .Y(_0474_),
    .D(_0473_));
 sg13g2_a21oi_1 _2849_ (.A1(_0420_),
    .A2(_0467_),
    .Y(_0475_),
    .B1(_0474_));
 sg13g2_o21ai_1 _2850_ (.B1(net541),
    .Y(_0476_),
    .A1(_0421_),
    .A2(_0426_));
 sg13g2_nor2_1 _2851_ (.A(net600),
    .B(_0437_),
    .Y(_0477_));
 sg13g2_nand2b_1 _2852_ (.Y(_0478_),
    .B(_0675_),
    .A_N(_0437_));
 sg13g2_xnor2_1 _2853_ (.Y(_0479_),
    .A(_0680_),
    .B(_0444_));
 sg13g2_a22oi_1 _2854_ (.Y(_0481_),
    .B1(_0460_),
    .B2(_0479_),
    .A2(_0444_),
    .A1(net555));
 sg13g2_o21ai_1 _2855_ (.B1(_0476_),
    .Y(_0482_),
    .A1(_0477_),
    .A2(_0481_));
 sg13g2_xnor2_1 _2856_ (.Y(_0483_),
    .A(net610),
    .B(_0451_));
 sg13g2_xnor2_1 _2857_ (.Y(_0484_),
    .A(net594),
    .B(_0427_));
 sg13g2_nand4_1 _2858_ (.B(_0479_),
    .C(_0483_),
    .A(_0478_),
    .Y(_0485_),
    .D(_0484_));
 sg13g2_a22oi_1 _2859_ (.Y(_0486_),
    .B1(_0482_),
    .B2(_0485_),
    .A2(_0437_),
    .A1(net600));
 sg13g2_nor2b_1 _2860_ (.A(_0484_),
    .B_N(_0476_),
    .Y(_0487_));
 sg13g2_o21ai_1 _2861_ (.B1(_0429_),
    .Y(_0488_),
    .A1(_0486_),
    .A2(_0487_));
 sg13g2_nor2b_1 _2862_ (.A(_0466_),
    .B_N(_0430_),
    .Y(_0489_));
 sg13g2_xnor2_1 _2863_ (.Y(_0490_),
    .A(_1443_),
    .B(_0402_));
 sg13g2_nor2_1 _2864_ (.A(net592),
    .B(_0398_),
    .Y(_0492_));
 sg13g2_xnor2_1 _2865_ (.Y(_0493_),
    .A(net594),
    .B(_0398_));
 sg13g2_o21ai_1 _2866_ (.B1(_0493_),
    .Y(_0494_),
    .A1(net600),
    .A2(_0375_));
 sg13g2_xnor2_1 _2867_ (.Y(_0495_),
    .A(net605),
    .B(_0383_));
 sg13g2_o21ai_1 _2868_ (.B1(_0495_),
    .Y(_0496_),
    .A1(net556),
    .A2(_0390_));
 sg13g2_a21oi_1 _2869_ (.A1(net600),
    .A2(_0375_),
    .Y(_0497_),
    .B1(_0384_));
 sg13g2_a21oi_1 _2870_ (.A1(_0496_),
    .A2(_0497_),
    .Y(_0498_),
    .B1(_0494_));
 sg13g2_o21ai_1 _2871_ (.B1(_0490_),
    .Y(_0499_),
    .A1(_0492_),
    .A2(_0498_));
 sg13g2_o21ai_1 _2872_ (.B1(_0499_),
    .Y(_0500_),
    .A1(_1442_),
    .A2(_0402_));
 sg13g2_a21oi_1 _2873_ (.A1(net600),
    .A2(_0375_),
    .Y(_0501_),
    .B1(_0494_));
 sg13g2_xnor2_1 _2874_ (.Y(_0503_),
    .A(_0392_),
    .B(_0390_));
 sg13g2_nand4_1 _2875_ (.B(_0495_),
    .C(_0501_),
    .A(_0490_),
    .Y(_0504_),
    .D(_0503_));
 sg13g2_nor2b_1 _2876_ (.A(_0418_),
    .B_N(_0504_),
    .Y(_0505_));
 sg13g2_a22oi_1 _2877_ (.Y(_0506_),
    .B1(_0500_),
    .B2(_0505_),
    .A2(_0489_),
    .A1(_0488_));
 sg13g2_nand2_1 _2878_ (.Y(_0507_),
    .A(_0447_),
    .B(_0267_));
 sg13g2_nand2_2 _2879_ (.Y(_0508_),
    .A(net577),
    .B(_0507_));
 sg13g2_nand2_1 _2880_ (.Y(_0509_),
    .A(_0699_),
    .B(_0508_));
 sg13g2_xnor2_1 _2881_ (.Y(_0510_),
    .A(_0028_),
    .B(_0509_));
 sg13g2_nand2_1 _2882_ (.Y(_0511_),
    .A(net573),
    .B(_0508_));
 sg13g2_xnor2_1 _2883_ (.Y(_0512_),
    .A(_0622_),
    .B(_0511_));
 sg13g2_o21ai_1 _2884_ (.B1(_0347_),
    .Y(_0514_),
    .A1(_0030_),
    .A2(_0508_));
 sg13g2_a21oi_1 _2885_ (.A1(net569),
    .A2(_0508_),
    .Y(_0515_),
    .B1(_0352_));
 sg13g2_nand2b_1 _2886_ (.Y(_0516_),
    .B(_0515_),
    .A_N(_0514_));
 sg13g2_nor4_1 _2887_ (.A(_0506_),
    .B(_0510_),
    .C(_0512_),
    .D(_0516_),
    .Y(_0517_));
 sg13g2_or2_1 _2888_ (.X(_0518_),
    .B(_0517_),
    .A(_0475_));
 sg13g2_mux2_1 _2889_ (.A0(_0019_),
    .A1(net8),
    .S(net529),
    .X(_0519_));
 sg13g2_nand2b_1 _2890_ (.Y(_0520_),
    .B(net529),
    .A_N(net6));
 sg13g2_o21ai_1 _2891_ (.B1(_0520_),
    .Y(_0521_),
    .A1(net529),
    .A2(_0017_));
 sg13g2_nand2b_1 _2892_ (.Y(_0522_),
    .B(net528),
    .A_N(net5));
 sg13g2_o21ai_1 _2893_ (.B1(_0522_),
    .Y(_0523_),
    .A1(net528),
    .A2(_0016_));
 sg13g2_nand2_1 _2894_ (.Y(_0525_),
    .A(_0714_),
    .B(_0802_));
 sg13g2_nand2_2 _2895_ (.Y(_0526_),
    .A(_0715_),
    .B(_0802_));
 sg13g2_nor4_1 _2896_ (.A(_0090_),
    .B(_0226_),
    .C(_0523_),
    .D(_0526_),
    .Y(_0527_));
 sg13g2_nor3_1 _2897_ (.A(_0299_),
    .B(_0521_),
    .C(_0526_),
    .Y(_0528_));
 sg13g2_and3_1 _2898_ (.X(_0529_),
    .A(_1469_),
    .B(_0294_),
    .C(_0528_));
 sg13g2_o21ai_1 _2899_ (.B1(_0525_),
    .Y(_0530_),
    .A1(_0527_),
    .A2(_0529_));
 sg13g2_nor3_1 _2900_ (.A(_0226_),
    .B(_0228_),
    .C(_0235_),
    .Y(_0531_));
 sg13g2_a221oi_1 _2901_ (.B2(_0028_),
    .C1(_0160_),
    .B1(_0232_),
    .A1(net589),
    .Y(_0532_),
    .A2(_0231_));
 sg13g2_a22oi_1 _2902_ (.Y(_0533_),
    .B1(_0531_),
    .B2(_0532_),
    .A2(_0519_),
    .A1(_0518_));
 sg13g2_nand4_1 _2903_ (.B(_0367_),
    .C(_0530_),
    .A(_0165_),
    .Y(_0534_),
    .D(_0533_));
 sg13g2_xnor2_1 _2904_ (.Y(_0536_),
    .A(net571),
    .B(net570));
 sg13g2_xnor2_1 _2905_ (.Y(_0537_),
    .A(net566),
    .B(_1070_));
 sg13g2_a221oi_1 _2906_ (.B2(net536),
    .C1(_0537_),
    .B1(_0536_),
    .A1(net571),
    .Y(_0538_),
    .A2(_0975_));
 sg13g2_xnor2_1 _2907_ (.Y(_0539_),
    .A(net562),
    .B(_1073_));
 sg13g2_a21oi_2 _2908_ (.B1(_1074_),
    .Y(_0540_),
    .A2(_0539_),
    .A1(_0538_));
 sg13g2_nand2_1 _2909_ (.Y(_0541_),
    .A(net610),
    .B(net595));
 sg13g2_a22oi_1 _2910_ (.Y(_0542_),
    .B1(_0541_),
    .B2(_0704_),
    .A2(_0233_),
    .A1(net541));
 sg13g2_nor3_1 _2911_ (.A(net610),
    .B(net552),
    .C(net591),
    .Y(_0543_));
 sg13g2_a22oi_1 _2912_ (.Y(_0544_),
    .B1(net595),
    .B2(_0543_),
    .A2(net555),
    .A1(net612));
 sg13g2_o21ai_1 _2913_ (.B1(net535),
    .Y(_0545_),
    .A1(_0542_),
    .A2(_0544_));
 sg13g2_a21oi_1 _2914_ (.A1(net585),
    .A2(net593),
    .Y(_0547_),
    .B1(net555));
 sg13g2_nor2_1 _2915_ (.A(_0928_),
    .B(_0940_),
    .Y(_0548_));
 sg13g2_nor3_1 _2916_ (.A(_1089_),
    .B(_0547_),
    .C(_0548_),
    .Y(_0549_));
 sg13g2_o21ai_1 _2917_ (.B1(_0818_),
    .Y(_0550_),
    .A1(net611),
    .A2(_0549_));
 sg13g2_a21oi_1 _2918_ (.A1(_0938_),
    .A2(_0233_),
    .Y(_0551_),
    .B1(_0543_));
 sg13g2_nand2b_1 _2919_ (.Y(_0552_),
    .B(net602),
    .A_N(net595));
 sg13g2_nand3_1 _2920_ (.B(_0930_),
    .C(_0552_),
    .A(_0928_),
    .Y(_0553_));
 sg13g2_a21oi_1 _2921_ (.A1(\hy0[0] ),
    .A2(net536),
    .Y(_0554_),
    .B1(_1176_));
 sg13g2_a22oi_1 _2922_ (.Y(_0555_),
    .B1(_0553_),
    .B2(_0554_),
    .A2(_0551_),
    .A1(_1173_));
 sg13g2_and4_1 _2923_ (.A(_0985_),
    .B(_0545_),
    .C(_0550_),
    .D(_0555_),
    .X(_0556_));
 sg13g2_and2_1 _2924_ (.A(_1076_),
    .B(_0556_),
    .X(_0558_));
 sg13g2_nand2_1 _2925_ (.Y(_0559_),
    .A(_0458_),
    .B(_0927_));
 sg13g2_a221oi_1 _2926_ (.B2(_0540_),
    .C1(_0558_),
    .B1(_1077_),
    .A1(_0458_),
    .Y(_0560_),
    .A2(_0927_));
 sg13g2_a22oi_1 _2927_ (.Y(_0561_),
    .B1(_1175_),
    .B2(_0080_),
    .A2(_1173_),
    .A1(_0079_));
 sg13g2_a22oi_1 _2928_ (.Y(_0562_),
    .B1(net535),
    .B2(_0081_),
    .A2(net540),
    .A1(_0078_));
 sg13g2_a21oi_1 _2929_ (.A1(_0561_),
    .A2(_0562_),
    .Y(_0563_),
    .B1(_0559_));
 sg13g2_xor2_1 _2930_ (.B(net638),
    .A(net581),
    .X(_0564_));
 sg13g2_inv_1 _2931_ (.Y(_0565_),
    .A(_0564_));
 sg13g2_nand4_1 _2932_ (.B(_0828_),
    .C(_0931_),
    .A(_0704_),
    .Y(_0566_),
    .D(_0564_));
 sg13g2_nor3_1 _2933_ (.A(_0824_),
    .B(_0540_),
    .C(_0566_),
    .Y(_0567_));
 sg13g2_nand4_1 _2934_ (.B(_0823_),
    .C(_0828_),
    .A(_0704_),
    .Y(_0569_),
    .D(_0931_));
 sg13g2_nor3_1 _2935_ (.A(_0540_),
    .B(_0565_),
    .C(_0569_),
    .Y(_0570_));
 sg13g2_nor4_1 _2936_ (.A(_0534_),
    .B(_0560_),
    .C(_0563_),
    .D(_0567_),
    .Y(_0571_));
 sg13g2_a21oi_2 _2937_ (.B1(_0720_),
    .Y(uo_out[6]),
    .A2(_0571_),
    .A1(_1395_));
 sg13g2_nor2_1 _2938_ (.A(_1067_),
    .B(_0534_),
    .Y(_0572_));
 sg13g2_o21ai_1 _2939_ (.B1(_1394_),
    .Y(_0573_),
    .A1(_0558_),
    .A2(_0567_));
 sg13g2_a21oi_2 _2940_ (.B1(_0720_),
    .Y(uo_out[2]),
    .A2(_0573_),
    .A1(_0572_));
 sg13g2_a21oi_1 _2941_ (.A1(net556),
    .A2(net608),
    .Y(_0574_),
    .B1(_0931_));
 sg13g2_nor2_1 _2942_ (.A(_0234_),
    .B(_0574_),
    .Y(_0575_));
 sg13g2_a21oi_1 _2943_ (.A1(net610),
    .A2(_1090_),
    .Y(_0576_),
    .B1(_0575_));
 sg13g2_nor2_1 _2944_ (.A(net595),
    .B(_0480_),
    .Y(_0578_));
 sg13g2_a22oi_1 _2945_ (.Y(_0579_),
    .B1(_0578_),
    .B2(net614),
    .A2(_1443_),
    .A1(_0938_));
 sg13g2_nor3_1 _2946_ (.A(_0819_),
    .B(_0206_),
    .C(_0579_),
    .Y(_0580_));
 sg13g2_nand2_1 _2947_ (.Y(_0581_),
    .A(net542),
    .B(_1175_));
 sg13g2_nor4_1 _2948_ (.A(net556),
    .B(net609),
    .C(_1089_),
    .D(_0581_),
    .Y(_0582_));
 sg13g2_and2_1 _2949_ (.A(net595),
    .B(_0233_),
    .X(_0583_));
 sg13g2_a21oi_1 _2950_ (.A1(_0704_),
    .A2(_0940_),
    .Y(_0584_),
    .B1(_0583_));
 sg13g2_nor2b_1 _2951_ (.A(_0584_),
    .B_N(_0930_),
    .Y(_0585_));
 sg13g2_nor3_1 _2952_ (.A(_0392_),
    .B(_0704_),
    .C(_0583_),
    .Y(_0586_));
 sg13g2_o21ai_1 _2953_ (.B1(net535),
    .Y(_0587_),
    .A1(_0585_),
    .A2(_0586_));
 sg13g2_o21ai_1 _2954_ (.B1(_0587_),
    .Y(_0589_),
    .A1(_1174_),
    .A2(_0576_));
 sg13g2_nor4_1 _2955_ (.A(_0985_),
    .B(_0580_),
    .C(_0582_),
    .D(_0589_),
    .Y(_0590_));
 sg13g2_or2_1 _2956_ (.X(_0591_),
    .B(_0590_),
    .A(_0556_));
 sg13g2_a21o_1 _2957_ (.A2(_0591_),
    .A1(_1076_),
    .B1(_1394_),
    .X(_0592_));
 sg13g2_a21oi_2 _2958_ (.B1(_0720_),
    .Y(uo_out[5]),
    .A2(_0592_),
    .A1(_0572_));
 sg13g2_nor2_1 _2959_ (.A(_1076_),
    .B(_0591_),
    .Y(_0593_));
 sg13g2_mux2_1 _2960_ (.A0(_0570_),
    .A1(_0593_),
    .S(_1393_),
    .X(_0594_));
 sg13g2_a21oi_1 _2961_ (.A1(_1068_),
    .A2(_0594_),
    .Y(_0595_),
    .B1(_0534_));
 sg13g2_nor2_2 _2962_ (.A(_0720_),
    .B(_0595_),
    .Y(uo_out[1]));
 sg13g2_or2_1 _2963_ (.X(_0596_),
    .B(_0534_),
    .A(_0720_));
 sg13g2_nor2_2 _2964_ (.A(_1395_),
    .B(_0596_),
    .Y(uo_out[4]));
 sg13g2_nand2b_1 _2965_ (.Y(_0598_),
    .B(_0558_),
    .A_N(_0567_));
 sg13g2_a21oi_2 _2966_ (.B1(_0596_),
    .Y(uo_out[0]),
    .A2(_0598_),
    .A1(_1395_));
 sg13g2_nand3_1 _2967_ (.B(net533),
    .C(_1051_),
    .A(net532),
    .Y(_0599_));
 sg13g2_nor2_1 _2968_ (.A(_0697_),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_nand2_1 _2969_ (.Y(_0601_),
    .A(net531),
    .B(_0600_));
 sg13g2_nand2_1 _2970_ (.Y(_0602_),
    .A(_0022_),
    .B(_0601_));
 sg13g2_or2_1 _2971_ (.X(_0603_),
    .B(_0601_),
    .A(_0022_));
 sg13g2_nand3_1 _2972_ (.B(_0602_),
    .C(_0603_),
    .A(net690),
    .Y(_0604_));
 sg13g2_inv_2 _2973_ (.Y(_0052_),
    .A(_0604_));
 sg13g2_nand4_1 _2974_ (.B(net531),
    .C(\counter[7] ),
    .A(\counter[6] ),
    .Y(_0606_),
    .D(_0600_));
 sg13g2_nand2_1 _2975_ (.Y(_0607_),
    .A(_0034_),
    .B(_0606_));
 sg13g2_nor2_1 _2976_ (.A(_0034_),
    .B(_0606_),
    .Y(_0608_));
 sg13g2_nand3b_1 _2977_ (.B(net691),
    .C(_0607_),
    .Y(_0609_),
    .A_N(_0608_));
 sg13g2_inv_1 _2978_ (.Y(_0054_),
    .A(_0609_));
 sg13g2_xnor2_1 _2979_ (.Y(_0610_),
    .A(\counter[7] ),
    .B(_0603_));
 sg13g2_nand2_2 _2980_ (.Y(_0611_),
    .A(net691),
    .B(_0610_));
 sg13g2_inv_1 _2981_ (.Y(_0053_),
    .A(_0611_));
 sg13g2_nand2_1 _2982_ (.Y(_0612_),
    .A(_0609_),
    .B(_0611_));
 sg13g2_nand3_1 _2983_ (.B(_0609_),
    .C(_0611_),
    .A(_0052_),
    .Y(_0613_));
 sg13g2_o21ai_1 _2984_ (.B1(net691),
    .Y(_0615_),
    .A1(\counter[9] ),
    .A2(_0608_));
 sg13g2_a21oi_2 _2985_ (.B1(_0615_),
    .Y(_0055_),
    .A2(_0608_),
    .A1(\counter[9] ));
 sg13g2_a21oi_1 _2986_ (.A1(_0052_),
    .A2(_0611_),
    .Y(_0616_),
    .B1(_0055_));
 sg13g2_inv_1 _2987_ (.Y(_0617_),
    .A(_0616_));
 sg13g2_nand2_1 _2988_ (.Y(_0000_),
    .A(_0613_),
    .B(_0617_));
 sg13g2_nor2_1 _2989_ (.A(_0052_),
    .B(_0611_),
    .Y(_0618_));
 sg13g2_nor2_1 _2990_ (.A(_0054_),
    .B(_0618_),
    .Y(_0619_));
 sg13g2_nor2_1 _2991_ (.A(_0055_),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_o21ai_1 _2992_ (.B1(_0620_),
    .Y(_0621_),
    .A1(_0052_),
    .A2(_0053_));
 sg13g2_nand2_1 _2993_ (.Y(_0001_),
    .A(_0612_),
    .B(_0621_));
 sg13g2_nand2_1 _2994_ (.Y(_0623_),
    .A(_0052_),
    .B(_0053_));
 sg13g2_nor2_1 _2995_ (.A(_0609_),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_a21oi_1 _2996_ (.A1(_0612_),
    .A2(_0055_),
    .Y(_0002_),
    .B1(_0624_));
 sg13g2_a22oi_1 _2997_ (.Y(_0003_),
    .B1(_0612_),
    .B2(_0617_),
    .A2(_0609_),
    .A1(_0604_));
 sg13g2_o21ai_1 _2998_ (.B1(_0613_),
    .Y(_0004_),
    .A1(_0055_),
    .A2(_0623_));
 sg13g2_a22oi_1 _2999_ (.Y(_0005_),
    .B1(_0620_),
    .B2(_0610_),
    .A2(_0055_),
    .A1(_0613_));
 sg13g2_nand4_1 _3000_ (.B(net624),
    .C(_0782_),
    .A(net619),
    .Y(_0625_),
    .D(_0406_));
 sg13g2_and2_2 _3001_ (.A(net691),
    .B(_0625_),
    .X(_0626_));
 sg13g2_nand2_1 _3002_ (.Y(_0627_),
    .A(net691),
    .B(_0625_));
 sg13g2_nand2b_1 _3003_ (.Y(_0628_),
    .B(_0975_),
    .A_N(net525));
 sg13g2_o21ai_1 _3004_ (.B1(net578),
    .Y(_0630_),
    .A1(net536),
    .A2(net525));
 sg13g2_nor2_1 _3005_ (.A(_0940_),
    .B(_0971_),
    .Y(_0631_));
 sg13g2_nand4_1 _3006_ (.B(_0930_),
    .C(_0932_),
    .A(net562),
    .Y(_0632_),
    .D(_0631_));
 sg13g2_o21ai_1 _3007_ (.B1(net690),
    .Y(_0633_),
    .A1(net567),
    .A2(_0632_));
 sg13g2_nor2_2 _3008_ (.A(_0625_),
    .B(_0633_),
    .Y(_0634_));
 sg13g2_or2_2 _3009_ (.X(_0635_),
    .B(_0633_),
    .A(_0625_));
 sg13g2_nand3_1 _3010_ (.B(_0630_),
    .C(_0634_),
    .A(_0628_),
    .Y(_0636_));
 sg13g2_o21ai_1 _3011_ (.B1(_0636_),
    .Y(_0637_),
    .A1(net578),
    .A2(net521));
 sg13g2_a22oi_1 _3012_ (.Y(_0638_),
    .B1(_0634_),
    .B2(net610),
    .A2(net523),
    .A1(net611));
 sg13g2_inv_1 _3013_ (.Y(_0067_),
    .A(_0638_));
 sg13g2_nand2b_1 _3014_ (.Y(_0640_),
    .B(_0638_),
    .A_N(_0637_));
 sg13g2_nor2_1 _3015_ (.A(net587),
    .B(net524),
    .Y(_0641_));
 sg13g2_xnor2_1 _3016_ (.Y(_0642_),
    .A(net584),
    .B(_0641_));
 sg13g2_a22oi_1 _3017_ (.Y(_0643_),
    .B1(_0634_),
    .B2(_0642_),
    .A2(net523),
    .A1(net585));
 sg13g2_inv_1 _3018_ (.Y(_0072_),
    .A(_0643_));
 sg13g2_xor2_1 _3019_ (.B(net609),
    .A(net611),
    .X(_0644_));
 sg13g2_nand2_1 _3020_ (.Y(_0645_),
    .A(_0634_),
    .B(_0644_));
 sg13g2_o21ai_1 _3021_ (.B1(_0645_),
    .Y(_0068_),
    .A1(net555),
    .A2(net521));
 sg13g2_nand2_1 _3022_ (.Y(_0646_),
    .A(net595),
    .B(net523));
 sg13g2_xnor2_1 _3023_ (.Y(_0647_),
    .A(net593),
    .B(_0939_));
 sg13g2_o21ai_1 _3024_ (.B1(_0646_),
    .Y(_0070_),
    .A1(_0635_),
    .A2(_0647_));
 sg13g2_nand2_1 _3025_ (.Y(_0649_),
    .A(net603),
    .B(net523));
 sg13g2_o21ai_1 _3026_ (.B1(_0649_),
    .Y(_0069_),
    .A1(_0316_),
    .A2(_0635_));
 sg13g2_a21oi_1 _3027_ (.A1(_0070_),
    .A2(_0069_),
    .Y(_0650_),
    .B1(_0068_));
 sg13g2_nand2_1 _3028_ (.Y(_0651_),
    .A(net588),
    .B(net523));
 sg13g2_xnor2_1 _3029_ (.Y(_0652_),
    .A(net587),
    .B(net524));
 sg13g2_o21ai_1 _3030_ (.B1(_0651_),
    .Y(_0071_),
    .A1(_0635_),
    .A2(_0652_));
 sg13g2_or2_1 _3031_ (.X(_0653_),
    .B(_0071_),
    .A(_0067_));
 sg13g2_a21oi_1 _3032_ (.A1(_0644_),
    .A2(_0070_),
    .Y(_0654_),
    .B1(_0653_));
 sg13g2_nor2_1 _3033_ (.A(_0650_),
    .B(_0654_),
    .Y(_0655_));
 sg13g2_nor2_1 _3034_ (.A(_0072_),
    .B(_0655_),
    .Y(_0657_));
 sg13g2_nand2_1 _3035_ (.Y(_0658_),
    .A(_0067_),
    .B(_0643_));
 sg13g2_nand2b_1 _3036_ (.Y(_0659_),
    .B(_0068_),
    .A_N(_0070_));
 sg13g2_nor2b_1 _3037_ (.A(_0068_),
    .B_N(_0070_),
    .Y(_0660_));
 sg13g2_a21o_1 _3038_ (.A2(_0659_),
    .A1(_0071_),
    .B1(_0660_),
    .X(_0661_));
 sg13g2_o21ai_1 _3039_ (.B1(_0637_),
    .Y(_0662_),
    .A1(_0658_),
    .A2(_0661_));
 sg13g2_o21ai_1 _3040_ (.B1(_0662_),
    .Y(_0006_),
    .A1(_0640_),
    .A2(_0657_));
 sg13g2_or2_1 _3041_ (.X(_0663_),
    .B(_0071_),
    .A(_0068_));
 sg13g2_nor3_1 _3042_ (.A(_0637_),
    .B(_0638_),
    .C(_0643_),
    .Y(_0664_));
 sg13g2_nand2_1 _3043_ (.Y(_0665_),
    .A(_0663_),
    .B(_0664_));
 sg13g2_nor2b_1 _3044_ (.A(_0068_),
    .B_N(_0069_),
    .Y(_0667_));
 sg13g2_nor3_1 _3045_ (.A(_0653_),
    .B(_0660_),
    .C(_0667_),
    .Y(_0668_));
 sg13g2_o21ai_1 _3046_ (.B1(_0637_),
    .Y(_0669_),
    .A1(_0067_),
    .A2(_0072_));
 sg13g2_o21ai_1 _3047_ (.B1(_0665_),
    .Y(_0007_),
    .A1(_0668_),
    .A2(_0669_));
 sg13g2_o21ai_1 _3048_ (.B1(_0637_),
    .Y(_0670_),
    .A1(_0658_),
    .A2(_0663_));
 sg13g2_and2_1 _3049_ (.A(_0643_),
    .B(_0668_),
    .X(_0671_));
 sg13g2_o21ai_1 _3050_ (.B1(_0670_),
    .Y(_0008_),
    .A1(_0640_),
    .A2(_0671_));
 sg13g2_nand2_1 _3051_ (.Y(_0672_),
    .A(_0661_),
    .B(_0664_));
 sg13g2_a21oi_1 _3052_ (.A1(_0638_),
    .A2(_0071_),
    .Y(_0673_),
    .B1(_0654_));
 sg13g2_nor3_1 _3053_ (.A(_0643_),
    .B(_0655_),
    .C(_0673_),
    .Y(_0674_));
 sg13g2_o21ai_1 _3054_ (.B1(_0672_),
    .Y(_0009_),
    .A1(_0669_),
    .A2(_0674_));
 sg13g2_a21oi_1 _3055_ (.A1(_0609_),
    .A2(_0618_),
    .Y(_0045_),
    .B1(_0055_));
 sg13g2_and2_1 _3056_ (.A(net690),
    .B(_0044_),
    .X(_0046_));
 sg13g2_and2_1 _3057_ (.A(net690),
    .B(_1052_),
    .X(_0047_));
 sg13g2_o21ai_1 _3058_ (.B1(net690),
    .Y(_0676_),
    .A1(net533),
    .A2(_1051_));
 sg13g2_a21oi_1 _3059_ (.A1(net533),
    .A2(_1051_),
    .Y(_0048_),
    .B1(_0676_));
 sg13g2_nor2b_1 _3060_ (.A(_0027_),
    .B_N(_1051_),
    .Y(_0677_));
 sg13g2_o21ai_1 _3061_ (.B1(net690),
    .Y(_0678_),
    .A1(net532),
    .A2(_0677_));
 sg13g2_a21oi_1 _3062_ (.A1(net532),
    .A2(_0677_),
    .Y(_0049_),
    .B1(_0678_));
 sg13g2_o21ai_1 _3063_ (.B1(net690),
    .Y(_0679_),
    .A1(_0697_),
    .A2(_0599_));
 sg13g2_a21oi_1 _3064_ (.A1(_0697_),
    .A2(_0599_),
    .Y(_0050_),
    .B1(_0679_));
 sg13g2_nor2_1 _3065_ (.A(_0024_),
    .B(_0599_),
    .Y(_0681_));
 sg13g2_o21ai_1 _3066_ (.B1(net690),
    .Y(_0682_),
    .A1(net530),
    .A2(_0681_));
 sg13g2_a21oi_1 _3067_ (.A1(net530),
    .A2(_0681_),
    .Y(_0051_),
    .B1(_0682_));
 sg13g2_and2_1 _3068_ (.A(net70),
    .B(net523),
    .X(_0056_));
 sg13g2_nor2_1 _3069_ (.A(_1123_),
    .B(net521),
    .Y(_0057_));
 sg13g2_nor2_1 _3070_ (.A(_1327_),
    .B(net521),
    .Y(_0058_));
 sg13g2_nor2_1 _3071_ (.A(_0372_),
    .B(net521),
    .Y(_0059_));
 sg13g2_nor2_1 _3072_ (.A(_0370_),
    .B(net521),
    .Y(_0060_));
 sg13g2_and2_1 _3073_ (.A(_0412_),
    .B(_0626_),
    .X(_0061_));
 sg13g2_nor2_1 _3074_ (.A(_0413_),
    .B(net522),
    .Y(_0062_));
 sg13g2_nor2_1 _3075_ (.A(_0417_),
    .B(net522),
    .Y(_0063_));
 sg13g2_nor2_1 _3076_ (.A(_0411_),
    .B(net522),
    .Y(_0064_));
 sg13g2_and2_1 _3077_ (.A(_0410_),
    .B(_0626_),
    .X(_0065_));
 sg13g2_nor3_1 _3078_ (.A(net6),
    .B(net7),
    .C(net8),
    .Y(_0684_));
 sg13g2_nor2_1 _3079_ (.A(net1),
    .B(net528),
    .Y(_0685_));
 sg13g2_nor4_1 _3080_ (.A(net2),
    .B(net3),
    .C(net4),
    .D(net5),
    .Y(_0686_));
 sg13g2_nand3_1 _3081_ (.B(_0685_),
    .C(_0686_),
    .A(_0684_),
    .Y(_0687_));
 sg13g2_and2_1 _3082_ (.A(net691),
    .B(_0687_),
    .X(_0066_));
 sg13g2_o21ai_1 _3083_ (.B1(_0636_),
    .Y(_0073_),
    .A1(_0447_),
    .A2(net521));
 sg13g2_nor4_1 _3084_ (.A(net578),
    .B(net536),
    .C(net524),
    .D(net523),
    .Y(_0689_));
 sg13g2_and2_1 _3085_ (.A(net522),
    .B(_0633_),
    .X(_0690_));
 sg13g2_xnor2_1 _3086_ (.Y(_0691_),
    .A(net571),
    .B(_0689_));
 sg13g2_nor2_1 _3087_ (.A(_0690_),
    .B(_0691_),
    .Y(_0074_));
 sg13g2_nor3_1 _3088_ (.A(net524),
    .B(_1069_),
    .C(net523),
    .Y(_0692_));
 sg13g2_xnor2_1 _3089_ (.Y(_0693_),
    .A(net567),
    .B(_0692_));
 sg13g2_nor2_1 _3090_ (.A(_0690_),
    .B(_0693_),
    .Y(_0075_));
 sg13g2_nor3_1 _3091_ (.A(net566),
    .B(net524),
    .C(_1069_),
    .Y(_0694_));
 sg13g2_a21oi_1 _3092_ (.A1(net562),
    .A2(_0694_),
    .Y(_0695_),
    .B1(_0635_));
 sg13g2_o21ai_1 _3093_ (.B1(_0695_),
    .Y(_0696_),
    .A1(net562),
    .A2(_0694_));
 sg13g2_o21ai_1 _3094_ (.B1(_0696_),
    .Y(_0076_),
    .A1(_0502_),
    .A2(net521));
 sg13g2_and3_1 _3095_ (.X(_0077_),
    .A(_0604_),
    .B(_0612_),
    .C(_0055_));
 sg13g2_dfrbp_1 _3096_ (.CLK(net557),
    .RESET_B(net36),
    .D(_0045_),
    .Q_N(_1538_),
    .Q(_0018_));
 sg13g2_dfrbp_1 _3097_ (.CLK(net559),
    .RESET_B(net60),
    .D(_0046_),
    .Q_N(_0044_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _3098_ (.CLK(net559),
    .RESET_B(net59),
    .D(_0047_),
    .Q_N(_1537_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _3099_ (.CLK(net559),
    .RESET_B(net58),
    .D(_0048_),
    .Q_N(_0027_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _3100_ (.CLK(net559),
    .RESET_B(net57),
    .D(_0049_),
    .Q_N(_0025_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _3101_ (.CLK(net559),
    .RESET_B(net56),
    .D(_0050_),
    .Q_N(_0024_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _3102_ (.CLK(net559),
    .RESET_B(net55),
    .D(_0051_),
    .Q_N(_0023_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _3103_ (.CLK(net558),
    .RESET_B(net54),
    .D(_0052_),
    .Q_N(_0022_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _3104_ (.CLK(net558),
    .RESET_B(net52),
    .D(_0053_),
    .Q_N(_1536_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _3105_ (.CLK(net557),
    .RESET_B(net51),
    .D(_0054_),
    .Q_N(_0034_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _3106_ (.CLK(net558),
    .RESET_B(net37),
    .D(_0055_),
    .Q_N(_1539_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _3107_ (.CLK(net557),
    .RESET_B(net38),
    .D(_0000_),
    .Q_N(_1540_),
    .Q(_0012_));
 sg13g2_dfrbp_1 _3108_ (.CLK(net557),
    .RESET_B(net39),
    .D(_0001_),
    .Q_N(_1541_),
    .Q(_0013_));
 sg13g2_dfrbp_1 _3109_ (.CLK(net558),
    .RESET_B(net40),
    .D(_0002_),
    .Q_N(_1542_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _3110_ (.CLK(net557),
    .RESET_B(net41),
    .D(_0003_),
    .Q_N(_1543_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _3111_ (.CLK(net557),
    .RESET_B(net53),
    .D(_0004_),
    .Q_N(_1544_),
    .Q(_0016_));
 sg13g2_dfrbp_1 _3112_ (.CLK(net557),
    .RESET_B(net50),
    .D(_0005_),
    .Q_N(_1535_),
    .Q(_0017_));
 sg13g2_dfrbp_1 _3113_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net49),
    .D(_0056_),
    .Q_N(\hx0[0] ),
    .Q(\gradient_sky.x[0] ));
 sg13g2_dfrbp_1 _3114_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net48),
    .D(_0057_),
    .Q_N(_0021_),
    .Q(\gradient_sky.x[1] ));
 sg13g2_dfrbp_1 _3115_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net47),
    .D(_0058_),
    .Q_N(_0040_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _3116_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net46),
    .D(_0059_),
    .Q_N(_0043_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _3117_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net45),
    .D(_0060_),
    .Q_N(_0037_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _3118_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net44),
    .D(_0061_),
    .Q_N(_0036_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _3119_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net43),
    .D(_0062_),
    .Q_N(_0035_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _3120_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net42),
    .D(_0063_),
    .Q_N(_0042_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _3121_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net35),
    .D(_0064_),
    .Q_N(_0031_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _3122_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net34),
    .D(_0065_),
    .Q_N(_0026_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _3123_ (.CLK(net557),
    .RESET_B(net64),
    .D(_0066_),
    .Q_N(_1545_),
    .Q(show));
 sg13g2_dfrbp_1 _3124_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net33),
    .D(_0010_),
    .Q_N(_1534_),
    .Q(hsync));
 sg13g2_dfrbp_1 _3125_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net32),
    .D(_0067_),
    .Q_N(\hy0[0] ),
    .Q(\gradient_sky.y[0] ));
 sg13g2_dfrbp_1 _3126_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net30),
    .D(_0068_),
    .Q_N(_0020_),
    .Q(\gradient_sky.y[1] ));
 sg13g2_dfrbp_1 _3127_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net28),
    .D(_0069_),
    .Q_N(_0041_),
    .Q(\gradient_sky.y[2] ));
 sg13g2_dfrbp_1 _3128_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net26),
    .D(_0070_),
    .Q_N(_0039_),
    .Q(\gradient_sky.y[3] ));
 sg13g2_dfrbp_1 _3129_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net69),
    .D(_0071_),
    .Q_N(_0038_),
    .Q(\gradient_sky.y[4] ));
 sg13g2_dfrbp_1 _3130_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net62),
    .D(_0072_),
    .Q_N(_0033_),
    .Q(\gradient_sky.y[5] ));
 sg13g2_dfrbp_1 _3131_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net31),
    .D(_0073_),
    .Q_N(_0032_),
    .Q(\gradient_sky.y[6] ));
 sg13g2_dfrbp_1 _3132_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net27),
    .D(_0074_),
    .Q_N(_0030_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _3133_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net63),
    .D(_0075_),
    .Q_N(_0029_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _3134_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net65),
    .D(_0076_),
    .Q_N(_0028_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _3135_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net66),
    .D(net72),
    .Q_N(_1546_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 _3136_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net67),
    .D(_0006_),
    .Q_N(_1547_),
    .Q(_0078_));
 sg13g2_dfrbp_1 _3137_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net68),
    .D(_0007_),
    .Q_N(_1548_),
    .Q(_0079_));
 sg13g2_dfrbp_1 _3138_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net25),
    .D(_0008_),
    .Q_N(_1549_),
    .Q(_0080_));
 sg13g2_dfrbp_1 _3139_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net29),
    .D(_0009_),
    .Q_N(_1533_),
    .Q(_0081_));
 sg13g2_dfrbp_1 _3140_ (.CLK(net558),
    .RESET_B(net61),
    .D(_0077_),
    .Q_N(_1532_),
    .Q(_0019_));
 sg13g2_tiehi _3128__26 (.L_HI(net26));
 sg13g2_tiehi _3132__27 (.L_HI(net27));
 sg13g2_tiehi _3127__28 (.L_HI(net28));
 sg13g2_tiehi _3139__29 (.L_HI(net29));
 sg13g2_tiehi _3126__30 (.L_HI(net30));
 sg13g2_tiehi _3131__31 (.L_HI(net31));
 sg13g2_tiehi _3125__32 (.L_HI(net32));
 sg13g2_tiehi _3124__33 (.L_HI(net33));
 sg13g2_tiehi _3122__34 (.L_HI(net34));
 sg13g2_tiehi _3121__35 (.L_HI(net35));
 sg13g2_tiehi _3096__36 (.L_HI(net36));
 sg13g2_tiehi _3106__37 (.L_HI(net37));
 sg13g2_tiehi _3107__38 (.L_HI(net38));
 sg13g2_tiehi _3108__39 (.L_HI(net39));
 sg13g2_tiehi _3109__40 (.L_HI(net40));
 sg13g2_tiehi _3110__41 (.L_HI(net41));
 sg13g2_tiehi _3120__42 (.L_HI(net42));
 sg13g2_tiehi _3119__43 (.L_HI(net43));
 sg13g2_tiehi _3118__44 (.L_HI(net44));
 sg13g2_tiehi _3117__45 (.L_HI(net45));
 sg13g2_tiehi _3116__46 (.L_HI(net46));
 sg13g2_tiehi _3115__47 (.L_HI(net47));
 sg13g2_tiehi _3114__48 (.L_HI(net48));
 sg13g2_tiehi _3113__49 (.L_HI(net49));
 sg13g2_tiehi _3112__50 (.L_HI(net50));
 sg13g2_tiehi _3105__51 (.L_HI(net51));
 sg13g2_tiehi _3104__52 (.L_HI(net52));
 sg13g2_tiehi _3111__53 (.L_HI(net53));
 sg13g2_tiehi _3103__54 (.L_HI(net54));
 sg13g2_tiehi _3102__55 (.L_HI(net55));
 sg13g2_tiehi _3101__56 (.L_HI(net56));
 sg13g2_tiehi _3100__57 (.L_HI(net57));
 sg13g2_tiehi _3099__58 (.L_HI(net58));
 sg13g2_tiehi _3098__59 (.L_HI(net59));
 sg13g2_tiehi _3097__60 (.L_HI(net60));
 sg13g2_tiehi _3140__61 (.L_HI(net61));
 sg13g2_tiehi _3130__62 (.L_HI(net62));
 sg13g2_tiehi _3133__63 (.L_HI(net63));
 sg13g2_tiehi _3123__64 (.L_HI(net64));
 sg13g2_tiehi _3134__65 (.L_HI(net65));
 sg13g2_tiehi _3135__66 (.L_HI(net66));
 sg13g2_tiehi _3136__67 (.L_HI(net67));
 sg13g2_tiehi _3137__68 (.L_HI(net68));
 sg13g2_tiehi _3129__69 (.L_HI(net69));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_nvious_graphics_10 (.L_LO(net10));
 sg13g2_tielo tt_um_nvious_graphics_11 (.L_LO(net11));
 sg13g2_tielo tt_um_nvious_graphics_12 (.L_LO(net12));
 sg13g2_tielo tt_um_nvious_graphics_13 (.L_LO(net13));
 sg13g2_tielo tt_um_nvious_graphics_14 (.L_LO(net14));
 sg13g2_tielo tt_um_nvious_graphics_15 (.L_LO(net15));
 sg13g2_tielo tt_um_nvious_graphics_16 (.L_LO(net16));
 sg13g2_tielo tt_um_nvious_graphics_17 (.L_LO(net17));
 sg13g2_tielo tt_um_nvious_graphics_18 (.L_LO(net18));
 sg13g2_tielo tt_um_nvious_graphics_19 (.L_LO(net19));
 sg13g2_tielo tt_um_nvious_graphics_20 (.L_LO(net20));
 sg13g2_tielo tt_um_nvious_graphics_21 (.L_LO(net21));
 sg13g2_tielo tt_um_nvious_graphics_22 (.L_LO(net22));
 sg13g2_tielo tt_um_nvious_graphics_23 (.L_LO(net23));
 sg13g2_tielo tt_um_nvious_graphics_24 (.L_LO(net24));
 sg13g2_tiehi _3138__25 (.L_HI(net25));
 sg13g2_buf_1 _3202_ (.A(net558),
    .X(uo_out[3]));
 sg13g2_buf_1 _3203_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(_0627_));
 sg13g2_buf_2 fanout522 (.A(_0627_),
    .X(net522));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(_0626_));
 sg13g2_buf_2 fanout524 (.A(_0941_),
    .X(net524));
 sg13g2_buf_1 fanout525 (.A(_0941_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_0856_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_0712_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net529),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(show),
    .X(net529));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(net531));
 sg13g2_buf_2 fanout531 (.A(\counter[5] ),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(\counter[3] ),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(\counter[2] ),
    .X(net533));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(net535));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(_1098_));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(_0929_));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(_0844_));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(_0825_));
 sg13g2_buf_2 fanout539 (.A(_0825_),
    .X(net539));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(_0818_));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(_0666_));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(_0648_));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(_0588_));
 sg13g2_buf_2 fanout544 (.A(_0588_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net547),
    .X(net545));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(net547));
 sg13g2_buf_2 fanout547 (.A(_0568_),
    .X(net547));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(_0535_));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(_0524_));
 sg13g2_buf_1 fanout550 (.A(_0524_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_0524_),
    .X(net551));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(_0469_));
 sg13g2_buf_2 fanout553 (.A(_0469_),
    .X(net553));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(_0436_));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(_0425_));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(_0414_));
 sg13g2_buf_2 fanout557 (.A(net558),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(\hvsync_gen.vsync ),
    .X(net559));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(net561));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(net562));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(net71));
 sg13g2_buf_4 fanout563 (.X(net563),
    .A(net565));
 sg13g2_buf_2 fanout564 (.A(net565),
    .X(net564));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(net566));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(_0029_));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(net73));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(\hvsync_gen.vpos[8] ));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(_0030_));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(_0030_));
 sg13g2_buf_4 fanout571 (.X(net571),
    .A(net574));
 sg13g2_buf_2 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(\hvsync_gen.vpos[7] ),
    .X(net574));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(net577));
 sg13g2_buf_2 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_4 fanout577 (.X(net577),
    .A(net578));
 sg13g2_buf_2 fanout578 (.A(net75),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(\gradient_sky.y[6] ),
    .X(net579));
 sg13g2_buf_4 fanout580 (.X(net580),
    .A(\gradient_sky.y[6] ));
 sg13g2_buf_4 fanout581 (.X(net581),
    .A(\gradient_sky.y[6] ));
 sg13g2_buf_4 fanout582 (.X(net582),
    .A(net583));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(net584));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(_0033_));
 sg13g2_buf_2 fanout585 (.A(\gradient_sky.y[5] ),
    .X(net585));
 sg13g2_buf_4 fanout586 (.X(net586),
    .A(\gradient_sky.y[5] ));
 sg13g2_buf_4 fanout587 (.X(net587),
    .A(_0038_));
 sg13g2_buf_2 fanout588 (.A(net591),
    .X(net588));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(net591));
 sg13g2_buf_2 fanout590 (.A(net591),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(\gradient_sky.y[4] ),
    .X(net591));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(net593));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(_0039_));
 sg13g2_buf_2 fanout594 (.A(net599),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(net599),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(net599),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(net599),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(\gradient_sky.y[3] ),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(net601),
    .X(net600));
 sg13g2_buf_4 fanout601 (.X(net601),
    .A(_0041_));
 sg13g2_buf_2 fanout602 (.A(_0041_),
    .X(net602));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(\gradient_sky.y[2] ));
 sg13g2_buf_2 fanout604 (.A(\gradient_sky.y[2] ),
    .X(net604));
 sg13g2_buf_4 fanout605 (.X(net605),
    .A(net606));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(_0020_));
 sg13g2_buf_4 fanout607 (.X(net607),
    .A(net609));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(net609));
 sg13g2_buf_2 fanout609 (.A(\gradient_sky.y[1] ),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(\hy0[0] ),
    .X(net610));
 sg13g2_buf_4 fanout611 (.X(net611),
    .A(net612));
 sg13g2_buf_4 fanout612 (.X(net612),
    .A(\gradient_sky.y[0] ));
 sg13g2_buf_4 fanout613 (.X(net613),
    .A(\gradient_sky.y[0] ));
 sg13g2_buf_2 fanout614 (.A(\gradient_sky.y[0] ),
    .X(net614));
 sg13g2_buf_4 fanout615 (.X(net615),
    .A(net74));
 sg13g2_buf_2 fanout616 (.A(_0026_),
    .X(net616));
 sg13g2_buf_4 fanout617 (.X(net617),
    .A(net619));
 sg13g2_buf_2 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_4 fanout619 (.X(net619),
    .A(\hvsync_gen.hpos[9] ));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(net623));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(net622));
 sg13g2_buf_2 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_0031_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(net626),
    .X(net624));
 sg13g2_buf_4 fanout625 (.X(net625),
    .A(net626));
 sg13g2_buf_2 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(\hvsync_gen.hpos[8] ));
 sg13g2_buf_4 fanout628 (.X(net628),
    .A(_0042_));
 sg13g2_buf_2 fanout629 (.A(_0042_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(net631),
    .X(net630));
 sg13g2_buf_4 fanout631 (.X(net631),
    .A(net76));
 sg13g2_buf_2 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(\hvsync_gen.hpos[7] ),
    .X(net633));
 sg13g2_buf_4 fanout634 (.X(net634),
    .A(_0035_));
 sg13g2_buf_2 fanout635 (.A(_0035_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net637),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_buf_2 fanout639 (.A(net642),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(net642),
    .X(net640));
 sg13g2_buf_4 fanout641 (.X(net641),
    .A(net642));
 sg13g2_buf_2 fanout642 (.A(\hvsync_gen.hpos[6] ),
    .X(net642));
 sg13g2_buf_4 fanout643 (.X(net643),
    .A(_0036_));
 sg13g2_buf_4 fanout644 (.X(net644),
    .A(net646));
 sg13g2_buf_2 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(net649),
    .X(net646));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(net648));
 sg13g2_buf_2 fanout648 (.A(net649),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(\hvsync_gen.hpos[5] ),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_4 fanout651 (.X(net651),
    .A(_0037_));
 sg13g2_buf_4 fanout652 (.X(net652),
    .A(net654));
 sg13g2_buf_2 fanout653 (.A(net654),
    .X(net653));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(net657));
 sg13g2_buf_2 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(net657),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(\hvsync_gen.hpos[4] ),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(net659),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_0043_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(net665),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(net664),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(net664),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_1 fanout665 (.A(net668),
    .X(net665));
 sg13g2_buf_4 fanout666 (.X(net666),
    .A(net667));
 sg13g2_buf_2 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(\hvsync_gen.hpos[3] ),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net671),
    .X(net669));
 sg13g2_buf_1 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_1 fanout671 (.A(_0040_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net675),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(net674),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(net675),
    .X(net674));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(\hvsync_gen.hpos[2] ));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(net678));
 sg13g2_buf_1 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(\hvsync_gen.hpos[2] ));
 sg13g2_buf_2 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(net681),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(net684),
    .X(net681));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(net684));
 sg13g2_buf_2 fanout683 (.A(net684),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(\gradient_sky.x[1] ),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(net686),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_1 fanout687 (.A(\gradient_sky.x[0] ),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(\gradient_sky.x[0] ),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(\gradient_sky.x[0] ),
    .X(net689));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(rst_n));
 sg13g2_buf_2 fanout691 (.A(rst_n),
    .X(net691));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_nvious_graphics_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\hx0[0] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold2 (.A(\hvsync_gen.vpos[9] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0011_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold4 (.A(\hvsync_gen.vpos[8] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0026_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0032_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold7 (.A(\hvsync_gen.hpos[7] ),
    .X(net76));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_fill_1 FILLER_4_56 ();
 sg13g2_fill_2 FILLER_4_66 ();
 sg13g2_fill_1 FILLER_4_68 ();
 sg13g2_decap_8 FILLER_4_75 ();
 sg13g2_decap_8 FILLER_4_82 ();
 sg13g2_decap_8 FILLER_4_89 ();
 sg13g2_fill_2 FILLER_4_96 ();
 sg13g2_fill_1 FILLER_4_98 ();
 sg13g2_fill_2 FILLER_4_108 ();
 sg13g2_fill_1 FILLER_4_110 ();
 sg13g2_decap_8 FILLER_4_115 ();
 sg13g2_decap_8 FILLER_4_122 ();
 sg13g2_decap_8 FILLER_4_129 ();
 sg13g2_fill_1 FILLER_4_136 ();
 sg13g2_decap_8 FILLER_4_142 ();
 sg13g2_decap_8 FILLER_4_149 ();
 sg13g2_decap_8 FILLER_4_187 ();
 sg13g2_decap_8 FILLER_4_194 ();
 sg13g2_fill_2 FILLER_4_201 ();
 sg13g2_fill_1 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_230 ();
 sg13g2_decap_8 FILLER_4_237 ();
 sg13g2_decap_8 FILLER_4_244 ();
 sg13g2_decap_8 FILLER_4_251 ();
 sg13g2_decap_8 FILLER_4_258 ();
 sg13g2_decap_8 FILLER_4_265 ();
 sg13g2_decap_8 FILLER_4_272 ();
 sg13g2_decap_8 FILLER_4_279 ();
 sg13g2_decap_8 FILLER_4_286 ();
 sg13g2_decap_8 FILLER_4_293 ();
 sg13g2_decap_4 FILLER_4_300 ();
 sg13g2_decap_8 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_344 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_11 ();
 sg13g2_decap_4 FILLER_5_17 ();
 sg13g2_fill_2 FILLER_5_55 ();
 sg13g2_fill_1 FILLER_5_57 ();
 sg13g2_fill_1 FILLER_5_133 ();
 sg13g2_fill_2 FILLER_5_141 ();
 sg13g2_fill_2 FILLER_5_151 ();
 sg13g2_fill_1 FILLER_5_153 ();
 sg13g2_fill_2 FILLER_5_207 ();
 sg13g2_decap_4 FILLER_5_234 ();
 sg13g2_fill_1 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_decap_8 FILLER_5_251 ();
 sg13g2_decap_4 FILLER_5_266 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_fill_2 FILLER_5_280 ();
 sg13g2_fill_1 FILLER_5_282 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_4 FILLER_5_298 ();
 sg13g2_fill_2 FILLER_5_302 ();
 sg13g2_fill_2 FILLER_5_308 ();
 sg13g2_fill_1 FILLER_5_310 ();
 sg13g2_decap_4 FILLER_5_320 ();
 sg13g2_fill_2 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_37 ();
 sg13g2_fill_2 FILLER_6_43 ();
 sg13g2_fill_2 FILLER_6_53 ();
 sg13g2_fill_2 FILLER_6_62 ();
 sg13g2_fill_2 FILLER_6_69 ();
 sg13g2_fill_1 FILLER_6_71 ();
 sg13g2_fill_2 FILLER_6_77 ();
 sg13g2_fill_2 FILLER_6_87 ();
 sg13g2_fill_1 FILLER_6_89 ();
 sg13g2_fill_1 FILLER_6_94 ();
 sg13g2_fill_2 FILLER_6_99 ();
 sg13g2_fill_1 FILLER_6_101 ();
 sg13g2_fill_2 FILLER_6_107 ();
 sg13g2_fill_2 FILLER_6_129 ();
 sg13g2_fill_1 FILLER_6_131 ();
 sg13g2_decap_4 FILLER_6_136 ();
 sg13g2_fill_2 FILLER_6_145 ();
 sg13g2_decap_4 FILLER_6_155 ();
 sg13g2_fill_2 FILLER_6_159 ();
 sg13g2_fill_2 FILLER_6_167 ();
 sg13g2_decap_4 FILLER_6_177 ();
 sg13g2_fill_1 FILLER_6_181 ();
 sg13g2_fill_2 FILLER_6_191 ();
 sg13g2_decap_4 FILLER_6_202 ();
 sg13g2_decap_4 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_fill_1 FILLER_6_252 ();
 sg13g2_fill_2 FILLER_6_271 ();
 sg13g2_fill_1 FILLER_6_273 ();
 sg13g2_fill_2 FILLER_6_295 ();
 sg13g2_fill_1 FILLER_6_297 ();
 sg13g2_fill_1 FILLER_6_320 ();
 sg13g2_fill_2 FILLER_6_338 ();
 sg13g2_fill_1 FILLER_6_340 ();
 sg13g2_fill_2 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_4 ();
 sg13g2_fill_1 FILLER_7_13 ();
 sg13g2_fill_2 FILLER_7_26 ();
 sg13g2_fill_1 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_39 ();
 sg13g2_fill_1 FILLER_7_41 ();
 sg13g2_fill_2 FILLER_7_49 ();
 sg13g2_fill_1 FILLER_7_83 ();
 sg13g2_fill_1 FILLER_7_89 ();
 sg13g2_fill_2 FILLER_7_105 ();
 sg13g2_decap_4 FILLER_7_117 ();
 sg13g2_fill_2 FILLER_7_141 ();
 sg13g2_fill_1 FILLER_7_143 ();
 sg13g2_decap_4 FILLER_7_189 ();
 sg13g2_fill_2 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_246 ();
 sg13g2_fill_1 FILLER_7_255 ();
 sg13g2_fill_2 FILLER_7_265 ();
 sg13g2_decap_4 FILLER_7_277 ();
 sg13g2_fill_2 FILLER_7_281 ();
 sg13g2_decap_4 FILLER_7_287 ();
 sg13g2_decap_4 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_fill_2 FILLER_7_320 ();
 sg13g2_decap_4 FILLER_7_342 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_fill_1 FILLER_7_365 ();
 sg13g2_decap_4 FILLER_7_397 ();
 sg13g2_fill_2 FILLER_7_401 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_4 ();
 sg13g2_decap_4 FILLER_8_36 ();
 sg13g2_fill_2 FILLER_8_69 ();
 sg13g2_fill_2 FILLER_8_80 ();
 sg13g2_fill_1 FILLER_8_82 ();
 sg13g2_fill_2 FILLER_8_88 ();
 sg13g2_fill_2 FILLER_8_94 ();
 sg13g2_decap_4 FILLER_8_116 ();
 sg13g2_fill_2 FILLER_8_124 ();
 sg13g2_fill_1 FILLER_8_126 ();
 sg13g2_fill_2 FILLER_8_147 ();
 sg13g2_fill_2 FILLER_8_162 ();
 sg13g2_fill_1 FILLER_8_181 ();
 sg13g2_fill_1 FILLER_8_206 ();
 sg13g2_decap_4 FILLER_8_211 ();
 sg13g2_fill_1 FILLER_8_215 ();
 sg13g2_decap_4 FILLER_8_236 ();
 sg13g2_fill_1 FILLER_8_240 ();
 sg13g2_decap_4 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_271 ();
 sg13g2_decap_8 FILLER_8_303 ();
 sg13g2_fill_2 FILLER_8_310 ();
 sg13g2_fill_1 FILLER_8_312 ();
 sg13g2_fill_2 FILLER_8_319 ();
 sg13g2_fill_2 FILLER_8_341 ();
 sg13g2_decap_4 FILLER_8_377 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_27 ();
 sg13g2_fill_1 FILLER_9_34 ();
 sg13g2_decap_4 FILLER_9_59 ();
 sg13g2_fill_1 FILLER_9_87 ();
 sg13g2_fill_1 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_123 ();
 sg13g2_fill_1 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_131 ();
 sg13g2_decap_8 FILLER_9_138 ();
 sg13g2_fill_1 FILLER_9_145 ();
 sg13g2_fill_2 FILLER_9_162 ();
 sg13g2_fill_1 FILLER_9_164 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_fill_1 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_fill_2 FILLER_9_214 ();
 sg13g2_fill_1 FILLER_9_216 ();
 sg13g2_decap_4 FILLER_9_227 ();
 sg13g2_decap_4 FILLER_9_239 ();
 sg13g2_decap_4 FILLER_9_256 ();
 sg13g2_fill_2 FILLER_9_260 ();
 sg13g2_fill_2 FILLER_9_284 ();
 sg13g2_fill_2 FILLER_9_331 ();
 sg13g2_fill_1 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_4 FILLER_9_357 ();
 sg13g2_fill_2 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_374 ();
 sg13g2_decap_4 FILLER_9_381 ();
 sg13g2_fill_2 FILLER_9_393 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_fill_2 FILLER_10_23 ();
 sg13g2_fill_1 FILLER_10_25 ();
 sg13g2_fill_1 FILLER_10_36 ();
 sg13g2_fill_2 FILLER_10_58 ();
 sg13g2_decap_8 FILLER_10_85 ();
 sg13g2_fill_1 FILLER_10_111 ();
 sg13g2_fill_2 FILLER_10_137 ();
 sg13g2_fill_1 FILLER_10_152 ();
 sg13g2_fill_2 FILLER_10_166 ();
 sg13g2_fill_2 FILLER_10_181 ();
 sg13g2_fill_1 FILLER_10_203 ();
 sg13g2_fill_1 FILLER_10_216 ();
 sg13g2_fill_1 FILLER_10_225 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_fill_1 FILLER_10_233 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_fill_2 FILLER_10_259 ();
 sg13g2_fill_1 FILLER_10_261 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_decap_4 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_fill_2 FILLER_10_321 ();
 sg13g2_fill_2 FILLER_10_329 ();
 sg13g2_fill_2 FILLER_10_335 ();
 sg13g2_fill_1 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_369 ();
 sg13g2_fill_1 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_45 ();
 sg13g2_decap_4 FILLER_11_57 ();
 sg13g2_fill_2 FILLER_11_79 ();
 sg13g2_fill_2 FILLER_11_86 ();
 sg13g2_fill_2 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_113 ();
 sg13g2_fill_2 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_131 ();
 sg13g2_fill_1 FILLER_11_136 ();
 sg13g2_fill_2 FILLER_11_141 ();
 sg13g2_fill_1 FILLER_11_143 ();
 sg13g2_fill_2 FILLER_11_149 ();
 sg13g2_fill_1 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_fill_2 FILLER_11_172 ();
 sg13g2_fill_1 FILLER_11_174 ();
 sg13g2_fill_2 FILLER_11_200 ();
 sg13g2_fill_1 FILLER_11_207 ();
 sg13g2_fill_2 FILLER_11_213 ();
 sg13g2_decap_4 FILLER_11_220 ();
 sg13g2_fill_2 FILLER_11_255 ();
 sg13g2_fill_1 FILLER_11_257 ();
 sg13g2_decap_4 FILLER_11_320 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_decap_4 FILLER_11_337 ();
 sg13g2_fill_1 FILLER_11_341 ();
 sg13g2_fill_1 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_356 ();
 sg13g2_decap_4 FILLER_11_363 ();
 sg13g2_fill_1 FILLER_11_382 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_9 ();
 sg13g2_fill_1 FILLER_12_26 ();
 sg13g2_fill_2 FILLER_12_46 ();
 sg13g2_fill_2 FILLER_12_54 ();
 sg13g2_fill_2 FILLER_12_66 ();
 sg13g2_fill_1 FILLER_12_68 ();
 sg13g2_decap_4 FILLER_12_73 ();
 sg13g2_fill_2 FILLER_12_93 ();
 sg13g2_fill_2 FILLER_12_123 ();
 sg13g2_fill_1 FILLER_12_125 ();
 sg13g2_fill_2 FILLER_12_147 ();
 sg13g2_fill_1 FILLER_12_164 ();
 sg13g2_decap_4 FILLER_12_182 ();
 sg13g2_fill_2 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_215 ();
 sg13g2_fill_2 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_230 ();
 sg13g2_fill_1 FILLER_12_243 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_4 FILLER_12_259 ();
 sg13g2_fill_1 FILLER_12_263 ();
 sg13g2_decap_4 FILLER_12_286 ();
 sg13g2_decap_4 FILLER_12_310 ();
 sg13g2_fill_1 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_13 ();
 sg13g2_fill_1 FILLER_13_24 ();
 sg13g2_fill_1 FILLER_13_31 ();
 sg13g2_fill_2 FILLER_13_37 ();
 sg13g2_fill_1 FILLER_13_39 ();
 sg13g2_decap_4 FILLER_13_54 ();
 sg13g2_fill_2 FILLER_13_58 ();
 sg13g2_decap_4 FILLER_13_72 ();
 sg13g2_fill_2 FILLER_13_76 ();
 sg13g2_decap_8 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_106 ();
 sg13g2_fill_1 FILLER_13_108 ();
 sg13g2_fill_1 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_125 ();
 sg13g2_decap_4 FILLER_13_131 ();
 sg13g2_fill_2 FILLER_13_135 ();
 sg13g2_fill_2 FILLER_13_156 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_fill_2 FILLER_13_170 ();
 sg13g2_fill_1 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_185 ();
 sg13g2_decap_8 FILLER_13_192 ();
 sg13g2_fill_2 FILLER_13_218 ();
 sg13g2_fill_2 FILLER_13_239 ();
 sg13g2_fill_1 FILLER_13_241 ();
 sg13g2_fill_2 FILLER_13_247 ();
 sg13g2_fill_2 FILLER_13_272 ();
 sg13g2_fill_1 FILLER_13_274 ();
 sg13g2_fill_2 FILLER_13_280 ();
 sg13g2_fill_1 FILLER_13_282 ();
 sg13g2_decap_4 FILLER_13_293 ();
 sg13g2_fill_2 FILLER_13_312 ();
 sg13g2_fill_1 FILLER_13_327 ();
 sg13g2_fill_2 FILLER_13_337 ();
 sg13g2_fill_2 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_fill_2 FILLER_13_377 ();
 sg13g2_fill_1 FILLER_13_379 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_54 ();
 sg13g2_decap_4 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_130 ();
 sg13g2_fill_2 FILLER_14_177 ();
 sg13g2_fill_2 FILLER_14_193 ();
 sg13g2_fill_1 FILLER_14_195 ();
 sg13g2_fill_2 FILLER_14_200 ();
 sg13g2_fill_2 FILLER_14_216 ();
 sg13g2_decap_4 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_250 ();
 sg13g2_fill_2 FILLER_14_269 ();
 sg13g2_fill_2 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_278 ();
 sg13g2_decap_4 FILLER_14_294 ();
 sg13g2_fill_2 FILLER_14_311 ();
 sg13g2_fill_2 FILLER_14_327 ();
 sg13g2_fill_1 FILLER_14_341 ();
 sg13g2_fill_2 FILLER_14_361 ();
 sg13g2_decap_4 FILLER_14_381 ();
 sg13g2_fill_1 FILLER_14_385 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_31 ();
 sg13g2_fill_2 FILLER_15_53 ();
 sg13g2_fill_1 FILLER_15_55 ();
 sg13g2_decap_8 FILLER_15_69 ();
 sg13g2_fill_2 FILLER_15_76 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_fill_1 FILLER_15_87 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_fill_2 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_125 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_fill_2 FILLER_15_140 ();
 sg13g2_fill_1 FILLER_15_142 ();
 sg13g2_decap_8 FILLER_15_153 ();
 sg13g2_decap_8 FILLER_15_169 ();
 sg13g2_fill_2 FILLER_15_176 ();
 sg13g2_fill_1 FILLER_15_178 ();
 sg13g2_fill_1 FILLER_15_184 ();
 sg13g2_decap_4 FILLER_15_190 ();
 sg13g2_fill_1 FILLER_15_194 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_221 ();
 sg13g2_fill_1 FILLER_15_223 ();
 sg13g2_fill_2 FILLER_15_229 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_decap_4 FILLER_15_274 ();
 sg13g2_fill_2 FILLER_15_278 ();
 sg13g2_fill_2 FILLER_15_292 ();
 sg13g2_fill_1 FILLER_15_294 ();
 sg13g2_fill_1 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_fill_2 FILLER_15_318 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_fill_2 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_4 FILLER_15_341 ();
 sg13g2_fill_2 FILLER_15_345 ();
 sg13g2_fill_2 FILLER_15_364 ();
 sg13g2_fill_1 FILLER_15_383 ();
 sg13g2_fill_2 FILLER_15_389 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_16 ();
 sg13g2_decap_8 FILLER_16_27 ();
 sg13g2_fill_1 FILLER_16_34 ();
 sg13g2_fill_2 FILLER_16_73 ();
 sg13g2_fill_1 FILLER_16_75 ();
 sg13g2_fill_1 FILLER_16_82 ();
 sg13g2_fill_2 FILLER_16_93 ();
 sg13g2_fill_1 FILLER_16_95 ();
 sg13g2_decap_4 FILLER_16_100 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_fill_1 FILLER_16_129 ();
 sg13g2_fill_1 FILLER_16_149 ();
 sg13g2_fill_2 FILLER_16_174 ();
 sg13g2_fill_1 FILLER_16_176 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_decap_4 FILLER_16_198 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_decap_4 FILLER_16_208 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_decap_8 FILLER_16_241 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_fill_1 FILLER_16_255 ();
 sg13g2_fill_2 FILLER_16_271 ();
 sg13g2_fill_1 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_299 ();
 sg13g2_fill_1 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_fill_2 FILLER_16_323 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_decap_4 FILLER_16_366 ();
 sg13g2_fill_2 FILLER_16_383 ();
 sg13g2_fill_1 FILLER_16_385 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_25 ();
 sg13g2_fill_1 FILLER_17_27 ();
 sg13g2_fill_2 FILLER_17_33 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_fill_1 FILLER_17_58 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_4 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_104 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_fill_2 FILLER_17_120 ();
 sg13g2_fill_1 FILLER_17_122 ();
 sg13g2_fill_2 FILLER_17_146 ();
 sg13g2_fill_1 FILLER_17_148 ();
 sg13g2_fill_1 FILLER_17_186 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_fill_2 FILLER_17_200 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_fill_1 FILLER_17_208 ();
 sg13g2_fill_2 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_fill_2 FILLER_17_225 ();
 sg13g2_fill_1 FILLER_17_244 ();
 sg13g2_fill_2 FILLER_17_253 ();
 sg13g2_fill_2 FILLER_17_278 ();
 sg13g2_fill_2 FILLER_17_284 ();
 sg13g2_fill_1 FILLER_17_286 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_fill_2 FILLER_17_312 ();
 sg13g2_fill_2 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_332 ();
 sg13g2_decap_4 FILLER_17_339 ();
 sg13g2_fill_1 FILLER_17_343 ();
 sg13g2_fill_1 FILLER_17_354 ();
 sg13g2_fill_2 FILLER_17_375 ();
 sg13g2_fill_1 FILLER_17_377 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_19 ();
 sg13g2_decap_4 FILLER_18_36 ();
 sg13g2_decap_4 FILLER_18_52 ();
 sg13g2_fill_2 FILLER_18_56 ();
 sg13g2_fill_2 FILLER_18_84 ();
 sg13g2_decap_4 FILLER_18_94 ();
 sg13g2_fill_1 FILLER_18_98 ();
 sg13g2_fill_2 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_122 ();
 sg13g2_decap_4 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_135 ();
 sg13g2_fill_1 FILLER_18_141 ();
 sg13g2_decap_8 FILLER_18_146 ();
 sg13g2_decap_4 FILLER_18_153 ();
 sg13g2_fill_1 FILLER_18_157 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_fill_2 FILLER_18_170 ();
 sg13g2_fill_1 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_fill_1 FILLER_18_195 ();
 sg13g2_fill_2 FILLER_18_201 ();
 sg13g2_fill_1 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_214 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_251 ();
 sg13g2_fill_2 FILLER_18_256 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_fill_2 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_4 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_323 ();
 sg13g2_fill_1 FILLER_18_335 ();
 sg13g2_fill_2 FILLER_18_353 ();
 sg13g2_fill_2 FILLER_18_371 ();
 sg13g2_fill_1 FILLER_18_373 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_decap_4 FILLER_19_31 ();
 sg13g2_decap_8 FILLER_19_43 ();
 sg13g2_decap_4 FILLER_19_50 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_fill_1 FILLER_19_73 ();
 sg13g2_decap_4 FILLER_19_92 ();
 sg13g2_fill_2 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_138 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_decap_4 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_198 ();
 sg13g2_decap_4 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_249 ();
 sg13g2_fill_1 FILLER_19_259 ();
 sg13g2_fill_2 FILLER_19_271 ();
 sg13g2_fill_2 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_294 ();
 sg13g2_decap_4 FILLER_19_303 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_fill_2 FILLER_19_333 ();
 sg13g2_fill_2 FILLER_19_350 ();
 sg13g2_fill_1 FILLER_19_352 ();
 sg13g2_fill_2 FILLER_19_384 ();
 sg13g2_fill_1 FILLER_19_386 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_15 ();
 sg13g2_fill_1 FILLER_20_17 ();
 sg13g2_decap_8 FILLER_20_26 ();
 sg13g2_decap_8 FILLER_20_33 ();
 sg13g2_fill_2 FILLER_20_40 ();
 sg13g2_fill_1 FILLER_20_47 ();
 sg13g2_fill_2 FILLER_20_61 ();
 sg13g2_fill_2 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_74 ();
 sg13g2_fill_1 FILLER_20_83 ();
 sg13g2_fill_2 FILLER_20_102 ();
 sg13g2_fill_1 FILLER_20_104 ();
 sg13g2_decap_8 FILLER_20_113 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_125 ();
 sg13g2_decap_8 FILLER_20_134 ();
 sg13g2_decap_8 FILLER_20_141 ();
 sg13g2_decap_4 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_152 ();
 sg13g2_fill_2 FILLER_20_159 ();
 sg13g2_fill_1 FILLER_20_161 ();
 sg13g2_fill_1 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_195 ();
 sg13g2_decap_8 FILLER_20_211 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_4 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_246 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_fill_2 FILLER_20_271 ();
 sg13g2_fill_1 FILLER_20_281 ();
 sg13g2_fill_2 FILLER_20_291 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_decap_8 FILLER_20_334 ();
 sg13g2_fill_1 FILLER_20_341 ();
 sg13g2_fill_2 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_352 ();
 sg13g2_decap_4 FILLER_20_374 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_53 ();
 sg13g2_fill_1 FILLER_21_55 ();
 sg13g2_fill_2 FILLER_21_136 ();
 sg13g2_fill_1 FILLER_21_170 ();
 sg13g2_fill_2 FILLER_21_179 ();
 sg13g2_fill_2 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_205 ();
 sg13g2_fill_1 FILLER_21_246 ();
 sg13g2_fill_2 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_decap_4 FILLER_21_267 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_300 ();
 sg13g2_decap_8 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_360 ();
 sg13g2_decap_4 FILLER_21_383 ();
 sg13g2_fill_2 FILLER_21_387 ();
 sg13g2_fill_1 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_16 ();
 sg13g2_fill_1 FILLER_22_18 ();
 sg13g2_fill_2 FILLER_22_34 ();
 sg13g2_decap_8 FILLER_22_71 ();
 sg13g2_decap_4 FILLER_22_78 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_fill_1 FILLER_22_97 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_fill_1 FILLER_22_108 ();
 sg13g2_fill_1 FILLER_22_124 ();
 sg13g2_fill_2 FILLER_22_130 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_142 ();
 sg13g2_fill_2 FILLER_22_148 ();
 sg13g2_fill_1 FILLER_22_150 ();
 sg13g2_fill_2 FILLER_22_155 ();
 sg13g2_decap_4 FILLER_22_162 ();
 sg13g2_fill_1 FILLER_22_166 ();
 sg13g2_fill_1 FILLER_22_181 ();
 sg13g2_decap_8 FILLER_22_192 ();
 sg13g2_decap_8 FILLER_22_211 ();
 sg13g2_decap_8 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_decap_8 FILLER_22_239 ();
 sg13g2_fill_1 FILLER_22_287 ();
 sg13g2_fill_2 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_296 ();
 sg13g2_fill_1 FILLER_22_307 ();
 sg13g2_fill_1 FILLER_22_313 ();
 sg13g2_fill_2 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_4 FILLER_22_349 ();
 sg13g2_decap_4 FILLER_22_357 ();
 sg13g2_fill_2 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_367 ();
 sg13g2_fill_2 FILLER_22_389 ();
 sg13g2_fill_1 FILLER_22_391 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_2 FILLER_23_35 ();
 sg13g2_decap_4 FILLER_23_84 ();
 sg13g2_fill_1 FILLER_23_88 ();
 sg13g2_decap_4 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_115 ();
 sg13g2_fill_2 FILLER_23_130 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_158 ();
 sg13g2_fill_2 FILLER_23_174 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_4 FILLER_23_217 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_decap_8 FILLER_23_265 ();
 sg13g2_fill_1 FILLER_23_272 ();
 sg13g2_decap_4 FILLER_23_289 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_decap_4 FILLER_23_302 ();
 sg13g2_fill_1 FILLER_23_306 ();
 sg13g2_decap_4 FILLER_23_318 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_fill_2 FILLER_23_374 ();
 sg13g2_fill_1 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_36 ();
 sg13g2_fill_2 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_65 ();
 sg13g2_fill_1 FILLER_24_71 ();
 sg13g2_decap_4 FILLER_24_103 ();
 sg13g2_fill_2 FILLER_24_141 ();
 sg13g2_decap_4 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_169 ();
 sg13g2_decap_4 FILLER_24_195 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_fill_2 FILLER_24_264 ();
 sg13g2_decap_4 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_decap_4 FILLER_24_387 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_26 ();
 sg13g2_decap_8 FILLER_25_33 ();
 sg13g2_decap_8 FILLER_25_40 ();
 sg13g2_fill_2 FILLER_25_47 ();
 sg13g2_decap_4 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_fill_2 FILLER_25_72 ();
 sg13g2_fill_1 FILLER_25_74 ();
 sg13g2_fill_1 FILLER_25_84 ();
 sg13g2_fill_2 FILLER_25_108 ();
 sg13g2_fill_2 FILLER_25_132 ();
 sg13g2_fill_1 FILLER_25_139 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_167 ();
 sg13g2_decap_4 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_239 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_289 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_decap_4 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_31 ();
 sg13g2_decap_4 FILLER_26_38 ();
 sg13g2_fill_1 FILLER_26_42 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_decap_8 FILLER_26_99 ();
 sg13g2_decap_4 FILLER_26_106 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_fill_2 FILLER_26_134 ();
 sg13g2_decap_4 FILLER_26_147 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_fill_1 FILLER_26_156 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_173 ();
 sg13g2_fill_2 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_221 ();
 sg13g2_decap_4 FILLER_26_244 ();
 sg13g2_fill_1 FILLER_26_248 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_decap_4 FILLER_26_311 ();
 sg13g2_fill_2 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_fill_2 FILLER_26_373 ();
 sg13g2_fill_1 FILLER_26_375 ();
 sg13g2_fill_2 FILLER_26_390 ();
 sg13g2_fill_1 FILLER_26_392 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_51 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_100 ();
 sg13g2_fill_1 FILLER_27_102 ();
 sg13g2_fill_1 FILLER_27_111 ();
 sg13g2_fill_1 FILLER_27_122 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_decap_4 FILLER_27_147 ();
 sg13g2_fill_2 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_157 ();
 sg13g2_decap_8 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_176 ();
 sg13g2_fill_2 FILLER_27_181 ();
 sg13g2_decap_4 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_192 ();
 sg13g2_decap_4 FILLER_27_210 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_221 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_4 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_265 ();
 sg13g2_decap_4 FILLER_27_290 ();
 sg13g2_fill_1 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_319 ();
 sg13g2_fill_2 FILLER_27_332 ();
 sg13g2_decap_4 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_fill_2 FILLER_27_364 ();
 sg13g2_fill_1 FILLER_27_371 ();
 sg13g2_decap_4 FILLER_27_377 ();
 sg13g2_fill_1 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_fill_1 FILLER_27_393 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_27 ();
 sg13g2_fill_1 FILLER_28_29 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_125 ();
 sg13g2_fill_2 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_197 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_decap_4 FILLER_28_239 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_decap_4 FILLER_28_257 ();
 sg13g2_fill_1 FILLER_28_261 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_4 FILLER_28_315 ();
 sg13g2_fill_1 FILLER_28_319 ();
 sg13g2_fill_2 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_decap_4 FILLER_28_353 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_fill_2 FILLER_28_369 ();
 sg13g2_fill_1 FILLER_28_371 ();
 sg13g2_fill_2 FILLER_28_395 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_34 ();
 sg13g2_decap_4 FILLER_29_43 ();
 sg13g2_decap_4 FILLER_29_59 ();
 sg13g2_fill_2 FILLER_29_63 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_fill_2 FILLER_29_79 ();
 sg13g2_fill_1 FILLER_29_81 ();
 sg13g2_fill_2 FILLER_29_87 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_decap_4 FILLER_29_124 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_decap_4 FILLER_29_142 ();
 sg13g2_fill_2 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_153 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_fill_2 FILLER_29_176 ();
 sg13g2_decap_8 FILLER_29_194 ();
 sg13g2_fill_2 FILLER_29_201 ();
 sg13g2_fill_2 FILLER_29_216 ();
 sg13g2_fill_1 FILLER_29_218 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_decap_8 FILLER_29_274 ();
 sg13g2_fill_2 FILLER_29_281 ();
 sg13g2_decap_4 FILLER_29_306 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_350 ();
 sg13g2_fill_2 FILLER_29_366 ();
 sg13g2_fill_2 FILLER_29_389 ();
 sg13g2_fill_1 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_24 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_32 ();
 sg13g2_fill_1 FILLER_30_34 ();
 sg13g2_fill_1 FILLER_30_69 ();
 sg13g2_fill_2 FILLER_30_78 ();
 sg13g2_fill_1 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_92 ();
 sg13g2_decap_4 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_102 ();
 sg13g2_fill_2 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_137 ();
 sg13g2_decap_4 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_decap_8 FILLER_30_186 ();
 sg13g2_decap_4 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_235 ();
 sg13g2_fill_2 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_decap_4 FILLER_30_269 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_decap_4 FILLER_30_325 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_334 ();
 sg13g2_fill_2 FILLER_30_341 ();
 sg13g2_fill_1 FILLER_30_343 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_fill_1 FILLER_30_360 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_45 ();
 sg13g2_decap_4 FILLER_31_62 ();
 sg13g2_fill_2 FILLER_31_66 ();
 sg13g2_fill_2 FILLER_31_97 ();
 sg13g2_fill_1 FILLER_31_99 ();
 sg13g2_fill_1 FILLER_31_111 ();
 sg13g2_fill_2 FILLER_31_116 ();
 sg13g2_decap_4 FILLER_31_155 ();
 sg13g2_fill_1 FILLER_31_159 ();
 sg13g2_fill_2 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_decap_8 FILLER_31_207 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_2 FILLER_31_236 ();
 sg13g2_fill_1 FILLER_31_238 ();
 sg13g2_decap_4 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_349 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_decap_4 FILLER_31_367 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_24 ();
 sg13g2_fill_1 FILLER_32_28 ();
 sg13g2_fill_2 FILLER_32_34 ();
 sg13g2_fill_1 FILLER_32_36 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_78 ();
 sg13g2_fill_1 FILLER_32_80 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_decap_8 FILLER_32_100 ();
 sg13g2_fill_1 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_143 ();
 sg13g2_fill_2 FILLER_32_156 ();
 sg13g2_fill_1 FILLER_32_158 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_decap_4 FILLER_32_176 ();
 sg13g2_decap_4 FILLER_32_185 ();
 sg13g2_fill_2 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_215 ();
 sg13g2_fill_1 FILLER_32_217 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_235 ();
 sg13g2_fill_2 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_283 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_293 ();
 sg13g2_decap_4 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_11 ();
 sg13g2_fill_2 FILLER_33_24 ();
 sg13g2_fill_1 FILLER_33_26 ();
 sg13g2_decap_8 FILLER_33_59 ();
 sg13g2_decap_8 FILLER_33_66 ();
 sg13g2_fill_2 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_83 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_decap_4 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_decap_8 FILLER_33_125 ();
 sg13g2_decap_4 FILLER_33_132 ();
 sg13g2_fill_2 FILLER_33_154 ();
 sg13g2_fill_1 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_195 ();
 sg13g2_fill_1 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_fill_2 FILLER_33_214 ();
 sg13g2_fill_2 FILLER_33_221 ();
 sg13g2_fill_1 FILLER_33_223 ();
 sg13g2_fill_2 FILLER_33_235 ();
 sg13g2_fill_1 FILLER_33_267 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_2 FILLER_33_376 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_2 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_36 ();
 sg13g2_fill_2 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_104 ();
 sg13g2_decap_8 FILLER_34_125 ();
 sg13g2_fill_2 FILLER_34_132 ();
 sg13g2_fill_1 FILLER_34_134 ();
 sg13g2_decap_4 FILLER_34_149 ();
 sg13g2_fill_2 FILLER_34_174 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_decap_4 FILLER_34_234 ();
 sg13g2_decap_4 FILLER_34_247 ();
 sg13g2_decap_4 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_320 ();
 sg13g2_fill_2 FILLER_34_353 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_decap_4 FILLER_34_360 ();
 sg13g2_fill_2 FILLER_34_364 ();
 sg13g2_fill_2 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_15 ();
 sg13g2_decap_8 FILLER_35_22 ();
 sg13g2_decap_4 FILLER_35_29 ();
 sg13g2_fill_2 FILLER_35_38 ();
 sg13g2_decap_8 FILLER_35_66 ();
 sg13g2_fill_1 FILLER_35_73 ();
 sg13g2_fill_2 FILLER_35_90 ();
 sg13g2_fill_2 FILLER_35_124 ();
 sg13g2_fill_2 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_fill_1 FILLER_35_194 ();
 sg13g2_fill_2 FILLER_35_200 ();
 sg13g2_fill_1 FILLER_35_202 ();
 sg13g2_fill_1 FILLER_35_207 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_fill_2 FILLER_35_260 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_fill_1 FILLER_35_290 ();
 sg13g2_decap_8 FILLER_35_295 ();
 sg13g2_decap_4 FILLER_35_306 ();
 sg13g2_fill_1 FILLER_35_310 ();
 sg13g2_decap_8 FILLER_35_319 ();
 sg13g2_fill_2 FILLER_35_326 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_349 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_fill_1 FILLER_35_376 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_fill_1 FILLER_36_46 ();
 sg13g2_fill_2 FILLER_36_61 ();
 sg13g2_fill_1 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_68 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_136 ();
 sg13g2_fill_2 FILLER_36_145 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_decap_4 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_184 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_216 ();
 sg13g2_fill_2 FILLER_36_225 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_decap_4 FILLER_36_270 ();
 sg13g2_decap_4 FILLER_36_283 ();
 sg13g2_decap_4 FILLER_36_303 ();
 sg13g2_fill_2 FILLER_36_319 ();
 sg13g2_fill_1 FILLER_36_330 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_4 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_25 ();
 sg13g2_fill_2 FILLER_37_45 ();
 sg13g2_fill_1 FILLER_37_47 ();
 sg13g2_fill_2 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_96 ();
 sg13g2_fill_2 FILLER_37_105 ();
 sg13g2_fill_2 FILLER_37_125 ();
 sg13g2_fill_2 FILLER_37_132 ();
 sg13g2_fill_2 FILLER_37_156 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_fill_1 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_292 ();
 sg13g2_decap_4 FILLER_37_320 ();
 sg13g2_fill_1 FILLER_37_324 ();
 sg13g2_fill_2 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_fill_1 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_83 ();
 sg13g2_fill_1 FILLER_38_120 ();
 sg13g2_fill_2 FILLER_38_130 ();
 sg13g2_decap_8 FILLER_38_186 ();
 sg13g2_decap_4 FILLER_38_193 ();
 sg13g2_fill_1 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_211 ();
 sg13g2_decap_4 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_232 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_decap_8 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_251 ();
 sg13g2_decap_8 FILLER_38_258 ();
 sg13g2_decap_4 FILLER_38_265 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_decap_4 FILLER_38_281 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_fill_2 FILLER_38_296 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_fill_2 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule

module tt_um_drum_goekce (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire clknet_0_clk;
 wire \a[0] ;
 wire \a[1] ;
 wire \a[2] ;
 wire \a[3] ;
 wire \a[4] ;
 wire \a[5] ;
 wire \a[6] ;
 wire \a[7] ;
 wire \b[0] ;
 wire \b[1] ;
 wire \b[2] ;
 wire \b[3] ;
 wire \b[4] ;
 wire \b[5] ;
 wire \b[6] ;
 wire \b[7] ;
 wire \ram[0][0] ;
 wire \ram[0][1] ;
 wire \ram[0][2] ;
 wire \ram[0][3] ;
 wire \ram[0][4] ;
 wire \ram[0][5] ;
 wire \ram[0][6] ;
 wire \ram[0][7] ;
 wire \ram[10][0] ;
 wire \ram[10][1] ;
 wire \ram[10][2] ;
 wire \ram[10][3] ;
 wire \ram[10][4] ;
 wire \ram[10][5] ;
 wire \ram[10][6] ;
 wire \ram[10][7] ;
 wire \ram[11][0] ;
 wire \ram[11][1] ;
 wire \ram[11][2] ;
 wire \ram[11][3] ;
 wire \ram[11][4] ;
 wire \ram[11][5] ;
 wire \ram[11][6] ;
 wire \ram[11][7] ;
 wire \ram[12][0] ;
 wire \ram[12][1] ;
 wire \ram[12][2] ;
 wire \ram[12][3] ;
 wire \ram[12][4] ;
 wire \ram[12][5] ;
 wire \ram[12][6] ;
 wire \ram[12][7] ;
 wire \ram[13][0] ;
 wire \ram[13][1] ;
 wire \ram[13][2] ;
 wire \ram[13][3] ;
 wire \ram[13][4] ;
 wire \ram[13][5] ;
 wire \ram[13][6] ;
 wire \ram[13][7] ;
 wire \ram[14][0] ;
 wire \ram[14][1] ;
 wire \ram[14][2] ;
 wire \ram[14][3] ;
 wire \ram[14][4] ;
 wire \ram[14][5] ;
 wire \ram[14][6] ;
 wire \ram[14][7] ;
 wire \ram[15][0] ;
 wire \ram[15][1] ;
 wire \ram[15][2] ;
 wire \ram[15][3] ;
 wire \ram[15][4] ;
 wire \ram[15][5] ;
 wire \ram[15][6] ;
 wire \ram[15][7] ;
 wire \ram[1][0] ;
 wire \ram[1][1] ;
 wire \ram[1][2] ;
 wire \ram[1][3] ;
 wire \ram[1][4] ;
 wire \ram[1][5] ;
 wire \ram[1][6] ;
 wire \ram[1][7] ;
 wire \ram[2][0] ;
 wire \ram[2][1] ;
 wire \ram[2][2] ;
 wire \ram[2][3] ;
 wire \ram[2][4] ;
 wire \ram[2][5] ;
 wire \ram[2][6] ;
 wire \ram[2][7] ;
 wire \ram[3][0] ;
 wire \ram[3][1] ;
 wire \ram[3][2] ;
 wire \ram[3][3] ;
 wire \ram[3][4] ;
 wire \ram[3][5] ;
 wire \ram[3][6] ;
 wire \ram[3][7] ;
 wire \ram[4][0] ;
 wire \ram[4][1] ;
 wire \ram[4][2] ;
 wire \ram[4][3] ;
 wire \ram[4][4] ;
 wire \ram[4][5] ;
 wire \ram[4][6] ;
 wire \ram[4][7] ;
 wire \ram[5][0] ;
 wire \ram[5][1] ;
 wire \ram[5][2] ;
 wire \ram[5][3] ;
 wire \ram[5][4] ;
 wire \ram[5][5] ;
 wire \ram[5][6] ;
 wire \ram[5][7] ;
 wire \ram[6][0] ;
 wire \ram[6][1] ;
 wire \ram[6][2] ;
 wire \ram[6][3] ;
 wire \ram[6][4] ;
 wire \ram[6][5] ;
 wire \ram[6][6] ;
 wire \ram[6][7] ;
 wire \ram[7][0] ;
 wire \ram[7][1] ;
 wire \ram[7][2] ;
 wire \ram[7][3] ;
 wire \ram[7][4] ;
 wire \ram[7][5] ;
 wire \ram[7][6] ;
 wire \ram[7][7] ;
 wire \result_addr[0] ;
 wire \result_addr[1] ;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;

 sg13g2_inv_1 _0953_ (.Y(_0139_),
    .A(net311));
 sg13g2_inv_1 _0954_ (.Y(_0140_),
    .A(net295));
 sg13g2_inv_1 _0955_ (.Y(_0141_),
    .A(\result_addr[1] ));
 sg13g2_inv_1 _0956_ (.Y(_0142_),
    .A(\result_addr[0] ));
 sg13g2_inv_1 _0957_ (.Y(_0143_),
    .A(\ram[5][4] ));
 sg13g2_inv_1 _0958_ (.Y(_0144_),
    .A(\ram[5][5] ));
 sg13g2_inv_1 _0959_ (.Y(_0145_),
    .A(\ram[5][7] ));
 sg13g2_inv_1 _0960_ (.Y(_0146_),
    .A(\ram[7][7] ));
 sg13g2_or2_1 _0961_ (.X(_0147_),
    .B(\a[6] ),
    .A(net288));
 sg13g2_xor2_1 _0962_ (.B(\a[6] ),
    .A(net287),
    .X(_0148_));
 sg13g2_or2_1 _0963_ (.X(_0149_),
    .B(\b[6] ),
    .A(net286));
 sg13g2_xor2_1 _0964_ (.B(\b[6] ),
    .A(net285),
    .X(_0150_));
 sg13g2_nor2_1 _0965_ (.A(_0148_),
    .B(net284),
    .Y(_0151_));
 sg13g2_or2_1 _0966_ (.X(_0152_),
    .B(net284),
    .A(_0148_));
 sg13g2_nand3_1 _0967_ (.B(\a[0] ),
    .C(\a[6] ),
    .A(net287),
    .Y(_0153_));
 sg13g2_o21ai_1 _0968_ (.B1(_0153_),
    .Y(_0154_),
    .A1(\a[0] ),
    .A2(_0147_));
 sg13g2_nand3_1 _0969_ (.B(\b[0] ),
    .C(\b[6] ),
    .A(net286),
    .Y(_0155_));
 sg13g2_o21ai_1 _0970_ (.B1(_0155_),
    .Y(_0156_),
    .A1(\b[0] ),
    .A2(_0149_));
 sg13g2_or2_1 _0971_ (.X(_0157_),
    .B(_0156_),
    .A(_0154_));
 sg13g2_nor2_1 _0972_ (.A(_0152_),
    .B(_0157_),
    .Y(_0158_));
 sg13g2_xnor2_1 _0973_ (.Y(_0159_),
    .A(net288),
    .B(net286));
 sg13g2_xor2_1 _0974_ (.B(net281),
    .A(_0158_),
    .X(_0160_));
 sg13g2_inv_1 _0975_ (.Y(uio_out[0]),
    .A(_0160_));
 sg13g2_xnor2_1 _0976_ (.Y(_0161_),
    .A(net285),
    .B(\b[2] ));
 sg13g2_xor2_1 _0977_ (.B(\b[2] ),
    .A(net285),
    .X(_0162_));
 sg13g2_o21ai_1 _0978_ (.B1(\b[1] ),
    .Y(_0163_),
    .A1(net285),
    .A2(\b[6] ));
 sg13g2_a21o_1 _0979_ (.A2(\b[6] ),
    .A1(net285),
    .B1(\b[1] ),
    .X(_0164_));
 sg13g2_a22oi_1 _0980_ (.Y(_0165_),
    .B1(_0163_),
    .B2(_0164_),
    .A2(_0162_),
    .A1(net284));
 sg13g2_xnor2_1 _0981_ (.Y(_0166_),
    .A(net287),
    .B(\a[2] ));
 sg13g2_xor2_1 _0982_ (.B(\a[2] ),
    .A(net287),
    .X(_0167_));
 sg13g2_o21ai_1 _0983_ (.B1(\a[1] ),
    .Y(_0168_),
    .A1(net287),
    .A2(\a[6] ));
 sg13g2_a21o_1 _0984_ (.A2(\a[6] ),
    .A1(net287),
    .B1(\a[1] ),
    .X(_0169_));
 sg13g2_a22oi_1 _0985_ (.Y(_0170_),
    .B1(_0168_),
    .B2(_0169_),
    .A2(_0167_),
    .A1(_0148_));
 sg13g2_or2_1 _0986_ (.X(_0171_),
    .B(_0170_),
    .A(_0165_));
 sg13g2_nor2_1 _0987_ (.A(_0154_),
    .B(_0165_),
    .Y(_0172_));
 sg13g2_nor2_1 _0988_ (.A(_0156_),
    .B(_0170_),
    .Y(_0173_));
 sg13g2_nor2_1 _0989_ (.A(_0157_),
    .B(_0171_),
    .Y(_0174_));
 sg13g2_xnor2_1 _0990_ (.Y(_0175_),
    .A(_0172_),
    .B(_0173_));
 sg13g2_and2_1 _0991_ (.A(_0148_),
    .B(net284),
    .X(_0176_));
 sg13g2_inv_1 _0992_ (.Y(_0177_),
    .A(net275));
 sg13g2_nor2_1 _0993_ (.A(net276),
    .B(net274),
    .Y(_0178_));
 sg13g2_nand2b_1 _0994_ (.Y(_0179_),
    .B(net254),
    .A_N(_0157_));
 sg13g2_o21ai_1 _0995_ (.B1(_0179_),
    .Y(_0180_),
    .A1(_0152_),
    .A2(_0175_));
 sg13g2_xor2_1 _0996_ (.B(_0180_),
    .A(net281),
    .X(_0181_));
 sg13g2_inv_2 _0997_ (.Y(uio_out[1]),
    .A(_0181_));
 sg13g2_xnor2_1 _0998_ (.Y(_0182_),
    .A(net285),
    .B(\b[3] ));
 sg13g2_mux2_2 _0999_ (.A0(_0161_),
    .A1(_0182_),
    .S(net284),
    .X(_0183_));
 sg13g2_nor2_1 _1000_ (.A(_0170_),
    .B(_0183_),
    .Y(_0184_));
 sg13g2_nand2_1 _1001_ (.Y(_0185_),
    .A(_0172_),
    .B(_0184_));
 sg13g2_o21ai_1 _1002_ (.B1(_0171_),
    .Y(_0186_),
    .A1(_0154_),
    .A2(_0183_));
 sg13g2_nand2_1 _1003_ (.Y(_0187_),
    .A(_0185_),
    .B(_0186_));
 sg13g2_xnor2_1 _1004_ (.Y(_0188_),
    .A(net287),
    .B(\a[3] ));
 sg13g2_mux2_2 _1005_ (.A0(_0166_),
    .A1(_0188_),
    .S(_0148_),
    .X(_0189_));
 sg13g2_nor2_1 _1006_ (.A(_0156_),
    .B(_0189_),
    .Y(_0190_));
 sg13g2_nor2b_1 _1007_ (.A(_0187_),
    .B_N(_0190_),
    .Y(_0191_));
 sg13g2_xnor2_1 _1008_ (.Y(_0192_),
    .A(_0187_),
    .B(_0190_));
 sg13g2_xnor2_1 _1009_ (.Y(_0193_),
    .A(_0174_),
    .B(_0192_));
 sg13g2_a22oi_1 _1010_ (.Y(_0194_),
    .B1(_0193_),
    .B2(net276),
    .A2(net254),
    .A1(_0175_));
 sg13g2_xor2_1 _1011_ (.B(_0194_),
    .A(net281),
    .X(_0195_));
 sg13g2_inv_2 _1012_ (.Y(uio_out[2]),
    .A(_0195_));
 sg13g2_xnor2_1 _1013_ (.Y(_0196_),
    .A(net285),
    .B(\b[4] ));
 sg13g2_mux2_2 _1014_ (.A0(_0182_),
    .A1(_0196_),
    .S(net284),
    .X(_0197_));
 sg13g2_xnor2_1 _1015_ (.Y(_0198_),
    .A(net288),
    .B(\a[4] ));
 sg13g2_mux2_2 _1016_ (.A0(_0188_),
    .A1(_0198_),
    .S(_0148_),
    .X(_0199_));
 sg13g2_nor2_2 _1017_ (.A(_0197_),
    .B(_0199_),
    .Y(_0200_));
 sg13g2_nor2_1 _1018_ (.A(_0154_),
    .B(_0197_),
    .Y(_0201_));
 sg13g2_nor2_1 _1019_ (.A(_0156_),
    .B(_0199_),
    .Y(_0202_));
 sg13g2_nand2_1 _1020_ (.Y(_0203_),
    .A(_0201_),
    .B(_0202_));
 sg13g2_xnor2_1 _1021_ (.Y(_0204_),
    .A(_0201_),
    .B(_0202_));
 sg13g2_or2_1 _1022_ (.X(_0205_),
    .B(_0189_),
    .A(_0183_));
 sg13g2_or2_1 _1023_ (.X(_0206_),
    .B(_0189_),
    .A(_0165_));
 sg13g2_nor2_1 _1024_ (.A(_0171_),
    .B(_0205_),
    .Y(_0207_));
 sg13g2_nor2b_1 _1025_ (.A(_0184_),
    .B_N(_0206_),
    .Y(_0208_));
 sg13g2_nand3_1 _1026_ (.B(_0184_),
    .C(_0206_),
    .A(_0172_),
    .Y(_0209_));
 sg13g2_o21ai_1 _1027_ (.B1(_0185_),
    .Y(_0210_),
    .A1(_0207_),
    .A2(_0208_));
 sg13g2_nand2_1 _1028_ (.Y(_0211_),
    .A(_0209_),
    .B(_0210_));
 sg13g2_xnor2_1 _1029_ (.Y(_0212_),
    .A(_0204_),
    .B(_0211_));
 sg13g2_a21oi_1 _1030_ (.A1(_0174_),
    .A2(_0192_),
    .Y(_0213_),
    .B1(_0191_));
 sg13g2_nor2_1 _1031_ (.A(_0212_),
    .B(_0213_),
    .Y(_0214_));
 sg13g2_xnor2_1 _1032_ (.Y(_0215_),
    .A(_0212_),
    .B(_0213_));
 sg13g2_and2_1 _1033_ (.A(net254),
    .B(_0193_),
    .X(_0216_));
 sg13g2_a221oi_1 _1034_ (.B2(net276),
    .C1(_0216_),
    .B1(_0215_),
    .A1(_0175_),
    .Y(_0217_),
    .A2(net274));
 sg13g2_xor2_1 _1035_ (.B(_0217_),
    .A(net283),
    .X(_0218_));
 sg13g2_inv_2 _1036_ (.Y(uio_out[3]),
    .A(_0218_));
 sg13g2_o21ai_1 _1037_ (.B1(_0209_),
    .Y(_0219_),
    .A1(_0204_),
    .A2(_0211_));
 sg13g2_nor2_1 _1038_ (.A(_0183_),
    .B(_0199_),
    .Y(_0220_));
 sg13g2_nor2_1 _1039_ (.A(_0165_),
    .B(_0199_),
    .Y(_0221_));
 sg13g2_nor2b_1 _1040_ (.A(_0206_),
    .B_N(_0220_),
    .Y(_0222_));
 sg13g2_xnor2_1 _1041_ (.Y(_0223_),
    .A(_0205_),
    .B(_0221_));
 sg13g2_xnor2_1 _1042_ (.Y(_0224_),
    .A(_0207_),
    .B(_0223_));
 sg13g2_xnor2_1 _1043_ (.Y(_0225_),
    .A(net288),
    .B(\a[5] ));
 sg13g2_mux2_2 _1044_ (.A0(_0198_),
    .A1(_0225_),
    .S(_0148_),
    .X(_0226_));
 sg13g2_nor2_1 _1045_ (.A(_0156_),
    .B(_0226_),
    .Y(_0227_));
 sg13g2_xnor2_1 _1046_ (.Y(_0228_),
    .A(net286),
    .B(\b[5] ));
 sg13g2_mux2_2 _1047_ (.A0(_0196_),
    .A1(_0228_),
    .S(_0150_),
    .X(_0229_));
 sg13g2_nor2_1 _1048_ (.A(_0170_),
    .B(_0229_),
    .Y(_0230_));
 sg13g2_nor2_1 _1049_ (.A(_0154_),
    .B(_0229_),
    .Y(_0231_));
 sg13g2_nor2_1 _1050_ (.A(_0170_),
    .B(_0197_),
    .Y(_0232_));
 sg13g2_xor2_1 _1051_ (.B(_0232_),
    .A(_0231_),
    .X(_0233_));
 sg13g2_xnor2_1 _1052_ (.Y(_0234_),
    .A(_0227_),
    .B(_0233_));
 sg13g2_nor2_1 _1053_ (.A(_0224_),
    .B(_0234_),
    .Y(_0235_));
 sg13g2_xor2_1 _1054_ (.B(_0234_),
    .A(_0224_),
    .X(_0236_));
 sg13g2_nand2_1 _1055_ (.Y(_0237_),
    .A(_0219_),
    .B(_0236_));
 sg13g2_xnor2_1 _1056_ (.Y(_0238_),
    .A(_0219_),
    .B(_0236_));
 sg13g2_xor2_1 _1057_ (.B(_0238_),
    .A(_0203_),
    .X(_0239_));
 sg13g2_and2_1 _1058_ (.A(_0214_),
    .B(_0239_),
    .X(_0240_));
 sg13g2_xnor2_1 _1059_ (.Y(_0241_),
    .A(_0214_),
    .B(_0239_));
 sg13g2_and2_1 _1060_ (.A(net255),
    .B(_0215_),
    .X(_0242_));
 sg13g2_a221oi_1 _1061_ (.B2(net276),
    .C1(_0242_),
    .B1(_0241_),
    .A1(net274),
    .Y(_0243_),
    .A2(_0193_));
 sg13g2_xor2_1 _1062_ (.B(_0243_),
    .A(net283),
    .X(_0244_));
 sg13g2_inv_1 _1063_ (.Y(uio_out[4]),
    .A(_0244_));
 sg13g2_o21ai_1 _1064_ (.B1(_0237_),
    .Y(_0245_),
    .A1(_0203_),
    .A2(_0238_));
 sg13g2_a22oi_1 _1065_ (.Y(_0246_),
    .B1(_0233_),
    .B2(_0227_),
    .A2(_0230_),
    .A1(_0201_));
 sg13g2_a21oi_1 _1066_ (.A1(_0207_),
    .A2(_0223_),
    .Y(_0247_),
    .B1(_0235_));
 sg13g2_nor2b_2 _1067_ (.A(_0148_),
    .B_N(_0225_),
    .Y(_0248_));
 sg13g2_or2_1 _1068_ (.X(_0249_),
    .B(_0248_),
    .A(_0156_));
 sg13g2_nor2_1 _1069_ (.A(_0189_),
    .B(_0229_),
    .Y(_0250_));
 sg13g2_nor2_1 _1070_ (.A(_0189_),
    .B(_0197_),
    .Y(_0251_));
 sg13g2_nand2_1 _1071_ (.Y(_0252_),
    .A(_0232_),
    .B(_0250_));
 sg13g2_xnor2_1 _1072_ (.Y(_0253_),
    .A(_0230_),
    .B(_0251_));
 sg13g2_xor2_1 _1073_ (.B(_0253_),
    .A(_0249_),
    .X(_0254_));
 sg13g2_nor2b_2 _1074_ (.A(net284),
    .B_N(_0228_),
    .Y(_0255_));
 sg13g2_nand2b_1 _1075_ (.Y(_0256_),
    .B(_0228_),
    .A_N(net284));
 sg13g2_nor2_1 _1076_ (.A(_0154_),
    .B(_0255_),
    .Y(_0257_));
 sg13g2_nor2_1 _1077_ (.A(_0183_),
    .B(_0226_),
    .Y(_0258_));
 sg13g2_nor2_1 _1078_ (.A(_0165_),
    .B(_0226_),
    .Y(_0259_));
 sg13g2_and2_1 _1079_ (.A(_0220_),
    .B(_0259_),
    .X(_0260_));
 sg13g2_xor2_1 _1080_ (.B(_0259_),
    .A(_0220_),
    .X(_0261_));
 sg13g2_xor2_1 _1081_ (.B(_0261_),
    .A(_0257_),
    .X(_0262_));
 sg13g2_and2_1 _1082_ (.A(_0222_),
    .B(_0262_),
    .X(_0263_));
 sg13g2_xor2_1 _1083_ (.B(_0262_),
    .A(_0222_),
    .X(_0264_));
 sg13g2_xnor2_1 _1084_ (.Y(_0265_),
    .A(_0254_),
    .B(_0264_));
 sg13g2_nor2_1 _1085_ (.A(_0247_),
    .B(_0265_),
    .Y(_0266_));
 sg13g2_xnor2_1 _1086_ (.Y(_0267_),
    .A(_0247_),
    .B(_0265_));
 sg13g2_nor2_1 _1087_ (.A(_0246_),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_xor2_1 _1088_ (.B(_0267_),
    .A(_0246_),
    .X(_0269_));
 sg13g2_and2_1 _1089_ (.A(_0245_),
    .B(_0269_),
    .X(_0270_));
 sg13g2_xor2_1 _1090_ (.B(_0269_),
    .A(_0245_),
    .X(_0271_));
 sg13g2_xnor2_1 _1091_ (.Y(_0272_),
    .A(_0240_),
    .B(_0271_));
 sg13g2_and2_1 _1092_ (.A(net275),
    .B(_0215_),
    .X(_0273_));
 sg13g2_a221oi_1 _1093_ (.B2(_0151_),
    .C1(_0273_),
    .B1(_0272_),
    .A1(net255),
    .Y(_0274_),
    .A2(_0241_));
 sg13g2_xor2_1 _1094_ (.B(_0274_),
    .A(net283),
    .X(_0275_));
 sg13g2_inv_2 _1095_ (.Y(uio_out[5]),
    .A(_0275_));
 sg13g2_a21oi_1 _1096_ (.A1(_0240_),
    .A2(_0271_),
    .Y(_0276_),
    .B1(_0270_));
 sg13g2_nor2_1 _1097_ (.A(_0266_),
    .B(_0268_),
    .Y(_0277_));
 sg13g2_o21ai_1 _1098_ (.B1(_0252_),
    .Y(_0278_),
    .A1(_0249_),
    .A2(_0253_));
 sg13g2_a21oi_1 _1099_ (.A1(_0254_),
    .A2(_0264_),
    .Y(_0279_),
    .B1(_0263_));
 sg13g2_nand2_1 _1100_ (.Y(_0280_),
    .A(_0200_),
    .B(_0250_));
 sg13g2_xnor2_1 _1101_ (.Y(_0281_),
    .A(_0200_),
    .B(_0250_));
 sg13g2_a21o_1 _1102_ (.A2(_0261_),
    .A1(_0257_),
    .B1(_0260_),
    .X(_0282_));
 sg13g2_nor2_1 _1103_ (.A(_0170_),
    .B(_0255_),
    .Y(_0283_));
 sg13g2_nor2_1 _1104_ (.A(_0183_),
    .B(_0248_),
    .Y(_0284_));
 sg13g2_nor2_1 _1105_ (.A(_0165_),
    .B(_0248_),
    .Y(_0285_));
 sg13g2_xor2_1 _1106_ (.B(_0285_),
    .A(_0258_),
    .X(_0286_));
 sg13g2_xor2_1 _1107_ (.B(_0286_),
    .A(_0283_),
    .X(_0287_));
 sg13g2_nand2_1 _1108_ (.Y(_0288_),
    .A(_0282_),
    .B(_0287_));
 sg13g2_xnor2_1 _1109_ (.Y(_0289_),
    .A(_0282_),
    .B(_0287_));
 sg13g2_xnor2_1 _1110_ (.Y(_0290_),
    .A(_0281_),
    .B(_0289_));
 sg13g2_nor2_1 _1111_ (.A(_0279_),
    .B(_0290_),
    .Y(_0291_));
 sg13g2_xor2_1 _1112_ (.B(_0290_),
    .A(_0279_),
    .X(_0292_));
 sg13g2_xnor2_1 _1113_ (.Y(_0293_),
    .A(_0278_),
    .B(_0292_));
 sg13g2_or2_1 _1114_ (.X(_0294_),
    .B(_0293_),
    .A(_0277_));
 sg13g2_xnor2_1 _1115_ (.Y(_0295_),
    .A(_0277_),
    .B(_0293_));
 sg13g2_xnor2_1 _1116_ (.Y(_0296_),
    .A(_0276_),
    .B(_0295_));
 sg13g2_and2_1 _1117_ (.A(net274),
    .B(_0241_),
    .X(_0297_));
 sg13g2_a221oi_1 _1118_ (.B2(_0151_),
    .C1(_0297_),
    .B1(_0296_),
    .A1(net255),
    .Y(_0298_),
    .A2(_0272_));
 sg13g2_xor2_1 _1119_ (.B(_0298_),
    .A(net282),
    .X(_0299_));
 sg13g2_inv_1 _1120_ (.Y(uio_out[6]),
    .A(_0299_));
 sg13g2_o21ai_1 _1121_ (.B1(_0294_),
    .Y(_0300_),
    .A1(_0276_),
    .A2(_0295_));
 sg13g2_a21oi_1 _1122_ (.A1(_0278_),
    .A2(_0292_),
    .Y(_0301_),
    .B1(_0291_));
 sg13g2_o21ai_1 _1123_ (.B1(_0288_),
    .Y(_0302_),
    .A1(_0281_),
    .A2(_0289_));
 sg13g2_nand2b_1 _1124_ (.Y(_0303_),
    .B(_0256_),
    .A_N(_0248_));
 sg13g2_nor2_1 _1125_ (.A(_0189_),
    .B(_0255_),
    .Y(_0304_));
 sg13g2_nand2_1 _1126_ (.Y(_0305_),
    .A(_0284_),
    .B(_0304_));
 sg13g2_xnor2_1 _1127_ (.Y(_0306_),
    .A(_0284_),
    .B(_0304_));
 sg13g2_a22oi_1 _1128_ (.Y(_0307_),
    .B1(_0286_),
    .B2(_0283_),
    .A2(_0284_),
    .A1(_0259_));
 sg13g2_nor2_1 _1129_ (.A(_0306_),
    .B(_0307_),
    .Y(_0308_));
 sg13g2_xnor2_1 _1130_ (.Y(_0309_),
    .A(_0306_),
    .B(_0307_));
 sg13g2_inv_1 _1131_ (.Y(_0310_),
    .A(_0309_));
 sg13g2_nor2_2 _1132_ (.A(_0226_),
    .B(_0229_),
    .Y(_0311_));
 sg13g2_or2_1 _1133_ (.X(_0312_),
    .B(_0226_),
    .A(_0197_));
 sg13g2_nand2_2 _1134_ (.Y(_0313_),
    .A(_0200_),
    .B(_0311_));
 sg13g2_inv_1 _1135_ (.Y(_0314_),
    .A(_0313_));
 sg13g2_o21ai_1 _1136_ (.B1(_0312_),
    .Y(_0315_),
    .A1(_0199_),
    .A2(_0229_));
 sg13g2_and2_1 _1137_ (.A(_0313_),
    .B(_0315_),
    .X(_0316_));
 sg13g2_xnor2_1 _1138_ (.Y(_0317_),
    .A(_0309_),
    .B(_0316_));
 sg13g2_nand2_1 _1139_ (.Y(_0318_),
    .A(_0302_),
    .B(_0317_));
 sg13g2_xnor2_1 _1140_ (.Y(_0319_),
    .A(_0302_),
    .B(_0317_));
 sg13g2_xnor2_1 _1141_ (.Y(_0320_),
    .A(_0280_),
    .B(_0319_));
 sg13g2_nor2_1 _1142_ (.A(_0301_),
    .B(_0320_),
    .Y(_0321_));
 sg13g2_xor2_1 _1143_ (.B(_0320_),
    .A(_0301_),
    .X(_0322_));
 sg13g2_xnor2_1 _1144_ (.Y(_0323_),
    .A(_0300_),
    .B(_0322_));
 sg13g2_and2_1 _1145_ (.A(net274),
    .B(_0272_),
    .X(_0324_));
 sg13g2_a221oi_1 _1146_ (.B2(net276),
    .C1(_0324_),
    .B1(_0323_),
    .A1(net255),
    .Y(_0325_),
    .A2(_0296_));
 sg13g2_xor2_1 _1147_ (.B(_0325_),
    .A(net281),
    .X(_0326_));
 sg13g2_inv_1 _1148_ (.Y(uio_out[7]),
    .A(_0326_));
 sg13g2_nand2_1 _1149_ (.Y(_0327_),
    .A(net293),
    .B(net4));
 sg13g2_and3_1 _1150_ (.X(_0328_),
    .A(net293),
    .B(net4),
    .C(net321));
 sg13g2_inv_1 _1151_ (.Y(_0329_),
    .A(net289));
 sg13g2_nand2_1 _1152_ (.Y(_0330_),
    .A(net302),
    .B(net289));
 sg13g2_nand4_1 _1153_ (.B(net305),
    .C(net296),
    .A(net313),
    .Y(_0331_),
    .D(net289));
 sg13g2_nand2_2 _1154_ (.Y(_0332_),
    .A(net5),
    .B(net290));
 sg13g2_nand2_1 _1155_ (.Y(_0333_),
    .A(net215),
    .B(net279));
 sg13g2_o21ai_1 _1156_ (.B1(_0333_),
    .Y(_0001_),
    .A1(net279),
    .A2(_0332_));
 sg13g2_nand2_2 _1157_ (.Y(_0334_),
    .A(net6),
    .B(net290));
 sg13g2_nand2_1 _1158_ (.Y(_0335_),
    .A(net207),
    .B(net279));
 sg13g2_o21ai_1 _1159_ (.B1(_0335_),
    .Y(_0002_),
    .A1(net279),
    .A2(_0334_));
 sg13g2_nand2_2 _1160_ (.Y(_0336_),
    .A(net7),
    .B(net290));
 sg13g2_nand2_1 _1161_ (.Y(_0337_),
    .A(net182),
    .B(_0331_));
 sg13g2_o21ai_1 _1162_ (.B1(_0337_),
    .Y(_0003_),
    .A1(net279),
    .A2(_0336_));
 sg13g2_nand2_2 _1163_ (.Y(_0338_),
    .A(net8),
    .B(net290));
 sg13g2_nand2_1 _1164_ (.Y(_0339_),
    .A(net223),
    .B(net279));
 sg13g2_o21ai_1 _1165_ (.B1(_0339_),
    .Y(_0004_),
    .A1(net279),
    .A2(_0338_));
 sg13g2_nand2_2 _1166_ (.Y(_0340_),
    .A(net9),
    .B(net290));
 sg13g2_nand2_1 _1167_ (.Y(_0341_),
    .A(net222),
    .B(net280));
 sg13g2_o21ai_1 _1168_ (.B1(_0341_),
    .Y(_0005_),
    .A1(net280),
    .A2(_0340_));
 sg13g2_nand2_2 _1169_ (.Y(_0342_),
    .A(net10),
    .B(net289));
 sg13g2_nand2_1 _1170_ (.Y(_0343_),
    .A(net231),
    .B(net280));
 sg13g2_o21ai_1 _1171_ (.B1(_0343_),
    .Y(_0006_),
    .A1(net280),
    .A2(_0342_));
 sg13g2_nand2_2 _1172_ (.Y(_0344_),
    .A(net11),
    .B(net289));
 sg13g2_nand2_1 _1173_ (.Y(_0345_),
    .A(net218),
    .B(net279));
 sg13g2_o21ai_1 _1174_ (.B1(_0345_),
    .Y(_0007_),
    .A1(net280),
    .A2(_0344_));
 sg13g2_nand2_2 _1175_ (.Y(_0346_),
    .A(net12),
    .B(net289));
 sg13g2_nand2_1 _1176_ (.Y(_0347_),
    .A(net238),
    .B(net280));
 sg13g2_o21ai_1 _1177_ (.B1(_0347_),
    .Y(_0008_),
    .A1(net280),
    .A2(_0346_));
 sg13g2_and2_1 _1178_ (.A(net320),
    .B(net151),
    .X(_0009_));
 sg13g2_xor2_1 _1179_ (.B(net358),
    .A(\result_addr[1] ),
    .X(_0348_));
 sg13g2_and2_1 _1180_ (.A(net320),
    .B(net359),
    .X(_0010_));
 sg13g2_nand4_1 _1181_ (.B(_0141_),
    .C(_0142_),
    .A(net319),
    .Y(_0349_),
    .D(net3));
 sg13g2_and2_1 _1182_ (.A(net319),
    .B(net272),
    .X(_0350_));
 sg13g2_nand2_1 _1183_ (.Y(_0351_),
    .A(net178),
    .B(net253));
 sg13g2_o21ai_1 _1184_ (.B1(_0351_),
    .Y(_0011_),
    .A1(_0160_),
    .A2(net272));
 sg13g2_nand2_1 _1185_ (.Y(_0352_),
    .A(net153),
    .B(net252));
 sg13g2_o21ai_1 _1186_ (.B1(_0352_),
    .Y(_0012_),
    .A1(_0181_),
    .A2(net273));
 sg13g2_nand2_1 _1187_ (.Y(_0353_),
    .A(net328),
    .B(net252));
 sg13g2_o21ai_1 _1188_ (.B1(_0353_),
    .Y(_0013_),
    .A1(_0195_),
    .A2(net273));
 sg13g2_nand2_1 _1189_ (.Y(_0354_),
    .A(net156),
    .B(net252));
 sg13g2_o21ai_1 _1190_ (.B1(_0354_),
    .Y(_0014_),
    .A1(_0218_),
    .A2(net273));
 sg13g2_nand2_1 _1191_ (.Y(_0355_),
    .A(net175),
    .B(net252));
 sg13g2_o21ai_1 _1192_ (.B1(_0355_),
    .Y(_0015_),
    .A1(_0244_),
    .A2(net273));
 sg13g2_nand2_1 _1193_ (.Y(_0356_),
    .A(net154),
    .B(net253));
 sg13g2_o21ai_1 _1194_ (.B1(_0356_),
    .Y(_0016_),
    .A1(_0275_),
    .A2(net272));
 sg13g2_nand2_1 _1195_ (.Y(_0357_),
    .A(net183),
    .B(net253));
 sg13g2_o21ai_1 _1196_ (.B1(_0357_),
    .Y(_0017_),
    .A1(_0299_),
    .A2(net272));
 sg13g2_nand2_1 _1197_ (.Y(_0358_),
    .A(net160),
    .B(net253));
 sg13g2_o21ai_1 _1198_ (.B1(_0358_),
    .Y(_0018_),
    .A1(_0326_),
    .A2(_0349_));
 sg13g2_a21oi_1 _1199_ (.A1(_0300_),
    .A2(_0322_),
    .Y(_0359_),
    .B1(_0321_));
 sg13g2_o21ai_1 _1200_ (.B1(_0318_),
    .Y(_0360_),
    .A1(_0280_),
    .A2(_0319_));
 sg13g2_a21oi_2 _1201_ (.B1(_0308_),
    .Y(_0361_),
    .A2(_0316_),
    .A1(_0310_));
 sg13g2_nand2b_1 _1202_ (.Y(_0362_),
    .B(_0256_),
    .A_N(_0199_));
 sg13g2_nor2_1 _1203_ (.A(_0199_),
    .B(_0305_),
    .Y(_0363_));
 sg13g2_a21oi_1 _1204_ (.A1(_0305_),
    .A2(_0362_),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_nor2_1 _1205_ (.A(_0229_),
    .B(_0248_),
    .Y(_0365_));
 sg13g2_nor2_1 _1206_ (.A(_0197_),
    .B(_0248_),
    .Y(_0366_));
 sg13g2_and2_1 _1207_ (.A(_0311_),
    .B(_0366_),
    .X(_0367_));
 sg13g2_xor2_1 _1208_ (.B(_0366_),
    .A(_0311_),
    .X(_0368_));
 sg13g2_xnor2_1 _1209_ (.Y(_0369_),
    .A(_0364_),
    .B(_0368_));
 sg13g2_nor2_1 _1210_ (.A(_0361_),
    .B(_0369_),
    .Y(_0370_));
 sg13g2_xor2_1 _1211_ (.B(_0369_),
    .A(_0361_),
    .X(_0371_));
 sg13g2_xnor2_1 _1212_ (.Y(_0372_),
    .A(_0313_),
    .B(_0371_));
 sg13g2_nand2_1 _1213_ (.Y(_0373_),
    .A(_0360_),
    .B(_0372_));
 sg13g2_xnor2_1 _1214_ (.Y(_0374_),
    .A(_0360_),
    .B(_0372_));
 sg13g2_xnor2_1 _1215_ (.Y(_0375_),
    .A(_0359_),
    .B(_0374_));
 sg13g2_and2_1 _1216_ (.A(net254),
    .B(_0323_),
    .X(_0376_));
 sg13g2_a221oi_1 _1217_ (.B2(net276),
    .C1(_0376_),
    .B1(_0375_),
    .A1(net274),
    .Y(_0377_),
    .A2(_0296_));
 sg13g2_xor2_1 _1218_ (.B(_0377_),
    .A(net283),
    .X(_0378_));
 sg13g2_nand2_1 _1219_ (.Y(_0379_),
    .A(net210),
    .B(net253));
 sg13g2_o21ai_1 _1220_ (.B1(_0379_),
    .Y(_0019_),
    .A1(net272),
    .A2(_0378_));
 sg13g2_o21ai_1 _1221_ (.B1(_0373_),
    .Y(_0380_),
    .A1(_0359_),
    .A2(_0374_));
 sg13g2_a21oi_1 _1222_ (.A1(_0314_),
    .A2(_0371_),
    .Y(_0381_),
    .B1(_0370_));
 sg13g2_nor2_1 _1223_ (.A(_0226_),
    .B(_0255_),
    .Y(_0382_));
 sg13g2_xnor2_1 _1224_ (.Y(_0383_),
    .A(_0365_),
    .B(_0382_));
 sg13g2_a21oi_1 _1225_ (.A1(_0364_),
    .A2(_0368_),
    .Y(_0384_),
    .B1(_0363_));
 sg13g2_xor2_1 _1226_ (.B(_0384_),
    .A(_0383_),
    .X(_0385_));
 sg13g2_nand2_1 _1227_ (.Y(_0386_),
    .A(_0367_),
    .B(_0385_));
 sg13g2_xnor2_1 _1228_ (.Y(_0387_),
    .A(_0367_),
    .B(_0385_));
 sg13g2_nor2_1 _1229_ (.A(_0381_),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_xor2_1 _1230_ (.B(_0387_),
    .A(_0381_),
    .X(_0389_));
 sg13g2_xnor2_1 _1231_ (.Y(_0390_),
    .A(_0380_),
    .B(_0389_));
 sg13g2_and2_1 _1232_ (.A(net254),
    .B(_0375_),
    .X(_0391_));
 sg13g2_a221oi_1 _1233_ (.B2(net276),
    .C1(_0391_),
    .B1(_0390_),
    .A1(net274),
    .Y(_0392_),
    .A2(_0323_));
 sg13g2_xor2_1 _1234_ (.B(_0392_),
    .A(net281),
    .X(_0393_));
 sg13g2_nand2_1 _1235_ (.Y(_0394_),
    .A(net221),
    .B(net252));
 sg13g2_o21ai_1 _1236_ (.B1(_0394_),
    .Y(_0020_),
    .A1(net273),
    .A2(_0393_));
 sg13g2_a21oi_1 _1237_ (.A1(_0380_),
    .A2(_0389_),
    .Y(_0395_),
    .B1(_0388_));
 sg13g2_nor2_1 _1238_ (.A(_0303_),
    .B(_0311_),
    .Y(_0396_));
 sg13g2_o21ai_1 _1239_ (.B1(_0386_),
    .Y(_0397_),
    .A1(_0383_),
    .A2(_0384_));
 sg13g2_xnor2_1 _1240_ (.Y(_0398_),
    .A(_0396_),
    .B(_0397_));
 sg13g2_xor2_1 _1241_ (.B(_0398_),
    .A(_0395_),
    .X(_0399_));
 sg13g2_a22oi_1 _1242_ (.Y(_0400_),
    .B1(_0390_),
    .B2(net254),
    .A2(_0375_),
    .A1(net274));
 sg13g2_o21ai_1 _1243_ (.B1(_0400_),
    .Y(_0401_),
    .A1(_0152_),
    .A2(_0399_));
 sg13g2_xnor2_1 _1244_ (.Y(_0402_),
    .A(net283),
    .B(_0401_));
 sg13g2_nand2_1 _1245_ (.Y(_0403_),
    .A(net230),
    .B(net252));
 sg13g2_o21ai_1 _1246_ (.B1(_0403_),
    .Y(_0021_),
    .A1(net273),
    .A2(_0402_));
 sg13g2_a22oi_1 _1247_ (.Y(_0404_),
    .B1(_0396_),
    .B2(_0397_),
    .A2(_0382_),
    .A1(_0365_));
 sg13g2_o21ai_1 _1248_ (.B1(_0404_),
    .Y(_0405_),
    .A1(_0395_),
    .A2(_0398_));
 sg13g2_nor2_1 _1249_ (.A(_0177_),
    .B(_0390_),
    .Y(_0406_));
 sg13g2_a221oi_1 _1250_ (.B2(net276),
    .C1(_0406_),
    .B1(_0405_),
    .A1(net254),
    .Y(_0407_),
    .A2(_0399_));
 sg13g2_xnor2_1 _1251_ (.Y(_0408_),
    .A(net281),
    .B(_0407_));
 sg13g2_nand2_1 _1252_ (.Y(_0409_),
    .A(net172),
    .B(net252));
 sg13g2_o21ai_1 _1253_ (.B1(_0409_),
    .Y(_0022_),
    .A1(net273),
    .A2(_0408_));
 sg13g2_a22oi_1 _1254_ (.Y(_0410_),
    .B1(_0405_),
    .B2(net254),
    .A2(_0399_),
    .A1(net275));
 sg13g2_xnor2_1 _1255_ (.Y(_0411_),
    .A(net281),
    .B(_0410_));
 sg13g2_nand2_1 _1256_ (.Y(_0412_),
    .A(net181),
    .B(net252));
 sg13g2_o21ai_1 _1257_ (.B1(_0412_),
    .Y(_0023_),
    .A1(net273),
    .A2(_0411_));
 sg13g2_nand2_1 _1258_ (.Y(_0413_),
    .A(net275),
    .B(_0405_));
 sg13g2_xnor2_1 _1259_ (.Y(_0414_),
    .A(net281),
    .B(_0413_));
 sg13g2_nand2_1 _1260_ (.Y(_0415_),
    .A(net224),
    .B(net253));
 sg13g2_o21ai_1 _1261_ (.B1(_0415_),
    .Y(_0024_),
    .A1(net272),
    .A2(_0414_));
 sg13g2_nand2_1 _1262_ (.Y(_0416_),
    .A(net232),
    .B(net253));
 sg13g2_o21ai_1 _1263_ (.B1(_0416_),
    .Y(_0025_),
    .A1(net282),
    .A2(net272));
 sg13g2_nand2_1 _1264_ (.Y(_0417_),
    .A(net196),
    .B(net253));
 sg13g2_o21ai_1 _1265_ (.B1(_0417_),
    .Y(_0026_),
    .A1(net282),
    .A2(net272));
 sg13g2_nand4_1 _1266_ (.B(\result_addr[1] ),
    .C(_0142_),
    .A(net319),
    .Y(_0418_),
    .D(net3));
 sg13g2_and2_1 _1267_ (.A(net319),
    .B(_0418_),
    .X(_0419_));
 sg13g2_nand2_1 _1268_ (.Y(_0420_),
    .A(net158),
    .B(net250));
 sg13g2_o21ai_1 _1269_ (.B1(_0420_),
    .Y(_0027_),
    .A1(_0378_),
    .A2(net270));
 sg13g2_nand2_1 _1270_ (.Y(_0421_),
    .A(net185),
    .B(net251));
 sg13g2_o21ai_1 _1271_ (.B1(_0421_),
    .Y(_0028_),
    .A1(_0393_),
    .A2(net271));
 sg13g2_nand2_1 _1272_ (.Y(_0422_),
    .A(net167),
    .B(net251));
 sg13g2_o21ai_1 _1273_ (.B1(_0422_),
    .Y(_0029_),
    .A1(_0402_),
    .A2(net271));
 sg13g2_nand2_1 _1274_ (.Y(_0423_),
    .A(net203),
    .B(net251));
 sg13g2_o21ai_1 _1275_ (.B1(_0423_),
    .Y(_0030_),
    .A1(_0408_),
    .A2(net271));
 sg13g2_nand2_1 _1276_ (.Y(_0424_),
    .A(net216),
    .B(net251));
 sg13g2_o21ai_1 _1277_ (.B1(_0424_),
    .Y(_0031_),
    .A1(_0411_),
    .A2(net271));
 sg13g2_nand2_1 _1278_ (.Y(_0425_),
    .A(net219),
    .B(net250));
 sg13g2_o21ai_1 _1279_ (.B1(_0425_),
    .Y(_0032_),
    .A1(_0414_),
    .A2(net270));
 sg13g2_nand2_1 _1280_ (.Y(_0426_),
    .A(net194),
    .B(net250));
 sg13g2_o21ai_1 _1281_ (.B1(_0426_),
    .Y(_0033_),
    .A1(net282),
    .A2(net270));
 sg13g2_nand2_1 _1282_ (.Y(_0427_),
    .A(net201),
    .B(_0419_));
 sg13g2_o21ai_1 _1283_ (.B1(_0427_),
    .Y(_0034_),
    .A1(net282),
    .A2(net270));
 sg13g2_nor3_1 _1284_ (.A(net313),
    .B(_0140_),
    .C(_0330_),
    .Y(_0428_));
 sg13g2_nor2_1 _1285_ (.A(net329),
    .B(net268),
    .Y(_0429_));
 sg13g2_a21oi_1 _1286_ (.A1(_0332_),
    .A2(net268),
    .Y(_0035_),
    .B1(_0429_));
 sg13g2_nor2_1 _1287_ (.A(net220),
    .B(net268),
    .Y(_0430_));
 sg13g2_a21oi_1 _1288_ (.A1(_0334_),
    .A2(net268),
    .Y(_0036_),
    .B1(_0430_));
 sg13g2_nor2_1 _1289_ (.A(net227),
    .B(net269),
    .Y(_0431_));
 sg13g2_a21oi_1 _1290_ (.A1(_0336_),
    .A2(_0428_),
    .Y(_0037_),
    .B1(_0431_));
 sg13g2_nor2_1 _1291_ (.A(net217),
    .B(net268),
    .Y(_0432_));
 sg13g2_a21oi_1 _1292_ (.A1(_0338_),
    .A2(net268),
    .Y(_0038_),
    .B1(_0432_));
 sg13g2_nor2_1 _1293_ (.A(net188),
    .B(net269),
    .Y(_0433_));
 sg13g2_a21oi_1 _1294_ (.A1(_0340_),
    .A2(net269),
    .Y(_0039_),
    .B1(_0433_));
 sg13g2_nor2_1 _1295_ (.A(net212),
    .B(net269),
    .Y(_0434_));
 sg13g2_a21oi_1 _1296_ (.A1(_0342_),
    .A2(net269),
    .Y(_0040_),
    .B1(_0434_));
 sg13g2_nor2_1 _1297_ (.A(net327),
    .B(net268),
    .Y(_0435_));
 sg13g2_a21oi_1 _1298_ (.A1(_0344_),
    .A2(net268),
    .Y(_0041_),
    .B1(_0435_));
 sg13g2_nor2_1 _1299_ (.A(net326),
    .B(net269),
    .Y(_0436_));
 sg13g2_a21oi_1 _1300_ (.A1(_0346_),
    .A2(net269),
    .Y(_0042_),
    .B1(_0436_));
 sg13g2_nand2_1 _1301_ (.Y(_0437_),
    .A(net173),
    .B(net250));
 sg13g2_o21ai_1 _1302_ (.B1(_0437_),
    .Y(_0043_),
    .A1(_0160_),
    .A2(net270));
 sg13g2_nand2_1 _1303_ (.Y(_0438_),
    .A(net164),
    .B(net251));
 sg13g2_o21ai_1 _1304_ (.B1(_0438_),
    .Y(_0044_),
    .A1(_0181_),
    .A2(net271));
 sg13g2_nand2_1 _1305_ (.Y(_0439_),
    .A(net189),
    .B(net251));
 sg13g2_o21ai_1 _1306_ (.B1(_0439_),
    .Y(_0045_),
    .A1(_0195_),
    .A2(net271));
 sg13g2_nand2_1 _1307_ (.Y(_0440_),
    .A(net228),
    .B(net251));
 sg13g2_o21ai_1 _1308_ (.B1(_0440_),
    .Y(_0046_),
    .A1(_0218_),
    .A2(net271));
 sg13g2_nand2_1 _1309_ (.Y(_0441_),
    .A(net235),
    .B(net250));
 sg13g2_o21ai_1 _1310_ (.B1(_0441_),
    .Y(_0047_),
    .A1(_0244_),
    .A2(net270));
 sg13g2_nand2_1 _1311_ (.Y(_0442_),
    .A(net174),
    .B(net250));
 sg13g2_o21ai_1 _1312_ (.B1(_0442_),
    .Y(_0048_),
    .A1(_0275_),
    .A2(net270));
 sg13g2_nand2_1 _1313_ (.Y(_0443_),
    .A(net186),
    .B(net250));
 sg13g2_o21ai_1 _1314_ (.B1(_0443_),
    .Y(_0049_),
    .A1(_0299_),
    .A2(net270));
 sg13g2_nand2_1 _1315_ (.Y(_0444_),
    .A(net179),
    .B(net250));
 sg13g2_o21ai_1 _1316_ (.B1(_0444_),
    .Y(_0050_),
    .A1(_0326_),
    .A2(_0418_));
 sg13g2_nor3_1 _1317_ (.A(net313),
    .B(net296),
    .C(_0330_),
    .Y(_0445_));
 sg13g2_nor2_1 _1318_ (.A(net234),
    .B(net266),
    .Y(_0446_));
 sg13g2_a21oi_1 _1319_ (.A1(_0332_),
    .A2(net266),
    .Y(_0051_),
    .B1(_0446_));
 sg13g2_nor2_1 _1320_ (.A(net240),
    .B(net266),
    .Y(_0447_));
 sg13g2_a21oi_1 _1321_ (.A1(_0334_),
    .A2(_0445_),
    .Y(_0052_),
    .B1(_0447_));
 sg13g2_nor2_1 _1322_ (.A(net239),
    .B(net266),
    .Y(_0448_));
 sg13g2_a21oi_1 _1323_ (.A1(_0336_),
    .A2(net266),
    .Y(_0053_),
    .B1(_0448_));
 sg13g2_nor2_1 _1324_ (.A(net241),
    .B(net266),
    .Y(_0449_));
 sg13g2_a21oi_1 _1325_ (.A1(_0338_),
    .A2(net266),
    .Y(_0054_),
    .B1(_0449_));
 sg13g2_nor2_1 _1326_ (.A(net324),
    .B(net267),
    .Y(_0450_));
 sg13g2_a21oi_1 _1327_ (.A1(_0340_),
    .A2(net267),
    .Y(_0055_),
    .B1(_0450_));
 sg13g2_nor2_1 _1328_ (.A(net244),
    .B(net267),
    .Y(_0451_));
 sg13g2_a21oi_1 _1329_ (.A1(_0342_),
    .A2(net267),
    .Y(_0056_),
    .B1(_0451_));
 sg13g2_nor2_1 _1330_ (.A(net334),
    .B(net266),
    .Y(_0452_));
 sg13g2_a21oi_1 _1331_ (.A1(_0344_),
    .A2(net267),
    .Y(_0057_),
    .B1(_0452_));
 sg13g2_nor2_1 _1332_ (.A(net338),
    .B(net267),
    .Y(_0453_));
 sg13g2_a21oi_1 _1333_ (.A1(_0346_),
    .A2(net267),
    .Y(_0058_),
    .B1(_0453_));
 sg13g2_nand4_1 _1334_ (.B(_0141_),
    .C(\result_addr[0] ),
    .A(net319),
    .Y(_0454_),
    .D(net3));
 sg13g2_and2_1 _1335_ (.A(net319),
    .B(net264),
    .X(_0455_));
 sg13g2_nand2_1 _1336_ (.Y(_0456_),
    .A(net192),
    .B(net249));
 sg13g2_o21ai_1 _1337_ (.B1(_0456_),
    .Y(_0059_),
    .A1(_0378_),
    .A2(net264));
 sg13g2_nand2_1 _1338_ (.Y(_0457_),
    .A(net242),
    .B(net248));
 sg13g2_o21ai_1 _1339_ (.B1(_0457_),
    .Y(_0060_),
    .A1(_0393_),
    .A2(net265));
 sg13g2_nand2_1 _1340_ (.Y(_0458_),
    .A(net184),
    .B(net248));
 sg13g2_o21ai_1 _1341_ (.B1(_0458_),
    .Y(_0061_),
    .A1(_0402_),
    .A2(net265));
 sg13g2_nand2_1 _1342_ (.Y(_0459_),
    .A(net193),
    .B(net248));
 sg13g2_o21ai_1 _1343_ (.B1(_0459_),
    .Y(_0062_),
    .A1(_0408_),
    .A2(net265));
 sg13g2_nand2_1 _1344_ (.Y(_0460_),
    .A(net197),
    .B(net248));
 sg13g2_o21ai_1 _1345_ (.B1(_0460_),
    .Y(_0063_),
    .A1(_0411_),
    .A2(net265));
 sg13g2_nand2_1 _1346_ (.Y(_0461_),
    .A(net199),
    .B(net249));
 sg13g2_o21ai_1 _1347_ (.B1(_0461_),
    .Y(_0064_),
    .A1(_0414_),
    .A2(net264));
 sg13g2_nand2_1 _1348_ (.Y(_0462_),
    .A(net208),
    .B(net249));
 sg13g2_o21ai_1 _1349_ (.B1(_0462_),
    .Y(_0065_),
    .A1(net282),
    .A2(net264));
 sg13g2_nand2_1 _1350_ (.Y(_0463_),
    .A(net213),
    .B(net249));
 sg13g2_o21ai_1 _1351_ (.B1(_0463_),
    .Y(_0066_),
    .A1(net282),
    .A2(_0454_));
 sg13g2_nor3_1 _1352_ (.A(net313),
    .B(net302),
    .C(_0329_),
    .Y(_0464_));
 sg13g2_nand2_1 _1353_ (.Y(_0465_),
    .A(_0140_),
    .B(_0464_));
 sg13g2_and2_2 _1354_ (.A(net321),
    .B(_0465_),
    .X(_0466_));
 sg13g2_nand2_1 _1355_ (.Y(_0467_),
    .A(net349),
    .B(_0466_));
 sg13g2_o21ai_1 _1356_ (.B1(_0467_),
    .Y(_0067_),
    .A1(_0332_),
    .A2(net247));
 sg13g2_nand2_1 _1357_ (.Y(_0468_),
    .A(net347),
    .B(_0466_));
 sg13g2_o21ai_1 _1358_ (.B1(_0468_),
    .Y(_0068_),
    .A1(_0334_),
    .A2(net247));
 sg13g2_nand2_1 _1359_ (.Y(_0469_),
    .A(net354),
    .B(_0466_));
 sg13g2_o21ai_1 _1360_ (.B1(_0469_),
    .Y(_0069_),
    .A1(_0336_),
    .A2(net247));
 sg13g2_nand2_1 _1361_ (.Y(_0470_),
    .A(net343),
    .B(_0466_));
 sg13g2_o21ai_1 _1362_ (.B1(_0470_),
    .Y(_0070_),
    .A1(_0338_),
    .A2(net247));
 sg13g2_nand2_1 _1363_ (.Y(_0471_),
    .A(net352),
    .B(_0466_));
 sg13g2_o21ai_1 _1364_ (.B1(_0471_),
    .Y(_0071_),
    .A1(_0340_),
    .A2(net247));
 sg13g2_nand2_1 _1365_ (.Y(_0472_),
    .A(net346),
    .B(_0466_));
 sg13g2_o21ai_1 _1366_ (.B1(_0472_),
    .Y(_0072_),
    .A1(_0342_),
    .A2(net247));
 sg13g2_nand2_1 _1367_ (.Y(_0473_),
    .A(net356),
    .B(_0466_));
 sg13g2_o21ai_1 _1368_ (.B1(_0473_),
    .Y(_0073_),
    .A1(_0344_),
    .A2(net247));
 sg13g2_nand2_1 _1369_ (.Y(_0474_),
    .A(net287),
    .B(_0466_));
 sg13g2_o21ai_1 _1370_ (.B1(_0474_),
    .Y(_0074_),
    .A1(_0346_),
    .A2(net247));
 sg13g2_nand4_1 _1371_ (.B(\result_addr[1] ),
    .C(net360),
    .A(net319),
    .Y(_0475_),
    .D(net3));
 sg13g2_and2_1 _1372_ (.A(net319),
    .B(net278),
    .X(_0476_));
 sg13g2_nand2_1 _1373_ (.Y(_0477_),
    .A(net211),
    .B(net263));
 sg13g2_o21ai_1 _1374_ (.B1(_0477_),
    .Y(_0075_),
    .A1(_0378_),
    .A2(net278));
 sg13g2_nand2_1 _1375_ (.Y(_0478_),
    .A(net187),
    .B(net262));
 sg13g2_o21ai_1 _1376_ (.B1(_0478_),
    .Y(_0076_),
    .A1(_0393_),
    .A2(net277));
 sg13g2_nand2_1 _1377_ (.Y(_0479_),
    .A(net171),
    .B(net262));
 sg13g2_o21ai_1 _1378_ (.B1(_0479_),
    .Y(_0077_),
    .A1(_0402_),
    .A2(net277));
 sg13g2_nand2_1 _1379_ (.Y(_0480_),
    .A(net177),
    .B(net262));
 sg13g2_o21ai_1 _1380_ (.B1(_0480_),
    .Y(_0078_),
    .A1(_0408_),
    .A2(net277));
 sg13g2_nand2_1 _1381_ (.Y(_0481_),
    .A(net202),
    .B(net262));
 sg13g2_o21ai_1 _1382_ (.B1(_0481_),
    .Y(_0079_),
    .A1(_0411_),
    .A2(net277));
 sg13g2_nand2_1 _1383_ (.Y(_0482_),
    .A(net165),
    .B(net263));
 sg13g2_o21ai_1 _1384_ (.B1(_0482_),
    .Y(_0080_),
    .A1(_0414_),
    .A2(net278));
 sg13g2_nor2_1 _1385_ (.A(net282),
    .B(net278),
    .Y(_0483_));
 sg13g2_a21o_1 _1386_ (.A2(net263),
    .A1(net344),
    .B1(_0483_),
    .X(_0081_));
 sg13g2_a21o_1 _1387_ (.A2(net263),
    .A1(net335),
    .B1(_0483_),
    .X(_0082_));
 sg13g2_nand2_1 _1388_ (.Y(_0484_),
    .A(net236),
    .B(net249));
 sg13g2_o21ai_1 _1389_ (.B1(_0484_),
    .Y(_0083_),
    .A1(_0160_),
    .A2(net264));
 sg13g2_nand2_1 _1390_ (.Y(_0485_),
    .A(net200),
    .B(net248));
 sg13g2_o21ai_1 _1391_ (.B1(_0485_),
    .Y(_0084_),
    .A1(_0181_),
    .A2(net265));
 sg13g2_nand2_1 _1392_ (.Y(_0486_),
    .A(net226),
    .B(net248));
 sg13g2_o21ai_1 _1393_ (.B1(_0486_),
    .Y(_0085_),
    .A1(_0195_),
    .A2(net265));
 sg13g2_nand2_1 _1394_ (.Y(_0487_),
    .A(net206),
    .B(net248));
 sg13g2_o21ai_1 _1395_ (.B1(_0487_),
    .Y(_0086_),
    .A1(_0218_),
    .A2(net265));
 sg13g2_nand2_1 _1396_ (.Y(_0488_),
    .A(net209),
    .B(net248));
 sg13g2_o21ai_1 _1397_ (.B1(_0488_),
    .Y(_0087_),
    .A1(_0244_),
    .A2(net265));
 sg13g2_nand2_1 _1398_ (.Y(_0489_),
    .A(net191),
    .B(net249));
 sg13g2_o21ai_1 _1399_ (.B1(_0489_),
    .Y(_0088_),
    .A1(_0275_),
    .A2(net264));
 sg13g2_nand2_1 _1400_ (.Y(_0490_),
    .A(net190),
    .B(net249));
 sg13g2_o21ai_1 _1401_ (.B1(_0490_),
    .Y(_0089_),
    .A1(_0299_),
    .A2(net264));
 sg13g2_nand2_1 _1402_ (.Y(_0491_),
    .A(net157),
    .B(net249));
 sg13g2_o21ai_1 _1403_ (.B1(_0491_),
    .Y(_0090_),
    .A1(_0326_),
    .A2(net264));
 sg13g2_nor3_1 _1404_ (.A(_0139_),
    .B(net296),
    .C(_0330_),
    .Y(_0492_));
 sg13g2_nor2_1 _1405_ (.A(net237),
    .B(net260),
    .Y(_0493_));
 sg13g2_a21oi_1 _1406_ (.A1(_0332_),
    .A2(net260),
    .Y(_0091_),
    .B1(_0493_));
 sg13g2_nor2_1 _1407_ (.A(net332),
    .B(_0492_),
    .Y(_0494_));
 sg13g2_a21oi_1 _1408_ (.A1(_0334_),
    .A2(net261),
    .Y(_0092_),
    .B1(_0494_));
 sg13g2_nor2_1 _1409_ (.A(net323),
    .B(net260),
    .Y(_0495_));
 sg13g2_a21oi_1 _1410_ (.A1(_0336_),
    .A2(net260),
    .Y(_0093_),
    .B1(_0495_));
 sg13g2_nor2_1 _1411_ (.A(net322),
    .B(net260),
    .Y(_0496_));
 sg13g2_a21oi_1 _1412_ (.A1(_0338_),
    .A2(net260),
    .Y(_0094_),
    .B1(_0496_));
 sg13g2_nor2_1 _1413_ (.A(net336),
    .B(net261),
    .Y(_0497_));
 sg13g2_a21oi_1 _1414_ (.A1(_0340_),
    .A2(net261),
    .Y(_0095_),
    .B1(_0497_));
 sg13g2_nor2_1 _1415_ (.A(net333),
    .B(net261),
    .Y(_0498_));
 sg13g2_a21oi_1 _1416_ (.A1(_0342_),
    .A2(net261),
    .Y(_0096_),
    .B1(_0498_));
 sg13g2_nor2_1 _1417_ (.A(net243),
    .B(net260),
    .Y(_0499_));
 sg13g2_a21oi_1 _1418_ (.A1(_0344_),
    .A2(net260),
    .Y(_0097_),
    .B1(_0499_));
 sg13g2_nor2_1 _1419_ (.A(net342),
    .B(net261),
    .Y(_0500_));
 sg13g2_a21oi_1 _1420_ (.A1(_0346_),
    .A2(net261),
    .Y(_0098_),
    .B1(_0500_));
 sg13g2_o21ai_1 _1421_ (.B1(net289),
    .Y(_0501_),
    .A1(net291),
    .A2(net302));
 sg13g2_nand3_1 _1422_ (.B(net289),
    .C(_0501_),
    .A(net298),
    .Y(_0502_));
 sg13g2_nand2_1 _1423_ (.Y(_0503_),
    .A(net162),
    .B(net258));
 sg13g2_o21ai_1 _1424_ (.B1(_0503_),
    .Y(_0099_),
    .A1(_0332_),
    .A2(net258));
 sg13g2_nand2_1 _1425_ (.Y(_0504_),
    .A(net205),
    .B(net258));
 sg13g2_o21ai_1 _1426_ (.B1(_0504_),
    .Y(_0100_),
    .A1(_0334_),
    .A2(net258));
 sg13g2_nand2_1 _1427_ (.Y(_0505_),
    .A(net163),
    .B(net258));
 sg13g2_o21ai_1 _1428_ (.B1(_0505_),
    .Y(_0101_),
    .A1(_0336_),
    .A2(net258));
 sg13g2_nand2_1 _1429_ (.Y(_0506_),
    .A(net169),
    .B(_0502_));
 sg13g2_o21ai_1 _1430_ (.B1(_0506_),
    .Y(_0102_),
    .A1(_0338_),
    .A2(net258));
 sg13g2_nand2_1 _1431_ (.Y(_0507_),
    .A(net159),
    .B(net259));
 sg13g2_o21ai_1 _1432_ (.B1(_0507_),
    .Y(_0103_),
    .A1(_0340_),
    .A2(net259));
 sg13g2_nand2_1 _1433_ (.Y(_0508_),
    .A(net195),
    .B(net259));
 sg13g2_o21ai_1 _1434_ (.B1(_0508_),
    .Y(_0104_),
    .A1(_0342_),
    .A2(net259));
 sg13g2_nand2_1 _1435_ (.Y(_0509_),
    .A(net152),
    .B(net258));
 sg13g2_o21ai_1 _1436_ (.B1(_0509_),
    .Y(_0105_),
    .A1(_0344_),
    .A2(net259));
 sg13g2_nand2_1 _1437_ (.Y(_0510_),
    .A(net166),
    .B(net259));
 sg13g2_o21ai_1 _1438_ (.B1(_0510_),
    .Y(_0106_),
    .A1(_0346_),
    .A2(net259));
 sg13g2_mux4_1 _1439_ (.S0(net317),
    .A0(\a[0] ),
    .A1(\b[0] ),
    .A2(\ram[10][0] ),
    .A3(\ram[11][0] ),
    .S1(net304),
    .X(_0511_));
 sg13g2_mux2_1 _1440_ (.A0(\ram[14][0] ),
    .A1(\ram[15][0] ),
    .S(net316),
    .X(_0512_));
 sg13g2_nand2b_1 _1441_ (.Y(_0513_),
    .B(net317),
    .A_N(\ram[13][0] ));
 sg13g2_o21ai_1 _1442_ (.B1(_0513_),
    .Y(_0514_),
    .A1(net317),
    .A2(\ram[12][0] ));
 sg13g2_o21ai_1 _1443_ (.B1(net298),
    .Y(_0515_),
    .A1(net303),
    .A2(_0514_));
 sg13g2_a21oi_1 _1444_ (.A1(net303),
    .A2(_0512_),
    .Y(_0516_),
    .B1(_0515_));
 sg13g2_nor2b_1 _1445_ (.A(_0516_),
    .B_N(net2),
    .Y(_0517_));
 sg13g2_o21ai_1 _1446_ (.B1(_0517_),
    .Y(_0518_),
    .A1(net297),
    .A2(_0511_));
 sg13g2_mux4_1 _1447_ (.S0(net312),
    .A0(\ram[0][0] ),
    .A1(\ram[1][0] ),
    .A2(\ram[2][0] ),
    .A3(\ram[3][0] ),
    .S1(net301),
    .X(_0519_));
 sg13g2_nand2b_1 _1448_ (.Y(_0520_),
    .B(net312),
    .A_N(\ram[5][0] ));
 sg13g2_o21ai_1 _1449_ (.B1(_0520_),
    .Y(_0521_),
    .A1(net312),
    .A2(\ram[4][0] ));
 sg13g2_nor2_1 _1450_ (.A(net312),
    .B(\ram[6][0] ),
    .Y(_0522_));
 sg13g2_o21ai_1 _1451_ (.B1(net301),
    .Y(_0523_),
    .A1(net291),
    .A2(\ram[7][0] ));
 sg13g2_o21ai_1 _1452_ (.B1(net1),
    .Y(_0524_),
    .A1(_0522_),
    .A2(_0523_));
 sg13g2_inv_1 _1453_ (.Y(_0525_),
    .A(_0524_));
 sg13g2_o21ai_1 _1454_ (.B1(_0525_),
    .Y(_0526_),
    .A1(net301),
    .A2(_0521_));
 sg13g2_o21ai_1 _1455_ (.B1(_0526_),
    .Y(_0527_),
    .A1(net295),
    .A2(_0519_));
 sg13g2_o21ai_1 _1456_ (.B1(_0518_),
    .Y(_0528_),
    .A1(net293),
    .A2(_0527_));
 sg13g2_and2_1 _1457_ (.A(net321),
    .B(_0528_),
    .X(_0107_));
 sg13g2_mux4_1 _1458_ (.S0(net317),
    .A0(\a[1] ),
    .A1(\b[1] ),
    .A2(\ram[10][1] ),
    .A3(\ram[11][1] ),
    .S1(net304),
    .X(_0529_));
 sg13g2_mux2_1 _1459_ (.A0(\ram[14][1] ),
    .A1(\ram[15][1] ),
    .S(net315),
    .X(_0530_));
 sg13g2_nand2b_1 _1460_ (.Y(_0531_),
    .B(net315),
    .A_N(\ram[13][1] ));
 sg13g2_o21ai_1 _1461_ (.B1(_0531_),
    .Y(_0532_),
    .A1(net315),
    .A2(\ram[12][1] ));
 sg13g2_o21ai_1 _1462_ (.B1(net298),
    .Y(_0533_),
    .A1(net304),
    .A2(_0532_));
 sg13g2_a21oi_1 _1463_ (.A1(net305),
    .A2(_0530_),
    .Y(_0534_),
    .B1(_0533_));
 sg13g2_nor2b_1 _1464_ (.A(_0534_),
    .B_N(net2),
    .Y(_0535_));
 sg13g2_o21ai_1 _1465_ (.B1(_0535_),
    .Y(_0536_),
    .A1(net297),
    .A2(_0529_));
 sg13g2_mux4_1 _1466_ (.S0(net311),
    .A0(\ram[0][1] ),
    .A1(\ram[1][1] ),
    .A2(\ram[2][1] ),
    .A3(\ram[3][1] ),
    .S1(net306),
    .X(_0537_));
 sg13g2_nand2b_1 _1467_ (.Y(_0538_),
    .B(net311),
    .A_N(\ram[5][1] ));
 sg13g2_o21ai_1 _1468_ (.B1(_0538_),
    .Y(_0539_),
    .A1(net311),
    .A2(\ram[4][1] ));
 sg13g2_nor2_1 _1469_ (.A(net311),
    .B(\ram[6][1] ),
    .Y(_0540_));
 sg13g2_o21ai_1 _1470_ (.B1(net301),
    .Y(_0541_),
    .A1(net291),
    .A2(\ram[7][1] ));
 sg13g2_o21ai_1 _1471_ (.B1(net295),
    .Y(_0542_),
    .A1(_0540_),
    .A2(_0541_));
 sg13g2_inv_1 _1472_ (.Y(_0543_),
    .A(_0542_));
 sg13g2_o21ai_1 _1473_ (.B1(_0543_),
    .Y(_0544_),
    .A1(net301),
    .A2(_0539_));
 sg13g2_o21ai_1 _1474_ (.B1(_0544_),
    .Y(_0545_),
    .A1(net295),
    .A2(_0537_));
 sg13g2_o21ai_1 _1475_ (.B1(_0536_),
    .Y(_0546_),
    .A1(net292),
    .A2(_0545_));
 sg13g2_and2_1 _1476_ (.A(net321),
    .B(_0546_),
    .X(_0108_));
 sg13g2_mux4_1 _1477_ (.S0(net317),
    .A0(\a[2] ),
    .A1(\b[2] ),
    .A2(\ram[10][2] ),
    .A3(\ram[11][2] ),
    .S1(net304),
    .X(_0547_));
 sg13g2_mux2_1 _1478_ (.A0(\ram[14][2] ),
    .A1(\ram[15][2] ),
    .S(net317),
    .X(_0548_));
 sg13g2_nand2b_1 _1479_ (.Y(_0549_),
    .B(net315),
    .A_N(\ram[13][2] ));
 sg13g2_o21ai_1 _1480_ (.B1(_0549_),
    .Y(_0550_),
    .A1(net315),
    .A2(\ram[12][2] ));
 sg13g2_o21ai_1 _1481_ (.B1(net297),
    .Y(_0551_),
    .A1(net303),
    .A2(_0550_));
 sg13g2_a21oi_1 _1482_ (.A1(net304),
    .A2(_0548_),
    .Y(_0552_),
    .B1(_0551_));
 sg13g2_nor2b_1 _1483_ (.A(_0552_),
    .B_N(net2),
    .Y(_0553_));
 sg13g2_o21ai_1 _1484_ (.B1(_0553_),
    .Y(_0554_),
    .A1(net297),
    .A2(_0547_));
 sg13g2_mux4_1 _1485_ (.S0(net308),
    .A0(\ram[0][2] ),
    .A1(\ram[1][2] ),
    .A2(\ram[2][2] ),
    .A3(\ram[3][2] ),
    .S1(net306),
    .X(_0555_));
 sg13g2_nand2b_1 _1486_ (.Y(_0556_),
    .B(net308),
    .A_N(\ram[5][2] ));
 sg13g2_o21ai_1 _1487_ (.B1(_0556_),
    .Y(_0557_),
    .A1(net308),
    .A2(\ram[4][2] ));
 sg13g2_nor2_1 _1488_ (.A(net308),
    .B(\ram[6][2] ),
    .Y(_0558_));
 sg13g2_o21ai_1 _1489_ (.B1(net299),
    .Y(_0559_),
    .A1(net291),
    .A2(\ram[7][2] ));
 sg13g2_o21ai_1 _1490_ (.B1(net294),
    .Y(_0560_),
    .A1(_0558_),
    .A2(_0559_));
 sg13g2_inv_1 _1491_ (.Y(_0561_),
    .A(_0560_));
 sg13g2_o21ai_1 _1492_ (.B1(_0561_),
    .Y(_0562_),
    .A1(net299),
    .A2(_0557_));
 sg13g2_o21ai_1 _1493_ (.B1(_0562_),
    .Y(_0563_),
    .A1(net294),
    .A2(_0555_));
 sg13g2_o21ai_1 _1494_ (.B1(_0554_),
    .Y(_0564_),
    .A1(net292),
    .A2(_0563_));
 sg13g2_and2_1 _1495_ (.A(net320),
    .B(_0564_),
    .X(_0109_));
 sg13g2_mux4_1 _1496_ (.S0(net317),
    .A0(\a[3] ),
    .A1(\b[3] ),
    .A2(\ram[10][3] ),
    .A3(\ram[11][3] ),
    .S1(net304),
    .X(_0565_));
 sg13g2_mux2_1 _1497_ (.A0(\ram[14][3] ),
    .A1(\ram[15][3] ),
    .S(net315),
    .X(_0566_));
 sg13g2_nand2b_1 _1498_ (.Y(_0567_),
    .B(net315),
    .A_N(\ram[13][3] ));
 sg13g2_o21ai_1 _1499_ (.B1(_0567_),
    .Y(_0568_),
    .A1(net315),
    .A2(\ram[12][3] ));
 sg13g2_o21ai_1 _1500_ (.B1(net298),
    .Y(_0569_),
    .A1(net305),
    .A2(_0568_));
 sg13g2_a21oi_1 _1501_ (.A1(net303),
    .A2(_0566_),
    .Y(_0570_),
    .B1(_0569_));
 sg13g2_nor2b_1 _1502_ (.A(_0570_),
    .B_N(net293),
    .Y(_0571_));
 sg13g2_o21ai_1 _1503_ (.B1(_0571_),
    .Y(_0572_),
    .A1(net297),
    .A2(_0565_));
 sg13g2_mux4_1 _1504_ (.S0(net307),
    .A0(\ram[0][3] ),
    .A1(\ram[1][3] ),
    .A2(\ram[2][3] ),
    .A3(\ram[3][3] ),
    .S1(net299),
    .X(_0573_));
 sg13g2_nand2b_1 _1505_ (.Y(_0574_),
    .B(net307),
    .A_N(\ram[5][3] ));
 sg13g2_o21ai_1 _1506_ (.B1(_0574_),
    .Y(_0575_),
    .A1(net307),
    .A2(\ram[4][3] ));
 sg13g2_nor2_1 _1507_ (.A(net307),
    .B(\ram[6][3] ),
    .Y(_0576_));
 sg13g2_o21ai_1 _1508_ (.B1(net299),
    .Y(_0577_),
    .A1(net291),
    .A2(\ram[7][3] ));
 sg13g2_o21ai_1 _1509_ (.B1(net294),
    .Y(_0578_),
    .A1(_0576_),
    .A2(_0577_));
 sg13g2_inv_1 _1510_ (.Y(_0579_),
    .A(_0578_));
 sg13g2_o21ai_1 _1511_ (.B1(_0579_),
    .Y(_0580_),
    .A1(net299),
    .A2(_0575_));
 sg13g2_o21ai_1 _1512_ (.B1(_0580_),
    .Y(_0581_),
    .A1(net294),
    .A2(_0573_));
 sg13g2_o21ai_1 _1513_ (.B1(_0572_),
    .Y(_0582_),
    .A1(net292),
    .A2(_0581_));
 sg13g2_and2_1 _1514_ (.A(net321),
    .B(_0582_),
    .X(_0110_));
 sg13g2_mux4_1 _1515_ (.S0(net314),
    .A0(\a[4] ),
    .A1(\b[4] ),
    .A2(\ram[10][4] ),
    .A3(\ram[11][4] ),
    .S1(net302),
    .X(_0583_));
 sg13g2_mux2_1 _1516_ (.A0(\ram[14][4] ),
    .A1(\ram[15][4] ),
    .S(net316),
    .X(_0584_));
 sg13g2_nand2b_1 _1517_ (.Y(_0585_),
    .B(net316),
    .A_N(\ram[13][4] ));
 sg13g2_o21ai_1 _1518_ (.B1(_0585_),
    .Y(_0586_),
    .A1(net316),
    .A2(\ram[12][4] ));
 sg13g2_o21ai_1 _1519_ (.B1(net297),
    .Y(_0587_),
    .A1(net303),
    .A2(_0586_));
 sg13g2_a21oi_1 _1520_ (.A1(net303),
    .A2(_0584_),
    .Y(_0588_),
    .B1(_0587_));
 sg13g2_nor2b_1 _1521_ (.A(_0588_),
    .B_N(net293),
    .Y(_0589_));
 sg13g2_o21ai_1 _1522_ (.B1(_0589_),
    .Y(_0590_),
    .A1(net296),
    .A2(_0583_));
 sg13g2_mux4_1 _1523_ (.S0(net307),
    .A0(\ram[0][4] ),
    .A1(\ram[1][4] ),
    .A2(\ram[2][4] ),
    .A3(\ram[3][4] ),
    .S1(net299),
    .X(_0591_));
 sg13g2_a21oi_1 _1524_ (.A1(net307),
    .A2(_0143_),
    .Y(_0592_),
    .B1(net299));
 sg13g2_o21ai_1 _1525_ (.B1(_0592_),
    .Y(_0593_),
    .A1(net307),
    .A2(\ram[4][4] ));
 sg13g2_nor2_1 _1526_ (.A(net307),
    .B(\ram[6][4] ),
    .Y(_0594_));
 sg13g2_o21ai_1 _1527_ (.B1(net299),
    .Y(_0595_),
    .A1(net291),
    .A2(\ram[7][4] ));
 sg13g2_o21ai_1 _1528_ (.B1(net294),
    .Y(_0596_),
    .A1(_0594_),
    .A2(_0595_));
 sg13g2_nand2b_1 _1529_ (.Y(_0597_),
    .B(_0593_),
    .A_N(_0596_));
 sg13g2_o21ai_1 _1530_ (.B1(_0597_),
    .Y(_0598_),
    .A1(net294),
    .A2(_0591_));
 sg13g2_o21ai_1 _1531_ (.B1(_0590_),
    .Y(_0599_),
    .A1(net292),
    .A2(_0598_));
 sg13g2_and2_1 _1532_ (.A(net320),
    .B(_0599_),
    .X(_0111_));
 sg13g2_mux4_1 _1533_ (.S0(net314),
    .A0(\a[5] ),
    .A1(\b[5] ),
    .A2(\ram[10][5] ),
    .A3(\ram[11][5] ),
    .S1(net302),
    .X(_0600_));
 sg13g2_mux2_1 _1534_ (.A0(\ram[14][5] ),
    .A1(\ram[15][5] ),
    .S(net313),
    .X(_0601_));
 sg13g2_nand2b_1 _1535_ (.Y(_0602_),
    .B(net313),
    .A_N(\ram[13][5] ));
 sg13g2_o21ai_1 _1536_ (.B1(_0602_),
    .Y(_0603_),
    .A1(net314),
    .A2(\ram[12][5] ));
 sg13g2_o21ai_1 _1537_ (.B1(net296),
    .Y(_0604_),
    .A1(net305),
    .A2(_0603_));
 sg13g2_a21oi_1 _1538_ (.A1(net305),
    .A2(_0601_),
    .Y(_0605_),
    .B1(_0604_));
 sg13g2_nor2b_1 _1539_ (.A(_0605_),
    .B_N(net292),
    .Y(_0606_));
 sg13g2_o21ai_1 _1540_ (.B1(_0606_),
    .Y(_0607_),
    .A1(net296),
    .A2(_0600_));
 sg13g2_mux4_1 _1541_ (.S0(net309),
    .A0(\ram[0][5] ),
    .A1(\ram[1][5] ),
    .A2(\ram[2][5] ),
    .A3(\ram[3][5] ),
    .S1(net300),
    .X(_0608_));
 sg13g2_a21oi_1 _1542_ (.A1(net309),
    .A2(_0144_),
    .Y(_0609_),
    .B1(net300));
 sg13g2_o21ai_1 _1543_ (.B1(_0609_),
    .Y(_0610_),
    .A1(net309),
    .A2(\ram[4][5] ));
 sg13g2_nor2_1 _1544_ (.A(net309),
    .B(\ram[6][5] ),
    .Y(_0611_));
 sg13g2_o21ai_1 _1545_ (.B1(net300),
    .Y(_0612_),
    .A1(net291),
    .A2(\ram[7][5] ));
 sg13g2_o21ai_1 _1546_ (.B1(net295),
    .Y(_0613_),
    .A1(_0611_),
    .A2(_0612_));
 sg13g2_nand2b_1 _1547_ (.Y(_0614_),
    .B(_0610_),
    .A_N(_0613_));
 sg13g2_o21ai_1 _1548_ (.B1(_0614_),
    .Y(_0615_),
    .A1(net294),
    .A2(_0608_));
 sg13g2_o21ai_1 _1549_ (.B1(_0607_),
    .Y(_0616_),
    .A1(net292),
    .A2(_0615_));
 sg13g2_and2_1 _1550_ (.A(net320),
    .B(_0616_),
    .X(_0112_));
 sg13g2_mux4_1 _1551_ (.S0(net314),
    .A0(\a[6] ),
    .A1(\b[6] ),
    .A2(\ram[10][6] ),
    .A3(\ram[11][6] ),
    .S1(net304),
    .X(_0617_));
 sg13g2_mux2_1 _1552_ (.A0(\ram[14][6] ),
    .A1(\ram[15][6] ),
    .S(net316),
    .X(_0618_));
 sg13g2_nand2b_1 _1553_ (.Y(_0619_),
    .B(net316),
    .A_N(\ram[13][6] ));
 sg13g2_o21ai_1 _1554_ (.B1(_0619_),
    .Y(_0620_),
    .A1(net316),
    .A2(\ram[12][6] ));
 sg13g2_o21ai_1 _1555_ (.B1(net297),
    .Y(_0621_),
    .A1(net303),
    .A2(_0620_));
 sg13g2_a21oi_1 _1556_ (.A1(net303),
    .A2(_0618_),
    .Y(_0622_),
    .B1(_0621_));
 sg13g2_nor2b_1 _1557_ (.A(_0622_),
    .B_N(net293),
    .Y(_0623_));
 sg13g2_o21ai_1 _1558_ (.B1(_0623_),
    .Y(_0624_),
    .A1(net297),
    .A2(_0617_));
 sg13g2_mux4_1 _1559_ (.S0(net309),
    .A0(\ram[0][6] ),
    .A1(\ram[1][6] ),
    .A2(\ram[2][6] ),
    .A3(\ram[3][6] ),
    .S1(net300),
    .X(_0625_));
 sg13g2_nand2b_1 _1560_ (.Y(_0626_),
    .B(net309),
    .A_N(\ram[5][6] ));
 sg13g2_o21ai_1 _1561_ (.B1(_0626_),
    .Y(_0627_),
    .A1(net309),
    .A2(\ram[4][6] ));
 sg13g2_nor2_1 _1562_ (.A(net309),
    .B(\ram[6][6] ),
    .Y(_0628_));
 sg13g2_o21ai_1 _1563_ (.B1(net300),
    .Y(_0629_),
    .A1(net291),
    .A2(\ram[7][6] ));
 sg13g2_o21ai_1 _1564_ (.B1(net294),
    .Y(_0630_),
    .A1(_0628_),
    .A2(_0629_));
 sg13g2_inv_1 _1565_ (.Y(_0631_),
    .A(_0630_));
 sg13g2_o21ai_1 _1566_ (.B1(_0631_),
    .Y(_0632_),
    .A1(net300),
    .A2(_0627_));
 sg13g2_o21ai_1 _1567_ (.B1(_0632_),
    .Y(_0633_),
    .A1(net295),
    .A2(_0625_));
 sg13g2_o21ai_1 _1568_ (.B1(_0624_),
    .Y(_0634_),
    .A1(net292),
    .A2(_0633_));
 sg13g2_and2_1 _1569_ (.A(net320),
    .B(_0634_),
    .X(_0113_));
 sg13g2_mux4_1 _1570_ (.S0(net310),
    .A0(\ram[0][7] ),
    .A1(\ram[1][7] ),
    .A2(\ram[2][7] ),
    .A3(\ram[3][7] ),
    .S1(net300),
    .X(_0635_));
 sg13g2_a21oi_1 _1571_ (.A1(net311),
    .A2(_0145_),
    .Y(_0636_),
    .B1(net301));
 sg13g2_o21ai_1 _1572_ (.B1(_0636_),
    .Y(_0637_),
    .A1(net311),
    .A2(\ram[4][7] ));
 sg13g2_o21ai_1 _1573_ (.B1(net300),
    .Y(_0638_),
    .A1(net311),
    .A2(\ram[6][7] ));
 sg13g2_a21oi_1 _1574_ (.A1(net312),
    .A2(_0146_),
    .Y(_0639_),
    .B1(_0638_));
 sg13g2_nor2_1 _1575_ (.A(_0140_),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_a21oi_1 _1576_ (.A1(_0637_),
    .A2(_0640_),
    .Y(_0641_),
    .B1(net292));
 sg13g2_o21ai_1 _1577_ (.B1(_0641_),
    .Y(_0642_),
    .A1(net295),
    .A2(_0635_));
 sg13g2_mux2_1 _1578_ (.A0(\ram[14][7] ),
    .A1(\ram[15][7] ),
    .S(net313),
    .X(_0643_));
 sg13g2_nand2b_1 _1579_ (.Y(_0644_),
    .B(net313),
    .A_N(\ram[13][7] ));
 sg13g2_o21ai_1 _1580_ (.B1(_0644_),
    .Y(_0645_),
    .A1(net314),
    .A2(\ram[12][7] ));
 sg13g2_o21ai_1 _1581_ (.B1(net298),
    .Y(_0646_),
    .A1(net302),
    .A2(_0645_));
 sg13g2_a21oi_1 _1582_ (.A1(net302),
    .A2(_0643_),
    .Y(_0647_),
    .B1(_0646_));
 sg13g2_mux4_1 _1583_ (.S0(net314),
    .A0(net288),
    .A1(net286),
    .A2(\ram[10][7] ),
    .A3(\ram[11][7] ),
    .S1(net302),
    .X(_0648_));
 sg13g2_o21ai_1 _1584_ (.B1(net293),
    .Y(_0649_),
    .A1(net296),
    .A2(_0648_));
 sg13g2_o21ai_1 _1585_ (.B1(_0642_),
    .Y(_0650_),
    .A1(_0647_),
    .A2(_0649_));
 sg13g2_and2_1 _1586_ (.A(net320),
    .B(_0650_),
    .X(_0114_));
 sg13g2_and2_1 _1587_ (.A(net296),
    .B(_0464_),
    .X(_0651_));
 sg13g2_nor2_1 _1588_ (.A(net337),
    .B(net245),
    .Y(_0652_));
 sg13g2_a21oi_1 _1589_ (.A1(_0332_),
    .A2(net245),
    .Y(_0115_),
    .B1(_0652_));
 sg13g2_nor2_1 _1590_ (.A(net325),
    .B(net245),
    .Y(_0653_));
 sg13g2_a21oi_1 _1591_ (.A1(_0334_),
    .A2(net245),
    .Y(_0116_),
    .B1(_0653_));
 sg13g2_nor2_1 _1592_ (.A(net339),
    .B(net245),
    .Y(_0654_));
 sg13g2_a21oi_1 _1593_ (.A1(_0336_),
    .A2(net245),
    .Y(_0117_),
    .B1(_0654_));
 sg13g2_nor2_1 _1594_ (.A(net331),
    .B(_0651_),
    .Y(_0655_));
 sg13g2_a21oi_1 _1595_ (.A1(_0338_),
    .A2(net245),
    .Y(_0118_),
    .B1(_0655_));
 sg13g2_nor2_1 _1596_ (.A(net233),
    .B(net246),
    .Y(_0656_));
 sg13g2_a21oi_1 _1597_ (.A1(_0340_),
    .A2(net246),
    .Y(_0119_),
    .B1(_0656_));
 sg13g2_nor2_1 _1598_ (.A(net341),
    .B(net246),
    .Y(_0657_));
 sg13g2_a21oi_1 _1599_ (.A1(_0342_),
    .A2(net246),
    .Y(_0120_),
    .B1(_0657_));
 sg13g2_nor2_1 _1600_ (.A(net340),
    .B(net245),
    .Y(_0658_));
 sg13g2_a21oi_1 _1601_ (.A1(_0344_),
    .A2(net246),
    .Y(_0121_),
    .B1(_0658_));
 sg13g2_nor2_1 _1602_ (.A(net330),
    .B(net246),
    .Y(_0659_));
 sg13g2_a21oi_1 _1603_ (.A1(_0346_),
    .A2(net246),
    .Y(_0122_),
    .B1(_0659_));
 sg13g2_o21ai_1 _1604_ (.B1(net321),
    .Y(_0660_),
    .A1(net298),
    .A2(_0327_));
 sg13g2_nand2_1 _1605_ (.Y(_0661_),
    .A(_0501_),
    .B(_0660_));
 sg13g2_nand2_1 _1606_ (.Y(_0662_),
    .A(net351),
    .B(net256));
 sg13g2_o21ai_1 _1607_ (.B1(_0662_),
    .Y(_0123_),
    .A1(_0332_),
    .A2(net256));
 sg13g2_nand2_1 _1608_ (.Y(_0663_),
    .A(net350),
    .B(net256));
 sg13g2_o21ai_1 _1609_ (.B1(_0663_),
    .Y(_0124_),
    .A1(_0334_),
    .A2(_0661_));
 sg13g2_nand2_1 _1610_ (.Y(_0664_),
    .A(net355),
    .B(net256));
 sg13g2_o21ai_1 _1611_ (.B1(_0664_),
    .Y(_0125_),
    .A1(_0336_),
    .A2(net256));
 sg13g2_nand2_1 _1612_ (.Y(_0665_),
    .A(net345),
    .B(net256));
 sg13g2_o21ai_1 _1613_ (.B1(_0665_),
    .Y(_0126_),
    .A1(_0338_),
    .A2(net256));
 sg13g2_nand2_1 _1614_ (.Y(_0666_),
    .A(net353),
    .B(net257));
 sg13g2_o21ai_1 _1615_ (.B1(_0666_),
    .Y(_0127_),
    .A1(_0340_),
    .A2(net257));
 sg13g2_nand2_1 _1616_ (.Y(_0667_),
    .A(net348),
    .B(net257));
 sg13g2_o21ai_1 _1617_ (.B1(_0667_),
    .Y(_0128_),
    .A1(_0342_),
    .A2(net257));
 sg13g2_nand2_1 _1618_ (.Y(_0668_),
    .A(net357),
    .B(net256));
 sg13g2_o21ai_1 _1619_ (.B1(_0668_),
    .Y(_0129_),
    .A1(_0344_),
    .A2(net257));
 sg13g2_nand2_1 _1620_ (.Y(_0669_),
    .A(net285),
    .B(net257));
 sg13g2_o21ai_1 _1621_ (.B1(_0669_),
    .Y(_0130_),
    .A1(_0346_),
    .A2(net257));
 sg13g2_nand2_1 _1622_ (.Y(_0670_),
    .A(net198),
    .B(net263));
 sg13g2_o21ai_1 _1623_ (.B1(_0670_),
    .Y(_0131_),
    .A1(_0160_),
    .A2(net278));
 sg13g2_nand2_1 _1624_ (.Y(_0671_),
    .A(net155),
    .B(net262));
 sg13g2_o21ai_1 _1625_ (.B1(_0671_),
    .Y(_0132_),
    .A1(_0181_),
    .A2(net277));
 sg13g2_nand2_1 _1626_ (.Y(_0672_),
    .A(net170),
    .B(net262));
 sg13g2_o21ai_1 _1627_ (.B1(_0672_),
    .Y(_0133_),
    .A1(_0195_),
    .A2(net277));
 sg13g2_nand2_1 _1628_ (.Y(_0673_),
    .A(net229),
    .B(net262));
 sg13g2_o21ai_1 _1629_ (.B1(_0673_),
    .Y(_0134_),
    .A1(_0218_),
    .A2(net277));
 sg13g2_nand2_1 _1630_ (.Y(_0674_),
    .A(net204),
    .B(net262));
 sg13g2_o21ai_1 _1631_ (.B1(_0674_),
    .Y(_0135_),
    .A1(_0244_),
    .A2(net277));
 sg13g2_nand2_1 _1632_ (.Y(_0675_),
    .A(net225),
    .B(net263));
 sg13g2_o21ai_1 _1633_ (.B1(_0675_),
    .Y(_0136_),
    .A1(_0275_),
    .A2(net278));
 sg13g2_nand2_1 _1634_ (.Y(_0676_),
    .A(net176),
    .B(net263));
 sg13g2_o21ai_1 _1635_ (.B1(_0676_),
    .Y(_0137_),
    .A1(_0299_),
    .A2(net278));
 sg13g2_nand2_1 _1636_ (.Y(_0677_),
    .A(net168),
    .B(net263));
 sg13g2_o21ai_1 _1637_ (.B1(_0677_),
    .Y(_0138_),
    .A1(_0326_),
    .A2(net278));
 sg13g2_dfrbp_1 _1638_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net149),
    .D(_0001_),
    .Q_N(_0814_),
    .Q(\ram[15][0] ));
 sg13g2_dfrbp_1 _1639_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net91),
    .D(_0002_),
    .Q_N(_0813_),
    .Q(\ram[15][1] ));
 sg13g2_dfrbp_1 _1640_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net90),
    .D(_0003_),
    .Q_N(_0812_),
    .Q(\ram[15][2] ));
 sg13g2_dfrbp_1 _1641_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net89),
    .D(_0004_),
    .Q_N(_0811_),
    .Q(\ram[15][3] ));
 sg13g2_dfrbp_1 _1642_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net88),
    .D(_0005_),
    .Q_N(_0810_),
    .Q(\ram[15][4] ));
 sg13g2_dfrbp_1 _1643_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net87),
    .D(_0006_),
    .Q_N(_0809_),
    .Q(\ram[15][5] ));
 sg13g2_dfrbp_1 _1644_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net86),
    .D(_0007_),
    .Q_N(_0808_),
    .Q(\ram[15][6] ));
 sg13g2_dfrbp_1 _1645_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net85),
    .D(_0008_),
    .Q_N(_0807_),
    .Q(\ram[15][7] ));
 sg13g2_dfrbp_1 _1646_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net84),
    .D(_0009_),
    .Q_N(_0000_),
    .Q(\result_addr[0] ));
 sg13g2_dfrbp_1 _1647_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net83),
    .D(_0010_),
    .Q_N(_0806_),
    .Q(\result_addr[1] ));
 sg13g2_dfrbp_1 _1648_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net82),
    .D(_0011_),
    .Q_N(_0805_),
    .Q(\ram[0][0] ));
 sg13g2_dfrbp_1 _1649_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net81),
    .D(_0012_),
    .Q_N(_0804_),
    .Q(\ram[0][1] ));
 sg13g2_dfrbp_1 _1650_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net80),
    .D(_0013_),
    .Q_N(_0803_),
    .Q(\ram[0][2] ));
 sg13g2_dfrbp_1 _1651_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net79),
    .D(_0014_),
    .Q_N(_0802_),
    .Q(\ram[0][3] ));
 sg13g2_dfrbp_1 _1652_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net78),
    .D(_0015_),
    .Q_N(_0801_),
    .Q(\ram[0][4] ));
 sg13g2_dfrbp_1 _1653_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net77),
    .D(_0016_),
    .Q_N(_0800_),
    .Q(\ram[0][5] ));
 sg13g2_dfrbp_1 _1654_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net76),
    .D(_0017_),
    .Q_N(_0799_),
    .Q(\ram[0][6] ));
 sg13g2_dfrbp_1 _1655_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net75),
    .D(net161),
    .Q_N(_0798_),
    .Q(\ram[0][7] ));
 sg13g2_dfrbp_1 _1656_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net74),
    .D(_0019_),
    .Q_N(_0797_),
    .Q(\ram[1][0] ));
 sg13g2_dfrbp_1 _1657_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net73),
    .D(_0020_),
    .Q_N(_0796_),
    .Q(\ram[1][1] ));
 sg13g2_dfrbp_1 _1658_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net72),
    .D(_0021_),
    .Q_N(_0795_),
    .Q(\ram[1][2] ));
 sg13g2_dfrbp_1 _1659_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net71),
    .D(_0022_),
    .Q_N(_0794_),
    .Q(\ram[1][3] ));
 sg13g2_dfrbp_1 _1660_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net70),
    .D(_0023_),
    .Q_N(_0793_),
    .Q(\ram[1][4] ));
 sg13g2_dfrbp_1 _1661_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net69),
    .D(_0024_),
    .Q_N(_0792_),
    .Q(\ram[1][5] ));
 sg13g2_dfrbp_1 _1662_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net68),
    .D(_0025_),
    .Q_N(_0791_),
    .Q(\ram[1][6] ));
 sg13g2_dfrbp_1 _1663_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net67),
    .D(_0026_),
    .Q_N(_0790_),
    .Q(\ram[1][7] ));
 sg13g2_dfrbp_1 _1664_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net66),
    .D(_0027_),
    .Q_N(_0789_),
    .Q(\ram[5][0] ));
 sg13g2_dfrbp_1 _1665_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net65),
    .D(_0028_),
    .Q_N(_0788_),
    .Q(\ram[5][1] ));
 sg13g2_dfrbp_1 _1666_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net64),
    .D(_0029_),
    .Q_N(_0787_),
    .Q(\ram[5][2] ));
 sg13g2_dfrbp_1 _1667_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net63),
    .D(_0030_),
    .Q_N(_0786_),
    .Q(\ram[5][3] ));
 sg13g2_dfrbp_1 _1668_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net62),
    .D(_0031_),
    .Q_N(_0785_),
    .Q(\ram[5][4] ));
 sg13g2_dfrbp_1 _1669_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net61),
    .D(_0032_),
    .Q_N(_0784_),
    .Q(\ram[5][5] ));
 sg13g2_dfrbp_1 _1670_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net60),
    .D(_0033_),
    .Q_N(_0783_),
    .Q(\ram[5][6] ));
 sg13g2_dfrbp_1 _1671_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net59),
    .D(_0034_),
    .Q_N(_0782_),
    .Q(\ram[5][7] ));
 sg13g2_dfrbp_1 _1672_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net58),
    .D(_0035_),
    .Q_N(_0781_),
    .Q(\ram[14][0] ));
 sg13g2_dfrbp_1 _1673_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net57),
    .D(_0036_),
    .Q_N(_0780_),
    .Q(\ram[14][1] ));
 sg13g2_dfrbp_1 _1674_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net56),
    .D(_0037_),
    .Q_N(_0779_),
    .Q(\ram[14][2] ));
 sg13g2_dfrbp_1 _1675_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net55),
    .D(_0038_),
    .Q_N(_0778_),
    .Q(\ram[14][3] ));
 sg13g2_dfrbp_1 _1676_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net54),
    .D(_0039_),
    .Q_N(_0777_),
    .Q(\ram[14][4] ));
 sg13g2_dfrbp_1 _1677_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net53),
    .D(_0040_),
    .Q_N(_0776_),
    .Q(\ram[14][5] ));
 sg13g2_dfrbp_1 _1678_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net52),
    .D(_0041_),
    .Q_N(_0775_),
    .Q(\ram[14][6] ));
 sg13g2_dfrbp_1 _1679_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net51),
    .D(_0042_),
    .Q_N(_0774_),
    .Q(\ram[14][7] ));
 sg13g2_dfrbp_1 _1680_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net50),
    .D(_0043_),
    .Q_N(_0773_),
    .Q(\ram[4][0] ));
 sg13g2_dfrbp_1 _1681_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net49),
    .D(_0044_),
    .Q_N(_0772_),
    .Q(\ram[4][1] ));
 sg13g2_dfrbp_1 _1682_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net48),
    .D(_0045_),
    .Q_N(_0771_),
    .Q(\ram[4][2] ));
 sg13g2_dfrbp_1 _1683_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net47),
    .D(_0046_),
    .Q_N(_0770_),
    .Q(\ram[4][3] ));
 sg13g2_dfrbp_1 _1684_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net46),
    .D(_0047_),
    .Q_N(_0769_),
    .Q(\ram[4][4] ));
 sg13g2_dfrbp_1 _1685_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net45),
    .D(_0048_),
    .Q_N(_0768_),
    .Q(\ram[4][5] ));
 sg13g2_dfrbp_1 _1686_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net44),
    .D(_0049_),
    .Q_N(_0767_),
    .Q(\ram[4][6] ));
 sg13g2_dfrbp_1 _1687_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net43),
    .D(net180),
    .Q_N(_0766_),
    .Q(\ram[4][7] ));
 sg13g2_dfrbp_1 _1688_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net42),
    .D(_0051_),
    .Q_N(_0765_),
    .Q(\ram[10][0] ));
 sg13g2_dfrbp_1 _1689_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net41),
    .D(_0052_),
    .Q_N(_0764_),
    .Q(\ram[10][1] ));
 sg13g2_dfrbp_1 _1690_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net40),
    .D(_0053_),
    .Q_N(_0763_),
    .Q(\ram[10][2] ));
 sg13g2_dfrbp_1 _1691_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net39),
    .D(_0054_),
    .Q_N(_0762_),
    .Q(\ram[10][3] ));
 sg13g2_dfrbp_1 _1692_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net38),
    .D(_0055_),
    .Q_N(_0761_),
    .Q(\ram[10][4] ));
 sg13g2_dfrbp_1 _1693_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net37),
    .D(_0056_),
    .Q_N(_0760_),
    .Q(\ram[10][5] ));
 sg13g2_dfrbp_1 _1694_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net36),
    .D(_0057_),
    .Q_N(_0759_),
    .Q(\ram[10][6] ));
 sg13g2_dfrbp_1 _1695_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net35),
    .D(_0058_),
    .Q_N(_0758_),
    .Q(\ram[10][7] ));
 sg13g2_dfrbp_1 _1696_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net34),
    .D(_0059_),
    .Q_N(_0757_),
    .Q(\ram[3][0] ));
 sg13g2_dfrbp_1 _1697_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net33),
    .D(_0060_),
    .Q_N(_0756_),
    .Q(\ram[3][1] ));
 sg13g2_dfrbp_1 _1698_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net32),
    .D(_0061_),
    .Q_N(_0755_),
    .Q(\ram[3][2] ));
 sg13g2_dfrbp_1 _1699_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net31),
    .D(_0062_),
    .Q_N(_0754_),
    .Q(\ram[3][3] ));
 sg13g2_dfrbp_1 _1700_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net30),
    .D(_0063_),
    .Q_N(_0753_),
    .Q(\ram[3][4] ));
 sg13g2_dfrbp_1 _1701_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net29),
    .D(_0064_),
    .Q_N(_0752_),
    .Q(\ram[3][5] ));
 sg13g2_dfrbp_1 _1702_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net28),
    .D(_0065_),
    .Q_N(_0751_),
    .Q(\ram[3][6] ));
 sg13g2_dfrbp_1 _1703_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net27),
    .D(net214),
    .Q_N(_0750_),
    .Q(\ram[3][7] ));
 sg13g2_dfrbp_1 _1704_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net26),
    .D(_0067_),
    .Q_N(_0749_),
    .Q(\a[0] ));
 sg13g2_dfrbp_1 _1705_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net24),
    .D(_0068_),
    .Q_N(_0748_),
    .Q(\a[1] ));
 sg13g2_dfrbp_1 _1706_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net22),
    .D(_0069_),
    .Q_N(_0747_),
    .Q(\a[2] ));
 sg13g2_dfrbp_1 _1707_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net20),
    .D(_0070_),
    .Q_N(_0746_),
    .Q(\a[3] ));
 sg13g2_dfrbp_1 _1708_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net18),
    .D(_0071_),
    .Q_N(_0745_),
    .Q(\a[4] ));
 sg13g2_dfrbp_1 _1709_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net16),
    .D(_0072_),
    .Q_N(_0744_),
    .Q(\a[5] ));
 sg13g2_dfrbp_1 _1710_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net14),
    .D(_0073_),
    .Q_N(_0743_),
    .Q(\a[6] ));
 sg13g2_dfrbp_1 _1711_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net150),
    .D(_0074_),
    .Q_N(_0742_),
    .Q(\a[7] ));
 sg13g2_dfrbp_1 _1712_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net148),
    .D(_0075_),
    .Q_N(_0741_),
    .Q(\ram[7][0] ));
 sg13g2_dfrbp_1 _1713_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net147),
    .D(_0076_),
    .Q_N(_0740_),
    .Q(\ram[7][1] ));
 sg13g2_dfrbp_1 _1714_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net146),
    .D(_0077_),
    .Q_N(_0739_),
    .Q(\ram[7][2] ));
 sg13g2_dfrbp_1 _1715_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net145),
    .D(_0078_),
    .Q_N(_0738_),
    .Q(\ram[7][3] ));
 sg13g2_dfrbp_1 _1716_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net144),
    .D(_0079_),
    .Q_N(_0737_),
    .Q(\ram[7][4] ));
 sg13g2_dfrbp_1 _1717_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net143),
    .D(_0080_),
    .Q_N(_0736_),
    .Q(\ram[7][5] ));
 sg13g2_dfrbp_1 _1718_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net142),
    .D(_0081_),
    .Q_N(_0735_),
    .Q(\ram[7][6] ));
 sg13g2_dfrbp_1 _1719_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net141),
    .D(_0082_),
    .Q_N(_0734_),
    .Q(\ram[7][7] ));
 sg13g2_dfrbp_1 _1720_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net140),
    .D(_0083_),
    .Q_N(_0733_),
    .Q(\ram[2][0] ));
 sg13g2_dfrbp_1 _1721_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net139),
    .D(_0084_),
    .Q_N(_0732_),
    .Q(\ram[2][1] ));
 sg13g2_dfrbp_1 _1722_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net138),
    .D(_0085_),
    .Q_N(_0731_),
    .Q(\ram[2][2] ));
 sg13g2_dfrbp_1 _1723_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net137),
    .D(_0086_),
    .Q_N(_0730_),
    .Q(\ram[2][3] ));
 sg13g2_dfrbp_1 _1724_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net136),
    .D(_0087_),
    .Q_N(_0729_),
    .Q(\ram[2][4] ));
 sg13g2_dfrbp_1 _1725_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net135),
    .D(_0088_),
    .Q_N(_0728_),
    .Q(\ram[2][5] ));
 sg13g2_dfrbp_1 _1726_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net134),
    .D(_0089_),
    .Q_N(_0727_),
    .Q(\ram[2][6] ));
 sg13g2_dfrbp_1 _1727_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net133),
    .D(_0090_),
    .Q_N(_0726_),
    .Q(\ram[2][7] ));
 sg13g2_dfrbp_1 _1728_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net132),
    .D(_0091_),
    .Q_N(_0725_),
    .Q(\ram[11][0] ));
 sg13g2_dfrbp_1 _1729_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net131),
    .D(_0092_),
    .Q_N(_0724_),
    .Q(\ram[11][1] ));
 sg13g2_dfrbp_1 _1730_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net130),
    .D(_0093_),
    .Q_N(_0723_),
    .Q(\ram[11][2] ));
 sg13g2_dfrbp_1 _1731_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net129),
    .D(_0094_),
    .Q_N(_0722_),
    .Q(\ram[11][3] ));
 sg13g2_dfrbp_1 _1732_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net128),
    .D(_0095_),
    .Q_N(_0721_),
    .Q(\ram[11][4] ));
 sg13g2_dfrbp_1 _1733_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net127),
    .D(_0096_),
    .Q_N(_0720_),
    .Q(\ram[11][5] ));
 sg13g2_dfrbp_1 _1734_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net126),
    .D(_0097_),
    .Q_N(_0719_),
    .Q(\ram[11][6] ));
 sg13g2_dfrbp_1 _1735_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net125),
    .D(_0098_),
    .Q_N(_0718_),
    .Q(\ram[11][7] ));
 sg13g2_dfrbp_1 _1736_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net124),
    .D(_0099_),
    .Q_N(_0717_),
    .Q(\ram[13][0] ));
 sg13g2_dfrbp_1 _1737_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net123),
    .D(_0100_),
    .Q_N(_0716_),
    .Q(\ram[13][1] ));
 sg13g2_dfrbp_1 _1738_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net122),
    .D(_0101_),
    .Q_N(_0715_),
    .Q(\ram[13][2] ));
 sg13g2_dfrbp_1 _1739_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net121),
    .D(_0102_),
    .Q_N(_0714_),
    .Q(\ram[13][3] ));
 sg13g2_dfrbp_1 _1740_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net120),
    .D(_0103_),
    .Q_N(_0713_),
    .Q(\ram[13][4] ));
 sg13g2_dfrbp_1 _1741_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net119),
    .D(_0104_),
    .Q_N(_0712_),
    .Q(\ram[13][5] ));
 sg13g2_dfrbp_1 _1742_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net118),
    .D(_0105_),
    .Q_N(_0711_),
    .Q(\ram[13][6] ));
 sg13g2_dfrbp_1 _1743_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net117),
    .D(_0106_),
    .Q_N(_0710_),
    .Q(\ram[13][7] ));
 sg13g2_dfrbp_1 _1744_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net116),
    .D(_0107_),
    .Q_N(_0709_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1745_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net115),
    .D(_0108_),
    .Q_N(_0708_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1746_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net114),
    .D(_0109_),
    .Q_N(_0707_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1747_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net113),
    .D(_0110_),
    .Q_N(_0706_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1748_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net112),
    .D(_0111_),
    .Q_N(_0705_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1749_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net111),
    .D(_0112_),
    .Q_N(_0704_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1750_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net110),
    .D(_0113_),
    .Q_N(_0703_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1751_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net109),
    .D(_0114_),
    .Q_N(_0702_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _1752_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net108),
    .D(_0115_),
    .Q_N(_0701_),
    .Q(\ram[12][0] ));
 sg13g2_dfrbp_1 _1753_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net107),
    .D(_0116_),
    .Q_N(_0700_),
    .Q(\ram[12][1] ));
 sg13g2_dfrbp_1 _1754_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net106),
    .D(_0117_),
    .Q_N(_0699_),
    .Q(\ram[12][2] ));
 sg13g2_dfrbp_1 _1755_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net105),
    .D(_0118_),
    .Q_N(_0698_),
    .Q(\ram[12][3] ));
 sg13g2_dfrbp_1 _1756_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net104),
    .D(_0119_),
    .Q_N(_0697_),
    .Q(\ram[12][4] ));
 sg13g2_dfrbp_1 _1757_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net103),
    .D(_0120_),
    .Q_N(_0696_),
    .Q(\ram[12][5] ));
 sg13g2_dfrbp_1 _1758_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net102),
    .D(_0121_),
    .Q_N(_0695_),
    .Q(\ram[12][6] ));
 sg13g2_dfrbp_1 _1759_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net101),
    .D(_0122_),
    .Q_N(_0694_),
    .Q(\ram[12][7] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net100),
    .D(_0123_),
    .Q_N(_0693_),
    .Q(\b[0] ));
 sg13g2_dfrbp_1 _1761_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net99),
    .D(_0124_),
    .Q_N(_0692_),
    .Q(\b[1] ));
 sg13g2_dfrbp_1 _1762_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net98),
    .D(_0125_),
    .Q_N(_0691_),
    .Q(\b[2] ));
 sg13g2_dfrbp_1 _1763_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net97),
    .D(_0126_),
    .Q_N(_0690_),
    .Q(\b[3] ));
 sg13g2_dfrbp_1 _1764_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net96),
    .D(_0127_),
    .Q_N(_0689_),
    .Q(\b[4] ));
 sg13g2_dfrbp_1 _1765_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net95),
    .D(_0128_),
    .Q_N(_0688_),
    .Q(\b[5] ));
 sg13g2_dfrbp_1 _1766_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net94),
    .D(_0129_),
    .Q_N(_0687_),
    .Q(\b[6] ));
 sg13g2_dfrbp_1 _1767_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net93),
    .D(_0130_),
    .Q_N(_0686_),
    .Q(\b[7] ));
 sg13g2_dfrbp_1 _1768_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net92),
    .D(_0131_),
    .Q_N(_0685_),
    .Q(\ram[6][0] ));
 sg13g2_dfrbp_1 _1769_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net25),
    .D(_0132_),
    .Q_N(_0684_),
    .Q(\ram[6][1] ));
 sg13g2_dfrbp_1 _1770_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net23),
    .D(_0133_),
    .Q_N(_0683_),
    .Q(\ram[6][2] ));
 sg13g2_dfrbp_1 _1771_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net21),
    .D(_0134_),
    .Q_N(_0682_),
    .Q(\ram[6][3] ));
 sg13g2_dfrbp_1 _1772_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net19),
    .D(_0135_),
    .Q_N(_0681_),
    .Q(\ram[6][4] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net17),
    .D(_0136_),
    .Q_N(_0680_),
    .Q(\ram[6][5] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net15),
    .D(_0137_),
    .Q_N(_0679_),
    .Q(\ram[6][6] ));
 sg13g2_dfrbp_1 _1775_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net13),
    .D(_0138_),
    .Q_N(_0678_),
    .Q(\ram[6][7] ));
 sg13g2_tiehi _1710__14 (.L_HI(net14));
 sg13g2_tiehi _1774__15 (.L_HI(net15));
 sg13g2_tiehi _1709__16 (.L_HI(net16));
 sg13g2_tiehi _1773__17 (.L_HI(net17));
 sg13g2_tiehi _1708__18 (.L_HI(net18));
 sg13g2_tiehi _1772__19 (.L_HI(net19));
 sg13g2_tiehi _1707__20 (.L_HI(net20));
 sg13g2_tiehi _1771__21 (.L_HI(net21));
 sg13g2_tiehi _1706__22 (.L_HI(net22));
 sg13g2_tiehi _1770__23 (.L_HI(net23));
 sg13g2_tiehi _1705__24 (.L_HI(net24));
 sg13g2_tiehi _1769__25 (.L_HI(net25));
 sg13g2_tiehi _1704__26 (.L_HI(net26));
 sg13g2_tiehi _1703__27 (.L_HI(net27));
 sg13g2_tiehi _1702__28 (.L_HI(net28));
 sg13g2_tiehi _1701__29 (.L_HI(net29));
 sg13g2_tiehi _1700__30 (.L_HI(net30));
 sg13g2_tiehi _1699__31 (.L_HI(net31));
 sg13g2_tiehi _1698__32 (.L_HI(net32));
 sg13g2_tiehi _1697__33 (.L_HI(net33));
 sg13g2_tiehi _1696__34 (.L_HI(net34));
 sg13g2_tiehi _1695__35 (.L_HI(net35));
 sg13g2_tiehi _1694__36 (.L_HI(net36));
 sg13g2_tiehi _1693__37 (.L_HI(net37));
 sg13g2_tiehi _1692__38 (.L_HI(net38));
 sg13g2_tiehi _1691__39 (.L_HI(net39));
 sg13g2_tiehi _1690__40 (.L_HI(net40));
 sg13g2_tiehi _1689__41 (.L_HI(net41));
 sg13g2_tiehi _1688__42 (.L_HI(net42));
 sg13g2_tiehi _1687__43 (.L_HI(net43));
 sg13g2_tiehi _1686__44 (.L_HI(net44));
 sg13g2_tiehi _1685__45 (.L_HI(net45));
 sg13g2_tiehi _1684__46 (.L_HI(net46));
 sg13g2_tiehi _1683__47 (.L_HI(net47));
 sg13g2_tiehi _1682__48 (.L_HI(net48));
 sg13g2_tiehi _1681__49 (.L_HI(net49));
 sg13g2_tiehi _1680__50 (.L_HI(net50));
 sg13g2_tiehi _1679__51 (.L_HI(net51));
 sg13g2_tiehi _1678__52 (.L_HI(net52));
 sg13g2_tiehi _1677__53 (.L_HI(net53));
 sg13g2_tiehi _1676__54 (.L_HI(net54));
 sg13g2_tiehi _1675__55 (.L_HI(net55));
 sg13g2_tiehi _1674__56 (.L_HI(net56));
 sg13g2_tiehi _1673__57 (.L_HI(net57));
 sg13g2_tiehi _1672__58 (.L_HI(net58));
 sg13g2_tiehi _1671__59 (.L_HI(net59));
 sg13g2_tiehi _1670__60 (.L_HI(net60));
 sg13g2_tiehi _1669__61 (.L_HI(net61));
 sg13g2_tiehi _1668__62 (.L_HI(net62));
 sg13g2_tiehi _1667__63 (.L_HI(net63));
 sg13g2_tiehi _1666__64 (.L_HI(net64));
 sg13g2_tiehi _1665__65 (.L_HI(net65));
 sg13g2_tiehi _1664__66 (.L_HI(net66));
 sg13g2_tiehi _1663__67 (.L_HI(net67));
 sg13g2_tiehi _1662__68 (.L_HI(net68));
 sg13g2_tiehi _1661__69 (.L_HI(net69));
 sg13g2_tiehi _1660__70 (.L_HI(net70));
 sg13g2_tiehi _1659__71 (.L_HI(net71));
 sg13g2_tiehi _1658__72 (.L_HI(net72));
 sg13g2_tiehi _1657__73 (.L_HI(net73));
 sg13g2_tiehi _1656__74 (.L_HI(net74));
 sg13g2_tiehi _1655__75 (.L_HI(net75));
 sg13g2_tiehi _1654__76 (.L_HI(net76));
 sg13g2_tiehi _1653__77 (.L_HI(net77));
 sg13g2_tiehi _1652__78 (.L_HI(net78));
 sg13g2_tiehi _1651__79 (.L_HI(net79));
 sg13g2_tiehi _1650__80 (.L_HI(net80));
 sg13g2_tiehi _1649__81 (.L_HI(net81));
 sg13g2_tiehi _1648__82 (.L_HI(net82));
 sg13g2_tiehi _1647__83 (.L_HI(net83));
 sg13g2_tiehi _1646__84 (.L_HI(net84));
 sg13g2_tiehi _1645__85 (.L_HI(net85));
 sg13g2_tiehi _1644__86 (.L_HI(net86));
 sg13g2_tiehi _1643__87 (.L_HI(net87));
 sg13g2_tiehi _1642__88 (.L_HI(net88));
 sg13g2_tiehi _1641__89 (.L_HI(net89));
 sg13g2_tiehi _1640__90 (.L_HI(net90));
 sg13g2_tiehi _1639__91 (.L_HI(net91));
 sg13g2_tiehi _1768__92 (.L_HI(net92));
 sg13g2_tiehi _1767__93 (.L_HI(net93));
 sg13g2_tiehi _1766__94 (.L_HI(net94));
 sg13g2_tiehi _1765__95 (.L_HI(net95));
 sg13g2_tiehi _1764__96 (.L_HI(net96));
 sg13g2_tiehi _1763__97 (.L_HI(net97));
 sg13g2_tiehi _1762__98 (.L_HI(net98));
 sg13g2_tiehi _1761__99 (.L_HI(net99));
 sg13g2_tiehi _1760__100 (.L_HI(net100));
 sg13g2_tiehi _1759__101 (.L_HI(net101));
 sg13g2_tiehi _1758__102 (.L_HI(net102));
 sg13g2_tiehi _1757__103 (.L_HI(net103));
 sg13g2_tiehi _1756__104 (.L_HI(net104));
 sg13g2_tiehi _1755__105 (.L_HI(net105));
 sg13g2_tiehi _1754__106 (.L_HI(net106));
 sg13g2_tiehi _1753__107 (.L_HI(net107));
 sg13g2_tiehi _1752__108 (.L_HI(net108));
 sg13g2_tiehi _1751__109 (.L_HI(net109));
 sg13g2_tiehi _1750__110 (.L_HI(net110));
 sg13g2_tiehi _1749__111 (.L_HI(net111));
 sg13g2_tiehi _1748__112 (.L_HI(net112));
 sg13g2_tiehi _1747__113 (.L_HI(net113));
 sg13g2_tiehi _1746__114 (.L_HI(net114));
 sg13g2_tiehi _1745__115 (.L_HI(net115));
 sg13g2_tiehi _1744__116 (.L_HI(net116));
 sg13g2_tiehi _1743__117 (.L_HI(net117));
 sg13g2_tiehi _1742__118 (.L_HI(net118));
 sg13g2_tiehi _1741__119 (.L_HI(net119));
 sg13g2_tiehi _1740__120 (.L_HI(net120));
 sg13g2_tiehi _1739__121 (.L_HI(net121));
 sg13g2_tiehi _1738__122 (.L_HI(net122));
 sg13g2_tiehi _1737__123 (.L_HI(net123));
 sg13g2_tiehi _1736__124 (.L_HI(net124));
 sg13g2_tiehi _1735__125 (.L_HI(net125));
 sg13g2_tiehi _1734__126 (.L_HI(net126));
 sg13g2_tiehi _1733__127 (.L_HI(net127));
 sg13g2_tiehi _1732__128 (.L_HI(net128));
 sg13g2_tiehi _1731__129 (.L_HI(net129));
 sg13g2_tiehi _1730__130 (.L_HI(net130));
 sg13g2_tiehi _1729__131 (.L_HI(net131));
 sg13g2_tiehi _1728__132 (.L_HI(net132));
 sg13g2_tiehi _1727__133 (.L_HI(net133));
 sg13g2_tiehi _1726__134 (.L_HI(net134));
 sg13g2_tiehi _1725__135 (.L_HI(net135));
 sg13g2_tiehi _1724__136 (.L_HI(net136));
 sg13g2_tiehi _1723__137 (.L_HI(net137));
 sg13g2_tiehi _1722__138 (.L_HI(net138));
 sg13g2_tiehi _1721__139 (.L_HI(net139));
 sg13g2_tiehi _1720__140 (.L_HI(net140));
 sg13g2_tiehi _1719__141 (.L_HI(net141));
 sg13g2_tiehi _1718__142 (.L_HI(net142));
 sg13g2_tiehi _1717__143 (.L_HI(net143));
 sg13g2_tiehi _1716__144 (.L_HI(net144));
 sg13g2_tiehi _1715__145 (.L_HI(net145));
 sg13g2_tiehi _1714__146 (.L_HI(net146));
 sg13g2_tiehi _1713__147 (.L_HI(net147));
 sg13g2_tiehi _1712__148 (.L_HI(net148));
 sg13g2_tiehi _1638__149 (.L_HI(net149));
 sg13g2_tiehi _1711__150 (.L_HI(net150));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _1914_ (.A(ui_in[6]),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1915_ (.A(ui_in[6]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1916_ (.A(ui_in[6]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1917_ (.A(ui_in[6]),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1918_ (.A(ui_in[6]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1919_ (.A(ui_in[6]),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1920_ (.A(ui_in[6]),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1921_ (.A(ui_in[6]),
    .X(uio_oe[7]));
 sg13g2_buf_2 fanout245 (.A(net246),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_0651_),
    .X(net246));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(_0465_));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(_0455_));
 sg13g2_buf_2 fanout249 (.A(_0455_),
    .X(net249));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(net251));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(_0419_));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(_0350_));
 sg13g2_buf_2 fanout253 (.A(_0350_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_0178_),
    .X(net254));
 sg13g2_buf_1 fanout255 (.A(_0178_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(net257),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_0661_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net259),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_0502_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(net261),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_0492_),
    .X(net261));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(_0476_));
 sg13g2_buf_2 fanout263 (.A(_0476_),
    .X(net263));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_0454_));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_0454_));
 sg13g2_buf_2 fanout266 (.A(net267),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_0445_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(net269),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_0428_),
    .X(net269));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(net271));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_0418_));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(_0349_));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_0349_));
 sg13g2_buf_2 fanout274 (.A(net275),
    .X(net274));
 sg13g2_buf_1 fanout275 (.A(_0176_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_0151_),
    .X(net276));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(_0475_));
 sg13g2_buf_2 fanout278 (.A(_0475_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_0331_),
    .X(net280));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(net283));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(net283));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_0159_));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_0150_));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(net286));
 sg13g2_buf_2 fanout286 (.A(\b[7] ),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(\a[7] ),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_0328_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_0328_),
    .X(net290));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(_0139_));
 sg13g2_buf_2 fanout292 (.A(net293),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net2),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(net295),
    .X(net294));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(net1));
 sg13g2_buf_2 fanout296 (.A(net298),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(net298),
    .X(net297));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(net1));
 sg13g2_buf_4 fanout299 (.X(net299),
    .A(net301));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(net301));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(net306));
 sg13g2_buf_4 fanout302 (.X(net302),
    .A(net305));
 sg13g2_buf_2 fanout303 (.A(net304),
    .X(net303));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(net305));
 sg13g2_buf_2 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(ui_in[1]),
    .X(net306));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(net310));
 sg13g2_buf_2 fanout308 (.A(net310),
    .X(net308));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(net310));
 sg13g2_buf_2 fanout310 (.A(net318),
    .X(net310));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(net318));
 sg13g2_buf_2 fanout312 (.A(net318),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net314),
    .X(net313));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(net318));
 sg13g2_buf_2 fanout315 (.A(net316),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(net318));
 sg13g2_buf_2 fanout318 (.A(ui_in[0]),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net320),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(net321),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(rst_n),
    .X(net321));
 sg13g2_buf_2 input1 (.A(ui_in[2]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[7]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[0]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[1]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[2]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[3]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[4]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[5]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[6]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[7]),
    .X(net12));
 sg13g2_tiehi _1775__13 (.L_HI(net13));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_29__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0000_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ram[13][6] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold3 (.A(\ram[0][1] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold4 (.A(\ram[0][5] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold5 (.A(\ram[6][1] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold6 (.A(\ram[0][3] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold7 (.A(\ram[2][7] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold8 (.A(\ram[5][0] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold9 (.A(\ram[13][4] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold10 (.A(\ram[0][7] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0018_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold12 (.A(\ram[13][0] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold13 (.A(\ram[13][2] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold14 (.A(\ram[4][1] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold15 (.A(\ram[7][5] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold16 (.A(\ram[13][7] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold17 (.A(\ram[5][2] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold18 (.A(\ram[6][7] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold19 (.A(\ram[13][3] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold20 (.A(\ram[6][2] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold21 (.A(\ram[7][2] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold22 (.A(\ram[1][3] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold23 (.A(\ram[4][0] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold24 (.A(\ram[4][5] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold25 (.A(\ram[0][4] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ram[6][6] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold27 (.A(\ram[7][3] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold28 (.A(\ram[0][0] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold29 (.A(\ram[4][7] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0050_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold31 (.A(\ram[1][4] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold32 (.A(\ram[15][2] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold33 (.A(\ram[0][6] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ram[3][2] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold35 (.A(\ram[5][1] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold36 (.A(\ram[4][6] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold37 (.A(\ram[7][1] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold38 (.A(\ram[14][4] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold39 (.A(\ram[4][2] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold40 (.A(\ram[2][6] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold41 (.A(\ram[2][5] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold42 (.A(\ram[3][0] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold43 (.A(\ram[3][3] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold44 (.A(\ram[5][6] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold45 (.A(\ram[13][5] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold46 (.A(\ram[1][7] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold47 (.A(\ram[3][4] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold48 (.A(\ram[6][0] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold49 (.A(\ram[3][5] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold50 (.A(\ram[2][1] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold51 (.A(\ram[5][7] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ram[7][4] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold53 (.A(\ram[5][3] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ram[6][4] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold55 (.A(\ram[13][1] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold56 (.A(\ram[2][3] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold57 (.A(\ram[15][1] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold58 (.A(\ram[3][6] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold59 (.A(\ram[2][4] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold60 (.A(\ram[1][0] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold61 (.A(\ram[7][0] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ram[14][5] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold63 (.A(\ram[3][7] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0066_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold65 (.A(\ram[15][0] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold66 (.A(\ram[5][4] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold67 (.A(\ram[14][3] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold68 (.A(\ram[15][6] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold69 (.A(\ram[5][5] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold70 (.A(\ram[14][1] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ram[1][1] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold72 (.A(\ram[15][4] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ram[15][3] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold74 (.A(\ram[1][5] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold75 (.A(\ram[6][5] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold76 (.A(\ram[2][2] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold77 (.A(\ram[14][2] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold78 (.A(\ram[4][3] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold79 (.A(\ram[6][3] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold80 (.A(\ram[1][2] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold81 (.A(\ram[15][5] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold82 (.A(\ram[1][6] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold83 (.A(\ram[12][4] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold84 (.A(\ram[10][0] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold85 (.A(\ram[4][4] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold86 (.A(\ram[2][0] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold87 (.A(\ram[11][0] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold88 (.A(\ram[15][7] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold89 (.A(\ram[10][2] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold90 (.A(\ram[10][1] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold91 (.A(\ram[10][3] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold92 (.A(\ram[3][1] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold93 (.A(\ram[11][6] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold94 (.A(\ram[10][5] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold95 (.A(\ram[11][3] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold96 (.A(\ram[11][2] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold97 (.A(\ram[10][4] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold98 (.A(\ram[12][1] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold99 (.A(\ram[14][7] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold100 (.A(\ram[14][6] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold101 (.A(\ram[0][2] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold102 (.A(\ram[14][0] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold103 (.A(\ram[12][7] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold104 (.A(\ram[12][3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold105 (.A(\ram[11][1] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold106 (.A(\ram[11][5] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold107 (.A(\ram[10][6] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold108 (.A(\ram[7][7] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold109 (.A(\ram[11][4] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold110 (.A(\ram[12][0] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold111 (.A(\ram[10][7] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold112 (.A(\ram[12][2] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold113 (.A(\ram[12][6] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold114 (.A(\ram[12][5] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold115 (.A(\ram[11][7] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold116 (.A(\a[3] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold117 (.A(\ram[7][6] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold118 (.A(\b[3] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold119 (.A(\a[5] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold120 (.A(\a[1] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold121 (.A(\b[5] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold122 (.A(\a[0] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold123 (.A(\b[1] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold124 (.A(\b[0] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold125 (.A(\a[4] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold126 (.A(\b[4] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold127 (.A(\a[2] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold128 (.A(\b[2] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold129 (.A(\a[6] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold130 (.A(\b[6] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold131 (.A(\result_addr[0] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0348_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold133 (.A(\result_addr[0] ),
    .X(net360));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_fill_2 FILLER_7_175 ();
 sg13g2_fill_1 FILLER_7_177 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_fill_2 FILLER_7_245 ();
 sg13g2_fill_1 FILLER_7_247 ();
 sg13g2_decap_8 FILLER_7_253 ();
 sg13g2_decap_8 FILLER_7_260 ();
 sg13g2_decap_4 FILLER_7_267 ();
 sg13g2_fill_2 FILLER_7_271 ();
 sg13g2_decap_8 FILLER_7_281 ();
 sg13g2_decap_8 FILLER_7_288 ();
 sg13g2_decap_8 FILLER_7_295 ();
 sg13g2_decap_8 FILLER_7_302 ();
 sg13g2_decap_8 FILLER_7_309 ();
 sg13g2_decap_8 FILLER_7_316 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_decap_8 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_351 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_4 FILLER_8_162 ();
 sg13g2_fill_2 FILLER_8_166 ();
 sg13g2_decap_4 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_201 ();
 sg13g2_decap_4 FILLER_8_208 ();
 sg13g2_fill_1 FILLER_8_212 ();
 sg13g2_decap_8 FILLER_8_229 ();
 sg13g2_fill_1 FILLER_8_236 ();
 sg13g2_fill_1 FILLER_8_243 ();
 sg13g2_decap_4 FILLER_8_264 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_176 ();
 sg13g2_decap_8 FILLER_9_180 ();
 sg13g2_fill_2 FILLER_9_187 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_fill_1 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_28 ();
 sg13g2_fill_1 FILLER_10_33 ();
 sg13g2_decap_8 FILLER_10_38 ();
 sg13g2_decap_8 FILLER_10_45 ();
 sg13g2_decap_8 FILLER_10_52 ();
 sg13g2_fill_2 FILLER_10_59 ();
 sg13g2_decap_4 FILLER_10_87 ();
 sg13g2_decap_4 FILLER_10_95 ();
 sg13g2_fill_2 FILLER_10_99 ();
 sg13g2_fill_1 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_114 ();
 sg13g2_decap_8 FILLER_10_121 ();
 sg13g2_decap_8 FILLER_10_132 ();
 sg13g2_decap_8 FILLER_10_139 ();
 sg13g2_fill_1 FILLER_10_146 ();
 sg13g2_decap_4 FILLER_10_155 ();
 sg13g2_decap_4 FILLER_10_172 ();
 sg13g2_fill_2 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_183 ();
 sg13g2_decap_8 FILLER_10_206 ();
 sg13g2_fill_2 FILLER_10_213 ();
 sg13g2_fill_1 FILLER_10_215 ();
 sg13g2_decap_4 FILLER_10_229 ();
 sg13g2_fill_2 FILLER_10_233 ();
 sg13g2_decap_4 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_245 ();
 sg13g2_decap_4 FILLER_10_266 ();
 sg13g2_fill_1 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_4 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_44 ();
 sg13g2_fill_2 FILLER_11_51 ();
 sg13g2_fill_1 FILLER_11_53 ();
 sg13g2_fill_2 FILLER_11_63 ();
 sg13g2_decap_4 FILLER_11_156 ();
 sg13g2_decap_8 FILLER_11_192 ();
 sg13g2_fill_2 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_201 ();
 sg13g2_fill_1 FILLER_11_215 ();
 sg13g2_decap_4 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_244 ();
 sg13g2_fill_2 FILLER_11_250 ();
 sg13g2_fill_1 FILLER_11_257 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_fill_1 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_289 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_fill_1 FILLER_12_26 ();
 sg13g2_fill_2 FILLER_12_94 ();
 sg13g2_fill_1 FILLER_12_101 ();
 sg13g2_fill_2 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_113 ();
 sg13g2_fill_2 FILLER_12_128 ();
 sg13g2_decap_4 FILLER_12_156 ();
 sg13g2_fill_2 FILLER_12_160 ();
 sg13g2_fill_2 FILLER_12_170 ();
 sg13g2_fill_1 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_178 ();
 sg13g2_fill_1 FILLER_12_210 ();
 sg13g2_decap_4 FILLER_12_216 ();
 sg13g2_fill_1 FILLER_12_220 ();
 sg13g2_fill_2 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_235 ();
 sg13g2_fill_1 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_293 ();
 sg13g2_decap_8 FILLER_12_300 ();
 sg13g2_decap_8 FILLER_12_307 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_19 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_fill_1 FILLER_13_53 ();
 sg13g2_decap_4 FILLER_13_59 ();
 sg13g2_fill_1 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_74 ();
 sg13g2_fill_1 FILLER_13_76 ();
 sg13g2_fill_2 FILLER_13_96 ();
 sg13g2_decap_4 FILLER_13_160 ();
 sg13g2_fill_1 FILLER_13_164 ();
 sg13g2_fill_1 FILLER_13_170 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_fill_2 FILLER_13_207 ();
 sg13g2_fill_1 FILLER_13_209 ();
 sg13g2_decap_8 FILLER_13_241 ();
 sg13g2_fill_2 FILLER_13_248 ();
 sg13g2_decap_4 FILLER_13_254 ();
 sg13g2_fill_1 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_fill_2 FILLER_13_281 ();
 sg13g2_fill_1 FILLER_13_283 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_41 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_fill_1 FILLER_14_113 ();
 sg13g2_fill_2 FILLER_14_128 ();
 sg13g2_decap_8 FILLER_14_134 ();
 sg13g2_fill_1 FILLER_14_141 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_fill_1 FILLER_14_158 ();
 sg13g2_decap_4 FILLER_14_164 ();
 sg13g2_fill_2 FILLER_14_176 ();
 sg13g2_fill_1 FILLER_14_178 ();
 sg13g2_decap_4 FILLER_14_197 ();
 sg13g2_fill_2 FILLER_14_201 ();
 sg13g2_decap_4 FILLER_14_212 ();
 sg13g2_fill_1 FILLER_14_216 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_fill_2 FILLER_14_244 ();
 sg13g2_fill_1 FILLER_14_246 ();
 sg13g2_decap_8 FILLER_14_256 ();
 sg13g2_fill_2 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_283 ();
 sg13g2_decap_8 FILLER_14_316 ();
 sg13g2_decap_4 FILLER_14_323 ();
 sg13g2_fill_2 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_24 ();
 sg13g2_decap_4 FILLER_15_30 ();
 sg13g2_fill_2 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_77 ();
 sg13g2_fill_2 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_85 ();
 sg13g2_fill_2 FILLER_15_103 ();
 sg13g2_fill_1 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_128 ();
 sg13g2_fill_2 FILLER_15_135 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_176 ();
 sg13g2_fill_1 FILLER_15_194 ();
 sg13g2_decap_8 FILLER_15_227 ();
 sg13g2_fill_1 FILLER_15_243 ();
 sg13g2_fill_2 FILLER_15_261 ();
 sg13g2_fill_1 FILLER_15_263 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_fill_2 FILLER_15_293 ();
 sg13g2_fill_2 FILLER_15_300 ();
 sg13g2_fill_2 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_32 ();
 sg13g2_fill_1 FILLER_16_37 ();
 sg13g2_fill_1 FILLER_16_58 ();
 sg13g2_fill_1 FILLER_16_81 ();
 sg13g2_fill_1 FILLER_16_136 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_fill_1 FILLER_16_172 ();
 sg13g2_fill_2 FILLER_16_187 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_195 ();
 sg13g2_decap_8 FILLER_16_202 ();
 sg13g2_fill_2 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_211 ();
 sg13g2_decap_8 FILLER_16_225 ();
 sg13g2_fill_1 FILLER_16_232 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_decap_4 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_311 ();
 sg13g2_fill_1 FILLER_16_317 ();
 sg13g2_fill_1 FILLER_16_353 ();
 sg13g2_fill_2 FILLER_16_394 ();
 sg13g2_fill_1 FILLER_16_396 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_15 ();
 sg13g2_fill_2 FILLER_17_22 ();
 sg13g2_fill_1 FILLER_17_24 ();
 sg13g2_fill_2 FILLER_17_51 ();
 sg13g2_fill_1 FILLER_17_79 ();
 sg13g2_decap_8 FILLER_17_136 ();
 sg13g2_fill_1 FILLER_17_143 ();
 sg13g2_decap_4 FILLER_17_158 ();
 sg13g2_fill_2 FILLER_17_166 ();
 sg13g2_fill_1 FILLER_17_186 ();
 sg13g2_decap_8 FILLER_17_229 ();
 sg13g2_decap_8 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_4 FILLER_17_294 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_fill_1 FILLER_17_308 ();
 sg13g2_fill_1 FILLER_17_313 ();
 sg13g2_fill_1 FILLER_17_332 ();
 sg13g2_fill_2 FILLER_17_380 ();
 sg13g2_fill_1 FILLER_17_382 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_44 ();
 sg13g2_decap_8 FILLER_18_75 ();
 sg13g2_fill_1 FILLER_18_82 ();
 sg13g2_fill_2 FILLER_18_97 ();
 sg13g2_fill_2 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_127 ();
 sg13g2_fill_1 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_4 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_239 ();
 sg13g2_fill_2 FILLER_18_251 ();
 sg13g2_decap_8 FILLER_18_257 ();
 sg13g2_fill_2 FILLER_18_264 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_fill_2 FILLER_18_285 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_fill_2 FILLER_18_376 ();
 sg13g2_fill_1 FILLER_18_378 ();
 sg13g2_fill_1 FILLER_18_392 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_35 ();
 sg13g2_fill_1 FILLER_19_84 ();
 sg13g2_fill_2 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_122 ();
 sg13g2_fill_1 FILLER_19_124 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_4 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_185 ();
 sg13g2_decap_8 FILLER_19_192 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_decap_4 FILLER_19_204 ();
 sg13g2_fill_1 FILLER_19_208 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_310 ();
 sg13g2_fill_1 FILLER_19_312 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_fill_2 FILLER_19_366 ();
 sg13g2_fill_1 FILLER_19_368 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_decap_4 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_170 ();
 sg13g2_fill_1 FILLER_20_188 ();
 sg13g2_fill_1 FILLER_20_215 ();
 sg13g2_decap_4 FILLER_20_237 ();
 sg13g2_fill_2 FILLER_20_241 ();
 sg13g2_decap_8 FILLER_20_247 ();
 sg13g2_decap_4 FILLER_20_254 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_decap_4 FILLER_20_280 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_decap_4 FILLER_20_289 ();
 sg13g2_fill_1 FILLER_20_293 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_fill_1 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_342 ();
 sg13g2_fill_2 FILLER_20_374 ();
 sg13g2_fill_1 FILLER_20_376 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_21_47 ();
 sg13g2_fill_1 FILLER_21_49 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_fill_2 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_fill_2 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_decap_4 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_decap_4 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_240 ();
 sg13g2_decap_8 FILLER_21_260 ();
 sg13g2_decap_8 FILLER_21_267 ();
 sg13g2_decap_4 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_336 ();
 sg13g2_fill_1 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_26 ();
 sg13g2_fill_1 FILLER_22_32 ();
 sg13g2_fill_2 FILLER_22_51 ();
 sg13g2_fill_2 FILLER_22_115 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_decap_4 FILLER_22_132 ();
 sg13g2_fill_2 FILLER_22_145 ();
 sg13g2_fill_2 FILLER_22_151 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_decap_8 FILLER_22_181 ();
 sg13g2_decap_8 FILLER_22_188 ();
 sg13g2_fill_2 FILLER_22_195 ();
 sg13g2_decap_4 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_205 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_fill_2 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_fill_2 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_296 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_fill_2 FILLER_22_370 ();
 sg13g2_fill_2 FILLER_22_381 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_30 ();
 sg13g2_decap_8 FILLER_23_62 ();
 sg13g2_fill_2 FILLER_23_69 ();
 sg13g2_decap_4 FILLER_23_75 ();
 sg13g2_decap_8 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_115 ();
 sg13g2_decap_4 FILLER_23_121 ();
 sg13g2_fill_2 FILLER_23_138 ();
 sg13g2_fill_1 FILLER_23_140 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_174 ();
 sg13g2_decap_4 FILLER_23_206 ();
 sg13g2_fill_1 FILLER_23_236 ();
 sg13g2_decap_4 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_2 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_311 ();
 sg13g2_fill_2 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_31 ();
 sg13g2_fill_2 FILLER_24_40 ();
 sg13g2_fill_1 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_47 ();
 sg13g2_fill_2 FILLER_24_52 ();
 sg13g2_fill_1 FILLER_24_54 ();
 sg13g2_fill_1 FILLER_24_108 ();
 sg13g2_fill_2 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_decap_8 FILLER_24_148 ();
 sg13g2_fill_2 FILLER_24_155 ();
 sg13g2_decap_4 FILLER_24_161 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_fill_1 FILLER_24_177 ();
 sg13g2_decap_4 FILLER_24_183 ();
 sg13g2_fill_1 FILLER_24_187 ();
 sg13g2_fill_2 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_279 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_301 ();
 sg13g2_fill_2 FILLER_24_342 ();
 sg13g2_fill_2 FILLER_24_374 ();
 sg13g2_fill_1 FILLER_24_376 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_4 FILLER_25_39 ();
 sg13g2_fill_1 FILLER_25_48 ();
 sg13g2_decap_4 FILLER_25_62 ();
 sg13g2_fill_1 FILLER_25_73 ();
 sg13g2_decap_4 FILLER_25_114 ();
 sg13g2_fill_2 FILLER_25_118 ();
 sg13g2_fill_2 FILLER_25_124 ();
 sg13g2_decap_4 FILLER_25_160 ();
 sg13g2_fill_2 FILLER_25_164 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_242 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_decap_4 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_337 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_fill_2 FILLER_25_359 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_fill_2 FILLER_25_367 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_9 ();
 sg13g2_fill_1 FILLER_26_49 ();
 sg13g2_fill_1 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_82 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_fill_2 FILLER_26_195 ();
 sg13g2_decap_8 FILLER_26_202 ();
 sg13g2_decap_4 FILLER_26_209 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_fill_2 FILLER_26_222 ();
 sg13g2_fill_2 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_decap_8 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_decap_4 FILLER_26_334 ();
 sg13g2_fill_1 FILLER_26_338 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_31 ();
 sg13g2_fill_2 FILLER_27_45 ();
 sg13g2_fill_1 FILLER_27_56 ();
 sg13g2_fill_2 FILLER_27_76 ();
 sg13g2_fill_2 FILLER_27_83 ();
 sg13g2_decap_8 FILLER_27_101 ();
 sg13g2_fill_2 FILLER_27_108 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_146 ();
 sg13g2_fill_2 FILLER_27_152 ();
 sg13g2_fill_2 FILLER_27_171 ();
 sg13g2_fill_2 FILLER_27_186 ();
 sg13g2_decap_4 FILLER_27_192 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_decap_4 FILLER_27_307 ();
 sg13g2_fill_2 FILLER_27_317 ();
 sg13g2_fill_1 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_fill_1 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_fill_1 FILLER_28_72 ();
 sg13g2_fill_2 FILLER_28_119 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_176 ();
 sg13g2_decap_4 FILLER_28_203 ();
 sg13g2_fill_1 FILLER_28_207 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_fill_2 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_230 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_decap_4 FILLER_28_238 ();
 sg13g2_fill_2 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_fill_2 FILLER_28_387 ();
 sg13g2_fill_1 FILLER_28_389 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_160 ();
 sg13g2_decap_8 FILLER_29_166 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_fill_2 FILLER_29_184 ();
 sg13g2_fill_1 FILLER_29_186 ();
 sg13g2_decap_4 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_195 ();
 sg13g2_decap_4 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_fill_1 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_fill_1 FILLER_29_294 ();
 sg13g2_fill_1 FILLER_29_371 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_30_39 ();
 sg13g2_fill_2 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_59 ();
 sg13g2_fill_1 FILLER_30_109 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_2 FILLER_30_138 ();
 sg13g2_fill_1 FILLER_30_140 ();
 sg13g2_decap_4 FILLER_30_172 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_decap_8 FILLER_30_218 ();
 sg13g2_decap_4 FILLER_30_225 ();
 sg13g2_fill_2 FILLER_30_255 ();
 sg13g2_fill_1 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_276 ();
 sg13g2_fill_1 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_343 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_392 ();
 sg13g2_fill_1 FILLER_30_398 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_fill_2 FILLER_31_80 ();
 sg13g2_fill_1 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_fill_2 FILLER_31_149 ();
 sg13g2_fill_2 FILLER_31_164 ();
 sg13g2_decap_8 FILLER_31_187 ();
 sg13g2_fill_2 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_196 ();
 sg13g2_decap_4 FILLER_31_227 ();
 sg13g2_decap_4 FILLER_31_236 ();
 sg13g2_fill_2 FILLER_31_240 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_fill_2 FILLER_31_332 ();
 sg13g2_fill_2 FILLER_31_360 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_fill_1 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_89 ();
 sg13g2_decap_4 FILLER_32_131 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_fill_2 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_decap_4 FILLER_32_210 ();
 sg13g2_decap_4 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_268 ();
 sg13g2_fill_2 FILLER_32_295 ();
 sg13g2_fill_2 FILLER_32_315 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_31 ();
 sg13g2_fill_1 FILLER_33_41 ();
 sg13g2_fill_1 FILLER_33_47 ();
 sg13g2_fill_2 FILLER_33_57 ();
 sg13g2_fill_1 FILLER_33_59 ();
 sg13g2_fill_2 FILLER_33_65 ();
 sg13g2_fill_1 FILLER_33_67 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_fill_1 FILLER_33_130 ();
 sg13g2_decap_4 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_decap_4 FILLER_33_234 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_fill_1 FILLER_33_315 ();
 sg13g2_fill_2 FILLER_33_361 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_fill_2 FILLER_33_384 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_48 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_152 ();
 sg13g2_fill_1 FILLER_34_208 ();
 sg13g2_fill_1 FILLER_34_218 ();
 sg13g2_decap_4 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_fill_2 FILLER_34_242 ();
 sg13g2_fill_1 FILLER_34_244 ();
 sg13g2_fill_2 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_280 ();
 sg13g2_fill_2 FILLER_34_337 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_fill_2 FILLER_35_43 ();
 sg13g2_fill_1 FILLER_35_45 ();
 sg13g2_fill_2 FILLER_35_56 ();
 sg13g2_fill_1 FILLER_35_58 ();
 sg13g2_fill_1 FILLER_35_93 ();
 sg13g2_fill_1 FILLER_35_120 ();
 sg13g2_decap_4 FILLER_35_152 ();
 sg13g2_fill_1 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_2 FILLER_35_353 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_86 ();
 sg13g2_fill_1 FILLER_36_88 ();
 sg13g2_fill_2 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_136 ();
 sg13g2_decap_4 FILLER_36_141 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_4 FILLER_36_203 ();
 sg13g2_fill_2 FILLER_36_229 ();
 sg13g2_decap_4 FILLER_36_235 ();
 sg13g2_fill_2 FILLER_36_239 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_fill_2 FILLER_36_281 ();
 sg13g2_fill_2 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_fill_1 FILLER_36_386 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_1 FILLER_37_15 ();
 sg13g2_fill_1 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_66 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_100 ();
 sg13g2_fill_2 FILLER_37_162 ();
 sg13g2_fill_1 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_187 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_fill_1 FILLER_37_295 ();
 sg13g2_fill_2 FILLER_37_320 ();
 sg13g2_fill_1 FILLER_37_322 ();
 sg13g2_fill_2 FILLER_37_357 ();
 sg13g2_fill_1 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_15 ();
 sg13g2_fill_2 FILLER_38_19 ();
 sg13g2_fill_1 FILLER_38_26 ();
 sg13g2_fill_1 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_71 ();
 sg13g2_fill_1 FILLER_38_137 ();
 sg13g2_fill_2 FILLER_38_151 ();
 sg13g2_decap_4 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_218 ();
 sg13g2_decap_4 FILLER_38_225 ();
 sg13g2_fill_1 FILLER_38_229 ();
 sg13g2_fill_2 FILLER_38_238 ();
 sg13g2_fill_2 FILLER_38_260 ();
 sg13g2_fill_1 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_407 ();
endmodule

module tt_um_algofoogle_tt09_ring_osc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire dummy;
 wire \myring.inv_in[0] ;
 wire \myring.inv_in[1000] ;
 wire \myring.inv_in[100] ;
 wire \myring.inv_in[101] ;
 wire \myring.inv_in[102] ;
 wire \myring.inv_in[103] ;
 wire \myring.inv_in[104] ;
 wire \myring.inv_in[105] ;
 wire \myring.inv_in[106] ;
 wire \myring.inv_in[107] ;
 wire \myring.inv_in[108] ;
 wire \myring.inv_in[109] ;
 wire \myring.inv_in[10] ;
 wire \myring.inv_in[110] ;
 wire \myring.inv_in[111] ;
 wire \myring.inv_in[112] ;
 wire \myring.inv_in[113] ;
 wire \myring.inv_in[114] ;
 wire \myring.inv_in[115] ;
 wire \myring.inv_in[116] ;
 wire \myring.inv_in[117] ;
 wire \myring.inv_in[118] ;
 wire \myring.inv_in[119] ;
 wire \myring.inv_in[11] ;
 wire \myring.inv_in[120] ;
 wire \myring.inv_in[121] ;
 wire \myring.inv_in[122] ;
 wire \myring.inv_in[123] ;
 wire \myring.inv_in[124] ;
 wire \myring.inv_in[125] ;
 wire \myring.inv_in[126] ;
 wire \myring.inv_in[127] ;
 wire \myring.inv_in[128] ;
 wire \myring.inv_in[129] ;
 wire \myring.inv_in[12] ;
 wire \myring.inv_in[130] ;
 wire \myring.inv_in[131] ;
 wire \myring.inv_in[132] ;
 wire \myring.inv_in[133] ;
 wire \myring.inv_in[134] ;
 wire \myring.inv_in[135] ;
 wire \myring.inv_in[136] ;
 wire \myring.inv_in[137] ;
 wire \myring.inv_in[138] ;
 wire \myring.inv_in[139] ;
 wire \myring.inv_in[13] ;
 wire \myring.inv_in[140] ;
 wire \myring.inv_in[141] ;
 wire \myring.inv_in[142] ;
 wire \myring.inv_in[143] ;
 wire \myring.inv_in[144] ;
 wire \myring.inv_in[145] ;
 wire \myring.inv_in[146] ;
 wire \myring.inv_in[147] ;
 wire \myring.inv_in[148] ;
 wire \myring.inv_in[149] ;
 wire \myring.inv_in[14] ;
 wire \myring.inv_in[150] ;
 wire \myring.inv_in[151] ;
 wire \myring.inv_in[152] ;
 wire \myring.inv_in[153] ;
 wire \myring.inv_in[154] ;
 wire \myring.inv_in[155] ;
 wire \myring.inv_in[156] ;
 wire \myring.inv_in[157] ;
 wire \myring.inv_in[158] ;
 wire \myring.inv_in[159] ;
 wire \myring.inv_in[15] ;
 wire \myring.inv_in[160] ;
 wire \myring.inv_in[161] ;
 wire \myring.inv_in[162] ;
 wire \myring.inv_in[163] ;
 wire \myring.inv_in[164] ;
 wire \myring.inv_in[165] ;
 wire \myring.inv_in[166] ;
 wire \myring.inv_in[167] ;
 wire \myring.inv_in[168] ;
 wire \myring.inv_in[169] ;
 wire \myring.inv_in[16] ;
 wire \myring.inv_in[170] ;
 wire \myring.inv_in[171] ;
 wire \myring.inv_in[172] ;
 wire \myring.inv_in[173] ;
 wire \myring.inv_in[174] ;
 wire \myring.inv_in[175] ;
 wire \myring.inv_in[176] ;
 wire \myring.inv_in[177] ;
 wire \myring.inv_in[178] ;
 wire \myring.inv_in[179] ;
 wire \myring.inv_in[17] ;
 wire \myring.inv_in[180] ;
 wire \myring.inv_in[181] ;
 wire \myring.inv_in[182] ;
 wire \myring.inv_in[183] ;
 wire \myring.inv_in[184] ;
 wire \myring.inv_in[185] ;
 wire \myring.inv_in[186] ;
 wire \myring.inv_in[187] ;
 wire \myring.inv_in[188] ;
 wire \myring.inv_in[189] ;
 wire \myring.inv_in[18] ;
 wire \myring.inv_in[190] ;
 wire \myring.inv_in[191] ;
 wire \myring.inv_in[192] ;
 wire \myring.inv_in[193] ;
 wire \myring.inv_in[194] ;
 wire \myring.inv_in[195] ;
 wire \myring.inv_in[196] ;
 wire \myring.inv_in[197] ;
 wire \myring.inv_in[198] ;
 wire \myring.inv_in[199] ;
 wire \myring.inv_in[19] ;
 wire \myring.inv_in[1] ;
 wire \myring.inv_in[200] ;
 wire \myring.inv_in[201] ;
 wire \myring.inv_in[202] ;
 wire \myring.inv_in[203] ;
 wire \myring.inv_in[204] ;
 wire \myring.inv_in[205] ;
 wire \myring.inv_in[206] ;
 wire \myring.inv_in[207] ;
 wire \myring.inv_in[208] ;
 wire \myring.inv_in[209] ;
 wire \myring.inv_in[20] ;
 wire \myring.inv_in[210] ;
 wire \myring.inv_in[211] ;
 wire \myring.inv_in[212] ;
 wire \myring.inv_in[213] ;
 wire \myring.inv_in[214] ;
 wire \myring.inv_in[215] ;
 wire \myring.inv_in[216] ;
 wire \myring.inv_in[217] ;
 wire \myring.inv_in[218] ;
 wire \myring.inv_in[219] ;
 wire \myring.inv_in[21] ;
 wire \myring.inv_in[220] ;
 wire \myring.inv_in[221] ;
 wire \myring.inv_in[222] ;
 wire \myring.inv_in[223] ;
 wire \myring.inv_in[224] ;
 wire \myring.inv_in[225] ;
 wire \myring.inv_in[226] ;
 wire \myring.inv_in[227] ;
 wire \myring.inv_in[228] ;
 wire \myring.inv_in[229] ;
 wire \myring.inv_in[22] ;
 wire \myring.inv_in[230] ;
 wire \myring.inv_in[231] ;
 wire \myring.inv_in[232] ;
 wire \myring.inv_in[233] ;
 wire \myring.inv_in[234] ;
 wire \myring.inv_in[235] ;
 wire \myring.inv_in[236] ;
 wire \myring.inv_in[237] ;
 wire \myring.inv_in[238] ;
 wire \myring.inv_in[239] ;
 wire \myring.inv_in[23] ;
 wire \myring.inv_in[240] ;
 wire \myring.inv_in[241] ;
 wire \myring.inv_in[242] ;
 wire \myring.inv_in[243] ;
 wire \myring.inv_in[244] ;
 wire \myring.inv_in[245] ;
 wire \myring.inv_in[246] ;
 wire \myring.inv_in[247] ;
 wire \myring.inv_in[248] ;
 wire \myring.inv_in[249] ;
 wire \myring.inv_in[24] ;
 wire \myring.inv_in[250] ;
 wire \myring.inv_in[251] ;
 wire \myring.inv_in[252] ;
 wire \myring.inv_in[253] ;
 wire \myring.inv_in[254] ;
 wire \myring.inv_in[255] ;
 wire \myring.inv_in[256] ;
 wire \myring.inv_in[257] ;
 wire \myring.inv_in[258] ;
 wire \myring.inv_in[259] ;
 wire \myring.inv_in[25] ;
 wire \myring.inv_in[260] ;
 wire \myring.inv_in[261] ;
 wire \myring.inv_in[262] ;
 wire \myring.inv_in[263] ;
 wire \myring.inv_in[264] ;
 wire \myring.inv_in[265] ;
 wire \myring.inv_in[266] ;
 wire \myring.inv_in[267] ;
 wire \myring.inv_in[268] ;
 wire \myring.inv_in[269] ;
 wire \myring.inv_in[26] ;
 wire \myring.inv_in[270] ;
 wire \myring.inv_in[271] ;
 wire \myring.inv_in[272] ;
 wire \myring.inv_in[273] ;
 wire \myring.inv_in[274] ;
 wire \myring.inv_in[275] ;
 wire \myring.inv_in[276] ;
 wire \myring.inv_in[277] ;
 wire \myring.inv_in[278] ;
 wire \myring.inv_in[279] ;
 wire \myring.inv_in[27] ;
 wire \myring.inv_in[280] ;
 wire \myring.inv_in[281] ;
 wire \myring.inv_in[282] ;
 wire \myring.inv_in[283] ;
 wire \myring.inv_in[284] ;
 wire \myring.inv_in[285] ;
 wire \myring.inv_in[286] ;
 wire \myring.inv_in[287] ;
 wire \myring.inv_in[288] ;
 wire \myring.inv_in[289] ;
 wire \myring.inv_in[28] ;
 wire \myring.inv_in[290] ;
 wire \myring.inv_in[291] ;
 wire \myring.inv_in[292] ;
 wire \myring.inv_in[293] ;
 wire \myring.inv_in[294] ;
 wire \myring.inv_in[295] ;
 wire \myring.inv_in[296] ;
 wire \myring.inv_in[297] ;
 wire \myring.inv_in[298] ;
 wire \myring.inv_in[299] ;
 wire \myring.inv_in[29] ;
 wire \myring.inv_in[2] ;
 wire \myring.inv_in[300] ;
 wire \myring.inv_in[301] ;
 wire \myring.inv_in[302] ;
 wire \myring.inv_in[303] ;
 wire \myring.inv_in[304] ;
 wire \myring.inv_in[305] ;
 wire \myring.inv_in[306] ;
 wire \myring.inv_in[307] ;
 wire \myring.inv_in[308] ;
 wire \myring.inv_in[309] ;
 wire \myring.inv_in[30] ;
 wire \myring.inv_in[310] ;
 wire \myring.inv_in[311] ;
 wire \myring.inv_in[312] ;
 wire \myring.inv_in[313] ;
 wire \myring.inv_in[314] ;
 wire \myring.inv_in[315] ;
 wire \myring.inv_in[316] ;
 wire \myring.inv_in[317] ;
 wire \myring.inv_in[318] ;
 wire \myring.inv_in[319] ;
 wire \myring.inv_in[31] ;
 wire \myring.inv_in[320] ;
 wire \myring.inv_in[321] ;
 wire \myring.inv_in[322] ;
 wire \myring.inv_in[323] ;
 wire \myring.inv_in[324] ;
 wire \myring.inv_in[325] ;
 wire \myring.inv_in[326] ;
 wire \myring.inv_in[327] ;
 wire \myring.inv_in[328] ;
 wire \myring.inv_in[329] ;
 wire \myring.inv_in[32] ;
 wire \myring.inv_in[330] ;
 wire \myring.inv_in[331] ;
 wire \myring.inv_in[332] ;
 wire \myring.inv_in[333] ;
 wire \myring.inv_in[334] ;
 wire \myring.inv_in[335] ;
 wire \myring.inv_in[336] ;
 wire \myring.inv_in[337] ;
 wire \myring.inv_in[338] ;
 wire \myring.inv_in[339] ;
 wire \myring.inv_in[33] ;
 wire \myring.inv_in[340] ;
 wire \myring.inv_in[341] ;
 wire \myring.inv_in[342] ;
 wire \myring.inv_in[343] ;
 wire \myring.inv_in[344] ;
 wire \myring.inv_in[345] ;
 wire \myring.inv_in[346] ;
 wire \myring.inv_in[347] ;
 wire \myring.inv_in[348] ;
 wire \myring.inv_in[349] ;
 wire \myring.inv_in[34] ;
 wire \myring.inv_in[350] ;
 wire \myring.inv_in[351] ;
 wire \myring.inv_in[352] ;
 wire \myring.inv_in[353] ;
 wire \myring.inv_in[354] ;
 wire \myring.inv_in[355] ;
 wire \myring.inv_in[356] ;
 wire \myring.inv_in[357] ;
 wire \myring.inv_in[358] ;
 wire \myring.inv_in[359] ;
 wire \myring.inv_in[35] ;
 wire \myring.inv_in[360] ;
 wire \myring.inv_in[361] ;
 wire \myring.inv_in[362] ;
 wire \myring.inv_in[363] ;
 wire \myring.inv_in[364] ;
 wire \myring.inv_in[365] ;
 wire \myring.inv_in[366] ;
 wire \myring.inv_in[367] ;
 wire \myring.inv_in[368] ;
 wire \myring.inv_in[369] ;
 wire \myring.inv_in[36] ;
 wire \myring.inv_in[370] ;
 wire \myring.inv_in[371] ;
 wire \myring.inv_in[372] ;
 wire \myring.inv_in[373] ;
 wire \myring.inv_in[374] ;
 wire \myring.inv_in[375] ;
 wire \myring.inv_in[376] ;
 wire \myring.inv_in[377] ;
 wire \myring.inv_in[378] ;
 wire \myring.inv_in[379] ;
 wire \myring.inv_in[37] ;
 wire \myring.inv_in[380] ;
 wire \myring.inv_in[381] ;
 wire \myring.inv_in[382] ;
 wire \myring.inv_in[383] ;
 wire \myring.inv_in[384] ;
 wire \myring.inv_in[385] ;
 wire \myring.inv_in[386] ;
 wire \myring.inv_in[387] ;
 wire \myring.inv_in[388] ;
 wire \myring.inv_in[389] ;
 wire \myring.inv_in[38] ;
 wire \myring.inv_in[390] ;
 wire \myring.inv_in[391] ;
 wire \myring.inv_in[392] ;
 wire \myring.inv_in[393] ;
 wire \myring.inv_in[394] ;
 wire \myring.inv_in[395] ;
 wire \myring.inv_in[396] ;
 wire \myring.inv_in[397] ;
 wire \myring.inv_in[398] ;
 wire \myring.inv_in[399] ;
 wire \myring.inv_in[39] ;
 wire \myring.inv_in[3] ;
 wire \myring.inv_in[400] ;
 wire \myring.inv_in[401] ;
 wire \myring.inv_in[402] ;
 wire \myring.inv_in[403] ;
 wire \myring.inv_in[404] ;
 wire \myring.inv_in[405] ;
 wire \myring.inv_in[406] ;
 wire \myring.inv_in[407] ;
 wire \myring.inv_in[408] ;
 wire \myring.inv_in[409] ;
 wire \myring.inv_in[40] ;
 wire \myring.inv_in[410] ;
 wire \myring.inv_in[411] ;
 wire \myring.inv_in[412] ;
 wire \myring.inv_in[413] ;
 wire \myring.inv_in[414] ;
 wire \myring.inv_in[415] ;
 wire \myring.inv_in[416] ;
 wire \myring.inv_in[417] ;
 wire \myring.inv_in[418] ;
 wire \myring.inv_in[419] ;
 wire \myring.inv_in[41] ;
 wire \myring.inv_in[420] ;
 wire \myring.inv_in[421] ;
 wire \myring.inv_in[422] ;
 wire \myring.inv_in[423] ;
 wire \myring.inv_in[424] ;
 wire \myring.inv_in[425] ;
 wire \myring.inv_in[426] ;
 wire \myring.inv_in[427] ;
 wire \myring.inv_in[428] ;
 wire \myring.inv_in[429] ;
 wire \myring.inv_in[42] ;
 wire \myring.inv_in[430] ;
 wire \myring.inv_in[431] ;
 wire \myring.inv_in[432] ;
 wire \myring.inv_in[433] ;
 wire \myring.inv_in[434] ;
 wire \myring.inv_in[435] ;
 wire \myring.inv_in[436] ;
 wire \myring.inv_in[437] ;
 wire \myring.inv_in[438] ;
 wire \myring.inv_in[439] ;
 wire \myring.inv_in[43] ;
 wire \myring.inv_in[440] ;
 wire \myring.inv_in[441] ;
 wire \myring.inv_in[442] ;
 wire \myring.inv_in[443] ;
 wire \myring.inv_in[444] ;
 wire \myring.inv_in[445] ;
 wire \myring.inv_in[446] ;
 wire \myring.inv_in[447] ;
 wire \myring.inv_in[448] ;
 wire \myring.inv_in[449] ;
 wire \myring.inv_in[44] ;
 wire \myring.inv_in[450] ;
 wire \myring.inv_in[451] ;
 wire \myring.inv_in[452] ;
 wire \myring.inv_in[453] ;
 wire \myring.inv_in[454] ;
 wire \myring.inv_in[455] ;
 wire \myring.inv_in[456] ;
 wire \myring.inv_in[457] ;
 wire \myring.inv_in[458] ;
 wire \myring.inv_in[459] ;
 wire \myring.inv_in[45] ;
 wire \myring.inv_in[460] ;
 wire \myring.inv_in[461] ;
 wire \myring.inv_in[462] ;
 wire \myring.inv_in[463] ;
 wire \myring.inv_in[464] ;
 wire \myring.inv_in[465] ;
 wire \myring.inv_in[466] ;
 wire \myring.inv_in[467] ;
 wire \myring.inv_in[468] ;
 wire \myring.inv_in[469] ;
 wire \myring.inv_in[46] ;
 wire \myring.inv_in[470] ;
 wire \myring.inv_in[471] ;
 wire \myring.inv_in[472] ;
 wire \myring.inv_in[473] ;
 wire \myring.inv_in[474] ;
 wire \myring.inv_in[475] ;
 wire \myring.inv_in[476] ;
 wire \myring.inv_in[477] ;
 wire \myring.inv_in[478] ;
 wire \myring.inv_in[479] ;
 wire \myring.inv_in[47] ;
 wire \myring.inv_in[480] ;
 wire \myring.inv_in[481] ;
 wire \myring.inv_in[482] ;
 wire \myring.inv_in[483] ;
 wire \myring.inv_in[484] ;
 wire \myring.inv_in[485] ;
 wire \myring.inv_in[486] ;
 wire \myring.inv_in[487] ;
 wire \myring.inv_in[488] ;
 wire \myring.inv_in[489] ;
 wire \myring.inv_in[48] ;
 wire \myring.inv_in[490] ;
 wire \myring.inv_in[491] ;
 wire \myring.inv_in[492] ;
 wire \myring.inv_in[493] ;
 wire \myring.inv_in[494] ;
 wire \myring.inv_in[495] ;
 wire \myring.inv_in[496] ;
 wire \myring.inv_in[497] ;
 wire \myring.inv_in[498] ;
 wire \myring.inv_in[499] ;
 wire \myring.inv_in[49] ;
 wire \myring.inv_in[4] ;
 wire \myring.inv_in[500] ;
 wire \myring.inv_in[501] ;
 wire \myring.inv_in[502] ;
 wire \myring.inv_in[503] ;
 wire \myring.inv_in[504] ;
 wire \myring.inv_in[505] ;
 wire \myring.inv_in[506] ;
 wire \myring.inv_in[507] ;
 wire \myring.inv_in[508] ;
 wire \myring.inv_in[509] ;
 wire \myring.inv_in[50] ;
 wire \myring.inv_in[510] ;
 wire \myring.inv_in[511] ;
 wire \myring.inv_in[512] ;
 wire \myring.inv_in[513] ;
 wire \myring.inv_in[514] ;
 wire \myring.inv_in[515] ;
 wire \myring.inv_in[516] ;
 wire \myring.inv_in[517] ;
 wire \myring.inv_in[518] ;
 wire \myring.inv_in[519] ;
 wire \myring.inv_in[51] ;
 wire \myring.inv_in[520] ;
 wire \myring.inv_in[521] ;
 wire \myring.inv_in[522] ;
 wire \myring.inv_in[523] ;
 wire \myring.inv_in[524] ;
 wire \myring.inv_in[525] ;
 wire \myring.inv_in[526] ;
 wire \myring.inv_in[527] ;
 wire \myring.inv_in[528] ;
 wire \myring.inv_in[529] ;
 wire \myring.inv_in[52] ;
 wire \myring.inv_in[530] ;
 wire \myring.inv_in[531] ;
 wire \myring.inv_in[532] ;
 wire \myring.inv_in[533] ;
 wire \myring.inv_in[534] ;
 wire \myring.inv_in[535] ;
 wire \myring.inv_in[536] ;
 wire \myring.inv_in[537] ;
 wire \myring.inv_in[538] ;
 wire \myring.inv_in[539] ;
 wire \myring.inv_in[53] ;
 wire \myring.inv_in[540] ;
 wire \myring.inv_in[541] ;
 wire \myring.inv_in[542] ;
 wire \myring.inv_in[543] ;
 wire \myring.inv_in[544] ;
 wire \myring.inv_in[545] ;
 wire \myring.inv_in[546] ;
 wire \myring.inv_in[547] ;
 wire \myring.inv_in[548] ;
 wire \myring.inv_in[549] ;
 wire \myring.inv_in[54] ;
 wire \myring.inv_in[550] ;
 wire \myring.inv_in[551] ;
 wire \myring.inv_in[552] ;
 wire \myring.inv_in[553] ;
 wire \myring.inv_in[554] ;
 wire \myring.inv_in[555] ;
 wire \myring.inv_in[556] ;
 wire \myring.inv_in[557] ;
 wire \myring.inv_in[558] ;
 wire \myring.inv_in[559] ;
 wire \myring.inv_in[55] ;
 wire \myring.inv_in[560] ;
 wire \myring.inv_in[561] ;
 wire \myring.inv_in[562] ;
 wire \myring.inv_in[563] ;
 wire \myring.inv_in[564] ;
 wire \myring.inv_in[565] ;
 wire \myring.inv_in[566] ;
 wire \myring.inv_in[567] ;
 wire \myring.inv_in[568] ;
 wire \myring.inv_in[569] ;
 wire \myring.inv_in[56] ;
 wire \myring.inv_in[570] ;
 wire \myring.inv_in[571] ;
 wire \myring.inv_in[572] ;
 wire \myring.inv_in[573] ;
 wire \myring.inv_in[574] ;
 wire \myring.inv_in[575] ;
 wire \myring.inv_in[576] ;
 wire \myring.inv_in[577] ;
 wire \myring.inv_in[578] ;
 wire \myring.inv_in[579] ;
 wire \myring.inv_in[57] ;
 wire \myring.inv_in[580] ;
 wire \myring.inv_in[581] ;
 wire \myring.inv_in[582] ;
 wire \myring.inv_in[583] ;
 wire \myring.inv_in[584] ;
 wire \myring.inv_in[585] ;
 wire \myring.inv_in[586] ;
 wire \myring.inv_in[587] ;
 wire \myring.inv_in[588] ;
 wire \myring.inv_in[589] ;
 wire \myring.inv_in[58] ;
 wire \myring.inv_in[590] ;
 wire \myring.inv_in[591] ;
 wire \myring.inv_in[592] ;
 wire \myring.inv_in[593] ;
 wire \myring.inv_in[594] ;
 wire \myring.inv_in[595] ;
 wire \myring.inv_in[596] ;
 wire \myring.inv_in[597] ;
 wire \myring.inv_in[598] ;
 wire \myring.inv_in[599] ;
 wire \myring.inv_in[59] ;
 wire \myring.inv_in[5] ;
 wire \myring.inv_in[600] ;
 wire \myring.inv_in[601] ;
 wire \myring.inv_in[602] ;
 wire \myring.inv_in[603] ;
 wire \myring.inv_in[604] ;
 wire \myring.inv_in[605] ;
 wire \myring.inv_in[606] ;
 wire \myring.inv_in[607] ;
 wire \myring.inv_in[608] ;
 wire \myring.inv_in[609] ;
 wire \myring.inv_in[60] ;
 wire \myring.inv_in[610] ;
 wire \myring.inv_in[611] ;
 wire \myring.inv_in[612] ;
 wire \myring.inv_in[613] ;
 wire \myring.inv_in[614] ;
 wire \myring.inv_in[615] ;
 wire \myring.inv_in[616] ;
 wire \myring.inv_in[617] ;
 wire \myring.inv_in[618] ;
 wire \myring.inv_in[619] ;
 wire \myring.inv_in[61] ;
 wire \myring.inv_in[620] ;
 wire \myring.inv_in[621] ;
 wire \myring.inv_in[622] ;
 wire \myring.inv_in[623] ;
 wire \myring.inv_in[624] ;
 wire \myring.inv_in[625] ;
 wire \myring.inv_in[626] ;
 wire \myring.inv_in[627] ;
 wire \myring.inv_in[628] ;
 wire \myring.inv_in[629] ;
 wire \myring.inv_in[62] ;
 wire \myring.inv_in[630] ;
 wire \myring.inv_in[631] ;
 wire \myring.inv_in[632] ;
 wire \myring.inv_in[633] ;
 wire \myring.inv_in[634] ;
 wire \myring.inv_in[635] ;
 wire \myring.inv_in[636] ;
 wire \myring.inv_in[637] ;
 wire \myring.inv_in[638] ;
 wire \myring.inv_in[639] ;
 wire \myring.inv_in[63] ;
 wire \myring.inv_in[640] ;
 wire \myring.inv_in[641] ;
 wire \myring.inv_in[642] ;
 wire \myring.inv_in[643] ;
 wire \myring.inv_in[644] ;
 wire \myring.inv_in[645] ;
 wire \myring.inv_in[646] ;
 wire \myring.inv_in[647] ;
 wire \myring.inv_in[648] ;
 wire \myring.inv_in[649] ;
 wire \myring.inv_in[64] ;
 wire \myring.inv_in[650] ;
 wire \myring.inv_in[651] ;
 wire \myring.inv_in[652] ;
 wire \myring.inv_in[653] ;
 wire \myring.inv_in[654] ;
 wire \myring.inv_in[655] ;
 wire \myring.inv_in[656] ;
 wire \myring.inv_in[657] ;
 wire \myring.inv_in[658] ;
 wire \myring.inv_in[659] ;
 wire \myring.inv_in[65] ;
 wire \myring.inv_in[660] ;
 wire \myring.inv_in[661] ;
 wire \myring.inv_in[662] ;
 wire \myring.inv_in[663] ;
 wire \myring.inv_in[664] ;
 wire \myring.inv_in[665] ;
 wire \myring.inv_in[666] ;
 wire \myring.inv_in[667] ;
 wire \myring.inv_in[668] ;
 wire \myring.inv_in[669] ;
 wire \myring.inv_in[66] ;
 wire \myring.inv_in[670] ;
 wire \myring.inv_in[671] ;
 wire \myring.inv_in[672] ;
 wire \myring.inv_in[673] ;
 wire \myring.inv_in[674] ;
 wire \myring.inv_in[675] ;
 wire \myring.inv_in[676] ;
 wire \myring.inv_in[677] ;
 wire \myring.inv_in[678] ;
 wire \myring.inv_in[679] ;
 wire \myring.inv_in[67] ;
 wire \myring.inv_in[680] ;
 wire \myring.inv_in[681] ;
 wire \myring.inv_in[682] ;
 wire \myring.inv_in[683] ;
 wire \myring.inv_in[684] ;
 wire \myring.inv_in[685] ;
 wire \myring.inv_in[686] ;
 wire \myring.inv_in[687] ;
 wire \myring.inv_in[688] ;
 wire \myring.inv_in[689] ;
 wire \myring.inv_in[68] ;
 wire \myring.inv_in[690] ;
 wire \myring.inv_in[691] ;
 wire \myring.inv_in[692] ;
 wire \myring.inv_in[693] ;
 wire \myring.inv_in[694] ;
 wire \myring.inv_in[695] ;
 wire \myring.inv_in[696] ;
 wire \myring.inv_in[697] ;
 wire \myring.inv_in[698] ;
 wire \myring.inv_in[699] ;
 wire \myring.inv_in[69] ;
 wire \myring.inv_in[6] ;
 wire \myring.inv_in[700] ;
 wire \myring.inv_in[701] ;
 wire \myring.inv_in[702] ;
 wire \myring.inv_in[703] ;
 wire \myring.inv_in[704] ;
 wire \myring.inv_in[705] ;
 wire \myring.inv_in[706] ;
 wire \myring.inv_in[707] ;
 wire \myring.inv_in[708] ;
 wire \myring.inv_in[709] ;
 wire \myring.inv_in[70] ;
 wire \myring.inv_in[710] ;
 wire \myring.inv_in[711] ;
 wire \myring.inv_in[712] ;
 wire \myring.inv_in[713] ;
 wire \myring.inv_in[714] ;
 wire \myring.inv_in[715] ;
 wire \myring.inv_in[716] ;
 wire \myring.inv_in[717] ;
 wire \myring.inv_in[718] ;
 wire \myring.inv_in[719] ;
 wire \myring.inv_in[71] ;
 wire \myring.inv_in[720] ;
 wire \myring.inv_in[721] ;
 wire \myring.inv_in[722] ;
 wire \myring.inv_in[723] ;
 wire \myring.inv_in[724] ;
 wire \myring.inv_in[725] ;
 wire \myring.inv_in[726] ;
 wire \myring.inv_in[727] ;
 wire \myring.inv_in[728] ;
 wire \myring.inv_in[729] ;
 wire \myring.inv_in[72] ;
 wire \myring.inv_in[730] ;
 wire \myring.inv_in[731] ;
 wire \myring.inv_in[732] ;
 wire \myring.inv_in[733] ;
 wire \myring.inv_in[734] ;
 wire \myring.inv_in[735] ;
 wire \myring.inv_in[736] ;
 wire \myring.inv_in[737] ;
 wire \myring.inv_in[738] ;
 wire \myring.inv_in[739] ;
 wire \myring.inv_in[73] ;
 wire \myring.inv_in[740] ;
 wire \myring.inv_in[741] ;
 wire \myring.inv_in[742] ;
 wire \myring.inv_in[743] ;
 wire \myring.inv_in[744] ;
 wire \myring.inv_in[745] ;
 wire \myring.inv_in[746] ;
 wire \myring.inv_in[747] ;
 wire \myring.inv_in[748] ;
 wire \myring.inv_in[749] ;
 wire \myring.inv_in[74] ;
 wire \myring.inv_in[750] ;
 wire \myring.inv_in[751] ;
 wire \myring.inv_in[752] ;
 wire \myring.inv_in[753] ;
 wire \myring.inv_in[754] ;
 wire \myring.inv_in[755] ;
 wire \myring.inv_in[756] ;
 wire \myring.inv_in[757] ;
 wire \myring.inv_in[758] ;
 wire \myring.inv_in[759] ;
 wire \myring.inv_in[75] ;
 wire \myring.inv_in[760] ;
 wire \myring.inv_in[761] ;
 wire \myring.inv_in[762] ;
 wire \myring.inv_in[763] ;
 wire \myring.inv_in[764] ;
 wire \myring.inv_in[765] ;
 wire \myring.inv_in[766] ;
 wire \myring.inv_in[767] ;
 wire \myring.inv_in[768] ;
 wire \myring.inv_in[769] ;
 wire \myring.inv_in[76] ;
 wire \myring.inv_in[770] ;
 wire \myring.inv_in[771] ;
 wire \myring.inv_in[772] ;
 wire \myring.inv_in[773] ;
 wire \myring.inv_in[774] ;
 wire \myring.inv_in[775] ;
 wire \myring.inv_in[776] ;
 wire \myring.inv_in[777] ;
 wire \myring.inv_in[778] ;
 wire \myring.inv_in[779] ;
 wire \myring.inv_in[77] ;
 wire \myring.inv_in[780] ;
 wire \myring.inv_in[781] ;
 wire \myring.inv_in[782] ;
 wire \myring.inv_in[783] ;
 wire \myring.inv_in[784] ;
 wire \myring.inv_in[785] ;
 wire \myring.inv_in[786] ;
 wire \myring.inv_in[787] ;
 wire \myring.inv_in[788] ;
 wire \myring.inv_in[789] ;
 wire \myring.inv_in[78] ;
 wire \myring.inv_in[790] ;
 wire \myring.inv_in[791] ;
 wire \myring.inv_in[792] ;
 wire \myring.inv_in[793] ;
 wire \myring.inv_in[794] ;
 wire \myring.inv_in[795] ;
 wire \myring.inv_in[796] ;
 wire \myring.inv_in[797] ;
 wire \myring.inv_in[798] ;
 wire \myring.inv_in[799] ;
 wire \myring.inv_in[79] ;
 wire \myring.inv_in[7] ;
 wire \myring.inv_in[800] ;
 wire \myring.inv_in[801] ;
 wire \myring.inv_in[802] ;
 wire \myring.inv_in[803] ;
 wire \myring.inv_in[804] ;
 wire \myring.inv_in[805] ;
 wire \myring.inv_in[806] ;
 wire \myring.inv_in[807] ;
 wire \myring.inv_in[808] ;
 wire \myring.inv_in[809] ;
 wire \myring.inv_in[80] ;
 wire \myring.inv_in[810] ;
 wire \myring.inv_in[811] ;
 wire \myring.inv_in[812] ;
 wire \myring.inv_in[813] ;
 wire \myring.inv_in[814] ;
 wire \myring.inv_in[815] ;
 wire \myring.inv_in[816] ;
 wire \myring.inv_in[817] ;
 wire \myring.inv_in[818] ;
 wire \myring.inv_in[819] ;
 wire \myring.inv_in[81] ;
 wire \myring.inv_in[820] ;
 wire \myring.inv_in[821] ;
 wire \myring.inv_in[822] ;
 wire \myring.inv_in[823] ;
 wire \myring.inv_in[824] ;
 wire \myring.inv_in[825] ;
 wire \myring.inv_in[826] ;
 wire \myring.inv_in[827] ;
 wire \myring.inv_in[828] ;
 wire \myring.inv_in[829] ;
 wire \myring.inv_in[82] ;
 wire \myring.inv_in[830] ;
 wire \myring.inv_in[831] ;
 wire \myring.inv_in[832] ;
 wire \myring.inv_in[833] ;
 wire \myring.inv_in[834] ;
 wire \myring.inv_in[835] ;
 wire \myring.inv_in[836] ;
 wire \myring.inv_in[837] ;
 wire \myring.inv_in[838] ;
 wire \myring.inv_in[839] ;
 wire \myring.inv_in[83] ;
 wire \myring.inv_in[840] ;
 wire \myring.inv_in[841] ;
 wire \myring.inv_in[842] ;
 wire \myring.inv_in[843] ;
 wire \myring.inv_in[844] ;
 wire \myring.inv_in[845] ;
 wire \myring.inv_in[846] ;
 wire \myring.inv_in[847] ;
 wire \myring.inv_in[848] ;
 wire \myring.inv_in[849] ;
 wire \myring.inv_in[84] ;
 wire \myring.inv_in[850] ;
 wire \myring.inv_in[851] ;
 wire \myring.inv_in[852] ;
 wire \myring.inv_in[853] ;
 wire \myring.inv_in[854] ;
 wire \myring.inv_in[855] ;
 wire \myring.inv_in[856] ;
 wire \myring.inv_in[857] ;
 wire \myring.inv_in[858] ;
 wire \myring.inv_in[859] ;
 wire \myring.inv_in[85] ;
 wire \myring.inv_in[860] ;
 wire \myring.inv_in[861] ;
 wire \myring.inv_in[862] ;
 wire \myring.inv_in[863] ;
 wire \myring.inv_in[864] ;
 wire \myring.inv_in[865] ;
 wire \myring.inv_in[866] ;
 wire \myring.inv_in[867] ;
 wire \myring.inv_in[868] ;
 wire \myring.inv_in[869] ;
 wire \myring.inv_in[86] ;
 wire \myring.inv_in[870] ;
 wire \myring.inv_in[871] ;
 wire \myring.inv_in[872] ;
 wire \myring.inv_in[873] ;
 wire \myring.inv_in[874] ;
 wire \myring.inv_in[875] ;
 wire \myring.inv_in[876] ;
 wire \myring.inv_in[877] ;
 wire \myring.inv_in[878] ;
 wire \myring.inv_in[879] ;
 wire \myring.inv_in[87] ;
 wire \myring.inv_in[880] ;
 wire \myring.inv_in[881] ;
 wire \myring.inv_in[882] ;
 wire \myring.inv_in[883] ;
 wire \myring.inv_in[884] ;
 wire \myring.inv_in[885] ;
 wire \myring.inv_in[886] ;
 wire \myring.inv_in[887] ;
 wire \myring.inv_in[888] ;
 wire \myring.inv_in[889] ;
 wire \myring.inv_in[88] ;
 wire \myring.inv_in[890] ;
 wire \myring.inv_in[891] ;
 wire \myring.inv_in[892] ;
 wire \myring.inv_in[893] ;
 wire \myring.inv_in[894] ;
 wire \myring.inv_in[895] ;
 wire \myring.inv_in[896] ;
 wire \myring.inv_in[897] ;
 wire \myring.inv_in[898] ;
 wire \myring.inv_in[899] ;
 wire \myring.inv_in[89] ;
 wire \myring.inv_in[8] ;
 wire \myring.inv_in[900] ;
 wire \myring.inv_in[901] ;
 wire \myring.inv_in[902] ;
 wire \myring.inv_in[903] ;
 wire \myring.inv_in[904] ;
 wire \myring.inv_in[905] ;
 wire \myring.inv_in[906] ;
 wire \myring.inv_in[907] ;
 wire \myring.inv_in[908] ;
 wire \myring.inv_in[909] ;
 wire \myring.inv_in[90] ;
 wire \myring.inv_in[910] ;
 wire \myring.inv_in[911] ;
 wire \myring.inv_in[912] ;
 wire \myring.inv_in[913] ;
 wire \myring.inv_in[914] ;
 wire \myring.inv_in[915] ;
 wire \myring.inv_in[916] ;
 wire \myring.inv_in[917] ;
 wire \myring.inv_in[918] ;
 wire \myring.inv_in[919] ;
 wire \myring.inv_in[91] ;
 wire \myring.inv_in[920] ;
 wire \myring.inv_in[921] ;
 wire \myring.inv_in[922] ;
 wire \myring.inv_in[923] ;
 wire \myring.inv_in[924] ;
 wire \myring.inv_in[925] ;
 wire \myring.inv_in[926] ;
 wire \myring.inv_in[927] ;
 wire \myring.inv_in[928] ;
 wire \myring.inv_in[929] ;
 wire \myring.inv_in[92] ;
 wire \myring.inv_in[930] ;
 wire \myring.inv_in[931] ;
 wire \myring.inv_in[932] ;
 wire \myring.inv_in[933] ;
 wire \myring.inv_in[934] ;
 wire \myring.inv_in[935] ;
 wire \myring.inv_in[936] ;
 wire \myring.inv_in[937] ;
 wire \myring.inv_in[938] ;
 wire \myring.inv_in[939] ;
 wire \myring.inv_in[93] ;
 wire \myring.inv_in[940] ;
 wire \myring.inv_in[941] ;
 wire \myring.inv_in[942] ;
 wire \myring.inv_in[943] ;
 wire \myring.inv_in[944] ;
 wire \myring.inv_in[945] ;
 wire \myring.inv_in[946] ;
 wire \myring.inv_in[947] ;
 wire \myring.inv_in[948] ;
 wire \myring.inv_in[949] ;
 wire \myring.inv_in[94] ;
 wire \myring.inv_in[950] ;
 wire \myring.inv_in[951] ;
 wire \myring.inv_in[952] ;
 wire \myring.inv_in[953] ;
 wire \myring.inv_in[954] ;
 wire \myring.inv_in[955] ;
 wire \myring.inv_in[956] ;
 wire \myring.inv_in[957] ;
 wire \myring.inv_in[958] ;
 wire \myring.inv_in[959] ;
 wire \myring.inv_in[95] ;
 wire \myring.inv_in[960] ;
 wire \myring.inv_in[961] ;
 wire \myring.inv_in[962] ;
 wire \myring.inv_in[963] ;
 wire \myring.inv_in[964] ;
 wire \myring.inv_in[965] ;
 wire \myring.inv_in[966] ;
 wire \myring.inv_in[967] ;
 wire \myring.inv_in[968] ;
 wire \myring.inv_in[969] ;
 wire \myring.inv_in[96] ;
 wire \myring.inv_in[970] ;
 wire \myring.inv_in[971] ;
 wire \myring.inv_in[972] ;
 wire \myring.inv_in[973] ;
 wire \myring.inv_in[974] ;
 wire \myring.inv_in[975] ;
 wire \myring.inv_in[976] ;
 wire \myring.inv_in[977] ;
 wire \myring.inv_in[978] ;
 wire \myring.inv_in[979] ;
 wire \myring.inv_in[97] ;
 wire \myring.inv_in[980] ;
 wire \myring.inv_in[981] ;
 wire \myring.inv_in[982] ;
 wire \myring.inv_in[983] ;
 wire \myring.inv_in[984] ;
 wire \myring.inv_in[985] ;
 wire \myring.inv_in[986] ;
 wire \myring.inv_in[987] ;
 wire \myring.inv_in[988] ;
 wire \myring.inv_in[989] ;
 wire \myring.inv_in[98] ;
 wire \myring.inv_in[990] ;
 wire \myring.inv_in[991] ;
 wire \myring.inv_in[992] ;
 wire \myring.inv_in[993] ;
 wire \myring.inv_in[994] ;
 wire \myring.inv_in[995] ;
 wire \myring.inv_in[996] ;
 wire \myring.inv_in[997] ;
 wire \myring.inv_in[998] ;
 wire \myring.inv_in[999] ;
 wire \myring.inv_in[99] ;
 wire \myring.inv_in[9] ;
 wire \myring.inv_out[1000] ;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;

 sg13g2_and4_1 _05_ (.A(net6),
    .B(net5),
    .C(net8),
    .D(net7),
    .X(_00_));
 sg13g2_nand3_1 _06_ (.B(net3),
    .C(_00_),
    .A(net4),
    .Y(_01_));
 sg13g2_nand4_1 _07_ (.B(net17),
    .C(net2),
    .A(net18),
    .Y(_02_),
    .D(net1));
 sg13g2_nand4_1 _08_ (.B(net13),
    .C(net16),
    .A(net14),
    .Y(_03_),
    .D(net15));
 sg13g2_nand4_1 _09_ (.B(net9),
    .C(net12),
    .A(net10),
    .Y(_04_),
    .D(net11));
 sg13g2_nor4_1 _10_ (.A(_01_),
    .B(_02_),
    .C(_03_),
    .D(_04_),
    .Y(dummy));
 sg13g2_and2_1 _11_ (.A(net1),
    .B(\myring.inv_out[1000] ),
    .X(\myring.inv_in[0] ));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_20 (.L_LO(net20));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_21 (.L_LO(net21));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_22 (.L_LO(net22));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_23 (.L_LO(net23));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_24 (.L_LO(net24));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_25 (.L_LO(net25));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_26 (.L_LO(net26));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_27 (.L_LO(net27));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_28 (.L_LO(net28));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_29 (.L_LO(net29));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_30 (.L_LO(net30));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_31 (.L_LO(net31));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_32 (.L_LO(net32));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_33 (.L_LO(net33));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_34 (.L_LO(net34));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_35 (.L_LO(net35));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_36 (.L_LO(net36));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_37 (.L_LO(net37));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_38 (.L_LO(net38));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_39 (.L_LO(net39));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_40 (.L_LO(net40));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 _34_ (.A(\myring.inv_in[0] ),
    .X(uo_out[0]));
 sg13g2_buf_1 _35_ (.A(dummy),
    .X(uo_out[1]));
 sg13g2_inv_1 \myring.inv_array[0]/sky_inverter/_0_  (.Y(\myring.inv_in[1] ),
    .A(\myring.inv_in[0] ));
 sg13g2_inv_1 \myring.inv_array[1000]/sky_inverter/_0_  (.Y(\myring.inv_out[1000] ),
    .A(\myring.inv_in[1000] ));
 sg13g2_inv_1 \myring.inv_array[100]/sky_inverter/_0_  (.Y(\myring.inv_in[101] ),
    .A(\myring.inv_in[100] ));
 sg13g2_inv_1 \myring.inv_array[101]/sky_inverter/_0_  (.Y(\myring.inv_in[102] ),
    .A(\myring.inv_in[101] ));
 sg13g2_inv_1 \myring.inv_array[102]/sky_inverter/_0_  (.Y(\myring.inv_in[103] ),
    .A(\myring.inv_in[102] ));
 sg13g2_inv_1 \myring.inv_array[103]/sky_inverter/_0_  (.Y(\myring.inv_in[104] ),
    .A(\myring.inv_in[103] ));
 sg13g2_inv_1 \myring.inv_array[104]/sky_inverter/_0_  (.Y(\myring.inv_in[105] ),
    .A(\myring.inv_in[104] ));
 sg13g2_inv_1 \myring.inv_array[105]/sky_inverter/_0_  (.Y(\myring.inv_in[106] ),
    .A(\myring.inv_in[105] ));
 sg13g2_inv_1 \myring.inv_array[106]/sky_inverter/_0_  (.Y(\myring.inv_in[107] ),
    .A(\myring.inv_in[106] ));
 sg13g2_inv_1 \myring.inv_array[107]/sky_inverter/_0_  (.Y(\myring.inv_in[108] ),
    .A(\myring.inv_in[107] ));
 sg13g2_inv_1 \myring.inv_array[108]/sky_inverter/_0_  (.Y(\myring.inv_in[109] ),
    .A(\myring.inv_in[108] ));
 sg13g2_inv_1 \myring.inv_array[109]/sky_inverter/_0_  (.Y(\myring.inv_in[110] ),
    .A(\myring.inv_in[109] ));
 sg13g2_inv_1 \myring.inv_array[10]/sky_inverter/_0_  (.Y(\myring.inv_in[11] ),
    .A(\myring.inv_in[10] ));
 sg13g2_inv_1 \myring.inv_array[110]/sky_inverter/_0_  (.Y(\myring.inv_in[111] ),
    .A(\myring.inv_in[110] ));
 sg13g2_inv_1 \myring.inv_array[111]/sky_inverter/_0_  (.Y(\myring.inv_in[112] ),
    .A(\myring.inv_in[111] ));
 sg13g2_inv_1 \myring.inv_array[112]/sky_inverter/_0_  (.Y(\myring.inv_in[113] ),
    .A(\myring.inv_in[112] ));
 sg13g2_inv_1 \myring.inv_array[113]/sky_inverter/_0_  (.Y(\myring.inv_in[114] ),
    .A(\myring.inv_in[113] ));
 sg13g2_inv_1 \myring.inv_array[114]/sky_inverter/_0_  (.Y(\myring.inv_in[115] ),
    .A(\myring.inv_in[114] ));
 sg13g2_inv_1 \myring.inv_array[115]/sky_inverter/_0_  (.Y(\myring.inv_in[116] ),
    .A(\myring.inv_in[115] ));
 sg13g2_inv_1 \myring.inv_array[116]/sky_inverter/_0_  (.Y(\myring.inv_in[117] ),
    .A(\myring.inv_in[116] ));
 sg13g2_inv_1 \myring.inv_array[117]/sky_inverter/_0_  (.Y(\myring.inv_in[118] ),
    .A(\myring.inv_in[117] ));
 sg13g2_inv_1 \myring.inv_array[118]/sky_inverter/_0_  (.Y(\myring.inv_in[119] ),
    .A(\myring.inv_in[118] ));
 sg13g2_inv_1 \myring.inv_array[119]/sky_inverter/_0_  (.Y(\myring.inv_in[120] ),
    .A(\myring.inv_in[119] ));
 sg13g2_inv_1 \myring.inv_array[11]/sky_inverter/_0_  (.Y(\myring.inv_in[12] ),
    .A(\myring.inv_in[11] ));
 sg13g2_inv_1 \myring.inv_array[120]/sky_inverter/_0_  (.Y(\myring.inv_in[121] ),
    .A(\myring.inv_in[120] ));
 sg13g2_inv_1 \myring.inv_array[121]/sky_inverter/_0_  (.Y(\myring.inv_in[122] ),
    .A(\myring.inv_in[121] ));
 sg13g2_inv_1 \myring.inv_array[122]/sky_inverter/_0_  (.Y(\myring.inv_in[123] ),
    .A(\myring.inv_in[122] ));
 sg13g2_inv_1 \myring.inv_array[123]/sky_inverter/_0_  (.Y(\myring.inv_in[124] ),
    .A(\myring.inv_in[123] ));
 sg13g2_inv_1 \myring.inv_array[124]/sky_inverter/_0_  (.Y(\myring.inv_in[125] ),
    .A(\myring.inv_in[124] ));
 sg13g2_inv_1 \myring.inv_array[125]/sky_inverter/_0_  (.Y(\myring.inv_in[126] ),
    .A(\myring.inv_in[125] ));
 sg13g2_inv_1 \myring.inv_array[126]/sky_inverter/_0_  (.Y(\myring.inv_in[127] ),
    .A(\myring.inv_in[126] ));
 sg13g2_inv_1 \myring.inv_array[127]/sky_inverter/_0_  (.Y(\myring.inv_in[128] ),
    .A(\myring.inv_in[127] ));
 sg13g2_inv_1 \myring.inv_array[128]/sky_inverter/_0_  (.Y(\myring.inv_in[129] ),
    .A(\myring.inv_in[128] ));
 sg13g2_inv_1 \myring.inv_array[129]/sky_inverter/_0_  (.Y(\myring.inv_in[130] ),
    .A(\myring.inv_in[129] ));
 sg13g2_inv_1 \myring.inv_array[12]/sky_inverter/_0_  (.Y(\myring.inv_in[13] ),
    .A(\myring.inv_in[12] ));
 sg13g2_inv_1 \myring.inv_array[130]/sky_inverter/_0_  (.Y(\myring.inv_in[131] ),
    .A(\myring.inv_in[130] ));
 sg13g2_inv_1 \myring.inv_array[131]/sky_inverter/_0_  (.Y(\myring.inv_in[132] ),
    .A(\myring.inv_in[131] ));
 sg13g2_inv_1 \myring.inv_array[132]/sky_inverter/_0_  (.Y(\myring.inv_in[133] ),
    .A(\myring.inv_in[132] ));
 sg13g2_inv_1 \myring.inv_array[133]/sky_inverter/_0_  (.Y(\myring.inv_in[134] ),
    .A(\myring.inv_in[133] ));
 sg13g2_inv_1 \myring.inv_array[134]/sky_inverter/_0_  (.Y(\myring.inv_in[135] ),
    .A(\myring.inv_in[134] ));
 sg13g2_inv_1 \myring.inv_array[135]/sky_inverter/_0_  (.Y(\myring.inv_in[136] ),
    .A(\myring.inv_in[135] ));
 sg13g2_inv_1 \myring.inv_array[136]/sky_inverter/_0_  (.Y(\myring.inv_in[137] ),
    .A(\myring.inv_in[136] ));
 sg13g2_inv_1 \myring.inv_array[137]/sky_inverter/_0_  (.Y(\myring.inv_in[138] ),
    .A(\myring.inv_in[137] ));
 sg13g2_inv_1 \myring.inv_array[138]/sky_inverter/_0_  (.Y(\myring.inv_in[139] ),
    .A(\myring.inv_in[138] ));
 sg13g2_inv_1 \myring.inv_array[139]/sky_inverter/_0_  (.Y(\myring.inv_in[140] ),
    .A(\myring.inv_in[139] ));
 sg13g2_inv_1 \myring.inv_array[13]/sky_inverter/_0_  (.Y(\myring.inv_in[14] ),
    .A(\myring.inv_in[13] ));
 sg13g2_inv_1 \myring.inv_array[140]/sky_inverter/_0_  (.Y(\myring.inv_in[141] ),
    .A(\myring.inv_in[140] ));
 sg13g2_inv_1 \myring.inv_array[141]/sky_inverter/_0_  (.Y(\myring.inv_in[142] ),
    .A(\myring.inv_in[141] ));
 sg13g2_inv_1 \myring.inv_array[142]/sky_inverter/_0_  (.Y(\myring.inv_in[143] ),
    .A(\myring.inv_in[142] ));
 sg13g2_inv_1 \myring.inv_array[143]/sky_inverter/_0_  (.Y(\myring.inv_in[144] ),
    .A(\myring.inv_in[143] ));
 sg13g2_inv_1 \myring.inv_array[144]/sky_inverter/_0_  (.Y(\myring.inv_in[145] ),
    .A(\myring.inv_in[144] ));
 sg13g2_inv_1 \myring.inv_array[145]/sky_inverter/_0_  (.Y(\myring.inv_in[146] ),
    .A(\myring.inv_in[145] ));
 sg13g2_inv_1 \myring.inv_array[146]/sky_inverter/_0_  (.Y(\myring.inv_in[147] ),
    .A(\myring.inv_in[146] ));
 sg13g2_inv_1 \myring.inv_array[147]/sky_inverter/_0_  (.Y(\myring.inv_in[148] ),
    .A(\myring.inv_in[147] ));
 sg13g2_inv_1 \myring.inv_array[148]/sky_inverter/_0_  (.Y(\myring.inv_in[149] ),
    .A(\myring.inv_in[148] ));
 sg13g2_inv_1 \myring.inv_array[149]/sky_inverter/_0_  (.Y(\myring.inv_in[150] ),
    .A(\myring.inv_in[149] ));
 sg13g2_inv_1 \myring.inv_array[14]/sky_inverter/_0_  (.Y(\myring.inv_in[15] ),
    .A(\myring.inv_in[14] ));
 sg13g2_inv_1 \myring.inv_array[150]/sky_inverter/_0_  (.Y(\myring.inv_in[151] ),
    .A(\myring.inv_in[150] ));
 sg13g2_inv_1 \myring.inv_array[151]/sky_inverter/_0_  (.Y(\myring.inv_in[152] ),
    .A(\myring.inv_in[151] ));
 sg13g2_inv_1 \myring.inv_array[152]/sky_inverter/_0_  (.Y(\myring.inv_in[153] ),
    .A(\myring.inv_in[152] ));
 sg13g2_inv_1 \myring.inv_array[153]/sky_inverter/_0_  (.Y(\myring.inv_in[154] ),
    .A(\myring.inv_in[153] ));
 sg13g2_inv_1 \myring.inv_array[154]/sky_inverter/_0_  (.Y(\myring.inv_in[155] ),
    .A(\myring.inv_in[154] ));
 sg13g2_inv_1 \myring.inv_array[155]/sky_inverter/_0_  (.Y(\myring.inv_in[156] ),
    .A(\myring.inv_in[155] ));
 sg13g2_inv_1 \myring.inv_array[156]/sky_inverter/_0_  (.Y(\myring.inv_in[157] ),
    .A(\myring.inv_in[156] ));
 sg13g2_inv_1 \myring.inv_array[157]/sky_inverter/_0_  (.Y(\myring.inv_in[158] ),
    .A(\myring.inv_in[157] ));
 sg13g2_inv_1 \myring.inv_array[158]/sky_inverter/_0_  (.Y(\myring.inv_in[159] ),
    .A(\myring.inv_in[158] ));
 sg13g2_inv_1 \myring.inv_array[159]/sky_inverter/_0_  (.Y(\myring.inv_in[160] ),
    .A(\myring.inv_in[159] ));
 sg13g2_inv_1 \myring.inv_array[15]/sky_inverter/_0_  (.Y(\myring.inv_in[16] ),
    .A(\myring.inv_in[15] ));
 sg13g2_inv_1 \myring.inv_array[160]/sky_inverter/_0_  (.Y(\myring.inv_in[161] ),
    .A(\myring.inv_in[160] ));
 sg13g2_inv_1 \myring.inv_array[161]/sky_inverter/_0_  (.Y(\myring.inv_in[162] ),
    .A(\myring.inv_in[161] ));
 sg13g2_inv_1 \myring.inv_array[162]/sky_inverter/_0_  (.Y(\myring.inv_in[163] ),
    .A(\myring.inv_in[162] ));
 sg13g2_inv_1 \myring.inv_array[163]/sky_inverter/_0_  (.Y(\myring.inv_in[164] ),
    .A(\myring.inv_in[163] ));
 sg13g2_inv_1 \myring.inv_array[164]/sky_inverter/_0_  (.Y(\myring.inv_in[165] ),
    .A(\myring.inv_in[164] ));
 sg13g2_inv_1 \myring.inv_array[165]/sky_inverter/_0_  (.Y(\myring.inv_in[166] ),
    .A(\myring.inv_in[165] ));
 sg13g2_inv_1 \myring.inv_array[166]/sky_inverter/_0_  (.Y(\myring.inv_in[167] ),
    .A(\myring.inv_in[166] ));
 sg13g2_inv_1 \myring.inv_array[167]/sky_inverter/_0_  (.Y(\myring.inv_in[168] ),
    .A(\myring.inv_in[167] ));
 sg13g2_inv_1 \myring.inv_array[168]/sky_inverter/_0_  (.Y(\myring.inv_in[169] ),
    .A(\myring.inv_in[168] ));
 sg13g2_inv_1 \myring.inv_array[169]/sky_inverter/_0_  (.Y(\myring.inv_in[170] ),
    .A(\myring.inv_in[169] ));
 sg13g2_inv_1 \myring.inv_array[16]/sky_inverter/_0_  (.Y(\myring.inv_in[17] ),
    .A(\myring.inv_in[16] ));
 sg13g2_inv_1 \myring.inv_array[170]/sky_inverter/_0_  (.Y(\myring.inv_in[171] ),
    .A(\myring.inv_in[170] ));
 sg13g2_inv_1 \myring.inv_array[171]/sky_inverter/_0_  (.Y(\myring.inv_in[172] ),
    .A(\myring.inv_in[171] ));
 sg13g2_inv_1 \myring.inv_array[172]/sky_inverter/_0_  (.Y(\myring.inv_in[173] ),
    .A(\myring.inv_in[172] ));
 sg13g2_inv_1 \myring.inv_array[173]/sky_inverter/_0_  (.Y(\myring.inv_in[174] ),
    .A(\myring.inv_in[173] ));
 sg13g2_inv_1 \myring.inv_array[174]/sky_inverter/_0_  (.Y(\myring.inv_in[175] ),
    .A(\myring.inv_in[174] ));
 sg13g2_inv_1 \myring.inv_array[175]/sky_inverter/_0_  (.Y(\myring.inv_in[176] ),
    .A(\myring.inv_in[175] ));
 sg13g2_inv_1 \myring.inv_array[176]/sky_inverter/_0_  (.Y(\myring.inv_in[177] ),
    .A(\myring.inv_in[176] ));
 sg13g2_inv_1 \myring.inv_array[177]/sky_inverter/_0_  (.Y(\myring.inv_in[178] ),
    .A(\myring.inv_in[177] ));
 sg13g2_inv_1 \myring.inv_array[178]/sky_inverter/_0_  (.Y(\myring.inv_in[179] ),
    .A(\myring.inv_in[178] ));
 sg13g2_inv_1 \myring.inv_array[179]/sky_inverter/_0_  (.Y(\myring.inv_in[180] ),
    .A(\myring.inv_in[179] ));
 sg13g2_inv_1 \myring.inv_array[17]/sky_inverter/_0_  (.Y(\myring.inv_in[18] ),
    .A(\myring.inv_in[17] ));
 sg13g2_inv_1 \myring.inv_array[180]/sky_inverter/_0_  (.Y(\myring.inv_in[181] ),
    .A(\myring.inv_in[180] ));
 sg13g2_inv_1 \myring.inv_array[181]/sky_inverter/_0_  (.Y(\myring.inv_in[182] ),
    .A(\myring.inv_in[181] ));
 sg13g2_inv_1 \myring.inv_array[182]/sky_inverter/_0_  (.Y(\myring.inv_in[183] ),
    .A(\myring.inv_in[182] ));
 sg13g2_inv_1 \myring.inv_array[183]/sky_inverter/_0_  (.Y(\myring.inv_in[184] ),
    .A(\myring.inv_in[183] ));
 sg13g2_inv_1 \myring.inv_array[184]/sky_inverter/_0_  (.Y(\myring.inv_in[185] ),
    .A(\myring.inv_in[184] ));
 sg13g2_inv_1 \myring.inv_array[185]/sky_inverter/_0_  (.Y(\myring.inv_in[186] ),
    .A(\myring.inv_in[185] ));
 sg13g2_inv_1 \myring.inv_array[186]/sky_inverter/_0_  (.Y(\myring.inv_in[187] ),
    .A(\myring.inv_in[186] ));
 sg13g2_inv_1 \myring.inv_array[187]/sky_inverter/_0_  (.Y(\myring.inv_in[188] ),
    .A(\myring.inv_in[187] ));
 sg13g2_inv_1 \myring.inv_array[188]/sky_inverter/_0_  (.Y(\myring.inv_in[189] ),
    .A(\myring.inv_in[188] ));
 sg13g2_inv_1 \myring.inv_array[189]/sky_inverter/_0_  (.Y(\myring.inv_in[190] ),
    .A(\myring.inv_in[189] ));
 sg13g2_inv_1 \myring.inv_array[18]/sky_inverter/_0_  (.Y(\myring.inv_in[19] ),
    .A(\myring.inv_in[18] ));
 sg13g2_inv_1 \myring.inv_array[190]/sky_inverter/_0_  (.Y(\myring.inv_in[191] ),
    .A(\myring.inv_in[190] ));
 sg13g2_inv_1 \myring.inv_array[191]/sky_inverter/_0_  (.Y(\myring.inv_in[192] ),
    .A(\myring.inv_in[191] ));
 sg13g2_inv_1 \myring.inv_array[192]/sky_inverter/_0_  (.Y(\myring.inv_in[193] ),
    .A(\myring.inv_in[192] ));
 sg13g2_inv_1 \myring.inv_array[193]/sky_inverter/_0_  (.Y(\myring.inv_in[194] ),
    .A(\myring.inv_in[193] ));
 sg13g2_inv_1 \myring.inv_array[194]/sky_inverter/_0_  (.Y(\myring.inv_in[195] ),
    .A(\myring.inv_in[194] ));
 sg13g2_inv_1 \myring.inv_array[195]/sky_inverter/_0_  (.Y(\myring.inv_in[196] ),
    .A(\myring.inv_in[195] ));
 sg13g2_inv_1 \myring.inv_array[196]/sky_inverter/_0_  (.Y(\myring.inv_in[197] ),
    .A(\myring.inv_in[196] ));
 sg13g2_inv_1 \myring.inv_array[197]/sky_inverter/_0_  (.Y(\myring.inv_in[198] ),
    .A(\myring.inv_in[197] ));
 sg13g2_inv_1 \myring.inv_array[198]/sky_inverter/_0_  (.Y(\myring.inv_in[199] ),
    .A(\myring.inv_in[198] ));
 sg13g2_inv_1 \myring.inv_array[199]/sky_inverter/_0_  (.Y(\myring.inv_in[200] ),
    .A(\myring.inv_in[199] ));
 sg13g2_inv_1 \myring.inv_array[19]/sky_inverter/_0_  (.Y(\myring.inv_in[20] ),
    .A(\myring.inv_in[19] ));
 sg13g2_inv_1 \myring.inv_array[1]/sky_inverter/_0_  (.Y(\myring.inv_in[2] ),
    .A(\myring.inv_in[1] ));
 sg13g2_inv_1 \myring.inv_array[200]/sky_inverter/_0_  (.Y(\myring.inv_in[201] ),
    .A(\myring.inv_in[200] ));
 sg13g2_inv_1 \myring.inv_array[201]/sky_inverter/_0_  (.Y(\myring.inv_in[202] ),
    .A(\myring.inv_in[201] ));
 sg13g2_inv_1 \myring.inv_array[202]/sky_inverter/_0_  (.Y(\myring.inv_in[203] ),
    .A(\myring.inv_in[202] ));
 sg13g2_inv_1 \myring.inv_array[203]/sky_inverter/_0_  (.Y(\myring.inv_in[204] ),
    .A(\myring.inv_in[203] ));
 sg13g2_inv_1 \myring.inv_array[204]/sky_inverter/_0_  (.Y(\myring.inv_in[205] ),
    .A(\myring.inv_in[204] ));
 sg13g2_inv_1 \myring.inv_array[205]/sky_inverter/_0_  (.Y(\myring.inv_in[206] ),
    .A(\myring.inv_in[205] ));
 sg13g2_inv_1 \myring.inv_array[206]/sky_inverter/_0_  (.Y(\myring.inv_in[207] ),
    .A(\myring.inv_in[206] ));
 sg13g2_inv_1 \myring.inv_array[207]/sky_inverter/_0_  (.Y(\myring.inv_in[208] ),
    .A(\myring.inv_in[207] ));
 sg13g2_inv_1 \myring.inv_array[208]/sky_inverter/_0_  (.Y(\myring.inv_in[209] ),
    .A(\myring.inv_in[208] ));
 sg13g2_inv_1 \myring.inv_array[209]/sky_inverter/_0_  (.Y(\myring.inv_in[210] ),
    .A(\myring.inv_in[209] ));
 sg13g2_inv_1 \myring.inv_array[20]/sky_inverter/_0_  (.Y(\myring.inv_in[21] ),
    .A(\myring.inv_in[20] ));
 sg13g2_inv_1 \myring.inv_array[210]/sky_inverter/_0_  (.Y(\myring.inv_in[211] ),
    .A(\myring.inv_in[210] ));
 sg13g2_inv_1 \myring.inv_array[211]/sky_inverter/_0_  (.Y(\myring.inv_in[212] ),
    .A(\myring.inv_in[211] ));
 sg13g2_inv_1 \myring.inv_array[212]/sky_inverter/_0_  (.Y(\myring.inv_in[213] ),
    .A(\myring.inv_in[212] ));
 sg13g2_inv_1 \myring.inv_array[213]/sky_inverter/_0_  (.Y(\myring.inv_in[214] ),
    .A(\myring.inv_in[213] ));
 sg13g2_inv_1 \myring.inv_array[214]/sky_inverter/_0_  (.Y(\myring.inv_in[215] ),
    .A(\myring.inv_in[214] ));
 sg13g2_inv_1 \myring.inv_array[215]/sky_inverter/_0_  (.Y(\myring.inv_in[216] ),
    .A(\myring.inv_in[215] ));
 sg13g2_inv_1 \myring.inv_array[216]/sky_inverter/_0_  (.Y(\myring.inv_in[217] ),
    .A(\myring.inv_in[216] ));
 sg13g2_inv_1 \myring.inv_array[217]/sky_inverter/_0_  (.Y(\myring.inv_in[218] ),
    .A(\myring.inv_in[217] ));
 sg13g2_inv_1 \myring.inv_array[218]/sky_inverter/_0_  (.Y(\myring.inv_in[219] ),
    .A(\myring.inv_in[218] ));
 sg13g2_inv_1 \myring.inv_array[219]/sky_inverter/_0_  (.Y(\myring.inv_in[220] ),
    .A(\myring.inv_in[219] ));
 sg13g2_inv_1 \myring.inv_array[21]/sky_inverter/_0_  (.Y(\myring.inv_in[22] ),
    .A(\myring.inv_in[21] ));
 sg13g2_inv_1 \myring.inv_array[220]/sky_inverter/_0_  (.Y(\myring.inv_in[221] ),
    .A(\myring.inv_in[220] ));
 sg13g2_inv_1 \myring.inv_array[221]/sky_inverter/_0_  (.Y(\myring.inv_in[222] ),
    .A(\myring.inv_in[221] ));
 sg13g2_inv_1 \myring.inv_array[222]/sky_inverter/_0_  (.Y(\myring.inv_in[223] ),
    .A(\myring.inv_in[222] ));
 sg13g2_inv_1 \myring.inv_array[223]/sky_inverter/_0_  (.Y(\myring.inv_in[224] ),
    .A(\myring.inv_in[223] ));
 sg13g2_inv_1 \myring.inv_array[224]/sky_inverter/_0_  (.Y(\myring.inv_in[225] ),
    .A(\myring.inv_in[224] ));
 sg13g2_inv_1 \myring.inv_array[225]/sky_inverter/_0_  (.Y(\myring.inv_in[226] ),
    .A(\myring.inv_in[225] ));
 sg13g2_inv_1 \myring.inv_array[226]/sky_inverter/_0_  (.Y(\myring.inv_in[227] ),
    .A(\myring.inv_in[226] ));
 sg13g2_inv_1 \myring.inv_array[227]/sky_inverter/_0_  (.Y(\myring.inv_in[228] ),
    .A(\myring.inv_in[227] ));
 sg13g2_inv_1 \myring.inv_array[228]/sky_inverter/_0_  (.Y(\myring.inv_in[229] ),
    .A(\myring.inv_in[228] ));
 sg13g2_inv_1 \myring.inv_array[229]/sky_inverter/_0_  (.Y(\myring.inv_in[230] ),
    .A(\myring.inv_in[229] ));
 sg13g2_inv_1 \myring.inv_array[22]/sky_inverter/_0_  (.Y(\myring.inv_in[23] ),
    .A(\myring.inv_in[22] ));
 sg13g2_inv_1 \myring.inv_array[230]/sky_inverter/_0_  (.Y(\myring.inv_in[231] ),
    .A(\myring.inv_in[230] ));
 sg13g2_inv_1 \myring.inv_array[231]/sky_inverter/_0_  (.Y(\myring.inv_in[232] ),
    .A(\myring.inv_in[231] ));
 sg13g2_inv_1 \myring.inv_array[232]/sky_inverter/_0_  (.Y(\myring.inv_in[233] ),
    .A(\myring.inv_in[232] ));
 sg13g2_inv_1 \myring.inv_array[233]/sky_inverter/_0_  (.Y(\myring.inv_in[234] ),
    .A(\myring.inv_in[233] ));
 sg13g2_inv_1 \myring.inv_array[234]/sky_inverter/_0_  (.Y(\myring.inv_in[235] ),
    .A(\myring.inv_in[234] ));
 sg13g2_inv_1 \myring.inv_array[235]/sky_inverter/_0_  (.Y(\myring.inv_in[236] ),
    .A(\myring.inv_in[235] ));
 sg13g2_inv_1 \myring.inv_array[236]/sky_inverter/_0_  (.Y(\myring.inv_in[237] ),
    .A(\myring.inv_in[236] ));
 sg13g2_inv_1 \myring.inv_array[237]/sky_inverter/_0_  (.Y(\myring.inv_in[238] ),
    .A(\myring.inv_in[237] ));
 sg13g2_inv_1 \myring.inv_array[238]/sky_inverter/_0_  (.Y(\myring.inv_in[239] ),
    .A(\myring.inv_in[238] ));
 sg13g2_inv_1 \myring.inv_array[239]/sky_inverter/_0_  (.Y(\myring.inv_in[240] ),
    .A(\myring.inv_in[239] ));
 sg13g2_inv_1 \myring.inv_array[23]/sky_inverter/_0_  (.Y(\myring.inv_in[24] ),
    .A(\myring.inv_in[23] ));
 sg13g2_inv_1 \myring.inv_array[240]/sky_inverter/_0_  (.Y(\myring.inv_in[241] ),
    .A(\myring.inv_in[240] ));
 sg13g2_inv_1 \myring.inv_array[241]/sky_inverter/_0_  (.Y(\myring.inv_in[242] ),
    .A(\myring.inv_in[241] ));
 sg13g2_inv_1 \myring.inv_array[242]/sky_inverter/_0_  (.Y(\myring.inv_in[243] ),
    .A(\myring.inv_in[242] ));
 sg13g2_inv_1 \myring.inv_array[243]/sky_inverter/_0_  (.Y(\myring.inv_in[244] ),
    .A(\myring.inv_in[243] ));
 sg13g2_inv_1 \myring.inv_array[244]/sky_inverter/_0_  (.Y(\myring.inv_in[245] ),
    .A(\myring.inv_in[244] ));
 sg13g2_inv_1 \myring.inv_array[245]/sky_inverter/_0_  (.Y(\myring.inv_in[246] ),
    .A(\myring.inv_in[245] ));
 sg13g2_inv_1 \myring.inv_array[246]/sky_inverter/_0_  (.Y(\myring.inv_in[247] ),
    .A(\myring.inv_in[246] ));
 sg13g2_inv_1 \myring.inv_array[247]/sky_inverter/_0_  (.Y(\myring.inv_in[248] ),
    .A(\myring.inv_in[247] ));
 sg13g2_inv_1 \myring.inv_array[248]/sky_inverter/_0_  (.Y(\myring.inv_in[249] ),
    .A(\myring.inv_in[248] ));
 sg13g2_inv_1 \myring.inv_array[249]/sky_inverter/_0_  (.Y(\myring.inv_in[250] ),
    .A(\myring.inv_in[249] ));
 sg13g2_inv_1 \myring.inv_array[24]/sky_inverter/_0_  (.Y(\myring.inv_in[25] ),
    .A(\myring.inv_in[24] ));
 sg13g2_inv_1 \myring.inv_array[250]/sky_inverter/_0_  (.Y(\myring.inv_in[251] ),
    .A(\myring.inv_in[250] ));
 sg13g2_inv_1 \myring.inv_array[251]/sky_inverter/_0_  (.Y(\myring.inv_in[252] ),
    .A(\myring.inv_in[251] ));
 sg13g2_inv_1 \myring.inv_array[252]/sky_inverter/_0_  (.Y(\myring.inv_in[253] ),
    .A(\myring.inv_in[252] ));
 sg13g2_inv_1 \myring.inv_array[253]/sky_inverter/_0_  (.Y(\myring.inv_in[254] ),
    .A(\myring.inv_in[253] ));
 sg13g2_inv_1 \myring.inv_array[254]/sky_inverter/_0_  (.Y(\myring.inv_in[255] ),
    .A(\myring.inv_in[254] ));
 sg13g2_inv_1 \myring.inv_array[255]/sky_inverter/_0_  (.Y(\myring.inv_in[256] ),
    .A(\myring.inv_in[255] ));
 sg13g2_inv_1 \myring.inv_array[256]/sky_inverter/_0_  (.Y(\myring.inv_in[257] ),
    .A(\myring.inv_in[256] ));
 sg13g2_inv_1 \myring.inv_array[257]/sky_inverter/_0_  (.Y(\myring.inv_in[258] ),
    .A(\myring.inv_in[257] ));
 sg13g2_inv_1 \myring.inv_array[258]/sky_inverter/_0_  (.Y(\myring.inv_in[259] ),
    .A(\myring.inv_in[258] ));
 sg13g2_inv_1 \myring.inv_array[259]/sky_inverter/_0_  (.Y(\myring.inv_in[260] ),
    .A(\myring.inv_in[259] ));
 sg13g2_inv_1 \myring.inv_array[25]/sky_inverter/_0_  (.Y(\myring.inv_in[26] ),
    .A(\myring.inv_in[25] ));
 sg13g2_inv_1 \myring.inv_array[260]/sky_inverter/_0_  (.Y(\myring.inv_in[261] ),
    .A(\myring.inv_in[260] ));
 sg13g2_inv_1 \myring.inv_array[261]/sky_inverter/_0_  (.Y(\myring.inv_in[262] ),
    .A(\myring.inv_in[261] ));
 sg13g2_inv_1 \myring.inv_array[262]/sky_inverter/_0_  (.Y(\myring.inv_in[263] ),
    .A(\myring.inv_in[262] ));
 sg13g2_inv_1 \myring.inv_array[263]/sky_inverter/_0_  (.Y(\myring.inv_in[264] ),
    .A(\myring.inv_in[263] ));
 sg13g2_inv_1 \myring.inv_array[264]/sky_inverter/_0_  (.Y(\myring.inv_in[265] ),
    .A(\myring.inv_in[264] ));
 sg13g2_inv_1 \myring.inv_array[265]/sky_inverter/_0_  (.Y(\myring.inv_in[266] ),
    .A(\myring.inv_in[265] ));
 sg13g2_inv_1 \myring.inv_array[266]/sky_inverter/_0_  (.Y(\myring.inv_in[267] ),
    .A(\myring.inv_in[266] ));
 sg13g2_inv_1 \myring.inv_array[267]/sky_inverter/_0_  (.Y(\myring.inv_in[268] ),
    .A(\myring.inv_in[267] ));
 sg13g2_inv_1 \myring.inv_array[268]/sky_inverter/_0_  (.Y(\myring.inv_in[269] ),
    .A(\myring.inv_in[268] ));
 sg13g2_inv_1 \myring.inv_array[269]/sky_inverter/_0_  (.Y(\myring.inv_in[270] ),
    .A(\myring.inv_in[269] ));
 sg13g2_inv_1 \myring.inv_array[26]/sky_inverter/_0_  (.Y(\myring.inv_in[27] ),
    .A(\myring.inv_in[26] ));
 sg13g2_inv_1 \myring.inv_array[270]/sky_inverter/_0_  (.Y(\myring.inv_in[271] ),
    .A(\myring.inv_in[270] ));
 sg13g2_inv_1 \myring.inv_array[271]/sky_inverter/_0_  (.Y(\myring.inv_in[272] ),
    .A(\myring.inv_in[271] ));
 sg13g2_inv_1 \myring.inv_array[272]/sky_inverter/_0_  (.Y(\myring.inv_in[273] ),
    .A(\myring.inv_in[272] ));
 sg13g2_inv_1 \myring.inv_array[273]/sky_inverter/_0_  (.Y(\myring.inv_in[274] ),
    .A(\myring.inv_in[273] ));
 sg13g2_inv_1 \myring.inv_array[274]/sky_inverter/_0_  (.Y(\myring.inv_in[275] ),
    .A(\myring.inv_in[274] ));
 sg13g2_inv_1 \myring.inv_array[275]/sky_inverter/_0_  (.Y(\myring.inv_in[276] ),
    .A(\myring.inv_in[275] ));
 sg13g2_inv_1 \myring.inv_array[276]/sky_inverter/_0_  (.Y(\myring.inv_in[277] ),
    .A(\myring.inv_in[276] ));
 sg13g2_inv_1 \myring.inv_array[277]/sky_inverter/_0_  (.Y(\myring.inv_in[278] ),
    .A(\myring.inv_in[277] ));
 sg13g2_inv_1 \myring.inv_array[278]/sky_inverter/_0_  (.Y(\myring.inv_in[279] ),
    .A(\myring.inv_in[278] ));
 sg13g2_inv_1 \myring.inv_array[279]/sky_inverter/_0_  (.Y(\myring.inv_in[280] ),
    .A(\myring.inv_in[279] ));
 sg13g2_inv_1 \myring.inv_array[27]/sky_inverter/_0_  (.Y(\myring.inv_in[28] ),
    .A(\myring.inv_in[27] ));
 sg13g2_inv_1 \myring.inv_array[280]/sky_inverter/_0_  (.Y(\myring.inv_in[281] ),
    .A(\myring.inv_in[280] ));
 sg13g2_inv_1 \myring.inv_array[281]/sky_inverter/_0_  (.Y(\myring.inv_in[282] ),
    .A(\myring.inv_in[281] ));
 sg13g2_inv_1 \myring.inv_array[282]/sky_inverter/_0_  (.Y(\myring.inv_in[283] ),
    .A(\myring.inv_in[282] ));
 sg13g2_inv_1 \myring.inv_array[283]/sky_inverter/_0_  (.Y(\myring.inv_in[284] ),
    .A(\myring.inv_in[283] ));
 sg13g2_inv_1 \myring.inv_array[284]/sky_inverter/_0_  (.Y(\myring.inv_in[285] ),
    .A(\myring.inv_in[284] ));
 sg13g2_inv_1 \myring.inv_array[285]/sky_inverter/_0_  (.Y(\myring.inv_in[286] ),
    .A(\myring.inv_in[285] ));
 sg13g2_inv_1 \myring.inv_array[286]/sky_inverter/_0_  (.Y(\myring.inv_in[287] ),
    .A(\myring.inv_in[286] ));
 sg13g2_inv_1 \myring.inv_array[287]/sky_inverter/_0_  (.Y(\myring.inv_in[288] ),
    .A(\myring.inv_in[287] ));
 sg13g2_inv_1 \myring.inv_array[288]/sky_inverter/_0_  (.Y(\myring.inv_in[289] ),
    .A(\myring.inv_in[288] ));
 sg13g2_inv_1 \myring.inv_array[289]/sky_inverter/_0_  (.Y(\myring.inv_in[290] ),
    .A(\myring.inv_in[289] ));
 sg13g2_inv_1 \myring.inv_array[28]/sky_inverter/_0_  (.Y(\myring.inv_in[29] ),
    .A(\myring.inv_in[28] ));
 sg13g2_inv_1 \myring.inv_array[290]/sky_inverter/_0_  (.Y(\myring.inv_in[291] ),
    .A(\myring.inv_in[290] ));
 sg13g2_inv_1 \myring.inv_array[291]/sky_inverter/_0_  (.Y(\myring.inv_in[292] ),
    .A(\myring.inv_in[291] ));
 sg13g2_inv_1 \myring.inv_array[292]/sky_inverter/_0_  (.Y(\myring.inv_in[293] ),
    .A(\myring.inv_in[292] ));
 sg13g2_inv_1 \myring.inv_array[293]/sky_inverter/_0_  (.Y(\myring.inv_in[294] ),
    .A(\myring.inv_in[293] ));
 sg13g2_inv_1 \myring.inv_array[294]/sky_inverter/_0_  (.Y(\myring.inv_in[295] ),
    .A(\myring.inv_in[294] ));
 sg13g2_inv_1 \myring.inv_array[295]/sky_inverter/_0_  (.Y(\myring.inv_in[296] ),
    .A(\myring.inv_in[295] ));
 sg13g2_inv_1 \myring.inv_array[296]/sky_inverter/_0_  (.Y(\myring.inv_in[297] ),
    .A(\myring.inv_in[296] ));
 sg13g2_inv_1 \myring.inv_array[297]/sky_inverter/_0_  (.Y(\myring.inv_in[298] ),
    .A(\myring.inv_in[297] ));
 sg13g2_inv_1 \myring.inv_array[298]/sky_inverter/_0_  (.Y(\myring.inv_in[299] ),
    .A(\myring.inv_in[298] ));
 sg13g2_inv_1 \myring.inv_array[299]/sky_inverter/_0_  (.Y(\myring.inv_in[300] ),
    .A(\myring.inv_in[299] ));
 sg13g2_inv_1 \myring.inv_array[29]/sky_inverter/_0_  (.Y(\myring.inv_in[30] ),
    .A(\myring.inv_in[29] ));
 sg13g2_inv_1 \myring.inv_array[2]/sky_inverter/_0_  (.Y(\myring.inv_in[3] ),
    .A(\myring.inv_in[2] ));
 sg13g2_inv_1 \myring.inv_array[300]/sky_inverter/_0_  (.Y(\myring.inv_in[301] ),
    .A(\myring.inv_in[300] ));
 sg13g2_inv_1 \myring.inv_array[301]/sky_inverter/_0_  (.Y(\myring.inv_in[302] ),
    .A(\myring.inv_in[301] ));
 sg13g2_inv_1 \myring.inv_array[302]/sky_inverter/_0_  (.Y(\myring.inv_in[303] ),
    .A(\myring.inv_in[302] ));
 sg13g2_inv_1 \myring.inv_array[303]/sky_inverter/_0_  (.Y(\myring.inv_in[304] ),
    .A(\myring.inv_in[303] ));
 sg13g2_inv_1 \myring.inv_array[304]/sky_inverter/_0_  (.Y(\myring.inv_in[305] ),
    .A(\myring.inv_in[304] ));
 sg13g2_inv_1 \myring.inv_array[305]/sky_inverter/_0_  (.Y(\myring.inv_in[306] ),
    .A(\myring.inv_in[305] ));
 sg13g2_inv_1 \myring.inv_array[306]/sky_inverter/_0_  (.Y(\myring.inv_in[307] ),
    .A(\myring.inv_in[306] ));
 sg13g2_inv_1 \myring.inv_array[307]/sky_inverter/_0_  (.Y(\myring.inv_in[308] ),
    .A(\myring.inv_in[307] ));
 sg13g2_inv_1 \myring.inv_array[308]/sky_inverter/_0_  (.Y(\myring.inv_in[309] ),
    .A(\myring.inv_in[308] ));
 sg13g2_inv_1 \myring.inv_array[309]/sky_inverter/_0_  (.Y(\myring.inv_in[310] ),
    .A(\myring.inv_in[309] ));
 sg13g2_inv_1 \myring.inv_array[30]/sky_inverter/_0_  (.Y(\myring.inv_in[31] ),
    .A(\myring.inv_in[30] ));
 sg13g2_inv_1 \myring.inv_array[310]/sky_inverter/_0_  (.Y(\myring.inv_in[311] ),
    .A(\myring.inv_in[310] ));
 sg13g2_inv_1 \myring.inv_array[311]/sky_inverter/_0_  (.Y(\myring.inv_in[312] ),
    .A(\myring.inv_in[311] ));
 sg13g2_inv_1 \myring.inv_array[312]/sky_inverter/_0_  (.Y(\myring.inv_in[313] ),
    .A(\myring.inv_in[312] ));
 sg13g2_inv_1 \myring.inv_array[313]/sky_inverter/_0_  (.Y(\myring.inv_in[314] ),
    .A(\myring.inv_in[313] ));
 sg13g2_inv_1 \myring.inv_array[314]/sky_inverter/_0_  (.Y(\myring.inv_in[315] ),
    .A(\myring.inv_in[314] ));
 sg13g2_inv_1 \myring.inv_array[315]/sky_inverter/_0_  (.Y(\myring.inv_in[316] ),
    .A(\myring.inv_in[315] ));
 sg13g2_inv_1 \myring.inv_array[316]/sky_inverter/_0_  (.Y(\myring.inv_in[317] ),
    .A(\myring.inv_in[316] ));
 sg13g2_inv_1 \myring.inv_array[317]/sky_inverter/_0_  (.Y(\myring.inv_in[318] ),
    .A(\myring.inv_in[317] ));
 sg13g2_inv_1 \myring.inv_array[318]/sky_inverter/_0_  (.Y(\myring.inv_in[319] ),
    .A(\myring.inv_in[318] ));
 sg13g2_inv_1 \myring.inv_array[319]/sky_inverter/_0_  (.Y(\myring.inv_in[320] ),
    .A(\myring.inv_in[319] ));
 sg13g2_inv_1 \myring.inv_array[31]/sky_inverter/_0_  (.Y(\myring.inv_in[32] ),
    .A(\myring.inv_in[31] ));
 sg13g2_inv_1 \myring.inv_array[320]/sky_inverter/_0_  (.Y(\myring.inv_in[321] ),
    .A(\myring.inv_in[320] ));
 sg13g2_inv_1 \myring.inv_array[321]/sky_inverter/_0_  (.Y(\myring.inv_in[322] ),
    .A(\myring.inv_in[321] ));
 sg13g2_inv_1 \myring.inv_array[322]/sky_inverter/_0_  (.Y(\myring.inv_in[323] ),
    .A(\myring.inv_in[322] ));
 sg13g2_inv_1 \myring.inv_array[323]/sky_inverter/_0_  (.Y(\myring.inv_in[324] ),
    .A(\myring.inv_in[323] ));
 sg13g2_inv_1 \myring.inv_array[324]/sky_inverter/_0_  (.Y(\myring.inv_in[325] ),
    .A(\myring.inv_in[324] ));
 sg13g2_inv_1 \myring.inv_array[325]/sky_inverter/_0_  (.Y(\myring.inv_in[326] ),
    .A(\myring.inv_in[325] ));
 sg13g2_inv_1 \myring.inv_array[326]/sky_inverter/_0_  (.Y(\myring.inv_in[327] ),
    .A(\myring.inv_in[326] ));
 sg13g2_inv_1 \myring.inv_array[327]/sky_inverter/_0_  (.Y(\myring.inv_in[328] ),
    .A(\myring.inv_in[327] ));
 sg13g2_inv_1 \myring.inv_array[328]/sky_inverter/_0_  (.Y(\myring.inv_in[329] ),
    .A(\myring.inv_in[328] ));
 sg13g2_inv_1 \myring.inv_array[329]/sky_inverter/_0_  (.Y(\myring.inv_in[330] ),
    .A(\myring.inv_in[329] ));
 sg13g2_inv_1 \myring.inv_array[32]/sky_inverter/_0_  (.Y(\myring.inv_in[33] ),
    .A(\myring.inv_in[32] ));
 sg13g2_inv_1 \myring.inv_array[330]/sky_inverter/_0_  (.Y(\myring.inv_in[331] ),
    .A(\myring.inv_in[330] ));
 sg13g2_inv_1 \myring.inv_array[331]/sky_inverter/_0_  (.Y(\myring.inv_in[332] ),
    .A(\myring.inv_in[331] ));
 sg13g2_inv_1 \myring.inv_array[332]/sky_inverter/_0_  (.Y(\myring.inv_in[333] ),
    .A(\myring.inv_in[332] ));
 sg13g2_inv_1 \myring.inv_array[333]/sky_inverter/_0_  (.Y(\myring.inv_in[334] ),
    .A(\myring.inv_in[333] ));
 sg13g2_inv_1 \myring.inv_array[334]/sky_inverter/_0_  (.Y(\myring.inv_in[335] ),
    .A(\myring.inv_in[334] ));
 sg13g2_inv_1 \myring.inv_array[335]/sky_inverter/_0_  (.Y(\myring.inv_in[336] ),
    .A(\myring.inv_in[335] ));
 sg13g2_inv_1 \myring.inv_array[336]/sky_inverter/_0_  (.Y(\myring.inv_in[337] ),
    .A(\myring.inv_in[336] ));
 sg13g2_inv_1 \myring.inv_array[337]/sky_inverter/_0_  (.Y(\myring.inv_in[338] ),
    .A(\myring.inv_in[337] ));
 sg13g2_inv_1 \myring.inv_array[338]/sky_inverter/_0_  (.Y(\myring.inv_in[339] ),
    .A(\myring.inv_in[338] ));
 sg13g2_inv_1 \myring.inv_array[339]/sky_inverter/_0_  (.Y(\myring.inv_in[340] ),
    .A(\myring.inv_in[339] ));
 sg13g2_inv_1 \myring.inv_array[33]/sky_inverter/_0_  (.Y(\myring.inv_in[34] ),
    .A(\myring.inv_in[33] ));
 sg13g2_inv_1 \myring.inv_array[340]/sky_inverter/_0_  (.Y(\myring.inv_in[341] ),
    .A(\myring.inv_in[340] ));
 sg13g2_inv_1 \myring.inv_array[341]/sky_inverter/_0_  (.Y(\myring.inv_in[342] ),
    .A(\myring.inv_in[341] ));
 sg13g2_inv_1 \myring.inv_array[342]/sky_inverter/_0_  (.Y(\myring.inv_in[343] ),
    .A(\myring.inv_in[342] ));
 sg13g2_inv_1 \myring.inv_array[343]/sky_inverter/_0_  (.Y(\myring.inv_in[344] ),
    .A(\myring.inv_in[343] ));
 sg13g2_inv_1 \myring.inv_array[344]/sky_inverter/_0_  (.Y(\myring.inv_in[345] ),
    .A(\myring.inv_in[344] ));
 sg13g2_inv_1 \myring.inv_array[345]/sky_inverter/_0_  (.Y(\myring.inv_in[346] ),
    .A(\myring.inv_in[345] ));
 sg13g2_inv_1 \myring.inv_array[346]/sky_inverter/_0_  (.Y(\myring.inv_in[347] ),
    .A(\myring.inv_in[346] ));
 sg13g2_inv_1 \myring.inv_array[347]/sky_inverter/_0_  (.Y(\myring.inv_in[348] ),
    .A(\myring.inv_in[347] ));
 sg13g2_inv_1 \myring.inv_array[348]/sky_inverter/_0_  (.Y(\myring.inv_in[349] ),
    .A(\myring.inv_in[348] ));
 sg13g2_inv_1 \myring.inv_array[349]/sky_inverter/_0_  (.Y(\myring.inv_in[350] ),
    .A(\myring.inv_in[349] ));
 sg13g2_inv_1 \myring.inv_array[34]/sky_inverter/_0_  (.Y(\myring.inv_in[35] ),
    .A(\myring.inv_in[34] ));
 sg13g2_inv_1 \myring.inv_array[350]/sky_inverter/_0_  (.Y(\myring.inv_in[351] ),
    .A(\myring.inv_in[350] ));
 sg13g2_inv_1 \myring.inv_array[351]/sky_inverter/_0_  (.Y(\myring.inv_in[352] ),
    .A(\myring.inv_in[351] ));
 sg13g2_inv_1 \myring.inv_array[352]/sky_inverter/_0_  (.Y(\myring.inv_in[353] ),
    .A(\myring.inv_in[352] ));
 sg13g2_inv_1 \myring.inv_array[353]/sky_inverter/_0_  (.Y(\myring.inv_in[354] ),
    .A(\myring.inv_in[353] ));
 sg13g2_inv_1 \myring.inv_array[354]/sky_inverter/_0_  (.Y(\myring.inv_in[355] ),
    .A(\myring.inv_in[354] ));
 sg13g2_inv_1 \myring.inv_array[355]/sky_inverter/_0_  (.Y(\myring.inv_in[356] ),
    .A(\myring.inv_in[355] ));
 sg13g2_inv_1 \myring.inv_array[356]/sky_inverter/_0_  (.Y(\myring.inv_in[357] ),
    .A(\myring.inv_in[356] ));
 sg13g2_inv_1 \myring.inv_array[357]/sky_inverter/_0_  (.Y(\myring.inv_in[358] ),
    .A(\myring.inv_in[357] ));
 sg13g2_inv_1 \myring.inv_array[358]/sky_inverter/_0_  (.Y(\myring.inv_in[359] ),
    .A(\myring.inv_in[358] ));
 sg13g2_inv_1 \myring.inv_array[359]/sky_inverter/_0_  (.Y(\myring.inv_in[360] ),
    .A(\myring.inv_in[359] ));
 sg13g2_inv_1 \myring.inv_array[35]/sky_inverter/_0_  (.Y(\myring.inv_in[36] ),
    .A(\myring.inv_in[35] ));
 sg13g2_inv_1 \myring.inv_array[360]/sky_inverter/_0_  (.Y(\myring.inv_in[361] ),
    .A(\myring.inv_in[360] ));
 sg13g2_inv_1 \myring.inv_array[361]/sky_inverter/_0_  (.Y(\myring.inv_in[362] ),
    .A(\myring.inv_in[361] ));
 sg13g2_inv_1 \myring.inv_array[362]/sky_inverter/_0_  (.Y(\myring.inv_in[363] ),
    .A(\myring.inv_in[362] ));
 sg13g2_inv_1 \myring.inv_array[363]/sky_inverter/_0_  (.Y(\myring.inv_in[364] ),
    .A(\myring.inv_in[363] ));
 sg13g2_inv_1 \myring.inv_array[364]/sky_inverter/_0_  (.Y(\myring.inv_in[365] ),
    .A(\myring.inv_in[364] ));
 sg13g2_inv_1 \myring.inv_array[365]/sky_inverter/_0_  (.Y(\myring.inv_in[366] ),
    .A(\myring.inv_in[365] ));
 sg13g2_inv_1 \myring.inv_array[366]/sky_inverter/_0_  (.Y(\myring.inv_in[367] ),
    .A(\myring.inv_in[366] ));
 sg13g2_inv_1 \myring.inv_array[367]/sky_inverter/_0_  (.Y(\myring.inv_in[368] ),
    .A(\myring.inv_in[367] ));
 sg13g2_inv_1 \myring.inv_array[368]/sky_inverter/_0_  (.Y(\myring.inv_in[369] ),
    .A(\myring.inv_in[368] ));
 sg13g2_inv_1 \myring.inv_array[369]/sky_inverter/_0_  (.Y(\myring.inv_in[370] ),
    .A(\myring.inv_in[369] ));
 sg13g2_inv_1 \myring.inv_array[36]/sky_inverter/_0_  (.Y(\myring.inv_in[37] ),
    .A(\myring.inv_in[36] ));
 sg13g2_inv_1 \myring.inv_array[370]/sky_inverter/_0_  (.Y(\myring.inv_in[371] ),
    .A(\myring.inv_in[370] ));
 sg13g2_inv_1 \myring.inv_array[371]/sky_inverter/_0_  (.Y(\myring.inv_in[372] ),
    .A(\myring.inv_in[371] ));
 sg13g2_inv_1 \myring.inv_array[372]/sky_inverter/_0_  (.Y(\myring.inv_in[373] ),
    .A(\myring.inv_in[372] ));
 sg13g2_inv_1 \myring.inv_array[373]/sky_inverter/_0_  (.Y(\myring.inv_in[374] ),
    .A(\myring.inv_in[373] ));
 sg13g2_inv_1 \myring.inv_array[374]/sky_inverter/_0_  (.Y(\myring.inv_in[375] ),
    .A(\myring.inv_in[374] ));
 sg13g2_inv_1 \myring.inv_array[375]/sky_inverter/_0_  (.Y(\myring.inv_in[376] ),
    .A(\myring.inv_in[375] ));
 sg13g2_inv_1 \myring.inv_array[376]/sky_inverter/_0_  (.Y(\myring.inv_in[377] ),
    .A(\myring.inv_in[376] ));
 sg13g2_inv_1 \myring.inv_array[377]/sky_inverter/_0_  (.Y(\myring.inv_in[378] ),
    .A(\myring.inv_in[377] ));
 sg13g2_inv_1 \myring.inv_array[378]/sky_inverter/_0_  (.Y(\myring.inv_in[379] ),
    .A(\myring.inv_in[378] ));
 sg13g2_inv_1 \myring.inv_array[379]/sky_inverter/_0_  (.Y(\myring.inv_in[380] ),
    .A(\myring.inv_in[379] ));
 sg13g2_inv_1 \myring.inv_array[37]/sky_inverter/_0_  (.Y(\myring.inv_in[38] ),
    .A(\myring.inv_in[37] ));
 sg13g2_inv_1 \myring.inv_array[380]/sky_inverter/_0_  (.Y(\myring.inv_in[381] ),
    .A(\myring.inv_in[380] ));
 sg13g2_inv_1 \myring.inv_array[381]/sky_inverter/_0_  (.Y(\myring.inv_in[382] ),
    .A(\myring.inv_in[381] ));
 sg13g2_inv_1 \myring.inv_array[382]/sky_inverter/_0_  (.Y(\myring.inv_in[383] ),
    .A(\myring.inv_in[382] ));
 sg13g2_inv_1 \myring.inv_array[383]/sky_inverter/_0_  (.Y(\myring.inv_in[384] ),
    .A(\myring.inv_in[383] ));
 sg13g2_inv_1 \myring.inv_array[384]/sky_inverter/_0_  (.Y(\myring.inv_in[385] ),
    .A(\myring.inv_in[384] ));
 sg13g2_inv_1 \myring.inv_array[385]/sky_inverter/_0_  (.Y(\myring.inv_in[386] ),
    .A(\myring.inv_in[385] ));
 sg13g2_inv_1 \myring.inv_array[386]/sky_inverter/_0_  (.Y(\myring.inv_in[387] ),
    .A(\myring.inv_in[386] ));
 sg13g2_inv_1 \myring.inv_array[387]/sky_inverter/_0_  (.Y(\myring.inv_in[388] ),
    .A(\myring.inv_in[387] ));
 sg13g2_inv_1 \myring.inv_array[388]/sky_inverter/_0_  (.Y(\myring.inv_in[389] ),
    .A(\myring.inv_in[388] ));
 sg13g2_inv_1 \myring.inv_array[389]/sky_inverter/_0_  (.Y(\myring.inv_in[390] ),
    .A(\myring.inv_in[389] ));
 sg13g2_inv_1 \myring.inv_array[38]/sky_inverter/_0_  (.Y(\myring.inv_in[39] ),
    .A(\myring.inv_in[38] ));
 sg13g2_inv_1 \myring.inv_array[390]/sky_inverter/_0_  (.Y(\myring.inv_in[391] ),
    .A(\myring.inv_in[390] ));
 sg13g2_inv_1 \myring.inv_array[391]/sky_inverter/_0_  (.Y(\myring.inv_in[392] ),
    .A(\myring.inv_in[391] ));
 sg13g2_inv_1 \myring.inv_array[392]/sky_inverter/_0_  (.Y(\myring.inv_in[393] ),
    .A(\myring.inv_in[392] ));
 sg13g2_inv_1 \myring.inv_array[393]/sky_inverter/_0_  (.Y(\myring.inv_in[394] ),
    .A(\myring.inv_in[393] ));
 sg13g2_inv_1 \myring.inv_array[394]/sky_inverter/_0_  (.Y(\myring.inv_in[395] ),
    .A(\myring.inv_in[394] ));
 sg13g2_inv_1 \myring.inv_array[395]/sky_inverter/_0_  (.Y(\myring.inv_in[396] ),
    .A(\myring.inv_in[395] ));
 sg13g2_inv_1 \myring.inv_array[396]/sky_inverter/_0_  (.Y(\myring.inv_in[397] ),
    .A(\myring.inv_in[396] ));
 sg13g2_inv_1 \myring.inv_array[397]/sky_inverter/_0_  (.Y(\myring.inv_in[398] ),
    .A(\myring.inv_in[397] ));
 sg13g2_inv_1 \myring.inv_array[398]/sky_inverter/_0_  (.Y(\myring.inv_in[399] ),
    .A(\myring.inv_in[398] ));
 sg13g2_inv_1 \myring.inv_array[399]/sky_inverter/_0_  (.Y(\myring.inv_in[400] ),
    .A(\myring.inv_in[399] ));
 sg13g2_inv_1 \myring.inv_array[39]/sky_inverter/_0_  (.Y(\myring.inv_in[40] ),
    .A(\myring.inv_in[39] ));
 sg13g2_inv_1 \myring.inv_array[3]/sky_inverter/_0_  (.Y(\myring.inv_in[4] ),
    .A(\myring.inv_in[3] ));
 sg13g2_inv_1 \myring.inv_array[400]/sky_inverter/_0_  (.Y(\myring.inv_in[401] ),
    .A(\myring.inv_in[400] ));
 sg13g2_inv_1 \myring.inv_array[401]/sky_inverter/_0_  (.Y(\myring.inv_in[402] ),
    .A(\myring.inv_in[401] ));
 sg13g2_inv_1 \myring.inv_array[402]/sky_inverter/_0_  (.Y(\myring.inv_in[403] ),
    .A(\myring.inv_in[402] ));
 sg13g2_inv_1 \myring.inv_array[403]/sky_inverter/_0_  (.Y(\myring.inv_in[404] ),
    .A(\myring.inv_in[403] ));
 sg13g2_inv_1 \myring.inv_array[404]/sky_inverter/_0_  (.Y(\myring.inv_in[405] ),
    .A(\myring.inv_in[404] ));
 sg13g2_inv_1 \myring.inv_array[405]/sky_inverter/_0_  (.Y(\myring.inv_in[406] ),
    .A(\myring.inv_in[405] ));
 sg13g2_inv_1 \myring.inv_array[406]/sky_inverter/_0_  (.Y(\myring.inv_in[407] ),
    .A(\myring.inv_in[406] ));
 sg13g2_inv_1 \myring.inv_array[407]/sky_inverter/_0_  (.Y(\myring.inv_in[408] ),
    .A(\myring.inv_in[407] ));
 sg13g2_inv_1 \myring.inv_array[408]/sky_inverter/_0_  (.Y(\myring.inv_in[409] ),
    .A(\myring.inv_in[408] ));
 sg13g2_inv_1 \myring.inv_array[409]/sky_inverter/_0_  (.Y(\myring.inv_in[410] ),
    .A(\myring.inv_in[409] ));
 sg13g2_inv_1 \myring.inv_array[40]/sky_inverter/_0_  (.Y(\myring.inv_in[41] ),
    .A(\myring.inv_in[40] ));
 sg13g2_inv_1 \myring.inv_array[410]/sky_inverter/_0_  (.Y(\myring.inv_in[411] ),
    .A(\myring.inv_in[410] ));
 sg13g2_inv_1 \myring.inv_array[411]/sky_inverter/_0_  (.Y(\myring.inv_in[412] ),
    .A(\myring.inv_in[411] ));
 sg13g2_inv_1 \myring.inv_array[412]/sky_inverter/_0_  (.Y(\myring.inv_in[413] ),
    .A(\myring.inv_in[412] ));
 sg13g2_inv_1 \myring.inv_array[413]/sky_inverter/_0_  (.Y(\myring.inv_in[414] ),
    .A(\myring.inv_in[413] ));
 sg13g2_inv_1 \myring.inv_array[414]/sky_inverter/_0_  (.Y(\myring.inv_in[415] ),
    .A(\myring.inv_in[414] ));
 sg13g2_inv_1 \myring.inv_array[415]/sky_inverter/_0_  (.Y(\myring.inv_in[416] ),
    .A(\myring.inv_in[415] ));
 sg13g2_inv_1 \myring.inv_array[416]/sky_inverter/_0_  (.Y(\myring.inv_in[417] ),
    .A(\myring.inv_in[416] ));
 sg13g2_inv_1 \myring.inv_array[417]/sky_inverter/_0_  (.Y(\myring.inv_in[418] ),
    .A(\myring.inv_in[417] ));
 sg13g2_inv_1 \myring.inv_array[418]/sky_inverter/_0_  (.Y(\myring.inv_in[419] ),
    .A(\myring.inv_in[418] ));
 sg13g2_inv_1 \myring.inv_array[419]/sky_inverter/_0_  (.Y(\myring.inv_in[420] ),
    .A(\myring.inv_in[419] ));
 sg13g2_inv_1 \myring.inv_array[41]/sky_inverter/_0_  (.Y(\myring.inv_in[42] ),
    .A(\myring.inv_in[41] ));
 sg13g2_inv_1 \myring.inv_array[420]/sky_inverter/_0_  (.Y(\myring.inv_in[421] ),
    .A(\myring.inv_in[420] ));
 sg13g2_inv_1 \myring.inv_array[421]/sky_inverter/_0_  (.Y(\myring.inv_in[422] ),
    .A(\myring.inv_in[421] ));
 sg13g2_inv_1 \myring.inv_array[422]/sky_inverter/_0_  (.Y(\myring.inv_in[423] ),
    .A(\myring.inv_in[422] ));
 sg13g2_inv_1 \myring.inv_array[423]/sky_inverter/_0_  (.Y(\myring.inv_in[424] ),
    .A(\myring.inv_in[423] ));
 sg13g2_inv_1 \myring.inv_array[424]/sky_inverter/_0_  (.Y(\myring.inv_in[425] ),
    .A(\myring.inv_in[424] ));
 sg13g2_inv_1 \myring.inv_array[425]/sky_inverter/_0_  (.Y(\myring.inv_in[426] ),
    .A(\myring.inv_in[425] ));
 sg13g2_inv_1 \myring.inv_array[426]/sky_inverter/_0_  (.Y(\myring.inv_in[427] ),
    .A(\myring.inv_in[426] ));
 sg13g2_inv_1 \myring.inv_array[427]/sky_inverter/_0_  (.Y(\myring.inv_in[428] ),
    .A(\myring.inv_in[427] ));
 sg13g2_inv_1 \myring.inv_array[428]/sky_inverter/_0_  (.Y(\myring.inv_in[429] ),
    .A(\myring.inv_in[428] ));
 sg13g2_inv_1 \myring.inv_array[429]/sky_inverter/_0_  (.Y(\myring.inv_in[430] ),
    .A(\myring.inv_in[429] ));
 sg13g2_inv_1 \myring.inv_array[42]/sky_inverter/_0_  (.Y(\myring.inv_in[43] ),
    .A(\myring.inv_in[42] ));
 sg13g2_inv_1 \myring.inv_array[430]/sky_inverter/_0_  (.Y(\myring.inv_in[431] ),
    .A(\myring.inv_in[430] ));
 sg13g2_inv_1 \myring.inv_array[431]/sky_inverter/_0_  (.Y(\myring.inv_in[432] ),
    .A(\myring.inv_in[431] ));
 sg13g2_inv_1 \myring.inv_array[432]/sky_inverter/_0_  (.Y(\myring.inv_in[433] ),
    .A(\myring.inv_in[432] ));
 sg13g2_inv_1 \myring.inv_array[433]/sky_inverter/_0_  (.Y(\myring.inv_in[434] ),
    .A(\myring.inv_in[433] ));
 sg13g2_inv_1 \myring.inv_array[434]/sky_inverter/_0_  (.Y(\myring.inv_in[435] ),
    .A(\myring.inv_in[434] ));
 sg13g2_inv_1 \myring.inv_array[435]/sky_inverter/_0_  (.Y(\myring.inv_in[436] ),
    .A(\myring.inv_in[435] ));
 sg13g2_inv_1 \myring.inv_array[436]/sky_inverter/_0_  (.Y(\myring.inv_in[437] ),
    .A(\myring.inv_in[436] ));
 sg13g2_inv_1 \myring.inv_array[437]/sky_inverter/_0_  (.Y(\myring.inv_in[438] ),
    .A(\myring.inv_in[437] ));
 sg13g2_inv_1 \myring.inv_array[438]/sky_inverter/_0_  (.Y(\myring.inv_in[439] ),
    .A(\myring.inv_in[438] ));
 sg13g2_inv_1 \myring.inv_array[439]/sky_inverter/_0_  (.Y(\myring.inv_in[440] ),
    .A(\myring.inv_in[439] ));
 sg13g2_inv_1 \myring.inv_array[43]/sky_inverter/_0_  (.Y(\myring.inv_in[44] ),
    .A(\myring.inv_in[43] ));
 sg13g2_inv_1 \myring.inv_array[440]/sky_inverter/_0_  (.Y(\myring.inv_in[441] ),
    .A(\myring.inv_in[440] ));
 sg13g2_inv_1 \myring.inv_array[441]/sky_inverter/_0_  (.Y(\myring.inv_in[442] ),
    .A(\myring.inv_in[441] ));
 sg13g2_inv_1 \myring.inv_array[442]/sky_inverter/_0_  (.Y(\myring.inv_in[443] ),
    .A(\myring.inv_in[442] ));
 sg13g2_inv_1 \myring.inv_array[443]/sky_inverter/_0_  (.Y(\myring.inv_in[444] ),
    .A(\myring.inv_in[443] ));
 sg13g2_inv_1 \myring.inv_array[444]/sky_inverter/_0_  (.Y(\myring.inv_in[445] ),
    .A(\myring.inv_in[444] ));
 sg13g2_inv_1 \myring.inv_array[445]/sky_inverter/_0_  (.Y(\myring.inv_in[446] ),
    .A(\myring.inv_in[445] ));
 sg13g2_inv_1 \myring.inv_array[446]/sky_inverter/_0_  (.Y(\myring.inv_in[447] ),
    .A(\myring.inv_in[446] ));
 sg13g2_inv_1 \myring.inv_array[447]/sky_inverter/_0_  (.Y(\myring.inv_in[448] ),
    .A(\myring.inv_in[447] ));
 sg13g2_inv_1 \myring.inv_array[448]/sky_inverter/_0_  (.Y(\myring.inv_in[449] ),
    .A(\myring.inv_in[448] ));
 sg13g2_inv_1 \myring.inv_array[449]/sky_inverter/_0_  (.Y(\myring.inv_in[450] ),
    .A(\myring.inv_in[449] ));
 sg13g2_inv_1 \myring.inv_array[44]/sky_inverter/_0_  (.Y(\myring.inv_in[45] ),
    .A(\myring.inv_in[44] ));
 sg13g2_inv_1 \myring.inv_array[450]/sky_inverter/_0_  (.Y(\myring.inv_in[451] ),
    .A(\myring.inv_in[450] ));
 sg13g2_inv_1 \myring.inv_array[451]/sky_inverter/_0_  (.Y(\myring.inv_in[452] ),
    .A(\myring.inv_in[451] ));
 sg13g2_inv_1 \myring.inv_array[452]/sky_inverter/_0_  (.Y(\myring.inv_in[453] ),
    .A(\myring.inv_in[452] ));
 sg13g2_inv_1 \myring.inv_array[453]/sky_inverter/_0_  (.Y(\myring.inv_in[454] ),
    .A(\myring.inv_in[453] ));
 sg13g2_inv_1 \myring.inv_array[454]/sky_inverter/_0_  (.Y(\myring.inv_in[455] ),
    .A(\myring.inv_in[454] ));
 sg13g2_inv_1 \myring.inv_array[455]/sky_inverter/_0_  (.Y(\myring.inv_in[456] ),
    .A(\myring.inv_in[455] ));
 sg13g2_inv_1 \myring.inv_array[456]/sky_inverter/_0_  (.Y(\myring.inv_in[457] ),
    .A(\myring.inv_in[456] ));
 sg13g2_inv_1 \myring.inv_array[457]/sky_inverter/_0_  (.Y(\myring.inv_in[458] ),
    .A(\myring.inv_in[457] ));
 sg13g2_inv_1 \myring.inv_array[458]/sky_inverter/_0_  (.Y(\myring.inv_in[459] ),
    .A(\myring.inv_in[458] ));
 sg13g2_inv_1 \myring.inv_array[459]/sky_inverter/_0_  (.Y(\myring.inv_in[460] ),
    .A(\myring.inv_in[459] ));
 sg13g2_inv_1 \myring.inv_array[45]/sky_inverter/_0_  (.Y(\myring.inv_in[46] ),
    .A(\myring.inv_in[45] ));
 sg13g2_inv_1 \myring.inv_array[460]/sky_inverter/_0_  (.Y(\myring.inv_in[461] ),
    .A(\myring.inv_in[460] ));
 sg13g2_inv_1 \myring.inv_array[461]/sky_inverter/_0_  (.Y(\myring.inv_in[462] ),
    .A(\myring.inv_in[461] ));
 sg13g2_inv_1 \myring.inv_array[462]/sky_inverter/_0_  (.Y(\myring.inv_in[463] ),
    .A(\myring.inv_in[462] ));
 sg13g2_inv_1 \myring.inv_array[463]/sky_inverter/_0_  (.Y(\myring.inv_in[464] ),
    .A(\myring.inv_in[463] ));
 sg13g2_inv_1 \myring.inv_array[464]/sky_inverter/_0_  (.Y(\myring.inv_in[465] ),
    .A(\myring.inv_in[464] ));
 sg13g2_inv_1 \myring.inv_array[465]/sky_inverter/_0_  (.Y(\myring.inv_in[466] ),
    .A(\myring.inv_in[465] ));
 sg13g2_inv_1 \myring.inv_array[466]/sky_inverter/_0_  (.Y(\myring.inv_in[467] ),
    .A(\myring.inv_in[466] ));
 sg13g2_inv_1 \myring.inv_array[467]/sky_inverter/_0_  (.Y(\myring.inv_in[468] ),
    .A(\myring.inv_in[467] ));
 sg13g2_inv_1 \myring.inv_array[468]/sky_inverter/_0_  (.Y(\myring.inv_in[469] ),
    .A(\myring.inv_in[468] ));
 sg13g2_inv_1 \myring.inv_array[469]/sky_inverter/_0_  (.Y(\myring.inv_in[470] ),
    .A(\myring.inv_in[469] ));
 sg13g2_inv_1 \myring.inv_array[46]/sky_inverter/_0_  (.Y(\myring.inv_in[47] ),
    .A(\myring.inv_in[46] ));
 sg13g2_inv_1 \myring.inv_array[470]/sky_inverter/_0_  (.Y(\myring.inv_in[471] ),
    .A(\myring.inv_in[470] ));
 sg13g2_inv_1 \myring.inv_array[471]/sky_inverter/_0_  (.Y(\myring.inv_in[472] ),
    .A(\myring.inv_in[471] ));
 sg13g2_inv_1 \myring.inv_array[472]/sky_inverter/_0_  (.Y(\myring.inv_in[473] ),
    .A(\myring.inv_in[472] ));
 sg13g2_inv_1 \myring.inv_array[473]/sky_inverter/_0_  (.Y(\myring.inv_in[474] ),
    .A(\myring.inv_in[473] ));
 sg13g2_inv_1 \myring.inv_array[474]/sky_inverter/_0_  (.Y(\myring.inv_in[475] ),
    .A(\myring.inv_in[474] ));
 sg13g2_inv_1 \myring.inv_array[475]/sky_inverter/_0_  (.Y(\myring.inv_in[476] ),
    .A(\myring.inv_in[475] ));
 sg13g2_inv_1 \myring.inv_array[476]/sky_inverter/_0_  (.Y(\myring.inv_in[477] ),
    .A(\myring.inv_in[476] ));
 sg13g2_inv_1 \myring.inv_array[477]/sky_inverter/_0_  (.Y(\myring.inv_in[478] ),
    .A(\myring.inv_in[477] ));
 sg13g2_inv_1 \myring.inv_array[478]/sky_inverter/_0_  (.Y(\myring.inv_in[479] ),
    .A(\myring.inv_in[478] ));
 sg13g2_inv_1 \myring.inv_array[479]/sky_inverter/_0_  (.Y(\myring.inv_in[480] ),
    .A(\myring.inv_in[479] ));
 sg13g2_inv_1 \myring.inv_array[47]/sky_inverter/_0_  (.Y(\myring.inv_in[48] ),
    .A(\myring.inv_in[47] ));
 sg13g2_inv_1 \myring.inv_array[480]/sky_inverter/_0_  (.Y(\myring.inv_in[481] ),
    .A(\myring.inv_in[480] ));
 sg13g2_inv_1 \myring.inv_array[481]/sky_inverter/_0_  (.Y(\myring.inv_in[482] ),
    .A(\myring.inv_in[481] ));
 sg13g2_inv_1 \myring.inv_array[482]/sky_inverter/_0_  (.Y(\myring.inv_in[483] ),
    .A(\myring.inv_in[482] ));
 sg13g2_inv_1 \myring.inv_array[483]/sky_inverter/_0_  (.Y(\myring.inv_in[484] ),
    .A(\myring.inv_in[483] ));
 sg13g2_inv_1 \myring.inv_array[484]/sky_inverter/_0_  (.Y(\myring.inv_in[485] ),
    .A(\myring.inv_in[484] ));
 sg13g2_inv_1 \myring.inv_array[485]/sky_inverter/_0_  (.Y(\myring.inv_in[486] ),
    .A(\myring.inv_in[485] ));
 sg13g2_inv_1 \myring.inv_array[486]/sky_inverter/_0_  (.Y(\myring.inv_in[487] ),
    .A(\myring.inv_in[486] ));
 sg13g2_inv_1 \myring.inv_array[487]/sky_inverter/_0_  (.Y(\myring.inv_in[488] ),
    .A(\myring.inv_in[487] ));
 sg13g2_inv_1 \myring.inv_array[488]/sky_inverter/_0_  (.Y(\myring.inv_in[489] ),
    .A(\myring.inv_in[488] ));
 sg13g2_inv_1 \myring.inv_array[489]/sky_inverter/_0_  (.Y(\myring.inv_in[490] ),
    .A(\myring.inv_in[489] ));
 sg13g2_inv_1 \myring.inv_array[48]/sky_inverter/_0_  (.Y(\myring.inv_in[49] ),
    .A(\myring.inv_in[48] ));
 sg13g2_inv_1 \myring.inv_array[490]/sky_inverter/_0_  (.Y(\myring.inv_in[491] ),
    .A(\myring.inv_in[490] ));
 sg13g2_inv_1 \myring.inv_array[491]/sky_inverter/_0_  (.Y(\myring.inv_in[492] ),
    .A(\myring.inv_in[491] ));
 sg13g2_inv_1 \myring.inv_array[492]/sky_inverter/_0_  (.Y(\myring.inv_in[493] ),
    .A(\myring.inv_in[492] ));
 sg13g2_inv_1 \myring.inv_array[493]/sky_inverter/_0_  (.Y(\myring.inv_in[494] ),
    .A(\myring.inv_in[493] ));
 sg13g2_inv_1 \myring.inv_array[494]/sky_inverter/_0_  (.Y(\myring.inv_in[495] ),
    .A(\myring.inv_in[494] ));
 sg13g2_inv_1 \myring.inv_array[495]/sky_inverter/_0_  (.Y(\myring.inv_in[496] ),
    .A(\myring.inv_in[495] ));
 sg13g2_inv_1 \myring.inv_array[496]/sky_inverter/_0_  (.Y(\myring.inv_in[497] ),
    .A(\myring.inv_in[496] ));
 sg13g2_inv_1 \myring.inv_array[497]/sky_inverter/_0_  (.Y(\myring.inv_in[498] ),
    .A(\myring.inv_in[497] ));
 sg13g2_inv_1 \myring.inv_array[498]/sky_inverter/_0_  (.Y(\myring.inv_in[499] ),
    .A(\myring.inv_in[498] ));
 sg13g2_inv_1 \myring.inv_array[499]/sky_inverter/_0_  (.Y(\myring.inv_in[500] ),
    .A(\myring.inv_in[499] ));
 sg13g2_inv_1 \myring.inv_array[49]/sky_inverter/_0_  (.Y(\myring.inv_in[50] ),
    .A(\myring.inv_in[49] ));
 sg13g2_inv_1 \myring.inv_array[4]/sky_inverter/_0_  (.Y(\myring.inv_in[5] ),
    .A(\myring.inv_in[4] ));
 sg13g2_inv_1 \myring.inv_array[500]/sky_inverter/_0_  (.Y(\myring.inv_in[501] ),
    .A(\myring.inv_in[500] ));
 sg13g2_inv_1 \myring.inv_array[501]/sky_inverter/_0_  (.Y(\myring.inv_in[502] ),
    .A(\myring.inv_in[501] ));
 sg13g2_inv_1 \myring.inv_array[502]/sky_inverter/_0_  (.Y(\myring.inv_in[503] ),
    .A(\myring.inv_in[502] ));
 sg13g2_inv_1 \myring.inv_array[503]/sky_inverter/_0_  (.Y(\myring.inv_in[504] ),
    .A(\myring.inv_in[503] ));
 sg13g2_inv_1 \myring.inv_array[504]/sky_inverter/_0_  (.Y(\myring.inv_in[505] ),
    .A(\myring.inv_in[504] ));
 sg13g2_inv_1 \myring.inv_array[505]/sky_inverter/_0_  (.Y(\myring.inv_in[506] ),
    .A(\myring.inv_in[505] ));
 sg13g2_inv_1 \myring.inv_array[506]/sky_inverter/_0_  (.Y(\myring.inv_in[507] ),
    .A(\myring.inv_in[506] ));
 sg13g2_inv_1 \myring.inv_array[507]/sky_inverter/_0_  (.Y(\myring.inv_in[508] ),
    .A(\myring.inv_in[507] ));
 sg13g2_inv_1 \myring.inv_array[508]/sky_inverter/_0_  (.Y(\myring.inv_in[509] ),
    .A(\myring.inv_in[508] ));
 sg13g2_inv_1 \myring.inv_array[509]/sky_inverter/_0_  (.Y(\myring.inv_in[510] ),
    .A(\myring.inv_in[509] ));
 sg13g2_inv_1 \myring.inv_array[50]/sky_inverter/_0_  (.Y(\myring.inv_in[51] ),
    .A(\myring.inv_in[50] ));
 sg13g2_inv_1 \myring.inv_array[510]/sky_inverter/_0_  (.Y(\myring.inv_in[511] ),
    .A(\myring.inv_in[510] ));
 sg13g2_inv_1 \myring.inv_array[511]/sky_inverter/_0_  (.Y(\myring.inv_in[512] ),
    .A(\myring.inv_in[511] ));
 sg13g2_inv_1 \myring.inv_array[512]/sky_inverter/_0_  (.Y(\myring.inv_in[513] ),
    .A(\myring.inv_in[512] ));
 sg13g2_inv_1 \myring.inv_array[513]/sky_inverter/_0_  (.Y(\myring.inv_in[514] ),
    .A(\myring.inv_in[513] ));
 sg13g2_inv_1 \myring.inv_array[514]/sky_inverter/_0_  (.Y(\myring.inv_in[515] ),
    .A(\myring.inv_in[514] ));
 sg13g2_inv_1 \myring.inv_array[515]/sky_inverter/_0_  (.Y(\myring.inv_in[516] ),
    .A(\myring.inv_in[515] ));
 sg13g2_inv_1 \myring.inv_array[516]/sky_inverter/_0_  (.Y(\myring.inv_in[517] ),
    .A(\myring.inv_in[516] ));
 sg13g2_inv_1 \myring.inv_array[517]/sky_inverter/_0_  (.Y(\myring.inv_in[518] ),
    .A(\myring.inv_in[517] ));
 sg13g2_inv_1 \myring.inv_array[518]/sky_inverter/_0_  (.Y(\myring.inv_in[519] ),
    .A(\myring.inv_in[518] ));
 sg13g2_inv_1 \myring.inv_array[519]/sky_inverter/_0_  (.Y(\myring.inv_in[520] ),
    .A(\myring.inv_in[519] ));
 sg13g2_inv_1 \myring.inv_array[51]/sky_inverter/_0_  (.Y(\myring.inv_in[52] ),
    .A(\myring.inv_in[51] ));
 sg13g2_inv_1 \myring.inv_array[520]/sky_inverter/_0_  (.Y(\myring.inv_in[521] ),
    .A(\myring.inv_in[520] ));
 sg13g2_inv_1 \myring.inv_array[521]/sky_inverter/_0_  (.Y(\myring.inv_in[522] ),
    .A(\myring.inv_in[521] ));
 sg13g2_inv_1 \myring.inv_array[522]/sky_inverter/_0_  (.Y(\myring.inv_in[523] ),
    .A(\myring.inv_in[522] ));
 sg13g2_inv_1 \myring.inv_array[523]/sky_inverter/_0_  (.Y(\myring.inv_in[524] ),
    .A(\myring.inv_in[523] ));
 sg13g2_inv_1 \myring.inv_array[524]/sky_inverter/_0_  (.Y(\myring.inv_in[525] ),
    .A(\myring.inv_in[524] ));
 sg13g2_inv_1 \myring.inv_array[525]/sky_inverter/_0_  (.Y(\myring.inv_in[526] ),
    .A(\myring.inv_in[525] ));
 sg13g2_inv_1 \myring.inv_array[526]/sky_inverter/_0_  (.Y(\myring.inv_in[527] ),
    .A(\myring.inv_in[526] ));
 sg13g2_inv_1 \myring.inv_array[527]/sky_inverter/_0_  (.Y(\myring.inv_in[528] ),
    .A(\myring.inv_in[527] ));
 sg13g2_inv_1 \myring.inv_array[528]/sky_inverter/_0_  (.Y(\myring.inv_in[529] ),
    .A(\myring.inv_in[528] ));
 sg13g2_inv_1 \myring.inv_array[529]/sky_inverter/_0_  (.Y(\myring.inv_in[530] ),
    .A(\myring.inv_in[529] ));
 sg13g2_inv_1 \myring.inv_array[52]/sky_inverter/_0_  (.Y(\myring.inv_in[53] ),
    .A(\myring.inv_in[52] ));
 sg13g2_inv_1 \myring.inv_array[530]/sky_inverter/_0_  (.Y(\myring.inv_in[531] ),
    .A(\myring.inv_in[530] ));
 sg13g2_inv_1 \myring.inv_array[531]/sky_inverter/_0_  (.Y(\myring.inv_in[532] ),
    .A(\myring.inv_in[531] ));
 sg13g2_inv_1 \myring.inv_array[532]/sky_inverter/_0_  (.Y(\myring.inv_in[533] ),
    .A(\myring.inv_in[532] ));
 sg13g2_inv_1 \myring.inv_array[533]/sky_inverter/_0_  (.Y(\myring.inv_in[534] ),
    .A(\myring.inv_in[533] ));
 sg13g2_inv_1 \myring.inv_array[534]/sky_inverter/_0_  (.Y(\myring.inv_in[535] ),
    .A(\myring.inv_in[534] ));
 sg13g2_inv_1 \myring.inv_array[535]/sky_inverter/_0_  (.Y(\myring.inv_in[536] ),
    .A(\myring.inv_in[535] ));
 sg13g2_inv_1 \myring.inv_array[536]/sky_inverter/_0_  (.Y(\myring.inv_in[537] ),
    .A(\myring.inv_in[536] ));
 sg13g2_inv_1 \myring.inv_array[537]/sky_inverter/_0_  (.Y(\myring.inv_in[538] ),
    .A(\myring.inv_in[537] ));
 sg13g2_inv_1 \myring.inv_array[538]/sky_inverter/_0_  (.Y(\myring.inv_in[539] ),
    .A(\myring.inv_in[538] ));
 sg13g2_inv_1 \myring.inv_array[539]/sky_inverter/_0_  (.Y(\myring.inv_in[540] ),
    .A(\myring.inv_in[539] ));
 sg13g2_inv_1 \myring.inv_array[53]/sky_inverter/_0_  (.Y(\myring.inv_in[54] ),
    .A(\myring.inv_in[53] ));
 sg13g2_inv_1 \myring.inv_array[540]/sky_inverter/_0_  (.Y(\myring.inv_in[541] ),
    .A(\myring.inv_in[540] ));
 sg13g2_inv_1 \myring.inv_array[541]/sky_inverter/_0_  (.Y(\myring.inv_in[542] ),
    .A(\myring.inv_in[541] ));
 sg13g2_inv_1 \myring.inv_array[542]/sky_inverter/_0_  (.Y(\myring.inv_in[543] ),
    .A(\myring.inv_in[542] ));
 sg13g2_inv_1 \myring.inv_array[543]/sky_inverter/_0_  (.Y(\myring.inv_in[544] ),
    .A(\myring.inv_in[543] ));
 sg13g2_inv_1 \myring.inv_array[544]/sky_inverter/_0_  (.Y(\myring.inv_in[545] ),
    .A(\myring.inv_in[544] ));
 sg13g2_inv_1 \myring.inv_array[545]/sky_inverter/_0_  (.Y(\myring.inv_in[546] ),
    .A(\myring.inv_in[545] ));
 sg13g2_inv_1 \myring.inv_array[546]/sky_inverter/_0_  (.Y(\myring.inv_in[547] ),
    .A(\myring.inv_in[546] ));
 sg13g2_inv_1 \myring.inv_array[547]/sky_inverter/_0_  (.Y(\myring.inv_in[548] ),
    .A(\myring.inv_in[547] ));
 sg13g2_inv_1 \myring.inv_array[548]/sky_inverter/_0_  (.Y(\myring.inv_in[549] ),
    .A(\myring.inv_in[548] ));
 sg13g2_inv_1 \myring.inv_array[549]/sky_inverter/_0_  (.Y(\myring.inv_in[550] ),
    .A(\myring.inv_in[549] ));
 sg13g2_inv_1 \myring.inv_array[54]/sky_inverter/_0_  (.Y(\myring.inv_in[55] ),
    .A(\myring.inv_in[54] ));
 sg13g2_inv_1 \myring.inv_array[550]/sky_inverter/_0_  (.Y(\myring.inv_in[551] ),
    .A(\myring.inv_in[550] ));
 sg13g2_inv_1 \myring.inv_array[551]/sky_inverter/_0_  (.Y(\myring.inv_in[552] ),
    .A(\myring.inv_in[551] ));
 sg13g2_inv_1 \myring.inv_array[552]/sky_inverter/_0_  (.Y(\myring.inv_in[553] ),
    .A(\myring.inv_in[552] ));
 sg13g2_inv_1 \myring.inv_array[553]/sky_inverter/_0_  (.Y(\myring.inv_in[554] ),
    .A(\myring.inv_in[553] ));
 sg13g2_inv_1 \myring.inv_array[554]/sky_inverter/_0_  (.Y(\myring.inv_in[555] ),
    .A(\myring.inv_in[554] ));
 sg13g2_inv_1 \myring.inv_array[555]/sky_inverter/_0_  (.Y(\myring.inv_in[556] ),
    .A(\myring.inv_in[555] ));
 sg13g2_inv_1 \myring.inv_array[556]/sky_inverter/_0_  (.Y(\myring.inv_in[557] ),
    .A(\myring.inv_in[556] ));
 sg13g2_inv_1 \myring.inv_array[557]/sky_inverter/_0_  (.Y(\myring.inv_in[558] ),
    .A(\myring.inv_in[557] ));
 sg13g2_inv_1 \myring.inv_array[558]/sky_inverter/_0_  (.Y(\myring.inv_in[559] ),
    .A(\myring.inv_in[558] ));
 sg13g2_inv_1 \myring.inv_array[559]/sky_inverter/_0_  (.Y(\myring.inv_in[560] ),
    .A(\myring.inv_in[559] ));
 sg13g2_inv_1 \myring.inv_array[55]/sky_inverter/_0_  (.Y(\myring.inv_in[56] ),
    .A(\myring.inv_in[55] ));
 sg13g2_inv_1 \myring.inv_array[560]/sky_inverter/_0_  (.Y(\myring.inv_in[561] ),
    .A(\myring.inv_in[560] ));
 sg13g2_inv_1 \myring.inv_array[561]/sky_inverter/_0_  (.Y(\myring.inv_in[562] ),
    .A(\myring.inv_in[561] ));
 sg13g2_inv_1 \myring.inv_array[562]/sky_inverter/_0_  (.Y(\myring.inv_in[563] ),
    .A(\myring.inv_in[562] ));
 sg13g2_inv_1 \myring.inv_array[563]/sky_inverter/_0_  (.Y(\myring.inv_in[564] ),
    .A(\myring.inv_in[563] ));
 sg13g2_inv_1 \myring.inv_array[564]/sky_inverter/_0_  (.Y(\myring.inv_in[565] ),
    .A(\myring.inv_in[564] ));
 sg13g2_inv_1 \myring.inv_array[565]/sky_inverter/_0_  (.Y(\myring.inv_in[566] ),
    .A(\myring.inv_in[565] ));
 sg13g2_inv_1 \myring.inv_array[566]/sky_inverter/_0_  (.Y(\myring.inv_in[567] ),
    .A(\myring.inv_in[566] ));
 sg13g2_inv_1 \myring.inv_array[567]/sky_inverter/_0_  (.Y(\myring.inv_in[568] ),
    .A(\myring.inv_in[567] ));
 sg13g2_inv_1 \myring.inv_array[568]/sky_inverter/_0_  (.Y(\myring.inv_in[569] ),
    .A(\myring.inv_in[568] ));
 sg13g2_inv_1 \myring.inv_array[569]/sky_inverter/_0_  (.Y(\myring.inv_in[570] ),
    .A(\myring.inv_in[569] ));
 sg13g2_inv_1 \myring.inv_array[56]/sky_inverter/_0_  (.Y(\myring.inv_in[57] ),
    .A(\myring.inv_in[56] ));
 sg13g2_inv_1 \myring.inv_array[570]/sky_inverter/_0_  (.Y(\myring.inv_in[571] ),
    .A(\myring.inv_in[570] ));
 sg13g2_inv_1 \myring.inv_array[571]/sky_inverter/_0_  (.Y(\myring.inv_in[572] ),
    .A(\myring.inv_in[571] ));
 sg13g2_inv_1 \myring.inv_array[572]/sky_inverter/_0_  (.Y(\myring.inv_in[573] ),
    .A(\myring.inv_in[572] ));
 sg13g2_inv_1 \myring.inv_array[573]/sky_inverter/_0_  (.Y(\myring.inv_in[574] ),
    .A(\myring.inv_in[573] ));
 sg13g2_inv_1 \myring.inv_array[574]/sky_inverter/_0_  (.Y(\myring.inv_in[575] ),
    .A(\myring.inv_in[574] ));
 sg13g2_inv_1 \myring.inv_array[575]/sky_inverter/_0_  (.Y(\myring.inv_in[576] ),
    .A(\myring.inv_in[575] ));
 sg13g2_inv_1 \myring.inv_array[576]/sky_inverter/_0_  (.Y(\myring.inv_in[577] ),
    .A(\myring.inv_in[576] ));
 sg13g2_inv_1 \myring.inv_array[577]/sky_inverter/_0_  (.Y(\myring.inv_in[578] ),
    .A(\myring.inv_in[577] ));
 sg13g2_inv_1 \myring.inv_array[578]/sky_inverter/_0_  (.Y(\myring.inv_in[579] ),
    .A(\myring.inv_in[578] ));
 sg13g2_inv_1 \myring.inv_array[579]/sky_inverter/_0_  (.Y(\myring.inv_in[580] ),
    .A(\myring.inv_in[579] ));
 sg13g2_inv_1 \myring.inv_array[57]/sky_inverter/_0_  (.Y(\myring.inv_in[58] ),
    .A(\myring.inv_in[57] ));
 sg13g2_inv_1 \myring.inv_array[580]/sky_inverter/_0_  (.Y(\myring.inv_in[581] ),
    .A(\myring.inv_in[580] ));
 sg13g2_inv_1 \myring.inv_array[581]/sky_inverter/_0_  (.Y(\myring.inv_in[582] ),
    .A(\myring.inv_in[581] ));
 sg13g2_inv_1 \myring.inv_array[582]/sky_inverter/_0_  (.Y(\myring.inv_in[583] ),
    .A(\myring.inv_in[582] ));
 sg13g2_inv_1 \myring.inv_array[583]/sky_inverter/_0_  (.Y(\myring.inv_in[584] ),
    .A(\myring.inv_in[583] ));
 sg13g2_inv_1 \myring.inv_array[584]/sky_inverter/_0_  (.Y(\myring.inv_in[585] ),
    .A(\myring.inv_in[584] ));
 sg13g2_inv_1 \myring.inv_array[585]/sky_inverter/_0_  (.Y(\myring.inv_in[586] ),
    .A(\myring.inv_in[585] ));
 sg13g2_inv_1 \myring.inv_array[586]/sky_inverter/_0_  (.Y(\myring.inv_in[587] ),
    .A(\myring.inv_in[586] ));
 sg13g2_inv_1 \myring.inv_array[587]/sky_inverter/_0_  (.Y(\myring.inv_in[588] ),
    .A(\myring.inv_in[587] ));
 sg13g2_inv_1 \myring.inv_array[588]/sky_inverter/_0_  (.Y(\myring.inv_in[589] ),
    .A(\myring.inv_in[588] ));
 sg13g2_inv_1 \myring.inv_array[589]/sky_inverter/_0_  (.Y(\myring.inv_in[590] ),
    .A(\myring.inv_in[589] ));
 sg13g2_inv_1 \myring.inv_array[58]/sky_inverter/_0_  (.Y(\myring.inv_in[59] ),
    .A(\myring.inv_in[58] ));
 sg13g2_inv_1 \myring.inv_array[590]/sky_inverter/_0_  (.Y(\myring.inv_in[591] ),
    .A(\myring.inv_in[590] ));
 sg13g2_inv_1 \myring.inv_array[591]/sky_inverter/_0_  (.Y(\myring.inv_in[592] ),
    .A(\myring.inv_in[591] ));
 sg13g2_inv_1 \myring.inv_array[592]/sky_inverter/_0_  (.Y(\myring.inv_in[593] ),
    .A(\myring.inv_in[592] ));
 sg13g2_inv_1 \myring.inv_array[593]/sky_inverter/_0_  (.Y(\myring.inv_in[594] ),
    .A(\myring.inv_in[593] ));
 sg13g2_inv_1 \myring.inv_array[594]/sky_inverter/_0_  (.Y(\myring.inv_in[595] ),
    .A(\myring.inv_in[594] ));
 sg13g2_inv_1 \myring.inv_array[595]/sky_inverter/_0_  (.Y(\myring.inv_in[596] ),
    .A(\myring.inv_in[595] ));
 sg13g2_inv_1 \myring.inv_array[596]/sky_inverter/_0_  (.Y(\myring.inv_in[597] ),
    .A(\myring.inv_in[596] ));
 sg13g2_inv_1 \myring.inv_array[597]/sky_inverter/_0_  (.Y(\myring.inv_in[598] ),
    .A(\myring.inv_in[597] ));
 sg13g2_inv_1 \myring.inv_array[598]/sky_inverter/_0_  (.Y(\myring.inv_in[599] ),
    .A(\myring.inv_in[598] ));
 sg13g2_inv_1 \myring.inv_array[599]/sky_inverter/_0_  (.Y(\myring.inv_in[600] ),
    .A(\myring.inv_in[599] ));
 sg13g2_inv_1 \myring.inv_array[59]/sky_inverter/_0_  (.Y(\myring.inv_in[60] ),
    .A(\myring.inv_in[59] ));
 sg13g2_inv_1 \myring.inv_array[5]/sky_inverter/_0_  (.Y(\myring.inv_in[6] ),
    .A(\myring.inv_in[5] ));
 sg13g2_inv_1 \myring.inv_array[600]/sky_inverter/_0_  (.Y(\myring.inv_in[601] ),
    .A(\myring.inv_in[600] ));
 sg13g2_inv_1 \myring.inv_array[601]/sky_inverter/_0_  (.Y(\myring.inv_in[602] ),
    .A(\myring.inv_in[601] ));
 sg13g2_inv_1 \myring.inv_array[602]/sky_inverter/_0_  (.Y(\myring.inv_in[603] ),
    .A(\myring.inv_in[602] ));
 sg13g2_inv_1 \myring.inv_array[603]/sky_inverter/_0_  (.Y(\myring.inv_in[604] ),
    .A(\myring.inv_in[603] ));
 sg13g2_inv_1 \myring.inv_array[604]/sky_inverter/_0_  (.Y(\myring.inv_in[605] ),
    .A(\myring.inv_in[604] ));
 sg13g2_inv_1 \myring.inv_array[605]/sky_inverter/_0_  (.Y(\myring.inv_in[606] ),
    .A(\myring.inv_in[605] ));
 sg13g2_inv_1 \myring.inv_array[606]/sky_inverter/_0_  (.Y(\myring.inv_in[607] ),
    .A(\myring.inv_in[606] ));
 sg13g2_inv_1 \myring.inv_array[607]/sky_inverter/_0_  (.Y(\myring.inv_in[608] ),
    .A(\myring.inv_in[607] ));
 sg13g2_inv_1 \myring.inv_array[608]/sky_inverter/_0_  (.Y(\myring.inv_in[609] ),
    .A(\myring.inv_in[608] ));
 sg13g2_inv_1 \myring.inv_array[609]/sky_inverter/_0_  (.Y(\myring.inv_in[610] ),
    .A(\myring.inv_in[609] ));
 sg13g2_inv_1 \myring.inv_array[60]/sky_inverter/_0_  (.Y(\myring.inv_in[61] ),
    .A(\myring.inv_in[60] ));
 sg13g2_inv_1 \myring.inv_array[610]/sky_inverter/_0_  (.Y(\myring.inv_in[611] ),
    .A(\myring.inv_in[610] ));
 sg13g2_inv_1 \myring.inv_array[611]/sky_inverter/_0_  (.Y(\myring.inv_in[612] ),
    .A(\myring.inv_in[611] ));
 sg13g2_inv_1 \myring.inv_array[612]/sky_inverter/_0_  (.Y(\myring.inv_in[613] ),
    .A(\myring.inv_in[612] ));
 sg13g2_inv_1 \myring.inv_array[613]/sky_inverter/_0_  (.Y(\myring.inv_in[614] ),
    .A(\myring.inv_in[613] ));
 sg13g2_inv_1 \myring.inv_array[614]/sky_inverter/_0_  (.Y(\myring.inv_in[615] ),
    .A(\myring.inv_in[614] ));
 sg13g2_inv_1 \myring.inv_array[615]/sky_inverter/_0_  (.Y(\myring.inv_in[616] ),
    .A(\myring.inv_in[615] ));
 sg13g2_inv_1 \myring.inv_array[616]/sky_inverter/_0_  (.Y(\myring.inv_in[617] ),
    .A(\myring.inv_in[616] ));
 sg13g2_inv_1 \myring.inv_array[617]/sky_inverter/_0_  (.Y(\myring.inv_in[618] ),
    .A(\myring.inv_in[617] ));
 sg13g2_inv_1 \myring.inv_array[618]/sky_inverter/_0_  (.Y(\myring.inv_in[619] ),
    .A(\myring.inv_in[618] ));
 sg13g2_inv_1 \myring.inv_array[619]/sky_inverter/_0_  (.Y(\myring.inv_in[620] ),
    .A(\myring.inv_in[619] ));
 sg13g2_inv_1 \myring.inv_array[61]/sky_inverter/_0_  (.Y(\myring.inv_in[62] ),
    .A(\myring.inv_in[61] ));
 sg13g2_inv_1 \myring.inv_array[620]/sky_inverter/_0_  (.Y(\myring.inv_in[621] ),
    .A(\myring.inv_in[620] ));
 sg13g2_inv_1 \myring.inv_array[621]/sky_inverter/_0_  (.Y(\myring.inv_in[622] ),
    .A(\myring.inv_in[621] ));
 sg13g2_inv_1 \myring.inv_array[622]/sky_inverter/_0_  (.Y(\myring.inv_in[623] ),
    .A(\myring.inv_in[622] ));
 sg13g2_inv_1 \myring.inv_array[623]/sky_inverter/_0_  (.Y(\myring.inv_in[624] ),
    .A(\myring.inv_in[623] ));
 sg13g2_inv_1 \myring.inv_array[624]/sky_inverter/_0_  (.Y(\myring.inv_in[625] ),
    .A(\myring.inv_in[624] ));
 sg13g2_inv_1 \myring.inv_array[625]/sky_inverter/_0_  (.Y(\myring.inv_in[626] ),
    .A(\myring.inv_in[625] ));
 sg13g2_inv_1 \myring.inv_array[626]/sky_inverter/_0_  (.Y(\myring.inv_in[627] ),
    .A(\myring.inv_in[626] ));
 sg13g2_inv_1 \myring.inv_array[627]/sky_inverter/_0_  (.Y(\myring.inv_in[628] ),
    .A(\myring.inv_in[627] ));
 sg13g2_inv_1 \myring.inv_array[628]/sky_inverter/_0_  (.Y(\myring.inv_in[629] ),
    .A(\myring.inv_in[628] ));
 sg13g2_inv_1 \myring.inv_array[629]/sky_inverter/_0_  (.Y(\myring.inv_in[630] ),
    .A(\myring.inv_in[629] ));
 sg13g2_inv_1 \myring.inv_array[62]/sky_inverter/_0_  (.Y(\myring.inv_in[63] ),
    .A(\myring.inv_in[62] ));
 sg13g2_inv_1 \myring.inv_array[630]/sky_inverter/_0_  (.Y(\myring.inv_in[631] ),
    .A(\myring.inv_in[630] ));
 sg13g2_inv_1 \myring.inv_array[631]/sky_inverter/_0_  (.Y(\myring.inv_in[632] ),
    .A(\myring.inv_in[631] ));
 sg13g2_inv_1 \myring.inv_array[632]/sky_inverter/_0_  (.Y(\myring.inv_in[633] ),
    .A(\myring.inv_in[632] ));
 sg13g2_inv_1 \myring.inv_array[633]/sky_inverter/_0_  (.Y(\myring.inv_in[634] ),
    .A(\myring.inv_in[633] ));
 sg13g2_inv_1 \myring.inv_array[634]/sky_inverter/_0_  (.Y(\myring.inv_in[635] ),
    .A(\myring.inv_in[634] ));
 sg13g2_inv_1 \myring.inv_array[635]/sky_inverter/_0_  (.Y(\myring.inv_in[636] ),
    .A(\myring.inv_in[635] ));
 sg13g2_inv_1 \myring.inv_array[636]/sky_inverter/_0_  (.Y(\myring.inv_in[637] ),
    .A(\myring.inv_in[636] ));
 sg13g2_inv_1 \myring.inv_array[637]/sky_inverter/_0_  (.Y(\myring.inv_in[638] ),
    .A(\myring.inv_in[637] ));
 sg13g2_inv_1 \myring.inv_array[638]/sky_inverter/_0_  (.Y(\myring.inv_in[639] ),
    .A(\myring.inv_in[638] ));
 sg13g2_inv_1 \myring.inv_array[639]/sky_inverter/_0_  (.Y(\myring.inv_in[640] ),
    .A(\myring.inv_in[639] ));
 sg13g2_inv_1 \myring.inv_array[63]/sky_inverter/_0_  (.Y(\myring.inv_in[64] ),
    .A(\myring.inv_in[63] ));
 sg13g2_inv_1 \myring.inv_array[640]/sky_inverter/_0_  (.Y(\myring.inv_in[641] ),
    .A(\myring.inv_in[640] ));
 sg13g2_inv_1 \myring.inv_array[641]/sky_inverter/_0_  (.Y(\myring.inv_in[642] ),
    .A(\myring.inv_in[641] ));
 sg13g2_inv_1 \myring.inv_array[642]/sky_inverter/_0_  (.Y(\myring.inv_in[643] ),
    .A(\myring.inv_in[642] ));
 sg13g2_inv_1 \myring.inv_array[643]/sky_inverter/_0_  (.Y(\myring.inv_in[644] ),
    .A(\myring.inv_in[643] ));
 sg13g2_inv_1 \myring.inv_array[644]/sky_inverter/_0_  (.Y(\myring.inv_in[645] ),
    .A(\myring.inv_in[644] ));
 sg13g2_inv_1 \myring.inv_array[645]/sky_inverter/_0_  (.Y(\myring.inv_in[646] ),
    .A(\myring.inv_in[645] ));
 sg13g2_inv_1 \myring.inv_array[646]/sky_inverter/_0_  (.Y(\myring.inv_in[647] ),
    .A(\myring.inv_in[646] ));
 sg13g2_inv_1 \myring.inv_array[647]/sky_inverter/_0_  (.Y(\myring.inv_in[648] ),
    .A(\myring.inv_in[647] ));
 sg13g2_inv_1 \myring.inv_array[648]/sky_inverter/_0_  (.Y(\myring.inv_in[649] ),
    .A(\myring.inv_in[648] ));
 sg13g2_inv_1 \myring.inv_array[649]/sky_inverter/_0_  (.Y(\myring.inv_in[650] ),
    .A(\myring.inv_in[649] ));
 sg13g2_inv_1 \myring.inv_array[64]/sky_inverter/_0_  (.Y(\myring.inv_in[65] ),
    .A(\myring.inv_in[64] ));
 sg13g2_inv_1 \myring.inv_array[650]/sky_inverter/_0_  (.Y(\myring.inv_in[651] ),
    .A(\myring.inv_in[650] ));
 sg13g2_inv_1 \myring.inv_array[651]/sky_inverter/_0_  (.Y(\myring.inv_in[652] ),
    .A(\myring.inv_in[651] ));
 sg13g2_inv_1 \myring.inv_array[652]/sky_inverter/_0_  (.Y(\myring.inv_in[653] ),
    .A(\myring.inv_in[652] ));
 sg13g2_inv_1 \myring.inv_array[653]/sky_inverter/_0_  (.Y(\myring.inv_in[654] ),
    .A(\myring.inv_in[653] ));
 sg13g2_inv_1 \myring.inv_array[654]/sky_inverter/_0_  (.Y(\myring.inv_in[655] ),
    .A(\myring.inv_in[654] ));
 sg13g2_inv_1 \myring.inv_array[655]/sky_inverter/_0_  (.Y(\myring.inv_in[656] ),
    .A(\myring.inv_in[655] ));
 sg13g2_inv_1 \myring.inv_array[656]/sky_inverter/_0_  (.Y(\myring.inv_in[657] ),
    .A(\myring.inv_in[656] ));
 sg13g2_inv_1 \myring.inv_array[657]/sky_inverter/_0_  (.Y(\myring.inv_in[658] ),
    .A(\myring.inv_in[657] ));
 sg13g2_inv_1 \myring.inv_array[658]/sky_inverter/_0_  (.Y(\myring.inv_in[659] ),
    .A(\myring.inv_in[658] ));
 sg13g2_inv_1 \myring.inv_array[659]/sky_inverter/_0_  (.Y(\myring.inv_in[660] ),
    .A(\myring.inv_in[659] ));
 sg13g2_inv_1 \myring.inv_array[65]/sky_inverter/_0_  (.Y(\myring.inv_in[66] ),
    .A(\myring.inv_in[65] ));
 sg13g2_inv_1 \myring.inv_array[660]/sky_inverter/_0_  (.Y(\myring.inv_in[661] ),
    .A(\myring.inv_in[660] ));
 sg13g2_inv_1 \myring.inv_array[661]/sky_inverter/_0_  (.Y(\myring.inv_in[662] ),
    .A(\myring.inv_in[661] ));
 sg13g2_inv_1 \myring.inv_array[662]/sky_inverter/_0_  (.Y(\myring.inv_in[663] ),
    .A(\myring.inv_in[662] ));
 sg13g2_inv_1 \myring.inv_array[663]/sky_inverter/_0_  (.Y(\myring.inv_in[664] ),
    .A(\myring.inv_in[663] ));
 sg13g2_inv_1 \myring.inv_array[664]/sky_inverter/_0_  (.Y(\myring.inv_in[665] ),
    .A(\myring.inv_in[664] ));
 sg13g2_inv_1 \myring.inv_array[665]/sky_inverter/_0_  (.Y(\myring.inv_in[666] ),
    .A(\myring.inv_in[665] ));
 sg13g2_inv_1 \myring.inv_array[666]/sky_inverter/_0_  (.Y(\myring.inv_in[667] ),
    .A(\myring.inv_in[666] ));
 sg13g2_inv_1 \myring.inv_array[667]/sky_inverter/_0_  (.Y(\myring.inv_in[668] ),
    .A(\myring.inv_in[667] ));
 sg13g2_inv_1 \myring.inv_array[668]/sky_inverter/_0_  (.Y(\myring.inv_in[669] ),
    .A(\myring.inv_in[668] ));
 sg13g2_inv_1 \myring.inv_array[669]/sky_inverter/_0_  (.Y(\myring.inv_in[670] ),
    .A(\myring.inv_in[669] ));
 sg13g2_inv_1 \myring.inv_array[66]/sky_inverter/_0_  (.Y(\myring.inv_in[67] ),
    .A(\myring.inv_in[66] ));
 sg13g2_inv_1 \myring.inv_array[670]/sky_inverter/_0_  (.Y(\myring.inv_in[671] ),
    .A(\myring.inv_in[670] ));
 sg13g2_inv_1 \myring.inv_array[671]/sky_inverter/_0_  (.Y(\myring.inv_in[672] ),
    .A(\myring.inv_in[671] ));
 sg13g2_inv_1 \myring.inv_array[672]/sky_inverter/_0_  (.Y(\myring.inv_in[673] ),
    .A(\myring.inv_in[672] ));
 sg13g2_inv_1 \myring.inv_array[673]/sky_inverter/_0_  (.Y(\myring.inv_in[674] ),
    .A(\myring.inv_in[673] ));
 sg13g2_inv_1 \myring.inv_array[674]/sky_inverter/_0_  (.Y(\myring.inv_in[675] ),
    .A(\myring.inv_in[674] ));
 sg13g2_inv_1 \myring.inv_array[675]/sky_inverter/_0_  (.Y(\myring.inv_in[676] ),
    .A(\myring.inv_in[675] ));
 sg13g2_inv_1 \myring.inv_array[676]/sky_inverter/_0_  (.Y(\myring.inv_in[677] ),
    .A(\myring.inv_in[676] ));
 sg13g2_inv_1 \myring.inv_array[677]/sky_inverter/_0_  (.Y(\myring.inv_in[678] ),
    .A(\myring.inv_in[677] ));
 sg13g2_inv_1 \myring.inv_array[678]/sky_inverter/_0_  (.Y(\myring.inv_in[679] ),
    .A(\myring.inv_in[678] ));
 sg13g2_inv_1 \myring.inv_array[679]/sky_inverter/_0_  (.Y(\myring.inv_in[680] ),
    .A(\myring.inv_in[679] ));
 sg13g2_inv_1 \myring.inv_array[67]/sky_inverter/_0_  (.Y(\myring.inv_in[68] ),
    .A(\myring.inv_in[67] ));
 sg13g2_inv_1 \myring.inv_array[680]/sky_inverter/_0_  (.Y(\myring.inv_in[681] ),
    .A(\myring.inv_in[680] ));
 sg13g2_inv_1 \myring.inv_array[681]/sky_inverter/_0_  (.Y(\myring.inv_in[682] ),
    .A(\myring.inv_in[681] ));
 sg13g2_inv_1 \myring.inv_array[682]/sky_inverter/_0_  (.Y(\myring.inv_in[683] ),
    .A(\myring.inv_in[682] ));
 sg13g2_inv_1 \myring.inv_array[683]/sky_inverter/_0_  (.Y(\myring.inv_in[684] ),
    .A(\myring.inv_in[683] ));
 sg13g2_inv_1 \myring.inv_array[684]/sky_inverter/_0_  (.Y(\myring.inv_in[685] ),
    .A(\myring.inv_in[684] ));
 sg13g2_inv_1 \myring.inv_array[685]/sky_inverter/_0_  (.Y(\myring.inv_in[686] ),
    .A(\myring.inv_in[685] ));
 sg13g2_inv_1 \myring.inv_array[686]/sky_inverter/_0_  (.Y(\myring.inv_in[687] ),
    .A(\myring.inv_in[686] ));
 sg13g2_inv_1 \myring.inv_array[687]/sky_inverter/_0_  (.Y(\myring.inv_in[688] ),
    .A(\myring.inv_in[687] ));
 sg13g2_inv_1 \myring.inv_array[688]/sky_inverter/_0_  (.Y(\myring.inv_in[689] ),
    .A(\myring.inv_in[688] ));
 sg13g2_inv_1 \myring.inv_array[689]/sky_inverter/_0_  (.Y(\myring.inv_in[690] ),
    .A(\myring.inv_in[689] ));
 sg13g2_inv_1 \myring.inv_array[68]/sky_inverter/_0_  (.Y(\myring.inv_in[69] ),
    .A(\myring.inv_in[68] ));
 sg13g2_inv_1 \myring.inv_array[690]/sky_inverter/_0_  (.Y(\myring.inv_in[691] ),
    .A(\myring.inv_in[690] ));
 sg13g2_inv_1 \myring.inv_array[691]/sky_inverter/_0_  (.Y(\myring.inv_in[692] ),
    .A(\myring.inv_in[691] ));
 sg13g2_inv_1 \myring.inv_array[692]/sky_inverter/_0_  (.Y(\myring.inv_in[693] ),
    .A(\myring.inv_in[692] ));
 sg13g2_inv_1 \myring.inv_array[693]/sky_inverter/_0_  (.Y(\myring.inv_in[694] ),
    .A(\myring.inv_in[693] ));
 sg13g2_inv_1 \myring.inv_array[694]/sky_inverter/_0_  (.Y(\myring.inv_in[695] ),
    .A(\myring.inv_in[694] ));
 sg13g2_inv_1 \myring.inv_array[695]/sky_inverter/_0_  (.Y(\myring.inv_in[696] ),
    .A(\myring.inv_in[695] ));
 sg13g2_inv_1 \myring.inv_array[696]/sky_inverter/_0_  (.Y(\myring.inv_in[697] ),
    .A(\myring.inv_in[696] ));
 sg13g2_inv_1 \myring.inv_array[697]/sky_inverter/_0_  (.Y(\myring.inv_in[698] ),
    .A(\myring.inv_in[697] ));
 sg13g2_inv_1 \myring.inv_array[698]/sky_inverter/_0_  (.Y(\myring.inv_in[699] ),
    .A(\myring.inv_in[698] ));
 sg13g2_inv_1 \myring.inv_array[699]/sky_inverter/_0_  (.Y(\myring.inv_in[700] ),
    .A(\myring.inv_in[699] ));
 sg13g2_inv_1 \myring.inv_array[69]/sky_inverter/_0_  (.Y(\myring.inv_in[70] ),
    .A(\myring.inv_in[69] ));
 sg13g2_inv_1 \myring.inv_array[6]/sky_inverter/_0_  (.Y(\myring.inv_in[7] ),
    .A(\myring.inv_in[6] ));
 sg13g2_inv_1 \myring.inv_array[700]/sky_inverter/_0_  (.Y(\myring.inv_in[701] ),
    .A(\myring.inv_in[700] ));
 sg13g2_inv_1 \myring.inv_array[701]/sky_inverter/_0_  (.Y(\myring.inv_in[702] ),
    .A(\myring.inv_in[701] ));
 sg13g2_inv_1 \myring.inv_array[702]/sky_inverter/_0_  (.Y(\myring.inv_in[703] ),
    .A(\myring.inv_in[702] ));
 sg13g2_inv_1 \myring.inv_array[703]/sky_inverter/_0_  (.Y(\myring.inv_in[704] ),
    .A(\myring.inv_in[703] ));
 sg13g2_inv_1 \myring.inv_array[704]/sky_inverter/_0_  (.Y(\myring.inv_in[705] ),
    .A(\myring.inv_in[704] ));
 sg13g2_inv_1 \myring.inv_array[705]/sky_inverter/_0_  (.Y(\myring.inv_in[706] ),
    .A(\myring.inv_in[705] ));
 sg13g2_inv_1 \myring.inv_array[706]/sky_inverter/_0_  (.Y(\myring.inv_in[707] ),
    .A(\myring.inv_in[706] ));
 sg13g2_inv_1 \myring.inv_array[707]/sky_inverter/_0_  (.Y(\myring.inv_in[708] ),
    .A(\myring.inv_in[707] ));
 sg13g2_inv_1 \myring.inv_array[708]/sky_inverter/_0_  (.Y(\myring.inv_in[709] ),
    .A(\myring.inv_in[708] ));
 sg13g2_inv_1 \myring.inv_array[709]/sky_inverter/_0_  (.Y(\myring.inv_in[710] ),
    .A(\myring.inv_in[709] ));
 sg13g2_inv_1 \myring.inv_array[70]/sky_inverter/_0_  (.Y(\myring.inv_in[71] ),
    .A(\myring.inv_in[70] ));
 sg13g2_inv_1 \myring.inv_array[710]/sky_inverter/_0_  (.Y(\myring.inv_in[711] ),
    .A(\myring.inv_in[710] ));
 sg13g2_inv_1 \myring.inv_array[711]/sky_inverter/_0_  (.Y(\myring.inv_in[712] ),
    .A(\myring.inv_in[711] ));
 sg13g2_inv_1 \myring.inv_array[712]/sky_inverter/_0_  (.Y(\myring.inv_in[713] ),
    .A(\myring.inv_in[712] ));
 sg13g2_inv_1 \myring.inv_array[713]/sky_inverter/_0_  (.Y(\myring.inv_in[714] ),
    .A(\myring.inv_in[713] ));
 sg13g2_inv_1 \myring.inv_array[714]/sky_inverter/_0_  (.Y(\myring.inv_in[715] ),
    .A(\myring.inv_in[714] ));
 sg13g2_inv_1 \myring.inv_array[715]/sky_inverter/_0_  (.Y(\myring.inv_in[716] ),
    .A(\myring.inv_in[715] ));
 sg13g2_inv_1 \myring.inv_array[716]/sky_inverter/_0_  (.Y(\myring.inv_in[717] ),
    .A(\myring.inv_in[716] ));
 sg13g2_inv_1 \myring.inv_array[717]/sky_inverter/_0_  (.Y(\myring.inv_in[718] ),
    .A(\myring.inv_in[717] ));
 sg13g2_inv_1 \myring.inv_array[718]/sky_inverter/_0_  (.Y(\myring.inv_in[719] ),
    .A(\myring.inv_in[718] ));
 sg13g2_inv_1 \myring.inv_array[719]/sky_inverter/_0_  (.Y(\myring.inv_in[720] ),
    .A(\myring.inv_in[719] ));
 sg13g2_inv_1 \myring.inv_array[71]/sky_inverter/_0_  (.Y(\myring.inv_in[72] ),
    .A(\myring.inv_in[71] ));
 sg13g2_inv_1 \myring.inv_array[720]/sky_inverter/_0_  (.Y(\myring.inv_in[721] ),
    .A(\myring.inv_in[720] ));
 sg13g2_inv_1 \myring.inv_array[721]/sky_inverter/_0_  (.Y(\myring.inv_in[722] ),
    .A(\myring.inv_in[721] ));
 sg13g2_inv_1 \myring.inv_array[722]/sky_inverter/_0_  (.Y(\myring.inv_in[723] ),
    .A(\myring.inv_in[722] ));
 sg13g2_inv_1 \myring.inv_array[723]/sky_inverter/_0_  (.Y(\myring.inv_in[724] ),
    .A(\myring.inv_in[723] ));
 sg13g2_inv_1 \myring.inv_array[724]/sky_inverter/_0_  (.Y(\myring.inv_in[725] ),
    .A(\myring.inv_in[724] ));
 sg13g2_inv_1 \myring.inv_array[725]/sky_inverter/_0_  (.Y(\myring.inv_in[726] ),
    .A(\myring.inv_in[725] ));
 sg13g2_inv_1 \myring.inv_array[726]/sky_inverter/_0_  (.Y(\myring.inv_in[727] ),
    .A(\myring.inv_in[726] ));
 sg13g2_inv_1 \myring.inv_array[727]/sky_inverter/_0_  (.Y(\myring.inv_in[728] ),
    .A(\myring.inv_in[727] ));
 sg13g2_inv_1 \myring.inv_array[728]/sky_inverter/_0_  (.Y(\myring.inv_in[729] ),
    .A(\myring.inv_in[728] ));
 sg13g2_inv_1 \myring.inv_array[729]/sky_inverter/_0_  (.Y(\myring.inv_in[730] ),
    .A(\myring.inv_in[729] ));
 sg13g2_inv_1 \myring.inv_array[72]/sky_inverter/_0_  (.Y(\myring.inv_in[73] ),
    .A(\myring.inv_in[72] ));
 sg13g2_inv_1 \myring.inv_array[730]/sky_inverter/_0_  (.Y(\myring.inv_in[731] ),
    .A(\myring.inv_in[730] ));
 sg13g2_inv_1 \myring.inv_array[731]/sky_inverter/_0_  (.Y(\myring.inv_in[732] ),
    .A(\myring.inv_in[731] ));
 sg13g2_inv_1 \myring.inv_array[732]/sky_inverter/_0_  (.Y(\myring.inv_in[733] ),
    .A(\myring.inv_in[732] ));
 sg13g2_inv_1 \myring.inv_array[733]/sky_inverter/_0_  (.Y(\myring.inv_in[734] ),
    .A(\myring.inv_in[733] ));
 sg13g2_inv_1 \myring.inv_array[734]/sky_inverter/_0_  (.Y(\myring.inv_in[735] ),
    .A(\myring.inv_in[734] ));
 sg13g2_inv_1 \myring.inv_array[735]/sky_inverter/_0_  (.Y(\myring.inv_in[736] ),
    .A(\myring.inv_in[735] ));
 sg13g2_inv_1 \myring.inv_array[736]/sky_inverter/_0_  (.Y(\myring.inv_in[737] ),
    .A(\myring.inv_in[736] ));
 sg13g2_inv_1 \myring.inv_array[737]/sky_inverter/_0_  (.Y(\myring.inv_in[738] ),
    .A(\myring.inv_in[737] ));
 sg13g2_inv_1 \myring.inv_array[738]/sky_inverter/_0_  (.Y(\myring.inv_in[739] ),
    .A(\myring.inv_in[738] ));
 sg13g2_inv_1 \myring.inv_array[739]/sky_inverter/_0_  (.Y(\myring.inv_in[740] ),
    .A(\myring.inv_in[739] ));
 sg13g2_inv_1 \myring.inv_array[73]/sky_inverter/_0_  (.Y(\myring.inv_in[74] ),
    .A(\myring.inv_in[73] ));
 sg13g2_inv_1 \myring.inv_array[740]/sky_inverter/_0_  (.Y(\myring.inv_in[741] ),
    .A(\myring.inv_in[740] ));
 sg13g2_inv_1 \myring.inv_array[741]/sky_inverter/_0_  (.Y(\myring.inv_in[742] ),
    .A(\myring.inv_in[741] ));
 sg13g2_inv_1 \myring.inv_array[742]/sky_inverter/_0_  (.Y(\myring.inv_in[743] ),
    .A(\myring.inv_in[742] ));
 sg13g2_inv_1 \myring.inv_array[743]/sky_inverter/_0_  (.Y(\myring.inv_in[744] ),
    .A(\myring.inv_in[743] ));
 sg13g2_inv_1 \myring.inv_array[744]/sky_inverter/_0_  (.Y(\myring.inv_in[745] ),
    .A(\myring.inv_in[744] ));
 sg13g2_inv_1 \myring.inv_array[745]/sky_inverter/_0_  (.Y(\myring.inv_in[746] ),
    .A(\myring.inv_in[745] ));
 sg13g2_inv_1 \myring.inv_array[746]/sky_inverter/_0_  (.Y(\myring.inv_in[747] ),
    .A(\myring.inv_in[746] ));
 sg13g2_inv_1 \myring.inv_array[747]/sky_inverter/_0_  (.Y(\myring.inv_in[748] ),
    .A(\myring.inv_in[747] ));
 sg13g2_inv_1 \myring.inv_array[748]/sky_inverter/_0_  (.Y(\myring.inv_in[749] ),
    .A(\myring.inv_in[748] ));
 sg13g2_inv_1 \myring.inv_array[749]/sky_inverter/_0_  (.Y(\myring.inv_in[750] ),
    .A(\myring.inv_in[749] ));
 sg13g2_inv_1 \myring.inv_array[74]/sky_inverter/_0_  (.Y(\myring.inv_in[75] ),
    .A(\myring.inv_in[74] ));
 sg13g2_inv_1 \myring.inv_array[750]/sky_inverter/_0_  (.Y(\myring.inv_in[751] ),
    .A(\myring.inv_in[750] ));
 sg13g2_inv_1 \myring.inv_array[751]/sky_inverter/_0_  (.Y(\myring.inv_in[752] ),
    .A(\myring.inv_in[751] ));
 sg13g2_inv_1 \myring.inv_array[752]/sky_inverter/_0_  (.Y(\myring.inv_in[753] ),
    .A(\myring.inv_in[752] ));
 sg13g2_inv_1 \myring.inv_array[753]/sky_inverter/_0_  (.Y(\myring.inv_in[754] ),
    .A(\myring.inv_in[753] ));
 sg13g2_inv_1 \myring.inv_array[754]/sky_inverter/_0_  (.Y(\myring.inv_in[755] ),
    .A(\myring.inv_in[754] ));
 sg13g2_inv_1 \myring.inv_array[755]/sky_inverter/_0_  (.Y(\myring.inv_in[756] ),
    .A(\myring.inv_in[755] ));
 sg13g2_inv_1 \myring.inv_array[756]/sky_inverter/_0_  (.Y(\myring.inv_in[757] ),
    .A(\myring.inv_in[756] ));
 sg13g2_inv_1 \myring.inv_array[757]/sky_inverter/_0_  (.Y(\myring.inv_in[758] ),
    .A(\myring.inv_in[757] ));
 sg13g2_inv_1 \myring.inv_array[758]/sky_inverter/_0_  (.Y(\myring.inv_in[759] ),
    .A(\myring.inv_in[758] ));
 sg13g2_inv_1 \myring.inv_array[759]/sky_inverter/_0_  (.Y(\myring.inv_in[760] ),
    .A(\myring.inv_in[759] ));
 sg13g2_inv_1 \myring.inv_array[75]/sky_inverter/_0_  (.Y(\myring.inv_in[76] ),
    .A(\myring.inv_in[75] ));
 sg13g2_inv_1 \myring.inv_array[760]/sky_inverter/_0_  (.Y(\myring.inv_in[761] ),
    .A(\myring.inv_in[760] ));
 sg13g2_inv_1 \myring.inv_array[761]/sky_inverter/_0_  (.Y(\myring.inv_in[762] ),
    .A(\myring.inv_in[761] ));
 sg13g2_inv_1 \myring.inv_array[762]/sky_inverter/_0_  (.Y(\myring.inv_in[763] ),
    .A(\myring.inv_in[762] ));
 sg13g2_inv_1 \myring.inv_array[763]/sky_inverter/_0_  (.Y(\myring.inv_in[764] ),
    .A(\myring.inv_in[763] ));
 sg13g2_inv_1 \myring.inv_array[764]/sky_inverter/_0_  (.Y(\myring.inv_in[765] ),
    .A(\myring.inv_in[764] ));
 sg13g2_inv_1 \myring.inv_array[765]/sky_inverter/_0_  (.Y(\myring.inv_in[766] ),
    .A(\myring.inv_in[765] ));
 sg13g2_inv_1 \myring.inv_array[766]/sky_inverter/_0_  (.Y(\myring.inv_in[767] ),
    .A(\myring.inv_in[766] ));
 sg13g2_inv_1 \myring.inv_array[767]/sky_inverter/_0_  (.Y(\myring.inv_in[768] ),
    .A(\myring.inv_in[767] ));
 sg13g2_inv_1 \myring.inv_array[768]/sky_inverter/_0_  (.Y(\myring.inv_in[769] ),
    .A(\myring.inv_in[768] ));
 sg13g2_inv_1 \myring.inv_array[769]/sky_inverter/_0_  (.Y(\myring.inv_in[770] ),
    .A(\myring.inv_in[769] ));
 sg13g2_inv_1 \myring.inv_array[76]/sky_inverter/_0_  (.Y(\myring.inv_in[77] ),
    .A(\myring.inv_in[76] ));
 sg13g2_inv_1 \myring.inv_array[770]/sky_inverter/_0_  (.Y(\myring.inv_in[771] ),
    .A(\myring.inv_in[770] ));
 sg13g2_inv_1 \myring.inv_array[771]/sky_inverter/_0_  (.Y(\myring.inv_in[772] ),
    .A(\myring.inv_in[771] ));
 sg13g2_inv_1 \myring.inv_array[772]/sky_inverter/_0_  (.Y(\myring.inv_in[773] ),
    .A(\myring.inv_in[772] ));
 sg13g2_inv_1 \myring.inv_array[773]/sky_inverter/_0_  (.Y(\myring.inv_in[774] ),
    .A(\myring.inv_in[773] ));
 sg13g2_inv_1 \myring.inv_array[774]/sky_inverter/_0_  (.Y(\myring.inv_in[775] ),
    .A(\myring.inv_in[774] ));
 sg13g2_inv_1 \myring.inv_array[775]/sky_inverter/_0_  (.Y(\myring.inv_in[776] ),
    .A(\myring.inv_in[775] ));
 sg13g2_inv_1 \myring.inv_array[776]/sky_inverter/_0_  (.Y(\myring.inv_in[777] ),
    .A(\myring.inv_in[776] ));
 sg13g2_inv_1 \myring.inv_array[777]/sky_inverter/_0_  (.Y(\myring.inv_in[778] ),
    .A(\myring.inv_in[777] ));
 sg13g2_inv_1 \myring.inv_array[778]/sky_inverter/_0_  (.Y(\myring.inv_in[779] ),
    .A(\myring.inv_in[778] ));
 sg13g2_inv_1 \myring.inv_array[779]/sky_inverter/_0_  (.Y(\myring.inv_in[780] ),
    .A(\myring.inv_in[779] ));
 sg13g2_inv_1 \myring.inv_array[77]/sky_inverter/_0_  (.Y(\myring.inv_in[78] ),
    .A(\myring.inv_in[77] ));
 sg13g2_inv_1 \myring.inv_array[780]/sky_inverter/_0_  (.Y(\myring.inv_in[781] ),
    .A(\myring.inv_in[780] ));
 sg13g2_inv_1 \myring.inv_array[781]/sky_inverter/_0_  (.Y(\myring.inv_in[782] ),
    .A(\myring.inv_in[781] ));
 sg13g2_inv_1 \myring.inv_array[782]/sky_inverter/_0_  (.Y(\myring.inv_in[783] ),
    .A(\myring.inv_in[782] ));
 sg13g2_inv_1 \myring.inv_array[783]/sky_inverter/_0_  (.Y(\myring.inv_in[784] ),
    .A(\myring.inv_in[783] ));
 sg13g2_inv_1 \myring.inv_array[784]/sky_inverter/_0_  (.Y(\myring.inv_in[785] ),
    .A(\myring.inv_in[784] ));
 sg13g2_inv_1 \myring.inv_array[785]/sky_inverter/_0_  (.Y(\myring.inv_in[786] ),
    .A(\myring.inv_in[785] ));
 sg13g2_inv_1 \myring.inv_array[786]/sky_inverter/_0_  (.Y(\myring.inv_in[787] ),
    .A(\myring.inv_in[786] ));
 sg13g2_inv_1 \myring.inv_array[787]/sky_inverter/_0_  (.Y(\myring.inv_in[788] ),
    .A(\myring.inv_in[787] ));
 sg13g2_inv_1 \myring.inv_array[788]/sky_inverter/_0_  (.Y(\myring.inv_in[789] ),
    .A(\myring.inv_in[788] ));
 sg13g2_inv_1 \myring.inv_array[789]/sky_inverter/_0_  (.Y(\myring.inv_in[790] ),
    .A(\myring.inv_in[789] ));
 sg13g2_inv_1 \myring.inv_array[78]/sky_inverter/_0_  (.Y(\myring.inv_in[79] ),
    .A(\myring.inv_in[78] ));
 sg13g2_inv_1 \myring.inv_array[790]/sky_inverter/_0_  (.Y(\myring.inv_in[791] ),
    .A(\myring.inv_in[790] ));
 sg13g2_inv_1 \myring.inv_array[791]/sky_inverter/_0_  (.Y(\myring.inv_in[792] ),
    .A(\myring.inv_in[791] ));
 sg13g2_inv_1 \myring.inv_array[792]/sky_inverter/_0_  (.Y(\myring.inv_in[793] ),
    .A(\myring.inv_in[792] ));
 sg13g2_inv_1 \myring.inv_array[793]/sky_inverter/_0_  (.Y(\myring.inv_in[794] ),
    .A(\myring.inv_in[793] ));
 sg13g2_inv_1 \myring.inv_array[794]/sky_inverter/_0_  (.Y(\myring.inv_in[795] ),
    .A(\myring.inv_in[794] ));
 sg13g2_inv_1 \myring.inv_array[795]/sky_inverter/_0_  (.Y(\myring.inv_in[796] ),
    .A(\myring.inv_in[795] ));
 sg13g2_inv_1 \myring.inv_array[796]/sky_inverter/_0_  (.Y(\myring.inv_in[797] ),
    .A(\myring.inv_in[796] ));
 sg13g2_inv_1 \myring.inv_array[797]/sky_inverter/_0_  (.Y(\myring.inv_in[798] ),
    .A(\myring.inv_in[797] ));
 sg13g2_inv_1 \myring.inv_array[798]/sky_inverter/_0_  (.Y(\myring.inv_in[799] ),
    .A(\myring.inv_in[798] ));
 sg13g2_inv_1 \myring.inv_array[799]/sky_inverter/_0_  (.Y(\myring.inv_in[800] ),
    .A(\myring.inv_in[799] ));
 sg13g2_inv_1 \myring.inv_array[79]/sky_inverter/_0_  (.Y(\myring.inv_in[80] ),
    .A(\myring.inv_in[79] ));
 sg13g2_inv_1 \myring.inv_array[7]/sky_inverter/_0_  (.Y(\myring.inv_in[8] ),
    .A(\myring.inv_in[7] ));
 sg13g2_inv_1 \myring.inv_array[800]/sky_inverter/_0_  (.Y(\myring.inv_in[801] ),
    .A(\myring.inv_in[800] ));
 sg13g2_inv_1 \myring.inv_array[801]/sky_inverter/_0_  (.Y(\myring.inv_in[802] ),
    .A(\myring.inv_in[801] ));
 sg13g2_inv_1 \myring.inv_array[802]/sky_inverter/_0_  (.Y(\myring.inv_in[803] ),
    .A(\myring.inv_in[802] ));
 sg13g2_inv_1 \myring.inv_array[803]/sky_inverter/_0_  (.Y(\myring.inv_in[804] ),
    .A(\myring.inv_in[803] ));
 sg13g2_inv_1 \myring.inv_array[804]/sky_inverter/_0_  (.Y(\myring.inv_in[805] ),
    .A(\myring.inv_in[804] ));
 sg13g2_inv_1 \myring.inv_array[805]/sky_inverter/_0_  (.Y(\myring.inv_in[806] ),
    .A(\myring.inv_in[805] ));
 sg13g2_inv_1 \myring.inv_array[806]/sky_inverter/_0_  (.Y(\myring.inv_in[807] ),
    .A(\myring.inv_in[806] ));
 sg13g2_inv_1 \myring.inv_array[807]/sky_inverter/_0_  (.Y(\myring.inv_in[808] ),
    .A(\myring.inv_in[807] ));
 sg13g2_inv_1 \myring.inv_array[808]/sky_inverter/_0_  (.Y(\myring.inv_in[809] ),
    .A(\myring.inv_in[808] ));
 sg13g2_inv_1 \myring.inv_array[809]/sky_inverter/_0_  (.Y(\myring.inv_in[810] ),
    .A(\myring.inv_in[809] ));
 sg13g2_inv_1 \myring.inv_array[80]/sky_inverter/_0_  (.Y(\myring.inv_in[81] ),
    .A(\myring.inv_in[80] ));
 sg13g2_inv_1 \myring.inv_array[810]/sky_inverter/_0_  (.Y(\myring.inv_in[811] ),
    .A(\myring.inv_in[810] ));
 sg13g2_inv_1 \myring.inv_array[811]/sky_inverter/_0_  (.Y(\myring.inv_in[812] ),
    .A(\myring.inv_in[811] ));
 sg13g2_inv_1 \myring.inv_array[812]/sky_inverter/_0_  (.Y(\myring.inv_in[813] ),
    .A(\myring.inv_in[812] ));
 sg13g2_inv_1 \myring.inv_array[813]/sky_inverter/_0_  (.Y(\myring.inv_in[814] ),
    .A(\myring.inv_in[813] ));
 sg13g2_inv_1 \myring.inv_array[814]/sky_inverter/_0_  (.Y(\myring.inv_in[815] ),
    .A(\myring.inv_in[814] ));
 sg13g2_inv_1 \myring.inv_array[815]/sky_inverter/_0_  (.Y(\myring.inv_in[816] ),
    .A(\myring.inv_in[815] ));
 sg13g2_inv_1 \myring.inv_array[816]/sky_inverter/_0_  (.Y(\myring.inv_in[817] ),
    .A(\myring.inv_in[816] ));
 sg13g2_inv_1 \myring.inv_array[817]/sky_inverter/_0_  (.Y(\myring.inv_in[818] ),
    .A(\myring.inv_in[817] ));
 sg13g2_inv_1 \myring.inv_array[818]/sky_inverter/_0_  (.Y(\myring.inv_in[819] ),
    .A(\myring.inv_in[818] ));
 sg13g2_inv_1 \myring.inv_array[819]/sky_inverter/_0_  (.Y(\myring.inv_in[820] ),
    .A(\myring.inv_in[819] ));
 sg13g2_inv_1 \myring.inv_array[81]/sky_inverter/_0_  (.Y(\myring.inv_in[82] ),
    .A(\myring.inv_in[81] ));
 sg13g2_inv_1 \myring.inv_array[820]/sky_inverter/_0_  (.Y(\myring.inv_in[821] ),
    .A(\myring.inv_in[820] ));
 sg13g2_inv_1 \myring.inv_array[821]/sky_inverter/_0_  (.Y(\myring.inv_in[822] ),
    .A(\myring.inv_in[821] ));
 sg13g2_inv_1 \myring.inv_array[822]/sky_inverter/_0_  (.Y(\myring.inv_in[823] ),
    .A(\myring.inv_in[822] ));
 sg13g2_inv_1 \myring.inv_array[823]/sky_inverter/_0_  (.Y(\myring.inv_in[824] ),
    .A(\myring.inv_in[823] ));
 sg13g2_inv_1 \myring.inv_array[824]/sky_inverter/_0_  (.Y(\myring.inv_in[825] ),
    .A(\myring.inv_in[824] ));
 sg13g2_inv_1 \myring.inv_array[825]/sky_inverter/_0_  (.Y(\myring.inv_in[826] ),
    .A(\myring.inv_in[825] ));
 sg13g2_inv_1 \myring.inv_array[826]/sky_inverter/_0_  (.Y(\myring.inv_in[827] ),
    .A(\myring.inv_in[826] ));
 sg13g2_inv_1 \myring.inv_array[827]/sky_inverter/_0_  (.Y(\myring.inv_in[828] ),
    .A(\myring.inv_in[827] ));
 sg13g2_inv_1 \myring.inv_array[828]/sky_inverter/_0_  (.Y(\myring.inv_in[829] ),
    .A(\myring.inv_in[828] ));
 sg13g2_inv_1 \myring.inv_array[829]/sky_inverter/_0_  (.Y(\myring.inv_in[830] ),
    .A(\myring.inv_in[829] ));
 sg13g2_inv_1 \myring.inv_array[82]/sky_inverter/_0_  (.Y(\myring.inv_in[83] ),
    .A(\myring.inv_in[82] ));
 sg13g2_inv_1 \myring.inv_array[830]/sky_inverter/_0_  (.Y(\myring.inv_in[831] ),
    .A(\myring.inv_in[830] ));
 sg13g2_inv_1 \myring.inv_array[831]/sky_inverter/_0_  (.Y(\myring.inv_in[832] ),
    .A(\myring.inv_in[831] ));
 sg13g2_inv_1 \myring.inv_array[832]/sky_inverter/_0_  (.Y(\myring.inv_in[833] ),
    .A(\myring.inv_in[832] ));
 sg13g2_inv_1 \myring.inv_array[833]/sky_inverter/_0_  (.Y(\myring.inv_in[834] ),
    .A(\myring.inv_in[833] ));
 sg13g2_inv_1 \myring.inv_array[834]/sky_inverter/_0_  (.Y(\myring.inv_in[835] ),
    .A(\myring.inv_in[834] ));
 sg13g2_inv_1 \myring.inv_array[835]/sky_inverter/_0_  (.Y(\myring.inv_in[836] ),
    .A(\myring.inv_in[835] ));
 sg13g2_inv_1 \myring.inv_array[836]/sky_inverter/_0_  (.Y(\myring.inv_in[837] ),
    .A(\myring.inv_in[836] ));
 sg13g2_inv_1 \myring.inv_array[837]/sky_inverter/_0_  (.Y(\myring.inv_in[838] ),
    .A(\myring.inv_in[837] ));
 sg13g2_inv_1 \myring.inv_array[838]/sky_inverter/_0_  (.Y(\myring.inv_in[839] ),
    .A(\myring.inv_in[838] ));
 sg13g2_inv_1 \myring.inv_array[839]/sky_inverter/_0_  (.Y(\myring.inv_in[840] ),
    .A(\myring.inv_in[839] ));
 sg13g2_inv_1 \myring.inv_array[83]/sky_inverter/_0_  (.Y(\myring.inv_in[84] ),
    .A(\myring.inv_in[83] ));
 sg13g2_inv_1 \myring.inv_array[840]/sky_inverter/_0_  (.Y(\myring.inv_in[841] ),
    .A(\myring.inv_in[840] ));
 sg13g2_inv_1 \myring.inv_array[841]/sky_inverter/_0_  (.Y(\myring.inv_in[842] ),
    .A(\myring.inv_in[841] ));
 sg13g2_inv_1 \myring.inv_array[842]/sky_inverter/_0_  (.Y(\myring.inv_in[843] ),
    .A(\myring.inv_in[842] ));
 sg13g2_inv_1 \myring.inv_array[843]/sky_inverter/_0_  (.Y(\myring.inv_in[844] ),
    .A(\myring.inv_in[843] ));
 sg13g2_inv_1 \myring.inv_array[844]/sky_inverter/_0_  (.Y(\myring.inv_in[845] ),
    .A(\myring.inv_in[844] ));
 sg13g2_inv_1 \myring.inv_array[845]/sky_inverter/_0_  (.Y(\myring.inv_in[846] ),
    .A(\myring.inv_in[845] ));
 sg13g2_inv_1 \myring.inv_array[846]/sky_inverter/_0_  (.Y(\myring.inv_in[847] ),
    .A(\myring.inv_in[846] ));
 sg13g2_inv_1 \myring.inv_array[847]/sky_inverter/_0_  (.Y(\myring.inv_in[848] ),
    .A(\myring.inv_in[847] ));
 sg13g2_inv_1 \myring.inv_array[848]/sky_inverter/_0_  (.Y(\myring.inv_in[849] ),
    .A(\myring.inv_in[848] ));
 sg13g2_inv_1 \myring.inv_array[849]/sky_inverter/_0_  (.Y(\myring.inv_in[850] ),
    .A(\myring.inv_in[849] ));
 sg13g2_inv_1 \myring.inv_array[84]/sky_inverter/_0_  (.Y(\myring.inv_in[85] ),
    .A(\myring.inv_in[84] ));
 sg13g2_inv_1 \myring.inv_array[850]/sky_inverter/_0_  (.Y(\myring.inv_in[851] ),
    .A(\myring.inv_in[850] ));
 sg13g2_inv_1 \myring.inv_array[851]/sky_inverter/_0_  (.Y(\myring.inv_in[852] ),
    .A(\myring.inv_in[851] ));
 sg13g2_inv_1 \myring.inv_array[852]/sky_inverter/_0_  (.Y(\myring.inv_in[853] ),
    .A(\myring.inv_in[852] ));
 sg13g2_inv_1 \myring.inv_array[853]/sky_inverter/_0_  (.Y(\myring.inv_in[854] ),
    .A(\myring.inv_in[853] ));
 sg13g2_inv_1 \myring.inv_array[854]/sky_inverter/_0_  (.Y(\myring.inv_in[855] ),
    .A(\myring.inv_in[854] ));
 sg13g2_inv_1 \myring.inv_array[855]/sky_inverter/_0_  (.Y(\myring.inv_in[856] ),
    .A(\myring.inv_in[855] ));
 sg13g2_inv_1 \myring.inv_array[856]/sky_inverter/_0_  (.Y(\myring.inv_in[857] ),
    .A(\myring.inv_in[856] ));
 sg13g2_inv_1 \myring.inv_array[857]/sky_inverter/_0_  (.Y(\myring.inv_in[858] ),
    .A(\myring.inv_in[857] ));
 sg13g2_inv_1 \myring.inv_array[858]/sky_inverter/_0_  (.Y(\myring.inv_in[859] ),
    .A(\myring.inv_in[858] ));
 sg13g2_inv_1 \myring.inv_array[859]/sky_inverter/_0_  (.Y(\myring.inv_in[860] ),
    .A(\myring.inv_in[859] ));
 sg13g2_inv_1 \myring.inv_array[85]/sky_inverter/_0_  (.Y(\myring.inv_in[86] ),
    .A(\myring.inv_in[85] ));
 sg13g2_inv_1 \myring.inv_array[860]/sky_inverter/_0_  (.Y(\myring.inv_in[861] ),
    .A(\myring.inv_in[860] ));
 sg13g2_inv_1 \myring.inv_array[861]/sky_inverter/_0_  (.Y(\myring.inv_in[862] ),
    .A(\myring.inv_in[861] ));
 sg13g2_inv_1 \myring.inv_array[862]/sky_inverter/_0_  (.Y(\myring.inv_in[863] ),
    .A(\myring.inv_in[862] ));
 sg13g2_inv_1 \myring.inv_array[863]/sky_inverter/_0_  (.Y(\myring.inv_in[864] ),
    .A(\myring.inv_in[863] ));
 sg13g2_inv_1 \myring.inv_array[864]/sky_inverter/_0_  (.Y(\myring.inv_in[865] ),
    .A(\myring.inv_in[864] ));
 sg13g2_inv_1 \myring.inv_array[865]/sky_inverter/_0_  (.Y(\myring.inv_in[866] ),
    .A(\myring.inv_in[865] ));
 sg13g2_inv_1 \myring.inv_array[866]/sky_inverter/_0_  (.Y(\myring.inv_in[867] ),
    .A(\myring.inv_in[866] ));
 sg13g2_inv_1 \myring.inv_array[867]/sky_inverter/_0_  (.Y(\myring.inv_in[868] ),
    .A(\myring.inv_in[867] ));
 sg13g2_inv_1 \myring.inv_array[868]/sky_inverter/_0_  (.Y(\myring.inv_in[869] ),
    .A(\myring.inv_in[868] ));
 sg13g2_inv_1 \myring.inv_array[869]/sky_inverter/_0_  (.Y(\myring.inv_in[870] ),
    .A(\myring.inv_in[869] ));
 sg13g2_inv_1 \myring.inv_array[86]/sky_inverter/_0_  (.Y(\myring.inv_in[87] ),
    .A(\myring.inv_in[86] ));
 sg13g2_inv_1 \myring.inv_array[870]/sky_inverter/_0_  (.Y(\myring.inv_in[871] ),
    .A(\myring.inv_in[870] ));
 sg13g2_inv_1 \myring.inv_array[871]/sky_inverter/_0_  (.Y(\myring.inv_in[872] ),
    .A(\myring.inv_in[871] ));
 sg13g2_inv_1 \myring.inv_array[872]/sky_inverter/_0_  (.Y(\myring.inv_in[873] ),
    .A(\myring.inv_in[872] ));
 sg13g2_inv_1 \myring.inv_array[873]/sky_inverter/_0_  (.Y(\myring.inv_in[874] ),
    .A(\myring.inv_in[873] ));
 sg13g2_inv_1 \myring.inv_array[874]/sky_inverter/_0_  (.Y(\myring.inv_in[875] ),
    .A(\myring.inv_in[874] ));
 sg13g2_inv_1 \myring.inv_array[875]/sky_inverter/_0_  (.Y(\myring.inv_in[876] ),
    .A(\myring.inv_in[875] ));
 sg13g2_inv_1 \myring.inv_array[876]/sky_inverter/_0_  (.Y(\myring.inv_in[877] ),
    .A(\myring.inv_in[876] ));
 sg13g2_inv_1 \myring.inv_array[877]/sky_inverter/_0_  (.Y(\myring.inv_in[878] ),
    .A(\myring.inv_in[877] ));
 sg13g2_inv_1 \myring.inv_array[878]/sky_inverter/_0_  (.Y(\myring.inv_in[879] ),
    .A(\myring.inv_in[878] ));
 sg13g2_inv_1 \myring.inv_array[879]/sky_inverter/_0_  (.Y(\myring.inv_in[880] ),
    .A(\myring.inv_in[879] ));
 sg13g2_inv_1 \myring.inv_array[87]/sky_inverter/_0_  (.Y(\myring.inv_in[88] ),
    .A(\myring.inv_in[87] ));
 sg13g2_inv_1 \myring.inv_array[880]/sky_inverter/_0_  (.Y(\myring.inv_in[881] ),
    .A(\myring.inv_in[880] ));
 sg13g2_inv_1 \myring.inv_array[881]/sky_inverter/_0_  (.Y(\myring.inv_in[882] ),
    .A(\myring.inv_in[881] ));
 sg13g2_inv_1 \myring.inv_array[882]/sky_inverter/_0_  (.Y(\myring.inv_in[883] ),
    .A(\myring.inv_in[882] ));
 sg13g2_inv_1 \myring.inv_array[883]/sky_inverter/_0_  (.Y(\myring.inv_in[884] ),
    .A(\myring.inv_in[883] ));
 sg13g2_inv_1 \myring.inv_array[884]/sky_inverter/_0_  (.Y(\myring.inv_in[885] ),
    .A(\myring.inv_in[884] ));
 sg13g2_inv_1 \myring.inv_array[885]/sky_inverter/_0_  (.Y(\myring.inv_in[886] ),
    .A(\myring.inv_in[885] ));
 sg13g2_inv_1 \myring.inv_array[886]/sky_inverter/_0_  (.Y(\myring.inv_in[887] ),
    .A(\myring.inv_in[886] ));
 sg13g2_inv_1 \myring.inv_array[887]/sky_inverter/_0_  (.Y(\myring.inv_in[888] ),
    .A(\myring.inv_in[887] ));
 sg13g2_inv_1 \myring.inv_array[888]/sky_inverter/_0_  (.Y(\myring.inv_in[889] ),
    .A(\myring.inv_in[888] ));
 sg13g2_inv_1 \myring.inv_array[889]/sky_inverter/_0_  (.Y(\myring.inv_in[890] ),
    .A(\myring.inv_in[889] ));
 sg13g2_inv_1 \myring.inv_array[88]/sky_inverter/_0_  (.Y(\myring.inv_in[89] ),
    .A(\myring.inv_in[88] ));
 sg13g2_inv_1 \myring.inv_array[890]/sky_inverter/_0_  (.Y(\myring.inv_in[891] ),
    .A(\myring.inv_in[890] ));
 sg13g2_inv_1 \myring.inv_array[891]/sky_inverter/_0_  (.Y(\myring.inv_in[892] ),
    .A(\myring.inv_in[891] ));
 sg13g2_inv_1 \myring.inv_array[892]/sky_inverter/_0_  (.Y(\myring.inv_in[893] ),
    .A(\myring.inv_in[892] ));
 sg13g2_inv_1 \myring.inv_array[893]/sky_inverter/_0_  (.Y(\myring.inv_in[894] ),
    .A(\myring.inv_in[893] ));
 sg13g2_inv_1 \myring.inv_array[894]/sky_inverter/_0_  (.Y(\myring.inv_in[895] ),
    .A(\myring.inv_in[894] ));
 sg13g2_inv_1 \myring.inv_array[895]/sky_inverter/_0_  (.Y(\myring.inv_in[896] ),
    .A(\myring.inv_in[895] ));
 sg13g2_inv_1 \myring.inv_array[896]/sky_inverter/_0_  (.Y(\myring.inv_in[897] ),
    .A(\myring.inv_in[896] ));
 sg13g2_inv_1 \myring.inv_array[897]/sky_inverter/_0_  (.Y(\myring.inv_in[898] ),
    .A(\myring.inv_in[897] ));
 sg13g2_inv_1 \myring.inv_array[898]/sky_inverter/_0_  (.Y(\myring.inv_in[899] ),
    .A(\myring.inv_in[898] ));
 sg13g2_inv_1 \myring.inv_array[899]/sky_inverter/_0_  (.Y(\myring.inv_in[900] ),
    .A(\myring.inv_in[899] ));
 sg13g2_inv_1 \myring.inv_array[89]/sky_inverter/_0_  (.Y(\myring.inv_in[90] ),
    .A(\myring.inv_in[89] ));
 sg13g2_inv_1 \myring.inv_array[8]/sky_inverter/_0_  (.Y(\myring.inv_in[9] ),
    .A(\myring.inv_in[8] ));
 sg13g2_inv_1 \myring.inv_array[900]/sky_inverter/_0_  (.Y(\myring.inv_in[901] ),
    .A(\myring.inv_in[900] ));
 sg13g2_inv_1 \myring.inv_array[901]/sky_inverter/_0_  (.Y(\myring.inv_in[902] ),
    .A(\myring.inv_in[901] ));
 sg13g2_inv_1 \myring.inv_array[902]/sky_inverter/_0_  (.Y(\myring.inv_in[903] ),
    .A(\myring.inv_in[902] ));
 sg13g2_inv_1 \myring.inv_array[903]/sky_inverter/_0_  (.Y(\myring.inv_in[904] ),
    .A(\myring.inv_in[903] ));
 sg13g2_inv_1 \myring.inv_array[904]/sky_inverter/_0_  (.Y(\myring.inv_in[905] ),
    .A(\myring.inv_in[904] ));
 sg13g2_inv_1 \myring.inv_array[905]/sky_inverter/_0_  (.Y(\myring.inv_in[906] ),
    .A(\myring.inv_in[905] ));
 sg13g2_inv_1 \myring.inv_array[906]/sky_inverter/_0_  (.Y(\myring.inv_in[907] ),
    .A(\myring.inv_in[906] ));
 sg13g2_inv_1 \myring.inv_array[907]/sky_inverter/_0_  (.Y(\myring.inv_in[908] ),
    .A(\myring.inv_in[907] ));
 sg13g2_inv_1 \myring.inv_array[908]/sky_inverter/_0_  (.Y(\myring.inv_in[909] ),
    .A(\myring.inv_in[908] ));
 sg13g2_inv_1 \myring.inv_array[909]/sky_inverter/_0_  (.Y(\myring.inv_in[910] ),
    .A(\myring.inv_in[909] ));
 sg13g2_inv_1 \myring.inv_array[90]/sky_inverter/_0_  (.Y(\myring.inv_in[91] ),
    .A(\myring.inv_in[90] ));
 sg13g2_inv_1 \myring.inv_array[910]/sky_inverter/_0_  (.Y(\myring.inv_in[911] ),
    .A(\myring.inv_in[910] ));
 sg13g2_inv_1 \myring.inv_array[911]/sky_inverter/_0_  (.Y(\myring.inv_in[912] ),
    .A(\myring.inv_in[911] ));
 sg13g2_inv_1 \myring.inv_array[912]/sky_inverter/_0_  (.Y(\myring.inv_in[913] ),
    .A(\myring.inv_in[912] ));
 sg13g2_inv_1 \myring.inv_array[913]/sky_inverter/_0_  (.Y(\myring.inv_in[914] ),
    .A(\myring.inv_in[913] ));
 sg13g2_inv_1 \myring.inv_array[914]/sky_inverter/_0_  (.Y(\myring.inv_in[915] ),
    .A(\myring.inv_in[914] ));
 sg13g2_inv_1 \myring.inv_array[915]/sky_inverter/_0_  (.Y(\myring.inv_in[916] ),
    .A(\myring.inv_in[915] ));
 sg13g2_inv_1 \myring.inv_array[916]/sky_inverter/_0_  (.Y(\myring.inv_in[917] ),
    .A(\myring.inv_in[916] ));
 sg13g2_inv_1 \myring.inv_array[917]/sky_inverter/_0_  (.Y(\myring.inv_in[918] ),
    .A(\myring.inv_in[917] ));
 sg13g2_inv_1 \myring.inv_array[918]/sky_inverter/_0_  (.Y(\myring.inv_in[919] ),
    .A(\myring.inv_in[918] ));
 sg13g2_inv_1 \myring.inv_array[919]/sky_inverter/_0_  (.Y(\myring.inv_in[920] ),
    .A(\myring.inv_in[919] ));
 sg13g2_inv_1 \myring.inv_array[91]/sky_inverter/_0_  (.Y(\myring.inv_in[92] ),
    .A(\myring.inv_in[91] ));
 sg13g2_inv_1 \myring.inv_array[920]/sky_inverter/_0_  (.Y(\myring.inv_in[921] ),
    .A(\myring.inv_in[920] ));
 sg13g2_inv_1 \myring.inv_array[921]/sky_inverter/_0_  (.Y(\myring.inv_in[922] ),
    .A(\myring.inv_in[921] ));
 sg13g2_inv_1 \myring.inv_array[922]/sky_inverter/_0_  (.Y(\myring.inv_in[923] ),
    .A(\myring.inv_in[922] ));
 sg13g2_inv_1 \myring.inv_array[923]/sky_inverter/_0_  (.Y(\myring.inv_in[924] ),
    .A(\myring.inv_in[923] ));
 sg13g2_inv_1 \myring.inv_array[924]/sky_inverter/_0_  (.Y(\myring.inv_in[925] ),
    .A(\myring.inv_in[924] ));
 sg13g2_inv_1 \myring.inv_array[925]/sky_inverter/_0_  (.Y(\myring.inv_in[926] ),
    .A(\myring.inv_in[925] ));
 sg13g2_inv_1 \myring.inv_array[926]/sky_inverter/_0_  (.Y(\myring.inv_in[927] ),
    .A(\myring.inv_in[926] ));
 sg13g2_inv_1 \myring.inv_array[927]/sky_inverter/_0_  (.Y(\myring.inv_in[928] ),
    .A(\myring.inv_in[927] ));
 sg13g2_inv_1 \myring.inv_array[928]/sky_inverter/_0_  (.Y(\myring.inv_in[929] ),
    .A(\myring.inv_in[928] ));
 sg13g2_inv_1 \myring.inv_array[929]/sky_inverter/_0_  (.Y(\myring.inv_in[930] ),
    .A(\myring.inv_in[929] ));
 sg13g2_inv_1 \myring.inv_array[92]/sky_inverter/_0_  (.Y(\myring.inv_in[93] ),
    .A(\myring.inv_in[92] ));
 sg13g2_inv_1 \myring.inv_array[930]/sky_inverter/_0_  (.Y(\myring.inv_in[931] ),
    .A(\myring.inv_in[930] ));
 sg13g2_inv_1 \myring.inv_array[931]/sky_inverter/_0_  (.Y(\myring.inv_in[932] ),
    .A(\myring.inv_in[931] ));
 sg13g2_inv_1 \myring.inv_array[932]/sky_inverter/_0_  (.Y(\myring.inv_in[933] ),
    .A(\myring.inv_in[932] ));
 sg13g2_inv_1 \myring.inv_array[933]/sky_inverter/_0_  (.Y(\myring.inv_in[934] ),
    .A(\myring.inv_in[933] ));
 sg13g2_inv_1 \myring.inv_array[934]/sky_inverter/_0_  (.Y(\myring.inv_in[935] ),
    .A(\myring.inv_in[934] ));
 sg13g2_inv_1 \myring.inv_array[935]/sky_inverter/_0_  (.Y(\myring.inv_in[936] ),
    .A(\myring.inv_in[935] ));
 sg13g2_inv_1 \myring.inv_array[936]/sky_inverter/_0_  (.Y(\myring.inv_in[937] ),
    .A(\myring.inv_in[936] ));
 sg13g2_inv_1 \myring.inv_array[937]/sky_inverter/_0_  (.Y(\myring.inv_in[938] ),
    .A(\myring.inv_in[937] ));
 sg13g2_inv_1 \myring.inv_array[938]/sky_inverter/_0_  (.Y(\myring.inv_in[939] ),
    .A(\myring.inv_in[938] ));
 sg13g2_inv_1 \myring.inv_array[939]/sky_inverter/_0_  (.Y(\myring.inv_in[940] ),
    .A(\myring.inv_in[939] ));
 sg13g2_inv_1 \myring.inv_array[93]/sky_inverter/_0_  (.Y(\myring.inv_in[94] ),
    .A(\myring.inv_in[93] ));
 sg13g2_inv_1 \myring.inv_array[940]/sky_inverter/_0_  (.Y(\myring.inv_in[941] ),
    .A(\myring.inv_in[940] ));
 sg13g2_inv_1 \myring.inv_array[941]/sky_inverter/_0_  (.Y(\myring.inv_in[942] ),
    .A(\myring.inv_in[941] ));
 sg13g2_inv_1 \myring.inv_array[942]/sky_inverter/_0_  (.Y(\myring.inv_in[943] ),
    .A(\myring.inv_in[942] ));
 sg13g2_inv_1 \myring.inv_array[943]/sky_inverter/_0_  (.Y(\myring.inv_in[944] ),
    .A(\myring.inv_in[943] ));
 sg13g2_inv_1 \myring.inv_array[944]/sky_inverter/_0_  (.Y(\myring.inv_in[945] ),
    .A(\myring.inv_in[944] ));
 sg13g2_inv_1 \myring.inv_array[945]/sky_inverter/_0_  (.Y(\myring.inv_in[946] ),
    .A(\myring.inv_in[945] ));
 sg13g2_inv_1 \myring.inv_array[946]/sky_inverter/_0_  (.Y(\myring.inv_in[947] ),
    .A(\myring.inv_in[946] ));
 sg13g2_inv_1 \myring.inv_array[947]/sky_inverter/_0_  (.Y(\myring.inv_in[948] ),
    .A(\myring.inv_in[947] ));
 sg13g2_inv_1 \myring.inv_array[948]/sky_inverter/_0_  (.Y(\myring.inv_in[949] ),
    .A(\myring.inv_in[948] ));
 sg13g2_inv_1 \myring.inv_array[949]/sky_inverter/_0_  (.Y(\myring.inv_in[950] ),
    .A(\myring.inv_in[949] ));
 sg13g2_inv_1 \myring.inv_array[94]/sky_inverter/_0_  (.Y(\myring.inv_in[95] ),
    .A(\myring.inv_in[94] ));
 sg13g2_inv_1 \myring.inv_array[950]/sky_inverter/_0_  (.Y(\myring.inv_in[951] ),
    .A(\myring.inv_in[950] ));
 sg13g2_inv_1 \myring.inv_array[951]/sky_inverter/_0_  (.Y(\myring.inv_in[952] ),
    .A(\myring.inv_in[951] ));
 sg13g2_inv_1 \myring.inv_array[952]/sky_inverter/_0_  (.Y(\myring.inv_in[953] ),
    .A(\myring.inv_in[952] ));
 sg13g2_inv_1 \myring.inv_array[953]/sky_inverter/_0_  (.Y(\myring.inv_in[954] ),
    .A(\myring.inv_in[953] ));
 sg13g2_inv_1 \myring.inv_array[954]/sky_inverter/_0_  (.Y(\myring.inv_in[955] ),
    .A(\myring.inv_in[954] ));
 sg13g2_inv_1 \myring.inv_array[955]/sky_inverter/_0_  (.Y(\myring.inv_in[956] ),
    .A(\myring.inv_in[955] ));
 sg13g2_inv_1 \myring.inv_array[956]/sky_inverter/_0_  (.Y(\myring.inv_in[957] ),
    .A(\myring.inv_in[956] ));
 sg13g2_inv_1 \myring.inv_array[957]/sky_inverter/_0_  (.Y(\myring.inv_in[958] ),
    .A(\myring.inv_in[957] ));
 sg13g2_inv_1 \myring.inv_array[958]/sky_inverter/_0_  (.Y(\myring.inv_in[959] ),
    .A(\myring.inv_in[958] ));
 sg13g2_inv_1 \myring.inv_array[959]/sky_inverter/_0_  (.Y(\myring.inv_in[960] ),
    .A(\myring.inv_in[959] ));
 sg13g2_inv_1 \myring.inv_array[95]/sky_inverter/_0_  (.Y(\myring.inv_in[96] ),
    .A(\myring.inv_in[95] ));
 sg13g2_inv_1 \myring.inv_array[960]/sky_inverter/_0_  (.Y(\myring.inv_in[961] ),
    .A(\myring.inv_in[960] ));
 sg13g2_inv_1 \myring.inv_array[961]/sky_inverter/_0_  (.Y(\myring.inv_in[962] ),
    .A(\myring.inv_in[961] ));
 sg13g2_inv_1 \myring.inv_array[962]/sky_inverter/_0_  (.Y(\myring.inv_in[963] ),
    .A(\myring.inv_in[962] ));
 sg13g2_inv_1 \myring.inv_array[963]/sky_inverter/_0_  (.Y(\myring.inv_in[964] ),
    .A(\myring.inv_in[963] ));
 sg13g2_inv_1 \myring.inv_array[964]/sky_inverter/_0_  (.Y(\myring.inv_in[965] ),
    .A(\myring.inv_in[964] ));
 sg13g2_inv_1 \myring.inv_array[965]/sky_inverter/_0_  (.Y(\myring.inv_in[966] ),
    .A(\myring.inv_in[965] ));
 sg13g2_inv_1 \myring.inv_array[966]/sky_inverter/_0_  (.Y(\myring.inv_in[967] ),
    .A(\myring.inv_in[966] ));
 sg13g2_inv_1 \myring.inv_array[967]/sky_inverter/_0_  (.Y(\myring.inv_in[968] ),
    .A(\myring.inv_in[967] ));
 sg13g2_inv_1 \myring.inv_array[968]/sky_inverter/_0_  (.Y(\myring.inv_in[969] ),
    .A(\myring.inv_in[968] ));
 sg13g2_inv_1 \myring.inv_array[969]/sky_inverter/_0_  (.Y(\myring.inv_in[970] ),
    .A(\myring.inv_in[969] ));
 sg13g2_inv_1 \myring.inv_array[96]/sky_inverter/_0_  (.Y(\myring.inv_in[97] ),
    .A(\myring.inv_in[96] ));
 sg13g2_inv_1 \myring.inv_array[970]/sky_inverter/_0_  (.Y(\myring.inv_in[971] ),
    .A(\myring.inv_in[970] ));
 sg13g2_inv_1 \myring.inv_array[971]/sky_inverter/_0_  (.Y(\myring.inv_in[972] ),
    .A(\myring.inv_in[971] ));
 sg13g2_inv_1 \myring.inv_array[972]/sky_inverter/_0_  (.Y(\myring.inv_in[973] ),
    .A(\myring.inv_in[972] ));
 sg13g2_inv_1 \myring.inv_array[973]/sky_inverter/_0_  (.Y(\myring.inv_in[974] ),
    .A(\myring.inv_in[973] ));
 sg13g2_inv_1 \myring.inv_array[974]/sky_inverter/_0_  (.Y(\myring.inv_in[975] ),
    .A(\myring.inv_in[974] ));
 sg13g2_inv_1 \myring.inv_array[975]/sky_inverter/_0_  (.Y(\myring.inv_in[976] ),
    .A(\myring.inv_in[975] ));
 sg13g2_inv_1 \myring.inv_array[976]/sky_inverter/_0_  (.Y(\myring.inv_in[977] ),
    .A(\myring.inv_in[976] ));
 sg13g2_inv_1 \myring.inv_array[977]/sky_inverter/_0_  (.Y(\myring.inv_in[978] ),
    .A(\myring.inv_in[977] ));
 sg13g2_inv_1 \myring.inv_array[978]/sky_inverter/_0_  (.Y(\myring.inv_in[979] ),
    .A(\myring.inv_in[978] ));
 sg13g2_inv_1 \myring.inv_array[979]/sky_inverter/_0_  (.Y(\myring.inv_in[980] ),
    .A(\myring.inv_in[979] ));
 sg13g2_inv_1 \myring.inv_array[97]/sky_inverter/_0_  (.Y(\myring.inv_in[98] ),
    .A(\myring.inv_in[97] ));
 sg13g2_inv_1 \myring.inv_array[980]/sky_inverter/_0_  (.Y(\myring.inv_in[981] ),
    .A(\myring.inv_in[980] ));
 sg13g2_inv_1 \myring.inv_array[981]/sky_inverter/_0_  (.Y(\myring.inv_in[982] ),
    .A(\myring.inv_in[981] ));
 sg13g2_inv_1 \myring.inv_array[982]/sky_inverter/_0_  (.Y(\myring.inv_in[983] ),
    .A(\myring.inv_in[982] ));
 sg13g2_inv_1 \myring.inv_array[983]/sky_inverter/_0_  (.Y(\myring.inv_in[984] ),
    .A(\myring.inv_in[983] ));
 sg13g2_inv_1 \myring.inv_array[984]/sky_inverter/_0_  (.Y(\myring.inv_in[985] ),
    .A(\myring.inv_in[984] ));
 sg13g2_inv_1 \myring.inv_array[985]/sky_inverter/_0_  (.Y(\myring.inv_in[986] ),
    .A(\myring.inv_in[985] ));
 sg13g2_inv_1 \myring.inv_array[986]/sky_inverter/_0_  (.Y(\myring.inv_in[987] ),
    .A(\myring.inv_in[986] ));
 sg13g2_inv_1 \myring.inv_array[987]/sky_inverter/_0_  (.Y(\myring.inv_in[988] ),
    .A(\myring.inv_in[987] ));
 sg13g2_inv_1 \myring.inv_array[988]/sky_inverter/_0_  (.Y(\myring.inv_in[989] ),
    .A(\myring.inv_in[988] ));
 sg13g2_inv_1 \myring.inv_array[989]/sky_inverter/_0_  (.Y(\myring.inv_in[990] ),
    .A(\myring.inv_in[989] ));
 sg13g2_inv_1 \myring.inv_array[98]/sky_inverter/_0_  (.Y(\myring.inv_in[99] ),
    .A(\myring.inv_in[98] ));
 sg13g2_inv_1 \myring.inv_array[990]/sky_inverter/_0_  (.Y(\myring.inv_in[991] ),
    .A(\myring.inv_in[990] ));
 sg13g2_inv_1 \myring.inv_array[991]/sky_inverter/_0_  (.Y(\myring.inv_in[992] ),
    .A(\myring.inv_in[991] ));
 sg13g2_inv_1 \myring.inv_array[992]/sky_inverter/_0_  (.Y(\myring.inv_in[993] ),
    .A(\myring.inv_in[992] ));
 sg13g2_inv_1 \myring.inv_array[993]/sky_inverter/_0_  (.Y(\myring.inv_in[994] ),
    .A(\myring.inv_in[993] ));
 sg13g2_inv_1 \myring.inv_array[994]/sky_inverter/_0_  (.Y(\myring.inv_in[995] ),
    .A(\myring.inv_in[994] ));
 sg13g2_inv_1 \myring.inv_array[995]/sky_inverter/_0_  (.Y(\myring.inv_in[996] ),
    .A(\myring.inv_in[995] ));
 sg13g2_inv_1 \myring.inv_array[996]/sky_inverter/_0_  (.Y(\myring.inv_in[997] ),
    .A(\myring.inv_in[996] ));
 sg13g2_inv_1 \myring.inv_array[997]/sky_inverter/_0_  (.Y(\myring.inv_in[998] ),
    .A(\myring.inv_in[997] ));
 sg13g2_inv_1 \myring.inv_array[998]/sky_inverter/_0_  (.Y(\myring.inv_in[999] ),
    .A(\myring.inv_in[998] ));
 sg13g2_inv_1 \myring.inv_array[999]/sky_inverter/_0_  (.Y(\myring.inv_in[1000] ),
    .A(\myring.inv_in[999] ));
 sg13g2_inv_1 \myring.inv_array[99]/sky_inverter/_0_  (.Y(\myring.inv_in[100] ),
    .A(\myring.inv_in[99] ));
 sg13g2_inv_1 \myring.inv_array[9]/sky_inverter/_0_  (.Y(\myring.inv_in[10] ),
    .A(\myring.inv_in[9] ));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[0]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[2]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[3]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[4]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[5]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[6]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(ui_in[7]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[0]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[1]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[2]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[3]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[4]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[5]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(uio_in[6]),
    .X(net17));
 sg13g2_buf_1 input18 (.A(uio_in[7]),
    .X(net18));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc_19 (.L_LO(net19));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_4 FILLER_9_147 ();
 sg13g2_fill_2 FILLER_9_151 ();
 sg13g2_fill_1 FILLER_9_159 ();
 sg13g2_decap_4 FILLER_9_163 ();
 sg13g2_fill_2 FILLER_9_167 ();
 sg13g2_fill_1 FILLER_9_172 ();
 sg13g2_fill_1 FILLER_9_176 ();
 sg13g2_decap_4 FILLER_9_180 ();
 sg13g2_decap_4 FILLER_9_190 ();
 sg13g2_fill_2 FILLER_9_194 ();
 sg13g2_decap_8 FILLER_9_199 ();
 sg13g2_decap_8 FILLER_9_206 ();
 sg13g2_decap_8 FILLER_9_213 ();
 sg13g2_decap_8 FILLER_9_220 ();
 sg13g2_decap_8 FILLER_9_227 ();
 sg13g2_decap_8 FILLER_9_234 ();
 sg13g2_decap_8 FILLER_9_241 ();
 sg13g2_decap_8 FILLER_9_248 ();
 sg13g2_decap_8 FILLER_9_255 ();
 sg13g2_decap_8 FILLER_9_262 ();
 sg13g2_decap_8 FILLER_9_269 ();
 sg13g2_decap_8 FILLER_9_276 ();
 sg13g2_decap_8 FILLER_9_283 ();
 sg13g2_decap_8 FILLER_9_290 ();
 sg13g2_decap_8 FILLER_9_297 ();
 sg13g2_decap_8 FILLER_9_304 ();
 sg13g2_decap_8 FILLER_9_311 ();
 sg13g2_decap_8 FILLER_9_318 ();
 sg13g2_decap_8 FILLER_9_325 ();
 sg13g2_decap_8 FILLER_9_332 ();
 sg13g2_decap_8 FILLER_9_339 ();
 sg13g2_decap_8 FILLER_9_346 ();
 sg13g2_decap_8 FILLER_9_353 ();
 sg13g2_decap_8 FILLER_9_360 ();
 sg13g2_decap_8 FILLER_9_367 ();
 sg13g2_decap_8 FILLER_9_374 ();
 sg13g2_decap_8 FILLER_9_381 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_4 FILLER_10_140 ();
 sg13g2_fill_2 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_227 ();
 sg13g2_decap_8 FILLER_10_234 ();
 sg13g2_decap_8 FILLER_10_241 ();
 sg13g2_decap_8 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_255 ();
 sg13g2_decap_8 FILLER_10_262 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_decap_8 FILLER_10_290 ();
 sg13g2_decap_8 FILLER_10_297 ();
 sg13g2_decap_8 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_311 ();
 sg13g2_decap_8 FILLER_10_318 ();
 sg13g2_decap_8 FILLER_10_325 ();
 sg13g2_decap_8 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_4 FILLER_11_140 ();
 sg13g2_decap_4 FILLER_11_165 ();
 sg13g2_fill_2 FILLER_11_169 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_176 ();
 sg13g2_decap_8 FILLER_11_180 ();
 sg13g2_decap_8 FILLER_11_187 ();
 sg13g2_decap_8 FILLER_11_194 ();
 sg13g2_decap_8 FILLER_11_201 ();
 sg13g2_decap_4 FILLER_11_208 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_decap_8 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_241 ();
 sg13g2_decap_8 FILLER_11_248 ();
 sg13g2_decap_8 FILLER_11_255 ();
 sg13g2_decap_8 FILLER_11_262 ();
 sg13g2_decap_8 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_283 ();
 sg13g2_decap_8 FILLER_11_290 ();
 sg13g2_decap_8 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_4 FILLER_12_140 ();
 sg13g2_fill_1 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_208 ();
 sg13g2_fill_2 FILLER_12_215 ();
 sg13g2_fill_1 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_4 FILLER_13_147 ();
 sg13g2_fill_2 FILLER_13_151 ();
 sg13g2_decap_8 FILLER_13_156 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_fill_1 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_169 ();
 sg13g2_decap_8 FILLER_13_176 ();
 sg13g2_decap_8 FILLER_13_183 ();
 sg13g2_decap_8 FILLER_13_190 ();
 sg13g2_fill_1 FILLER_13_197 ();
 sg13g2_decap_8 FILLER_13_213 ();
 sg13g2_fill_2 FILLER_13_220 ();
 sg13g2_decap_8 FILLER_13_240 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_decap_8 FILLER_13_254 ();
 sg13g2_decap_8 FILLER_13_261 ();
 sg13g2_decap_8 FILLER_13_268 ();
 sg13g2_decap_8 FILLER_13_275 ();
 sg13g2_decap_8 FILLER_13_282 ();
 sg13g2_decap_8 FILLER_13_289 ();
 sg13g2_decap_8 FILLER_13_296 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_310 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_fill_2 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_216 ();
 sg13g2_fill_1 FILLER_14_223 ();
 sg13g2_decap_8 FILLER_14_242 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_decap_8 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_4 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_215 ();
 sg13g2_decap_8 FILLER_15_243 ();
 sg13g2_decap_8 FILLER_15_250 ();
 sg13g2_decap_8 FILLER_15_257 ();
 sg13g2_decap_8 FILLER_15_264 ();
 sg13g2_decap_8 FILLER_15_271 ();
 sg13g2_decap_8 FILLER_15_278 ();
 sg13g2_decap_8 FILLER_15_285 ();
 sg13g2_decap_8 FILLER_15_292 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_161 ();
 sg13g2_fill_2 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_168 ();
 sg13g2_fill_1 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_176 ();
 sg13g2_fill_2 FILLER_16_183 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_fill_1 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_194 ();
 sg13g2_decap_8 FILLER_17_201 ();
 sg13g2_decap_4 FILLER_17_208 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_4 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_159 ();
 sg13g2_fill_2 FILLER_18_166 ();
 sg13g2_fill_1 FILLER_18_168 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_decap_4 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_181 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_decap_4 FILLER_18_206 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_4 FILLER_18_242 ();
 sg13g2_fill_2 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_251 ();
 sg13g2_decap_4 FILLER_18_255 ();
 sg13g2_fill_2 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_264 ();
 sg13g2_decap_8 FILLER_18_271 ();
 sg13g2_decap_8 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_292 ();
 sg13g2_decap_8 FILLER_18_299 ();
 sg13g2_decap_8 FILLER_18_306 ();
 sg13g2_decap_8 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_4 FILLER_19_133 ();
 sg13g2_fill_2 FILLER_19_137 ();
 sg13g2_fill_2 FILLER_19_160 ();
 sg13g2_fill_1 FILLER_19_162 ();
 sg13g2_fill_1 FILLER_19_205 ();
 sg13g2_decap_4 FILLER_19_212 ();
 sg13g2_decap_8 FILLER_19_219 ();
 sg13g2_fill_2 FILLER_19_229 ();
 sg13g2_fill_1 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_309 ();
 sg13g2_decap_8 FILLER_19_316 ();
 sg13g2_decap_8 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_4 FILLER_20_112 ();
 sg13g2_fill_1 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_fill_2 FILLER_20_137 ();
 sg13g2_fill_2 FILLER_20_154 ();
 sg13g2_fill_2 FILLER_20_171 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_fill_1 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_1 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_139 ();
 sg13g2_decap_8 FILLER_21_146 ();
 sg13g2_decap_4 FILLER_21_153 ();
 sg13g2_fill_2 FILLER_21_157 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_4 FILLER_21_210 ();
 sg13g2_fill_1 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_decap_8 FILLER_21_237 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_fill_2 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_100 ();
 sg13g2_decap_8 FILLER_22_122 ();
 sg13g2_decap_8 FILLER_22_129 ();
 sg13g2_fill_1 FILLER_22_136 ();
 sg13g2_fill_1 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_4 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_190 ();
 sg13g2_fill_1 FILLER_22_197 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_fill_2 FILLER_22_242 ();
 sg13g2_decap_4 FILLER_22_259 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_267 ();
 sg13g2_decap_8 FILLER_22_274 ();
 sg13g2_decap_8 FILLER_22_281 ();
 sg13g2_decap_8 FILLER_22_288 ();
 sg13g2_decap_8 FILLER_22_295 ();
 sg13g2_decap_8 FILLER_22_302 ();
 sg13g2_decap_8 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_98 ();
 sg13g2_fill_2 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_126 ();
 sg13g2_fill_1 FILLER_23_128 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_151 ();
 sg13g2_fill_1 FILLER_23_153 ();
 sg13g2_decap_8 FILLER_23_181 ();
 sg13g2_decap_4 FILLER_23_188 ();
 sg13g2_fill_2 FILLER_23_192 ();
 sg13g2_decap_8 FILLER_23_212 ();
 sg13g2_decap_4 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_267 ();
 sg13g2_fill_1 FILLER_23_272 ();
 sg13g2_decap_8 FILLER_23_276 ();
 sg13g2_decap_8 FILLER_23_283 ();
 sg13g2_decap_8 FILLER_23_290 ();
 sg13g2_decap_8 FILLER_23_297 ();
 sg13g2_decap_8 FILLER_23_304 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_decap_8 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_fill_2 FILLER_24_115 ();
 sg13g2_fill_1 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_decap_8 FILLER_24_152 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_decap_8 FILLER_24_191 ();
 sg13g2_decap_8 FILLER_24_213 ();
 sg13g2_decap_4 FILLER_24_220 ();
 sg13g2_fill_2 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_244 ();
 sg13g2_decap_4 FILLER_24_251 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_328 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_114 ();
 sg13g2_fill_1 FILLER_25_131 ();
 sg13g2_decap_8 FILLER_25_138 ();
 sg13g2_decap_4 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_160 ();
 sg13g2_fill_2 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_decap_4 FILLER_25_191 ();
 sg13g2_fill_2 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_252 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_fill_1 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_4 FILLER_25_272 ();
 sg13g2_decap_4 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_4 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_192 ();
 sg13g2_decap_8 FILLER_26_199 ();
 sg13g2_decap_8 FILLER_26_206 ();
 sg13g2_fill_2 FILLER_26_213 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_decap_4 FILLER_26_225 ();
 sg13g2_fill_2 FILLER_26_229 ();
 sg13g2_decap_8 FILLER_26_234 ();
 sg13g2_fill_1 FILLER_26_241 ();
 sg13g2_decap_4 FILLER_26_275 ();
 sg13g2_fill_2 FILLER_26_279 ();
 sg13g2_fill_2 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_303 ();
 sg13g2_fill_2 FILLER_26_310 ();
 sg13g2_fill_1 FILLER_26_312 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_173 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_decap_8 FILLER_27_256 ();
 sg13g2_fill_1 FILLER_27_263 ();
 sg13g2_decap_8 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_fill_2 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_135 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_165 ();
 sg13g2_fill_2 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_181 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_4 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_250 ();
 sg13g2_decap_8 FILLER_28_257 ();
 sg13g2_fill_1 FILLER_28_264 ();
 sg13g2_fill_1 FILLER_28_286 ();
 sg13g2_decap_8 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_319 ();
 sg13g2_decap_8 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_28_333 ();
 sg13g2_decap_8 FILLER_28_340 ();
 sg13g2_decap_8 FILLER_28_347 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_361 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_4 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_decap_4 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_218 ();
 sg13g2_decap_8 FILLER_29_246 ();
 sg13g2_decap_8 FILLER_29_253 ();
 sg13g2_decap_8 FILLER_29_260 ();
 sg13g2_decap_4 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_296 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_decap_8 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_decap_8 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_29_352 ();
 sg13g2_decap_8 FILLER_29_359 ();
 sg13g2_decap_8 FILLER_29_366 ();
 sg13g2_decap_8 FILLER_29_373 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_4 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_158 ();
 sg13g2_fill_2 FILLER_30_163 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_4 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_190 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_fill_1 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_240 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_267 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_1 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_283 ();
 sg13g2_decap_8 FILLER_30_290 ();
 sg13g2_decap_8 FILLER_30_297 ();
 sg13g2_decap_8 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_311 ();
 sg13g2_decap_8 FILLER_30_318 ();
 sg13g2_decap_8 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_fill_2 FILLER_31_189 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_fill_2 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_decap_4 FILLER_31_290 ();
 sg13g2_fill_1 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_4 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_340 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_351 ();
 sg13g2_decap_8 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_365 ();
 sg13g2_decap_8 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_31_400 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_4 FILLER_32_182 ();
 sg13g2_fill_1 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_208 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_decap_8 FILLER_32_225 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_234 ();
 sg13g2_decap_8 FILLER_32_241 ();
 sg13g2_decap_8 FILLER_32_248 ();
 sg13g2_decap_4 FILLER_32_255 ();
 sg13g2_decap_8 FILLER_32_264 ();
 sg13g2_decap_8 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_311 ();
 sg13g2_decap_4 FILLER_32_318 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_fill_1 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_174 ();
 sg13g2_decap_8 FILLER_33_181 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_decap_4 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_decap_4 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_300 ();
 sg13g2_decap_8 FILLER_33_332 ();
 sg13g2_decap_8 FILLER_33_339 ();
 sg13g2_decap_4 FILLER_33_346 ();
 sg13g2_fill_1 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_133 ();
 sg13g2_decap_4 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_decap_4 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_209 ();
 sg13g2_decap_8 FILLER_34_225 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_decap_8 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_282 ();
 sg13g2_fill_1 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_303 ();
 sg13g2_decap_4 FILLER_34_310 ();
 sg13g2_decap_4 FILLER_34_317 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_decap_4 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_fill_2 FILLER_34_338 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_4 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_133 ();
 sg13g2_fill_1 FILLER_35_135 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_174 ();
 sg13g2_decap_4 FILLER_35_181 ();
 sg13g2_fill_2 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_190 ();
 sg13g2_decap_8 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_1 FILLER_35_206 ();
 sg13g2_decap_8 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_251 ();
 sg13g2_fill_2 FILLER_35_258 ();
 sg13g2_fill_1 FILLER_35_260 ();
 sg13g2_fill_1 FILLER_35_267 ();
 sg13g2_decap_4 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_288 ();
 sg13g2_fill_2 FILLER_35_307 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_205 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_decap_4 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_275 ();
 sg13g2_decap_4 FILLER_36_282 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_330 ();
 sg13g2_decap_4 FILLER_36_337 ();
 sg13g2_decap_8 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_351 ();
 sg13g2_decap_8 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_4 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_123 ();
 sg13g2_fill_1 FILLER_37_142 ();
 sg13g2_decap_8 FILLER_37_176 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_fill_2 FILLER_37_205 ();
 sg13g2_fill_2 FILLER_37_213 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_4 FILLER_37_231 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_decap_8 FILLER_37_281 ();
 sg13g2_fill_2 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_1 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_fill_1 FILLER_38_196 ();
 sg13g2_fill_1 FILLER_38_204 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_decap_4 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_235 ();
 sg13g2_fill_1 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_263 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_decap_4 FILLER_38_276 ();
 sg13g2_decap_4 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_decap_4 FILLER_38_332 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_decap_4 FILLER_38_348 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_4 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_4 FILLER_38_387 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net19;
 assign uio_oe[1] = net20;
 assign uio_oe[2] = net21;
 assign uio_oe[3] = net22;
 assign uio_oe[4] = net23;
 assign uio_oe[5] = net24;
 assign uio_oe[6] = net25;
 assign uio_oe[7] = net26;
 assign uio_out[0] = net27;
 assign uio_out[1] = net28;
 assign uio_out[2] = net29;
 assign uio_out[3] = net30;
 assign uio_out[4] = net31;
 assign uio_out[5] = net32;
 assign uio_out[6] = net33;
 assign uio_out[7] = net34;
 assign uo_out[2] = net35;
 assign uo_out[3] = net36;
 assign uo_out[4] = net37;
 assign uo_out[5] = net38;
 assign uo_out[6] = net39;
 assign uo_out[7] = net40;
endmodule

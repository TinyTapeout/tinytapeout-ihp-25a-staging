module tt_um_UartMain (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire clknet_0_clk;
 wire \e.buf_.dataReg[0] ;
 wire \e.buf_.dataReg[1] ;
 wire \e.buf_.dataReg[2] ;
 wire \e.buf_.dataReg[3] ;
 wire \e.buf_.dataReg[4] ;
 wire \e.buf_.dataReg[5] ;
 wire \e.buf_.dataReg[6] ;
 wire \e.buf_.dataReg[7] ;
 wire \e.buf_.io_in_bits[0] ;
 wire \e.buf_.io_in_bits[1] ;
 wire \e.buf_.io_in_bits[2] ;
 wire \e.buf_.io_in_bits[3] ;
 wire \e.buf_.io_in_bits[4] ;
 wire \e.buf_.io_in_bits[5] ;
 wire \e.buf_.io_in_bits[6] ;
 wire \e.buf_.io_in_bits[7] ;
 wire \e.buf_.io_in_valid ;
 wire \e.buf_.io_out_valid ;
 wire \e.io_txd ;
 wire \e.key[0] ;
 wire \e.key[1] ;
 wire \e.key[2] ;
 wire \e.key[3] ;
 wire \e.key[4] ;
 wire \e.key[5] ;
 wire \e.key[6] ;
 wire \e.key[7] ;
 wire \e.rx.bitsReg[0] ;
 wire \e.rx.bitsReg[1] ;
 wire \e.rx.bitsReg[2] ;
 wire \e.rx.bitsReg[3] ;
 wire \e.rx.cntReg[0] ;
 wire \e.rx.cntReg[10] ;
 wire \e.rx.cntReg[11] ;
 wire \e.rx.cntReg[12] ;
 wire \e.rx.cntReg[13] ;
 wire \e.rx.cntReg[14] ;
 wire \e.rx.cntReg[15] ;
 wire \e.rx.cntReg[16] ;
 wire \e.rx.cntReg[17] ;
 wire \e.rx.cntReg[18] ;
 wire \e.rx.cntReg[19] ;
 wire \e.rx.cntReg[1] ;
 wire \e.rx.cntReg[2] ;
 wire \e.rx.cntReg[3] ;
 wire \e.rx.cntReg[4] ;
 wire \e.rx.cntReg[5] ;
 wire \e.rx.cntReg[6] ;
 wire \e.rx.cntReg[7] ;
 wire \e.rx.cntReg[8] ;
 wire \e.rx.cntReg[9] ;
 wire \e.rx.rxReg ;
 wire \e.rx.rxReg_REG ;
 wire \e.tx._shiftReg_T_1[0] ;
 wire \e.tx._shiftReg_T_1[1] ;
 wire \e.tx._shiftReg_T_1[2] ;
 wire \e.tx._shiftReg_T_1[3] ;
 wire \e.tx._shiftReg_T_1[4] ;
 wire \e.tx._shiftReg_T_1[5] ;
 wire \e.tx._shiftReg_T_1[6] ;
 wire \e.tx._shiftReg_T_1[7] ;
 wire \e.tx.bitsReg[0] ;
 wire \e.tx.bitsReg[1] ;
 wire \e.tx.bitsReg[2] ;
 wire \e.tx.bitsReg[3] ;
 wire \e.tx.cntReg[0] ;
 wire \e.tx.cntReg[10] ;
 wire \e.tx.cntReg[11] ;
 wire \e.tx.cntReg[12] ;
 wire \e.tx.cntReg[13] ;
 wire \e.tx.cntReg[14] ;
 wire \e.tx.cntReg[15] ;
 wire \e.tx.cntReg[16] ;
 wire \e.tx.cntReg[17] ;
 wire \e.tx.cntReg[18] ;
 wire \e.tx.cntReg[19] ;
 wire \e.tx.cntReg[1] ;
 wire \e.tx.cntReg[2] ;
 wire \e.tx.cntReg[3] ;
 wire \e.tx.cntReg[4] ;
 wire \e.tx.cntReg[5] ;
 wire \e.tx.cntReg[6] ;
 wire \e.tx.cntReg[7] ;
 wire \e.tx.cntReg[8] ;
 wire \e.tx.cntReg[9] ;
 wire \e.updateKey ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;

 sg13g2_inv_1 _0500_ (.Y(_0093_),
    .A(net192));
 sg13g2_inv_1 _0501_ (.Y(_0094_),
    .A(net205));
 sg13g2_inv_1 _0502_ (.Y(_0095_),
    .A(net182));
 sg13g2_inv_1 _0503_ (.Y(_0096_),
    .A(net185));
 sg13g2_inv_1 _0504_ (.Y(_0097_),
    .A(net233));
 sg13g2_inv_1 _0505_ (.Y(_0098_),
    .A(\e.rx.cntReg[18] ));
 sg13g2_inv_1 _0506_ (.Y(_0099_),
    .A(net249));
 sg13g2_inv_1 _0507_ (.Y(_0100_),
    .A(\e.rx.cntReg[8] ));
 sg13g2_inv_1 _0508_ (.Y(_0101_),
    .A(net158));
 sg13g2_inv_1 _0509_ (.Y(_0102_),
    .A(net166));
 sg13g2_inv_1 _0510_ (.Y(_0103_),
    .A(net285));
 sg13g2_inv_1 _0511_ (.Y(_0104_),
    .A(net142));
 sg13g2_inv_1 _0512_ (.Y(_0105_),
    .A(net152));
 sg13g2_or2_1 _0513_ (.X(_0001_),
    .B(net2),
    .A(net116));
 sg13g2_or2_1 _0514_ (.X(_0000_),
    .B(net144),
    .A(net111));
 sg13g2_nor2_1 _0515_ (.A(net143),
    .B(net111),
    .Y(_0009_));
 sg13g2_or2_1 _0516_ (.X(_0106_),
    .B(net229),
    .A(net143));
 sg13g2_nand2_1 _0517_ (.Y(_0107_),
    .A(net143),
    .B(net229));
 sg13g2_a21oi_1 _0518_ (.A1(_0106_),
    .A2(_0107_),
    .Y(_0010_),
    .B1(net111));
 sg13g2_xor2_1 _0519_ (.B(_0106_),
    .A(net270),
    .X(_0108_));
 sg13g2_nor2_1 _0520_ (.A(net111),
    .B(_0108_),
    .Y(_0011_));
 sg13g2_nor4_2 _0521_ (.A(net143),
    .B(net229),
    .C(net224),
    .Y(_0109_),
    .D(\e.tx.cntReg[2] ));
 sg13g2_or3_1 _0522_ (.A(net224),
    .B(\e.tx.cntReg[2] ),
    .C(_0106_),
    .X(_0110_));
 sg13g2_xnor2_1 _0523_ (.Y(_0111_),
    .A(net230),
    .B(_0109_));
 sg13g2_nor2_1 _0524_ (.A(net111),
    .B(net231),
    .Y(_0012_));
 sg13g2_nor2_1 _0525_ (.A(net155),
    .B(\e.tx.cntReg[4] ),
    .Y(_0112_));
 sg13g2_nand2_1 _0526_ (.Y(_0113_),
    .A(_0109_),
    .B(_0112_));
 sg13g2_xor2_1 _0527_ (.B(_0113_),
    .A(net263),
    .X(_0114_));
 sg13g2_nor2_1 _0528_ (.A(net111),
    .B(_0114_),
    .Y(_0013_));
 sg13g2_nor2_1 _0529_ (.A(net164),
    .B(net295),
    .Y(_0115_));
 sg13g2_and3_1 _0530_ (.X(_0116_),
    .A(_0109_),
    .B(_0112_),
    .C(_0115_));
 sg13g2_nand3_1 _0531_ (.B(_0112_),
    .C(_0115_),
    .A(_0109_),
    .Y(_0117_));
 sg13g2_or2_1 _0532_ (.X(_0118_),
    .B(\e.tx.cntReg[8] ),
    .A(net293));
 sg13g2_nor2_1 _0533_ (.A(\e.tx.cntReg[8] ),
    .B(net104),
    .Y(_0119_));
 sg13g2_nor3_1 _0534_ (.A(_0105_),
    .B(net104),
    .C(net294),
    .Y(_0120_));
 sg13g2_o21ai_1 _0535_ (.B1(_0105_),
    .Y(_0121_),
    .A1(net104),
    .A2(_0118_));
 sg13g2_nor4_1 _0536_ (.A(\e.tx.cntReg[9] ),
    .B(\e.tx.cntReg[8] ),
    .C(\e.tx.cntReg[11] ),
    .D(\e.tx.cntReg[10] ),
    .Y(_0122_));
 sg13g2_or3_1 _0537_ (.A(\e.tx.cntReg[11] ),
    .B(\e.tx.cntReg[10] ),
    .C(_0118_),
    .X(_0123_));
 sg13g2_nor4_1 _0538_ (.A(\e.tx.cntReg[13] ),
    .B(\e.tx.cntReg[12] ),
    .C(\e.tx.cntReg[14] ),
    .D(\e.tx.cntReg[15] ),
    .Y(_0124_));
 sg13g2_and2_1 _0539_ (.A(_0122_),
    .B(_0124_),
    .X(_0125_));
 sg13g2_nand2_1 _0540_ (.Y(_0126_),
    .A(_0122_),
    .B(_0124_));
 sg13g2_nor4_2 _0541_ (.A(\e.tx.cntReg[16] ),
    .B(\e.tx.cntReg[17] ),
    .C(\e.tx.cntReg[18] ),
    .Y(_0127_),
    .D(\e.tx.cntReg[19] ));
 sg13g2_and3_2 _0542_ (.X(_0128_),
    .A(_0116_),
    .B(_0125_),
    .C(_0127_));
 sg13g2_nand3_1 _0543_ (.B(_0125_),
    .C(_0127_),
    .A(_0116_),
    .Y(_0129_));
 sg13g2_nor2_1 _0544_ (.A(_0120_),
    .B(_0128_),
    .Y(_0130_));
 sg13g2_a21oi_1 _0545_ (.A1(_0121_),
    .A2(_0130_),
    .Y(_0014_),
    .B1(net109));
 sg13g2_nor3_1 _0546_ (.A(net288),
    .B(_0117_),
    .C(_0123_),
    .Y(_0131_));
 sg13g2_o21ai_1 _0547_ (.B1(net288),
    .Y(_0132_),
    .A1(_0117_),
    .A2(_0123_));
 sg13g2_nor2b_1 _0548_ (.A(net289),
    .B_N(_0132_),
    .Y(_0133_));
 sg13g2_nor2_1 _0549_ (.A(net109),
    .B(_0133_),
    .Y(_0015_));
 sg13g2_nor2_1 _0550_ (.A(net109),
    .B(_0128_),
    .Y(_0134_));
 sg13g2_nand2b_1 _0551_ (.Y(_0135_),
    .B(net99),
    .A_N(net109));
 sg13g2_o21ai_1 _0552_ (.B1(net224),
    .Y(_0136_),
    .A1(\e.tx.cntReg[2] ),
    .A2(_0106_));
 sg13g2_a21oi_1 _0553_ (.A1(_0110_),
    .A2(net225),
    .Y(_0016_),
    .B1(net92));
 sg13g2_o21ai_1 _0554_ (.B1(net155),
    .Y(_0137_),
    .A1(\e.tx.cntReg[4] ),
    .A2(_0110_));
 sg13g2_a21oi_1 _0555_ (.A1(_0113_),
    .A2(net156),
    .Y(_0017_),
    .B1(net92));
 sg13g2_o21ai_1 _0556_ (.B1(net164),
    .Y(_0138_),
    .A1(\e.tx.cntReg[6] ),
    .A2(_0113_));
 sg13g2_a21oi_1 _0557_ (.A1(net104),
    .A2(net165),
    .Y(_0018_),
    .B1(net92));
 sg13g2_xnor2_1 _0558_ (.Y(_0139_),
    .A(net260),
    .B(_0116_));
 sg13g2_nor2_1 _0559_ (.A(net93),
    .B(_0139_),
    .Y(_0019_));
 sg13g2_xnor2_1 _0560_ (.Y(_0140_),
    .A(net247),
    .B(_0119_));
 sg13g2_nor2_1 _0561_ (.A(net92),
    .B(net248),
    .Y(_0020_));
 sg13g2_nor2_1 _0562_ (.A(net232),
    .B(_0120_),
    .Y(_0141_));
 sg13g2_and2_1 _0563_ (.A(net232),
    .B(_0120_),
    .X(_0142_));
 sg13g2_nor3_1 _0564_ (.A(net93),
    .B(_0141_),
    .C(_0142_),
    .Y(_0021_));
 sg13g2_nor4_2 _0565_ (.A(\e.tx.cntReg[13] ),
    .B(\e.tx.cntReg[12] ),
    .C(net104),
    .Y(_0143_),
    .D(_0123_));
 sg13g2_xnor2_1 _0566_ (.Y(_0144_),
    .A(net261),
    .B(_0131_));
 sg13g2_nor2_1 _0567_ (.A(net93),
    .B(net262),
    .Y(_0022_));
 sg13g2_xor2_1 _0568_ (.B(_0143_),
    .A(net210),
    .X(_0145_));
 sg13g2_nor2_1 _0569_ (.A(net93),
    .B(net211),
    .Y(_0023_));
 sg13g2_a21oi_1 _0570_ (.A1(_0007_),
    .A2(_0143_),
    .Y(_0146_),
    .B1(net149));
 sg13g2_and3_1 _0571_ (.X(_0147_),
    .A(net149),
    .B(_0007_),
    .C(_0143_));
 sg13g2_nor3_1 _0572_ (.A(net93),
    .B(net150),
    .C(_0147_),
    .Y(_0024_));
 sg13g2_nor3_1 _0573_ (.A(net290),
    .B(net104),
    .C(_0126_),
    .Y(_0148_));
 sg13g2_o21ai_1 _0574_ (.B1(net290),
    .Y(_0149_),
    .A1(net104),
    .A2(_0126_));
 sg13g2_nor2b_1 _0575_ (.A(net291),
    .B_N(_0149_),
    .Y(_0150_));
 sg13g2_nor2_1 _0576_ (.A(net92),
    .B(_0150_),
    .Y(_0025_));
 sg13g2_nor4_2 _0577_ (.A(\e.tx.cntReg[16] ),
    .B(\e.tx.cntReg[17] ),
    .C(net104),
    .Y(_0151_),
    .D(_0126_));
 sg13g2_xnor2_1 _0578_ (.Y(_0152_),
    .A(net276),
    .B(_0148_));
 sg13g2_nor2_1 _0579_ (.A(net92),
    .B(net277),
    .Y(_0026_));
 sg13g2_xor2_1 _0580_ (.B(_0151_),
    .A(net221),
    .X(_0153_));
 sg13g2_nor2_1 _0581_ (.A(net92),
    .B(net222),
    .Y(_0027_));
 sg13g2_a21oi_1 _0582_ (.A1(_0008_),
    .A2(_0151_),
    .Y(_0154_),
    .B1(net179));
 sg13g2_and3_1 _0583_ (.X(_0155_),
    .A(net179),
    .B(_0008_),
    .C(_0151_));
 sg13g2_nor3_1 _0584_ (.A(net92),
    .B(net180),
    .C(_0155_),
    .Y(_0028_));
 sg13g2_nor2_1 _0585_ (.A(net252),
    .B(\e.tx.bitsReg[0] ),
    .Y(_0156_));
 sg13g2_or2_1 _0586_ (.X(_0157_),
    .B(\e.tx.bitsReg[0] ),
    .A(\e.tx.bitsReg[1] ));
 sg13g2_nor3_2 _0587_ (.A(net170),
    .B(\e.tx.bitsReg[1] ),
    .C(\e.tx.bitsReg[0] ),
    .Y(_0158_));
 sg13g2_inv_1 _0588_ (.Y(_0159_),
    .A(_0158_));
 sg13g2_nor2b_1 _0589_ (.A(net206),
    .B_N(_0158_),
    .Y(_0160_));
 sg13g2_nand2b_1 _0590_ (.Y(_0161_),
    .B(_0158_),
    .A_N(\e.tx.bitsReg[3] ));
 sg13g2_nand2_2 _0591_ (.Y(_0162_),
    .A(net108),
    .B(net103));
 sg13g2_and2_1 _0592_ (.A(_0128_),
    .B(_0162_),
    .X(_0163_));
 sg13g2_a21oi_1 _0593_ (.A1(\e.tx._shiftReg_T_1[0] ),
    .A2(_0161_),
    .Y(_0164_),
    .B1(net110));
 sg13g2_a22oi_1 _0594_ (.Y(_0029_),
    .B1(_0163_),
    .B2(_0164_),
    .A2(_0134_),
    .A1(_0102_));
 sg13g2_nand2b_1 _0595_ (.Y(_0165_),
    .B(net185),
    .A_N(\e.buf_.dataReg[0] ));
 sg13g2_a21oi_1 _0596_ (.A1(_0096_),
    .A2(\e.buf_.dataReg[0] ),
    .Y(_0166_),
    .B1(net108));
 sg13g2_nand3_1 _0597_ (.B(_0165_),
    .C(_0166_),
    .A(net103),
    .Y(_0167_));
 sg13g2_o21ai_1 _0598_ (.B1(_0167_),
    .Y(_0168_),
    .A1(\e.tx._shiftReg_T_1[1] ),
    .A2(net103));
 sg13g2_a21oi_1 _0599_ (.A1(net214),
    .A2(net99),
    .Y(_0169_),
    .B1(net109));
 sg13g2_o21ai_1 _0600_ (.B1(_0169_),
    .Y(_0030_),
    .A1(net99),
    .A2(_0168_));
 sg13g2_xnor2_1 _0601_ (.Y(_0170_),
    .A(\e.key[1] ),
    .B(\e.buf_.dataReg[1] ));
 sg13g2_nand3b_1 _0602_ (.B(net102),
    .C(_0170_),
    .Y(_0171_),
    .A_N(_0002_));
 sg13g2_o21ai_1 _0603_ (.B1(_0171_),
    .Y(_0172_),
    .A1(net208),
    .A2(net102));
 sg13g2_a21oi_1 _0604_ (.A1(net227),
    .A2(net97),
    .Y(_0173_),
    .B1(net116));
 sg13g2_o21ai_1 _0605_ (.B1(_0173_),
    .Y(_0031_),
    .A1(net97),
    .A2(_0172_));
 sg13g2_nand2b_1 _0606_ (.Y(_0174_),
    .B(net182),
    .A_N(\e.buf_.dataReg[2] ));
 sg13g2_a21oi_1 _0607_ (.A1(_0095_),
    .A2(\e.buf_.dataReg[2] ),
    .Y(_0175_),
    .B1(net108));
 sg13g2_nand3_1 _0608_ (.B(_0174_),
    .C(_0175_),
    .A(net102),
    .Y(_0176_));
 sg13g2_o21ai_1 _0609_ (.B1(_0176_),
    .Y(_0177_),
    .A1(\e.tx._shiftReg_T_1[3] ),
    .A2(_0160_));
 sg13g2_a21oi_1 _0610_ (.A1(net208),
    .A2(net98),
    .Y(_0178_),
    .B1(net118));
 sg13g2_o21ai_1 _0611_ (.B1(_0178_),
    .Y(_0032_),
    .A1(net98),
    .A2(_0177_));
 sg13g2_xnor2_1 _0612_ (.Y(_0179_),
    .A(\e.key[3] ),
    .B(\e.buf_.dataReg[3] ));
 sg13g2_nand3b_1 _0613_ (.B(net102),
    .C(_0179_),
    .Y(_0180_),
    .A_N(net108));
 sg13g2_o21ai_1 _0614_ (.B1(_0180_),
    .Y(_0181_),
    .A1(net213),
    .A2(net103));
 sg13g2_a21oi_1 _0615_ (.A1(net223),
    .A2(net98),
    .Y(_0182_),
    .B1(net118));
 sg13g2_o21ai_1 _0616_ (.B1(_0182_),
    .Y(_0033_),
    .A1(net98),
    .A2(_0181_));
 sg13g2_nand2b_1 _0617_ (.Y(_0183_),
    .B(net205),
    .A_N(\e.buf_.dataReg[4] ));
 sg13g2_a21oi_1 _0618_ (.A1(_0094_),
    .A2(\e.buf_.dataReg[4] ),
    .Y(_0184_),
    .B1(net108));
 sg13g2_nand3_1 _0619_ (.B(_0183_),
    .C(_0184_),
    .A(net102),
    .Y(_0185_));
 sg13g2_o21ai_1 _0620_ (.B1(_0185_),
    .Y(_0186_),
    .A1(net200),
    .A2(net102));
 sg13g2_a21oi_1 _0621_ (.A1(net213),
    .A2(net97),
    .Y(_0187_),
    .B1(net118));
 sg13g2_o21ai_1 _0622_ (.B1(_0187_),
    .Y(_0034_),
    .A1(net98),
    .A2(_0186_));
 sg13g2_xnor2_1 _0623_ (.Y(_0188_),
    .A(\e.key[5] ),
    .B(\e.buf_.dataReg[5] ));
 sg13g2_nand3b_1 _0624_ (.B(net102),
    .C(_0188_),
    .Y(_0189_),
    .A_N(net108));
 sg13g2_o21ai_1 _0625_ (.B1(_0189_),
    .Y(_0190_),
    .A1(\e.tx._shiftReg_T_1[6] ),
    .A2(net102));
 sg13g2_a21oi_1 _0626_ (.A1(net200),
    .A2(net97),
    .Y(_0191_),
    .B1(net118));
 sg13g2_o21ai_1 _0627_ (.B1(_0191_),
    .Y(_0035_),
    .A1(net97),
    .A2(_0190_));
 sg13g2_nand2b_1 _0628_ (.Y(_0192_),
    .B(net192),
    .A_N(\e.buf_.dataReg[6] ));
 sg13g2_a21oi_1 _0629_ (.A1(_0093_),
    .A2(\e.buf_.dataReg[6] ),
    .Y(_0193_),
    .B1(net108));
 sg13g2_nand3_1 _0630_ (.B(_0192_),
    .C(_0193_),
    .A(net103),
    .Y(_0194_));
 sg13g2_o21ai_1 _0631_ (.B1(_0194_),
    .Y(_0195_),
    .A1(net158),
    .A2(net103));
 sg13g2_a21oi_1 _0632_ (.A1(net202),
    .A2(net97),
    .Y(_0196_),
    .B1(net116));
 sg13g2_o21ai_1 _0633_ (.B1(_0196_),
    .Y(_0036_),
    .A1(net97),
    .A2(_0195_));
 sg13g2_nor2_1 _0634_ (.A(net99),
    .B(_0161_),
    .Y(_0197_));
 sg13g2_xor2_1 _0635_ (.B(\e.buf_.dataReg[7] ),
    .A(\e.key[7] ),
    .X(_0198_));
 sg13g2_nor3_1 _0636_ (.A(_0103_),
    .B(net115),
    .C(_0198_),
    .Y(_0199_));
 sg13g2_a22oi_1 _0637_ (.Y(_0037_),
    .B1(_0197_),
    .B2(_0199_),
    .A2(_0134_),
    .A1(_0101_));
 sg13g2_nor2b_1 _0638_ (.A(net108),
    .B_N(net268),
    .Y(_0200_));
 sg13g2_nor2_1 _0639_ (.A(net268),
    .B(net1),
    .Y(_0201_));
 sg13g2_nor3_1 _0640_ (.A(net116),
    .B(_0200_),
    .C(_0201_),
    .Y(_0038_));
 sg13g2_nor2b_1 _0641_ (.A(\e.buf_.io_out_valid ),
    .B_N(net145),
    .Y(_0202_));
 sg13g2_nand2_1 _0642_ (.Y(_0203_),
    .A(net145),
    .B(_0103_));
 sg13g2_nor2_1 _0643_ (.A(net153),
    .B(net101),
    .Y(_0204_));
 sg13g2_nor2_1 _0644_ (.A(net184),
    .B(net107),
    .Y(_0205_));
 sg13g2_nor3_1 _0645_ (.A(net110),
    .B(_0204_),
    .C(_0205_),
    .Y(_0039_));
 sg13g2_nor2_1 _0646_ (.A(\e.buf_.io_in_bits[1] ),
    .B(net101),
    .Y(_0206_));
 sg13g2_nor2_1 _0647_ (.A(net241),
    .B(_0202_),
    .Y(_0207_));
 sg13g2_nor3_1 _0648_ (.A(net115),
    .B(_0206_),
    .C(net242),
    .Y(_0040_));
 sg13g2_nor2_1 _0649_ (.A(net194),
    .B(_0203_),
    .Y(_0208_));
 sg13g2_nor2_1 _0650_ (.A(net244),
    .B(net107),
    .Y(_0209_));
 sg13g2_nor3_1 _0651_ (.A(net117),
    .B(_0208_),
    .C(_0209_),
    .Y(_0041_));
 sg13g2_nor2_1 _0652_ (.A(net190),
    .B(net101),
    .Y(_0210_));
 sg13g2_nor2_1 _0653_ (.A(net197),
    .B(net107),
    .Y(_0211_));
 sg13g2_nor3_1 _0654_ (.A(net117),
    .B(_0210_),
    .C(_0211_),
    .Y(_0042_));
 sg13g2_nor2_1 _0655_ (.A(net173),
    .B(net101),
    .Y(_0212_));
 sg13g2_nor2_1 _0656_ (.A(net196),
    .B(net107),
    .Y(_0213_));
 sg13g2_nor3_1 _0657_ (.A(net117),
    .B(_0212_),
    .C(_0213_),
    .Y(_0043_));
 sg13g2_nor2_1 _0658_ (.A(net177),
    .B(net101),
    .Y(_0214_));
 sg13g2_nor2_1 _0659_ (.A(net178),
    .B(net107),
    .Y(_0215_));
 sg13g2_nor3_1 _0660_ (.A(net117),
    .B(_0214_),
    .C(_0215_),
    .Y(_0044_));
 sg13g2_nor2_1 _0661_ (.A(net168),
    .B(net101),
    .Y(_0216_));
 sg13g2_nor2_1 _0662_ (.A(net212),
    .B(net107),
    .Y(_0217_));
 sg13g2_nor3_1 _0663_ (.A(net115),
    .B(_0216_),
    .C(_0217_),
    .Y(_0045_));
 sg13g2_nor2_1 _0664_ (.A(net203),
    .B(net101),
    .Y(_0218_));
 sg13g2_nor2_1 _0665_ (.A(net234),
    .B(net107),
    .Y(_0219_));
 sg13g2_nor3_1 _0666_ (.A(net115),
    .B(_0218_),
    .C(_0219_),
    .Y(_0046_));
 sg13g2_nor2_1 _0667_ (.A(net292),
    .B(\e.rx.cntReg[0] ),
    .Y(_0220_));
 sg13g2_or2_1 _0668_ (.X(_0221_),
    .B(\e.rx.cntReg[0] ),
    .A(net264));
 sg13g2_nor4_2 _0669_ (.A(net238),
    .B(net245),
    .C(net264),
    .Y(_0222_),
    .D(\e.rx.cntReg[0] ));
 sg13g2_or4_2 _0670_ (.A(net238),
    .B(\e.rx.cntReg[2] ),
    .C(\e.rx.cntReg[1] ),
    .D(\e.rx.cntReg[0] ),
    .X(_0223_));
 sg13g2_nor4_2 _0671_ (.A(\e.rx.cntReg[7] ),
    .B(net296),
    .C(\e.rx.cntReg[5] ),
    .Y(_0224_),
    .D(\e.rx.cntReg[4] ));
 sg13g2_and2_1 _0672_ (.A(_0222_),
    .B(_0224_),
    .X(_0225_));
 sg13g2_nand2_2 _0673_ (.Y(_0226_),
    .A(_0222_),
    .B(_0224_));
 sg13g2_nor2_1 _0674_ (.A(\e.rx.cntReg[11] ),
    .B(\e.rx.cntReg[10] ),
    .Y(_0227_));
 sg13g2_nor3_2 _0675_ (.A(\e.rx.cntReg[12] ),
    .B(\e.rx.cntReg[9] ),
    .C(\e.rx.cntReg[8] ),
    .Y(_0228_));
 sg13g2_nand2_1 _0676_ (.Y(_0229_),
    .A(_0227_),
    .B(_0228_));
 sg13g2_nor3_1 _0677_ (.A(\e.rx.cntReg[15] ),
    .B(\e.rx.cntReg[14] ),
    .C(\e.rx.cntReg[13] ),
    .Y(_0230_));
 sg13g2_and3_1 _0678_ (.X(_0231_),
    .A(_0227_),
    .B(_0228_),
    .C(_0230_));
 sg13g2_nand3_1 _0679_ (.B(_0228_),
    .C(_0230_),
    .A(_0227_),
    .Y(_0232_));
 sg13g2_nor2_1 _0680_ (.A(net100),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_nor4_2 _0681_ (.A(\e.rx.cntReg[19] ),
    .B(\e.rx.cntReg[18] ),
    .C(\e.rx.cntReg[17] ),
    .Y(_0234_),
    .D(\e.rx.cntReg[16] ));
 sg13g2_or4_2 _0682_ (.A(\e.rx.cntReg[19] ),
    .B(\e.rx.cntReg[18] ),
    .C(\e.rx.cntReg[17] ),
    .D(\e.rx.cntReg[16] ),
    .X(_0235_));
 sg13g2_nor3_2 _0683_ (.A(_0226_),
    .B(_0232_),
    .C(_0235_),
    .Y(_0236_));
 sg13g2_nand3_1 _0684_ (.B(_0231_),
    .C(_0234_),
    .A(_0225_),
    .Y(_0237_));
 sg13g2_nor2_1 _0685_ (.A(\e.rx.bitsReg[1] ),
    .B(\e.rx.bitsReg[0] ),
    .Y(_0238_));
 sg13g2_nand2b_1 _0686_ (.Y(_0239_),
    .B(_0238_),
    .A_N(net218));
 sg13g2_nor4_2 _0687_ (.A(net257),
    .B(net218),
    .C(net237),
    .Y(_0240_),
    .D(net233));
 sg13g2_nor4_1 _0688_ (.A(net100),
    .B(_0232_),
    .C(_0235_),
    .D(_0240_),
    .Y(_0241_));
 sg13g2_nor2b_1 _0689_ (.A(\e.buf_.io_in_bits[1] ),
    .B_N(net96),
    .Y(_0242_));
 sg13g2_nor2_1 _0690_ (.A(net153),
    .B(net96),
    .Y(_0243_));
 sg13g2_nor3_1 _0691_ (.A(net113),
    .B(_0242_),
    .C(_0243_),
    .Y(_0047_));
 sg13g2_nor2b_1 _0692_ (.A(net194),
    .B_N(net94),
    .Y(_0244_));
 sg13g2_nor2_1 _0693_ (.A(\e.buf_.io_in_bits[1] ),
    .B(net94),
    .Y(_0245_));
 sg13g2_nor3_1 _0694_ (.A(net114),
    .B(_0244_),
    .C(_0245_),
    .Y(_0048_));
 sg13g2_nor2b_1 _0695_ (.A(net190),
    .B_N(net94),
    .Y(_0246_));
 sg13g2_nor2_1 _0696_ (.A(\e.buf_.io_in_bits[2] ),
    .B(net94),
    .Y(_0247_));
 sg13g2_nor3_1 _0697_ (.A(net114),
    .B(_0246_),
    .C(_0247_),
    .Y(_0049_));
 sg13g2_nor2b_1 _0698_ (.A(net173),
    .B_N(net94),
    .Y(_0248_));
 sg13g2_nor2_1 _0699_ (.A(\e.buf_.io_in_bits[3] ),
    .B(net95),
    .Y(_0249_));
 sg13g2_nor3_1 _0700_ (.A(net114),
    .B(_0248_),
    .C(_0249_),
    .Y(_0050_));
 sg13g2_nor2b_1 _0701_ (.A(net177),
    .B_N(net94),
    .Y(_0250_));
 sg13g2_nor2_1 _0702_ (.A(net173),
    .B(net94),
    .Y(_0251_));
 sg13g2_nor3_1 _0703_ (.A(net114),
    .B(_0250_),
    .C(_0251_),
    .Y(_0051_));
 sg13g2_nor2b_1 _0704_ (.A(net168),
    .B_N(net96),
    .Y(_0252_));
 sg13g2_nor2_1 _0705_ (.A(net177),
    .B(net94),
    .Y(_0253_));
 sg13g2_nor3_1 _0706_ (.A(net113),
    .B(_0252_),
    .C(_0253_),
    .Y(_0052_));
 sg13g2_nor2b_1 _0707_ (.A(\e.buf_.io_in_bits[7] ),
    .B_N(net96),
    .Y(_0254_));
 sg13g2_nor2_1 _0708_ (.A(net168),
    .B(net96),
    .Y(_0255_));
 sg13g2_nor3_1 _0709_ (.A(net113),
    .B(_0254_),
    .C(_0255_),
    .Y(_0053_));
 sg13g2_nor2b_1 _0710_ (.A(\e.rx.rxReg ),
    .B_N(net96),
    .Y(_0256_));
 sg13g2_nor2_1 _0711_ (.A(net203),
    .B(net96),
    .Y(_0257_));
 sg13g2_nor3_1 _0712_ (.A(net111),
    .B(_0256_),
    .C(_0257_),
    .Y(_0054_));
 sg13g2_a21o_1 _0713_ (.A2(_0240_),
    .A1(_0236_),
    .B1(net112),
    .X(_0258_));
 sg13g2_a21oi_1 _0714_ (.A1(_0104_),
    .A2(_0237_),
    .Y(_0055_),
    .B1(_0258_));
 sg13g2_nand2_1 _0715_ (.Y(_0259_),
    .A(net264),
    .B(\e.rx.cntReg[0] ));
 sg13g2_a21oi_1 _0716_ (.A1(_0221_),
    .A2(net265),
    .Y(_0056_),
    .B1(_0258_));
 sg13g2_and2_1 _0717_ (.A(\e.rx.rxReg ),
    .B(_0240_),
    .X(_0260_));
 sg13g2_nand2_1 _0718_ (.Y(_0261_),
    .A(\e.rx.rxReg ),
    .B(_0240_));
 sg13g2_nor4_1 _0719_ (.A(net100),
    .B(_0232_),
    .C(_0235_),
    .D(_0261_),
    .Y(_0262_));
 sg13g2_nand4_1 _0720_ (.B(_0231_),
    .C(_0234_),
    .A(_0225_),
    .Y(_0263_),
    .D(_0260_));
 sg13g2_and3_1 _0721_ (.X(_0264_),
    .A(net245),
    .B(_0220_),
    .C(_0263_));
 sg13g2_a21oi_1 _0722_ (.A1(_0220_),
    .A2(_0263_),
    .Y(_0265_),
    .B1(net245));
 sg13g2_nor3_1 _0723_ (.A(net114),
    .B(_0264_),
    .C(net246),
    .Y(_0057_));
 sg13g2_nand2b_1 _0724_ (.Y(_0266_),
    .B(_0237_),
    .A_N(net112));
 sg13g2_o21ai_1 _0725_ (.B1(net238),
    .Y(_0267_),
    .A1(\e.rx.cntReg[2] ),
    .A2(_0221_));
 sg13g2_a21oi_1 _0726_ (.A1(_0223_),
    .A2(net239),
    .Y(_0058_),
    .B1(_0266_));
 sg13g2_xnor2_1 _0727_ (.Y(_0268_),
    .A(net278),
    .B(_0222_));
 sg13g2_nor2_1 _0728_ (.A(_0258_),
    .B(net279),
    .Y(_0059_));
 sg13g2_nor3_2 _0729_ (.A(net286),
    .B(net278),
    .C(_0223_),
    .Y(_0269_));
 sg13g2_o21ai_1 _0730_ (.B1(net286),
    .Y(_0270_),
    .A1(net278),
    .A2(_0223_));
 sg13g2_nor2b_1 _0731_ (.A(net287),
    .B_N(_0270_),
    .Y(_0271_));
 sg13g2_nor2_1 _0732_ (.A(net91),
    .B(_0271_),
    .Y(_0060_));
 sg13g2_nand2_1 _0733_ (.Y(_0272_),
    .A(net255),
    .B(_0269_));
 sg13g2_xor2_1 _0734_ (.B(_0269_),
    .A(net255),
    .X(_0273_));
 sg13g2_a21oi_1 _0735_ (.A1(_0237_),
    .A2(net256),
    .Y(_0061_),
    .B1(_0258_));
 sg13g2_or3_1 _0736_ (.A(net112),
    .B(net96),
    .C(_0262_),
    .X(_0274_));
 sg13g2_xor2_1 _0737_ (.B(_0272_),
    .A(net282),
    .X(_0275_));
 sg13g2_a21oi_1 _0738_ (.A1(_0237_),
    .A2(_0275_),
    .Y(_0062_),
    .B1(_0274_));
 sg13g2_xnor2_1 _0739_ (.Y(_0276_),
    .A(net275),
    .B(_0225_));
 sg13g2_nor2_1 _0740_ (.A(net91),
    .B(_0276_),
    .Y(_0063_));
 sg13g2_and4_1 _0741_ (.A(_0099_),
    .B(_0100_),
    .C(_0222_),
    .D(_0224_),
    .X(_0277_));
 sg13g2_nand3_1 _0742_ (.B(_0100_),
    .C(_0225_),
    .A(_0099_),
    .Y(_0278_));
 sg13g2_o21ai_1 _0743_ (.B1(net249),
    .Y(_0279_),
    .A1(\e.rx.cntReg[8] ),
    .A2(_0226_));
 sg13g2_a21oi_1 _0744_ (.A1(_0278_),
    .A2(net250),
    .Y(_0064_),
    .B1(_0274_));
 sg13g2_nand2_1 _0745_ (.Y(_0280_),
    .A(net162),
    .B(_0277_));
 sg13g2_nor2_1 _0746_ (.A(net162),
    .B(_0277_),
    .Y(_0281_));
 sg13g2_nor2_1 _0747_ (.A(_0236_),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_a221oi_1 _0748_ (.B2(_0282_),
    .C1(net112),
    .B1(_0280_),
    .A1(_0236_),
    .Y(_0065_),
    .A2(_0260_));
 sg13g2_xor2_1 _0749_ (.B(_0280_),
    .A(net280),
    .X(_0283_));
 sg13g2_a21oi_1 _0750_ (.A1(_0237_),
    .A2(_0283_),
    .Y(_0066_),
    .B1(_0274_));
 sg13g2_and2_1 _0751_ (.A(_0227_),
    .B(_0277_),
    .X(_0284_));
 sg13g2_and3_1 _0752_ (.X(_0285_),
    .A(net160),
    .B(_0263_),
    .C(_0284_));
 sg13g2_a21oi_1 _0753_ (.A1(_0263_),
    .A2(_0284_),
    .Y(_0286_),
    .B1(net160));
 sg13g2_nor3_1 _0754_ (.A(net112),
    .B(_0285_),
    .C(net161),
    .Y(_0067_));
 sg13g2_nor3_1 _0755_ (.A(net283),
    .B(net100),
    .C(_0229_),
    .Y(_0287_));
 sg13g2_o21ai_1 _0756_ (.B1(net283),
    .Y(_0288_),
    .A1(net100),
    .A2(_0229_));
 sg13g2_nor2b_1 _0757_ (.A(net284),
    .B_N(_0288_),
    .Y(_0289_));
 sg13g2_nor2_1 _0758_ (.A(net91),
    .B(_0289_),
    .Y(_0068_));
 sg13g2_or4_1 _0759_ (.A(\e.rx.cntReg[14] ),
    .B(\e.rx.cntReg[13] ),
    .C(net100),
    .D(_0229_),
    .X(_0290_));
 sg13g2_xnor2_1 _0760_ (.Y(_0291_),
    .A(net235),
    .B(_0287_));
 sg13g2_nor2_1 _0761_ (.A(net91),
    .B(net236),
    .Y(_0069_));
 sg13g2_a21oi_1 _0762_ (.A1(net175),
    .A2(_0290_),
    .Y(_0292_),
    .B1(_0233_));
 sg13g2_nor2_1 _0763_ (.A(net91),
    .B(net176),
    .Y(_0070_));
 sg13g2_nor3_1 _0764_ (.A(\e.rx.cntReg[16] ),
    .B(net100),
    .C(_0232_),
    .Y(_0293_));
 sg13g2_xnor2_1 _0765_ (.Y(_0294_),
    .A(net281),
    .B(_0233_));
 sg13g2_nor2_1 _0766_ (.A(net91),
    .B(_0294_),
    .Y(_0071_));
 sg13g2_nor4_2 _0767_ (.A(\e.rx.cntReg[17] ),
    .B(\e.rx.cntReg[16] ),
    .C(net100),
    .Y(_0295_),
    .D(_0232_));
 sg13g2_xnor2_1 _0768_ (.Y(_0296_),
    .A(net273),
    .B(_0293_));
 sg13g2_nor2_1 _0769_ (.A(net91),
    .B(net274),
    .Y(_0072_));
 sg13g2_xnor2_1 _0770_ (.Y(_0297_),
    .A(net271),
    .B(_0295_));
 sg13g2_nor2_1 _0771_ (.A(net91),
    .B(net272),
    .Y(_0073_));
 sg13g2_nand2b_1 _0772_ (.Y(_0298_),
    .B(net147),
    .A_N(net111));
 sg13g2_a21oi_1 _0773_ (.A1(_0098_),
    .A2(_0295_),
    .Y(_0074_),
    .B1(_0298_));
 sg13g2_nand2_1 _0774_ (.Y(_0299_),
    .A(_0097_),
    .B(net95));
 sg13g2_nor4_1 _0775_ (.A(_0226_),
    .B(_0232_),
    .C(_0235_),
    .D(_0260_),
    .Y(_0300_));
 sg13g2_nand2_1 _0776_ (.Y(_0301_),
    .A(net233),
    .B(_0237_));
 sg13g2_a21oi_1 _0777_ (.A1(_0299_),
    .A2(_0301_),
    .Y(_0075_),
    .B1(net112));
 sg13g2_a21oi_1 _0778_ (.A1(_0097_),
    .A2(net95),
    .Y(_0302_),
    .B1(net237));
 sg13g2_and3_1 _0779_ (.X(_0303_),
    .A(net237),
    .B(_0097_),
    .C(net95));
 sg13g2_nor3_1 _0780_ (.A(net114),
    .B(_0302_),
    .C(_0303_),
    .Y(_0076_));
 sg13g2_nand2b_1 _0781_ (.Y(_0304_),
    .B(\e.rx.bitsReg[3] ),
    .A_N(\e.rx.bitsReg[2] ));
 sg13g2_and3_1 _0782_ (.X(_0305_),
    .A(_0238_),
    .B(_0300_),
    .C(_0304_));
 sg13g2_a21oi_1 _0783_ (.A1(_0238_),
    .A2(_0300_),
    .Y(_0306_),
    .B1(net218));
 sg13g2_nor3_1 _0784_ (.A(net112),
    .B(_0305_),
    .C(net219),
    .Y(_0077_));
 sg13g2_o21ai_1 _0785_ (.B1(net257),
    .Y(_0307_),
    .A1(_0237_),
    .A2(_0239_));
 sg13g2_nand3_1 _0786_ (.B(_0240_),
    .C(_0261_),
    .A(_0236_),
    .Y(_0308_));
 sg13g2_a21oi_1 _0787_ (.A1(net258),
    .A2(_0308_),
    .Y(_0078_),
    .B1(net112));
 sg13g2_nor4_1 _0788_ (.A(\e.rx.bitsReg[3] ),
    .B(\e.rx.bitsReg[2] ),
    .C(\e.rx.bitsReg[1] ),
    .D(_0097_),
    .Y(_0309_));
 sg13g2_a21oi_1 _0789_ (.A1(_0236_),
    .A2(_0309_),
    .Y(_0310_),
    .B1(net145));
 sg13g2_nor3_1 _0790_ (.A(net113),
    .B(net107),
    .C(net146),
    .Y(_0079_));
 sg13g2_nor2_1 _0791_ (.A(_0103_),
    .B(net268),
    .Y(_0311_));
 sg13g2_o21ai_1 _0792_ (.B1(_0311_),
    .Y(_0312_),
    .A1(net97),
    .A2(_0161_));
 sg13g2_a21oi_1 _0793_ (.A1(net101),
    .A2(_0312_),
    .Y(_0080_),
    .B1(net115));
 sg13g2_nand2_1 _0794_ (.Y(_0313_),
    .A(net267),
    .B(net99));
 sg13g2_nand3b_1 _0795_ (.B(_0128_),
    .C(_0162_),
    .Y(_0314_),
    .A_N(net267));
 sg13g2_a21oi_1 _0796_ (.A1(_0313_),
    .A2(_0314_),
    .Y(_0081_),
    .B1(net109));
 sg13g2_o21ai_1 _0797_ (.B1(net252),
    .Y(_0315_),
    .A1(\e.tx.bitsReg[0] ),
    .A2(net99));
 sg13g2_nand3_1 _0798_ (.B(_0156_),
    .C(_0162_),
    .A(_0128_),
    .Y(_0316_));
 sg13g2_a21oi_1 _0799_ (.A1(net253),
    .A2(_0316_),
    .Y(_0082_),
    .B1(net109));
 sg13g2_o21ai_1 _0800_ (.B1(net170),
    .Y(_0317_),
    .A1(net99),
    .A2(_0157_));
 sg13g2_nand3_1 _0801_ (.B(_0128_),
    .C(_0158_),
    .A(\e.tx.bitsReg[3] ),
    .Y(_0318_));
 sg13g2_a21oi_1 _0802_ (.A1(net171),
    .A2(_0318_),
    .Y(_0083_),
    .B1(net109));
 sg13g2_o21ai_1 _0803_ (.B1(net206),
    .Y(_0319_),
    .A1(net99),
    .A2(_0159_));
 sg13g2_nand3_1 _0804_ (.B(net103),
    .C(_0162_),
    .A(_0128_),
    .Y(_0320_));
 sg13g2_a21oi_1 _0805_ (.A1(net207),
    .A2(_0320_),
    .Y(_0084_),
    .B1(net110));
 sg13g2_and2_1 _0806_ (.A(\e.buf_.io_out_valid ),
    .B(\e.updateKey ),
    .X(_0321_));
 sg13g2_nand2_2 _0807_ (.Y(_0322_),
    .A(\e.buf_.io_out_valid ),
    .B(\e.updateKey ));
 sg13g2_a21oi_1 _0808_ (.A1(net184),
    .A2(net105),
    .Y(_0323_),
    .B1(net110));
 sg13g2_o21ai_1 _0809_ (.B1(_0323_),
    .Y(_0085_),
    .A1(_0096_),
    .A2(net105));
 sg13g2_nor2_1 _0810_ (.A(\e.buf_.dataReg[1] ),
    .B(_0322_),
    .Y(_0324_));
 sg13g2_nor2_1 _0811_ (.A(net188),
    .B(net106),
    .Y(_0325_));
 sg13g2_nor3_1 _0812_ (.A(net115),
    .B(_0324_),
    .C(_0325_),
    .Y(_0086_));
 sg13g2_a21oi_1 _0813_ (.A1(\e.buf_.dataReg[2] ),
    .A2(net106),
    .Y(_0326_),
    .B1(net117));
 sg13g2_o21ai_1 _0814_ (.B1(_0326_),
    .Y(_0087_),
    .A1(_0095_),
    .A2(net105));
 sg13g2_nor2_1 _0815_ (.A(net197),
    .B(_0322_),
    .Y(_0327_));
 sg13g2_nor2_1 _0816_ (.A(net198),
    .B(net106),
    .Y(_0328_));
 sg13g2_nor3_1 _0817_ (.A(net117),
    .B(_0327_),
    .C(_0328_),
    .Y(_0088_));
 sg13g2_a21oi_1 _0818_ (.A1(net196),
    .A2(net105),
    .Y(_0329_),
    .B1(net117));
 sg13g2_o21ai_1 _0819_ (.B1(_0329_),
    .Y(_0089_),
    .A1(_0094_),
    .A2(net105));
 sg13g2_nor2_1 _0820_ (.A(net178),
    .B(_0322_),
    .Y(_0330_));
 sg13g2_nor2_1 _0821_ (.A(net186),
    .B(net106),
    .Y(_0331_));
 sg13g2_nor3_1 _0822_ (.A(net117),
    .B(_0330_),
    .C(_0331_),
    .Y(_0090_));
 sg13g2_a21oi_1 _0823_ (.A1(\e.buf_.dataReg[6] ),
    .A2(net105),
    .Y(_0332_),
    .B1(net115));
 sg13g2_o21ai_1 _0824_ (.B1(_0332_),
    .Y(_0091_),
    .A1(_0093_),
    .A2(net105));
 sg13g2_nor2_1 _0825_ (.A(\e.buf_.dataReg[7] ),
    .B(_0322_),
    .Y(_0333_));
 sg13g2_nor2_1 _0826_ (.A(net216),
    .B(net105),
    .Y(_0334_));
 sg13g2_nor3_1 _0827_ (.A(net115),
    .B(_0333_),
    .C(_0334_),
    .Y(_0092_));
 sg13g2_dfrbp_1 _0828_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net64),
    .D(_0009_),
    .Q_N(_0411_),
    .Q(\e.tx.cntReg[0] ));
 sg13g2_dfrbp_1 _0829_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net27),
    .D(_0010_),
    .Q_N(_0410_),
    .Q(\e.tx.cntReg[1] ));
 sg13g2_dfrbp_1 _0830_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net26),
    .D(_0011_),
    .Q_N(_0409_),
    .Q(\e.tx.cntReg[2] ));
 sg13g2_dfrbp_1 _0831_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net141),
    .D(_0012_),
    .Q_N(_0408_),
    .Q(\e.tx.cntReg[4] ));
 sg13g2_dfrbp_1 _0832_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net140),
    .D(_0013_),
    .Q_N(_0407_),
    .Q(\e.tx.cntReg[6] ));
 sg13g2_dfrbp_1 _0833_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net139),
    .D(_0014_),
    .Q_N(_0006_),
    .Q(\e.tx.cntReg[10] ));
 sg13g2_dfrbp_1 _0834_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net138),
    .D(_0015_),
    .Q_N(_0406_),
    .Q(\e.tx.cntReg[12] ));
 sg13g2_dfrbp_1 _0835_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net137),
    .D(net226),
    .Q_N(_0405_),
    .Q(\e.tx.cntReg[3] ));
 sg13g2_dfrbp_1 _0836_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net136),
    .D(net157),
    .Q_N(_0404_),
    .Q(\e.tx.cntReg[5] ));
 sg13g2_dfrbp_1 _0837_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net135),
    .D(_0018_),
    .Q_N(_0403_),
    .Q(\e.tx.cntReg[7] ));
 sg13g2_dfrbp_1 _0838_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net134),
    .D(_0019_),
    .Q_N(_0402_),
    .Q(\e.tx.cntReg[8] ));
 sg13g2_dfrbp_1 _0839_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net133),
    .D(_0020_),
    .Q_N(_0401_),
    .Q(\e.tx.cntReg[9] ));
 sg13g2_dfrbp_1 _0840_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net132),
    .D(_0021_),
    .Q_N(_0400_),
    .Q(\e.tx.cntReg[11] ));
 sg13g2_dfrbp_1 _0841_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net131),
    .D(_0022_),
    .Q_N(_0399_),
    .Q(\e.tx.cntReg[13] ));
 sg13g2_dfrbp_1 _0842_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net130),
    .D(_0023_),
    .Q_N(_0007_),
    .Q(\e.tx.cntReg[14] ));
 sg13g2_dfrbp_1 _0843_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net129),
    .D(net151),
    .Q_N(_0398_),
    .Q(\e.tx.cntReg[15] ));
 sg13g2_dfrbp_1 _0844_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net128),
    .D(_0025_),
    .Q_N(_0397_),
    .Q(\e.tx.cntReg[16] ));
 sg13g2_dfrbp_1 _0845_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net127),
    .D(_0026_),
    .Q_N(_0396_),
    .Q(\e.tx.cntReg[17] ));
 sg13g2_dfrbp_1 _0846_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net126),
    .D(_0027_),
    .Q_N(_0008_),
    .Q(\e.tx.cntReg[18] ));
 sg13g2_dfrbp_1 _0847_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net125),
    .D(net181),
    .Q_N(_0395_),
    .Q(\e.tx.cntReg[19] ));
 sg13g2_dfrbp_1 _0848_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net124),
    .D(net167),
    .Q_N(_0394_),
    .Q(\e.io_txd ));
 sg13g2_dfrbp_1 _0849_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net122),
    .D(net215),
    .Q_N(_0393_),
    .Q(\e.tx._shiftReg_T_1[0] ));
 sg13g2_dfrbp_1 _0850_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net90),
    .D(net228),
    .Q_N(_0392_),
    .Q(\e.tx._shiftReg_T_1[1] ));
 sg13g2_dfrbp_1 _0851_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net88),
    .D(net209),
    .Q_N(_0391_),
    .Q(\e.tx._shiftReg_T_1[2] ));
 sg13g2_dfrbp_1 _0852_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net86),
    .D(_0033_),
    .Q_N(_0390_),
    .Q(\e.tx._shiftReg_T_1[3] ));
 sg13g2_dfrbp_1 _0853_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net84),
    .D(_0034_),
    .Q_N(_0389_),
    .Q(\e.tx._shiftReg_T_1[4] ));
 sg13g2_dfrbp_1 _0854_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net82),
    .D(net201),
    .Q_N(_0388_),
    .Q(\e.tx._shiftReg_T_1[5] ));
 sg13g2_dfrbp_1 _0855_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net80),
    .D(_0036_),
    .Q_N(_0387_),
    .Q(\e.tx._shiftReg_T_1[6] ));
 sg13g2_dfrbp_1 _0856_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net78),
    .D(net159),
    .Q_N(_0386_),
    .Q(\e.tx._shiftReg_T_1[7] ));
 sg13g2_dfrbp_1 _0857_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net76),
    .D(net269),
    .Q_N(_0385_),
    .Q(\e.updateKey ));
 sg13g2_dfrbp_1 _0858_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net75),
    .D(_0039_),
    .Q_N(_0384_),
    .Q(\e.buf_.dataReg[0] ));
 sg13g2_dfrbp_1 _0859_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net73),
    .D(net243),
    .Q_N(_0383_),
    .Q(\e.buf_.dataReg[1] ));
 sg13g2_dfrbp_1 _0860_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net71),
    .D(_0041_),
    .Q_N(_0382_),
    .Q(\e.buf_.dataReg[2] ));
 sg13g2_dfrbp_1 _0861_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net69),
    .D(_0042_),
    .Q_N(_0381_),
    .Q(\e.buf_.dataReg[3] ));
 sg13g2_dfrbp_1 _0862_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net67),
    .D(_0043_),
    .Q_N(_0380_),
    .Q(\e.buf_.dataReg[4] ));
 sg13g2_dfrbp_1 _0863_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net63),
    .D(_0044_),
    .Q_N(_0379_),
    .Q(\e.buf_.dataReg[5] ));
 sg13g2_dfrbp_1 _0864_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net61),
    .D(_0045_),
    .Q_N(_0378_),
    .Q(\e.buf_.dataReg[6] ));
 sg13g2_dfrbp_1 _0865_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net65),
    .D(_0046_),
    .Q_N(_0412_),
    .Q(\e.buf_.dataReg[7] ));
 sg13g2_dfrbp_1 _0866_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net32),
    .D(_0001_),
    .Q_N(_0413_),
    .Q(\e.rx.rxReg_REG ));
 sg13g2_dfrbp_1 _0867_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net59),
    .D(_0000_),
    .Q_N(_0377_),
    .Q(\e.rx.rxReg ));
 sg13g2_dfrbp_1 _0868_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net57),
    .D(net154),
    .Q_N(_0376_),
    .Q(\e.buf_.io_in_bits[0] ));
 sg13g2_dfrbp_1 _0869_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net55),
    .D(net195),
    .Q_N(_0375_),
    .Q(\e.buf_.io_in_bits[1] ));
 sg13g2_dfrbp_1 _0870_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net53),
    .D(net191),
    .Q_N(_0374_),
    .Q(\e.buf_.io_in_bits[2] ));
 sg13g2_dfrbp_1 _0871_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net51),
    .D(net174),
    .Q_N(_0373_),
    .Q(\e.buf_.io_in_bits[3] ));
 sg13g2_dfrbp_1 _0872_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net49),
    .D(_0051_),
    .Q_N(_0372_),
    .Q(\e.buf_.io_in_bits[4] ));
 sg13g2_dfrbp_1 _0873_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net47),
    .D(_0052_),
    .Q_N(_0371_),
    .Q(\e.buf_.io_in_bits[5] ));
 sg13g2_dfrbp_1 _0874_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net45),
    .D(net169),
    .Q_N(_0370_),
    .Q(\e.buf_.io_in_bits[6] ));
 sg13g2_dfrbp_1 _0875_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net43),
    .D(net204),
    .Q_N(_0369_),
    .Q(\e.buf_.io_in_bits[7] ));
 sg13g2_dfrbp_1 _0876_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net41),
    .D(_0055_),
    .Q_N(_0003_),
    .Q(\e.rx.cntReg[0] ));
 sg13g2_dfrbp_1 _0877_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net39),
    .D(net266),
    .Q_N(_0368_),
    .Q(\e.rx.cntReg[1] ));
 sg13g2_dfrbp_1 _0878_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net37),
    .D(_0057_),
    .Q_N(_0367_),
    .Q(\e.rx.cntReg[2] ));
 sg13g2_dfrbp_1 _0879_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net35),
    .D(net240),
    .Q_N(_0366_),
    .Q(\e.rx.cntReg[3] ));
 sg13g2_dfrbp_1 _0880_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net33),
    .D(_0059_),
    .Q_N(_0365_),
    .Q(\e.rx.cntReg[4] ));
 sg13g2_dfrbp_1 _0881_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net31),
    .D(_0060_),
    .Q_N(_0364_),
    .Q(\e.rx.cntReg[5] ));
 sg13g2_dfrbp_1 _0882_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net29),
    .D(_0061_),
    .Q_N(_0004_),
    .Q(\e.rx.cntReg[6] ));
 sg13g2_dfrbp_1 _0883_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net123),
    .D(_0062_),
    .Q_N(_0363_),
    .Q(\e.rx.cntReg[7] ));
 sg13g2_dfrbp_1 _0884_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(_0063_),
    .Q_N(_0362_),
    .Q(\e.rx.cntReg[8] ));
 sg13g2_dfrbp_1 _0885_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net85),
    .D(net251),
    .Q_N(_0361_),
    .Q(\e.rx.cntReg[9] ));
 sg13g2_dfrbp_1 _0886_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net81),
    .D(net163),
    .Q_N(_0005_),
    .Q(\e.rx.cntReg[10] ));
 sg13g2_dfrbp_1 _0887_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net77),
    .D(_0066_),
    .Q_N(_0360_),
    .Q(\e.rx.cntReg[11] ));
 sg13g2_dfrbp_1 _0888_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net72),
    .D(_0067_),
    .Q_N(_0359_),
    .Q(\e.rx.cntReg[12] ));
 sg13g2_dfrbp_1 _0889_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net68),
    .D(_0068_),
    .Q_N(_0358_),
    .Q(\e.rx.cntReg[13] ));
 sg13g2_dfrbp_1 _0890_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net62),
    .D(_0069_),
    .Q_N(_0357_),
    .Q(\e.rx.cntReg[14] ));
 sg13g2_dfrbp_1 _0891_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net58),
    .D(_0070_),
    .Q_N(_0356_),
    .Q(\e.rx.cntReg[15] ));
 sg13g2_dfrbp_1 _0892_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net54),
    .D(_0071_),
    .Q_N(_0355_),
    .Q(\e.rx.cntReg[16] ));
 sg13g2_dfrbp_1 _0893_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net50),
    .D(_0072_),
    .Q_N(_0354_),
    .Q(\e.rx.cntReg[17] ));
 sg13g2_dfrbp_1 _0894_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net46),
    .D(_0073_),
    .Q_N(_0353_),
    .Q(\e.rx.cntReg[18] ));
 sg13g2_dfrbp_1 _0895_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net42),
    .D(net148),
    .Q_N(_0352_),
    .Q(\e.rx.cntReg[19] ));
 sg13g2_dfrbp_1 _0896_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net38),
    .D(_0075_),
    .Q_N(_0351_),
    .Q(\e.rx.bitsReg[0] ));
 sg13g2_dfrbp_1 _0897_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net34),
    .D(_0076_),
    .Q_N(_0350_),
    .Q(\e.rx.bitsReg[1] ));
 sg13g2_dfrbp_1 _0898_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net30),
    .D(net220),
    .Q_N(_0349_),
    .Q(\e.rx.bitsReg[2] ));
 sg13g2_dfrbp_1 _0899_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net121),
    .D(net259),
    .Q_N(_0348_),
    .Q(\e.rx.bitsReg[3] ));
 sg13g2_dfrbp_1 _0900_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net83),
    .D(_0079_),
    .Q_N(_0347_),
    .Q(\e.buf_.io_in_valid ));
 sg13g2_dfrbp_1 _0901_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net74),
    .D(_0080_),
    .Q_N(_0002_),
    .Q(\e.buf_.io_out_valid ));
 sg13g2_dfrbp_1 _0902_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net70),
    .D(_0081_),
    .Q_N(_0346_),
    .Q(\e.tx.bitsReg[0] ));
 sg13g2_dfrbp_1 _0903_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net60),
    .D(net254),
    .Q_N(_0345_),
    .Q(\e.tx.bitsReg[1] ));
 sg13g2_dfrbp_1 _0904_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net52),
    .D(net172),
    .Q_N(_0344_),
    .Q(\e.tx.bitsReg[2] ));
 sg13g2_dfrbp_1 _0905_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net44),
    .D(_0084_),
    .Q_N(_0343_),
    .Q(\e.tx.bitsReg[3] ));
 sg13g2_dfrbp_1 _0906_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net36),
    .D(_0085_),
    .Q_N(_0342_),
    .Q(\e.key[0] ));
 sg13g2_dfrbp_1 _0907_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net28),
    .D(net189),
    .Q_N(_0341_),
    .Q(\e.key[1] ));
 sg13g2_dfrbp_1 _0908_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net79),
    .D(net183),
    .Q_N(_0340_),
    .Q(\e.key[2] ));
 sg13g2_dfrbp_1 _0909_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net56),
    .D(net199),
    .Q_N(_0339_),
    .Q(\e.key[3] ));
 sg13g2_dfrbp_1 _0910_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net40),
    .D(_0089_),
    .Q_N(_0338_),
    .Q(\e.key[4] ));
 sg13g2_dfrbp_1 _0911_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net87),
    .D(net187),
    .Q_N(_0337_),
    .Q(\e.key[5] ));
 sg13g2_dfrbp_1 _0912_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net48),
    .D(net193),
    .Q_N(_0336_),
    .Q(\e.key[6] ));
 sg13g2_dfrbp_1 _0913_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net66),
    .D(net217),
    .Q_N(_0335_),
    .Q(\e.key[7] ));
 sg13g2_tiehi _0829__27 (.L_HI(net27));
 sg13g2_tiehi _0907__28 (.L_HI(net28));
 sg13g2_tiehi _0882__29 (.L_HI(net29));
 sg13g2_tiehi _0898__30 (.L_HI(net30));
 sg13g2_tiehi _0881__31 (.L_HI(net31));
 sg13g2_tiehi _0866__32 (.L_HI(net32));
 sg13g2_tiehi _0880__33 (.L_HI(net33));
 sg13g2_tiehi _0897__34 (.L_HI(net34));
 sg13g2_tiehi _0879__35 (.L_HI(net35));
 sg13g2_tiehi _0906__36 (.L_HI(net36));
 sg13g2_tiehi _0878__37 (.L_HI(net37));
 sg13g2_tiehi _0896__38 (.L_HI(net38));
 sg13g2_tiehi _0877__39 (.L_HI(net39));
 sg13g2_tiehi _0910__40 (.L_HI(net40));
 sg13g2_tiehi _0876__41 (.L_HI(net41));
 sg13g2_tiehi _0895__42 (.L_HI(net42));
 sg13g2_tiehi _0875__43 (.L_HI(net43));
 sg13g2_tiehi _0905__44 (.L_HI(net44));
 sg13g2_tiehi _0874__45 (.L_HI(net45));
 sg13g2_tiehi _0894__46 (.L_HI(net46));
 sg13g2_tiehi _0873__47 (.L_HI(net47));
 sg13g2_tiehi _0912__48 (.L_HI(net48));
 sg13g2_tiehi _0872__49 (.L_HI(net49));
 sg13g2_tiehi _0893__50 (.L_HI(net50));
 sg13g2_tiehi _0871__51 (.L_HI(net51));
 sg13g2_tiehi _0904__52 (.L_HI(net52));
 sg13g2_tiehi _0870__53 (.L_HI(net53));
 sg13g2_tiehi _0892__54 (.L_HI(net54));
 sg13g2_tiehi _0869__55 (.L_HI(net55));
 sg13g2_tiehi _0909__56 (.L_HI(net56));
 sg13g2_tiehi _0868__57 (.L_HI(net57));
 sg13g2_tiehi _0891__58 (.L_HI(net58));
 sg13g2_tiehi _0867__59 (.L_HI(net59));
 sg13g2_tiehi _0903__60 (.L_HI(net60));
 sg13g2_tiehi _0864__61 (.L_HI(net61));
 sg13g2_tiehi _0890__62 (.L_HI(net62));
 sg13g2_tiehi _0863__63 (.L_HI(net63));
 sg13g2_tiehi _0828__64 (.L_HI(net64));
 sg13g2_tiehi _0865__65 (.L_HI(net65));
 sg13g2_tiehi _0913__66 (.L_HI(net66));
 sg13g2_tiehi _0862__67 (.L_HI(net67));
 sg13g2_tiehi _0889__68 (.L_HI(net68));
 sg13g2_tiehi _0861__69 (.L_HI(net69));
 sg13g2_tiehi _0902__70 (.L_HI(net70));
 sg13g2_tiehi _0860__71 (.L_HI(net71));
 sg13g2_tiehi _0888__72 (.L_HI(net72));
 sg13g2_tiehi _0859__73 (.L_HI(net73));
 sg13g2_tiehi _0901__74 (.L_HI(net74));
 sg13g2_tiehi _0858__75 (.L_HI(net75));
 sg13g2_tiehi _0857__76 (.L_HI(net76));
 sg13g2_tiehi _0887__77 (.L_HI(net77));
 sg13g2_tiehi _0856__78 (.L_HI(net78));
 sg13g2_tiehi _0908__79 (.L_HI(net79));
 sg13g2_tiehi _0855__80 (.L_HI(net80));
 sg13g2_tiehi _0886__81 (.L_HI(net81));
 sg13g2_tiehi _0854__82 (.L_HI(net82));
 sg13g2_tiehi _0900__83 (.L_HI(net83));
 sg13g2_tiehi _0853__84 (.L_HI(net84));
 sg13g2_tiehi _0885__85 (.L_HI(net85));
 sg13g2_tiehi _0852__86 (.L_HI(net86));
 sg13g2_tiehi _0911__87 (.L_HI(net87));
 sg13g2_tiehi _0851__88 (.L_HI(net88));
 sg13g2_tiehi _0884__89 (.L_HI(net89));
 sg13g2_tiehi _0850__90 (.L_HI(net90));
 sg13g2_tiehi _0899__91 (.L_HI(net121));
 sg13g2_tiehi _0849__92 (.L_HI(net122));
 sg13g2_tiehi _0883__93 (.L_HI(net123));
 sg13g2_tiehi _0848__94 (.L_HI(net124));
 sg13g2_tiehi _0847__95 (.L_HI(net125));
 sg13g2_tiehi _0846__96 (.L_HI(net126));
 sg13g2_tiehi _0845__97 (.L_HI(net127));
 sg13g2_tiehi _0844__98 (.L_HI(net128));
 sg13g2_tiehi _0843__99 (.L_HI(net129));
 sg13g2_tiehi _0842__100 (.L_HI(net130));
 sg13g2_tiehi _0841__101 (.L_HI(net131));
 sg13g2_tiehi _0840__102 (.L_HI(net132));
 sg13g2_tiehi _0839__103 (.L_HI(net133));
 sg13g2_tiehi _0838__104 (.L_HI(net134));
 sg13g2_tiehi _0837__105 (.L_HI(net135));
 sg13g2_tiehi _0836__106 (.L_HI(net136));
 sg13g2_tiehi _0835__107 (.L_HI(net137));
 sg13g2_tiehi _0834__108 (.L_HI(net138));
 sg13g2_tiehi _0833__109 (.L_HI(net139));
 sg13g2_tiehi _0832__110 (.L_HI(net140));
 sg13g2_tiehi _0831__111 (.L_HI(net141));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_UartMain_4 (.L_LO(net4));
 sg13g2_tielo tt_um_UartMain_5 (.L_LO(net5));
 sg13g2_tielo tt_um_UartMain_6 (.L_LO(net6));
 sg13g2_tielo tt_um_UartMain_7 (.L_LO(net7));
 sg13g2_tielo tt_um_UartMain_8 (.L_LO(net8));
 sg13g2_tielo tt_um_UartMain_9 (.L_LO(net9));
 sg13g2_tielo tt_um_UartMain_10 (.L_LO(net10));
 sg13g2_tielo tt_um_UartMain_11 (.L_LO(net11));
 sg13g2_tielo tt_um_UartMain_12 (.L_LO(net12));
 sg13g2_tielo tt_um_UartMain_13 (.L_LO(net13));
 sg13g2_tielo tt_um_UartMain_14 (.L_LO(net14));
 sg13g2_tielo tt_um_UartMain_15 (.L_LO(net15));
 sg13g2_tielo tt_um_UartMain_16 (.L_LO(net16));
 sg13g2_tielo tt_um_UartMain_17 (.L_LO(net17));
 sg13g2_tielo tt_um_UartMain_18 (.L_LO(net18));
 sg13g2_tielo tt_um_UartMain_19 (.L_LO(net19));
 sg13g2_tielo tt_um_UartMain_20 (.L_LO(net20));
 sg13g2_tielo tt_um_UartMain_21 (.L_LO(net21));
 sg13g2_tielo tt_um_UartMain_22 (.L_LO(net22));
 sg13g2_tielo tt_um_UartMain_23 (.L_LO(net23));
 sg13g2_tielo tt_um_UartMain_24 (.L_LO(net24));
 sg13g2_tielo tt_um_UartMain_25 (.L_LO(net25));
 sg13g2_tiehi _0830__26 (.L_HI(net26));
 sg13g2_buf_1 _1023_ (.A(\e.io_txd ),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout91 (.A(_0266_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0135_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0135_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(net95),
    .X(net94));
 sg13g2_buf_1 fanout95 (.A(_0241_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0241_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0129_),
    .X(net97));
 sg13g2_buf_1 fanout98 (.A(_0129_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0129_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0226_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_0203_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(net103),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0160_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0117_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_0321_),
    .X(net105));
 sg13g2_buf_1 fanout106 (.A(_0321_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0202_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_0002_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(net120),
    .X(net109));
 sg13g2_buf_1 fanout110 (.A(net120),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(net120),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(net114),
    .X(net112));
 sg13g2_buf_1 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(net120),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(net119),
    .X(net115));
 sg13g2_buf_1 fanout116 (.A(net119),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(net119),
    .X(net117));
 sg13g2_buf_1 fanout118 (.A(net119),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(net120),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(rst_n),
    .X(net120));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[7]),
    .X(net2));
 sg13g2_tielo tt_um_UartMain_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0003_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold2 (.A(\e.tx.cntReg[0] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold3 (.A(\e.rx.rxReg_REG ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold4 (.A(\e.buf_.io_in_valid ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0310_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold6 (.A(\e.rx.cntReg[19] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0074_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold8 (.A(\e.tx.cntReg[15] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0146_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0024_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0006_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold12 (.A(\e.buf_.io_in_bits[0] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0047_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold14 (.A(\e.tx.cntReg[5] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0137_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0017_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold17 (.A(\e.tx._shiftReg_T_1[7] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0037_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold19 (.A(\e.rx.cntReg[12] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0286_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0005_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0065_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold23 (.A(\e.tx.cntReg[7] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0138_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold25 (.A(\e.io_txd ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0029_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold27 (.A(\e.buf_.io_in_bits[6] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0053_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold29 (.A(\e.tx.bitsReg[2] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0317_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0083_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold32 (.A(\e.buf_.io_in_bits[4] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0050_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold34 (.A(\e.rx.cntReg[15] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0292_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold36 (.A(\e.buf_.io_in_bits[5] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold37 (.A(\e.buf_.dataReg[5] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold38 (.A(\e.tx.cntReg[19] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0154_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0028_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold41 (.A(\e.key[2] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0087_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold43 (.A(\e.buf_.dataReg[0] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold44 (.A(\e.key[0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold45 (.A(\e.key[5] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0090_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold47 (.A(\e.key[1] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0086_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold49 (.A(\e.buf_.io_in_bits[3] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0049_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold51 (.A(\e.key[6] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0091_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold53 (.A(\e.buf_.io_in_bits[2] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0048_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold55 (.A(\e.buf_.dataReg[4] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold56 (.A(\e.buf_.dataReg[3] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold57 (.A(\e.key[3] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0088_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold59 (.A(\e.tx._shiftReg_T_1[5] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0035_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold61 (.A(\e.tx._shiftReg_T_1[6] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold62 (.A(\e.buf_.io_in_bits[7] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0054_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold64 (.A(\e.key[4] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold65 (.A(\e.tx.bitsReg[3] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0319_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold67 (.A(\e.tx._shiftReg_T_1[2] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0032_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0007_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0145_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold71 (.A(\e.buf_.dataReg[6] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold72 (.A(\e.tx._shiftReg_T_1[4] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold73 (.A(\e.tx._shiftReg_T_1[0] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0030_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold75 (.A(\e.key[7] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0092_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold77 (.A(\e.rx.bitsReg[2] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0306_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0077_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0008_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0153_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold82 (.A(\e.tx._shiftReg_T_1[3] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold83 (.A(\e.tx.cntReg[3] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0136_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0016_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold86 (.A(\e.tx._shiftReg_T_1[1] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0031_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold88 (.A(\e.tx.cntReg[1] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold89 (.A(\e.tx.cntReg[4] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0111_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold91 (.A(\e.tx.cntReg[11] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold92 (.A(\e.rx.bitsReg[0] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold93 (.A(\e.buf_.dataReg[7] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold94 (.A(\e.rx.cntReg[14] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0291_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold96 (.A(\e.rx.bitsReg[1] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold97 (.A(\e.rx.cntReg[3] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0267_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0058_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold100 (.A(\e.buf_.dataReg[1] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0207_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0040_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold103 (.A(\e.buf_.dataReg[2] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold104 (.A(\e.rx.cntReg[2] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0265_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold106 (.A(\e.tx.cntReg[9] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0140_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold108 (.A(\e.rx.cntReg[9] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0279_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0064_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold111 (.A(\e.tx.bitsReg[1] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0315_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0082_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0004_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0273_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold116 (.A(\e.rx.bitsReg[3] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0307_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0078_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold119 (.A(\e.tx.cntReg[8] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold120 (.A(\e.tx.cntReg[13] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0144_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold122 (.A(\e.tx.cntReg[6] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold123 (.A(\e.rx.cntReg[1] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0259_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0056_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold126 (.A(\e.tx.bitsReg[0] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold127 (.A(\e.updateKey ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0038_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold129 (.A(\e.tx.cntReg[2] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold130 (.A(\e.rx.cntReg[18] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0297_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold132 (.A(\e.rx.cntReg[17] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0296_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold134 (.A(\e.rx.cntReg[8] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold135 (.A(\e.tx.cntReg[17] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0152_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold137 (.A(\e.rx.cntReg[4] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0268_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold139 (.A(\e.rx.cntReg[11] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold140 (.A(\e.rx.cntReg[16] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold141 (.A(\e.rx.cntReg[7] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold142 (.A(\e.rx.cntReg[13] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0287_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold144 (.A(\e.buf_.io_out_valid ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold145 (.A(\e.rx.cntReg[5] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0269_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold147 (.A(\e.tx.cntReg[12] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0131_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold149 (.A(\e.tx.cntReg[16] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0148_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold151 (.A(\e.rx.cntReg[1] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold152 (.A(\e.tx.cntReg[9] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0118_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold154 (.A(\e.tx.cntReg[6] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold155 (.A(\e.rx.cntReg[6] ),
    .X(net296));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_231 ();
 sg13g2_fill_2 FILLER_14_235 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_278 ();
 sg13g2_fill_1 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_decap_8 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_310 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_fill_2 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_225 ();
 sg13g2_fill_1 FILLER_15_232 ();
 sg13g2_decap_4 FILLER_15_259 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_decap_4 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_273 ();
 sg13g2_fill_1 FILLER_15_313 ();
 sg13g2_fill_2 FILLER_15_318 ();
 sg13g2_fill_1 FILLER_15_320 ();
 sg13g2_decap_4 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_359 ();
 sg13g2_decap_4 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_fill_2 FILLER_16_196 ();
 sg13g2_fill_1 FILLER_16_198 ();
 sg13g2_fill_1 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_252 ();
 sg13g2_fill_2 FILLER_16_300 ();
 sg13g2_decap_4 FILLER_16_325 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_fill_2 FILLER_17_222 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_fill_1 FILLER_17_238 ();
 sg13g2_fill_2 FILLER_17_262 ();
 sg13g2_fill_2 FILLER_17_268 ();
 sg13g2_fill_1 FILLER_17_270 ();
 sg13g2_fill_1 FILLER_17_334 ();
 sg13g2_fill_1 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_4 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_300 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_fill_2 FILLER_19_294 ();
 sg13g2_fill_1 FILLER_19_388 ();
 sg13g2_fill_1 FILLER_19_398 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_fill_1 FILLER_20_220 ();
 sg13g2_fill_1 FILLER_20_230 ();
 sg13g2_fill_1 FILLER_20_259 ();
 sg13g2_fill_2 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_fill_2 FILLER_20_320 ();
 sg13g2_fill_2 FILLER_20_348 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_4 FILLER_21_216 ();
 sg13g2_decap_8 FILLER_21_241 ();
 sg13g2_decap_4 FILLER_21_248 ();
 sg13g2_fill_2 FILLER_21_274 ();
 sg13g2_fill_1 FILLER_21_276 ();
 sg13g2_fill_2 FILLER_21_349 ();
 sg13g2_fill_2 FILLER_21_361 ();
 sg13g2_fill_1 FILLER_21_377 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_4 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_247 ();
 sg13g2_decap_4 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_258 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_fill_2 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_348 ();
 sg13g2_fill_1 FILLER_22_350 ();
 sg13g2_fill_2 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_4 FILLER_23_170 ();
 sg13g2_fill_1 FILLER_23_174 ();
 sg13g2_fill_2 FILLER_23_209 ();
 sg13g2_fill_1 FILLER_23_211 ();
 sg13g2_fill_2 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_decap_4 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_4 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_131 ();
 sg13g2_decap_4 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_fill_2 FILLER_24_147 ();
 sg13g2_decap_4 FILLER_24_209 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_fill_2 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_4 FILLER_25_121 ();
 sg13g2_fill_2 FILLER_25_125 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_327 ();
 sg13g2_fill_1 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_128 ();
 sg13g2_fill_1 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_4 FILLER_26_224 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_decap_4 FILLER_26_234 ();
 sg13g2_fill_1 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_fill_1 FILLER_26_327 ();
 sg13g2_fill_2 FILLER_26_336 ();
 sg13g2_fill_2 FILLER_26_347 ();
 sg13g2_fill_1 FILLER_26_349 ();
 sg13g2_fill_2 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_117 ();
 sg13g2_fill_2 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_379 ();
 sg13g2_fill_1 FILLER_27_381 ();
 sg13g2_fill_2 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_4 FILLER_28_91 ();
 sg13g2_fill_2 FILLER_28_121 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_142 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_fill_1 FILLER_28_264 ();
 sg13g2_fill_2 FILLER_28_292 ();
 sg13g2_fill_1 FILLER_28_350 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_fill_1 FILLER_28_365 ();
 sg13g2_fill_1 FILLER_28_370 ();
 sg13g2_fill_1 FILLER_28_380 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_184 ();
 sg13g2_fill_2 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_fill_2 FILLER_29_363 ();
 sg13g2_fill_2 FILLER_29_369 ();
 sg13g2_fill_1 FILLER_29_371 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_2 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_fill_2 FILLER_30_212 ();
 sg13g2_fill_1 FILLER_30_214 ();
 sg13g2_fill_2 FILLER_30_220 ();
 sg13g2_fill_2 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_fill_1 FILLER_30_269 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_338 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_136 ();
 sg13g2_fill_2 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_84 ();
 sg13g2_fill_1 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_fill_2 FILLER_32_340 ();
 sg13g2_fill_1 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_383 ();
 sg13g2_fill_2 FILLER_32_393 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_4 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_95 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_fill_1 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_187 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_2 FILLER_34_222 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_238 ();
 sg13g2_fill_2 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_288 ();
 sg13g2_fill_1 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_130 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_fill_2 FILLER_35_346 ();
 sg13g2_fill_1 FILLER_35_368 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_114 ();
 sg13g2_decap_4 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_141 ();
 sg13g2_fill_2 FILLER_36_184 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_196 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_fill_2 FILLER_36_252 ();
 sg13g2_fill_2 FILLER_36_277 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_363 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_132 ();
 sg13g2_fill_2 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_185 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_fill_1 FILLER_37_343 ();
 sg13g2_fill_1 FILLER_37_367 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_fill_2 FILLER_38_272 ();
 sg13g2_fill_2 FILLER_38_339 ();
 sg13g2_fill_1 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_373 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
 assign uo_out[1] = net19;
 assign uo_out[2] = net20;
 assign uo_out[3] = net21;
 assign uo_out[4] = net22;
 assign uo_out[5] = net23;
 assign uo_out[6] = net24;
 assign uo_out[7] = net25;
endmodule

module tt_um_wokwi_413387065339458561 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire clknet_leaf_0_clk;
 wire \pixel_0[0] ;
 wire \pixel_0[10] ;
 wire \pixel_0[11] ;
 wire \pixel_0[12] ;
 wire \pixel_0[13] ;
 wire \pixel_0[14] ;
 wire \pixel_0[15] ;
 wire \pixel_0[16] ;
 wire \pixel_0[17] ;
 wire \pixel_0[18] ;
 wire \pixel_0[19] ;
 wire \pixel_0[1] ;
 wire \pixel_0[20] ;
 wire \pixel_0[21] ;
 wire \pixel_0[22] ;
 wire \pixel_0[23] ;
 wire \pixel_0[2] ;
 wire \pixel_0[3] ;
 wire \pixel_0[4] ;
 wire \pixel_0[5] ;
 wire \pixel_0[6] ;
 wire \pixel_0[7] ;
 wire \pixel_0[8] ;
 wire \pixel_0[9] ;
 wire \pixel_1[0] ;
 wire \pixel_1[10] ;
 wire \pixel_1[11] ;
 wire \pixel_1[12] ;
 wire \pixel_1[13] ;
 wire \pixel_1[14] ;
 wire \pixel_1[15] ;
 wire \pixel_1[16] ;
 wire \pixel_1[17] ;
 wire \pixel_1[18] ;
 wire \pixel_1[19] ;
 wire \pixel_1[1] ;
 wire \pixel_1[20] ;
 wire \pixel_1[21] ;
 wire \pixel_1[22] ;
 wire \pixel_1[23] ;
 wire \pixel_1[2] ;
 wire \pixel_1[3] ;
 wire \pixel_1[4] ;
 wire \pixel_1[5] ;
 wire \pixel_1[6] ;
 wire \pixel_1[7] ;
 wire \pixel_1[8] ;
 wire \pixel_1[9] ;
 wire \pixel_2[0] ;
 wire \pixel_2[10] ;
 wire \pixel_2[11] ;
 wire \pixel_2[12] ;
 wire \pixel_2[13] ;
 wire \pixel_2[14] ;
 wire \pixel_2[15] ;
 wire \pixel_2[16] ;
 wire \pixel_2[17] ;
 wire \pixel_2[18] ;
 wire \pixel_2[19] ;
 wire \pixel_2[1] ;
 wire \pixel_2[20] ;
 wire \pixel_2[21] ;
 wire \pixel_2[22] ;
 wire \pixel_2[23] ;
 wire \pixel_2[2] ;
 wire \pixel_2[3] ;
 wire \pixel_2[4] ;
 wire \pixel_2[5] ;
 wire \pixel_2[6] ;
 wire \pixel_2[7] ;
 wire \pixel_2[8] ;
 wire \pixel_2[9] ;
 wire \pixel_3[0] ;
 wire \pixel_3[10] ;
 wire \pixel_3[11] ;
 wire \pixel_3[12] ;
 wire \pixel_3[13] ;
 wire \pixel_3[14] ;
 wire \pixel_3[15] ;
 wire \pixel_3[16] ;
 wire \pixel_3[17] ;
 wire \pixel_3[18] ;
 wire \pixel_3[19] ;
 wire \pixel_3[1] ;
 wire \pixel_3[20] ;
 wire \pixel_3[21] ;
 wire \pixel_3[22] ;
 wire \pixel_3[23] ;
 wire \pixel_3[2] ;
 wire \pixel_3[3] ;
 wire \pixel_3[4] ;
 wire \pixel_3[5] ;
 wire \pixel_3[6] ;
 wire \pixel_3[7] ;
 wire \pixel_3[8] ;
 wire \pixel_3[9] ;
 wire \pixel_4[0] ;
 wire \pixel_4[10] ;
 wire \pixel_4[11] ;
 wire \pixel_4[12] ;
 wire \pixel_4[13] ;
 wire \pixel_4[14] ;
 wire \pixel_4[15] ;
 wire \pixel_4[16] ;
 wire \pixel_4[17] ;
 wire \pixel_4[18] ;
 wire \pixel_4[19] ;
 wire \pixel_4[1] ;
 wire \pixel_4[20] ;
 wire \pixel_4[21] ;
 wire \pixel_4[22] ;
 wire \pixel_4[23] ;
 wire \pixel_4[2] ;
 wire \pixel_4[3] ;
 wire \pixel_4[4] ;
 wire \pixel_4[5] ;
 wire \pixel_4[6] ;
 wire \pixel_4[7] ;
 wire \pixel_4[8] ;
 wire \pixel_4[9] ;
 wire \pixel_5[0] ;
 wire \pixel_5[10] ;
 wire \pixel_5[11] ;
 wire \pixel_5[12] ;
 wire \pixel_5[13] ;
 wire \pixel_5[14] ;
 wire \pixel_5[15] ;
 wire \pixel_5[16] ;
 wire \pixel_5[17] ;
 wire \pixel_5[18] ;
 wire \pixel_5[19] ;
 wire \pixel_5[1] ;
 wire \pixel_5[20] ;
 wire \pixel_5[21] ;
 wire \pixel_5[22] ;
 wire \pixel_5[23] ;
 wire \pixel_5[2] ;
 wire \pixel_5[3] ;
 wire \pixel_5[4] ;
 wire \pixel_5[5] ;
 wire \pixel_5[6] ;
 wire \pixel_5[7] ;
 wire \pixel_5[8] ;
 wire \pixel_5[9] ;
 wire \pixel_6[0] ;
 wire \pixel_6[10] ;
 wire \pixel_6[11] ;
 wire \pixel_6[12] ;
 wire \pixel_6[13] ;
 wire \pixel_6[14] ;
 wire \pixel_6[15] ;
 wire \pixel_6[16] ;
 wire \pixel_6[17] ;
 wire \pixel_6[18] ;
 wire \pixel_6[19] ;
 wire \pixel_6[1] ;
 wire \pixel_6[20] ;
 wire \pixel_6[21] ;
 wire \pixel_6[22] ;
 wire \pixel_6[23] ;
 wire \pixel_6[2] ;
 wire \pixel_6[3] ;
 wire \pixel_6[4] ;
 wire \pixel_6[5] ;
 wire \pixel_6[6] ;
 wire \pixel_6[7] ;
 wire \pixel_6[8] ;
 wire \pixel_6[9] ;
 wire \spi_in.bit_count[0] ;
 wire \spi_in.bit_count[1] ;
 wire \spi_in.bit_count[2] ;
 wire \spi_in.bit_count[3] ;
 wire \spi_in.bit_count[4] ;
 wire \spi_in.bit_count[5] ;
 wire \spi_in.bit_count[6] ;
 wire \spi_in.bit_count[7] ;
 wire \spi_in.bit_count[8] ;
 wire \spi_in.index[0] ;
 wire \spi_in.index[1] ;
 wire \spi_in.index[2] ;
 wire \spi_in.index[3] ;
 wire \spi_in.index[4] ;
 wire \spi_in.index[5] ;
 wire \spi_in.index[6] ;
 wire \spi_in.index[7] ;
 wire \spi_in.last_sck ;
 wire \spi_in.state[0] ;
 wire \spi_in.state[1] ;
 wire \spi_in.state[2] ;
 wire \uart_output.count[0] ;
 wire \uart_output.count[1] ;
 wire \uart_output.count[2] ;
 wire \uart_output.count[3] ;
 wire \uart_output.count[4] ;
 wire \uart_output.count[5] ;
 wire \uart_output.count[6] ;
 wire \uart_output.count[7] ;
 wire \uart_output.index[0] ;
 wire \uart_output.index[1] ;
 wire \uart_output.index[2] ;
 wire \uart_output.index[3] ;
 wire \uart_output.index[4] ;
 wire \uart_output.index[5] ;
 wire \uart_output.index[6] ;
 wire \uart_output.index[7] ;
 wire \uart_output.uart_out ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire \ws2812_out.counter[0] ;
 wire \ws2812_out.counter[10] ;
 wire \ws2812_out.counter[1] ;
 wire \ws2812_out.counter[2] ;
 wire \ws2812_out.counter[3] ;
 wire \ws2812_out.counter[4] ;
 wire \ws2812_out.counter[5] ;
 wire \ws2812_out.counter[6] ;
 wire \ws2812_out.counter[7] ;
 wire \ws2812_out.counter[8] ;
 wire \ws2812_out.counter[9] ;
 wire \ws2812_out.datacounter[0] ;
 wire \ws2812_out.datacounter[1] ;
 wire \ws2812_out.datacounter[2] ;
 wire \ws2812_out.datacounter[3] ;
 wire \ws2812_out.datacounter[4] ;
 wire \ws2812_out.datacounter[5] ;
 wire \ws2812_out.datacounter[6] ;
 wire \ws2812_out.datacounter[7] ;
 wire \ws2812_out.led_o ;
 wire \ws2812_out.state ;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1;
 wire net2;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;

 sg13g2_inv_1 _1847_ (.Y(_0949_),
    .A(\pixel_3[15] ));
 sg13g2_inv_1 _1848_ (.Y(_0950_),
    .A(\pixel_3[13] ));
 sg13g2_inv_1 _1849_ (.Y(_0951_),
    .A(\pixel_3[9] ));
 sg13g2_inv_1 _1850_ (.Y(_0952_),
    .A(net483));
 sg13g2_inv_1 _1851_ (.Y(_0953_),
    .A(\pixel_5[23] ));
 sg13g2_inv_1 _1852_ (.Y(_0954_),
    .A(\pixel_5[7] ));
 sg13g2_inv_1 _1853_ (.Y(_0955_),
    .A(\pixel_5[5] ));
 sg13g2_inv_1 _1854_ (.Y(_0956_),
    .A(\pixel_5[3] ));
 sg13g2_inv_1 _1855_ (.Y(_0957_),
    .A(\pixel_6[23] ));
 sg13g2_inv_1 _1856_ (.Y(_0958_),
    .A(net284));
 sg13g2_inv_1 _1857_ (.Y(_0959_),
    .A(net355));
 sg13g2_inv_1 _1858_ (.Y(_0960_),
    .A(\uart_output.index[7] ));
 sg13g2_inv_1 _1859_ (.Y(_0961_),
    .A(\uart_output.index[6] ));
 sg13g2_inv_1 _1860_ (.Y(_0962_),
    .A(\uart_output.index[5] ));
 sg13g2_inv_1 _1861_ (.Y(_0963_),
    .A(net937));
 sg13g2_inv_2 _1862_ (.Y(_0964_),
    .A(net939));
 sg13g2_inv_1 _1863_ (.Y(_0965_),
    .A(\ws2812_out.datacounter[7] ));
 sg13g2_inv_1 _1864_ (.Y(_0966_),
    .A(\ws2812_out.datacounter[5] ));
 sg13g2_inv_4 _1865_ (.A(\ws2812_out.datacounter[4] ),
    .Y(_0967_));
 sg13g2_inv_4 _1866_ (.A(net947),
    .Y(_0968_));
 sg13g2_inv_4 _1867_ (.A(net949),
    .Y(_0969_));
 sg13g2_inv_1 _1868_ (.Y(_0970_),
    .A(\ws2812_out.counter[8] ));
 sg13g2_inv_1 _1869_ (.Y(_0971_),
    .A(\ws2812_out.counter[0] ));
 sg13g2_inv_1 _1870_ (.Y(_0972_),
    .A(net924));
 sg13g2_inv_1 _1871_ (.Y(_0973_),
    .A(\uart_output.count[5] ));
 sg13g2_inv_4 _1872_ (.A(net1006),
    .Y(_0974_));
 sg13g2_inv_4 _1873_ (.A(net1002),
    .Y(_0975_));
 sg13g2_inv_2 _1874_ (.Y(_0976_),
    .A(net908));
 sg13g2_inv_1 _1875_ (.Y(_0977_),
    .A(_0008_));
 sg13g2_inv_1 _1876_ (.Y(_0978_),
    .A(_0012_));
 sg13g2_nor4_1 _1877_ (.A(_0958_),
    .B(net423),
    .C(net473),
    .D(net467),
    .Y(_0979_));
 sg13g2_nor2b_2 _1878_ (.A(\spi_in.last_sck ),
    .B_N(net1),
    .Y(_0980_));
 sg13g2_nand2b_2 _1879_ (.Y(_0981_),
    .B(net1),
    .A_N(\spi_in.last_sck ));
 sg13g2_nor4_1 _1880_ (.A(net463),
    .B(net418),
    .C(net452),
    .D(net457),
    .Y(_0982_));
 sg13g2_and3_1 _1881_ (.X(_0983_),
    .A(\spi_in.bit_count[5] ),
    .B(_0979_),
    .C(_0982_));
 sg13g2_nand2_1 _1882_ (.Y(_0984_),
    .A(_0980_),
    .B(_0983_));
 sg13g2_nand3_1 _1883_ (.B(net1007),
    .C(_0984_),
    .A(net475),
    .Y(_0985_));
 sg13g2_nand2_1 _1884_ (.Y(_0986_),
    .A(net934),
    .B(net1007));
 sg13g2_nor2_1 _1885_ (.A(\spi_in.bit_count[5] ),
    .B(_0981_),
    .Y(_0987_));
 sg13g2_nand3_1 _1886_ (.B(_0982_),
    .C(_0987_),
    .A(_0979_),
    .Y(_0988_));
 sg13g2_o21ai_1 _1887_ (.B1(_0985_),
    .Y(_0001_),
    .A1(_0986_),
    .A2(_0988_));
 sg13g2_and3_1 _1888_ (.X(_0989_),
    .A(net452),
    .B(\spi_in.bit_count[0] ),
    .C(_0980_));
 sg13g2_and4_1 _1889_ (.A(net418),
    .B(net452),
    .C(net457),
    .D(_0980_),
    .X(_0990_));
 sg13g2_and2_1 _1890_ (.A(net463),
    .B(_0990_),
    .X(_0991_));
 sg13g2_and2_1 _1891_ (.A(net467),
    .B(_0991_),
    .X(_0992_));
 sg13g2_nor3_1 _1892_ (.A(net423),
    .B(\spi_in.bit_count[6] ),
    .C(\spi_in.bit_count[5] ),
    .Y(_0993_));
 sg13g2_nand3_1 _1893_ (.B(_0992_),
    .C(_0993_),
    .A(net446),
    .Y(_0994_));
 sg13g2_nor2_1 _1894_ (.A(_0975_),
    .B(_0981_),
    .Y(_0995_));
 sg13g2_o21ai_1 _1895_ (.B1(net490),
    .Y(_0996_),
    .A1(_0994_),
    .A2(_0995_));
 sg13g2_nand3_1 _1896_ (.B(_0980_),
    .C(_0983_),
    .A(net475),
    .Y(_0997_));
 sg13g2_nand3_1 _1897_ (.B(net491),
    .C(_0997_),
    .A(net1005),
    .Y(_0000_));
 sg13g2_nand2b_1 _1898_ (.Y(_0998_),
    .B(_0988_),
    .A_N(_0986_));
 sg13g2_nor2b_1 _1899_ (.A(net1002),
    .B_N(\spi_in.state[0] ),
    .Y(_0999_));
 sg13g2_nand2_1 _1900_ (.Y(_1000_),
    .A(net1005),
    .B(_0999_));
 sg13g2_o21ai_1 _1901_ (.B1(_0998_),
    .Y(_0002_),
    .A1(net447),
    .A2(_1000_));
 sg13g2_nor2_1 _1902_ (.A(\ws2812_out.counter[1] ),
    .B(_0978_),
    .Y(_1001_));
 sg13g2_o21ai_1 _1903_ (.B1(_0014_),
    .Y(_1002_),
    .A1(_0013_),
    .A2(_1001_));
 sg13g2_nor2b_1 _1904_ (.A(net949),
    .B_N(net952),
    .Y(_1003_));
 sg13g2_nand2b_1 _1905_ (.Y(_1004_),
    .B(net952),
    .A_N(net950));
 sg13g2_nand2_1 _1906_ (.Y(_1005_),
    .A(\pixel_3[19] ),
    .B(net886));
 sg13g2_nor2b_1 _1907_ (.A(net953),
    .B_N(net949),
    .Y(_1006_));
 sg13g2_nand2b_1 _1908_ (.Y(_1007_),
    .B(net950),
    .A_N(net952));
 sg13g2_nand2_1 _1909_ (.Y(_1008_),
    .A(\pixel_3[21] ),
    .B(net884));
 sg13g2_and2_2 _1910_ (.A(net949),
    .B(net953),
    .X(_1009_));
 sg13g2_nand2_2 _1911_ (.Y(_1010_),
    .A(net949),
    .B(net953));
 sg13g2_nor2_1 _1912_ (.A(net949),
    .B(net952),
    .Y(_1011_));
 sg13g2_or2_2 _1913_ (.X(_1012_),
    .B(net953),
    .A(net951));
 sg13g2_a22oi_1 _1914_ (.Y(_1013_),
    .B1(net881),
    .B2(\pixel_3[17] ),
    .A2(net882),
    .A1(\pixel_3[23] ));
 sg13g2_nand4_1 _1915_ (.B(_1005_),
    .C(_1008_),
    .A(net964),
    .Y(_1014_),
    .D(_1013_));
 sg13g2_a21oi_1 _1916_ (.A1(\pixel_3[18] ),
    .A2(net886),
    .Y(_1015_),
    .B1(net963));
 sg13g2_nand2_1 _1917_ (.Y(_1016_),
    .A(\pixel_3[22] ),
    .B(_1009_));
 sg13g2_a22oi_1 _1918_ (.Y(_1017_),
    .B1(net881),
    .B2(\pixel_3[16] ),
    .A2(net884),
    .A1(\pixel_3[20] ));
 sg13g2_nand3_1 _1919_ (.B(_1016_),
    .C(_1017_),
    .A(_1015_),
    .Y(_1018_));
 sg13g2_a21oi_1 _1920_ (.A1(_1014_),
    .A2(_1018_),
    .Y(_1019_),
    .B1(_0968_));
 sg13g2_mux4_1 _1921_ (.S0(net968),
    .A0(\pixel_4[12] ),
    .A1(\pixel_4[13] ),
    .A2(\pixel_4[14] ),
    .A3(\pixel_4[15] ),
    .S1(net954),
    .X(_1020_));
 sg13g2_mux4_1 _1922_ (.S0(net967),
    .A0(\pixel_4[8] ),
    .A1(\pixel_4[9] ),
    .A2(\pixel_4[10] ),
    .A3(\pixel_4[11] ),
    .S1(net954),
    .X(_1021_));
 sg13g2_mux2_2 _1923_ (.A0(_1020_),
    .A1(_1021_),
    .S(_0969_),
    .X(_1022_));
 sg13g2_o21ai_1 _1924_ (.B1(_0967_),
    .Y(_1023_),
    .A1(net948),
    .A2(_1022_));
 sg13g2_nor2b_1 _1925_ (.A(net967),
    .B_N(\pixel_3[6] ),
    .Y(_1024_));
 sg13g2_a21oi_1 _1926_ (.A1(\pixel_3[7] ),
    .A2(net967),
    .Y(_1025_),
    .B1(_1024_));
 sg13g2_nor2b_1 _1927_ (.A(net967),
    .B_N(\pixel_3[4] ),
    .Y(_1026_));
 sg13g2_a21oi_2 _1928_ (.B1(_1026_),
    .Y(_1027_),
    .A2(net969),
    .A1(\pixel_3[5] ));
 sg13g2_a22oi_1 _1929_ (.Y(_1028_),
    .B1(_1027_),
    .B2(net884),
    .A2(_1025_),
    .A1(net882));
 sg13g2_nor2b_1 _1930_ (.A(net966),
    .B_N(\pixel_3[0] ),
    .Y(_1029_));
 sg13g2_a21oi_1 _1931_ (.A1(\pixel_3[1] ),
    .A2(net966),
    .Y(_1030_),
    .B1(_1029_));
 sg13g2_nor2b_1 _1932_ (.A(net966),
    .B_N(\pixel_3[2] ),
    .Y(_1031_));
 sg13g2_a21oi_1 _1933_ (.A1(\pixel_3[3] ),
    .A2(net965),
    .Y(_1032_),
    .B1(_1031_));
 sg13g2_a22oi_1 _1934_ (.Y(_1033_),
    .B1(_1032_),
    .B2(net886),
    .A2(_1030_),
    .A1(net880));
 sg13g2_a21oi_1 _1935_ (.A1(_1028_),
    .A2(_1033_),
    .Y(_1034_),
    .B1(\ws2812_out.datacounter[3] ));
 sg13g2_o21ai_1 _1936_ (.B1(net879),
    .Y(_1035_),
    .A1(\pixel_3[8] ),
    .A2(net957));
 sg13g2_a21oi_1 _1937_ (.A1(_0951_),
    .A2(net956),
    .Y(_1036_),
    .B1(_1035_));
 sg13g2_o21ai_1 _1938_ (.B1(net882),
    .Y(_1037_),
    .A1(\pixel_3[14] ),
    .A2(net957));
 sg13g2_a21oi_1 _1939_ (.A1(_0949_),
    .A2(net956),
    .Y(_1038_),
    .B1(_1037_));
 sg13g2_nor2b_1 _1940_ (.A(\pixel_3[11] ),
    .B_N(net956),
    .Y(_1039_));
 sg13g2_o21ai_1 _1941_ (.B1(net885),
    .Y(_1040_),
    .A1(\pixel_3[10] ),
    .A2(net956));
 sg13g2_o21ai_1 _1942_ (.B1(net883),
    .Y(_1041_),
    .A1(\pixel_3[12] ),
    .A2(net956));
 sg13g2_a21oi_1 _1943_ (.A1(_0950_),
    .A2(net956),
    .Y(_1042_),
    .B1(_1041_));
 sg13g2_o21ai_1 _1944_ (.B1(net948),
    .Y(_1043_),
    .A1(_1039_),
    .A2(_1040_));
 sg13g2_nor4_2 _1945_ (.A(_1036_),
    .B(_1038_),
    .C(_1042_),
    .Y(_1044_),
    .D(_1043_));
 sg13g2_nor3_1 _1946_ (.A(_0967_),
    .B(_1034_),
    .C(_1044_),
    .Y(_1045_));
 sg13g2_o21ai_1 _1947_ (.B1(_0966_),
    .Y(_1046_),
    .A1(_1019_),
    .A2(_1023_));
 sg13g2_nor2_1 _1948_ (.A(_1045_),
    .B(_1046_),
    .Y(_1047_));
 sg13g2_nor2b_1 _1949_ (.A(net960),
    .B_N(\pixel_2[18] ),
    .Y(_1048_));
 sg13g2_a21oi_1 _1950_ (.A1(\pixel_2[19] ),
    .A2(net960),
    .Y(_1049_),
    .B1(_1048_));
 sg13g2_nor2b_1 _1951_ (.A(net961),
    .B_N(\pixel_2[16] ),
    .Y(_1050_));
 sg13g2_a21oi_1 _1952_ (.A1(\pixel_2[17] ),
    .A2(net960),
    .Y(_1051_),
    .B1(_1050_));
 sg13g2_mux4_1 _1953_ (.S0(net961),
    .A0(\pixel_2[20] ),
    .A1(\pixel_2[21] ),
    .A2(\pixel_2[22] ),
    .A3(\pixel_2[23] ),
    .S1(net953),
    .X(_1052_));
 sg13g2_nand2b_1 _1954_ (.Y(_1053_),
    .B(net950),
    .A_N(_1052_));
 sg13g2_a221oi_1 _1955_ (.B2(net879),
    .C1(net948),
    .B1(_1051_),
    .A1(net885),
    .Y(_1054_),
    .A2(_1049_));
 sg13g2_mux4_1 _1956_ (.S0(net959),
    .A0(\pixel_2[4] ),
    .A1(\pixel_2[5] ),
    .A2(\pixel_2[6] ),
    .A3(\pixel_2[7] ),
    .S1(net952),
    .X(_1055_));
 sg13g2_o21ai_1 _1957_ (.B1(net948),
    .Y(_1056_),
    .A1(_0969_),
    .A2(_1055_));
 sg13g2_mux4_1 _1958_ (.S0(net961),
    .A0(\pixel_2[0] ),
    .A1(\pixel_2[1] ),
    .A2(\pixel_2[2] ),
    .A3(\pixel_2[3] ),
    .S1(net955),
    .X(_1057_));
 sg13g2_nor2_1 _1959_ (.A(net950),
    .B(_1057_),
    .Y(_1058_));
 sg13g2_o21ai_1 _1960_ (.B1(_0967_),
    .Y(_1059_),
    .A1(_1056_),
    .A2(_1058_));
 sg13g2_a21oi_1 _1961_ (.A1(_1053_),
    .A2(_1054_),
    .Y(_1060_),
    .B1(_1059_));
 sg13g2_nor2b_1 _1962_ (.A(net965),
    .B_N(\pixel_2[8] ),
    .Y(_1061_));
 sg13g2_a21oi_1 _1963_ (.A1(\pixel_2[9] ),
    .A2(net965),
    .Y(_1062_),
    .B1(_1061_));
 sg13g2_nor2b_1 _1964_ (.A(net965),
    .B_N(\pixel_2[10] ),
    .Y(_1063_));
 sg13g2_a21oi_1 _1965_ (.A1(\pixel_2[11] ),
    .A2(net965),
    .Y(_1064_),
    .B1(_1063_));
 sg13g2_mux4_1 _1966_ (.S0(net968),
    .A0(\pixel_2[12] ),
    .A1(\pixel_2[13] ),
    .A2(\pixel_2[14] ),
    .A3(\pixel_2[15] ),
    .S1(net955),
    .X(_1065_));
 sg13g2_nand2b_1 _1967_ (.Y(_1066_),
    .B(net951),
    .A_N(_1065_));
 sg13g2_a221oi_1 _1968_ (.B2(net887),
    .C1(net948),
    .B1(_1064_),
    .A1(net880),
    .Y(_1067_),
    .A2(_1062_));
 sg13g2_mux4_1 _1969_ (.S0(net965),
    .A0(\pixel_1[16] ),
    .A1(\pixel_1[17] ),
    .A2(\pixel_1[18] ),
    .A3(\pixel_1[19] ),
    .S1(net954),
    .X(_1068_));
 sg13g2_nor2_1 _1970_ (.A(net951),
    .B(_1068_),
    .Y(_1069_));
 sg13g2_mux4_1 _1971_ (.S0(net969),
    .A0(\pixel_1[20] ),
    .A1(\pixel_1[21] ),
    .A2(\pixel_1[22] ),
    .A3(\pixel_1[23] ),
    .S1(net954),
    .X(_1070_));
 sg13g2_o21ai_1 _1972_ (.B1(net947),
    .Y(_1071_),
    .A1(_0969_),
    .A2(_1070_));
 sg13g2_o21ai_1 _1973_ (.B1(\ws2812_out.datacounter[4] ),
    .Y(_1072_),
    .A1(_1069_),
    .A2(_1071_));
 sg13g2_a21oi_1 _1974_ (.A1(_1066_),
    .A2(_1067_),
    .Y(_1073_),
    .B1(_1072_));
 sg13g2_o21ai_1 _1975_ (.B1(\ws2812_out.datacounter[5] ),
    .Y(_1074_),
    .A1(_1060_),
    .A2(_1073_));
 sg13g2_nand2_1 _1976_ (.Y(_1075_),
    .A(_0965_),
    .B(_1074_));
 sg13g2_o21ai_1 _1977_ (.B1(\ws2812_out.datacounter[6] ),
    .Y(_1076_),
    .A1(_1047_),
    .A2(_1075_));
 sg13g2_a21oi_1 _1978_ (.A1(_0978_),
    .A2(_0013_),
    .Y(_1077_),
    .B1(\ws2812_out.counter[3] ));
 sg13g2_nor2_1 _1979_ (.A(_0014_),
    .B(_1077_),
    .Y(_1078_));
 sg13g2_o21ai_1 _1980_ (.B1(net959),
    .Y(_1079_),
    .A1(\pixel_0[19] ),
    .A2(_1004_));
 sg13g2_nor2_1 _1981_ (.A(\pixel_0[17] ),
    .B(_1012_),
    .Y(_1080_));
 sg13g2_nor2_1 _1982_ (.A(\pixel_0[23] ),
    .B(_1010_),
    .Y(_1081_));
 sg13g2_nor2_1 _1983_ (.A(\pixel_0[21] ),
    .B(_1007_),
    .Y(_1082_));
 sg13g2_nor4_1 _1984_ (.A(_1079_),
    .B(_1080_),
    .C(_1081_),
    .D(_1082_),
    .Y(_1083_));
 sg13g2_nor2_1 _1985_ (.A(\pixel_0[18] ),
    .B(_1004_),
    .Y(_1084_));
 sg13g2_nand3b_1 _1986_ (.B(net950),
    .C(net952),
    .Y(_1085_),
    .A_N(\pixel_0[22] ));
 sg13g2_o21ai_1 _1987_ (.B1(_1085_),
    .Y(_1086_),
    .A1(\pixel_0[20] ),
    .A2(_1007_));
 sg13g2_nor2_1 _1988_ (.A(\pixel_0[16] ),
    .B(_1012_),
    .Y(_1087_));
 sg13g2_nor4_1 _1989_ (.A(net959),
    .B(_1084_),
    .C(_1086_),
    .D(_1087_),
    .Y(_1088_));
 sg13g2_o21ai_1 _1990_ (.B1(_0968_),
    .Y(_1089_),
    .A1(_1083_),
    .A2(_1088_));
 sg13g2_nor2b_1 _1991_ (.A(net960),
    .B_N(\pixel_0[0] ),
    .Y(_1090_));
 sg13g2_a21oi_1 _1992_ (.A1(\pixel_0[1] ),
    .A2(net960),
    .Y(_1091_),
    .B1(_1090_));
 sg13g2_nor2b_1 _1993_ (.A(net956),
    .B_N(\pixel_0[2] ),
    .Y(_1092_));
 sg13g2_a21oi_1 _1994_ (.A1(\pixel_0[3] ),
    .A2(net957),
    .Y(_1093_),
    .B1(_1092_));
 sg13g2_a221oi_1 _1995_ (.B2(net885),
    .C1(_0968_),
    .B1(_1093_),
    .A1(net879),
    .Y(_1094_),
    .A2(_1091_));
 sg13g2_mux4_1 _1996_ (.S0(net958),
    .A0(\pixel_0[4] ),
    .A1(\pixel_0[5] ),
    .A2(\pixel_0[6] ),
    .A3(\pixel_0[7] ),
    .S1(net952),
    .X(_1095_));
 sg13g2_nand2b_1 _1997_ (.Y(_1096_),
    .B(net949),
    .A_N(_1095_));
 sg13g2_a21oi_1 _1998_ (.A1(_1094_),
    .A2(_1096_),
    .Y(_1097_),
    .B1(_0967_));
 sg13g2_nor2b_1 _1999_ (.A(net967),
    .B_N(\pixel_1[2] ),
    .Y(_1098_));
 sg13g2_a21oi_2 _2000_ (.B1(_1098_),
    .Y(_1099_),
    .A2(net967),
    .A1(\pixel_1[3] ));
 sg13g2_nor2b_1 _2001_ (.A(net967),
    .B_N(\pixel_1[0] ),
    .Y(_1100_));
 sg13g2_a21oi_2 _2002_ (.B1(_1100_),
    .Y(_1101_),
    .A2(net967),
    .A1(\pixel_1[1] ));
 sg13g2_mux4_1 _2003_ (.S0(net968),
    .A0(\pixel_1[4] ),
    .A1(\pixel_1[5] ),
    .A2(\pixel_1[6] ),
    .A3(\pixel_1[7] ),
    .S1(net954),
    .X(_1102_));
 sg13g2_nand2b_1 _2004_ (.Y(_1103_),
    .B(net951),
    .A_N(_1102_));
 sg13g2_a221oi_1 _2005_ (.B2(net880),
    .C1(net947),
    .B1(_1101_),
    .A1(net886),
    .Y(_1104_),
    .A2(_1099_));
 sg13g2_mux4_1 _2006_ (.S0(net959),
    .A0(\pixel_1[12] ),
    .A1(\pixel_1[13] ),
    .A2(\pixel_1[14] ),
    .A3(\pixel_1[15] ),
    .S1(net953),
    .X(_1105_));
 sg13g2_mux4_1 _2007_ (.S0(net960),
    .A0(\pixel_1[8] ),
    .A1(\pixel_1[9] ),
    .A2(\pixel_1[10] ),
    .A3(\pixel_1[11] ),
    .S1(net953),
    .X(_1106_));
 sg13g2_nor2_1 _2008_ (.A(net949),
    .B(_1106_),
    .Y(_1107_));
 sg13g2_nor2_1 _2009_ (.A(_0968_),
    .B(_1107_),
    .Y(_1108_));
 sg13g2_o21ai_1 _2010_ (.B1(_1108_),
    .Y(_1109_),
    .A1(_0969_),
    .A2(_1105_));
 sg13g2_a21oi_2 _2011_ (.B1(\ws2812_out.datacounter[4] ),
    .Y(_1110_),
    .A2(_1104_),
    .A1(_1103_));
 sg13g2_a22oi_1 _2012_ (.Y(_1111_),
    .B1(_1109_),
    .B2(_1110_),
    .A2(_1097_),
    .A1(_1089_));
 sg13g2_nor2b_1 _2013_ (.A(net968),
    .B_N(\pixel_0[12] ),
    .Y(_1112_));
 sg13g2_a21oi_2 _2014_ (.B1(_1112_),
    .Y(_1113_),
    .A2(net968),
    .A1(\pixel_0[13] ));
 sg13g2_nand3_1 _2015_ (.B(_0010_),
    .C(_0017_),
    .A(\ws2812_out.datacounter[5] ),
    .Y(_1114_));
 sg13g2_nor2b_1 _2016_ (.A(net962),
    .B_N(\pixel_0[8] ),
    .Y(_1115_));
 sg13g2_a21oi_1 _2017_ (.A1(\pixel_0[9] ),
    .A2(net962),
    .Y(_1116_),
    .B1(_1115_));
 sg13g2_mux4_1 _2018_ (.S0(net963),
    .A0(\pixel_0[10] ),
    .A1(\pixel_0[11] ),
    .A2(\pixel_0[14] ),
    .A3(\pixel_0[15] ),
    .S1(net951),
    .X(_1117_));
 sg13g2_nand2b_1 _2019_ (.Y(_1118_),
    .B(net954),
    .A_N(_1117_));
 sg13g2_a221oi_1 _2020_ (.B2(net880),
    .C1(_1114_),
    .B1(_1116_),
    .A1(net884),
    .Y(_1119_),
    .A2(_1113_));
 sg13g2_a221oi_1 _2021_ (.B2(_1119_),
    .C1(_0965_),
    .B1(_1118_),
    .A1(_0966_),
    .Y(_1120_),
    .A2(_1111_));
 sg13g2_nor2_1 _2022_ (.A(_1078_),
    .B(_1120_),
    .Y(_1121_));
 sg13g2_nor2_1 _2023_ (.A(\ws2812_out.datacounter[7] ),
    .B(\ws2812_out.datacounter[6] ),
    .Y(_1122_));
 sg13g2_a21oi_1 _2024_ (.A1(\pixel_4[18] ),
    .A2(net885),
    .Y(_1123_),
    .B1(net957));
 sg13g2_nand2_1 _2025_ (.Y(_1124_),
    .A(\pixel_4[20] ),
    .B(net883));
 sg13g2_a22oi_1 _2026_ (.Y(_1125_),
    .B1(net879),
    .B2(\pixel_4[16] ),
    .A2(net882),
    .A1(\pixel_4[22] ));
 sg13g2_nand3_1 _2027_ (.B(_1124_),
    .C(_1125_),
    .A(_1123_),
    .Y(_1126_));
 sg13g2_nand2_1 _2028_ (.Y(_1127_),
    .A(\pixel_4[17] ),
    .B(net879));
 sg13g2_nand2_1 _2029_ (.Y(_1128_),
    .A(\pixel_4[21] ),
    .B(net883));
 sg13g2_a22oi_1 _2030_ (.Y(_1129_),
    .B1(net882),
    .B2(\pixel_4[23] ),
    .A2(net885),
    .A1(\pixel_4[19] ));
 sg13g2_nand4_1 _2031_ (.B(_1127_),
    .C(_1128_),
    .A(net959),
    .Y(_1130_),
    .D(_1129_));
 sg13g2_a21o_1 _2032_ (.A2(_1130_),
    .A1(_1126_),
    .B1(net948),
    .X(_1131_));
 sg13g2_mux2_1 _2033_ (.A0(\pixel_4[0] ),
    .A1(\pixel_4[1] ),
    .S(net960),
    .X(_1132_));
 sg13g2_mux2_1 _2034_ (.A0(\pixel_4[2] ),
    .A1(\pixel_4[3] ),
    .S(net961),
    .X(_1133_));
 sg13g2_a221oi_1 _2035_ (.B2(net885),
    .C1(_0968_),
    .B1(_1133_),
    .A1(net881),
    .Y(_1134_),
    .A2(_1132_));
 sg13g2_a22oi_1 _2036_ (.Y(_1135_),
    .B1(_1009_),
    .B2(\pixel_4[7] ),
    .A2(net883),
    .A1(\pixel_4[5] ));
 sg13g2_a22oi_1 _2037_ (.Y(_1136_),
    .B1(net882),
    .B2(\pixel_4[6] ),
    .A2(net883),
    .A1(\pixel_4[4] ));
 sg13g2_mux2_1 _2038_ (.A0(_1136_),
    .A1(_1135_),
    .S(net961),
    .X(_1137_));
 sg13g2_a21oi_1 _2039_ (.A1(_1134_),
    .A2(_1137_),
    .Y(_1138_),
    .B1(_0967_));
 sg13g2_o21ai_1 _2040_ (.B1(net886),
    .Y(_1139_),
    .A1(\pixel_5[2] ),
    .A2(net962));
 sg13g2_a21oi_1 _2041_ (.A1(_0956_),
    .A2(net962),
    .Y(_1140_),
    .B1(_1139_));
 sg13g2_o21ai_1 _2042_ (.B1(net884),
    .Y(_1141_),
    .A1(\pixel_5[4] ),
    .A2(net968));
 sg13g2_a21oi_1 _2043_ (.A1(_0955_),
    .A2(net963),
    .Y(_1142_),
    .B1(_1141_));
 sg13g2_nor2b_1 _2044_ (.A(net962),
    .B_N(\pixel_5[0] ),
    .Y(_1143_));
 sg13g2_a21oi_1 _2045_ (.A1(\pixel_5[1] ),
    .A2(net962),
    .Y(_1144_),
    .B1(_1143_));
 sg13g2_a21oi_1 _2046_ (.A1(_0954_),
    .A2(net964),
    .Y(_1145_),
    .B1(_1010_));
 sg13g2_o21ai_1 _2047_ (.B1(_1145_),
    .Y(_1146_),
    .A1(\pixel_5[6] ),
    .A2(net962));
 sg13g2_o21ai_1 _2048_ (.B1(_1146_),
    .Y(_1147_),
    .A1(_1012_),
    .A2(_1144_));
 sg13g2_or4_1 _2049_ (.A(net947),
    .B(_1140_),
    .C(_1142_),
    .D(_1147_),
    .X(_1148_));
 sg13g2_mux2_1 _2050_ (.A0(\pixel_5[8] ),
    .A1(\pixel_5[9] ),
    .S(net961),
    .X(_1149_));
 sg13g2_mux2_1 _2051_ (.A0(\pixel_5[10] ),
    .A1(\pixel_5[11] ),
    .S(net961),
    .X(_1150_));
 sg13g2_mux4_1 _2052_ (.S0(net959),
    .A0(\pixel_5[12] ),
    .A1(\pixel_5[13] ),
    .A2(\pixel_5[14] ),
    .A3(\pixel_5[15] ),
    .S1(net952),
    .X(_1151_));
 sg13g2_nand2_1 _2053_ (.Y(_1152_),
    .A(net950),
    .B(_1151_));
 sg13g2_a221oi_1 _2054_ (.B2(net887),
    .C1(_0968_),
    .B1(_1150_),
    .A1(net881),
    .Y(_1153_),
    .A2(_1149_));
 sg13g2_a21oi_1 _2055_ (.A1(_1152_),
    .A2(_1153_),
    .Y(_1154_),
    .B1(\ws2812_out.datacounter[4] ));
 sg13g2_a221oi_1 _2056_ (.B2(_1154_),
    .C1(_0966_),
    .B1(_1148_),
    .A1(_1131_),
    .Y(_1155_),
    .A2(_1138_));
 sg13g2_a21oi_1 _2057_ (.A1(\pixel_6[14] ),
    .A2(net882),
    .Y(_1156_),
    .B1(net965));
 sg13g2_nand2_1 _2058_ (.Y(_1157_),
    .A(\pixel_6[10] ),
    .B(net886));
 sg13g2_a22oi_1 _2059_ (.Y(_1158_),
    .B1(net880),
    .B2(\pixel_6[8] ),
    .A2(net884),
    .A1(\pixel_6[12] ));
 sg13g2_nand3_1 _2060_ (.B(_1157_),
    .C(_1158_),
    .A(_1156_),
    .Y(_1159_));
 sg13g2_nand2_1 _2061_ (.Y(_1160_),
    .A(\pixel_6[13] ),
    .B(net884));
 sg13g2_nand2_1 _2062_ (.Y(_1161_),
    .A(\pixel_6[9] ),
    .B(net880));
 sg13g2_a22oi_1 _2063_ (.Y(_1162_),
    .B1(_1009_),
    .B2(\pixel_6[15] ),
    .A2(net886),
    .A1(\pixel_6[11] ));
 sg13g2_nand4_1 _2064_ (.B(_1160_),
    .C(_1161_),
    .A(net966),
    .Y(_1163_),
    .D(_1162_));
 sg13g2_a21o_1 _2065_ (.A2(_1163_),
    .A1(_1159_),
    .B1(net947),
    .X(_1164_));
 sg13g2_nand2b_1 _2066_ (.Y(_1165_),
    .B(net968),
    .A_N(\pixel_5[21] ));
 sg13g2_or2_1 _2067_ (.X(_1166_),
    .B(net968),
    .A(\pixel_5[20] ));
 sg13g2_nand3_1 _2068_ (.B(_1165_),
    .C(_1166_),
    .A(net884),
    .Y(_1167_));
 sg13g2_a21oi_1 _2069_ (.A1(_0953_),
    .A2(net963),
    .Y(_1168_),
    .B1(_1010_));
 sg13g2_o21ai_1 _2070_ (.B1(_1168_),
    .Y(_1169_),
    .A1(\pixel_5[22] ),
    .A2(net963));
 sg13g2_a22oi_1 _2071_ (.Y(_1170_),
    .B1(net880),
    .B2(\pixel_5[17] ),
    .A2(net886),
    .A1(\pixel_5[19] ));
 sg13g2_a22oi_1 _2072_ (.Y(_1171_),
    .B1(net880),
    .B2(\pixel_5[16] ),
    .A2(net887),
    .A1(\pixel_5[18] ));
 sg13g2_mux2_1 _2073_ (.A0(_1171_),
    .A1(_1170_),
    .S(net965),
    .X(_1172_));
 sg13g2_nand4_1 _2074_ (.B(_1167_),
    .C(_1169_),
    .A(net947),
    .Y(_1173_),
    .D(_1172_));
 sg13g2_and2_1 _2075_ (.A(\ws2812_out.datacounter[4] ),
    .B(_1173_),
    .X(_1174_));
 sg13g2_mux2_1 _2076_ (.A0(\pixel_6[6] ),
    .A1(\pixel_6[7] ),
    .S(net958),
    .X(_1175_));
 sg13g2_mux2_1 _2077_ (.A0(\pixel_6[4] ),
    .A1(\pixel_6[5] ),
    .S(net959),
    .X(_1176_));
 sg13g2_mux2_1 _2078_ (.A0(\pixel_6[2] ),
    .A1(\pixel_6[3] ),
    .S(net957),
    .X(_1177_));
 sg13g2_a22oi_1 _2079_ (.Y(_1178_),
    .B1(_1177_),
    .B2(net885),
    .A2(_1176_),
    .A1(net883));
 sg13g2_mux2_1 _2080_ (.A0(\pixel_6[0] ),
    .A1(\pixel_6[1] ),
    .S(net960),
    .X(_1179_));
 sg13g2_a221oi_1 _2081_ (.B2(net879),
    .C1(_0968_),
    .B1(_1179_),
    .A1(net882),
    .Y(_1180_),
    .A2(_1175_));
 sg13g2_mux2_1 _2082_ (.A0(\pixel_6[18] ),
    .A1(\pixel_6[19] ),
    .S(net956),
    .X(_1181_));
 sg13g2_or2_1 _2083_ (.X(_1182_),
    .B(net958),
    .A(\pixel_6[22] ));
 sg13g2_a21oi_1 _2084_ (.A1(_0957_),
    .A2(net957),
    .Y(_1183_),
    .B1(_1010_));
 sg13g2_a221oi_1 _2085_ (.B2(_1183_),
    .C1(net948),
    .B1(_1182_),
    .A1(net885),
    .Y(_1184_),
    .A2(_1181_));
 sg13g2_a22oi_1 _2086_ (.Y(_1185_),
    .B1(net879),
    .B2(\pixel_6[17] ),
    .A2(net883),
    .A1(\pixel_6[21] ));
 sg13g2_a22oi_1 _2087_ (.Y(_1186_),
    .B1(net879),
    .B2(\pixel_6[16] ),
    .A2(net883),
    .A1(\pixel_6[20] ));
 sg13g2_mux2_1 _2088_ (.A0(_1186_),
    .A1(_1185_),
    .S(net957),
    .X(_1187_));
 sg13g2_a22oi_1 _2089_ (.Y(_1188_),
    .B1(_1184_),
    .B2(_1187_),
    .A2(_1180_),
    .A1(_1178_));
 sg13g2_a221oi_1 _2090_ (.B2(_0967_),
    .C1(\ws2812_out.datacounter[5] ),
    .B1(_1188_),
    .A1(_1164_),
    .Y(_1189_),
    .A2(_1174_));
 sg13g2_o21ai_1 _2091_ (.B1(_1122_),
    .Y(_1190_),
    .A1(_1155_),
    .A2(_1189_));
 sg13g2_nand3_1 _2092_ (.B(_1121_),
    .C(_1190_),
    .A(_1076_),
    .Y(_1191_));
 sg13g2_or2_1 _2093_ (.X(_1192_),
    .B(\ws2812_out.counter[8] ),
    .A(\ws2812_out.counter[9] ));
 sg13g2_nor4_2 _2094_ (.A(\ws2812_out.counter[7] ),
    .B(\ws2812_out.counter[6] ),
    .C(\ws2812_out.counter[5] ),
    .Y(_1193_),
    .D(_1192_));
 sg13g2_nand3b_1 _2095_ (.B(\ws2812_out.state ),
    .C(_1193_),
    .Y(_1194_),
    .A_N(\ws2812_out.counter[10] ));
 sg13g2_a21oi_1 _2096_ (.A1(_1002_),
    .A2(_1191_),
    .Y(\ws2812_out.led_o ),
    .B1(_1194_));
 sg13g2_nand4_1 _2097_ (.B(\ws2812_out.counter[2] ),
    .C(\ws2812_out.counter[3] ),
    .A(\ws2812_out.counter[4] ),
    .Y(_1195_),
    .D(\ws2812_out.counter[1] ));
 sg13g2_a21oi_1 _2098_ (.A1(\ws2812_out.counter[10] ),
    .A2(_0971_),
    .Y(_1196_),
    .B1(_1195_));
 sg13g2_nand2_1 _2099_ (.Y(_1197_),
    .A(_0018_),
    .B(_1193_));
 sg13g2_o21ai_1 _2100_ (.B1(\ws2812_out.state ),
    .Y(_1198_),
    .A1(_1196_),
    .A2(_1197_));
 sg13g2_and2_1 _2101_ (.A(net1003),
    .B(_1198_),
    .X(_1199_));
 sg13g2_nor4_1 _2102_ (.A(\ws2812_out.counter[4] ),
    .B(\ws2812_out.counter[2] ),
    .C(\ws2812_out.counter[3] ),
    .D(\ws2812_out.counter[1] ),
    .Y(_1200_));
 sg13g2_nand4_1 _2103_ (.B(\ws2812_out.counter[7] ),
    .C(\ws2812_out.counter[6] ),
    .A(_0970_),
    .Y(_1201_),
    .D(\ws2812_out.counter[5] ));
 sg13g2_o21ai_1 _2104_ (.B1(_0019_),
    .Y(_1202_),
    .A1(_1200_),
    .A2(_1201_));
 sg13g2_o21ai_1 _2105_ (.B1(\ws2812_out.counter[10] ),
    .Y(_1203_),
    .A1(\ws2812_out.counter[9] ),
    .A2(_1202_));
 sg13g2_o21ai_1 _2106_ (.B1(_1199_),
    .Y(_1204_),
    .A1(\ws2812_out.state ),
    .A2(_1203_));
 sg13g2_nor2_1 _2107_ (.A(net381),
    .B(_1204_),
    .Y(_0024_));
 sg13g2_nand2_1 _2108_ (.Y(_1205_),
    .A(\ws2812_out.counter[1] ),
    .B(\ws2812_out.counter[0] ));
 sg13g2_xnor2_1 _2109_ (.Y(_1206_),
    .A(net488),
    .B(net381));
 sg13g2_nor2_1 _2110_ (.A(_1204_),
    .B(_1206_),
    .Y(_0025_));
 sg13g2_nor2_1 _2111_ (.A(net369),
    .B(_1205_),
    .Y(_1207_));
 sg13g2_and2_1 _2112_ (.A(net369),
    .B(_1205_),
    .X(_1208_));
 sg13g2_nor3_1 _2113_ (.A(_1204_),
    .B(_1207_),
    .C(net370),
    .Y(_0026_));
 sg13g2_xor2_1 _2114_ (.B(_1207_),
    .A(net444),
    .X(_1209_));
 sg13g2_nor2_1 _2115_ (.A(_1204_),
    .B(net445),
    .Y(_0027_));
 sg13g2_and4_1 _2116_ (.A(\ws2812_out.counter[2] ),
    .B(\ws2812_out.counter[3] ),
    .C(\ws2812_out.counter[1] ),
    .D(\ws2812_out.counter[0] ),
    .X(_1210_));
 sg13g2_xor2_1 _2117_ (.B(_1210_),
    .A(net461),
    .X(_1211_));
 sg13g2_nor2_1 _2118_ (.A(_1204_),
    .B(net462),
    .Y(_0028_));
 sg13g2_nor2b_1 _2119_ (.A(net507),
    .B_N(_1203_),
    .Y(_1212_));
 sg13g2_nand2_2 _2120_ (.Y(_1213_),
    .A(net1003),
    .B(_1212_));
 sg13g2_and2_1 _2121_ (.A(\ws2812_out.counter[4] ),
    .B(_1210_),
    .X(_1214_));
 sg13g2_and2_1 _2122_ (.A(net468),
    .B(_1214_),
    .X(_1215_));
 sg13g2_nor2_1 _2123_ (.A(net468),
    .B(_1214_),
    .Y(_1216_));
 sg13g2_nor3_1 _2124_ (.A(_1213_),
    .B(_1215_),
    .C(net469),
    .Y(_0029_));
 sg13g2_and2_1 _2125_ (.A(net471),
    .B(_1215_),
    .X(_1217_));
 sg13g2_nor2_1 _2126_ (.A(net471),
    .B(_1215_),
    .Y(_1218_));
 sg13g2_nor3_1 _2127_ (.A(_1213_),
    .B(_1217_),
    .C(_1218_),
    .Y(_0030_));
 sg13g2_and2_1 _2128_ (.A(net480),
    .B(_1217_),
    .X(_1219_));
 sg13g2_nor2_1 _2129_ (.A(net480),
    .B(_1217_),
    .Y(_1220_));
 sg13g2_nor3_1 _2130_ (.A(_1213_),
    .B(_1219_),
    .C(_1220_),
    .Y(_0031_));
 sg13g2_xor2_1 _2131_ (.B(_1219_),
    .A(net343),
    .X(_1221_));
 sg13g2_nor2_1 _2132_ (.A(_1204_),
    .B(net344),
    .Y(_0032_));
 sg13g2_nand3_1 _2133_ (.B(\ws2812_out.counter[8] ),
    .C(_1219_),
    .A(net509),
    .Y(_1222_));
 sg13g2_a21oi_1 _2134_ (.A1(\ws2812_out.counter[8] ),
    .A2(_1219_),
    .Y(_1223_),
    .B1(net509));
 sg13g2_nor2_1 _2135_ (.A(_1213_),
    .B(net510),
    .Y(_1224_));
 sg13g2_and2_1 _2136_ (.A(_1222_),
    .B(_1224_),
    .X(_0033_));
 sg13g2_xnor2_1 _2137_ (.Y(_1225_),
    .A(net300),
    .B(_1222_));
 sg13g2_nor2_1 _2138_ (.A(_1213_),
    .B(net301),
    .Y(_0034_));
 sg13g2_nand4_1 _2139_ (.B(\uart_output.count[4] ),
    .C(\uart_output.count[6] ),
    .A(_0973_),
    .Y(_1226_),
    .D(\uart_output.count[7] ));
 sg13g2_nor3_1 _2140_ (.A(\uart_output.count[1] ),
    .B(\uart_output.count[2] ),
    .C(_1226_),
    .Y(_1227_));
 sg13g2_nand3_1 _2141_ (.B(\uart_output.count[3] ),
    .C(_1227_),
    .A(\uart_output.count[0] ),
    .Y(_1228_));
 sg13g2_and2_2 _2142_ (.A(net1006),
    .B(_1228_),
    .X(_1229_));
 sg13g2_nand2_2 _2143_ (.Y(_1230_),
    .A(net1006),
    .B(_1228_));
 sg13g2_and2_1 _2144_ (.A(net250),
    .B(_1229_),
    .X(_0035_));
 sg13g2_xnor2_1 _2145_ (.Y(_1231_),
    .A(\uart_output.count[0] ),
    .B(net465));
 sg13g2_nor2_1 _2146_ (.A(_1230_),
    .B(net466),
    .Y(_0036_));
 sg13g2_and3_1 _2147_ (.X(_1232_),
    .A(\uart_output.count[0] ),
    .B(\uart_output.count[1] ),
    .C(net384));
 sg13g2_a21oi_1 _2148_ (.A1(\uart_output.count[0] ),
    .A2(\uart_output.count[1] ),
    .Y(_1233_),
    .B1(net384));
 sg13g2_nor3_1 _2149_ (.A(_1230_),
    .B(_1232_),
    .C(net385),
    .Y(_0037_));
 sg13g2_and2_1 _2150_ (.A(net401),
    .B(_1232_),
    .X(_1234_));
 sg13g2_nor2_1 _2151_ (.A(net401),
    .B(_1232_),
    .Y(_1235_));
 sg13g2_nor3_1 _2152_ (.A(_1230_),
    .B(_1234_),
    .C(net402),
    .Y(_0038_));
 sg13g2_and2_1 _2153_ (.A(net411),
    .B(_1234_),
    .X(_1236_));
 sg13g2_nor2_1 _2154_ (.A(net411),
    .B(_1234_),
    .Y(_1237_));
 sg13g2_nor3_1 _2155_ (.A(_1230_),
    .B(_1236_),
    .C(_1237_),
    .Y(_0039_));
 sg13g2_nor2_1 _2156_ (.A(net456),
    .B(_1236_),
    .Y(_1238_));
 sg13g2_and2_1 _2157_ (.A(net456),
    .B(_1236_),
    .X(_1239_));
 sg13g2_nor3_1 _2158_ (.A(_1230_),
    .B(_1238_),
    .C(_1239_),
    .Y(_0040_));
 sg13g2_nor2_1 _2159_ (.A(net413),
    .B(_1239_),
    .Y(_1240_));
 sg13g2_and2_1 _2160_ (.A(net413),
    .B(_1239_),
    .X(_1241_));
 sg13g2_nor3_1 _2161_ (.A(_1230_),
    .B(net414),
    .C(_1241_),
    .Y(_0041_));
 sg13g2_a21oi_1 _2162_ (.A1(net459),
    .A2(_1241_),
    .Y(_1242_),
    .B1(_1230_));
 sg13g2_o21ai_1 _2163_ (.B1(_1242_),
    .Y(_1243_),
    .A1(net459),
    .A2(_1241_));
 sg13g2_inv_1 _2164_ (.Y(_0042_),
    .A(_1243_));
 sg13g2_nor2_1 _2165_ (.A(net963),
    .B(_1198_),
    .Y(_1244_));
 sg13g2_a21oi_1 _2166_ (.A1(net963),
    .A2(_1198_),
    .Y(_1245_),
    .B1(net986));
 sg13g2_nand2b_1 _2167_ (.Y(_0043_),
    .B(_1245_),
    .A_N(_1244_));
 sg13g2_o21ai_1 _2168_ (.B1(net954),
    .Y(_1246_),
    .A1(net963),
    .A2(_1198_));
 sg13g2_nand2b_1 _2169_ (.Y(_1247_),
    .B(_1244_),
    .A_N(net954));
 sg13g2_nand3_1 _2170_ (.B(_1246_),
    .C(_1247_),
    .A(net1004),
    .Y(_0044_));
 sg13g2_nor2_1 _2171_ (.A(net951),
    .B(_1247_),
    .Y(_1248_));
 sg13g2_a21oi_1 _2172_ (.A1(net951),
    .A2(_1247_),
    .Y(_1249_),
    .B1(net986));
 sg13g2_nand2b_1 _2173_ (.Y(_0045_),
    .B(_1249_),
    .A_N(_1248_));
 sg13g2_nor3_1 _2174_ (.A(net947),
    .B(net962),
    .C(_1012_),
    .Y(_1250_));
 sg13g2_and2_1 _2175_ (.A(_0967_),
    .B(_1250_),
    .X(_1251_));
 sg13g2_inv_1 _2176_ (.Y(_1252_),
    .A(_1251_));
 sg13g2_nor2_1 _2177_ (.A(\ws2812_out.datacounter[5] ),
    .B(_1252_),
    .Y(_1253_));
 sg13g2_nand2_1 _2178_ (.Y(_1254_),
    .A(_1122_),
    .B(_1253_));
 sg13g2_nand2_1 _2179_ (.Y(_1255_),
    .A(net1003),
    .B(_1254_));
 sg13g2_o21ai_1 _2180_ (.B1(net1003),
    .Y(_1256_),
    .A1(_1198_),
    .A2(_1254_));
 sg13g2_xnor2_1 _2181_ (.Y(_1257_),
    .A(net947),
    .B(_1248_));
 sg13g2_nor2_1 _2182_ (.A(_1256_),
    .B(_1257_),
    .Y(_0046_));
 sg13g2_nand2_1 _2183_ (.Y(_1258_),
    .A(\ws2812_out.datacounter[4] ),
    .B(_1199_));
 sg13g2_or2_1 _2184_ (.X(_1259_),
    .B(_1255_),
    .A(_1198_));
 sg13g2_xor2_1 _2185_ (.B(_1250_),
    .A(net481),
    .X(_1260_));
 sg13g2_o21ai_1 _2186_ (.B1(_1258_),
    .Y(_0047_),
    .A1(_1259_),
    .A2(_1260_));
 sg13g2_o21ai_1 _2187_ (.B1(net499),
    .Y(_1261_),
    .A1(_1198_),
    .A2(_1252_));
 sg13g2_nand2b_1 _2188_ (.Y(_1262_),
    .B(_1253_),
    .A_N(_1198_));
 sg13g2_nand3_1 _2189_ (.B(_1261_),
    .C(_1262_),
    .A(net1003),
    .Y(_0048_));
 sg13g2_nand2_1 _2190_ (.Y(_1263_),
    .A(\ws2812_out.datacounter[6] ),
    .B(_1199_));
 sg13g2_xor2_1 _2191_ (.B(_1253_),
    .A(net441),
    .X(_1264_));
 sg13g2_o21ai_1 _2192_ (.B1(_1263_),
    .Y(_0049_),
    .A1(_1259_),
    .A2(_1264_));
 sg13g2_o21ai_1 _2193_ (.B1(net387),
    .Y(_1265_),
    .A1(\ws2812_out.datacounter[6] ),
    .A2(_1262_));
 sg13g2_nand2b_1 _2194_ (.Y(_0050_),
    .B(net388),
    .A_N(_1256_));
 sg13g2_nor2_1 _2195_ (.A(net940),
    .B(net942),
    .Y(_1266_));
 sg13g2_nand2_1 _2196_ (.Y(_1267_),
    .A(\uart_output.index[5] ),
    .B(net938));
 sg13g2_o21ai_1 _2197_ (.B1(_0961_),
    .Y(_1268_),
    .A1(_1266_),
    .A2(_1267_));
 sg13g2_nand2_1 _2198_ (.Y(_1269_),
    .A(\uart_output.index[7] ),
    .B(_1268_));
 sg13g2_nor2b_1 _2199_ (.A(_1228_),
    .B_N(_1269_),
    .Y(_1270_));
 sg13g2_mux2_1 _2200_ (.A0(_1270_),
    .A1(_1228_),
    .S(net946),
    .X(_1271_));
 sg13g2_and2_1 _2201_ (.A(net1006),
    .B(_1271_),
    .X(_0051_));
 sg13g2_nand2b_2 _2202_ (.Y(_1272_),
    .B(net945),
    .A_N(net944));
 sg13g2_nand2b_2 _2203_ (.Y(_1273_),
    .B(net944),
    .A_N(net946));
 sg13g2_nand2_2 _2204_ (.Y(_1274_),
    .A(net1006),
    .B(_1270_));
 sg13g2_a21oi_1 _2205_ (.A1(_1272_),
    .A2(_1273_),
    .Y(_1275_),
    .B1(_1274_));
 sg13g2_a21o_1 _2206_ (.A2(_1229_),
    .A1(net422),
    .B1(_1275_),
    .X(_0052_));
 sg13g2_nand2_1 _2207_ (.Y(_1276_),
    .A(net943),
    .B(_1229_));
 sg13g2_nand2_1 _2208_ (.Y(_1277_),
    .A(net422),
    .B(net946));
 sg13g2_nor2_1 _2209_ (.A(_0007_),
    .B(_1277_),
    .Y(_1278_));
 sg13g2_xnor2_1 _2210_ (.Y(_1279_),
    .A(net478),
    .B(_1277_));
 sg13g2_o21ai_1 _2211_ (.B1(_1276_),
    .Y(_0053_),
    .A1(_1274_),
    .A2(_1279_));
 sg13g2_nand2_1 _2212_ (.Y(_1280_),
    .A(net398),
    .B(_1229_));
 sg13g2_xor2_1 _2213_ (.B(_1278_),
    .A(_0006_),
    .X(_1281_));
 sg13g2_o21ai_1 _2214_ (.B1(_1280_),
    .Y(_0054_),
    .A1(_1274_),
    .A2(_1281_));
 sg13g2_nand2_1 _2215_ (.Y(_1282_),
    .A(net943),
    .B(net944));
 sg13g2_nand3_1 _2216_ (.B(net944),
    .C(net945),
    .A(net941),
    .Y(_1283_));
 sg13g2_nor2_1 _2217_ (.A(_0964_),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_nand2_1 _2218_ (.Y(_1285_),
    .A(net938),
    .B(_1284_));
 sg13g2_a21oi_1 _2219_ (.A1(_1269_),
    .A2(_1285_),
    .Y(_1286_),
    .B1(_1228_));
 sg13g2_nor2b_1 _2220_ (.A(_1228_),
    .B_N(_1284_),
    .Y(_1287_));
 sg13g2_o21ai_1 _2221_ (.B1(net1006),
    .Y(_1288_),
    .A1(net938),
    .A2(_1287_));
 sg13g2_nor2_1 _2222_ (.A(_1286_),
    .B(_1288_),
    .Y(_0055_));
 sg13g2_nand2_1 _2223_ (.Y(_1289_),
    .A(\uart_output.index[5] ),
    .B(_1229_));
 sg13g2_xnor2_1 _2224_ (.Y(_1290_),
    .A(net394),
    .B(_1285_));
 sg13g2_o21ai_1 _2225_ (.B1(_1289_),
    .Y(_0056_),
    .A1(_1274_),
    .A2(_1290_));
 sg13g2_nand2b_1 _2226_ (.Y(_1291_),
    .B(_1284_),
    .A_N(_1267_));
 sg13g2_and2_1 _2227_ (.A(_0004_),
    .B(_1291_),
    .X(_1292_));
 sg13g2_nor2_1 _2228_ (.A(_0004_),
    .B(_1291_),
    .Y(_1293_));
 sg13g2_nor3_1 _2229_ (.A(_1274_),
    .B(_1292_),
    .C(_1293_),
    .Y(_1294_));
 sg13g2_a21o_1 _2230_ (.A2(_1229_),
    .A1(net435),
    .B1(_1294_),
    .X(_0057_));
 sg13g2_nand2_1 _2231_ (.Y(_1295_),
    .A(\uart_output.index[7] ),
    .B(_1229_));
 sg13g2_xor2_1 _2232_ (.B(_1293_),
    .A(net437),
    .X(_1296_));
 sg13g2_o21ai_1 _2233_ (.B1(_1295_),
    .Y(_0058_),
    .A1(_1274_),
    .A2(net438));
 sg13g2_nand2b_1 _2234_ (.Y(_0059_),
    .B(net1005),
    .A_N(net1));
 sg13g2_or2_2 _2235_ (.X(_1297_),
    .B(_1273_),
    .A(net941));
 sg13g2_nand2b_1 _2236_ (.Y(_1298_),
    .B(net943),
    .A_N(net945));
 sg13g2_nand3_1 _2237_ (.B(_1272_),
    .C(_1273_),
    .A(net941),
    .Y(_1299_));
 sg13g2_nand3_1 _2238_ (.B(_1297_),
    .C(_1299_),
    .A(net939),
    .Y(_1300_));
 sg13g2_nand2_1 _2239_ (.Y(_1301_),
    .A(_0964_),
    .B(net945));
 sg13g2_nand3_1 _2240_ (.B(_1300_),
    .C(_1301_),
    .A(net937),
    .Y(_1302_));
 sg13g2_a21oi_2 _2241_ (.B1(net939),
    .Y(_1303_),
    .A2(_1273_),
    .A1(net943));
 sg13g2_and2_1 _2242_ (.A(_1297_),
    .B(_1303_),
    .X(_1304_));
 sg13g2_nand2b_1 _2243_ (.Y(_1305_),
    .B(net945),
    .A_N(net941));
 sg13g2_o21ai_1 _2244_ (.B1(net940),
    .Y(_1306_),
    .A1(net942),
    .A2(_1272_));
 sg13g2_nor2b_1 _2245_ (.A(_1306_),
    .B_N(_1298_),
    .Y(_1307_));
 sg13g2_a22oi_1 _2246_ (.Y(_1308_),
    .B1(_1307_),
    .B2(_1282_),
    .A2(_1304_),
    .A1(_1272_));
 sg13g2_o21ai_1 _2247_ (.B1(_1302_),
    .Y(_1309_),
    .A1(net937),
    .A2(_1308_));
 sg13g2_nand2_1 _2248_ (.Y(_1310_),
    .A(net941),
    .B(_0009_));
 sg13g2_and2_1 _2249_ (.A(net939),
    .B(_1310_),
    .X(_1311_));
 sg13g2_nor2_1 _2250_ (.A(net944),
    .B(net945),
    .Y(_1312_));
 sg13g2_nand2b_1 _2251_ (.Y(_1313_),
    .B(_1312_),
    .A_N(net941));
 sg13g2_a22oi_1 _2252_ (.Y(_1314_),
    .B1(_1311_),
    .B2(_1313_),
    .A2(_1303_),
    .A1(_1297_));
 sg13g2_or2_1 _2253_ (.X(_1315_),
    .B(_1314_),
    .A(net937));
 sg13g2_o21ai_1 _2254_ (.B1(_1303_),
    .Y(_1316_),
    .A1(net943),
    .A2(_0977_));
 sg13g2_nand3_1 _2255_ (.B(_1277_),
    .C(_1298_),
    .A(\uart_output.index[3] ),
    .Y(_1317_));
 sg13g2_and2_1 _2256_ (.A(net938),
    .B(_1317_),
    .X(_1318_));
 sg13g2_a21oi_1 _2257_ (.A1(_1316_),
    .A2(_1318_),
    .Y(_1319_),
    .B1(_0961_));
 sg13g2_a221oi_1 _2258_ (.B2(_1319_),
    .C1(_0962_),
    .B1(_1315_),
    .A1(_0961_),
    .Y(_1320_),
    .A2(_1309_));
 sg13g2_o21ai_1 _2259_ (.B1(_1299_),
    .Y(_1321_),
    .A1(net942),
    .A2(_1272_));
 sg13g2_xnor2_1 _2260_ (.Y(_1322_),
    .A(net942),
    .B(net944));
 sg13g2_o21ai_1 _2261_ (.B1(net937),
    .Y(_1323_),
    .A1(_1312_),
    .A2(_1322_));
 sg13g2_o21ai_1 _2262_ (.B1(_1323_),
    .Y(_1324_),
    .A1(net939),
    .A2(net945));
 sg13g2_nand2_1 _2263_ (.Y(_1325_),
    .A(_0964_),
    .B(_1322_));
 sg13g2_o21ai_1 _2264_ (.B1(_1321_),
    .Y(_1326_),
    .A1(net939),
    .A2(net945));
 sg13g2_a22oi_1 _2265_ (.Y(_1327_),
    .B1(_1326_),
    .B2(_0963_),
    .A2(_1325_),
    .A1(_1324_));
 sg13g2_nor2_1 _2266_ (.A(\uart_output.index[6] ),
    .B(_1327_),
    .Y(_1328_));
 sg13g2_and2_1 _2267_ (.A(_0964_),
    .B(_1283_),
    .X(_1329_));
 sg13g2_a221oi_1 _2268_ (.B2(_1297_),
    .C1(_0963_),
    .B1(_1329_),
    .A1(net939),
    .Y(_1330_),
    .A2(_1305_));
 sg13g2_nand2_1 _2269_ (.Y(_1331_),
    .A(net944),
    .B(_0007_));
 sg13g2_and2_1 _2270_ (.A(_0964_),
    .B(_1272_),
    .X(_1332_));
 sg13g2_a221oi_1 _2271_ (.B2(_1332_),
    .C1(net937),
    .B1(_1331_),
    .A1(net940),
    .Y(_1333_),
    .A2(_1299_));
 sg13g2_nor3_1 _2272_ (.A(_0961_),
    .B(_1330_),
    .C(_1333_),
    .Y(_1334_));
 sg13g2_nor3_1 _2273_ (.A(\uart_output.index[5] ),
    .B(_1328_),
    .C(_1334_),
    .Y(_1335_));
 sg13g2_o21ai_1 _2274_ (.B1(_0960_),
    .Y(_1336_),
    .A1(_1320_),
    .A2(_1335_));
 sg13g2_nand2_1 _2275_ (.Y(_1337_),
    .A(\uart_output.index[7] ),
    .B(_0004_));
 sg13g2_nand2b_1 _2276_ (.Y(_1338_),
    .B(_0009_),
    .A_N(net941));
 sg13g2_a22oi_1 _2277_ (.Y(_1339_),
    .B1(_1338_),
    .B2(_1303_),
    .A2(_1311_),
    .A1(_1297_));
 sg13g2_nand2_1 _2278_ (.Y(_1340_),
    .A(_0963_),
    .B(_1339_));
 sg13g2_nand2b_1 _2279_ (.Y(_1341_),
    .B(_1273_),
    .A_N(_1306_));
 sg13g2_nand3_1 _2280_ (.B(_1310_),
    .C(_1313_),
    .A(_0964_),
    .Y(_1342_));
 sg13g2_nand3_1 _2281_ (.B(_1341_),
    .C(_1342_),
    .A(net937),
    .Y(_1343_));
 sg13g2_nand3_1 _2282_ (.B(_1340_),
    .C(_1343_),
    .A(_0962_),
    .Y(_1344_));
 sg13g2_o21ai_1 _2283_ (.B1(net941),
    .Y(_1345_),
    .A1(net944),
    .A2(net946));
 sg13g2_a21oi_1 _2284_ (.A1(_1338_),
    .A2(_1345_),
    .Y(_1346_),
    .B1(net939));
 sg13g2_nor3_1 _2285_ (.A(net937),
    .B(_1307_),
    .C(_1346_),
    .Y(_1347_));
 sg13g2_nor3_1 _2286_ (.A(_0963_),
    .B(_1301_),
    .C(_1331_),
    .Y(_1348_));
 sg13g2_o21ai_1 _2287_ (.B1(\uart_output.index[5] ),
    .Y(_1349_),
    .A1(_1347_),
    .A2(_1348_));
 sg13g2_a21oi_1 _2288_ (.A1(_1344_),
    .A2(_1349_),
    .Y(_1350_),
    .B1(_1337_));
 sg13g2_nor3_1 _2289_ (.A(net993),
    .B(_1228_),
    .C(_1350_),
    .Y(_1351_));
 sg13g2_a22oi_1 _2290_ (.Y(_0060_),
    .B1(_1336_),
    .B2(_1351_),
    .A2(_1229_),
    .A1(_0959_));
 sg13g2_nor3_1 _2291_ (.A(\spi_in.bit_count[4] ),
    .B(\spi_in.bit_count[3] ),
    .C(net897),
    .Y(_1352_));
 sg13g2_nor3_1 _2292_ (.A(\spi_in.state[0] ),
    .B(_0981_),
    .C(_1352_),
    .Y(_1353_));
 sg13g2_nand2b_1 _2293_ (.Y(_1354_),
    .B(\spi_in.state[1] ),
    .A_N(_0983_));
 sg13g2_nand2_1 _2294_ (.Y(_1355_),
    .A(_1353_),
    .B(_1354_));
 sg13g2_inv_1 _2295_ (.Y(_1356_),
    .A(net777));
 sg13g2_nor2b_1 _2296_ (.A(\spi_in.state[1] ),
    .B_N(_1353_),
    .Y(_1357_));
 sg13g2_nand2b_1 _2297_ (.Y(_1358_),
    .B(_1353_),
    .A_N(\spi_in.state[1] ));
 sg13g2_nor2_2 _2298_ (.A(net893),
    .B(net804),
    .Y(_1359_));
 sg13g2_nand2_2 _2299_ (.Y(_1360_),
    .A(net935),
    .B(net828));
 sg13g2_a21oi_1 _2300_ (.A1(net917),
    .A2(_1360_),
    .Y(_1361_),
    .B1(net989));
 sg13g2_o21ai_1 _2301_ (.B1(_1361_),
    .Y(_0061_),
    .A1(net917),
    .A2(net777));
 sg13g2_nor2_1 _2302_ (.A(\spi_in.index[1] ),
    .B(_1356_),
    .Y(_1362_));
 sg13g2_nor2b_1 _2303_ (.A(\spi_in.index[1] ),
    .B_N(net917),
    .Y(_1363_));
 sg13g2_nor2b_1 _2304_ (.A(net917),
    .B_N(\spi_in.index[1] ),
    .Y(_1364_));
 sg13g2_nor2_2 _2305_ (.A(\spi_in.index[1] ),
    .B(net917),
    .Y(_1365_));
 sg13g2_or2_2 _2306_ (.X(_1366_),
    .B(net917),
    .A(\spi_in.index[1] ));
 sg13g2_nand2_2 _2307_ (.Y(_1367_),
    .A(\spi_in.index[1] ),
    .B(\spi_in.index[0] ));
 sg13g2_inv_1 _2308_ (.Y(_1368_),
    .A(_1367_));
 sg13g2_nor4_1 _2309_ (.A(net503),
    .B(net777),
    .C(_1365_),
    .D(_1368_),
    .Y(_1369_));
 sg13g2_o21ai_1 _2310_ (.B1(net1004),
    .Y(_0062_),
    .A1(_1362_),
    .A2(net504));
 sg13g2_o21ai_1 _2311_ (.B1(net484),
    .Y(_1370_),
    .A1(net777),
    .A2(_1366_));
 sg13g2_nor2_1 _2312_ (.A(net484),
    .B(_1366_),
    .Y(_1371_));
 sg13g2_o21ai_1 _2313_ (.B1(_1356_),
    .Y(_1372_),
    .A1(_0016_),
    .A2(_1371_));
 sg13g2_nand3_1 _2314_ (.B(_1370_),
    .C(_1372_),
    .A(net1004),
    .Y(_0063_));
 sg13g2_nand2_2 _2315_ (.Y(_1373_),
    .A(net916),
    .B(_1365_));
 sg13g2_and3_1 _2316_ (.X(_1374_),
    .A(net911),
    .B(net915),
    .C(_1365_));
 sg13g2_nand3_1 _2317_ (.B(net915),
    .C(_1365_),
    .A(net911),
    .Y(_1375_));
 sg13g2_xnor2_1 _2318_ (.Y(_1376_),
    .A(net910),
    .B(_1373_));
 sg13g2_xor2_1 _2319_ (.B(_1373_),
    .A(net910),
    .X(_1377_));
 sg13g2_a22oi_1 _2320_ (.Y(_1378_),
    .B1(_1359_),
    .B2(net865),
    .A2(net777),
    .A1(net911));
 sg13g2_nor2_1 _2321_ (.A(net989),
    .B(_1378_),
    .Y(_0064_));
 sg13g2_nor4_2 _2322_ (.A(net913),
    .B(\spi_in.index[2] ),
    .C(\spi_in.index[1] ),
    .Y(_1379_),
    .D(net917));
 sg13g2_nand2_1 _2323_ (.Y(_1380_),
    .A(net908),
    .B(_1379_));
 sg13g2_xnor2_1 _2324_ (.Y(_1381_),
    .A(_0976_),
    .B(_1379_));
 sg13g2_xnor2_1 _2325_ (.Y(_1382_),
    .A(net908),
    .B(_1379_));
 sg13g2_a22oi_1 _2326_ (.Y(_1383_),
    .B1(net776),
    .B2(net871),
    .A2(_1355_),
    .A1(net428));
 sg13g2_nor2_1 _2327_ (.A(net994),
    .B(_1383_),
    .Y(_0065_));
 sg13g2_nand2b_1 _2328_ (.Y(_1384_),
    .B(_1379_),
    .A_N(net428));
 sg13g2_o21ai_1 _2329_ (.B1(net902),
    .Y(_1385_),
    .A1(net777),
    .A2(_1384_));
 sg13g2_nor2_1 _2330_ (.A(net902),
    .B(\spi_in.index[4] ),
    .Y(_1386_));
 sg13g2_nand2_1 _2331_ (.Y(_1387_),
    .A(_1379_),
    .B(_1386_));
 sg13g2_a21oi_1 _2332_ (.A1(_1379_),
    .A2(_1386_),
    .Y(_1388_),
    .B1(net503));
 sg13g2_o21ai_1 _2333_ (.B1(net1005),
    .Y(_1389_),
    .A1(net777),
    .A2(_1388_));
 sg13g2_nand2b_1 _2334_ (.Y(_0066_),
    .B(_1385_),
    .A_N(_1389_));
 sg13g2_nand3b_1 _2335_ (.B(_1379_),
    .C(_1386_),
    .Y(_1390_),
    .A_N(\spi_in.index[6] ));
 sg13g2_xor2_1 _2336_ (.B(_1387_),
    .A(\spi_in.index[6] ),
    .X(_1391_));
 sg13g2_xnor2_1 _2337_ (.Y(_1392_),
    .A(\spi_in.index[6] ),
    .B(_1387_));
 sg13g2_a22oi_1 _2338_ (.Y(_1393_),
    .B1(net776),
    .B2(net857),
    .A2(_1355_),
    .A1(net487));
 sg13g2_nor2_1 _2339_ (.A(net997),
    .B(_1393_),
    .Y(_0067_));
 sg13g2_nor2_1 _2340_ (.A(net496),
    .B(_1356_),
    .Y(_1394_));
 sg13g2_nor4_1 _2341_ (.A(\spi_in.index[7] ),
    .B(\spi_in.index[6] ),
    .C(net902),
    .D(\spi_in.index[4] ),
    .Y(_1395_));
 sg13g2_and2_2 _2342_ (.A(_1379_),
    .B(_1395_),
    .X(_1396_));
 sg13g2_a21oi_1 _2343_ (.A1(\spi_in.index[7] ),
    .A2(_1390_),
    .Y(_1397_),
    .B1(_1396_));
 sg13g2_a21o_2 _2344_ (.A2(_1390_),
    .A1(\spi_in.index[7] ),
    .B1(_1396_),
    .X(_1398_));
 sg13g2_nor3_1 _2345_ (.A(_0016_),
    .B(net777),
    .C(_1398_),
    .Y(_1399_));
 sg13g2_o21ai_1 _2346_ (.B1(net1005),
    .Y(_0068_),
    .A1(_1394_),
    .A2(_1399_));
 sg13g2_nor2_1 _2347_ (.A(net934),
    .B(_0999_),
    .Y(_1400_));
 sg13g2_a21oi_1 _2348_ (.A1(_1354_),
    .A2(_1400_),
    .Y(_1401_),
    .B1(_0981_));
 sg13g2_o21ai_1 _2349_ (.B1(net1005),
    .Y(_1402_),
    .A1(net457),
    .A2(_1401_));
 sg13g2_a21oi_1 _2350_ (.A1(net457),
    .A2(_0980_),
    .Y(_0069_),
    .B1(_1402_));
 sg13g2_nor2_1 _2351_ (.A(\spi_in.state[0] ),
    .B(\spi_in.state[1] ),
    .Y(_1403_));
 sg13g2_a22oi_1 _2352_ (.Y(_1404_),
    .B1(_1403_),
    .B2(net897),
    .A2(_1400_),
    .A1(_0015_));
 sg13g2_nor2_1 _2353_ (.A(_0981_),
    .B(_1404_),
    .Y(_1405_));
 sg13g2_o21ai_1 _2354_ (.B1(net1005),
    .Y(_1406_),
    .A1(_0981_),
    .A2(_1404_));
 sg13g2_a21oi_1 _2355_ (.A1(\spi_in.bit_count[0] ),
    .A2(_0980_),
    .Y(_1407_),
    .B1(net452));
 sg13g2_nor3_1 _2356_ (.A(_0989_),
    .B(_1406_),
    .C(net453),
    .Y(_0070_));
 sg13g2_nor2_1 _2357_ (.A(net418),
    .B(_0989_),
    .Y(_1408_));
 sg13g2_nor3_1 _2358_ (.A(_0990_),
    .B(_1406_),
    .C(net419),
    .Y(_0071_));
 sg13g2_nor2_1 _2359_ (.A(net463),
    .B(_0990_),
    .Y(_1409_));
 sg13g2_nor3_1 _2360_ (.A(_0991_),
    .B(_1406_),
    .C(_1409_),
    .Y(_0072_));
 sg13g2_nor2_1 _2361_ (.A(net467),
    .B(_0991_),
    .Y(_1410_));
 sg13g2_nor3_1 _2362_ (.A(_0992_),
    .B(_1406_),
    .C(_1410_),
    .Y(_0073_));
 sg13g2_nor2_1 _2363_ (.A(net489),
    .B(_0992_),
    .Y(_1411_));
 sg13g2_nand2_1 _2364_ (.Y(_1412_),
    .A(_0983_),
    .B(_1400_));
 sg13g2_nor2_1 _2365_ (.A(_0981_),
    .B(_1412_),
    .Y(_1413_));
 sg13g2_and2_1 _2366_ (.A(net489),
    .B(_0992_),
    .X(_1414_));
 sg13g2_nor4_1 _2367_ (.A(_1406_),
    .B(_1411_),
    .C(_1413_),
    .D(_1414_),
    .Y(_0074_));
 sg13g2_nor2_1 _2368_ (.A(net473),
    .B(_1414_),
    .Y(_1415_));
 sg13g2_and2_1 _2369_ (.A(net473),
    .B(_1414_),
    .X(_0247_));
 sg13g2_nor3_1 _2370_ (.A(_1406_),
    .B(net474),
    .C(_0247_),
    .Y(_0075_));
 sg13g2_a21oi_1 _2371_ (.A1(_1404_),
    .A2(_0247_),
    .Y(_0248_),
    .B1(net423));
 sg13g2_o21ai_1 _2372_ (.B1(net423),
    .Y(_0249_),
    .A1(_1405_),
    .A2(_0247_));
 sg13g2_nand2_1 _2373_ (.Y(_0250_),
    .A(net1005),
    .B(_0249_));
 sg13g2_nor2_1 _2374_ (.A(net424),
    .B(_0250_),
    .Y(_0076_));
 sg13g2_nand2_1 _2375_ (.Y(_0251_),
    .A(net284),
    .B(_0981_));
 sg13g2_nand4_1 _2376_ (.B(\spi_in.bit_count[2] ),
    .C(\spi_in.bit_count[1] ),
    .A(\spi_in.bit_count[3] ),
    .Y(_0252_),
    .D(\spi_in.bit_count[0] ));
 sg13g2_nand4_1 _2377_ (.B(\spi_in.bit_count[6] ),
    .C(\spi_in.bit_count[5] ),
    .A(\spi_in.bit_count[7] ),
    .Y(_0253_),
    .D(\spi_in.bit_count[4] ));
 sg13g2_nor2_1 _2378_ (.A(_0252_),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_xnor2_1 _2379_ (.Y(_0255_),
    .A(_0020_),
    .B(_0254_));
 sg13g2_nand4_1 _2380_ (.B(_1404_),
    .C(_1412_),
    .A(_0980_),
    .Y(_0256_),
    .D(_0255_));
 sg13g2_a21oi_1 _2381_ (.A1(_0251_),
    .A2(_0256_),
    .Y(_0077_),
    .B1(net996));
 sg13g2_xor2_1 _2382_ (.B(_1380_),
    .A(net902),
    .X(_0257_));
 sg13g2_xnor2_1 _2383_ (.Y(_0258_),
    .A(net902),
    .B(_1380_));
 sg13g2_nand3_1 _2384_ (.B(_1396_),
    .C(net835),
    .A(net865),
    .Y(_0259_));
 sg13g2_a21oi_1 _2385_ (.A1(net925),
    .A2(_0259_),
    .Y(_0260_),
    .B1(net804));
 sg13g2_nand2b_1 _2386_ (.Y(_0261_),
    .B(net506),
    .A_N(_0260_));
 sg13g2_nor2_1 _2387_ (.A(_0975_),
    .B(_1360_),
    .Y(_0262_));
 sg13g2_nand2_2 _2388_ (.Y(_0263_),
    .A(net1001),
    .B(net776));
 sg13g2_o21ai_1 _2389_ (.B1(_0261_),
    .Y(_0264_),
    .A1(_0259_),
    .A2(_0263_));
 sg13g2_and2_1 _2390_ (.A(net1004),
    .B(_0264_),
    .X(_0078_));
 sg13g2_and2_2 _2391_ (.A(net915),
    .B(_1363_),
    .X(_0265_));
 sg13g2_nor2b_2 _2392_ (.A(net910),
    .B_N(_0265_),
    .Y(_0266_));
 sg13g2_nand4_1 _2393_ (.B(net861),
    .C(net842),
    .A(net875),
    .Y(_0267_),
    .D(_0266_));
 sg13g2_o21ai_1 _2394_ (.B1(net924),
    .Y(_0268_),
    .A1(net848),
    .A2(_0267_));
 sg13g2_nand2_1 _2395_ (.Y(_0269_),
    .A(net815),
    .B(_0268_));
 sg13g2_nor2_2 _2396_ (.A(net857),
    .B(net849),
    .Y(_0270_));
 sg13g2_nand2_1 _2397_ (.Y(_0271_),
    .A(net861),
    .B(net853));
 sg13g2_nand2_2 _2398_ (.Y(_0272_),
    .A(net1001),
    .B(_0265_));
 sg13g2_nand2b_2 _2399_ (.Y(_0273_),
    .B(net776),
    .A_N(net905));
 sg13g2_nor4_2 _2400_ (.A(net864),
    .B(net868),
    .C(_0272_),
    .Y(_0274_),
    .D(_0273_));
 sg13g2_a22oi_1 _2401_ (.Y(_0275_),
    .B1(net798),
    .B2(_0274_),
    .A2(_0269_),
    .A1(net366));
 sg13g2_nor2_1 _2402_ (.A(net982),
    .B(_0275_),
    .Y(_0079_));
 sg13g2_nand2_2 _2403_ (.Y(_0276_),
    .A(net916),
    .B(_1364_));
 sg13g2_nor2_2 _2404_ (.A(net910),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_nand4_1 _2405_ (.B(net860),
    .C(net841),
    .A(net874),
    .Y(_0278_),
    .D(_0277_));
 sg13g2_o21ai_1 _2406_ (.B1(net922),
    .Y(_0279_),
    .A1(net847),
    .A2(_0278_));
 sg13g2_nand2_1 _2407_ (.Y(_0280_),
    .A(net810),
    .B(_0279_));
 sg13g2_nor3_2 _2408_ (.A(_0975_),
    .B(_1396_),
    .C(_0276_),
    .Y(_0281_));
 sg13g2_and2_2 _2409_ (.A(_1377_),
    .B(_0281_),
    .X(_0282_));
 sg13g2_nand2_2 _2410_ (.Y(_0283_),
    .A(net876),
    .B(_0282_));
 sg13g2_nor2_2 _2411_ (.A(net905),
    .B(_0283_),
    .Y(_0284_));
 sg13g2_nor2_2 _2412_ (.A(_1360_),
    .B(net796),
    .Y(_0285_));
 sg13g2_a22oi_1 _2413_ (.Y(_0286_),
    .B1(_0284_),
    .B2(net767),
    .A2(_0280_),
    .A1(net337));
 sg13g2_nor2_1 _2414_ (.A(net975),
    .B(net338),
    .Y(_0080_));
 sg13g2_and3_2 _2415_ (.X(_0287_),
    .A(\spi_in.index[1] ),
    .B(net917),
    .C(net915));
 sg13g2_nor2b_2 _2416_ (.A(net910),
    .B_N(_0287_),
    .Y(_0288_));
 sg13g2_nand4_1 _2417_ (.B(net861),
    .C(net845),
    .A(net876),
    .Y(_0289_),
    .D(_0288_));
 sg13g2_o21ai_1 _2418_ (.B1(net922),
    .Y(_0290_),
    .A1(net847),
    .A2(_0289_));
 sg13g2_nand2_1 _2419_ (.Y(_0291_),
    .A(net810),
    .B(_0290_));
 sg13g2_nand2_2 _2420_ (.Y(_0292_),
    .A(net1001),
    .B(_0287_));
 sg13g2_nor4_2 _2421_ (.A(net864),
    .B(net868),
    .C(_0273_),
    .Y(_0293_),
    .D(_0292_));
 sg13g2_a22oi_1 _2422_ (.Y(_0294_),
    .B1(_0293_),
    .B2(net798),
    .A2(_0291_),
    .A1(net410));
 sg13g2_nor2_1 _2423_ (.A(net975),
    .B(_0294_),
    .Y(_0081_));
 sg13g2_nor2_2 _2424_ (.A(net916),
    .B(_1366_),
    .Y(_0295_));
 sg13g2_nor4_2 _2425_ (.A(net914),
    .B(net915),
    .C(_1366_),
    .Y(_0296_),
    .D(_1396_));
 sg13g2_and3_1 _2426_ (.X(_0297_),
    .A(net872),
    .B(net838),
    .C(_0296_));
 sg13g2_nand2_1 _2427_ (.Y(_0298_),
    .A(net859),
    .B(_0297_));
 sg13g2_o21ai_1 _2428_ (.B1(net918),
    .Y(_0299_),
    .A1(net846),
    .A2(_0298_));
 sg13g2_nand2_1 _2429_ (.Y(_0300_),
    .A(net806),
    .B(_0299_));
 sg13g2_and2_1 _2430_ (.A(net1000),
    .B(_0297_),
    .X(_0301_));
 sg13g2_a22oi_1 _2431_ (.Y(_0302_),
    .B1(_0301_),
    .B2(net766),
    .A2(_0300_),
    .A1(net312));
 sg13g2_nor2_1 _2432_ (.A(net970),
    .B(_0302_),
    .Y(_0082_));
 sg13g2_nor2b_2 _2433_ (.A(net916),
    .B_N(_1363_),
    .Y(_0303_));
 sg13g2_nor2b_2 _2434_ (.A(net911),
    .B_N(_0303_),
    .Y(_0304_));
 sg13g2_nand4_1 _2435_ (.B(net860),
    .C(net838),
    .A(net873),
    .Y(_0305_),
    .D(net830));
 sg13g2_o21ai_1 _2436_ (.B1(net920),
    .Y(_0306_),
    .A1(net847),
    .A2(_0305_));
 sg13g2_nand2_1 _2437_ (.Y(_0307_),
    .A(net806),
    .B(_0306_));
 sg13g2_and4_2 _2438_ (.A(net1000),
    .B(net873),
    .C(net838),
    .D(net830),
    .X(_0308_));
 sg13g2_a22oi_1 _2439_ (.Y(_0309_),
    .B1(_0308_),
    .B2(net766),
    .A2(_0307_),
    .A1(net407));
 sg13g2_nor2_1 _2440_ (.A(net970),
    .B(_0309_),
    .Y(_0083_));
 sg13g2_nor2b_2 _2441_ (.A(net915),
    .B_N(_1364_),
    .Y(_0310_));
 sg13g2_nor2b_2 _2442_ (.A(net910),
    .B_N(_0310_),
    .Y(_0311_));
 sg13g2_nand4_1 _2443_ (.B(net859),
    .C(net838),
    .A(net872),
    .Y(_0312_),
    .D(_0311_));
 sg13g2_o21ai_1 _2444_ (.B1(net918),
    .Y(_0313_),
    .A1(net846),
    .A2(_0312_));
 sg13g2_nand2_1 _2445_ (.Y(_0314_),
    .A(net806),
    .B(_0313_));
 sg13g2_nand3b_1 _2446_ (.B(_0310_),
    .C(net1001),
    .Y(_0315_),
    .A_N(_1396_));
 sg13g2_nor2_2 _2447_ (.A(net865),
    .B(_0315_),
    .Y(_0316_));
 sg13g2_nand2_1 _2448_ (.Y(_0317_),
    .A(net874),
    .B(_0316_));
 sg13g2_nor2_2 _2449_ (.A(net905),
    .B(_0317_),
    .Y(_0318_));
 sg13g2_a22oi_1 _2450_ (.Y(_0319_),
    .B1(_0318_),
    .B2(net766),
    .A2(_0314_),
    .A1(net360));
 sg13g2_nor2_1 _2451_ (.A(net971),
    .B(_0319_),
    .Y(_0084_));
 sg13g2_nor2_1 _2452_ (.A(net916),
    .B(_1367_),
    .Y(_0320_));
 sg13g2_nor3_2 _2453_ (.A(net911),
    .B(net915),
    .C(_1367_),
    .Y(_0321_));
 sg13g2_and2_1 _2454_ (.A(net872),
    .B(_0321_),
    .X(_0322_));
 sg13g2_nand3_1 _2455_ (.B(net838),
    .C(_0322_),
    .A(net859),
    .Y(_0323_));
 sg13g2_o21ai_1 _2456_ (.B1(net918),
    .Y(_0324_),
    .A1(net846),
    .A2(_0323_));
 sg13g2_nand2_1 _2457_ (.Y(_0325_),
    .A(net807),
    .B(_0324_));
 sg13g2_and3_1 _2458_ (.X(_0326_),
    .A(net1000),
    .B(net838),
    .C(_0322_));
 sg13g2_a22oi_1 _2459_ (.Y(_0327_),
    .B1(_0326_),
    .B2(net766),
    .A2(_0325_),
    .A1(net376));
 sg13g2_nor2_1 _2460_ (.A(net970),
    .B(_0327_),
    .Y(_0085_));
 sg13g2_nand3_1 _2461_ (.B(_1374_),
    .C(net844),
    .A(net906),
    .Y(_0328_));
 sg13g2_nor2_1 _2462_ (.A(net796),
    .B(_0328_),
    .Y(_0329_));
 sg13g2_o21ai_1 _2463_ (.B1(net828),
    .Y(_0330_),
    .A1(net894),
    .A2(_0329_));
 sg13g2_a22oi_1 _2464_ (.Y(_0331_),
    .B1(_0330_),
    .B2(net259),
    .A2(_0329_),
    .A1(net775));
 sg13g2_nor2_1 _2465_ (.A(net989),
    .B(_0331_),
    .Y(_0086_));
 sg13g2_and2_1 _2466_ (.A(net914),
    .B(_0265_),
    .X(_0332_));
 sg13g2_nand3_1 _2467_ (.B(net844),
    .C(_0332_),
    .A(net906),
    .Y(_0333_));
 sg13g2_or2_1 _2468_ (.X(_0334_),
    .B(_0333_),
    .A(net857));
 sg13g2_o21ai_1 _2469_ (.B1(net927),
    .Y(_0335_),
    .A1(net850),
    .A2(_0334_));
 sg13g2_nand2_1 _2470_ (.Y(_0336_),
    .A(net819),
    .B(_0335_));
 sg13g2_nor4_2 _2471_ (.A(net863),
    .B(net870),
    .C(_0272_),
    .Y(_0337_),
    .D(_0273_));
 sg13g2_a22oi_1 _2472_ (.Y(_0338_),
    .B1(_0337_),
    .B2(net801),
    .A2(_0336_),
    .A1(net443));
 sg13g2_nor2_1 _2473_ (.A(net987),
    .B(_0338_),
    .Y(_0087_));
 sg13g2_and3_1 _2474_ (.X(_0339_),
    .A(net911),
    .B(net915),
    .C(_1364_));
 sg13g2_nand4_1 _2475_ (.B(net862),
    .C(net843),
    .A(net909),
    .Y(_0340_),
    .D(_0339_));
 sg13g2_o21ai_1 _2476_ (.B1(net928),
    .Y(_0341_),
    .A1(net850),
    .A2(_0340_));
 sg13g2_nand2_1 _2477_ (.Y(_0342_),
    .A(net819),
    .B(_0341_));
 sg13g2_nand3_1 _2478_ (.B(net877),
    .C(_0281_),
    .A(net865),
    .Y(_0343_));
 sg13g2_nor2_1 _2479_ (.A(net904),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_a22oi_1 _2480_ (.Y(_0345_),
    .B1(_0344_),
    .B2(net770),
    .A2(_0342_),
    .A1(net451));
 sg13g2_nor2_1 _2481_ (.A(net989),
    .B(_0345_),
    .Y(_0088_));
 sg13g2_and2_1 _2482_ (.A(net914),
    .B(_0287_),
    .X(_0346_));
 sg13g2_nand3_1 _2483_ (.B(net844),
    .C(_0346_),
    .A(net906),
    .Y(_0347_));
 sg13g2_or2_1 _2484_ (.X(_0348_),
    .B(_0347_),
    .A(net857));
 sg13g2_o21ai_1 _2485_ (.B1(net928),
    .Y(_0349_),
    .A1(net850),
    .A2(_0348_));
 sg13g2_nand2_1 _2486_ (.Y(_0350_),
    .A(net819),
    .B(_0349_));
 sg13g2_nor4_2 _2487_ (.A(net863),
    .B(net870),
    .C(_0273_),
    .Y(_0351_),
    .D(_0292_));
 sg13g2_a22oi_1 _2488_ (.Y(_0352_),
    .B1(_0351_),
    .B2(net801),
    .A2(_0350_),
    .A1(net391));
 sg13g2_nor2_1 _2489_ (.A(net989),
    .B(_0352_),
    .Y(_0089_));
 sg13g2_nand2_1 _2490_ (.Y(_0353_),
    .A(net912),
    .B(_0295_));
 sg13g2_nand4_1 _2491_ (.B(net908),
    .C(net843),
    .A(net913),
    .Y(_0354_),
    .D(_0295_));
 sg13g2_or2_1 _2492_ (.X(_0355_),
    .B(_0354_),
    .A(net858));
 sg13g2_o21ai_1 _2493_ (.B1(net933),
    .Y(_0356_),
    .A1(net850),
    .A2(_0355_));
 sg13g2_nand2_1 _2494_ (.Y(_0357_),
    .A(net826),
    .B(_0356_));
 sg13g2_nor2_1 _2495_ (.A(_0975_),
    .B(_0354_),
    .Y(_0358_));
 sg13g2_a22oi_1 _2496_ (.Y(_0359_),
    .B1(_0358_),
    .B2(net770),
    .A2(_0357_),
    .A1(net494));
 sg13g2_nor2_1 _2497_ (.A(net995),
    .B(_0359_),
    .Y(_0090_));
 sg13g2_nand4_1 _2498_ (.B(net907),
    .C(net844),
    .A(net912),
    .Y(_0360_),
    .D(_0303_));
 sg13g2_or2_1 _2499_ (.X(_0361_),
    .B(_0360_),
    .A(net858));
 sg13g2_o21ai_1 _2500_ (.B1(net933),
    .Y(_0362_),
    .A1(net849),
    .A2(_0361_));
 sg13g2_nand2_1 _2501_ (.Y(_0363_),
    .A(net826),
    .B(_0362_));
 sg13g2_nor2_1 _2502_ (.A(_0975_),
    .B(_0360_),
    .Y(_0364_));
 sg13g2_a22oi_1 _2503_ (.Y(_0365_),
    .B1(_0364_),
    .B2(net769),
    .A2(_0363_),
    .A1(net495));
 sg13g2_nor2_1 _2504_ (.A(net994),
    .B(_0365_),
    .Y(_0091_));
 sg13g2_nand4_1 _2505_ (.B(net907),
    .C(net843),
    .A(net912),
    .Y(_0366_),
    .D(_0310_));
 sg13g2_or2_1 _2506_ (.X(_0367_),
    .B(_0366_),
    .A(net858));
 sg13g2_o21ai_1 _2507_ (.B1(net932),
    .Y(_0368_),
    .A1(net849),
    .A2(_0367_));
 sg13g2_nand2_1 _2508_ (.Y(_0369_),
    .A(net822),
    .B(_0368_));
 sg13g2_nor2_2 _2509_ (.A(net863),
    .B(_0315_),
    .Y(_0370_));
 sg13g2_nand2_2 _2510_ (.Y(_0371_),
    .A(net878),
    .B(_0370_));
 sg13g2_nor2_2 _2511_ (.A(net901),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_a22oi_1 _2512_ (.Y(_0373_),
    .B1(_0372_),
    .B2(net769),
    .A2(_0369_),
    .A1(net455));
 sg13g2_nor2_1 _2513_ (.A(net994),
    .B(_0373_),
    .Y(_0092_));
 sg13g2_nand3_1 _2514_ (.B(net907),
    .C(_0320_),
    .A(net913),
    .Y(_0374_));
 sg13g2_nor2_1 _2515_ (.A(net836),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_nand2_1 _2516_ (.Y(_0376_),
    .A(net862),
    .B(_0375_));
 sg13g2_o21ai_1 _2517_ (.B1(net930),
    .Y(_0377_),
    .A1(net849),
    .A2(_0376_));
 sg13g2_nand2_1 _2518_ (.Y(_0378_),
    .A(net828),
    .B(_0377_));
 sg13g2_nor3_2 _2519_ (.A(_0975_),
    .B(net836),
    .C(_0374_),
    .Y(_0379_));
 sg13g2_a22oi_1 _2520_ (.Y(_0380_),
    .B1(_0379_),
    .B2(net769),
    .A2(_0378_),
    .A1(net440));
 sg13g2_nor2_1 _2521_ (.A(net994),
    .B(_0380_),
    .Y(_0093_));
 sg13g2_or4_1 _2522_ (.A(net910),
    .B(_1373_),
    .C(net870),
    .D(_1396_),
    .X(_0381_));
 sg13g2_or2_1 _2523_ (.X(_0382_),
    .B(_0381_),
    .A(net905));
 sg13g2_nor2_1 _2524_ (.A(net795),
    .B(_0382_),
    .Y(_0383_));
 sg13g2_o21ai_1 _2525_ (.B1(net815),
    .Y(_0384_),
    .A1(net893),
    .A2(_0383_));
 sg13g2_a22oi_1 _2526_ (.Y(_0385_),
    .B1(_0384_),
    .B2(net318),
    .A2(_0383_),
    .A1(net773));
 sg13g2_nor2_1 _2527_ (.A(net983),
    .B(_0385_),
    .Y(_0094_));
 sg13g2_nand4_1 _2528_ (.B(net861),
    .C(net842),
    .A(net868),
    .Y(_0386_),
    .D(_0266_));
 sg13g2_o21ai_1 _2529_ (.B1(net924),
    .Y(_0387_),
    .A1(net848),
    .A2(_0386_));
 sg13g2_nand2_1 _2530_ (.Y(_0388_),
    .A(net816),
    .B(_0387_));
 sg13g2_nand2_2 _2531_ (.Y(_0389_),
    .A(net776),
    .B(net844));
 sg13g2_nor4_2 _2532_ (.A(net864),
    .B(net875),
    .C(_0272_),
    .Y(_0390_),
    .D(_0389_));
 sg13g2_a22oi_1 _2533_ (.Y(_0391_),
    .B1(_0390_),
    .B2(net798),
    .A2(_0388_),
    .A1(net354));
 sg13g2_nor2_1 _2534_ (.A(net976),
    .B(_0391_),
    .Y(_0095_));
 sg13g2_nand4_1 _2535_ (.B(net860),
    .C(net840),
    .A(net866),
    .Y(_0392_),
    .D(_0277_));
 sg13g2_o21ai_1 _2536_ (.B1(net921),
    .Y(_0393_),
    .A1(net847),
    .A2(_0392_));
 sg13g2_nand2_1 _2537_ (.Y(_0394_),
    .A(net811),
    .B(_0393_));
 sg13g2_nand2_2 _2538_ (.Y(_0395_),
    .A(net868),
    .B(_0282_));
 sg13g2_nor2_1 _2539_ (.A(net832),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_a22oi_1 _2540_ (.Y(_0397_),
    .B1(_0396_),
    .B2(net767),
    .A2(_0394_),
    .A1(net363));
 sg13g2_nor2_1 _2541_ (.A(net975),
    .B(_0397_),
    .Y(_0096_));
 sg13g2_nand4_1 _2542_ (.B(net860),
    .C(net840),
    .A(net867),
    .Y(_0398_),
    .D(_0288_));
 sg13g2_o21ai_1 _2543_ (.B1(net922),
    .Y(_0399_),
    .A1(net848),
    .A2(_0398_));
 sg13g2_nand2_1 _2544_ (.Y(_0400_),
    .A(net810),
    .B(_0399_));
 sg13g2_nor4_2 _2545_ (.A(net864),
    .B(net876),
    .C(_0292_),
    .Y(_0401_),
    .D(_0389_));
 sg13g2_a22oi_1 _2546_ (.Y(_0402_),
    .B1(_0401_),
    .B2(net798),
    .A2(_0400_),
    .A1(net379));
 sg13g2_nor2_1 _2547_ (.A(net976),
    .B(_0402_),
    .Y(_0097_));
 sg13g2_and3_1 _2548_ (.X(_0403_),
    .A(net866),
    .B(net840),
    .C(_0296_));
 sg13g2_nand2_1 _2549_ (.Y(_0404_),
    .A(net860),
    .B(_0403_));
 sg13g2_o21ai_1 _2550_ (.B1(net921),
    .Y(_0405_),
    .A1(net847),
    .A2(_0404_));
 sg13g2_nand2_1 _2551_ (.Y(_0406_),
    .A(net809),
    .B(_0405_));
 sg13g2_and2_1 _2552_ (.A(net1001),
    .B(_0403_),
    .X(_0407_));
 sg13g2_a22oi_1 _2553_ (.Y(_0408_),
    .B1(_0407_),
    .B2(net767),
    .A2(_0406_),
    .A1(net450));
 sg13g2_nor2_1 _2554_ (.A(net974),
    .B(_0408_),
    .Y(_0098_));
 sg13g2_nand4_1 _2555_ (.B(net860),
    .C(net840),
    .A(net866),
    .Y(_0409_),
    .D(_0304_));
 sg13g2_o21ai_1 _2556_ (.B1(net921),
    .Y(_0410_),
    .A1(net847),
    .A2(_0409_));
 sg13g2_nand2_1 _2557_ (.Y(_0411_),
    .A(net811),
    .B(_0410_));
 sg13g2_and4_2 _2558_ (.A(net1000),
    .B(net866),
    .C(net840),
    .D(net830),
    .X(_0412_));
 sg13g2_a22oi_1 _2559_ (.Y(_0413_),
    .B1(_0412_),
    .B2(net767),
    .A2(_0411_),
    .A1(net460));
 sg13g2_nor2_1 _2560_ (.A(net974),
    .B(_0413_),
    .Y(_0099_));
 sg13g2_nand4_1 _2561_ (.B(net859),
    .C(net839),
    .A(net867),
    .Y(_0414_),
    .D(_0311_));
 sg13g2_o21ai_1 _2562_ (.B1(net920),
    .Y(_0415_),
    .A1(net846),
    .A2(_0414_));
 sg13g2_nand2_1 _2563_ (.Y(_0416_),
    .A(net809),
    .B(_0415_));
 sg13g2_nand2_2 _2564_ (.Y(_0417_),
    .A(net867),
    .B(_0316_));
 sg13g2_nor2_2 _2565_ (.A(net832),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_a22oi_1 _2566_ (.Y(_0419_),
    .B1(_0418_),
    .B2(net767),
    .A2(_0416_),
    .A1(net336));
 sg13g2_nor2_1 _2567_ (.A(net973),
    .B(_0419_),
    .Y(_0100_));
 sg13g2_and3_1 _2568_ (.X(_0420_),
    .A(net866),
    .B(net840),
    .C(_0321_));
 sg13g2_nand2_1 _2569_ (.Y(_0421_),
    .A(net860),
    .B(_0420_));
 sg13g2_o21ai_1 _2570_ (.B1(net921),
    .Y(_0422_),
    .A1(net847),
    .A2(_0421_));
 sg13g2_nand2_1 _2571_ (.Y(_0423_),
    .A(net809),
    .B(_0422_));
 sg13g2_and2_1 _2572_ (.A(net1000),
    .B(_0420_),
    .X(_0424_));
 sg13g2_a22oi_1 _2573_ (.Y(_0425_),
    .B1(_0424_),
    .B2(net767),
    .A2(_0423_),
    .A1(net390));
 sg13g2_nor2_1 _2574_ (.A(net973),
    .B(_0425_),
    .Y(_0101_));
 sg13g2_nor3_2 _2575_ (.A(net904),
    .B(net909),
    .C(_1375_),
    .Y(_0426_));
 sg13g2_and2_1 _2576_ (.A(net862),
    .B(_0426_),
    .X(_0427_));
 sg13g2_a21oi_1 _2577_ (.A1(net854),
    .A2(_0427_),
    .Y(_0428_),
    .B1(net894));
 sg13g2_o21ai_1 _2578_ (.B1(net498),
    .Y(_0429_),
    .A1(net802),
    .A2(_0428_));
 sg13g2_or4_2 _2579_ (.A(_0975_),
    .B(_1375_),
    .C(net878),
    .D(_0389_),
    .X(_0430_));
 sg13g2_o21ai_1 _2580_ (.B1(_0429_),
    .Y(_0431_),
    .A1(net795),
    .A2(_0430_));
 sg13g2_and2_1 _2581_ (.A(net1003),
    .B(_0431_),
    .X(_0102_));
 sg13g2_and3_1 _2582_ (.X(_0432_),
    .A(net911),
    .B(_0976_),
    .C(_0265_));
 sg13g2_nor2b_1 _2583_ (.A(net904),
    .B_N(_0432_),
    .Y(_0433_));
 sg13g2_nand2_1 _2584_ (.Y(_0434_),
    .A(net862),
    .B(_0433_));
 sg13g2_o21ai_1 _2585_ (.B1(net929),
    .Y(_0435_),
    .A1(net850),
    .A2(_0434_));
 sg13g2_nand2_1 _2586_ (.Y(_0436_),
    .A(net818),
    .B(_0435_));
 sg13g2_nor4_2 _2587_ (.A(net863),
    .B(net877),
    .C(_0272_),
    .Y(_0437_),
    .D(_0389_));
 sg13g2_a22oi_1 _2588_ (.Y(_0438_),
    .B1(_0437_),
    .B2(net798),
    .A2(_0436_),
    .A1(net392));
 sg13g2_nor2_1 _2589_ (.A(net985),
    .B(_0438_),
    .Y(_0103_));
 sg13g2_and2_1 _2590_ (.A(_0976_),
    .B(_0339_),
    .X(_0439_));
 sg13g2_nand2b_1 _2591_ (.Y(_0440_),
    .B(_0439_),
    .A_N(net904));
 sg13g2_or2_1 _2592_ (.X(_0441_),
    .B(_0440_),
    .A(net857));
 sg13g2_o21ai_1 _2593_ (.B1(net929),
    .Y(_0442_),
    .A1(net849),
    .A2(_0441_));
 sg13g2_nand2_1 _2594_ (.Y(_0443_),
    .A(net821),
    .B(_0442_));
 sg13g2_nand3_1 _2595_ (.B(net870),
    .C(_0281_),
    .A(net865),
    .Y(_0444_));
 sg13g2_nor2_2 _2596_ (.A(net836),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_a22oi_1 _2597_ (.Y(_0446_),
    .B1(_0445_),
    .B2(net770),
    .A2(_0443_),
    .A1(net425));
 sg13g2_nor2_1 _2598_ (.A(net986),
    .B(_0446_),
    .Y(_0104_));
 sg13g2_and2_1 _2599_ (.A(_0976_),
    .B(_0346_),
    .X(_0447_));
 sg13g2_nand2b_1 _2600_ (.Y(_0448_),
    .B(_0447_),
    .A_N(net904));
 sg13g2_or2_1 _2601_ (.X(_0449_),
    .B(_0448_),
    .A(net857));
 sg13g2_o21ai_1 _2602_ (.B1(net929),
    .Y(_0450_),
    .A1(net850),
    .A2(_0449_));
 sg13g2_nand2_1 _2603_ (.Y(_0451_),
    .A(net818),
    .B(_0450_));
 sg13g2_nor4_2 _2604_ (.A(net863),
    .B(net877),
    .C(_0292_),
    .Y(_0452_),
    .D(_0389_));
 sg13g2_a22oi_1 _2605_ (.Y(_0453_),
    .B1(_0452_),
    .B2(net799),
    .A2(_0451_),
    .A1(net346));
 sg13g2_nor2_1 _2606_ (.A(net986),
    .B(_0453_),
    .Y(_0105_));
 sg13g2_nor2_1 _2607_ (.A(net907),
    .B(_0353_),
    .Y(_0454_));
 sg13g2_nor3_2 _2608_ (.A(net900),
    .B(net907),
    .C(_0353_),
    .Y(_0455_));
 sg13g2_nand2_1 _2609_ (.Y(_0456_),
    .A(net862),
    .B(_0455_));
 sg13g2_o21ai_1 _2610_ (.B1(net930),
    .Y(_0457_),
    .A1(net849),
    .A2(_0456_));
 sg13g2_nand2_1 _2611_ (.Y(_0458_),
    .A(net823),
    .B(_0457_));
 sg13g2_and2_1 _2612_ (.A(net1002),
    .B(_0455_),
    .X(_0459_));
 sg13g2_a22oi_1 _2613_ (.Y(_0460_),
    .B1(_0459_),
    .B2(net769),
    .A2(_0458_),
    .A1(net432));
 sg13g2_nor2_1 _2614_ (.A(net991),
    .B(_0460_),
    .Y(_0106_));
 sg13g2_and3_1 _2615_ (.X(_0461_),
    .A(net912),
    .B(_0976_),
    .C(_0303_));
 sg13g2_nand2b_2 _2616_ (.Y(_0462_),
    .B(_0461_),
    .A_N(net901));
 sg13g2_nor2_1 _2617_ (.A(net796),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_o21ai_1 _2618_ (.B1(net822),
    .Y(_0464_),
    .A1(net896),
    .A2(_0463_));
 sg13g2_a22oi_1 _2619_ (.Y(_0465_),
    .B1(_0464_),
    .B2(net279),
    .A2(_0463_),
    .A1(net774));
 sg13g2_nor2_1 _2620_ (.A(net991),
    .B(_0465_),
    .Y(_0107_));
 sg13g2_and3_1 _2621_ (.X(_0466_),
    .A(net912),
    .B(_0976_),
    .C(_0310_));
 sg13g2_nand2b_1 _2622_ (.Y(_0467_),
    .B(_0466_),
    .A_N(net901));
 sg13g2_or2_1 _2623_ (.X(_0468_),
    .B(_0467_),
    .A(net858));
 sg13g2_o21ai_1 _2624_ (.B1(net930),
    .Y(_0469_),
    .A1(net849),
    .A2(_0468_));
 sg13g2_nand2_1 _2625_ (.Y(_0470_),
    .A(net822),
    .B(_0469_));
 sg13g2_nand2_2 _2626_ (.Y(_0471_),
    .A(net870),
    .B(_0370_));
 sg13g2_nor2_2 _2627_ (.A(net836),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_a22oi_1 _2628_ (.Y(_0473_),
    .B1(_0472_),
    .B2(net769),
    .A2(_0470_),
    .A1(net449));
 sg13g2_nor2_1 _2629_ (.A(net999),
    .B(_0473_),
    .Y(_0108_));
 sg13g2_and3_2 _2630_ (.X(_0474_),
    .A(net911),
    .B(_0976_),
    .C(_0320_));
 sg13g2_nand2b_2 _2631_ (.Y(_0475_),
    .B(_0474_),
    .A_N(net904));
 sg13g2_nor2_1 _2632_ (.A(net795),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_o21ai_1 _2633_ (.B1(net818),
    .Y(_0477_),
    .A1(net894),
    .A2(_0476_));
 sg13g2_a22oi_1 _2634_ (.Y(_0478_),
    .B1(_0477_),
    .B2(net288),
    .A2(_0476_),
    .A1(net772));
 sg13g2_nor2_1 _2635_ (.A(net985),
    .B(_0478_),
    .Y(_0109_));
 sg13g2_nor4_2 _2636_ (.A(net910),
    .B(_1373_),
    .C(net877),
    .Y(_0479_),
    .D(_1396_));
 sg13g2_nand2_1 _2637_ (.Y(_0480_),
    .A(net842),
    .B(_0479_));
 sg13g2_nor2_1 _2638_ (.A(net794),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_o21ai_1 _2639_ (.B1(net813),
    .Y(_0482_),
    .A1(net891),
    .A2(_0481_));
 sg13g2_a22oi_1 _2640_ (.Y(_0483_),
    .B1(_0482_),
    .B2(net252),
    .A2(_0481_),
    .A1(net771));
 sg13g2_nor2_1 _2641_ (.A(net984),
    .B(_0483_),
    .Y(_0110_));
 sg13g2_nand4_1 _2642_ (.B(net861),
    .C(net833),
    .A(net875),
    .Y(_0484_),
    .D(_0266_));
 sg13g2_o21ai_1 _2643_ (.B1(net926),
    .Y(_0485_),
    .A1(net848),
    .A2(_0484_));
 sg13g2_nand2_1 _2644_ (.Y(_0486_),
    .A(net814),
    .B(_0485_));
 sg13g2_nand2_1 _2645_ (.Y(_0487_),
    .A(net776),
    .B(net835));
 sg13g2_nor4_2 _2646_ (.A(net864),
    .B(net869),
    .C(_0272_),
    .Y(_0488_),
    .D(net765));
 sg13g2_a22oi_1 _2647_ (.Y(_0489_),
    .B1(_0488_),
    .B2(net799),
    .A2(_0486_),
    .A1(net400));
 sg13g2_nor2_1 _2648_ (.A(net981),
    .B(_0489_),
    .Y(_0111_));
 sg13g2_nand4_1 _2649_ (.B(net862),
    .C(net833),
    .A(net875),
    .Y(_0490_),
    .D(_0277_));
 sg13g2_o21ai_1 _2650_ (.B1(net926),
    .Y(_0491_),
    .A1(net848),
    .A2(_0490_));
 sg13g2_nand2_1 _2651_ (.Y(_0492_),
    .A(net814),
    .B(_0491_));
 sg13g2_nor2_2 _2652_ (.A(net842),
    .B(_0283_),
    .Y(_0493_));
 sg13g2_a22oi_1 _2653_ (.Y(_0494_),
    .B1(_0493_),
    .B2(net768),
    .A2(_0492_),
    .A1(net335));
 sg13g2_nor2_1 _2654_ (.A(net980),
    .B(_0494_),
    .Y(_0112_));
 sg13g2_nand4_1 _2655_ (.B(net861),
    .C(net833),
    .A(net875),
    .Y(_0495_),
    .D(_0288_));
 sg13g2_o21ai_1 _2656_ (.B1(net926),
    .Y(_0496_),
    .A1(net848),
    .A2(_0495_));
 sg13g2_nand2_1 _2657_ (.Y(_0497_),
    .A(net814),
    .B(_0496_));
 sg13g2_nor4_2 _2658_ (.A(net864),
    .B(net869),
    .C(_0292_),
    .Y(_0498_),
    .D(net765));
 sg13g2_a22oi_1 _2659_ (.Y(_0499_),
    .B1(_0498_),
    .B2(net798),
    .A2(_0497_),
    .A1(net404));
 sg13g2_nor2_1 _2660_ (.A(net979),
    .B(_0499_),
    .Y(_0113_));
 sg13g2_and3_1 _2661_ (.X(_0500_),
    .A(net872),
    .B(net831),
    .C(_0296_));
 sg13g2_nand2_1 _2662_ (.Y(_0501_),
    .A(net859),
    .B(_0500_));
 sg13g2_o21ai_1 _2663_ (.B1(net919),
    .Y(_0502_),
    .A1(net846),
    .A2(_0501_));
 sg13g2_nand2_1 _2664_ (.Y(_0503_),
    .A(net807),
    .B(_0502_));
 sg13g2_and2_1 _2665_ (.A(net1000),
    .B(_0500_),
    .X(_0504_));
 sg13g2_a22oi_1 _2666_ (.Y(_0505_),
    .B1(_0504_),
    .B2(net766),
    .A2(_0503_),
    .A1(net358));
 sg13g2_nor2_1 _2667_ (.A(net971),
    .B(_0505_),
    .Y(_0114_));
 sg13g2_nand4_1 _2668_ (.B(net859),
    .C(net832),
    .A(net873),
    .Y(_0506_),
    .D(net830));
 sg13g2_o21ai_1 _2669_ (.B1(net919),
    .Y(_0507_),
    .A1(net846),
    .A2(_0506_));
 sg13g2_nand2_1 _2670_ (.Y(_0508_),
    .A(net805),
    .B(_0507_));
 sg13g2_and4_2 _2671_ (.A(net1000),
    .B(net872),
    .C(net831),
    .D(net830),
    .X(_0509_));
 sg13g2_a22oi_1 _2672_ (.Y(_0510_),
    .B1(_0509_),
    .B2(net766),
    .A2(_0508_),
    .A1(net328));
 sg13g2_nor2_1 _2673_ (.A(net978),
    .B(_0510_),
    .Y(_0115_));
 sg13g2_nand4_1 _2674_ (.B(net859),
    .C(net831),
    .A(net873),
    .Y(_0511_),
    .D(_0311_));
 sg13g2_o21ai_1 _2675_ (.B1(net919),
    .Y(_0512_),
    .A1(net846),
    .A2(_0511_));
 sg13g2_nand2_1 _2676_ (.Y(_0513_),
    .A(net808),
    .B(_0512_));
 sg13g2_nor2_2 _2677_ (.A(net839),
    .B(_0317_),
    .Y(_0514_));
 sg13g2_a22oi_1 _2678_ (.Y(_0515_),
    .B1(_0514_),
    .B2(net766),
    .A2(_0513_),
    .A1(net368));
 sg13g2_nor2_1 _2679_ (.A(net972),
    .B(_0515_),
    .Y(_0116_));
 sg13g2_nand3_1 _2680_ (.B(net831),
    .C(_0322_),
    .A(net859),
    .Y(_0516_));
 sg13g2_o21ai_1 _2681_ (.B1(net918),
    .Y(_0517_),
    .A1(net846),
    .A2(_0516_));
 sg13g2_nand2_1 _2682_ (.Y(_0518_),
    .A(net805),
    .B(_0517_));
 sg13g2_and3_1 _2683_ (.X(_0519_),
    .A(net1000),
    .B(net831),
    .C(_0322_));
 sg13g2_a22oi_1 _2684_ (.Y(_0520_),
    .B1(_0519_),
    .B2(net766),
    .A2(_0518_),
    .A1(net408));
 sg13g2_nor2_1 _2685_ (.A(net971),
    .B(_0520_),
    .Y(_0117_));
 sg13g2_nand3_1 _2686_ (.B(_1374_),
    .C(net836),
    .A(net906),
    .Y(_0521_));
 sg13g2_nor2_1 _2687_ (.A(net795),
    .B(_0521_),
    .Y(_0522_));
 sg13g2_o21ai_1 _2688_ (.B1(net819),
    .Y(_0523_),
    .A1(net895),
    .A2(_0522_));
 sg13g2_a22oi_1 _2689_ (.Y(_0524_),
    .B1(_0523_),
    .B2(net348),
    .A2(_0522_),
    .A1(net775));
 sg13g2_nor2_1 _2690_ (.A(net987),
    .B(_0524_),
    .Y(_0118_));
 sg13g2_nand3_1 _2691_ (.B(net835),
    .C(_0332_),
    .A(net906),
    .Y(_0525_));
 sg13g2_o21ai_1 _2692_ (.B1(net927),
    .Y(_0526_),
    .A1(net795),
    .A2(_0525_));
 sg13g2_nand2_1 _2693_ (.Y(_0527_),
    .A(net820),
    .B(_0526_));
 sg13g2_nor4_2 _2694_ (.A(net863),
    .B(net870),
    .C(_0272_),
    .Y(_0528_),
    .D(_0487_));
 sg13g2_a22oi_1 _2695_ (.Y(_0529_),
    .B1(_0528_),
    .B2(net798),
    .A2(_0527_),
    .A1(net364));
 sg13g2_nor2_1 _2696_ (.A(net988),
    .B(_0529_),
    .Y(_0119_));
 sg13g2_nand3_1 _2697_ (.B(net835),
    .C(_0339_),
    .A(net906),
    .Y(_0530_));
 sg13g2_o21ai_1 _2698_ (.B1(net928),
    .Y(_0531_),
    .A1(net797),
    .A2(_0530_));
 sg13g2_nand2_1 _2699_ (.Y(_0532_),
    .A(net821),
    .B(_0531_));
 sg13g2_nor2_1 _2700_ (.A(net844),
    .B(_0343_),
    .Y(_0533_));
 sg13g2_a22oi_1 _2701_ (.Y(_0534_),
    .B1(_0533_),
    .B2(net770),
    .A2(_0532_),
    .A1(net464));
 sg13g2_nor2_1 _2702_ (.A(net988),
    .B(_0534_),
    .Y(_0120_));
 sg13g2_nand3_1 _2703_ (.B(net835),
    .C(_0346_),
    .A(net906),
    .Y(_0535_));
 sg13g2_o21ai_1 _2704_ (.B1(net927),
    .Y(_0536_),
    .A1(net797),
    .A2(_0535_));
 sg13g2_nand2_1 _2705_ (.Y(_0537_),
    .A(net820),
    .B(_0536_));
 sg13g2_nor4_2 _2706_ (.A(_1377_),
    .B(net870),
    .C(_0292_),
    .Y(_0538_),
    .D(net765));
 sg13g2_a22oi_1 _2707_ (.Y(_0539_),
    .B1(_0538_),
    .B2(net799),
    .A2(_0537_),
    .A1(net389));
 sg13g2_nor2_1 _2708_ (.A(net987),
    .B(_0539_),
    .Y(_0121_));
 sg13g2_nand4_1 _2709_ (.B(net912),
    .C(net907),
    .A(net900),
    .Y(_0540_),
    .D(_0295_));
 sg13g2_nor2_1 _2710_ (.A(net797),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_o21ai_1 _2711_ (.B1(net823),
    .Y(_0542_),
    .A1(net897),
    .A2(_0541_));
 sg13g2_a22oi_1 _2712_ (.Y(_0543_),
    .B1(_0542_),
    .B2(net403),
    .A2(_0541_),
    .A1(net774));
 sg13g2_nor2_1 _2713_ (.A(net993),
    .B(_0543_),
    .Y(_0122_));
 sg13g2_nand4_1 _2714_ (.B(net912),
    .C(net907),
    .A(net900),
    .Y(_0544_),
    .D(_0303_));
 sg13g2_nor2_1 _2715_ (.A(net796),
    .B(_0544_),
    .Y(_0545_));
 sg13g2_o21ai_1 _2716_ (.B1(net823),
    .Y(_0546_),
    .A1(net896),
    .A2(_0545_));
 sg13g2_a22oi_1 _2717_ (.Y(_0547_),
    .B1(_0546_),
    .B2(net330),
    .A2(_0545_),
    .A1(net774));
 sg13g2_nor2_1 _2718_ (.A(net992),
    .B(_0547_),
    .Y(_0123_));
 sg13g2_nand4_1 _2719_ (.B(net912),
    .C(net907),
    .A(net900),
    .Y(_0548_),
    .D(_0310_));
 sg13g2_o21ai_1 _2720_ (.B1(net931),
    .Y(_0549_),
    .A1(net796),
    .A2(_0548_));
 sg13g2_nand2_1 _2721_ (.Y(_0550_),
    .A(net823),
    .B(_0549_));
 sg13g2_nor2_1 _2722_ (.A(net843),
    .B(_0371_),
    .Y(_0551_));
 sg13g2_a22oi_1 _2723_ (.Y(_0552_),
    .B1(_0551_),
    .B2(net769),
    .A2(_0550_),
    .A1(net486));
 sg13g2_nor2_1 _2724_ (.A(net991),
    .B(_0552_),
    .Y(_0124_));
 sg13g2_nor2_2 _2725_ (.A(net843),
    .B(_0374_),
    .Y(_0553_));
 sg13g2_a21oi_1 _2726_ (.A1(net800),
    .A2(_0553_),
    .Y(_0554_),
    .B1(net896));
 sg13g2_o21ai_1 _2727_ (.B1(net373),
    .Y(_0555_),
    .A1(net803),
    .A2(_0554_));
 sg13g2_nand3_1 _2728_ (.B(net800),
    .C(_0553_),
    .A(net775),
    .Y(_0556_));
 sg13g2_a21oi_1 _2729_ (.A1(_0555_),
    .A2(_0556_),
    .Y(_0125_),
    .B1(net991));
 sg13g2_nand2b_1 _2730_ (.Y(_0557_),
    .B(net835),
    .A_N(_0381_));
 sg13g2_nor2_1 _2731_ (.A(net795),
    .B(_0557_),
    .Y(_0558_));
 sg13g2_o21ai_1 _2732_ (.B1(net816),
    .Y(_0559_),
    .A1(net893),
    .A2(_0558_));
 sg13g2_a22oi_1 _2733_ (.Y(_0560_),
    .B1(_0559_),
    .B2(net251),
    .A2(_0558_),
    .A1(net773));
 sg13g2_nor2_1 _2734_ (.A(net984),
    .B(_0560_),
    .Y(_0126_));
 sg13g2_nand3_1 _2735_ (.B(net834),
    .C(_0266_),
    .A(net868),
    .Y(_0561_));
 sg13g2_o21ai_1 _2736_ (.B1(net925),
    .Y(_0562_),
    .A1(net795),
    .A2(_0561_));
 sg13g2_nand2_1 _2737_ (.Y(_0563_),
    .A(net816),
    .B(_0562_));
 sg13g2_nor4_2 _2738_ (.A(net864),
    .B(net877),
    .C(_0272_),
    .Y(_0564_),
    .D(net765));
 sg13g2_a22oi_1 _2739_ (.Y(_0565_),
    .B1(_0564_),
    .B2(net799),
    .A2(_0563_),
    .A1(net380));
 sg13g2_nor2_1 _2740_ (.A(net983),
    .B(_0565_),
    .Y(_0127_));
 sg13g2_nand3_1 _2741_ (.B(net834),
    .C(_0277_),
    .A(net868),
    .Y(_0566_));
 sg13g2_o21ai_1 _2742_ (.B1(net924),
    .Y(_0567_),
    .A1(net794),
    .A2(_0566_));
 sg13g2_nand2_1 _2743_ (.Y(_0568_),
    .A(net816),
    .B(_0567_));
 sg13g2_nor2_1 _2744_ (.A(net842),
    .B(_0395_),
    .Y(_0569_));
 sg13g2_a22oi_1 _2745_ (.Y(_0570_),
    .B1(_0569_),
    .B2(net768),
    .A2(_0568_),
    .A1(net319));
 sg13g2_nor2_1 _2746_ (.A(net983),
    .B(_0570_),
    .Y(_0128_));
 sg13g2_nand3_1 _2747_ (.B(net834),
    .C(_0288_),
    .A(net868),
    .Y(_0571_));
 sg13g2_o21ai_1 _2748_ (.B1(net925),
    .Y(_0572_),
    .A1(net794),
    .A2(_0571_));
 sg13g2_nand2_1 _2749_ (.Y(_0573_),
    .A(net817),
    .B(_0572_));
 sg13g2_nor4_2 _2750_ (.A(net864),
    .B(net876),
    .C(_0292_),
    .Y(_0574_),
    .D(net765));
 sg13g2_a22oi_1 _2751_ (.Y(_0575_),
    .B1(_0574_),
    .B2(net798),
    .A2(_0573_),
    .A1(net367));
 sg13g2_nor2_1 _2752_ (.A(net984),
    .B(_0575_),
    .Y(_0129_));
 sg13g2_nand3_1 _2753_ (.B(net833),
    .C(_0296_),
    .A(net869),
    .Y(_0576_));
 sg13g2_nor2_1 _2754_ (.A(net794),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_o21ai_1 _2755_ (.B1(net813),
    .Y(_0578_),
    .A1(net892),
    .A2(_0577_));
 sg13g2_a22oi_1 _2756_ (.Y(_0579_),
    .B1(_0578_),
    .B2(net265),
    .A2(_0577_),
    .A1(net771));
 sg13g2_nor2_1 _2757_ (.A(net981),
    .B(_0579_),
    .Y(_0130_));
 sg13g2_nand3_1 _2758_ (.B(net835),
    .C(_0304_),
    .A(net870),
    .Y(_0580_));
 sg13g2_nor2_1 _2759_ (.A(net794),
    .B(_0580_),
    .Y(_0581_));
 sg13g2_o21ai_1 _2760_ (.B1(net813),
    .Y(_0582_),
    .A1(net892),
    .A2(_0581_));
 sg13g2_a22oi_1 _2761_ (.Y(_0583_),
    .B1(_0582_),
    .B2(net272),
    .A2(_0581_),
    .A1(net772));
 sg13g2_nor2_1 _2762_ (.A(net981),
    .B(_0583_),
    .Y(_0131_));
 sg13g2_nand3_1 _2763_ (.B(net833),
    .C(_0311_),
    .A(net869),
    .Y(_0584_));
 sg13g2_o21ai_1 _2764_ (.B1(net926),
    .Y(_0585_),
    .A1(net794),
    .A2(_0584_));
 sg13g2_nand2_1 _2765_ (.Y(_0586_),
    .A(net812),
    .B(_0585_));
 sg13g2_nor2_1 _2766_ (.A(net842),
    .B(_0417_),
    .Y(_0587_));
 sg13g2_a22oi_1 _2767_ (.Y(_0588_),
    .B1(_0587_),
    .B2(net768),
    .A2(_0586_),
    .A1(net416));
 sg13g2_nor2_1 _2768_ (.A(net979),
    .B(_0588_),
    .Y(_0132_));
 sg13g2_nand3_1 _2769_ (.B(net835),
    .C(_0321_),
    .A(net869),
    .Y(_0589_));
 sg13g2_nor2_1 _2770_ (.A(net794),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_o21ai_1 _2771_ (.B1(net813),
    .Y(_0591_),
    .A1(net892),
    .A2(_0590_));
 sg13g2_a22oi_1 _2772_ (.Y(_0592_),
    .B1(_0591_),
    .B2(net323),
    .A2(_0590_),
    .A1(net772));
 sg13g2_nor2_1 _2773_ (.A(net981),
    .B(_0592_),
    .Y(_0133_));
 sg13g2_nand3_1 _2774_ (.B(_0976_),
    .C(_1374_),
    .A(net902),
    .Y(_0593_));
 sg13g2_o21ai_1 _2775_ (.B1(net934),
    .Y(_0594_),
    .A1(net796),
    .A2(_0593_));
 sg13g2_nand2_1 _2776_ (.Y(_0595_),
    .A(net827),
    .B(_0594_));
 sg13g2_nor4_2 _2777_ (.A(_0975_),
    .B(_1375_),
    .C(net877),
    .Y(_0596_),
    .D(net765));
 sg13g2_a22oi_1 _2778_ (.Y(_0597_),
    .B1(_0596_),
    .B2(net801),
    .A2(_0595_),
    .A1(net396));
 sg13g2_nor2_1 _2779_ (.A(net996),
    .B(_0597_),
    .Y(_0134_));
 sg13g2_nand2_1 _2780_ (.Y(_0598_),
    .A(net903),
    .B(_0432_));
 sg13g2_o21ai_1 _2781_ (.B1(net933),
    .Y(_0599_),
    .A1(net796),
    .A2(_0598_));
 sg13g2_nand2_1 _2782_ (.Y(_0600_),
    .A(net827),
    .B(_0599_));
 sg13g2_nor4_2 _2783_ (.A(net863),
    .B(net877),
    .C(_0272_),
    .Y(_0601_),
    .D(net765));
 sg13g2_a22oi_1 _2784_ (.Y(_0602_),
    .B1(_0601_),
    .B2(net801),
    .A2(_0600_),
    .A1(net361));
 sg13g2_nor2_1 _2785_ (.A(net996),
    .B(_0602_),
    .Y(_0135_));
 sg13g2_and3_1 _2786_ (.X(_0603_),
    .A(net902),
    .B(net801),
    .C(_0439_));
 sg13g2_o21ai_1 _2787_ (.B1(net826),
    .Y(_0604_),
    .A1(net897),
    .A2(_0603_));
 sg13g2_nor2_2 _2788_ (.A(net843),
    .B(_0444_),
    .Y(_0605_));
 sg13g2_a22oi_1 _2789_ (.Y(_0606_),
    .B1(_0605_),
    .B2(net769),
    .A2(_0604_),
    .A1(net427));
 sg13g2_nor2_1 _2790_ (.A(net995),
    .B(_0606_),
    .Y(_0136_));
 sg13g2_and3_1 _2791_ (.X(_0607_),
    .A(net903),
    .B(net800),
    .C(_0447_));
 sg13g2_o21ai_1 _2792_ (.B1(net827),
    .Y(_0608_),
    .A1(net898),
    .A2(_0607_));
 sg13g2_nor4_2 _2793_ (.A(net863),
    .B(net877),
    .C(_0292_),
    .Y(_0609_),
    .D(net765));
 sg13g2_a22oi_1 _2794_ (.Y(_0610_),
    .B1(_0609_),
    .B2(net800),
    .A2(_0608_),
    .A1(net421));
 sg13g2_nor2_1 _2795_ (.A(net996),
    .B(_0610_),
    .Y(_0137_));
 sg13g2_nand3_1 _2796_ (.B(net800),
    .C(_0454_),
    .A(net901),
    .Y(_0611_));
 sg13g2_a21oi_1 _2797_ (.A1(net931),
    .A2(_0611_),
    .Y(_0612_),
    .B1(net802));
 sg13g2_nand2b_1 _2798_ (.Y(_0613_),
    .B(net508),
    .A_N(_0612_));
 sg13g2_o21ai_1 _2799_ (.B1(_0613_),
    .Y(_0614_),
    .A1(_0263_),
    .A2(_0611_));
 sg13g2_and2_1 _2800_ (.A(net1006),
    .B(_0614_),
    .X(_0138_));
 sg13g2_nand2_1 _2801_ (.Y(_0615_),
    .A(net900),
    .B(_0461_));
 sg13g2_o21ai_1 _2802_ (.B1(net931),
    .Y(_0616_),
    .A1(net797),
    .A2(_0615_));
 sg13g2_nand2_1 _2803_ (.Y(_0617_),
    .A(net824),
    .B(_0616_));
 sg13g2_nor2_1 _2804_ (.A(_0263_),
    .B(_0615_),
    .Y(_0618_));
 sg13g2_a22oi_1 _2805_ (.Y(_0619_),
    .B1(_0618_),
    .B2(net800),
    .A2(_0617_),
    .A1(net383));
 sg13g2_nor2_1 _2806_ (.A(net992),
    .B(_0619_),
    .Y(_0139_));
 sg13g2_nand3_1 _2807_ (.B(net800),
    .C(_0466_),
    .A(net900),
    .Y(_0620_));
 sg13g2_a21o_1 _2808_ (.A2(_0620_),
    .A1(net932),
    .B1(net803),
    .X(_0621_));
 sg13g2_nor2_2 _2809_ (.A(net843),
    .B(_0471_),
    .Y(_0622_));
 sg13g2_a22oi_1 _2810_ (.Y(_0623_),
    .B1(_0622_),
    .B2(net769),
    .A2(_0621_),
    .A1(net405));
 sg13g2_nor2_1 _2811_ (.A(net992),
    .B(_0623_),
    .Y(_0140_));
 sg13g2_nand2_1 _2812_ (.Y(_0624_),
    .A(net900),
    .B(_0474_));
 sg13g2_o21ai_1 _2813_ (.B1(net932),
    .Y(_0625_),
    .A1(net796),
    .A2(_0624_));
 sg13g2_nand2_1 _2814_ (.Y(_0626_),
    .A(net824),
    .B(_0625_));
 sg13g2_nor2_1 _2815_ (.A(_0263_),
    .B(_0624_),
    .Y(_0627_));
 sg13g2_a22oi_1 _2816_ (.Y(_0628_),
    .B1(_0627_),
    .B2(net800),
    .A2(_0626_),
    .A1(net406));
 sg13g2_nor2_1 _2817_ (.A(net992),
    .B(_0628_),
    .Y(_0141_));
 sg13g2_nand2_1 _2818_ (.Y(_0629_),
    .A(net833),
    .B(_0479_));
 sg13g2_nor2_1 _2819_ (.A(net794),
    .B(_0629_),
    .Y(_0630_));
 sg13g2_o21ai_1 _2820_ (.B1(net812),
    .Y(_0631_),
    .A1(net889),
    .A2(_0630_));
 sg13g2_a22oi_1 _2821_ (.Y(_0632_),
    .B1(_0631_),
    .B2(net276),
    .A2(_0630_),
    .A1(net771));
 sg13g2_nor2_1 _2822_ (.A(net972),
    .B(_0632_),
    .Y(_0142_));
 sg13g2_nor2_1 _2823_ (.A(net861),
    .B(net848),
    .Y(_0633_));
 sg13g2_nand2_1 _2824_ (.Y(_0634_),
    .A(net857),
    .B(net855));
 sg13g2_and4_1 _2825_ (.A(net876),
    .B(net842),
    .C(_0266_),
    .D(net789),
    .X(_0635_));
 sg13g2_o21ai_1 _2826_ (.B1(net815),
    .Y(_0636_),
    .A1(net899),
    .A2(_0635_));
 sg13g2_a22oi_1 _2827_ (.Y(_0637_),
    .B1(_0636_),
    .B2(net342),
    .A2(net789),
    .A1(_0274_));
 sg13g2_nor2_1 _2828_ (.A(net982),
    .B(_0637_),
    .Y(_0143_));
 sg13g2_and4_1 _2829_ (.A(net874),
    .B(net839),
    .C(_0277_),
    .D(net785),
    .X(_0638_));
 sg13g2_o21ai_1 _2830_ (.B1(net808),
    .Y(_0639_),
    .A1(net888),
    .A2(_0638_));
 sg13g2_nor2_2 _2831_ (.A(_1360_),
    .B(net783),
    .Y(_0640_));
 sg13g2_a22oi_1 _2832_ (.Y(_0641_),
    .B1(net761),
    .B2(_0284_),
    .A2(_0639_),
    .A1(net352));
 sg13g2_nor2_1 _2833_ (.A(net975),
    .B(net353),
    .Y(_0144_));
 sg13g2_and4_1 _2834_ (.A(net874),
    .B(net839),
    .C(_0288_),
    .D(net787),
    .X(_0642_));
 sg13g2_o21ai_1 _2835_ (.B1(net810),
    .Y(_0643_),
    .A1(net889),
    .A2(_0642_));
 sg13g2_a22oi_1 _2836_ (.Y(_0644_),
    .B1(_0643_),
    .B2(net270),
    .A2(net786),
    .A1(_0293_));
 sg13g2_nor2_1 _2837_ (.A(net975),
    .B(_0644_),
    .Y(_0145_));
 sg13g2_a21oi_1 _2838_ (.A1(_0297_),
    .A2(net785),
    .Y(_0645_),
    .B1(net888));
 sg13g2_o21ai_1 _2839_ (.B1(net347),
    .Y(_0646_),
    .A1(net804),
    .A2(_0645_));
 sg13g2_nand2_1 _2840_ (.Y(_0647_),
    .A(_0301_),
    .B(net760));
 sg13g2_a21oi_1 _2841_ (.A1(_0646_),
    .A2(_0647_),
    .Y(_0146_),
    .B1(net972));
 sg13g2_and4_1 _2842_ (.A(net873),
    .B(net839),
    .C(net830),
    .D(net787),
    .X(_0648_));
 sg13g2_o21ai_1 _2843_ (.B1(net806),
    .Y(_0649_),
    .A1(net889),
    .A2(_0648_));
 sg13g2_a22oi_1 _2844_ (.Y(_0650_),
    .B1(_0649_),
    .B2(net382),
    .A2(net760),
    .A1(_0308_));
 sg13g2_nor2_1 _2845_ (.A(net973),
    .B(_0650_),
    .Y(_0147_));
 sg13g2_and4_1 _2846_ (.A(net872),
    .B(net838),
    .C(_0311_),
    .D(net785),
    .X(_0651_));
 sg13g2_o21ai_1 _2847_ (.B1(net808),
    .Y(_0652_),
    .A1(net888),
    .A2(_0651_));
 sg13g2_a22oi_1 _2848_ (.Y(_0653_),
    .B1(_0652_),
    .B2(net290),
    .A2(net760),
    .A1(_0318_));
 sg13g2_nor2_1 _2849_ (.A(net972),
    .B(_0653_),
    .Y(_0148_));
 sg13g2_and3_1 _2850_ (.X(_0654_),
    .A(net838),
    .B(_0322_),
    .C(net785));
 sg13g2_o21ai_1 _2851_ (.B1(net806),
    .Y(_0655_),
    .A1(net889),
    .A2(_0654_));
 sg13g2_a22oi_1 _2852_ (.Y(_0656_),
    .B1(_0655_),
    .B2(net378),
    .A2(net760),
    .A1(_0326_));
 sg13g2_nor2_1 _2853_ (.A(net970),
    .B(_0656_),
    .Y(_0149_));
 sg13g2_nor2_1 _2854_ (.A(_0328_),
    .B(net783),
    .Y(_0657_));
 sg13g2_o21ai_1 _2855_ (.B1(net819),
    .Y(_0658_),
    .A1(net895),
    .A2(_0657_));
 sg13g2_a22oi_1 _2856_ (.Y(_0659_),
    .B1(_0658_),
    .B2(net273),
    .A2(_0657_),
    .A1(net775));
 sg13g2_nor2_1 _2857_ (.A(net989),
    .B(_0659_),
    .Y(_0150_));
 sg13g2_o21ai_1 _2858_ (.B1(net927),
    .Y(_0660_),
    .A1(_0333_),
    .A2(net780));
 sg13g2_nand2_1 _2859_ (.Y(_0661_),
    .A(net819),
    .B(_0660_));
 sg13g2_a22oi_1 _2860_ (.Y(_0662_),
    .B1(_0661_),
    .B2(net271),
    .A2(net793),
    .A1(_0337_));
 sg13g2_nor2_1 _2861_ (.A(net990),
    .B(_0662_),
    .Y(_0151_));
 sg13g2_and4_1 _2862_ (.A(net906),
    .B(net843),
    .C(_0339_),
    .D(net790),
    .X(_0663_));
 sg13g2_o21ai_1 _2863_ (.B1(net819),
    .Y(_0664_),
    .A1(net895),
    .A2(_0663_));
 sg13g2_a22oi_1 _2864_ (.Y(_0665_),
    .B1(_0664_),
    .B2(net267),
    .A2(net764),
    .A1(_0344_));
 sg13g2_nor2_1 _2865_ (.A(net989),
    .B(_0665_),
    .Y(_0152_));
 sg13g2_o21ai_1 _2866_ (.B1(net928),
    .Y(_0666_),
    .A1(_0347_),
    .A2(net783));
 sg13g2_nand2_1 _2867_ (.Y(_0667_),
    .A(net821),
    .B(_0666_));
 sg13g2_a22oi_1 _2868_ (.Y(_0668_),
    .B1(_0667_),
    .B2(net291),
    .A2(net790),
    .A1(_0351_));
 sg13g2_nor2_1 _2869_ (.A(net989),
    .B(_0668_),
    .Y(_0153_));
 sg13g2_o21ai_1 _2870_ (.B1(net933),
    .Y(_0669_),
    .A1(_0354_),
    .A2(net782));
 sg13g2_nand2_1 _2871_ (.Y(_0670_),
    .A(net826),
    .B(_0669_));
 sg13g2_a22oi_1 _2872_ (.Y(_0671_),
    .B1(_0670_),
    .B2(net339),
    .A2(net763),
    .A1(_0358_));
 sg13g2_nor2_1 _2873_ (.A(net995),
    .B(_0671_),
    .Y(_0154_));
 sg13g2_o21ai_1 _2874_ (.B1(net933),
    .Y(_0672_),
    .A1(_0360_),
    .A2(net782));
 sg13g2_nand2_1 _2875_ (.Y(_0673_),
    .A(net826),
    .B(_0672_));
 sg13g2_a22oi_1 _2876_ (.Y(_0674_),
    .B1(_0673_),
    .B2(net412),
    .A2(net763),
    .A1(_0364_));
 sg13g2_nor2_1 _2877_ (.A(net995),
    .B(_0674_),
    .Y(_0155_));
 sg13g2_o21ai_1 _2878_ (.B1(net930),
    .Y(_0675_),
    .A1(_0366_),
    .A2(net781));
 sg13g2_nand2_1 _2879_ (.Y(_0676_),
    .A(net825),
    .B(_0675_));
 sg13g2_a22oi_1 _2880_ (.Y(_0677_),
    .B1(_0676_),
    .B2(net334),
    .A2(net763),
    .A1(_0372_));
 sg13g2_nor2_1 _2881_ (.A(net994),
    .B(_0677_),
    .Y(_0156_));
 sg13g2_a21oi_1 _2882_ (.A1(_0375_),
    .A2(net792),
    .Y(_0678_),
    .B1(net896));
 sg13g2_o21ai_1 _2883_ (.B1(net362),
    .Y(_0679_),
    .A1(net802),
    .A2(_0678_));
 sg13g2_nand2_1 _2884_ (.Y(_0680_),
    .A(_0379_),
    .B(net764));
 sg13g2_a21oi_1 _2885_ (.A1(_0679_),
    .A2(_0680_),
    .Y(_0157_),
    .B1(net994));
 sg13g2_nand2b_1 _2886_ (.Y(_0681_),
    .B(net788),
    .A_N(_0382_));
 sg13g2_a22oi_1 _2887_ (.Y(_0682_),
    .B1(net776),
    .B2(_0681_),
    .A2(net804),
    .A1(net483));
 sg13g2_a221oi_1 _2888_ (.B2(_0263_),
    .C1(net983),
    .B1(_0682_),
    .A1(_0952_),
    .Y(_0158_),
    .A2(_0681_));
 sg13g2_and4_1 _2889_ (.A(net868),
    .B(net842),
    .C(_0266_),
    .D(net789),
    .X(_0683_));
 sg13g2_o21ai_1 _2890_ (.B1(net816),
    .Y(_0684_),
    .A1(net893),
    .A2(_0683_));
 sg13g2_a22oi_1 _2891_ (.Y(_0685_),
    .B1(_0684_),
    .B2(net257),
    .A2(net786),
    .A1(_0390_));
 sg13g2_nor2_1 _2892_ (.A(net982),
    .B(_0685_),
    .Y(_0159_));
 sg13g2_and4_1 _2893_ (.A(net866),
    .B(net840),
    .C(_0277_),
    .D(net786),
    .X(_0686_));
 sg13g2_o21ai_1 _2894_ (.B1(net810),
    .Y(_0687_),
    .A1(net890),
    .A2(_0686_));
 sg13g2_a22oi_1 _2895_ (.Y(_0688_),
    .B1(_0687_),
    .B2(net326),
    .A2(net761),
    .A1(_0396_));
 sg13g2_nor2_1 _2896_ (.A(net976),
    .B(_0688_),
    .Y(_0160_));
 sg13g2_and4_1 _2897_ (.A(net866),
    .B(net841),
    .C(_0288_),
    .D(net786),
    .X(_0689_));
 sg13g2_o21ai_1 _2898_ (.B1(net810),
    .Y(_0690_),
    .A1(net890),
    .A2(_0689_));
 sg13g2_a22oi_1 _2899_ (.Y(_0691_),
    .B1(_0690_),
    .B2(net324),
    .A2(net786),
    .A1(_0401_));
 sg13g2_nor2_1 _2900_ (.A(net976),
    .B(_0691_),
    .Y(_0161_));
 sg13g2_a21oi_1 _2901_ (.A1(_0403_),
    .A2(net786),
    .Y(_0692_),
    .B1(net890));
 sg13g2_o21ai_1 _2902_ (.B1(net433),
    .Y(_0693_),
    .A1(net804),
    .A2(_0692_));
 sg13g2_nand2_1 _2903_ (.Y(_0694_),
    .A(_0407_),
    .B(net761));
 sg13g2_a21oi_1 _2904_ (.A1(_0693_),
    .A2(_0694_),
    .Y(_0162_),
    .B1(net974));
 sg13g2_and4_1 _2905_ (.A(net866),
    .B(net840),
    .C(net830),
    .D(net786),
    .X(_0695_));
 sg13g2_o21ai_1 _2906_ (.B1(net809),
    .Y(_0696_),
    .A1(net890),
    .A2(_0695_));
 sg13g2_a22oi_1 _2907_ (.Y(_0697_),
    .B1(_0696_),
    .B2(net314),
    .A2(net761),
    .A1(_0412_));
 sg13g2_nor2_1 _2908_ (.A(net974),
    .B(_0697_),
    .Y(_0163_));
 sg13g2_and4_1 _2909_ (.A(net867),
    .B(net839),
    .C(_0311_),
    .D(net787),
    .X(_0698_));
 sg13g2_o21ai_1 _2910_ (.B1(net807),
    .Y(_0699_),
    .A1(net888),
    .A2(_0698_));
 sg13g2_a22oi_1 _2911_ (.Y(_0700_),
    .B1(_0699_),
    .B2(net397),
    .A2(net761),
    .A1(_0418_));
 sg13g2_nor2_1 _2912_ (.A(net973),
    .B(_0700_),
    .Y(_0164_));
 sg13g2_a21oi_1 _2913_ (.A1(_0420_),
    .A2(net786),
    .Y(_0701_),
    .B1(net890));
 sg13g2_o21ai_1 _2914_ (.B1(net377),
    .Y(_0702_),
    .A1(net804),
    .A2(_0701_));
 sg13g2_nand2_1 _2915_ (.Y(_0703_),
    .A(_0424_),
    .B(net761));
 sg13g2_a21oi_1 _2916_ (.A1(_0702_),
    .A2(_0703_),
    .Y(_0165_),
    .B1(net973));
 sg13g2_a21oi_1 _2917_ (.A1(_0426_),
    .A2(net790),
    .Y(_0704_),
    .B1(net894));
 sg13g2_o21ai_1 _2918_ (.B1(net502),
    .Y(_0705_),
    .A1(net802),
    .A2(_0704_));
 sg13g2_o21ai_1 _2919_ (.B1(_0705_),
    .Y(_0706_),
    .A1(_0430_),
    .A2(net783));
 sg13g2_and2_1 _2920_ (.A(net1003),
    .B(_0706_),
    .X(_0166_));
 sg13g2_a21oi_1 _2921_ (.A1(_0433_),
    .A2(net790),
    .Y(_0707_),
    .B1(net894));
 sg13g2_o21ai_1 _2922_ (.B1(net393),
    .Y(_0708_),
    .A1(net802),
    .A2(_0707_));
 sg13g2_nand2_1 _2923_ (.Y(_0709_),
    .A(_0437_),
    .B(net790));
 sg13g2_a21oi_1 _2924_ (.A1(_0708_),
    .A2(_0709_),
    .Y(_0167_),
    .B1(net985));
 sg13g2_o21ai_1 _2925_ (.B1(net929),
    .Y(_0710_),
    .A1(_0440_),
    .A2(net783));
 sg13g2_nand2_1 _2926_ (.Y(_0711_),
    .A(net822),
    .B(_0710_));
 sg13g2_a22oi_1 _2927_ (.Y(_0712_),
    .B1(_0711_),
    .B2(net299),
    .A2(net764),
    .A1(_0445_));
 sg13g2_nor2_1 _2928_ (.A(net986),
    .B(_0712_),
    .Y(_0168_));
 sg13g2_o21ai_1 _2929_ (.B1(net929),
    .Y(_0713_),
    .A1(_0448_),
    .A2(net784));
 sg13g2_nand2_1 _2930_ (.Y(_0714_),
    .A(net821),
    .B(_0713_));
 sg13g2_a22oi_1 _2931_ (.Y(_0715_),
    .B1(_0714_),
    .B2(net293),
    .A2(net790),
    .A1(_0452_));
 sg13g2_nor2_1 _2932_ (.A(net985),
    .B(_0715_),
    .Y(_0169_));
 sg13g2_a21oi_1 _2933_ (.A1(_0455_),
    .A2(net791),
    .Y(_0716_),
    .B1(net896));
 sg13g2_o21ai_1 _2934_ (.B1(net417),
    .Y(_0717_),
    .A1(net803),
    .A2(_0716_));
 sg13g2_nand2_1 _2935_ (.Y(_0718_),
    .A(_0459_),
    .B(net763));
 sg13g2_a21oi_1 _2936_ (.A1(_0717_),
    .A2(_0718_),
    .Y(_0170_),
    .B1(net991));
 sg13g2_nor2_1 _2937_ (.A(_0462_),
    .B(net781),
    .Y(_0719_));
 sg13g2_o21ai_1 _2938_ (.B1(net822),
    .Y(_0720_),
    .A1(net896),
    .A2(_0719_));
 sg13g2_a22oi_1 _2939_ (.Y(_0721_),
    .B1(_0720_),
    .B2(net420),
    .A2(_0719_),
    .A1(net774));
 sg13g2_nor2_1 _2940_ (.A(net991),
    .B(_0721_),
    .Y(_0171_));
 sg13g2_o21ai_1 _2941_ (.B1(net930),
    .Y(_0722_),
    .A1(_0467_),
    .A2(net781));
 sg13g2_nand2_1 _2942_ (.Y(_0723_),
    .A(net822),
    .B(_0722_));
 sg13g2_a22oi_1 _2943_ (.Y(_0724_),
    .B1(_0723_),
    .B2(net375),
    .A2(net763),
    .A1(_0472_));
 sg13g2_nor2_1 _2944_ (.A(net998),
    .B(_0724_),
    .Y(_0172_));
 sg13g2_nor2_1 _2945_ (.A(_0475_),
    .B(net780),
    .Y(_0725_));
 sg13g2_o21ai_1 _2946_ (.B1(net818),
    .Y(_0726_),
    .A1(net894),
    .A2(_0725_));
 sg13g2_a22oi_1 _2947_ (.Y(_0727_),
    .B1(_0726_),
    .B2(net275),
    .A2(_0725_),
    .A1(net772));
 sg13g2_nor2_1 _2948_ (.A(net985),
    .B(_0727_),
    .Y(_0173_));
 sg13g2_nor2_1 _2949_ (.A(_0480_),
    .B(net779),
    .Y(_0728_));
 sg13g2_o21ai_1 _2950_ (.B1(net812),
    .Y(_0729_),
    .A1(net891),
    .A2(_0728_));
 sg13g2_a22oi_1 _2951_ (.Y(_0730_),
    .B1(_0729_),
    .B2(net289),
    .A2(_0728_),
    .A1(net771));
 sg13g2_nor2_1 _2952_ (.A(net979),
    .B(_0730_),
    .Y(_0174_));
 sg13g2_and4_1 _2953_ (.A(net875),
    .B(net834),
    .C(_0266_),
    .D(net788),
    .X(_0731_));
 sg13g2_o21ai_1 _2954_ (.B1(net814),
    .Y(_0732_),
    .A1(net891),
    .A2(_0731_));
 sg13g2_a22oi_1 _2955_ (.Y(_0733_),
    .B1(_0732_),
    .B2(net322),
    .A2(net788),
    .A1(_0488_));
 sg13g2_nor2_1 _2956_ (.A(net984),
    .B(_0733_),
    .Y(_0175_));
 sg13g2_and4_1 _2957_ (.A(net875),
    .B(net833),
    .C(_0277_),
    .D(net788),
    .X(_0734_));
 sg13g2_o21ai_1 _2958_ (.B1(net812),
    .Y(_0735_),
    .A1(net891),
    .A2(_0734_));
 sg13g2_a22oi_1 _2959_ (.Y(_0736_),
    .B1(_0735_),
    .B2(net325),
    .A2(net762),
    .A1(_0493_));
 sg13g2_nor2_1 _2960_ (.A(net980),
    .B(_0736_),
    .Y(_0176_));
 sg13g2_and4_1 _2961_ (.A(net875),
    .B(net833),
    .C(_0288_),
    .D(net788),
    .X(_0737_));
 sg13g2_o21ai_1 _2962_ (.B1(net814),
    .Y(_0738_),
    .A1(net891),
    .A2(_0737_));
 sg13g2_a22oi_1 _2963_ (.Y(_0739_),
    .B1(_0738_),
    .B2(net264),
    .A2(net788),
    .A1(_0498_));
 sg13g2_nor2_1 _2964_ (.A(net979),
    .B(_0739_),
    .Y(_0177_));
 sg13g2_a21oi_1 _2965_ (.A1(_0500_),
    .A2(net785),
    .Y(_0740_),
    .B1(net888));
 sg13g2_o21ai_1 _2966_ (.B1(net329),
    .Y(_0741_),
    .A1(net804),
    .A2(_0740_));
 sg13g2_nand2_1 _2967_ (.Y(_0742_),
    .A(_0504_),
    .B(net760));
 sg13g2_a21oi_1 _2968_ (.A1(_0741_),
    .A2(_0742_),
    .Y(_0178_),
    .B1(net971));
 sg13g2_and4_1 _2969_ (.A(net872),
    .B(net831),
    .C(net830),
    .D(net785),
    .X(_0743_));
 sg13g2_o21ai_1 _2970_ (.B1(net805),
    .Y(_0744_),
    .A1(net888),
    .A2(_0743_));
 sg13g2_a22oi_1 _2971_ (.Y(_0745_),
    .B1(_0744_),
    .B2(net274),
    .A2(net760),
    .A1(_0509_));
 sg13g2_nor2_1 _2972_ (.A(net971),
    .B(_0745_),
    .Y(_0179_));
 sg13g2_and4_1 _2973_ (.A(net872),
    .B(net831),
    .C(_0311_),
    .D(net785),
    .X(_0746_));
 sg13g2_o21ai_1 _2974_ (.B1(net805),
    .Y(_0747_),
    .A1(net888),
    .A2(_0746_));
 sg13g2_a22oi_1 _2975_ (.Y(_0748_),
    .B1(_0747_),
    .B2(net255),
    .A2(net760),
    .A1(_0514_));
 sg13g2_nor2_1 _2976_ (.A(net971),
    .B(_0748_),
    .Y(_0180_));
 sg13g2_and3_1 _2977_ (.X(_0749_),
    .A(net831),
    .B(_0322_),
    .C(net785));
 sg13g2_o21ai_1 _2978_ (.B1(net805),
    .Y(_0750_),
    .A1(net888),
    .A2(_0749_));
 sg13g2_a22oi_1 _2979_ (.Y(_0751_),
    .B1(_0750_),
    .B2(net310),
    .A2(net760),
    .A1(_0519_));
 sg13g2_nor2_1 _2980_ (.A(net971),
    .B(_0751_),
    .Y(_0181_));
 sg13g2_nor2_1 _2981_ (.A(_0521_),
    .B(net780),
    .Y(_0752_));
 sg13g2_o21ai_1 _2982_ (.B1(net820),
    .Y(_0753_),
    .A1(net895),
    .A2(_0752_));
 sg13g2_a22oi_1 _2983_ (.Y(_0754_),
    .B1(_0753_),
    .B2(net256),
    .A2(_0752_),
    .A1(net773));
 sg13g2_nor2_1 _2984_ (.A(net987),
    .B(_0754_),
    .Y(_0182_));
 sg13g2_o21ai_1 _2985_ (.B1(net927),
    .Y(_0755_),
    .A1(_0525_),
    .A2(net780));
 sg13g2_nand2_1 _2986_ (.Y(_0756_),
    .A(net820),
    .B(_0755_));
 sg13g2_a22oi_1 _2987_ (.Y(_0757_),
    .B1(_0756_),
    .B2(net309),
    .A2(net790),
    .A1(_0528_));
 sg13g2_nor2_1 _2988_ (.A(net987),
    .B(_0757_),
    .Y(_0183_));
 sg13g2_o21ai_1 _2989_ (.B1(net928),
    .Y(_0758_),
    .A1(_0530_),
    .A2(net784));
 sg13g2_nand2_1 _2990_ (.Y(_0759_),
    .A(net821),
    .B(_0758_));
 sg13g2_a22oi_1 _2991_ (.Y(_0760_),
    .B1(_0759_),
    .B2(net374),
    .A2(net764),
    .A1(_0533_));
 sg13g2_nor2_1 _2992_ (.A(net988),
    .B(_0760_),
    .Y(_0184_));
 sg13g2_o21ai_1 _2993_ (.B1(net927),
    .Y(_0761_),
    .A1(_0535_),
    .A2(net780));
 sg13g2_nand2_1 _2994_ (.Y(_0762_),
    .A(net820),
    .B(_0761_));
 sg13g2_a22oi_1 _2995_ (.Y(_0763_),
    .B1(_0762_),
    .B2(net262),
    .A2(net790),
    .A1(_0538_));
 sg13g2_nor2_1 _2996_ (.A(net988),
    .B(_0763_),
    .Y(_0185_));
 sg13g2_nor2_1 _2997_ (.A(_0540_),
    .B(net781),
    .Y(_0764_));
 sg13g2_o21ai_1 _2998_ (.B1(net823),
    .Y(_0765_),
    .A1(net897),
    .A2(_0764_));
 sg13g2_a22oi_1 _2999_ (.Y(_0766_),
    .B1(_0765_),
    .B2(net313),
    .A2(_0764_),
    .A1(net774));
 sg13g2_nor2_1 _3000_ (.A(net993),
    .B(_0766_),
    .Y(_0186_));
 sg13g2_nor2_1 _3001_ (.A(_0544_),
    .B(net781),
    .Y(_0767_));
 sg13g2_o21ai_1 _3002_ (.B1(net823),
    .Y(_0768_),
    .A1(net897),
    .A2(_0767_));
 sg13g2_a22oi_1 _3003_ (.Y(_0769_),
    .B1(_0768_),
    .B2(net306),
    .A2(_0767_),
    .A1(net774));
 sg13g2_nor2_1 _3004_ (.A(net993),
    .B(_0769_),
    .Y(_0187_));
 sg13g2_o21ai_1 _3005_ (.B1(net931),
    .Y(_0770_),
    .A1(_0548_),
    .A2(net781));
 sg13g2_nand2_1 _3006_ (.Y(_0771_),
    .A(net823),
    .B(_0770_));
 sg13g2_a22oi_1 _3007_ (.Y(_0772_),
    .B1(_0771_),
    .B2(net307),
    .A2(net763),
    .A1(_0551_));
 sg13g2_nor2_1 _3008_ (.A(net993),
    .B(_0772_),
    .Y(_0188_));
 sg13g2_a21oi_1 _3009_ (.A1(_0553_),
    .A2(net791),
    .Y(_0773_),
    .B1(net896));
 sg13g2_o21ai_1 _3010_ (.B1(net409),
    .Y(_0774_),
    .A1(net803),
    .A2(_0773_));
 sg13g2_nand3_1 _3011_ (.B(_0553_),
    .C(net791),
    .A(net774),
    .Y(_0775_));
 sg13g2_a21oi_1 _3012_ (.A1(_0774_),
    .A2(_0775_),
    .Y(_0189_),
    .B1(net992));
 sg13g2_nor2_1 _3013_ (.A(_0557_),
    .B(net780),
    .Y(_0776_));
 sg13g2_o21ai_1 _3014_ (.B1(net816),
    .Y(_0777_),
    .A1(net893),
    .A2(_0776_));
 sg13g2_a22oi_1 _3015_ (.Y(_0778_),
    .B1(_0777_),
    .B2(net303),
    .A2(_0776_),
    .A1(net773));
 sg13g2_nor2_1 _3016_ (.A(net983),
    .B(_0778_),
    .Y(_0190_));
 sg13g2_o21ai_1 _3017_ (.B1(net925),
    .Y(_0779_),
    .A1(_0561_),
    .A2(net780));
 sg13g2_nand2_1 _3018_ (.Y(_0780_),
    .A(net816),
    .B(_0779_));
 sg13g2_a22oi_1 _3019_ (.Y(_0781_),
    .B1(_0780_),
    .B2(net277),
    .A2(net788),
    .A1(_0564_));
 sg13g2_nor2_1 _3020_ (.A(net983),
    .B(_0781_),
    .Y(_0191_));
 sg13g2_o21ai_1 _3021_ (.B1(net924),
    .Y(_0782_),
    .A1(_0566_),
    .A2(net779));
 sg13g2_nand2_1 _3022_ (.Y(_0783_),
    .A(net815),
    .B(_0782_));
 sg13g2_a22oi_1 _3023_ (.Y(_0784_),
    .B1(_0783_),
    .B2(net258),
    .A2(net762),
    .A1(_0569_));
 sg13g2_nor2_1 _3024_ (.A(net982),
    .B(_0784_),
    .Y(_0192_));
 sg13g2_o21ai_1 _3025_ (.B1(net925),
    .Y(_0785_),
    .A1(_0571_),
    .A2(net779));
 sg13g2_nand2_1 _3026_ (.Y(_0786_),
    .A(net817),
    .B(_0785_));
 sg13g2_a22oi_1 _3027_ (.Y(_0787_),
    .B1(_0786_),
    .B2(net295),
    .A2(net788),
    .A1(_0574_));
 sg13g2_nor2_1 _3028_ (.A(net984),
    .B(_0787_),
    .Y(_0193_));
 sg13g2_nor2_1 _3029_ (.A(_0576_),
    .B(net779),
    .Y(_0788_));
 sg13g2_o21ai_1 _3030_ (.B1(net813),
    .Y(_0789_),
    .A1(net891),
    .A2(_0788_));
 sg13g2_a22oi_1 _3031_ (.Y(_0790_),
    .B1(_0789_),
    .B2(net281),
    .A2(_0788_),
    .A1(net771));
 sg13g2_nor2_1 _3032_ (.A(net979),
    .B(_0790_),
    .Y(_0194_));
 sg13g2_nor2_1 _3033_ (.A(_0580_),
    .B(net779),
    .Y(_0791_));
 sg13g2_o21ai_1 _3034_ (.B1(net813),
    .Y(_0792_),
    .A1(net892),
    .A2(_0791_));
 sg13g2_a22oi_1 _3035_ (.Y(_0793_),
    .B1(_0792_),
    .B2(net316),
    .A2(_0791_),
    .A1(net771));
 sg13g2_nor2_1 _3036_ (.A(net981),
    .B(_0793_),
    .Y(_0195_));
 sg13g2_o21ai_1 _3037_ (.B1(net926),
    .Y(_0794_),
    .A1(_0584_),
    .A2(net779));
 sg13g2_nand2_1 _3038_ (.Y(_0795_),
    .A(net812),
    .B(_0794_));
 sg13g2_a22oi_1 _3039_ (.Y(_0796_),
    .B1(_0795_),
    .B2(net415),
    .A2(net762),
    .A1(_0587_));
 sg13g2_nor2_1 _3040_ (.A(net979),
    .B(_0796_),
    .Y(_0196_));
 sg13g2_nor2_1 _3041_ (.A(_0589_),
    .B(net779),
    .Y(_0797_));
 sg13g2_o21ai_1 _3042_ (.B1(net813),
    .Y(_0798_),
    .A1(net892),
    .A2(_0797_));
 sg13g2_a22oi_1 _3043_ (.Y(_0799_),
    .B1(_0798_),
    .B2(net304),
    .A2(_0797_),
    .A1(net771));
 sg13g2_nor2_1 _3044_ (.A(net981),
    .B(_0799_),
    .Y(_0197_));
 sg13g2_o21ai_1 _3045_ (.B1(net934),
    .Y(_0800_),
    .A1(_0593_),
    .A2(net782));
 sg13g2_nand2_1 _3046_ (.Y(_0801_),
    .A(net827),
    .B(_0800_));
 sg13g2_a22oi_1 _3047_ (.Y(_0802_),
    .B1(_0801_),
    .B2(net434),
    .A2(net792),
    .A1(_0596_));
 sg13g2_nor2_1 _3048_ (.A(net996),
    .B(_0802_),
    .Y(_0198_));
 sg13g2_o21ai_1 _3049_ (.B1(net933),
    .Y(_0803_),
    .A1(_0598_),
    .A2(net782));
 sg13g2_nand2_1 _3050_ (.Y(_0804_),
    .A(net827),
    .B(_0803_));
 sg13g2_a22oi_1 _3051_ (.Y(_0805_),
    .B1(_0804_),
    .B2(net372),
    .A2(net792),
    .A1(_0601_));
 sg13g2_nor2_1 _3052_ (.A(net996),
    .B(_0805_),
    .Y(_0199_));
 sg13g2_and3_1 _3053_ (.X(_0806_),
    .A(net902),
    .B(_0439_),
    .C(net792));
 sg13g2_o21ai_1 _3054_ (.B1(net826),
    .Y(_0807_),
    .A1(net897),
    .A2(_0806_));
 sg13g2_a22oi_1 _3055_ (.Y(_0808_),
    .B1(_0807_),
    .B2(net263),
    .A2(net763),
    .A1(_0605_));
 sg13g2_nor2_1 _3056_ (.A(net994),
    .B(_0808_),
    .Y(_0200_));
 sg13g2_and3_1 _3057_ (.X(_0809_),
    .A(net903),
    .B(_0447_),
    .C(net791));
 sg13g2_o21ai_1 _3058_ (.B1(net827),
    .Y(_0810_),
    .A1(net898),
    .A2(_0809_));
 sg13g2_a22oi_1 _3059_ (.Y(_0811_),
    .B1(_0810_),
    .B2(net283),
    .A2(net792),
    .A1(_0609_));
 sg13g2_nor2_1 _3060_ (.A(net994),
    .B(_0811_),
    .Y(_0201_));
 sg13g2_nand3_1 _3061_ (.B(_0454_),
    .C(net791),
    .A(net900),
    .Y(_0812_));
 sg13g2_a21oi_1 _3062_ (.A1(net931),
    .A2(_0812_),
    .Y(_0813_),
    .B1(net802));
 sg13g2_nand2b_1 _3063_ (.Y(_0814_),
    .B(net501),
    .A_N(_0813_));
 sg13g2_o21ai_1 _3064_ (.B1(_0814_),
    .Y(_0815_),
    .A1(_0263_),
    .A2(_0812_));
 sg13g2_and2_1 _3065_ (.A(net1006),
    .B(_0815_),
    .X(_0202_));
 sg13g2_o21ai_1 _3066_ (.B1(net931),
    .Y(_0816_),
    .A1(_0615_),
    .A2(net781));
 sg13g2_nand2_1 _3067_ (.Y(_0817_),
    .A(net824),
    .B(_0816_));
 sg13g2_a22oi_1 _3068_ (.Y(_0818_),
    .B1(_0817_),
    .B2(net296),
    .A2(net791),
    .A1(_0618_));
 sg13g2_nor2_1 _3069_ (.A(net992),
    .B(_0818_),
    .Y(_0203_));
 sg13g2_nand3_1 _3070_ (.B(_0466_),
    .C(net791),
    .A(net901),
    .Y(_0819_));
 sg13g2_a21o_1 _3071_ (.A2(_0819_),
    .A1(net931),
    .B1(net803),
    .X(_0820_));
 sg13g2_a22oi_1 _3072_ (.Y(_0821_),
    .B1(_0820_),
    .B2(net287),
    .A2(net763),
    .A1(_0622_));
 sg13g2_nor2_1 _3073_ (.A(net992),
    .B(_0821_),
    .Y(_0204_));
 sg13g2_o21ai_1 _3074_ (.B1(net931),
    .Y(_0822_),
    .A1(_0624_),
    .A2(net781));
 sg13g2_nand2_1 _3075_ (.Y(_0823_),
    .A(net824),
    .B(_0822_));
 sg13g2_a22oi_1 _3076_ (.Y(_0824_),
    .B1(_0823_),
    .B2(net331),
    .A2(net791),
    .A1(_0627_));
 sg13g2_nor2_1 _3077_ (.A(net992),
    .B(_0824_),
    .Y(_0205_));
 sg13g2_nor2_1 _3078_ (.A(_0629_),
    .B(net779),
    .Y(_0825_));
 sg13g2_o21ai_1 _3079_ (.B1(net812),
    .Y(_0826_),
    .A1(net891),
    .A2(_0825_));
 sg13g2_a22oi_1 _3080_ (.Y(_0827_),
    .B1(_0826_),
    .B2(net268),
    .A2(_0825_),
    .A1(net773));
 sg13g2_nor2_1 _3081_ (.A(net982),
    .B(_0827_),
    .Y(_0206_));
 sg13g2_o21ai_1 _3082_ (.B1(net924),
    .Y(_0828_),
    .A1(net853),
    .A2(_0267_));
 sg13g2_nand2_1 _3083_ (.Y(_0829_),
    .A(net815),
    .B(_0828_));
 sg13g2_nor2_1 _3084_ (.A(net857),
    .B(net854),
    .Y(_0830_));
 sg13g2_nand2_2 _3085_ (.Y(_0831_),
    .A(net862),
    .B(net849));
 sg13g2_a22oi_1 _3086_ (.Y(_0832_),
    .B1(net778),
    .B2(_0274_),
    .A2(_0829_),
    .A1(net359));
 sg13g2_nor2_1 _3087_ (.A(net982),
    .B(_0832_),
    .Y(_0207_));
 sg13g2_o21ai_1 _3088_ (.B1(net922),
    .Y(_0833_),
    .A1(net852),
    .A2(_0278_));
 sg13g2_nand2_1 _3089_ (.Y(_0834_),
    .A(net810),
    .B(_0833_));
 sg13g2_nor2_2 _3090_ (.A(_1360_),
    .B(_0831_),
    .Y(_0835_));
 sg13g2_a22oi_1 _3091_ (.Y(_0836_),
    .B1(net758),
    .B2(_0284_),
    .A2(_0834_),
    .A1(net430));
 sg13g2_nor2_1 _3092_ (.A(net975),
    .B(net431),
    .Y(_0208_));
 sg13g2_o21ai_1 _3093_ (.B1(net924),
    .Y(_0837_),
    .A1(net853),
    .A2(_0289_));
 sg13g2_nand2_1 _3094_ (.Y(_0838_),
    .A(net815),
    .B(_0837_));
 sg13g2_a22oi_1 _3095_ (.Y(_0839_),
    .B1(_0838_),
    .B2(net317),
    .A2(net778),
    .A1(_0293_));
 sg13g2_nor2_1 _3096_ (.A(net982),
    .B(_0839_),
    .Y(_0209_));
 sg13g2_o21ai_1 _3097_ (.B1(net918),
    .Y(_0840_),
    .A1(net851),
    .A2(_0298_));
 sg13g2_nand2_1 _3098_ (.Y(_0841_),
    .A(net805),
    .B(_0840_));
 sg13g2_a22oi_1 _3099_ (.Y(_0842_),
    .B1(_0841_),
    .B2(net254),
    .A2(net757),
    .A1(_0301_));
 sg13g2_nor2_1 _3100_ (.A(net970),
    .B(_0842_),
    .Y(_0210_));
 sg13g2_o21ai_1 _3101_ (.B1(net918),
    .Y(_0843_),
    .A1(net851),
    .A2(_0305_));
 sg13g2_nand2_1 _3102_ (.Y(_0844_),
    .A(net806),
    .B(_0843_));
 sg13g2_a22oi_1 _3103_ (.Y(_0845_),
    .B1(_0844_),
    .B2(net315),
    .A2(net757),
    .A1(_0308_));
 sg13g2_nor2_1 _3104_ (.A(net970),
    .B(_0845_),
    .Y(_0211_));
 sg13g2_o21ai_1 _3105_ (.B1(net919),
    .Y(_0846_),
    .A1(net851),
    .A2(_0312_));
 sg13g2_nand2_1 _3106_ (.Y(_0847_),
    .A(net806),
    .B(_0846_));
 sg13g2_a22oi_1 _3107_ (.Y(_0848_),
    .B1(_0847_),
    .B2(net286),
    .A2(net757),
    .A1(_0318_));
 sg13g2_nor2_1 _3108_ (.A(net970),
    .B(_0848_),
    .Y(_0212_));
 sg13g2_o21ai_1 _3109_ (.B1(net918),
    .Y(_0849_),
    .A1(net851),
    .A2(_0323_));
 sg13g2_nand2_1 _3110_ (.Y(_0850_),
    .A(net806),
    .B(_0849_));
 sg13g2_a22oi_1 _3111_ (.Y(_0851_),
    .B1(_0850_),
    .B2(net305),
    .A2(net757),
    .A1(_0326_));
 sg13g2_nor2_1 _3112_ (.A(net970),
    .B(_0851_),
    .Y(_0213_));
 sg13g2_nor2_1 _3113_ (.A(_0328_),
    .B(_0831_),
    .Y(_0852_));
 sg13g2_nand2b_1 _3114_ (.Y(_0853_),
    .B(net776),
    .A_N(_0852_));
 sg13g2_a21oi_1 _3115_ (.A1(net477),
    .A2(net802),
    .Y(_0854_),
    .B1(net775));
 sg13g2_o21ai_1 _3116_ (.B1(net1004),
    .Y(_0855_),
    .A1(net477),
    .A2(_0852_));
 sg13g2_a21oi_1 _3117_ (.A1(_0853_),
    .A2(_0854_),
    .Y(_0214_),
    .B1(_0855_));
 sg13g2_o21ai_1 _3118_ (.B1(net927),
    .Y(_0856_),
    .A1(net854),
    .A2(_0334_));
 sg13g2_nand2_1 _3119_ (.Y(_0857_),
    .A(net820),
    .B(_0856_));
 sg13g2_a22oi_1 _3120_ (.Y(_0858_),
    .B1(_0857_),
    .B2(net253),
    .A2(_0830_),
    .A1(_0337_));
 sg13g2_nor2_1 _3121_ (.A(net987),
    .B(_0858_),
    .Y(_0215_));
 sg13g2_o21ai_1 _3122_ (.B1(net928),
    .Y(_0859_),
    .A1(net854),
    .A2(_0340_));
 sg13g2_nand2_1 _3123_ (.Y(_0860_),
    .A(net819),
    .B(_0859_));
 sg13g2_a22oi_1 _3124_ (.Y(_0861_),
    .B1(_0860_),
    .B2(net349),
    .A2(_0835_),
    .A1(_0344_));
 sg13g2_nor2_1 _3125_ (.A(net987),
    .B(_0861_),
    .Y(_0216_));
 sg13g2_o21ai_1 _3126_ (.B1(net927),
    .Y(_0862_),
    .A1(net854),
    .A2(_0348_));
 sg13g2_nand2_1 _3127_ (.Y(_0863_),
    .A(net820),
    .B(_0862_));
 sg13g2_a22oi_1 _3128_ (.Y(_0864_),
    .B1(_0863_),
    .B2(net308),
    .A2(_0830_),
    .A1(_0351_));
 sg13g2_nor2_1 _3129_ (.A(net987),
    .B(_0864_),
    .Y(_0217_));
 sg13g2_o21ai_1 _3130_ (.B1(net933),
    .Y(_0865_),
    .A1(net855),
    .A2(_0355_));
 sg13g2_nand2_1 _3131_ (.Y(_0866_),
    .A(net827),
    .B(_0865_));
 sg13g2_a22oi_1 _3132_ (.Y(_0867_),
    .B1(_0866_),
    .B2(net294),
    .A2(_0835_),
    .A1(_0358_));
 sg13g2_nor2_1 _3133_ (.A(net995),
    .B(_0867_),
    .Y(_0218_));
 sg13g2_o21ai_1 _3134_ (.B1(net933),
    .Y(_0868_),
    .A1(net855),
    .A2(_0361_));
 sg13g2_nand2_1 _3135_ (.Y(_0869_),
    .A(net826),
    .B(_0868_));
 sg13g2_a22oi_1 _3136_ (.Y(_0870_),
    .B1(_0869_),
    .B2(net371),
    .A2(_0835_),
    .A1(_0364_));
 sg13g2_nor2_1 _3137_ (.A(net995),
    .B(_0870_),
    .Y(_0219_));
 sg13g2_o21ai_1 _3138_ (.B1(net932),
    .Y(_0871_),
    .A1(net855),
    .A2(_0367_));
 sg13g2_nand2_1 _3139_ (.Y(_0872_),
    .A(net824),
    .B(_0871_));
 sg13g2_a22oi_1 _3140_ (.Y(_0873_),
    .B1(_0872_),
    .B2(net426),
    .A2(net759),
    .A1(_0372_));
 sg13g2_nor2_1 _3141_ (.A(net995),
    .B(_0873_),
    .Y(_0220_));
 sg13g2_o21ai_1 _3142_ (.B1(net930),
    .Y(_0874_),
    .A1(net854),
    .A2(_0376_));
 sg13g2_nand2_1 _3143_ (.Y(_0875_),
    .A(net826),
    .B(_0874_));
 sg13g2_a22oi_1 _3144_ (.Y(_0876_),
    .B1(_0875_),
    .B2(net297),
    .A2(net759),
    .A1(_0379_));
 sg13g2_nor2_1 _3145_ (.A(net995),
    .B(_0876_),
    .Y(_0221_));
 sg13g2_nor2_1 _3146_ (.A(_0382_),
    .B(_0831_),
    .Y(_0877_));
 sg13g2_o21ai_1 _3147_ (.B1(net815),
    .Y(_0878_),
    .A1(net893),
    .A2(_0877_));
 sg13g2_a22oi_1 _3148_ (.Y(_0879_),
    .B1(_0878_),
    .B2(net261),
    .A2(_0877_),
    .A1(net773));
 sg13g2_nor2_1 _3149_ (.A(net982),
    .B(_0879_),
    .Y(_0222_));
 sg13g2_o21ai_1 _3150_ (.B1(net924),
    .Y(_0880_),
    .A1(net853),
    .A2(_0386_));
 sg13g2_nand2_1 _3151_ (.Y(_0881_),
    .A(net815),
    .B(_0880_));
 sg13g2_a22oi_1 _3152_ (.Y(_0882_),
    .B1(_0881_),
    .B2(net280),
    .A2(net778),
    .A1(_0390_));
 sg13g2_nor2_1 _3153_ (.A(net983),
    .B(_0882_),
    .Y(_0223_));
 sg13g2_o21ai_1 _3154_ (.B1(net921),
    .Y(_0883_),
    .A1(net852),
    .A2(_0392_));
 sg13g2_nand2_1 _3155_ (.Y(_0884_),
    .A(net811),
    .B(_0883_));
 sg13g2_a22oi_1 _3156_ (.Y(_0885_),
    .B1(_0884_),
    .B2(net340),
    .A2(net758),
    .A1(_0396_));
 sg13g2_nor2_1 _3157_ (.A(net975),
    .B(_0885_),
    .Y(_0224_));
 sg13g2_o21ai_1 _3158_ (.B1(net922),
    .Y(_0886_),
    .A1(net852),
    .A2(_0398_));
 sg13g2_nand2_1 _3159_ (.Y(_0887_),
    .A(net810),
    .B(_0886_));
 sg13g2_a22oi_1 _3160_ (.Y(_0888_),
    .B1(_0887_),
    .B2(net298),
    .A2(net778),
    .A1(_0401_));
 sg13g2_nor2_1 _3161_ (.A(net975),
    .B(_0888_),
    .Y(_0225_));
 sg13g2_o21ai_1 _3162_ (.B1(net921),
    .Y(_0889_),
    .A1(net852),
    .A2(_0404_));
 sg13g2_nand2_1 _3163_ (.Y(_0890_),
    .A(net809),
    .B(_0889_));
 sg13g2_a22oi_1 _3164_ (.Y(_0891_),
    .B1(_0890_),
    .B2(net266),
    .A2(net758),
    .A1(_0407_));
 sg13g2_nor2_1 _3165_ (.A(net974),
    .B(_0891_),
    .Y(_0226_));
 sg13g2_o21ai_1 _3166_ (.B1(net921),
    .Y(_0892_),
    .A1(net852),
    .A2(_0409_));
 sg13g2_nand2_1 _3167_ (.Y(_0893_),
    .A(net809),
    .B(_0892_));
 sg13g2_a22oi_1 _3168_ (.Y(_0894_),
    .B1(_0893_),
    .B2(net327),
    .A2(net758),
    .A1(_0412_));
 sg13g2_nor2_1 _3169_ (.A(net973),
    .B(_0894_),
    .Y(_0227_));
 sg13g2_o21ai_1 _3170_ (.B1(net920),
    .Y(_0895_),
    .A1(net852),
    .A2(_0414_));
 sg13g2_nand2_1 _3171_ (.Y(_0896_),
    .A(net809),
    .B(_0895_));
 sg13g2_a22oi_1 _3172_ (.Y(_0897_),
    .B1(_0896_),
    .B2(net345),
    .A2(net758),
    .A1(_0418_));
 sg13g2_nor2_1 _3173_ (.A(net973),
    .B(_0897_),
    .Y(_0228_));
 sg13g2_o21ai_1 _3174_ (.B1(net921),
    .Y(_0898_),
    .A1(net852),
    .A2(_0421_));
 sg13g2_nand2_1 _3175_ (.Y(_0899_),
    .A(net809),
    .B(_0898_));
 sg13g2_a22oi_1 _3176_ (.Y(_0900_),
    .B1(_0899_),
    .B2(net269),
    .A2(net758),
    .A1(_0424_));
 sg13g2_nor2_1 _3177_ (.A(net973),
    .B(_0900_),
    .Y(_0229_));
 sg13g2_a21oi_1 _3178_ (.A1(net850),
    .A2(_0427_),
    .Y(_0901_),
    .B1(net894));
 sg13g2_o21ai_1 _3179_ (.B1(net493),
    .Y(_0902_),
    .A1(net802),
    .A2(_0901_));
 sg13g2_o21ai_1 _3180_ (.B1(_0902_),
    .Y(_0903_),
    .A1(_0430_),
    .A2(_0831_));
 sg13g2_and2_1 _3181_ (.A(net1003),
    .B(_0903_),
    .X(_0230_));
 sg13g2_o21ai_1 _3182_ (.B1(net929),
    .Y(_0904_),
    .A1(net854),
    .A2(_0434_));
 sg13g2_nand2_1 _3183_ (.Y(_0905_),
    .A(net818),
    .B(_0904_));
 sg13g2_a22oi_1 _3184_ (.Y(_0906_),
    .B1(_0905_),
    .B2(net260),
    .A2(net778),
    .A1(_0437_));
 sg13g2_nor2_1 _3185_ (.A(net985),
    .B(_0906_),
    .Y(_0231_));
 sg13g2_o21ai_1 _3186_ (.B1(net929),
    .Y(_0907_),
    .A1(net855),
    .A2(_0441_));
 sg13g2_nand2_1 _3187_ (.Y(_0908_),
    .A(net818),
    .B(_0907_));
 sg13g2_a22oi_1 _3188_ (.Y(_0909_),
    .B1(_0908_),
    .B2(net311),
    .A2(net759),
    .A1(_0445_));
 sg13g2_nor2_1 _3189_ (.A(net986),
    .B(_0909_),
    .Y(_0232_));
 sg13g2_o21ai_1 _3190_ (.B1(net929),
    .Y(_0910_),
    .A1(net854),
    .A2(_0449_));
 sg13g2_nand2_1 _3191_ (.Y(_0911_),
    .A(net818),
    .B(_0910_));
 sg13g2_a22oi_1 _3192_ (.Y(_0912_),
    .B1(_0911_),
    .B2(net357),
    .A2(net778),
    .A1(_0452_));
 sg13g2_nor2_1 _3193_ (.A(net985),
    .B(_0912_),
    .Y(_0233_));
 sg13g2_o21ai_1 _3194_ (.B1(net930),
    .Y(_0913_),
    .A1(net855),
    .A2(_0456_));
 sg13g2_nand2_1 _3195_ (.Y(_0914_),
    .A(net823),
    .B(_0913_));
 sg13g2_a22oi_1 _3196_ (.Y(_0915_),
    .B1(_0914_),
    .B2(net351),
    .A2(net759),
    .A1(_0459_));
 sg13g2_nor2_1 _3197_ (.A(net991),
    .B(_0915_),
    .Y(_0234_));
 sg13g2_nor2_1 _3198_ (.A(_0462_),
    .B(_0831_),
    .Y(_0916_));
 sg13g2_o21ai_1 _3199_ (.B1(net822),
    .Y(_0917_),
    .A1(net896),
    .A2(_0916_));
 sg13g2_a22oi_1 _3200_ (.Y(_0918_),
    .B1(_0917_),
    .B2(net332),
    .A2(_0916_),
    .A1(net774));
 sg13g2_nor2_1 _3201_ (.A(net991),
    .B(_0918_),
    .Y(_0235_));
 sg13g2_o21ai_1 _3202_ (.B1(net930),
    .Y(_0919_),
    .A1(net855),
    .A2(_0468_));
 sg13g2_nand2_1 _3203_ (.Y(_0920_),
    .A(net822),
    .B(_0919_));
 sg13g2_a22oi_1 _3204_ (.Y(_0921_),
    .B1(_0920_),
    .B2(net341),
    .A2(net759),
    .A1(_0472_));
 sg13g2_nor2_1 _3205_ (.A(net986),
    .B(_0921_),
    .Y(_0236_));
 sg13g2_nor2_1 _3206_ (.A(_0475_),
    .B(_0831_),
    .Y(_0922_));
 sg13g2_o21ai_1 _3207_ (.B1(net818),
    .Y(_0923_),
    .A1(net894),
    .A2(_0922_));
 sg13g2_a22oi_1 _3208_ (.Y(_0924_),
    .B1(_0923_),
    .B2(net320),
    .A2(_0922_),
    .A1(net772));
 sg13g2_nor2_1 _3209_ (.A(net985),
    .B(_0924_),
    .Y(_0237_));
 sg13g2_nor2_1 _3210_ (.A(_0480_),
    .B(_0831_),
    .Y(_0925_));
 sg13g2_o21ai_1 _3211_ (.B1(net812),
    .Y(_0926_),
    .A1(net891),
    .A2(_0925_));
 sg13g2_a22oi_1 _3212_ (.Y(_0927_),
    .B1(_0926_),
    .B2(net333),
    .A2(_0925_),
    .A1(net771));
 sg13g2_nor2_1 _3213_ (.A(net979),
    .B(_0927_),
    .Y(_0238_));
 sg13g2_o21ai_1 _3214_ (.B1(net926),
    .Y(_0928_),
    .A1(net853),
    .A2(_0484_));
 sg13g2_nand2_1 _3215_ (.Y(_0929_),
    .A(net813),
    .B(_0928_));
 sg13g2_a22oi_1 _3216_ (.Y(_0930_),
    .B1(_0929_),
    .B2(net350),
    .A2(net778),
    .A1(_0488_));
 sg13g2_nor2_1 _3217_ (.A(net979),
    .B(_0930_),
    .Y(_0239_));
 sg13g2_o21ai_1 _3218_ (.B1(net926),
    .Y(_0931_),
    .A1(net856),
    .A2(_0490_));
 sg13g2_nand2_1 _3219_ (.Y(_0932_),
    .A(net812),
    .B(_0931_));
 sg13g2_a22oi_1 _3220_ (.Y(_0933_),
    .B1(_0932_),
    .B2(net321),
    .A2(net759),
    .A1(_0493_));
 sg13g2_nor2_1 _3221_ (.A(net980),
    .B(_0933_),
    .Y(_0240_));
 sg13g2_o21ai_1 _3222_ (.B1(net926),
    .Y(_0934_),
    .A1(net853),
    .A2(_0495_));
 sg13g2_nand2_1 _3223_ (.Y(_0935_),
    .A(net814),
    .B(_0934_));
 sg13g2_a22oi_1 _3224_ (.Y(_0936_),
    .B1(_0935_),
    .B2(net282),
    .A2(net778),
    .A1(_0498_));
 sg13g2_nor2_1 _3225_ (.A(net980),
    .B(_0936_),
    .Y(_0241_));
 sg13g2_o21ai_1 _3226_ (.B1(net919),
    .Y(_0937_),
    .A1(net851),
    .A2(_0501_));
 sg13g2_nand2_1 _3227_ (.Y(_0938_),
    .A(net805),
    .B(_0937_));
 sg13g2_a22oi_1 _3228_ (.Y(_0939_),
    .B1(_0938_),
    .B2(net365),
    .A2(net757),
    .A1(_0504_));
 sg13g2_nor2_1 _3229_ (.A(net978),
    .B(_0939_),
    .Y(_0242_));
 sg13g2_o21ai_1 _3230_ (.B1(net919),
    .Y(_0940_),
    .A1(net851),
    .A2(_0506_));
 sg13g2_nand2_1 _3231_ (.Y(_0941_),
    .A(net808),
    .B(_0940_));
 sg13g2_a22oi_1 _3232_ (.Y(_0942_),
    .B1(_0941_),
    .B2(net278),
    .A2(net757),
    .A1(_0509_));
 sg13g2_nor2_1 _3233_ (.A(net972),
    .B(_0942_),
    .Y(_0243_));
 sg13g2_o21ai_1 _3234_ (.B1(net923),
    .Y(_0943_),
    .A1(net851),
    .A2(_0511_));
 sg13g2_nand2_1 _3235_ (.Y(_0944_),
    .A(net808),
    .B(_0943_));
 sg13g2_a22oi_1 _3236_ (.Y(_0945_),
    .B1(_0944_),
    .B2(net292),
    .A2(net757),
    .A1(_0514_));
 sg13g2_nor2_1 _3237_ (.A(net972),
    .B(_0945_),
    .Y(_0244_));
 sg13g2_o21ai_1 _3238_ (.B1(net918),
    .Y(_0946_),
    .A1(net851),
    .A2(_0516_));
 sg13g2_nand2_1 _3239_ (.Y(_0947_),
    .A(net805),
    .B(_0946_));
 sg13g2_a22oi_1 _3240_ (.Y(_0948_),
    .B1(_0947_),
    .B2(net429),
    .A2(net757),
    .A1(_0519_));
 sg13g2_nor2_1 _3241_ (.A(net971),
    .B(_0948_),
    .Y(_0245_));
 sg13g2_nor2_1 _3242_ (.A(_1212_),
    .B(_1256_),
    .Y(_0246_));
 sg13g2_dfrbp_1 _3243_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net61),
    .D(_0024_),
    .Q_N(_1618_),
    .Q(\ws2812_out.counter[0] ));
 sg13g2_dfrbp_1 _3244_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net238),
    .D(_0025_),
    .Q_N(_1617_),
    .Q(\ws2812_out.counter[1] ));
 sg13g2_dfrbp_1 _3245_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net237),
    .D(_0026_),
    .Q_N(_0012_),
    .Q(\ws2812_out.counter[2] ));
 sg13g2_dfrbp_1 _3246_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net236),
    .D(_0027_),
    .Q_N(_0013_),
    .Q(\ws2812_out.counter[3] ));
 sg13g2_dfrbp_1 _3247_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net235),
    .D(_0028_),
    .Q_N(_0014_),
    .Q(\ws2812_out.counter[4] ));
 sg13g2_dfrbp_1 _3248_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net234),
    .D(net470),
    .Q_N(_1616_),
    .Q(\ws2812_out.counter[5] ));
 sg13g2_dfrbp_1 _3249_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net233),
    .D(net472),
    .Q_N(_1615_),
    .Q(\ws2812_out.counter[6] ));
 sg13g2_dfrbp_1 _3250_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net232),
    .D(_0031_),
    .Q_N(_1614_),
    .Q(\ws2812_out.counter[7] ));
 sg13g2_dfrbp_1 _3251_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net231),
    .D(_0032_),
    .Q_N(_0019_),
    .Q(\ws2812_out.counter[8] ));
 sg13g2_dfrbp_1 _3252_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net230),
    .D(net511),
    .Q_N(_1613_),
    .Q(\ws2812_out.counter[9] ));
 sg13g2_dfrbp_1 _3253_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net229),
    .D(net302),
    .Q_N(_0018_),
    .Q(\ws2812_out.counter[10] ));
 sg13g2_dfrbp_1 _3254_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net228),
    .D(_0035_),
    .Q_N(_0023_),
    .Q(\uart_output.count[0] ));
 sg13g2_dfrbp_1 _3255_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net227),
    .D(_0036_),
    .Q_N(_1612_),
    .Q(\uart_output.count[1] ));
 sg13g2_dfrbp_1 _3256_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net226),
    .D(net386),
    .Q_N(_1611_),
    .Q(\uart_output.count[2] ));
 sg13g2_dfrbp_1 _3257_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net225),
    .D(_0038_),
    .Q_N(_1610_),
    .Q(\uart_output.count[3] ));
 sg13g2_dfrbp_1 _3258_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net224),
    .D(_0039_),
    .Q_N(_1609_),
    .Q(\uart_output.count[4] ));
 sg13g2_dfrbp_1 _3259_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net223),
    .D(_0040_),
    .Q_N(_1608_),
    .Q(\uart_output.count[5] ));
 sg13g2_dfrbp_1 _3260_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net222),
    .D(_0041_),
    .Q_N(_1607_),
    .Q(\uart_output.count[6] ));
 sg13g2_dfrbp_1 _3261_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net221),
    .D(_0042_),
    .Q_N(_1606_),
    .Q(\uart_output.count[7] ));
 sg13g2_dfrbp_1 _3262_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net220),
    .D(_0043_),
    .Q_N(_1605_),
    .Q(\ws2812_out.datacounter[0] ));
 sg13g2_dfrbp_1 _3263_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net218),
    .D(_0044_),
    .Q_N(_1604_),
    .Q(\ws2812_out.datacounter[1] ));
 sg13g2_dfrbp_1 _3264_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net216),
    .D(_0045_),
    .Q_N(_1603_),
    .Q(\ws2812_out.datacounter[2] ));
 sg13g2_dfrbp_1 _3265_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net214),
    .D(_0046_),
    .Q_N(_0017_),
    .Q(\ws2812_out.datacounter[3] ));
 sg13g2_dfrbp_1 _3266_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net212),
    .D(net482),
    .Q_N(_0010_),
    .Q(\ws2812_out.datacounter[4] ));
 sg13g2_dfrbp_1 _3267_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net210),
    .D(net500),
    .Q_N(_1602_),
    .Q(\ws2812_out.datacounter[5] ));
 sg13g2_dfrbp_1 _3268_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net208),
    .D(net442),
    .Q_N(_0011_),
    .Q(\ws2812_out.datacounter[6] ));
 sg13g2_dfrbp_1 _3269_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net206),
    .D(_0050_),
    .Q_N(_1601_),
    .Q(\ws2812_out.datacounter[7] ));
 sg13g2_dfrbp_1 _3270_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net204),
    .D(_0051_),
    .Q_N(_0009_),
    .Q(\uart_output.index[0] ));
 sg13g2_dfrbp_1 _3271_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net202),
    .D(_0052_),
    .Q_N(_0008_),
    .Q(\uart_output.index[1] ));
 sg13g2_dfrbp_1 _3272_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net200),
    .D(net479),
    .Q_N(_0007_),
    .Q(\uart_output.index[2] ));
 sg13g2_dfrbp_1 _3273_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net198),
    .D(net399),
    .Q_N(_0006_),
    .Q(\uart_output.index[3] ));
 sg13g2_dfrbp_1 _3274_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net196),
    .D(net514),
    .Q_N(_1600_),
    .Q(\uart_output.index[4] ));
 sg13g2_dfrbp_1 _3275_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net194),
    .D(net395),
    .Q_N(_0005_),
    .Q(\uart_output.index[5] ));
 sg13g2_dfrbp_1 _3276_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net192),
    .D(net436),
    .Q_N(_0004_),
    .Q(\uart_output.index[6] ));
 sg13g2_dfrbp_1 _3277_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net190),
    .D(net439),
    .Q_N(_0003_),
    .Q(\uart_output.index[7] ));
 sg13g2_dfrbp_1 _3278_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net188),
    .D(_0059_),
    .Q_N(_1599_),
    .Q(\spi_in.last_sck ));
 sg13g2_dfrbp_1 _3279_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net62),
    .D(net356),
    .Q_N(_1619_),
    .Q(\uart_output.uart_out ));
 sg13g2_dfrbp_1 _3280_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net63),
    .D(net492),
    .Q_N(_1620_),
    .Q(\spi_in.state[0] ));
 sg13g2_dfrbp_1 _3281_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net68),
    .D(net476),
    .Q_N(_0015_),
    .Q(\spi_in.state[1] ));
 sg13g2_dfrbp_1 _3282_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net187),
    .D(net448),
    .Q_N(_0016_),
    .Q(\spi_in.state[2] ));
 sg13g2_dfrbp_1 _3283_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net185),
    .D(_0061_),
    .Q_N(_1598_),
    .Q(\spi_in.index[0] ));
 sg13g2_dfrbp_1 _3284_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net183),
    .D(net505),
    .Q_N(_1597_),
    .Q(\spi_in.index[1] ));
 sg13g2_dfrbp_1 _3285_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net181),
    .D(net485),
    .Q_N(_0021_),
    .Q(\spi_in.index[2] ));
 sg13g2_dfrbp_1 _3286_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net179),
    .D(_0064_),
    .Q_N(_1596_),
    .Q(\spi_in.index[3] ));
 sg13g2_dfrbp_1 _3287_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net177),
    .D(_0065_),
    .Q_N(_0022_),
    .Q(\spi_in.index[4] ));
 sg13g2_dfrbp_1 _3288_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net175),
    .D(_0066_),
    .Q_N(_1595_),
    .Q(\spi_in.index[5] ));
 sg13g2_dfrbp_1 _3289_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net173),
    .D(_0067_),
    .Q_N(_1594_),
    .Q(\spi_in.index[6] ));
 sg13g2_dfrbp_1 _3290_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net171),
    .D(net497),
    .Q_N(_1593_),
    .Q(\spi_in.index[7] ));
 sg13g2_dfrbp_1 _3291_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net169),
    .D(net458),
    .Q_N(_1592_),
    .Q(\spi_in.bit_count[0] ));
 sg13g2_dfrbp_1 _3292_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net167),
    .D(net454),
    .Q_N(_1591_),
    .Q(\spi_in.bit_count[1] ));
 sg13g2_dfrbp_1 _3293_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net165),
    .D(_0071_),
    .Q_N(_1590_),
    .Q(\spi_in.bit_count[2] ));
 sg13g2_dfrbp_1 _3294_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net163),
    .D(_0072_),
    .Q_N(_1589_),
    .Q(\spi_in.bit_count[3] ));
 sg13g2_dfrbp_1 _3295_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net161),
    .D(_0073_),
    .Q_N(_1588_),
    .Q(\spi_in.bit_count[4] ));
 sg13g2_dfrbp_1 _3296_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net159),
    .D(_0074_),
    .Q_N(_1587_),
    .Q(\spi_in.bit_count[5] ));
 sg13g2_dfrbp_1 _3297_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net157),
    .D(_0075_),
    .Q_N(_1586_),
    .Q(\spi_in.bit_count[6] ));
 sg13g2_dfrbp_1 _3298_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net155),
    .D(_0076_),
    .Q_N(_1585_),
    .Q(\spi_in.bit_count[7] ));
 sg13g2_dfrbp_1 _3299_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net153),
    .D(net285),
    .Q_N(_0020_),
    .Q(\spi_in.bit_count[8] ));
 sg13g2_dfrbp_1 _3300_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net151),
    .D(_0078_),
    .Q_N(_1584_),
    .Q(\pixel_6[0] ));
 sg13g2_dfrbp_1 _3301_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net149),
    .D(_0079_),
    .Q_N(_1583_),
    .Q(\pixel_6[1] ));
 sg13g2_dfrbp_1 _3302_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net147),
    .D(_0080_),
    .Q_N(_1582_),
    .Q(\pixel_6[2] ));
 sg13g2_dfrbp_1 _3303_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net145),
    .D(_0081_),
    .Q_N(_1581_),
    .Q(\pixel_6[3] ));
 sg13g2_dfrbp_1 _3304_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net143),
    .D(_0082_),
    .Q_N(_1580_),
    .Q(\pixel_6[4] ));
 sg13g2_dfrbp_1 _3305_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net141),
    .D(_0083_),
    .Q_N(_1579_),
    .Q(\pixel_6[5] ));
 sg13g2_dfrbp_1 _3306_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net139),
    .D(_0084_),
    .Q_N(_1578_),
    .Q(\pixel_6[6] ));
 sg13g2_dfrbp_1 _3307_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net137),
    .D(_0085_),
    .Q_N(_1577_),
    .Q(\pixel_6[7] ));
 sg13g2_dfrbp_1 _3308_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net135),
    .D(_0086_),
    .Q_N(_1576_),
    .Q(\pixel_6[8] ));
 sg13g2_dfrbp_1 _3309_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net133),
    .D(_0087_),
    .Q_N(_1575_),
    .Q(\pixel_6[9] ));
 sg13g2_dfrbp_1 _3310_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net131),
    .D(_0088_),
    .Q_N(_1574_),
    .Q(\pixel_6[10] ));
 sg13g2_dfrbp_1 _3311_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net129),
    .D(_0089_),
    .Q_N(_1573_),
    .Q(\pixel_6[11] ));
 sg13g2_dfrbp_1 _3312_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net127),
    .D(_0090_),
    .Q_N(_1572_),
    .Q(\pixel_6[12] ));
 sg13g2_dfrbp_1 _3313_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net125),
    .D(_0091_),
    .Q_N(_1571_),
    .Q(\pixel_6[13] ));
 sg13g2_dfrbp_1 _3314_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net123),
    .D(_0092_),
    .Q_N(_1570_),
    .Q(\pixel_6[14] ));
 sg13g2_dfrbp_1 _3315_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net121),
    .D(_0093_),
    .Q_N(_1569_),
    .Q(\pixel_6[15] ));
 sg13g2_dfrbp_1 _3316_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net119),
    .D(_0094_),
    .Q_N(_1568_),
    .Q(\pixel_6[16] ));
 sg13g2_dfrbp_1 _3317_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net117),
    .D(_0095_),
    .Q_N(_1567_),
    .Q(\pixel_6[17] ));
 sg13g2_dfrbp_1 _3318_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net115),
    .D(_0096_),
    .Q_N(_1566_),
    .Q(\pixel_6[18] ));
 sg13g2_dfrbp_1 _3319_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net113),
    .D(_0097_),
    .Q_N(_1565_),
    .Q(\pixel_6[19] ));
 sg13g2_dfrbp_1 _3320_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net111),
    .D(_0098_),
    .Q_N(_1564_),
    .Q(\pixel_6[20] ));
 sg13g2_dfrbp_1 _3321_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net109),
    .D(_0099_),
    .Q_N(_1563_),
    .Q(\pixel_6[21] ));
 sg13g2_dfrbp_1 _3322_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net107),
    .D(_0100_),
    .Q_N(_1562_),
    .Q(\pixel_6[22] ));
 sg13g2_dfrbp_1 _3323_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net105),
    .D(_0101_),
    .Q_N(_1561_),
    .Q(\pixel_6[23] ));
 sg13g2_dfrbp_1 _3324_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net103),
    .D(_0102_),
    .Q_N(_1560_),
    .Q(\pixel_5[0] ));
 sg13g2_dfrbp_1 _3325_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net101),
    .D(_0103_),
    .Q_N(_1559_),
    .Q(\pixel_5[1] ));
 sg13g2_dfrbp_1 _3326_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net99),
    .D(_0104_),
    .Q_N(_1558_),
    .Q(\pixel_5[2] ));
 sg13g2_dfrbp_1 _3327_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net97),
    .D(_0105_),
    .Q_N(_1557_),
    .Q(\pixel_5[3] ));
 sg13g2_dfrbp_1 _3328_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net95),
    .D(_0106_),
    .Q_N(_1556_),
    .Q(\pixel_5[4] ));
 sg13g2_dfrbp_1 _3329_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net93),
    .D(_0107_),
    .Q_N(_1555_),
    .Q(\pixel_5[5] ));
 sg13g2_dfrbp_1 _3330_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net91),
    .D(_0108_),
    .Q_N(_1554_),
    .Q(\pixel_5[6] ));
 sg13g2_dfrbp_1 _3331_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net89),
    .D(_0109_),
    .Q_N(_1553_),
    .Q(\pixel_5[7] ));
 sg13g2_dfrbp_1 _3332_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net87),
    .D(_0110_),
    .Q_N(_1552_),
    .Q(\pixel_5[8] ));
 sg13g2_dfrbp_1 _3333_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net85),
    .D(_0111_),
    .Q_N(_1551_),
    .Q(\pixel_5[9] ));
 sg13g2_dfrbp_1 _3334_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net83),
    .D(_0112_),
    .Q_N(_1550_),
    .Q(\pixel_5[10] ));
 sg13g2_dfrbp_1 _3335_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net81),
    .D(_0113_),
    .Q_N(_1549_),
    .Q(\pixel_5[11] ));
 sg13g2_dfrbp_1 _3336_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net79),
    .D(_0114_),
    .Q_N(_1548_),
    .Q(\pixel_5[12] ));
 sg13g2_dfrbp_1 _3337_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net77),
    .D(_0115_),
    .Q_N(_1547_),
    .Q(\pixel_5[13] ));
 sg13g2_dfrbp_1 _3338_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net75),
    .D(_0116_),
    .Q_N(_1546_),
    .Q(\pixel_5[14] ));
 sg13g2_dfrbp_1 _3339_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net73),
    .D(_0117_),
    .Q_N(_1545_),
    .Q(\pixel_5[15] ));
 sg13g2_dfrbp_1 _3340_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net71),
    .D(_0118_),
    .Q_N(_1544_),
    .Q(\pixel_5[16] ));
 sg13g2_dfrbp_1 _3341_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net69),
    .D(_0119_),
    .Q_N(_1543_),
    .Q(\pixel_5[17] ));
 sg13g2_dfrbp_1 _3342_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net67),
    .D(_0120_),
    .Q_N(_1542_),
    .Q(\pixel_5[18] ));
 sg13g2_dfrbp_1 _3343_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net65),
    .D(_0121_),
    .Q_N(_1541_),
    .Q(\pixel_5[19] ));
 sg13g2_dfrbp_1 _3344_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net60),
    .D(_0122_),
    .Q_N(_1540_),
    .Q(\pixel_5[20] ));
 sg13g2_dfrbp_1 _3345_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net58),
    .D(_0123_),
    .Q_N(_1539_),
    .Q(\pixel_5[21] ));
 sg13g2_dfrbp_1 _3346_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net56),
    .D(_0124_),
    .Q_N(_1538_),
    .Q(\pixel_5[22] ));
 sg13g2_dfrbp_1 _3347_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net54),
    .D(_0125_),
    .Q_N(_1537_),
    .Q(\pixel_5[23] ));
 sg13g2_dfrbp_1 _3348_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net52),
    .D(_0126_),
    .Q_N(_1536_),
    .Q(\pixel_4[0] ));
 sg13g2_dfrbp_1 _3349_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net50),
    .D(_0127_),
    .Q_N(_1535_),
    .Q(\pixel_4[1] ));
 sg13g2_dfrbp_1 _3350_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net48),
    .D(_0128_),
    .Q_N(_1534_),
    .Q(\pixel_4[2] ));
 sg13g2_dfrbp_1 _3351_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net46),
    .D(_0129_),
    .Q_N(_1533_),
    .Q(\pixel_4[3] ));
 sg13g2_dfrbp_1 _3352_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net44),
    .D(_0130_),
    .Q_N(_1532_),
    .Q(\pixel_4[4] ));
 sg13g2_dfrbp_1 _3353_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net42),
    .D(_0131_),
    .Q_N(_1531_),
    .Q(\pixel_4[5] ));
 sg13g2_dfrbp_1 _3354_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net40),
    .D(_0132_),
    .Q_N(_1530_),
    .Q(\pixel_4[6] ));
 sg13g2_dfrbp_1 _3355_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net38),
    .D(_0133_),
    .Q_N(_1529_),
    .Q(\pixel_4[7] ));
 sg13g2_dfrbp_1 _3356_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net36),
    .D(_0134_),
    .Q_N(_1528_),
    .Q(\pixel_4[8] ));
 sg13g2_dfrbp_1 _3357_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net34),
    .D(_0135_),
    .Q_N(_1527_),
    .Q(\pixel_4[9] ));
 sg13g2_dfrbp_1 _3358_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net32),
    .D(_0136_),
    .Q_N(_1526_),
    .Q(\pixel_4[10] ));
 sg13g2_dfrbp_1 _3359_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net30),
    .D(_0137_),
    .Q_N(_1525_),
    .Q(\pixel_4[11] ));
 sg13g2_dfrbp_1 _3360_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net28),
    .D(_0138_),
    .Q_N(_1524_),
    .Q(\pixel_4[12] ));
 sg13g2_dfrbp_1 _3361_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net26),
    .D(_0139_),
    .Q_N(_1523_),
    .Q(\pixel_4[13] ));
 sg13g2_dfrbp_1 _3362_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net24),
    .D(_0140_),
    .Q_N(_1522_),
    .Q(\pixel_4[14] ));
 sg13g2_dfrbp_1 _3363_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net248),
    .D(_0141_),
    .Q_N(_1521_),
    .Q(\pixel_4[15] ));
 sg13g2_dfrbp_1 _3364_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net246),
    .D(_0142_),
    .Q_N(_1520_),
    .Q(\pixel_4[16] ));
 sg13g2_dfrbp_1 _3365_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net244),
    .D(_0143_),
    .Q_N(_1519_),
    .Q(\pixel_4[17] ));
 sg13g2_dfrbp_1 _3366_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net242),
    .D(_0144_),
    .Q_N(_1518_),
    .Q(\pixel_4[18] ));
 sg13g2_dfrbp_1 _3367_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net240),
    .D(_0145_),
    .Q_N(_1517_),
    .Q(\pixel_4[19] ));
 sg13g2_dfrbp_1 _3368_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net219),
    .D(_0146_),
    .Q_N(_1516_),
    .Q(\pixel_4[20] ));
 sg13g2_dfrbp_1 _3369_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net215),
    .D(_0147_),
    .Q_N(_1515_),
    .Q(\pixel_4[21] ));
 sg13g2_dfrbp_1 _3370_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net211),
    .D(_0148_),
    .Q_N(_1514_),
    .Q(\pixel_4[22] ));
 sg13g2_dfrbp_1 _3371_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net207),
    .D(_0149_),
    .Q_N(_1513_),
    .Q(\pixel_4[23] ));
 sg13g2_dfrbp_1 _3372_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net203),
    .D(_0150_),
    .Q_N(_1512_),
    .Q(\pixel_3[0] ));
 sg13g2_dfrbp_1 _3373_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net199),
    .D(_0151_),
    .Q_N(_1511_),
    .Q(\pixel_3[1] ));
 sg13g2_dfrbp_1 _3374_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net195),
    .D(_0152_),
    .Q_N(_1510_),
    .Q(\pixel_3[2] ));
 sg13g2_dfrbp_1 _3375_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net191),
    .D(_0153_),
    .Q_N(_1509_),
    .Q(\pixel_3[3] ));
 sg13g2_dfrbp_1 _3376_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net186),
    .D(_0154_),
    .Q_N(_1508_),
    .Q(\pixel_3[4] ));
 sg13g2_dfrbp_1 _3377_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net182),
    .D(_0155_),
    .Q_N(_1507_),
    .Q(\pixel_3[5] ));
 sg13g2_dfrbp_1 _3378_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net178),
    .D(_0156_),
    .Q_N(_1506_),
    .Q(\pixel_3[6] ));
 sg13g2_dfrbp_1 _3379_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net174),
    .D(_0157_),
    .Q_N(_1505_),
    .Q(\pixel_3[7] ));
 sg13g2_dfrbp_1 _3380_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net170),
    .D(_0158_),
    .Q_N(_1504_),
    .Q(\pixel_3[8] ));
 sg13g2_dfrbp_1 _3381_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net166),
    .D(_0159_),
    .Q_N(_1503_),
    .Q(\pixel_3[9] ));
 sg13g2_dfrbp_1 _3382_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net162),
    .D(_0160_),
    .Q_N(_1502_),
    .Q(\pixel_3[10] ));
 sg13g2_dfrbp_1 _3383_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net158),
    .D(_0161_),
    .Q_N(_1501_),
    .Q(\pixel_3[11] ));
 sg13g2_dfrbp_1 _3384_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net154),
    .D(_0162_),
    .Q_N(_1500_),
    .Q(\pixel_3[12] ));
 sg13g2_dfrbp_1 _3385_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net150),
    .D(_0163_),
    .Q_N(_1499_),
    .Q(\pixel_3[13] ));
 sg13g2_dfrbp_1 _3386_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net146),
    .D(_0164_),
    .Q_N(_1498_),
    .Q(\pixel_3[14] ));
 sg13g2_dfrbp_1 _3387_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net142),
    .D(_0165_),
    .Q_N(_1497_),
    .Q(\pixel_3[15] ));
 sg13g2_dfrbp_1 _3388_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net138),
    .D(_0166_),
    .Q_N(_1496_),
    .Q(\pixel_3[16] ));
 sg13g2_dfrbp_1 _3389_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net134),
    .D(_0167_),
    .Q_N(_1495_),
    .Q(\pixel_3[17] ));
 sg13g2_dfrbp_1 _3390_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net130),
    .D(_0168_),
    .Q_N(_1494_),
    .Q(\pixel_3[18] ));
 sg13g2_dfrbp_1 _3391_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net126),
    .D(_0169_),
    .Q_N(_1493_),
    .Q(\pixel_3[19] ));
 sg13g2_dfrbp_1 _3392_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net122),
    .D(_0170_),
    .Q_N(_1492_),
    .Q(\pixel_3[20] ));
 sg13g2_dfrbp_1 _3393_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net118),
    .D(_0171_),
    .Q_N(_1491_),
    .Q(\pixel_3[21] ));
 sg13g2_dfrbp_1 _3394_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net114),
    .D(_0172_),
    .Q_N(_1490_),
    .Q(\pixel_3[22] ));
 sg13g2_dfrbp_1 _3395_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net110),
    .D(_0173_),
    .Q_N(_1489_),
    .Q(\pixel_3[23] ));
 sg13g2_dfrbp_1 _3396_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net106),
    .D(_0174_),
    .Q_N(_1488_),
    .Q(\pixel_2[0] ));
 sg13g2_dfrbp_1 _3397_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net102),
    .D(_0175_),
    .Q_N(_1487_),
    .Q(\pixel_2[1] ));
 sg13g2_dfrbp_1 _3398_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net98),
    .D(_0176_),
    .Q_N(_1486_),
    .Q(\pixel_2[2] ));
 sg13g2_dfrbp_1 _3399_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net94),
    .D(_0177_),
    .Q_N(_1485_),
    .Q(\pixel_2[3] ));
 sg13g2_dfrbp_1 _3400_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net90),
    .D(_0178_),
    .Q_N(_1484_),
    .Q(\pixel_2[4] ));
 sg13g2_dfrbp_1 _3401_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net86),
    .D(_0179_),
    .Q_N(_1483_),
    .Q(\pixel_2[5] ));
 sg13g2_dfrbp_1 _3402_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net82),
    .D(_0180_),
    .Q_N(_1482_),
    .Q(\pixel_2[6] ));
 sg13g2_dfrbp_1 _3403_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net78),
    .D(_0181_),
    .Q_N(_1481_),
    .Q(\pixel_2[7] ));
 sg13g2_dfrbp_1 _3404_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net74),
    .D(_0182_),
    .Q_N(_1480_),
    .Q(\pixel_2[8] ));
 sg13g2_dfrbp_1 _3405_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net70),
    .D(_0183_),
    .Q_N(_1479_),
    .Q(\pixel_2[9] ));
 sg13g2_dfrbp_1 _3406_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net66),
    .D(_0184_),
    .Q_N(_1478_),
    .Q(\pixel_2[10] ));
 sg13g2_dfrbp_1 _3407_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net59),
    .D(_0185_),
    .Q_N(_1477_),
    .Q(\pixel_2[11] ));
 sg13g2_dfrbp_1 _3408_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net55),
    .D(_0186_),
    .Q_N(_1476_),
    .Q(\pixel_2[12] ));
 sg13g2_dfrbp_1 _3409_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net51),
    .D(_0187_),
    .Q_N(_1475_),
    .Q(\pixel_2[13] ));
 sg13g2_dfrbp_1 _3410_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net47),
    .D(_0188_),
    .Q_N(_1474_),
    .Q(\pixel_2[14] ));
 sg13g2_dfrbp_1 _3411_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net43),
    .D(_0189_),
    .Q_N(_1473_),
    .Q(\pixel_2[15] ));
 sg13g2_dfrbp_1 _3412_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net39),
    .D(_0190_),
    .Q_N(_1472_),
    .Q(\pixel_2[16] ));
 sg13g2_dfrbp_1 _3413_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net35),
    .D(_0191_),
    .Q_N(_1471_),
    .Q(\pixel_2[17] ));
 sg13g2_dfrbp_1 _3414_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net31),
    .D(_0192_),
    .Q_N(_1470_),
    .Q(\pixel_2[18] ));
 sg13g2_dfrbp_1 _3415_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net27),
    .D(_0193_),
    .Q_N(_1469_),
    .Q(\pixel_2[19] ));
 sg13g2_dfrbp_1 _3416_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net249),
    .D(_0194_),
    .Q_N(_1468_),
    .Q(\pixel_2[20] ));
 sg13g2_dfrbp_1 _3417_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net245),
    .D(_0195_),
    .Q_N(_1467_),
    .Q(\pixel_2[21] ));
 sg13g2_dfrbp_1 _3418_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net241),
    .D(_0196_),
    .Q_N(_1466_),
    .Q(\pixel_2[22] ));
 sg13g2_dfrbp_1 _3419_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net217),
    .D(_0197_),
    .Q_N(_1465_),
    .Q(\pixel_2[23] ));
 sg13g2_dfrbp_1 _3420_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net209),
    .D(_0198_),
    .Q_N(_1464_),
    .Q(\pixel_1[0] ));
 sg13g2_dfrbp_1 _3421_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net201),
    .D(_0199_),
    .Q_N(_1463_),
    .Q(\pixel_1[1] ));
 sg13g2_dfrbp_1 _3422_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net193),
    .D(_0200_),
    .Q_N(_1462_),
    .Q(\pixel_1[2] ));
 sg13g2_dfrbp_1 _3423_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net184),
    .D(_0201_),
    .Q_N(_1461_),
    .Q(\pixel_1[3] ));
 sg13g2_dfrbp_1 _3424_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net176),
    .D(_0202_),
    .Q_N(_1460_),
    .Q(\pixel_1[4] ));
 sg13g2_dfrbp_1 _3425_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net168),
    .D(_0203_),
    .Q_N(_1459_),
    .Q(\pixel_1[5] ));
 sg13g2_dfrbp_1 _3426_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net160),
    .D(_0204_),
    .Q_N(_1458_),
    .Q(\pixel_1[6] ));
 sg13g2_dfrbp_1 _3427_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net152),
    .D(_0205_),
    .Q_N(_1457_),
    .Q(\pixel_1[7] ));
 sg13g2_dfrbp_1 _3428_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net144),
    .D(_0206_),
    .Q_N(_1456_),
    .Q(\pixel_1[8] ));
 sg13g2_dfrbp_1 _3429_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net136),
    .D(_0207_),
    .Q_N(_1455_),
    .Q(\pixel_1[9] ));
 sg13g2_dfrbp_1 _3430_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net128),
    .D(_0208_),
    .Q_N(_1454_),
    .Q(\pixel_1[10] ));
 sg13g2_dfrbp_1 _3431_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net120),
    .D(_0209_),
    .Q_N(_1453_),
    .Q(\pixel_1[11] ));
 sg13g2_dfrbp_1 _3432_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net112),
    .D(_0210_),
    .Q_N(_1452_),
    .Q(\pixel_1[12] ));
 sg13g2_dfrbp_1 _3433_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net104),
    .D(_0211_),
    .Q_N(_1451_),
    .Q(\pixel_1[13] ));
 sg13g2_dfrbp_1 _3434_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net96),
    .D(_0212_),
    .Q_N(_1450_),
    .Q(\pixel_1[14] ));
 sg13g2_dfrbp_1 _3435_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net88),
    .D(_0213_),
    .Q_N(_1449_),
    .Q(\pixel_1[15] ));
 sg13g2_dfrbp_1 _3436_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net80),
    .D(_0214_),
    .Q_N(_1448_),
    .Q(\pixel_1[16] ));
 sg13g2_dfrbp_1 _3437_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net72),
    .D(_0215_),
    .Q_N(_1447_),
    .Q(\pixel_1[17] ));
 sg13g2_dfrbp_1 _3438_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net64),
    .D(_0216_),
    .Q_N(_1446_),
    .Q(\pixel_1[18] ));
 sg13g2_dfrbp_1 _3439_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net53),
    .D(_0217_),
    .Q_N(_1445_),
    .Q(\pixel_1[19] ));
 sg13g2_dfrbp_1 _3440_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net45),
    .D(_0218_),
    .Q_N(_1444_),
    .Q(\pixel_1[20] ));
 sg13g2_dfrbp_1 _3441_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net37),
    .D(_0219_),
    .Q_N(_1443_),
    .Q(\pixel_1[21] ));
 sg13g2_dfrbp_1 _3442_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net29),
    .D(_0220_),
    .Q_N(_1442_),
    .Q(\pixel_1[22] ));
 sg13g2_dfrbp_1 _3443_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net247),
    .D(_0221_),
    .Q_N(_1441_),
    .Q(\pixel_1[23] ));
 sg13g2_dfrbp_1 _3444_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net239),
    .D(_0222_),
    .Q_N(_1440_),
    .Q(\pixel_0[0] ));
 sg13g2_dfrbp_1 _3445_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net205),
    .D(_0223_),
    .Q_N(_1439_),
    .Q(\pixel_0[1] ));
 sg13g2_dfrbp_1 _3446_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net189),
    .D(_0224_),
    .Q_N(_1438_),
    .Q(\pixel_0[2] ));
 sg13g2_dfrbp_1 _3447_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net172),
    .D(_0225_),
    .Q_N(_1437_),
    .Q(\pixel_0[3] ));
 sg13g2_dfrbp_1 _3448_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net156),
    .D(_0226_),
    .Q_N(_1436_),
    .Q(\pixel_0[4] ));
 sg13g2_dfrbp_1 _3449_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net140),
    .D(_0227_),
    .Q_N(_1435_),
    .Q(\pixel_0[5] ));
 sg13g2_dfrbp_1 _3450_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net124),
    .D(_0228_),
    .Q_N(_1434_),
    .Q(\pixel_0[6] ));
 sg13g2_dfrbp_1 _3451_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net108),
    .D(_0229_),
    .Q_N(_1433_),
    .Q(\pixel_0[7] ));
 sg13g2_dfrbp_1 _3452_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net92),
    .D(_0230_),
    .Q_N(_1432_),
    .Q(\pixel_0[8] ));
 sg13g2_dfrbp_1 _3453_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net76),
    .D(_0231_),
    .Q_N(_1431_),
    .Q(\pixel_0[9] ));
 sg13g2_dfrbp_1 _3454_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net57),
    .D(_0232_),
    .Q_N(_1430_),
    .Q(\pixel_0[10] ));
 sg13g2_dfrbp_1 _3455_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net41),
    .D(_0233_),
    .Q_N(_1429_),
    .Q(\pixel_0[11] ));
 sg13g2_dfrbp_1 _3456_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net25),
    .D(_0234_),
    .Q_N(_1428_),
    .Q(\pixel_0[12] ));
 sg13g2_dfrbp_1 _3457_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net213),
    .D(_0235_),
    .Q_N(_1427_),
    .Q(\pixel_0[13] ));
 sg13g2_dfrbp_1 _3458_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net180),
    .D(_0236_),
    .Q_N(_1426_),
    .Q(\pixel_0[14] ));
 sg13g2_dfrbp_1 _3459_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net148),
    .D(_0237_),
    .Q_N(_1425_),
    .Q(\pixel_0[15] ));
 sg13g2_dfrbp_1 _3460_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net116),
    .D(_0238_),
    .Q_N(_1424_),
    .Q(\pixel_0[16] ));
 sg13g2_dfrbp_1 _3461_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net84),
    .D(_0239_),
    .Q_N(_1423_),
    .Q(\pixel_0[17] ));
 sg13g2_dfrbp_1 _3462_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net49),
    .D(_0240_),
    .Q_N(_1422_),
    .Q(\pixel_0[18] ));
 sg13g2_dfrbp_1 _3463_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net243),
    .D(_0241_),
    .Q_N(_1421_),
    .Q(\pixel_0[19] ));
 sg13g2_dfrbp_1 _3464_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net164),
    .D(_0242_),
    .Q_N(_1420_),
    .Q(\pixel_0[20] ));
 sg13g2_dfrbp_1 _3465_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net100),
    .D(_0243_),
    .Q_N(_1419_),
    .Q(\pixel_0[21] ));
 sg13g2_dfrbp_1 _3466_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net33),
    .D(_0244_),
    .Q_N(_1418_),
    .Q(\pixel_0[22] ));
 sg13g2_dfrbp_1 _3467_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net132),
    .D(_0245_),
    .Q_N(_1417_),
    .Q(\pixel_0[23] ));
 sg13g2_dfrbp_1 _3468_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net197),
    .D(_0246_),
    .Q_N(_1416_),
    .Q(\ws2812_out.state ));
 sg13g2_tiehi _3456__25 (.L_HI(net25));
 sg13g2_tiehi _3361__26 (.L_HI(net26));
 sg13g2_tiehi _3415__27 (.L_HI(net27));
 sg13g2_tiehi _3360__28 (.L_HI(net28));
 sg13g2_tiehi _3442__29 (.L_HI(net29));
 sg13g2_tiehi _3359__30 (.L_HI(net30));
 sg13g2_tiehi _3414__31 (.L_HI(net31));
 sg13g2_tiehi _3358__32 (.L_HI(net32));
 sg13g2_tiehi _3466__33 (.L_HI(net33));
 sg13g2_tiehi _3357__34 (.L_HI(net34));
 sg13g2_tiehi _3413__35 (.L_HI(net35));
 sg13g2_tiehi _3356__36 (.L_HI(net36));
 sg13g2_tiehi _3441__37 (.L_HI(net37));
 sg13g2_tiehi _3355__38 (.L_HI(net38));
 sg13g2_tiehi _3412__39 (.L_HI(net39));
 sg13g2_tiehi _3354__40 (.L_HI(net40));
 sg13g2_tiehi _3455__41 (.L_HI(net41));
 sg13g2_tiehi _3353__42 (.L_HI(net42));
 sg13g2_tiehi _3411__43 (.L_HI(net43));
 sg13g2_tiehi _3352__44 (.L_HI(net44));
 sg13g2_tiehi _3440__45 (.L_HI(net45));
 sg13g2_tiehi _3351__46 (.L_HI(net46));
 sg13g2_tiehi _3410__47 (.L_HI(net47));
 sg13g2_tiehi _3350__48 (.L_HI(net48));
 sg13g2_tiehi _3462__49 (.L_HI(net49));
 sg13g2_tiehi _3349__50 (.L_HI(net50));
 sg13g2_tiehi _3409__51 (.L_HI(net51));
 sg13g2_tiehi _3348__52 (.L_HI(net52));
 sg13g2_tiehi _3439__53 (.L_HI(net53));
 sg13g2_tiehi _3347__54 (.L_HI(net54));
 sg13g2_tiehi _3408__55 (.L_HI(net55));
 sg13g2_tiehi _3346__56 (.L_HI(net56));
 sg13g2_tiehi _3454__57 (.L_HI(net57));
 sg13g2_tiehi _3345__58 (.L_HI(net58));
 sg13g2_tiehi _3407__59 (.L_HI(net59));
 sg13g2_tiehi _3344__60 (.L_HI(net60));
 sg13g2_tiehi _3243__61 (.L_HI(net61));
 sg13g2_tiehi _3279__62 (.L_HI(net62));
 sg13g2_tiehi _3280__63 (.L_HI(net63));
 sg13g2_tiehi _3438__64 (.L_HI(net64));
 sg13g2_tiehi _3343__65 (.L_HI(net65));
 sg13g2_tiehi _3406__66 (.L_HI(net66));
 sg13g2_tiehi _3342__67 (.L_HI(net67));
 sg13g2_tiehi _3281__68 (.L_HI(net68));
 sg13g2_tiehi _3341__69 (.L_HI(net69));
 sg13g2_tiehi _3405__70 (.L_HI(net70));
 sg13g2_tiehi _3340__71 (.L_HI(net71));
 sg13g2_tiehi _3437__72 (.L_HI(net72));
 sg13g2_tiehi _3339__73 (.L_HI(net73));
 sg13g2_tiehi _3404__74 (.L_HI(net74));
 sg13g2_tiehi _3338__75 (.L_HI(net75));
 sg13g2_tiehi _3453__76 (.L_HI(net76));
 sg13g2_tiehi _3337__77 (.L_HI(net77));
 sg13g2_tiehi _3403__78 (.L_HI(net78));
 sg13g2_tiehi _3336__79 (.L_HI(net79));
 sg13g2_tiehi _3436__80 (.L_HI(net80));
 sg13g2_tiehi _3335__81 (.L_HI(net81));
 sg13g2_tiehi _3402__82 (.L_HI(net82));
 sg13g2_tiehi _3334__83 (.L_HI(net83));
 sg13g2_tiehi _3461__84 (.L_HI(net84));
 sg13g2_tiehi _3333__85 (.L_HI(net85));
 sg13g2_tiehi _3401__86 (.L_HI(net86));
 sg13g2_tiehi _3332__87 (.L_HI(net87));
 sg13g2_tiehi _3435__88 (.L_HI(net88));
 sg13g2_tiehi _3331__89 (.L_HI(net89));
 sg13g2_tiehi _3400__90 (.L_HI(net90));
 sg13g2_tiehi _3330__91 (.L_HI(net91));
 sg13g2_tiehi _3452__92 (.L_HI(net92));
 sg13g2_tiehi _3329__93 (.L_HI(net93));
 sg13g2_tiehi _3399__94 (.L_HI(net94));
 sg13g2_tiehi _3328__95 (.L_HI(net95));
 sg13g2_tiehi _3434__96 (.L_HI(net96));
 sg13g2_tiehi _3327__97 (.L_HI(net97));
 sg13g2_tiehi _3398__98 (.L_HI(net98));
 sg13g2_tiehi _3326__99 (.L_HI(net99));
 sg13g2_tiehi _3465__100 (.L_HI(net100));
 sg13g2_tiehi _3325__101 (.L_HI(net101));
 sg13g2_tiehi _3397__102 (.L_HI(net102));
 sg13g2_tiehi _3324__103 (.L_HI(net103));
 sg13g2_tiehi _3433__104 (.L_HI(net104));
 sg13g2_tiehi _3323__105 (.L_HI(net105));
 sg13g2_tiehi _3396__106 (.L_HI(net106));
 sg13g2_tiehi _3322__107 (.L_HI(net107));
 sg13g2_tiehi _3451__108 (.L_HI(net108));
 sg13g2_tiehi _3321__109 (.L_HI(net109));
 sg13g2_tiehi _3395__110 (.L_HI(net110));
 sg13g2_tiehi _3320__111 (.L_HI(net111));
 sg13g2_tiehi _3432__112 (.L_HI(net112));
 sg13g2_tiehi _3319__113 (.L_HI(net113));
 sg13g2_tiehi _3394__114 (.L_HI(net114));
 sg13g2_tiehi _3318__115 (.L_HI(net115));
 sg13g2_tiehi _3460__116 (.L_HI(net116));
 sg13g2_tiehi _3317__117 (.L_HI(net117));
 sg13g2_tiehi _3393__118 (.L_HI(net118));
 sg13g2_tiehi _3316__119 (.L_HI(net119));
 sg13g2_tiehi _3431__120 (.L_HI(net120));
 sg13g2_tiehi _3315__121 (.L_HI(net121));
 sg13g2_tiehi _3392__122 (.L_HI(net122));
 sg13g2_tiehi _3314__123 (.L_HI(net123));
 sg13g2_tiehi _3450__124 (.L_HI(net124));
 sg13g2_tiehi _3313__125 (.L_HI(net125));
 sg13g2_tiehi _3391__126 (.L_HI(net126));
 sg13g2_tiehi _3312__127 (.L_HI(net127));
 sg13g2_tiehi _3430__128 (.L_HI(net128));
 sg13g2_tiehi _3311__129 (.L_HI(net129));
 sg13g2_tiehi _3390__130 (.L_HI(net130));
 sg13g2_tiehi _3310__131 (.L_HI(net131));
 sg13g2_tiehi _3467__132 (.L_HI(net132));
 sg13g2_tiehi _3309__133 (.L_HI(net133));
 sg13g2_tiehi _3389__134 (.L_HI(net134));
 sg13g2_tiehi _3308__135 (.L_HI(net135));
 sg13g2_tiehi _3429__136 (.L_HI(net136));
 sg13g2_tiehi _3307__137 (.L_HI(net137));
 sg13g2_tiehi _3388__138 (.L_HI(net138));
 sg13g2_tiehi _3306__139 (.L_HI(net139));
 sg13g2_tiehi _3449__140 (.L_HI(net140));
 sg13g2_tiehi _3305__141 (.L_HI(net141));
 sg13g2_tiehi _3387__142 (.L_HI(net142));
 sg13g2_tiehi _3304__143 (.L_HI(net143));
 sg13g2_tiehi _3428__144 (.L_HI(net144));
 sg13g2_tiehi _3303__145 (.L_HI(net145));
 sg13g2_tiehi _3386__146 (.L_HI(net146));
 sg13g2_tiehi _3302__147 (.L_HI(net147));
 sg13g2_tiehi _3459__148 (.L_HI(net148));
 sg13g2_tiehi _3301__149 (.L_HI(net149));
 sg13g2_tiehi _3385__150 (.L_HI(net150));
 sg13g2_tiehi _3300__151 (.L_HI(net151));
 sg13g2_tiehi _3427__152 (.L_HI(net152));
 sg13g2_tiehi _3299__153 (.L_HI(net153));
 sg13g2_tiehi _3384__154 (.L_HI(net154));
 sg13g2_tiehi _3298__155 (.L_HI(net155));
 sg13g2_tiehi _3448__156 (.L_HI(net156));
 sg13g2_tiehi _3297__157 (.L_HI(net157));
 sg13g2_tiehi _3383__158 (.L_HI(net158));
 sg13g2_tiehi _3296__159 (.L_HI(net159));
 sg13g2_tiehi _3426__160 (.L_HI(net160));
 sg13g2_tiehi _3295__161 (.L_HI(net161));
 sg13g2_tiehi _3382__162 (.L_HI(net162));
 sg13g2_tiehi _3294__163 (.L_HI(net163));
 sg13g2_tiehi _3464__164 (.L_HI(net164));
 sg13g2_tiehi _3293__165 (.L_HI(net165));
 sg13g2_tiehi _3381__166 (.L_HI(net166));
 sg13g2_tiehi _3292__167 (.L_HI(net167));
 sg13g2_tiehi _3425__168 (.L_HI(net168));
 sg13g2_tiehi _3291__169 (.L_HI(net169));
 sg13g2_tiehi _3380__170 (.L_HI(net170));
 sg13g2_tiehi _3290__171 (.L_HI(net171));
 sg13g2_tiehi _3447__172 (.L_HI(net172));
 sg13g2_tiehi _3289__173 (.L_HI(net173));
 sg13g2_tiehi _3379__174 (.L_HI(net174));
 sg13g2_tiehi _3288__175 (.L_HI(net175));
 sg13g2_tiehi _3424__176 (.L_HI(net176));
 sg13g2_tiehi _3287__177 (.L_HI(net177));
 sg13g2_tiehi _3378__178 (.L_HI(net178));
 sg13g2_tiehi _3286__179 (.L_HI(net179));
 sg13g2_tiehi _3458__180 (.L_HI(net180));
 sg13g2_tiehi _3285__181 (.L_HI(net181));
 sg13g2_tiehi _3377__182 (.L_HI(net182));
 sg13g2_tiehi _3284__183 (.L_HI(net183));
 sg13g2_tiehi _3423__184 (.L_HI(net184));
 sg13g2_tiehi _3283__185 (.L_HI(net185));
 sg13g2_tiehi _3376__186 (.L_HI(net186));
 sg13g2_tiehi _3282__187 (.L_HI(net187));
 sg13g2_tiehi _3278__188 (.L_HI(net188));
 sg13g2_tiehi _3446__189 (.L_HI(net189));
 sg13g2_tiehi _3277__190 (.L_HI(net190));
 sg13g2_tiehi _3375__191 (.L_HI(net191));
 sg13g2_tiehi _3276__192 (.L_HI(net192));
 sg13g2_tiehi _3422__193 (.L_HI(net193));
 sg13g2_tiehi _3275__194 (.L_HI(net194));
 sg13g2_tiehi _3374__195 (.L_HI(net195));
 sg13g2_tiehi _3274__196 (.L_HI(net196));
 sg13g2_tiehi _3468__197 (.L_HI(net197));
 sg13g2_tiehi _3273__198 (.L_HI(net198));
 sg13g2_tiehi _3373__199 (.L_HI(net199));
 sg13g2_tiehi _3272__200 (.L_HI(net200));
 sg13g2_tiehi _3421__201 (.L_HI(net201));
 sg13g2_tiehi _3271__202 (.L_HI(net202));
 sg13g2_tiehi _3372__203 (.L_HI(net203));
 sg13g2_tiehi _3270__204 (.L_HI(net204));
 sg13g2_tiehi _3445__205 (.L_HI(net205));
 sg13g2_tiehi _3269__206 (.L_HI(net206));
 sg13g2_tiehi _3371__207 (.L_HI(net207));
 sg13g2_tiehi _3268__208 (.L_HI(net208));
 sg13g2_tiehi _3420__209 (.L_HI(net209));
 sg13g2_tiehi _3267__210 (.L_HI(net210));
 sg13g2_tiehi _3370__211 (.L_HI(net211));
 sg13g2_tiehi _3266__212 (.L_HI(net212));
 sg13g2_tiehi _3457__213 (.L_HI(net213));
 sg13g2_tiehi _3265__214 (.L_HI(net214));
 sg13g2_tiehi _3369__215 (.L_HI(net215));
 sg13g2_tiehi _3264__216 (.L_HI(net216));
 sg13g2_tiehi _3419__217 (.L_HI(net217));
 sg13g2_tiehi _3263__218 (.L_HI(net218));
 sg13g2_tiehi _3368__219 (.L_HI(net219));
 sg13g2_tiehi _3262__220 (.L_HI(net220));
 sg13g2_tiehi _3261__221 (.L_HI(net221));
 sg13g2_tiehi _3260__222 (.L_HI(net222));
 sg13g2_tiehi _3259__223 (.L_HI(net223));
 sg13g2_tiehi _3258__224 (.L_HI(net224));
 sg13g2_tiehi _3257__225 (.L_HI(net225));
 sg13g2_tiehi _3256__226 (.L_HI(net226));
 sg13g2_tiehi _3255__227 (.L_HI(net227));
 sg13g2_tiehi _3254__228 (.L_HI(net228));
 sg13g2_tiehi _3253__229 (.L_HI(net229));
 sg13g2_tiehi _3252__230 (.L_HI(net230));
 sg13g2_tiehi _3251__231 (.L_HI(net231));
 sg13g2_tiehi _3250__232 (.L_HI(net232));
 sg13g2_tiehi _3249__233 (.L_HI(net233));
 sg13g2_tiehi _3248__234 (.L_HI(net234));
 sg13g2_tiehi _3247__235 (.L_HI(net235));
 sg13g2_tiehi _3246__236 (.L_HI(net236));
 sg13g2_tiehi _3245__237 (.L_HI(net237));
 sg13g2_tiehi _3244__238 (.L_HI(net238));
 sg13g2_tiehi _3444__239 (.L_HI(net239));
 sg13g2_tiehi _3367__240 (.L_HI(net240));
 sg13g2_tiehi _3418__241 (.L_HI(net241));
 sg13g2_tiehi _3366__242 (.L_HI(net242));
 sg13g2_tiehi _3463__243 (.L_HI(net243));
 sg13g2_tiehi _3365__244 (.L_HI(net244));
 sg13g2_tiehi _3417__245 (.L_HI(net245));
 sg13g2_tiehi _3364__246 (.L_HI(net246));
 sg13g2_tiehi _3443__247 (.L_HI(net247));
 sg13g2_tiehi _3363__248 (.L_HI(net248));
 sg13g2_tiehi _3416__249 (.L_HI(net249));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_wokwi_413387065339458561_3 (.L_LO(net3));
 sg13g2_tielo tt_um_wokwi_413387065339458561_4 (.L_LO(net4));
 sg13g2_tielo tt_um_wokwi_413387065339458561_5 (.L_LO(net5));
 sg13g2_tielo tt_um_wokwi_413387065339458561_6 (.L_LO(net6));
 sg13g2_tielo tt_um_wokwi_413387065339458561_7 (.L_LO(net7));
 sg13g2_tielo tt_um_wokwi_413387065339458561_8 (.L_LO(net8));
 sg13g2_tielo tt_um_wokwi_413387065339458561_9 (.L_LO(net9));
 sg13g2_tielo tt_um_wokwi_413387065339458561_10 (.L_LO(net10));
 sg13g2_tielo tt_um_wokwi_413387065339458561_11 (.L_LO(net11));
 sg13g2_tielo tt_um_wokwi_413387065339458561_12 (.L_LO(net12));
 sg13g2_tielo tt_um_wokwi_413387065339458561_13 (.L_LO(net13));
 sg13g2_tielo tt_um_wokwi_413387065339458561_14 (.L_LO(net14));
 sg13g2_tielo tt_um_wokwi_413387065339458561_15 (.L_LO(net15));
 sg13g2_tielo tt_um_wokwi_413387065339458561_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_413387065339458561_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_413387065339458561_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_413387065339458561_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_413387065339458561_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_413387065339458561_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_413387065339458561_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_413387065339458561_23 (.L_LO(net23));
 sg13g2_tiehi _3362__24 (.L_HI(net24));
 sg13g2_buf_4 _3717_ (.X(uo_out[0]),
    .A(\ws2812_out.led_o ));
 sg13g2_buf_1 _3718_ (.A(\uart_output.uart_out ),
    .X(uo_out[1]));
 sg13g2_buf_2 fanout757 (.A(net759),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_4 fanout759 (.X(net759),
    .A(_0835_));
 sg13g2_buf_2 fanout760 (.A(net761),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(net762),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_0640_),
    .X(net762));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(net764));
 sg13g2_buf_2 fanout764 (.A(_0640_),
    .X(net764));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(_0487_));
 sg13g2_buf_4 fanout766 (.X(net766),
    .A(net768));
 sg13g2_buf_2 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(_0285_));
 sg13g2_buf_4 fanout769 (.X(net769),
    .A(net770));
 sg13g2_buf_2 fanout770 (.A(_0285_),
    .X(net770));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(net773));
 sg13g2_buf_2 fanout772 (.A(net773),
    .X(net772));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(_0262_));
 sg13g2_buf_2 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_0262_),
    .X(net775));
 sg13g2_buf_4 fanout776 (.X(net776),
    .A(_1359_));
 sg13g2_buf_2 fanout777 (.A(_1355_),
    .X(net777));
 sg13g2_buf_4 fanout778 (.X(net778),
    .A(_0830_));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(net780));
 sg13g2_buf_4 fanout780 (.X(net780),
    .A(net784));
 sg13g2_buf_2 fanout781 (.A(net783),
    .X(net781));
 sg13g2_buf_1 fanout782 (.A(net783),
    .X(net782));
 sg13g2_buf_4 fanout783 (.X(net783),
    .A(net784));
 sg13g2_buf_2 fanout784 (.A(_0634_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(net787),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(net789),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(net789),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_0633_),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(net793));
 sg13g2_buf_4 fanout791 (.X(net791),
    .A(net793));
 sg13g2_buf_2 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_0633_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_4 fanout795 (.X(net795),
    .A(net797));
 sg13g2_buf_4 fanout796 (.X(net796),
    .A(net797));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(_0271_));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(_0270_));
 sg13g2_buf_2 fanout799 (.A(_0270_),
    .X(net799));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(net801));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(_0270_));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(_1358_));
 sg13g2_buf_2 fanout803 (.A(net804),
    .X(net803));
 sg13g2_buf_8 fanout804 (.A(_1358_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(net807),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(net807),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(net808),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(net829),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(net811),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(net811),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(net829),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(net814),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(net814),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(net817),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(net816),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(net817),
    .X(net816));
 sg13g2_buf_1 fanout817 (.A(net829),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(net821),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(net820),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(net821),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(net829),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(net825),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(net825),
    .X(net823));
 sg13g2_buf_1 fanout824 (.A(net825),
    .X(net824));
 sg13g2_buf_1 fanout825 (.A(net829),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(net827),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(net828),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(net829),
    .X(net828));
 sg13g2_buf_4 fanout829 (.X(net829),
    .A(_1357_));
 sg13g2_buf_2 fanout830 (.A(_0304_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(net837),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(net834),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(net837),
    .X(net834));
 sg13g2_buf_4 fanout835 (.X(net835),
    .A(net837));
 sg13g2_buf_2 fanout836 (.A(net837),
    .X(net836));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(_0258_));
 sg13g2_buf_2 fanout838 (.A(net839),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(net841),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_1 fanout841 (.A(net845),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(net845),
    .X(net842));
 sg13g2_buf_4 fanout843 (.X(net843),
    .A(net844));
 sg13g2_buf_2 fanout844 (.A(net845),
    .X(net844));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(_0257_));
 sg13g2_buf_2 fanout846 (.A(net847),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(net848),
    .X(net847));
 sg13g2_buf_4 fanout848 (.X(net848),
    .A(_1398_));
 sg13g2_buf_4 fanout849 (.X(net849),
    .A(net850));
 sg13g2_buf_4 fanout850 (.X(net850),
    .A(_1398_));
 sg13g2_buf_2 fanout851 (.A(net853),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_4 fanout853 (.X(net853),
    .A(net856));
 sg13g2_buf_4 fanout854 (.X(net854),
    .A(net856));
 sg13g2_buf_4 fanout855 (.X(net855),
    .A(net856));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(_1397_));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(_1392_));
 sg13g2_buf_1 fanout858 (.A(_1392_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(net862),
    .X(net861));
 sg13g2_buf_4 fanout862 (.X(net862),
    .A(_1391_));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(_1377_));
 sg13g2_buf_4 fanout864 (.X(net864),
    .A(net865));
 sg13g2_buf_2 fanout865 (.A(_1376_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(net867),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net871),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(net869),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(net871),
    .X(net869));
 sg13g2_buf_4 fanout870 (.X(net870),
    .A(net871));
 sg13g2_buf_4 fanout871 (.X(net871),
    .A(_1382_));
 sg13g2_buf_2 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(net874),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net878),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(net878),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(net878),
    .X(net876));
 sg13g2_buf_4 fanout877 (.X(net877),
    .A(net878));
 sg13g2_buf_4 fanout878 (.X(net878),
    .A(_1381_));
 sg13g2_buf_4 fanout879 (.X(net879),
    .A(net881));
 sg13g2_buf_4 fanout880 (.X(net880),
    .A(net881));
 sg13g2_buf_2 fanout881 (.A(_1011_),
    .X(net881));
 sg13g2_buf_4 fanout882 (.X(net882),
    .A(_1009_));
 sg13g2_buf_4 fanout883 (.X(net883),
    .A(_1006_));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(_1006_));
 sg13g2_buf_4 fanout885 (.X(net885),
    .A(net887));
 sg13g2_buf_4 fanout886 (.X(net886),
    .A(net887));
 sg13g2_buf_2 fanout887 (.A(_1003_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(net889),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(net899),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(net893),
    .X(net891));
 sg13g2_buf_1 fanout892 (.A(net893),
    .X(net892));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(net899));
 sg13g2_buf_2 fanout894 (.A(net898),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(net898),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(net897),
    .X(net896));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(net898));
 sg13g2_buf_4 fanout898 (.X(net898),
    .A(net899));
 sg13g2_buf_2 fanout899 (.A(_0972_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(net901),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(net903),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(net903),
    .X(net902));
 sg13g2_buf_1 fanout903 (.A(net904),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(net905),
    .X(net904));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(\spi_in.index[5] ));
 sg13g2_buf_2 fanout906 (.A(net909),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(net909),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(net909),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(_0022_),
    .X(net909));
 sg13g2_buf_4 fanout910 (.X(net910),
    .A(net914));
 sg13g2_buf_2 fanout911 (.A(net914),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(net913),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(net914),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(\spi_in.index[3] ),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(net916),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_0021_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(net512),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(net919),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(net920),
    .X(net919));
 sg13g2_buf_1 fanout920 (.A(net923),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(net923),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(net923),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(net936),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(net925),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(net936),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(net936),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(net928),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(net936),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(net936),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(net932),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(net932),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(net935),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(net935),
    .X(net933));
 sg13g2_buf_1 fanout934 (.A(net935),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(net936),
    .X(net935));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(\spi_in.state[2] ));
 sg13g2_buf_2 fanout937 (.A(net938),
    .X(net937));
 sg13g2_buf_1 fanout938 (.A(net513),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_1 fanout940 (.A(\uart_output.index[3] ),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(net942),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(net943),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(\uart_output.index[2] ),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(\uart_output.index[1] ),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(net946),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(\uart_output.index[0] ),
    .X(net946));
 sg13g2_buf_4 fanout947 (.X(net947),
    .A(net948));
 sg13g2_buf_4 fanout948 (.X(net948),
    .A(\ws2812_out.datacounter[3] ));
 sg13g2_buf_4 fanout949 (.X(net949),
    .A(net950));
 sg13g2_buf_2 fanout950 (.A(net951),
    .X(net950));
 sg13g2_buf_4 fanout951 (.X(net951),
    .A(net515));
 sg13g2_buf_4 fanout952 (.X(net952),
    .A(net953));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(net955));
 sg13g2_buf_4 fanout954 (.X(net954),
    .A(net955));
 sg13g2_buf_4 fanout955 (.X(net955),
    .A(\ws2812_out.datacounter[1] ));
 sg13g2_buf_2 fanout956 (.A(net957),
    .X(net956));
 sg13g2_buf_4 fanout957 (.X(net957),
    .A(net958));
 sg13g2_buf_2 fanout958 (.A(net959),
    .X(net958));
 sg13g2_buf_4 fanout959 (.X(net959),
    .A(\ws2812_out.datacounter[0] ));
 sg13g2_buf_4 fanout960 (.X(net960),
    .A(net961));
 sg13g2_buf_4 fanout961 (.X(net961),
    .A(\ws2812_out.datacounter[0] ));
 sg13g2_buf_2 fanout962 (.A(net964),
    .X(net962));
 sg13g2_buf_4 fanout963 (.X(net963),
    .A(net964));
 sg13g2_buf_1 fanout964 (.A(net969),
    .X(net964));
 sg13g2_buf_4 fanout965 (.X(net965),
    .A(net969));
 sg13g2_buf_1 fanout966 (.A(net969),
    .X(net966));
 sg13g2_buf_4 fanout967 (.X(net967),
    .A(net969));
 sg13g2_buf_4 fanout968 (.X(net968),
    .A(net969));
 sg13g2_buf_4 fanout969 (.X(net969),
    .A(\ws2812_out.datacounter[0] ));
 sg13g2_buf_2 fanout970 (.A(net972),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(net972),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(net978),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(net977),
    .X(net973));
 sg13g2_buf_1 fanout974 (.A(net977),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(net977),
    .X(net975));
 sg13g2_buf_1 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(net978),
    .X(net977));
 sg13g2_buf_1 fanout978 (.A(_0974_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(net981),
    .X(net979));
 sg13g2_buf_1 fanout980 (.A(net981),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(net984),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(net983),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(net984),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_0974_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(net986),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(net999),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(net990),
    .X(net987));
 sg13g2_buf_1 fanout988 (.A(net990),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(net990),
    .X(net989));
 sg13g2_buf_1 fanout990 (.A(net999),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(net998),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(net993),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(net998),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(net997),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(net997),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(net997),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(net998),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(net999),
    .X(net998));
 sg13g2_buf_1 fanout999 (.A(_0974_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(net1001),
    .X(net1000));
 sg13g2_buf_4 fanout1001 (.X(net1001),
    .A(net1002));
 sg13g2_buf_4 fanout1002 (.X(net1002),
    .A(ui_in[1]));
 sg13g2_buf_2 fanout1003 (.A(net1004),
    .X(net1003));
 sg13g2_buf_4 fanout1004 (.X(net1004),
    .A(net1007));
 sg13g2_buf_2 fanout1005 (.A(net1007),
    .X(net1005));
 sg13g2_buf_4 fanout1006 (.X(net1006),
    .A(net1007));
 sg13g2_buf_2 fanout1007 (.A(rst_n),
    .X(net1007));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_tielo tt_um_wokwi_413387065339458561_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_29_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_24_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_18_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_9_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_11_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0023_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold2 (.A(\pixel_4[0] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold3 (.A(\pixel_5[8] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold4 (.A(\pixel_1[17] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold5 (.A(\pixel_1[12] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold6 (.A(\pixel_2[6] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold7 (.A(\pixel_2[8] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold8 (.A(\pixel_3[9] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold9 (.A(\pixel_2[18] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold10 (.A(\pixel_6[8] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold11 (.A(\pixel_0[9] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold12 (.A(\pixel_0[0] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold13 (.A(\pixel_2[11] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold14 (.A(\pixel_1[2] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold15 (.A(\pixel_2[3] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold16 (.A(\pixel_4[4] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold17 (.A(\pixel_0[4] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold18 (.A(\pixel_3[2] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold19 (.A(\pixel_1[8] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold20 (.A(\pixel_0[7] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold21 (.A(\pixel_4[19] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold22 (.A(\pixel_3[1] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold23 (.A(\pixel_4[5] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold24 (.A(\pixel_3[0] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold25 (.A(\pixel_2[5] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold26 (.A(\pixel_3[23] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold27 (.A(\pixel_4[16] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold28 (.A(\pixel_2[17] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold29 (.A(\pixel_0[21] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold30 (.A(\pixel_5[5] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold31 (.A(\pixel_0[1] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold32 (.A(\pixel_2[20] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold33 (.A(\pixel_0[19] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold34 (.A(\pixel_1[3] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold35 (.A(\spi_in.bit_count[8] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0077_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold37 (.A(\pixel_1[14] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold38 (.A(\pixel_1[6] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold39 (.A(\pixel_5[7] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold40 (.A(\pixel_2[0] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold41 (.A(\pixel_4[22] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold42 (.A(\pixel_3[3] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold43 (.A(\pixel_0[22] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold44 (.A(\pixel_3[19] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold45 (.A(\pixel_1[20] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold46 (.A(\pixel_2[19] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold47 (.A(\pixel_1[5] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold48 (.A(\pixel_1[23] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold49 (.A(\pixel_0[3] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold50 (.A(\pixel_3[18] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0018_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold52 (.A(_1225_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0034_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold54 (.A(\pixel_2[16] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold55 (.A(\pixel_2[23] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold56 (.A(\pixel_1[15] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold57 (.A(\pixel_2[13] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold58 (.A(\pixel_2[14] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold59 (.A(\pixel_1[19] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold60 (.A(\pixel_2[9] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold61 (.A(\pixel_2[7] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold62 (.A(\pixel_0[10] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold63 (.A(\pixel_6[4] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold64 (.A(\pixel_2[12] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold65 (.A(\pixel_3[13] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold66 (.A(\pixel_1[13] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold67 (.A(\pixel_2[21] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold68 (.A(\pixel_1[11] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold69 (.A(\pixel_6[16] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold70 (.A(\pixel_4[2] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold71 (.A(\pixel_0[15] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold72 (.A(\pixel_0[18] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold73 (.A(\pixel_2[1] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold74 (.A(\pixel_4[7] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold75 (.A(\pixel_3[11] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold76 (.A(\pixel_2[2] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold77 (.A(\pixel_3[10] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold78 (.A(\pixel_0[5] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold79 (.A(\pixel_5[13] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold80 (.A(\pixel_2[4] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold81 (.A(\pixel_5[21] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold82 (.A(\pixel_1[7] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold83 (.A(\pixel_0[13] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold84 (.A(\pixel_0[16] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold85 (.A(\pixel_3[6] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold86 (.A(\pixel_5[10] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold87 (.A(\pixel_6[22] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold88 (.A(\pixel_6[2] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0286_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold90 (.A(\pixel_3[4] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold91 (.A(\pixel_0[2] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold92 (.A(\pixel_0[14] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold93 (.A(\pixel_4[17] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0019_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold95 (.A(_1221_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold96 (.A(\pixel_0[6] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold97 (.A(\pixel_5[3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold98 (.A(\pixel_4[20] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold99 (.A(\pixel_5[16] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold100 (.A(\pixel_1[18] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold101 (.A(\pixel_0[17] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold102 (.A(\pixel_0[12] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold103 (.A(\pixel_4[18] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0641_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold105 (.A(\pixel_6[17] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold106 (.A(\uart_output.uart_out ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0060_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold108 (.A(\pixel_0[11] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold109 (.A(\pixel_5[12] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold110 (.A(\pixel_1[9] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold111 (.A(\pixel_6[6] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold112 (.A(\pixel_4[9] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold113 (.A(\pixel_3[7] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold114 (.A(\pixel_6[18] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold115 (.A(\pixel_5[17] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold116 (.A(\pixel_0[20] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold117 (.A(\pixel_6[1] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold118 (.A(\pixel_4[3] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold119 (.A(\pixel_5[14] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0012_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold121 (.A(_1208_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold122 (.A(\pixel_1[21] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold123 (.A(\pixel_1[1] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold124 (.A(\pixel_5[23] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold125 (.A(\pixel_2[10] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold126 (.A(\pixel_3[22] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold127 (.A(\pixel_6[7] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold128 (.A(\pixel_3[15] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold129 (.A(\pixel_4[23] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold130 (.A(\pixel_6[19] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold131 (.A(\pixel_4[1] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold132 (.A(\ws2812_out.counter[0] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold133 (.A(\pixel_4[21] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold134 (.A(\pixel_4[13] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold135 (.A(\uart_output.count[2] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold136 (.A(_1233_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0037_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold138 (.A(\ws2812_out.datacounter[7] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold139 (.A(_1265_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold140 (.A(\pixel_5[19] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold141 (.A(\pixel_6[23] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold142 (.A(\pixel_6[11] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold143 (.A(\pixel_5[1] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold144 (.A(\pixel_3[17] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0005_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0056_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold147 (.A(\pixel_4[8] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold148 (.A(\pixel_3[14] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold149 (.A(\uart_output.index[3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0054_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold151 (.A(\pixel_5[9] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold152 (.A(\uart_output.count[3] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold153 (.A(_1235_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold154 (.A(\pixel_5[20] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold155 (.A(\pixel_5[11] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold156 (.A(\pixel_4[14] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold157 (.A(\pixel_4[15] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold158 (.A(\pixel_6[5] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold159 (.A(\pixel_5[15] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold160 (.A(\pixel_2[15] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold161 (.A(\pixel_6[3] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold162 (.A(\uart_output.count[4] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold163 (.A(\pixel_3[5] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold164 (.A(\uart_output.count[6] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold165 (.A(_1240_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold166 (.A(\pixel_2[22] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold167 (.A(\pixel_4[6] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold168 (.A(\pixel_3[20] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold169 (.A(\spi_in.bit_count[2] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold170 (.A(_1408_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold171 (.A(\pixel_3[21] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold172 (.A(\pixel_4[11] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold173 (.A(\uart_output.index[1] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold174 (.A(\spi_in.bit_count[7] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0248_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold176 (.A(\pixel_5[2] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold177 (.A(\pixel_1[22] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold178 (.A(\pixel_4[10] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold179 (.A(\spi_in.index[4] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold180 (.A(\pixel_0[23] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold181 (.A(\pixel_1[10] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0836_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold183 (.A(\pixel_5[4] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold184 (.A(\pixel_3[12] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold185 (.A(\pixel_1[0] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold186 (.A(\uart_output.index[6] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0057_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0003_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1296_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0058_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold191 (.A(\pixel_6[15] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0011_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0049_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold194 (.A(\pixel_6[9] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0013_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold196 (.A(_1209_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0020_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0994_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0002_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold200 (.A(\pixel_5[6] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold201 (.A(\pixel_6[20] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold202 (.A(\pixel_6[10] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold203 (.A(\spi_in.bit_count[1] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold204 (.A(_1407_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0070_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold206 (.A(\pixel_6[14] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold207 (.A(\uart_output.count[5] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold208 (.A(\spi_in.bit_count[0] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0069_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold210 (.A(\uart_output.count[7] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold211 (.A(\pixel_6[21] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0014_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold213 (.A(_1211_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold214 (.A(\spi_in.bit_count[3] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold215 (.A(\pixel_5[18] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold216 (.A(\uart_output.count[1] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold217 (.A(_1231_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold218 (.A(\spi_in.bit_count[4] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold219 (.A(\ws2812_out.counter[5] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold220 (.A(_1216_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0029_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold222 (.A(\ws2812_out.counter[6] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0030_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold224 (.A(\spi_in.bit_count[6] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold225 (.A(_1415_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold226 (.A(\spi_in.state[1] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0001_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold228 (.A(\pixel_1[16] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0007_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0053_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold231 (.A(\ws2812_out.counter[7] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0010_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0047_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold234 (.A(\pixel_3[8] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold235 (.A(\spi_in.index[2] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0063_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold237 (.A(\pixel_5[22] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold238 (.A(\spi_in.index[6] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold239 (.A(\ws2812_out.counter[1] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold240 (.A(\spi_in.bit_count[5] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold241 (.A(\spi_in.state[0] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0996_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0000_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold244 (.A(\pixel_0[8] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold245 (.A(\pixel_6[12] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold246 (.A(\pixel_6[13] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold247 (.A(\spi_in.index[7] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0068_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold249 (.A(\pixel_5[0] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold250 (.A(\ws2812_out.datacounter[5] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0048_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold252 (.A(\pixel_1[4] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold253 (.A(\pixel_3[16] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0016_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold255 (.A(_1369_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0062_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold257 (.A(\pixel_6[0] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold258 (.A(\ws2812_out.state ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold259 (.A(\pixel_4[12] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold260 (.A(\ws2812_out.counter[9] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold261 (.A(_1223_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0033_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold263 (.A(\spi_in.index[0] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold264 (.A(\uart_output.index[4] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0055_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold266 (.A(\ws2812_out.datacounter[2] ),
    .X(net515));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_fill_1 FILLER_0_231 ();
 sg13g2_fill_2 FILLER_0_236 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_fill_1 FILLER_0_289 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_fill_1 FILLER_1_189 ();
 sg13g2_fill_2 FILLER_1_220 ();
 sg13g2_decap_8 FILLER_1_304 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_fill_2 FILLER_2_196 ();
 sg13g2_fill_1 FILLER_2_232 ();
 sg13g2_fill_2 FILLER_2_241 ();
 sg13g2_fill_2 FILLER_2_273 ();
 sg13g2_fill_1 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_fill_2 FILLER_3_189 ();
 sg13g2_fill_2 FILLER_3_247 ();
 sg13g2_fill_1 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_356 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_175 ();
 sg13g2_fill_2 FILLER_4_202 ();
 sg13g2_fill_1 FILLER_4_230 ();
 sg13g2_fill_1 FILLER_4_244 ();
 sg13g2_fill_2 FILLER_4_260 ();
 sg13g2_fill_1 FILLER_4_298 ();
 sg13g2_fill_1 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_4 FILLER_5_168 ();
 sg13g2_fill_2 FILLER_5_172 ();
 sg13g2_fill_1 FILLER_5_213 ();
 sg13g2_fill_1 FILLER_5_260 ();
 sg13g2_fill_2 FILLER_5_270 ();
 sg13g2_fill_1 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_4 FILLER_6_168 ();
 sg13g2_fill_1 FILLER_6_202 ();
 sg13g2_fill_2 FILLER_6_250 ();
 sg13g2_fill_2 FILLER_6_269 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_175 ();
 sg13g2_fill_2 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_277 ();
 sg13g2_fill_1 FILLER_7_286 ();
 sg13g2_fill_1 FILLER_7_295 ();
 sg13g2_fill_1 FILLER_7_305 ();
 sg13g2_fill_1 FILLER_7_316 ();
 sg13g2_fill_2 FILLER_7_322 ();
 sg13g2_fill_1 FILLER_7_342 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_4 FILLER_8_168 ();
 sg13g2_decap_4 FILLER_8_202 ();
 sg13g2_fill_2 FILLER_8_206 ();
 sg13g2_decap_8 FILLER_8_212 ();
 sg13g2_decap_8 FILLER_8_219 ();
 sg13g2_fill_2 FILLER_8_226 ();
 sg13g2_fill_1 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_233 ();
 sg13g2_fill_2 FILLER_8_240 ();
 sg13g2_fill_2 FILLER_8_277 ();
 sg13g2_fill_1 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_4 FILLER_8_291 ();
 sg13g2_fill_2 FILLER_8_304 ();
 sg13g2_fill_2 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_163 ();
 sg13g2_fill_2 FILLER_9_190 ();
 sg13g2_fill_1 FILLER_9_247 ();
 sg13g2_fill_2 FILLER_9_266 ();
 sg13g2_fill_1 FILLER_9_286 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_4 FILLER_10_154 ();
 sg13g2_fill_2 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_4 FILLER_11_147 ();
 sg13g2_fill_1 FILLER_11_173 ();
 sg13g2_fill_1 FILLER_11_209 ();
 sg13g2_fill_1 FILLER_11_227 ();
 sg13g2_fill_2 FILLER_11_276 ();
 sg13g2_fill_2 FILLER_11_289 ();
 sg13g2_fill_1 FILLER_11_291 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_fill_1 FILLER_12_161 ();
 sg13g2_fill_1 FILLER_12_193 ();
 sg13g2_decap_4 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_fill_2 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_291 ();
 sg13g2_fill_2 FILLER_12_319 ();
 sg13g2_fill_1 FILLER_12_321 ();
 sg13g2_fill_1 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_fill_2 FILLER_13_161 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_fill_1 FILLER_13_174 ();
 sg13g2_fill_2 FILLER_13_180 ();
 sg13g2_decap_4 FILLER_13_204 ();
 sg13g2_fill_2 FILLER_13_208 ();
 sg13g2_fill_2 FILLER_13_218 ();
 sg13g2_decap_8 FILLER_13_237 ();
 sg13g2_decap_8 FILLER_13_244 ();
 sg13g2_decap_4 FILLER_13_251 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_decap_4 FILLER_13_271 ();
 sg13g2_fill_2 FILLER_13_275 ();
 sg13g2_decap_8 FILLER_13_283 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_2 FILLER_13_296 ();
 sg13g2_fill_1 FILLER_13_298 ();
 sg13g2_fill_2 FILLER_13_305 ();
 sg13g2_fill_1 FILLER_13_307 ();
 sg13g2_fill_2 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_161 ();
 sg13g2_fill_2 FILLER_14_188 ();
 sg13g2_decap_4 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_239 ();
 sg13g2_fill_2 FILLER_14_245 ();
 sg13g2_fill_1 FILLER_14_257 ();
 sg13g2_fill_1 FILLER_14_266 ();
 sg13g2_fill_1 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_277 ();
 sg13g2_fill_2 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_fill_2 FILLER_14_297 ();
 sg13g2_fill_1 FILLER_14_299 ();
 sg13g2_fill_1 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_154 ();
 sg13g2_fill_1 FILLER_15_240 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_decap_4 FILLER_15_254 ();
 sg13g2_fill_2 FILLER_15_267 ();
 sg13g2_fill_2 FILLER_15_307 ();
 sg13g2_fill_1 FILLER_15_309 ();
 sg13g2_fill_1 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_161 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_fill_1 FILLER_16_227 ();
 sg13g2_fill_1 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_295 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_4 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_172 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_4 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_decap_8 FILLER_17_215 ();
 sg13g2_fill_2 FILLER_17_222 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_fill_1 FILLER_17_304 ();
 sg13g2_fill_2 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_fill_2 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_fill_2 FILLER_18_175 ();
 sg13g2_decap_4 FILLER_18_181 ();
 sg13g2_fill_2 FILLER_18_185 ();
 sg13g2_fill_1 FILLER_18_249 ();
 sg13g2_fill_2 FILLER_18_254 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_fill_2 FILLER_18_272 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_4 FILLER_19_161 ();
 sg13g2_fill_1 FILLER_19_165 ();
 sg13g2_fill_2 FILLER_19_215 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_253 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_fill_2 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_fill_2 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_211 ();
 sg13g2_decap_8 FILLER_20_218 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_decap_4 FILLER_20_263 ();
 sg13g2_fill_1 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_4 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_186 ();
 sg13g2_fill_2 FILLER_21_192 ();
 sg13g2_fill_1 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_220 ();
 sg13g2_decap_8 FILLER_21_227 ();
 sg13g2_decap_4 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_fill_1 FILLER_21_300 ();
 sg13g2_decap_4 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_4 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_211 ();
 sg13g2_decap_8 FILLER_22_227 ();
 sg13g2_decap_8 FILLER_22_234 ();
 sg13g2_fill_1 FILLER_22_261 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_269 ();
 sg13g2_fill_1 FILLER_22_278 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_decap_4 FILLER_22_313 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_337 ();
 sg13g2_fill_2 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_260 ();
 sg13g2_fill_1 FILLER_23_266 ();
 sg13g2_fill_2 FILLER_23_272 ();
 sg13g2_fill_1 FILLER_23_274 ();
 sg13g2_decap_4 FILLER_23_285 ();
 sg13g2_fill_2 FILLER_23_289 ();
 sg13g2_fill_2 FILLER_23_317 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_fill_1 FILLER_23_327 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_fill_2 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_245 ();
 sg13g2_fill_2 FILLER_24_260 ();
 sg13g2_fill_1 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_300 ();
 sg13g2_fill_2 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_335 ();
 sg13g2_fill_2 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_241 ();
 sg13g2_fill_1 FILLER_25_252 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_fill_2 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_4 FILLER_26_112 ();
 sg13g2_fill_2 FILLER_26_120 ();
 sg13g2_fill_1 FILLER_26_122 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_decap_8 FILLER_26_134 ();
 sg13g2_decap_8 FILLER_26_141 ();
 sg13g2_decap_8 FILLER_26_148 ();
 sg13g2_decap_8 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_fill_2 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_194 ();
 sg13g2_decap_4 FILLER_26_199 ();
 sg13g2_fill_1 FILLER_26_203 ();
 sg13g2_fill_1 FILLER_26_221 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_fill_2 FILLER_26_239 ();
 sg13g2_fill_1 FILLER_26_302 ();
 sg13g2_fill_1 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_131 ();
 sg13g2_decap_8 FILLER_27_136 ();
 sg13g2_decap_4 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_147 ();
 sg13g2_fill_2 FILLER_27_201 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_fill_2 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_2 FILLER_27_261 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_fill_2 FILLER_27_300 ();
 sg13g2_fill_2 FILLER_27_323 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_fill_2 FILLER_27_330 ();
 sg13g2_fill_1 FILLER_27_332 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_decap_8 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_4 FILLER_28_91 ();
 sg13g2_fill_2 FILLER_28_95 ();
 sg13g2_fill_2 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_178 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_fill_2 FILLER_28_239 ();
 sg13g2_fill_2 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_84 ();
 sg13g2_fill_1 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_148 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_2 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_217 ();
 sg13g2_fill_2 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_282 ();
 sg13g2_fill_2 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_91 ();
 sg13g2_fill_2 FILLER_30_118 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_decap_4 FILLER_30_194 ();
 sg13g2_fill_2 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_281 ();
 sg13g2_fill_2 FILLER_30_293 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_320 ();
 sg13g2_fill_2 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_341 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_4 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_188 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_227 ();
 sg13g2_fill_2 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_286 ();
 sg13g2_fill_2 FILLER_31_293 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_fill_2 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_339 ();
 sg13g2_decap_8 FILLER_31_375 ();
 sg13g2_decap_8 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_31_389 ();
 sg13g2_decap_8 FILLER_31_396 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_fill_2 FILLER_32_139 ();
 sg13g2_fill_1 FILLER_32_141 ();
 sg13g2_fill_1 FILLER_32_167 ();
 sg13g2_decap_4 FILLER_32_194 ();
 sg13g2_decap_4 FILLER_32_209 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_decap_4 FILLER_32_225 ();
 sg13g2_decap_4 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_241 ();
 sg13g2_decap_8 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_255 ();
 sg13g2_decap_8 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_fill_2 FILLER_32_315 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_fill_1 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_156 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_decap_8 FILLER_33_171 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_decap_4 FILLER_33_188 ();
 sg13g2_fill_2 FILLER_33_192 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_fill_2 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_244 ();
 sg13g2_fill_2 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_fill_2 FILLER_33_275 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_fill_1 FILLER_33_362 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_4 FILLER_34_98 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_2 FILLER_34_117 ();
 sg13g2_fill_1 FILLER_34_124 ();
 sg13g2_fill_2 FILLER_34_150 ();
 sg13g2_fill_2 FILLER_34_178 ();
 sg13g2_fill_2 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_fill_1 FILLER_34_258 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_decap_4 FILLER_34_295 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_4 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_102 ();
 sg13g2_fill_1 FILLER_35_175 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_2 FILLER_35_283 ();
 sg13g2_decap_8 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_321 ();
 sg13g2_fill_1 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_349 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_4 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_202 ();
 sg13g2_fill_1 FILLER_36_209 ();
 sg13g2_fill_1 FILLER_36_216 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_fill_2 FILLER_36_236 ();
 sg13g2_fill_1 FILLER_36_238 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_decap_4 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_decap_4 FILLER_36_303 ();
 sg13g2_fill_2 FILLER_36_307 ();
 sg13g2_decap_4 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_86 ();
 sg13g2_fill_2 FILLER_37_108 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_fill_2 FILLER_37_219 ();
 sg13g2_fill_1 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_294 ();
 sg13g2_decap_4 FILLER_37_308 ();
 sg13g2_fill_1 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_136 ();
 sg13g2_fill_1 FILLER_38_138 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_4 FILLER_38_201 ();
 sg13g2_fill_1 FILLER_38_205 ();
 sg13g2_decap_4 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_fill_2 FILLER_38_247 ();
 sg13g2_fill_2 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_290 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_fill_2 FILLER_38_320 ();
 sg13g2_fill_1 FILLER_38_332 ();
 sg13g2_fill_2 FILLER_38_339 ();
 sg13g2_fill_2 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_fill_1 FILLER_39_121 ();
 sg13g2_fill_1 FILLER_39_127 ();
 sg13g2_fill_1 FILLER_39_158 ();
 sg13g2_fill_2 FILLER_39_187 ();
 sg13g2_decap_4 FILLER_39_204 ();
 sg13g2_decap_8 FILLER_39_233 ();
 sg13g2_decap_4 FILLER_39_240 ();
 sg13g2_fill_1 FILLER_39_244 ();
 sg13g2_decap_4 FILLER_39_249 ();
 sg13g2_fill_2 FILLER_39_253 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_fill_2 FILLER_39_267 ();
 sg13g2_fill_1 FILLER_39_269 ();
 sg13g2_decap_8 FILLER_39_375 ();
 sg13g2_decap_8 FILLER_39_382 ();
 sg13g2_decap_8 FILLER_39_389 ();
 sg13g2_decap_8 FILLER_39_396 ();
 sg13g2_decap_4 FILLER_39_403 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_fill_1 FILLER_40_91 ();
 sg13g2_fill_1 FILLER_40_124 ();
 sg13g2_fill_2 FILLER_40_155 ();
 sg13g2_decap_8 FILLER_40_202 ();
 sg13g2_fill_2 FILLER_40_209 ();
 sg13g2_fill_1 FILLER_40_211 ();
 sg13g2_decap_8 FILLER_40_225 ();
 sg13g2_decap_4 FILLER_40_232 ();
 sg13g2_fill_1 FILLER_40_236 ();
 sg13g2_decap_4 FILLER_40_242 ();
 sg13g2_fill_1 FILLER_40_246 ();
 sg13g2_decap_4 FILLER_40_260 ();
 sg13g2_fill_2 FILLER_40_264 ();
 sg13g2_fill_1 FILLER_40_338 ();
 sg13g2_fill_1 FILLER_40_344 ();
 sg13g2_fill_1 FILLER_40_350 ();
 sg13g2_fill_2 FILLER_40_359 ();
 sg13g2_fill_1 FILLER_40_361 ();
 sg13g2_decap_8 FILLER_40_366 ();
 sg13g2_decap_8 FILLER_40_373 ();
 sg13g2_decap_8 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_40_387 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_4 FILLER_41_91 ();
 sg13g2_fill_2 FILLER_41_95 ();
 sg13g2_fill_1 FILLER_41_131 ();
 sg13g2_fill_1 FILLER_41_158 ();
 sg13g2_decap_8 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_218 ();
 sg13g2_decap_4 FILLER_41_225 ();
 sg13g2_decap_8 FILLER_41_256 ();
 sg13g2_fill_1 FILLER_41_263 ();
 sg13g2_decap_8 FILLER_41_272 ();
 sg13g2_decap_8 FILLER_41_279 ();
 sg13g2_fill_1 FILLER_41_286 ();
 sg13g2_fill_1 FILLER_41_294 ();
 sg13g2_decap_4 FILLER_41_306 ();
 sg13g2_decap_8 FILLER_41_326 ();
 sg13g2_decap_8 FILLER_41_333 ();
 sg13g2_decap_8 FILLER_41_340 ();
 sg13g2_decap_8 FILLER_41_347 ();
 sg13g2_fill_2 FILLER_41_354 ();
 sg13g2_fill_1 FILLER_41_356 ();
 sg13g2_fill_2 FILLER_41_361 ();
 sg13g2_decap_8 FILLER_41_389 ();
 sg13g2_decap_8 FILLER_41_396 ();
 sg13g2_decap_4 FILLER_41_403 ();
 sg13g2_fill_2 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_4 FILLER_42_98 ();
 sg13g2_fill_2 FILLER_42_102 ();
 sg13g2_fill_2 FILLER_42_138 ();
 sg13g2_decap_8 FILLER_42_144 ();
 sg13g2_decap_8 FILLER_42_151 ();
 sg13g2_decap_8 FILLER_42_158 ();
 sg13g2_fill_2 FILLER_42_165 ();
 sg13g2_fill_1 FILLER_42_175 ();
 sg13g2_decap_4 FILLER_42_190 ();
 sg13g2_fill_2 FILLER_42_199 ();
 sg13g2_fill_2 FILLER_42_247 ();
 sg13g2_decap_8 FILLER_42_262 ();
 sg13g2_decap_8 FILLER_42_269 ();
 sg13g2_decap_8 FILLER_42_276 ();
 sg13g2_decap_8 FILLER_42_283 ();
 sg13g2_fill_2 FILLER_42_290 ();
 sg13g2_decap_4 FILLER_42_298 ();
 sg13g2_fill_1 FILLER_42_302 ();
 sg13g2_decap_8 FILLER_42_307 ();
 sg13g2_decap_8 FILLER_42_314 ();
 sg13g2_decap_8 FILLER_42_321 ();
 sg13g2_fill_1 FILLER_42_328 ();
 sg13g2_fill_2 FILLER_42_333 ();
 sg13g2_fill_1 FILLER_42_335 ();
 sg13g2_fill_1 FILLER_42_365 ();
 sg13g2_decap_8 FILLER_42_379 ();
 sg13g2_decap_8 FILLER_42_386 ();
 sg13g2_decap_8 FILLER_42_393 ();
 sg13g2_decap_8 FILLER_42_400 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_fill_2 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_137 ();
 sg13g2_decap_4 FILLER_43_144 ();
 sg13g2_fill_2 FILLER_43_148 ();
 sg13g2_decap_8 FILLER_43_158 ();
 sg13g2_decap_8 FILLER_43_165 ();
 sg13g2_decap_8 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_179 ();
 sg13g2_fill_1 FILLER_43_201 ();
 sg13g2_fill_2 FILLER_43_287 ();
 sg13g2_fill_1 FILLER_43_289 ();
 sg13g2_fill_2 FILLER_43_298 ();
 sg13g2_fill_1 FILLER_43_300 ();
 sg13g2_fill_2 FILLER_43_328 ();
 sg13g2_fill_1 FILLER_43_330 ();
 sg13g2_fill_2 FILLER_43_337 ();
 sg13g2_fill_1 FILLER_43_339 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_4 FILLER_44_112 ();
 sg13g2_fill_2 FILLER_44_120 ();
 sg13g2_fill_1 FILLER_44_122 ();
 sg13g2_fill_1 FILLER_44_127 ();
 sg13g2_decap_8 FILLER_44_164 ();
 sg13g2_fill_1 FILLER_44_209 ();
 sg13g2_fill_1 FILLER_44_229 ();
 sg13g2_fill_1 FILLER_44_314 ();
 sg13g2_fill_2 FILLER_44_339 ();
 sg13g2_fill_1 FILLER_44_341 ();
 sg13g2_fill_1 FILLER_44_351 ();
 sg13g2_decap_8 FILLER_44_400 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_4 FILLER_45_126 ();
 sg13g2_fill_1 FILLER_45_130 ();
 sg13g2_decap_8 FILLER_45_174 ();
 sg13g2_fill_1 FILLER_45_181 ();
 sg13g2_fill_1 FILLER_45_206 ();
 sg13g2_fill_2 FILLER_45_212 ();
 sg13g2_fill_2 FILLER_45_219 ();
 sg13g2_fill_2 FILLER_45_264 ();
 sg13g2_fill_2 FILLER_45_316 ();
 sg13g2_decap_4 FILLER_45_326 ();
 sg13g2_decap_8 FILLER_45_397 ();
 sg13g2_decap_4 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_fill_1 FILLER_46_126 ();
 sg13g2_fill_2 FILLER_46_132 ();
 sg13g2_fill_2 FILLER_46_166 ();
 sg13g2_fill_1 FILLER_46_199 ();
 sg13g2_decap_8 FILLER_46_209 ();
 sg13g2_decap_8 FILLER_46_216 ();
 sg13g2_fill_2 FILLER_46_223 ();
 sg13g2_fill_1 FILLER_46_262 ();
 sg13g2_fill_1 FILLER_46_282 ();
 sg13g2_decap_8 FILLER_46_307 ();
 sg13g2_fill_2 FILLER_46_314 ();
 sg13g2_fill_1 FILLER_46_325 ();
 sg13g2_fill_2 FILLER_46_331 ();
 sg13g2_fill_2 FILLER_46_368 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_fill_2 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_139 ();
 sg13g2_decap_4 FILLER_47_146 ();
 sg13g2_fill_2 FILLER_47_150 ();
 sg13g2_fill_2 FILLER_47_157 ();
 sg13g2_fill_1 FILLER_47_159 ();
 sg13g2_decap_4 FILLER_47_190 ();
 sg13g2_decap_4 FILLER_47_217 ();
 sg13g2_decap_4 FILLER_47_226 ();
 sg13g2_fill_2 FILLER_47_230 ();
 sg13g2_fill_1 FILLER_47_236 ();
 sg13g2_fill_1 FILLER_47_259 ();
 sg13g2_fill_2 FILLER_47_298 ();
 sg13g2_fill_1 FILLER_47_300 ();
 sg13g2_decap_8 FILLER_47_313 ();
 sg13g2_fill_1 FILLER_47_320 ();
 sg13g2_fill_2 FILLER_47_358 ();
 sg13g2_fill_1 FILLER_47_360 ();
 sg13g2_decap_8 FILLER_47_373 ();
 sg13g2_decap_8 FILLER_47_380 ();
 sg13g2_decap_8 FILLER_47_387 ();
 sg13g2_decap_8 FILLER_47_394 ();
 sg13g2_decap_8 FILLER_47_401 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_4 FILLER_48_147 ();
 sg13g2_fill_2 FILLER_48_151 ();
 sg13g2_decap_4 FILLER_48_162 ();
 sg13g2_fill_1 FILLER_48_180 ();
 sg13g2_fill_2 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_48_202 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_fill_2 FILLER_48_273 ();
 sg13g2_fill_1 FILLER_48_275 ();
 sg13g2_fill_1 FILLER_48_329 ();
 sg13g2_decap_4 FILLER_48_334 ();
 sg13g2_decap_8 FILLER_48_387 ();
 sg13g2_decap_8 FILLER_48_394 ();
 sg13g2_decap_8 FILLER_48_401 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_4 FILLER_49_140 ();
 sg13g2_fill_1 FILLER_49_144 ();
 sg13g2_fill_1 FILLER_49_171 ();
 sg13g2_fill_2 FILLER_49_177 ();
 sg13g2_fill_1 FILLER_49_179 ();
 sg13g2_fill_2 FILLER_49_184 ();
 sg13g2_decap_8 FILLER_49_263 ();
 sg13g2_fill_1 FILLER_49_283 ();
 sg13g2_decap_8 FILLER_49_292 ();
 sg13g2_fill_1 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_391 ();
 sg13g2_decap_8 FILLER_49_398 ();
 sg13g2_decap_4 FILLER_49_405 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_4 FILLER_50_147 ();
 sg13g2_fill_2 FILLER_50_203 ();
 sg13g2_fill_1 FILLER_50_205 ();
 sg13g2_decap_4 FILLER_50_246 ();
 sg13g2_fill_1 FILLER_50_250 ();
 sg13g2_decap_4 FILLER_50_260 ();
 sg13g2_decap_8 FILLER_50_269 ();
 sg13g2_fill_2 FILLER_50_276 ();
 sg13g2_fill_1 FILLER_50_278 ();
 sg13g2_decap_8 FILLER_50_288 ();
 sg13g2_fill_2 FILLER_50_295 ();
 sg13g2_decap_4 FILLER_50_303 ();
 sg13g2_decap_4 FILLER_50_312 ();
 sg13g2_fill_1 FILLER_50_336 ();
 sg13g2_decap_8 FILLER_50_393 ();
 sg13g2_decap_8 FILLER_50_400 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_fill_1 FILLER_51_166 ();
 sg13g2_decap_8 FILLER_51_200 ();
 sg13g2_decap_4 FILLER_51_207 ();
 sg13g2_fill_2 FILLER_51_211 ();
 sg13g2_fill_1 FILLER_51_254 ();
 sg13g2_decap_8 FILLER_51_271 ();
 sg13g2_decap_4 FILLER_51_278 ();
 sg13g2_fill_1 FILLER_51_282 ();
 sg13g2_fill_2 FILLER_51_304 ();
 sg13g2_fill_1 FILLER_51_306 ();
 sg13g2_fill_2 FILLER_51_337 ();
 sg13g2_fill_1 FILLER_51_362 ();
 sg13g2_decap_8 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_decap_4 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_4 FILLER_52_91 ();
 sg13g2_fill_2 FILLER_52_95 ();
 sg13g2_decap_8 FILLER_52_101 ();
 sg13g2_decap_4 FILLER_52_108 ();
 sg13g2_decap_8 FILLER_52_116 ();
 sg13g2_decap_8 FILLER_52_123 ();
 sg13g2_decap_8 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_173 ();
 sg13g2_fill_1 FILLER_52_198 ();
 sg13g2_fill_1 FILLER_52_203 ();
 sg13g2_decap_8 FILLER_52_208 ();
 sg13g2_fill_2 FILLER_52_215 ();
 sg13g2_fill_1 FILLER_52_217 ();
 sg13g2_fill_1 FILLER_52_224 ();
 sg13g2_decap_4 FILLER_52_235 ();
 sg13g2_fill_1 FILLER_52_239 ();
 sg13g2_fill_2 FILLER_52_251 ();
 sg13g2_decap_8 FILLER_52_277 ();
 sg13g2_fill_1 FILLER_52_284 ();
 sg13g2_fill_1 FILLER_52_311 ();
 sg13g2_fill_2 FILLER_52_321 ();
 sg13g2_fill_1 FILLER_52_323 ();
 sg13g2_decap_8 FILLER_52_387 ();
 sg13g2_decap_8 FILLER_52_394 ();
 sg13g2_decap_8 FILLER_52_401 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_fill_2 FILLER_53_84 ();
 sg13g2_fill_1 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_122 ();
 sg13g2_decap_8 FILLER_53_129 ();
 sg13g2_decap_4 FILLER_53_136 ();
 sg13g2_fill_2 FILLER_53_140 ();
 sg13g2_fill_1 FILLER_53_192 ();
 sg13g2_fill_2 FILLER_53_219 ();
 sg13g2_fill_2 FILLER_53_236 ();
 sg13g2_decap_4 FILLER_53_242 ();
 sg13g2_fill_2 FILLER_53_252 ();
 sg13g2_fill_1 FILLER_53_254 ();
 sg13g2_fill_2 FILLER_53_266 ();
 sg13g2_fill_2 FILLER_53_304 ();
 sg13g2_fill_2 FILLER_53_315 ();
 sg13g2_fill_2 FILLER_53_341 ();
 sg13g2_decap_8 FILLER_53_382 ();
 sg13g2_decap_8 FILLER_53_389 ();
 sg13g2_decap_8 FILLER_53_396 ();
 sg13g2_decap_4 FILLER_53_403 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_4 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_130 ();
 sg13g2_decap_8 FILLER_54_137 ();
 sg13g2_fill_2 FILLER_54_144 ();
 sg13g2_fill_2 FILLER_54_184 ();
 sg13g2_fill_1 FILLER_54_195 ();
 sg13g2_decap_4 FILLER_54_239 ();
 sg13g2_fill_1 FILLER_54_243 ();
 sg13g2_fill_2 FILLER_54_249 ();
 sg13g2_fill_1 FILLER_54_303 ();
 sg13g2_fill_2 FILLER_54_309 ();
 sg13g2_fill_1 FILLER_54_311 ();
 sg13g2_fill_2 FILLER_54_317 ();
 sg13g2_fill_1 FILLER_54_319 ();
 sg13g2_fill_2 FILLER_54_325 ();
 sg13g2_decap_8 FILLER_54_393 ();
 sg13g2_decap_8 FILLER_54_400 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_fill_1 FILLER_55_77 ();
 sg13g2_fill_2 FILLER_55_95 ();
 sg13g2_fill_2 FILLER_55_113 ();
 sg13g2_decap_4 FILLER_55_119 ();
 sg13g2_fill_2 FILLER_55_123 ();
 sg13g2_decap_4 FILLER_55_130 ();
 sg13g2_fill_2 FILLER_55_134 ();
 sg13g2_fill_2 FILLER_55_191 ();
 sg13g2_fill_2 FILLER_55_267 ();
 sg13g2_fill_1 FILLER_55_269 ();
 sg13g2_decap_4 FILLER_55_294 ();
 sg13g2_fill_1 FILLER_55_337 ();
 sg13g2_decap_8 FILLER_55_386 ();
 sg13g2_decap_8 FILLER_55_393 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_fill_1 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_111 ();
 sg13g2_decap_8 FILLER_56_118 ();
 sg13g2_decap_8 FILLER_56_125 ();
 sg13g2_decap_8 FILLER_56_132 ();
 sg13g2_fill_2 FILLER_56_139 ();
 sg13g2_fill_2 FILLER_56_171 ();
 sg13g2_fill_1 FILLER_56_173 ();
 sg13g2_fill_2 FILLER_56_191 ();
 sg13g2_fill_1 FILLER_56_193 ();
 sg13g2_fill_1 FILLER_56_208 ();
 sg13g2_decap_4 FILLER_56_280 ();
 sg13g2_fill_2 FILLER_56_284 ();
 sg13g2_decap_4 FILLER_56_291 ();
 sg13g2_fill_2 FILLER_56_310 ();
 sg13g2_fill_2 FILLER_56_322 ();
 sg13g2_fill_1 FILLER_56_348 ();
 sg13g2_fill_1 FILLER_56_358 ();
 sg13g2_decap_8 FILLER_56_393 ();
 sg13g2_decap_8 FILLER_56_400 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_fill_2 FILLER_57_110 ();
 sg13g2_fill_1 FILLER_57_112 ();
 sg13g2_decap_4 FILLER_57_117 ();
 sg13g2_decap_8 FILLER_57_130 ();
 sg13g2_decap_4 FILLER_57_137 ();
 sg13g2_fill_1 FILLER_57_141 ();
 sg13g2_fill_2 FILLER_57_150 ();
 sg13g2_decap_4 FILLER_57_160 ();
 sg13g2_fill_1 FILLER_57_196 ();
 sg13g2_fill_1 FILLER_57_211 ();
 sg13g2_fill_1 FILLER_57_236 ();
 sg13g2_fill_2 FILLER_57_251 ();
 sg13g2_fill_1 FILLER_57_253 ();
 sg13g2_fill_2 FILLER_57_260 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_decap_8 FILLER_57_278 ();
 sg13g2_decap_8 FILLER_57_285 ();
 sg13g2_fill_2 FILLER_57_292 ();
 sg13g2_fill_1 FILLER_57_300 ();
 sg13g2_decap_4 FILLER_57_310 ();
 sg13g2_fill_2 FILLER_57_323 ();
 sg13g2_fill_1 FILLER_57_325 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_8 FILLER_57_400 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_fill_2 FILLER_58_99 ();
 sg13g2_fill_1 FILLER_58_106 ();
 sg13g2_decap_8 FILLER_58_141 ();
 sg13g2_decap_8 FILLER_58_148 ();
 sg13g2_fill_2 FILLER_58_168 ();
 sg13g2_fill_1 FILLER_58_222 ();
 sg13g2_decap_8 FILLER_58_240 ();
 sg13g2_decap_4 FILLER_58_255 ();
 sg13g2_fill_2 FILLER_58_263 ();
 sg13g2_fill_1 FILLER_58_265 ();
 sg13g2_fill_1 FILLER_58_271 ();
 sg13g2_fill_1 FILLER_58_277 ();
 sg13g2_decap_4 FILLER_58_283 ();
 sg13g2_fill_2 FILLER_58_310 ();
 sg13g2_fill_1 FILLER_58_312 ();
 sg13g2_decap_4 FILLER_58_319 ();
 sg13g2_fill_2 FILLER_58_327 ();
 sg13g2_fill_1 FILLER_58_341 ();
 sg13g2_decap_8 FILLER_58_393 ();
 sg13g2_decap_8 FILLER_58_400 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_4 FILLER_59_56 ();
 sg13g2_fill_2 FILLER_59_137 ();
 sg13g2_fill_1 FILLER_59_139 ();
 sg13g2_fill_2 FILLER_59_172 ();
 sg13g2_fill_1 FILLER_59_174 ();
 sg13g2_fill_2 FILLER_59_198 ();
 sg13g2_fill_1 FILLER_59_200 ();
 sg13g2_fill_2 FILLER_59_211 ();
 sg13g2_decap_8 FILLER_59_227 ();
 sg13g2_decap_4 FILLER_59_234 ();
 sg13g2_fill_1 FILLER_59_238 ();
 sg13g2_fill_1 FILLER_59_251 ();
 sg13g2_fill_2 FILLER_59_256 ();
 sg13g2_decap_4 FILLER_59_266 ();
 sg13g2_fill_2 FILLER_59_270 ();
 sg13g2_decap_4 FILLER_59_286 ();
 sg13g2_fill_1 FILLER_59_297 ();
 sg13g2_fill_2 FILLER_59_325 ();
 sg13g2_fill_1 FILLER_59_332 ();
 sg13g2_decap_8 FILLER_59_375 ();
 sg13g2_decap_8 FILLER_59_382 ();
 sg13g2_decap_8 FILLER_59_389 ();
 sg13g2_decap_8 FILLER_59_396 ();
 sg13g2_decap_4 FILLER_59_403 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_fill_2 FILLER_60_63 ();
 sg13g2_fill_1 FILLER_60_91 ();
 sg13g2_fill_1 FILLER_60_102 ();
 sg13g2_fill_2 FILLER_60_165 ();
 sg13g2_fill_2 FILLER_60_176 ();
 sg13g2_fill_2 FILLER_60_193 ();
 sg13g2_fill_1 FILLER_60_195 ();
 sg13g2_fill_1 FILLER_60_206 ();
 sg13g2_decap_8 FILLER_60_215 ();
 sg13g2_decap_4 FILLER_60_222 ();
 sg13g2_fill_2 FILLER_60_226 ();
 sg13g2_fill_2 FILLER_60_281 ();
 sg13g2_fill_1 FILLER_60_283 ();
 sg13g2_fill_1 FILLER_60_317 ();
 sg13g2_fill_2 FILLER_60_349 ();
 sg13g2_fill_1 FILLER_60_351 ();
 sg13g2_decap_8 FILLER_60_369 ();
 sg13g2_decap_8 FILLER_60_376 ();
 sg13g2_decap_8 FILLER_60_383 ();
 sg13g2_decap_8 FILLER_60_390 ();
 sg13g2_decap_8 FILLER_60_397 ();
 sg13g2_decap_4 FILLER_60_404 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_fill_2 FILLER_61_63 ();
 sg13g2_fill_2 FILLER_61_96 ();
 sg13g2_fill_1 FILLER_61_106 ();
 sg13g2_fill_1 FILLER_61_117 ();
 sg13g2_decap_8 FILLER_61_136 ();
 sg13g2_fill_1 FILLER_61_143 ();
 sg13g2_fill_2 FILLER_61_210 ();
 sg13g2_fill_1 FILLER_61_212 ();
 sg13g2_fill_2 FILLER_61_223 ();
 sg13g2_fill_1 FILLER_61_225 ();
 sg13g2_fill_2 FILLER_61_238 ();
 sg13g2_fill_1 FILLER_61_240 ();
 sg13g2_fill_2 FILLER_61_250 ();
 sg13g2_fill_1 FILLER_61_252 ();
 sg13g2_fill_1 FILLER_61_270 ();
 sg13g2_fill_1 FILLER_61_284 ();
 sg13g2_fill_2 FILLER_61_296 ();
 sg13g2_fill_2 FILLER_61_303 ();
 sg13g2_fill_1 FILLER_61_327 ();
 sg13g2_decap_8 FILLER_61_363 ();
 sg13g2_decap_8 FILLER_61_370 ();
 sg13g2_decap_8 FILLER_61_377 ();
 sg13g2_decap_8 FILLER_61_384 ();
 sg13g2_decap_8 FILLER_61_391 ();
 sg13g2_decap_8 FILLER_61_398 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_4 FILLER_62_70 ();
 sg13g2_fill_1 FILLER_62_74 ();
 sg13g2_fill_2 FILLER_62_86 ();
 sg13g2_decap_8 FILLER_62_129 ();
 sg13g2_fill_2 FILLER_62_136 ();
 sg13g2_fill_1 FILLER_62_164 ();
 sg13g2_fill_2 FILLER_62_190 ();
 sg13g2_fill_1 FILLER_62_202 ();
 sg13g2_fill_2 FILLER_62_247 ();
 sg13g2_fill_1 FILLER_62_249 ();
 sg13g2_fill_2 FILLER_62_256 ();
 sg13g2_decap_8 FILLER_62_292 ();
 sg13g2_decap_4 FILLER_62_299 ();
 sg13g2_fill_2 FILLER_62_303 ();
 sg13g2_fill_1 FILLER_62_310 ();
 sg13g2_fill_2 FILLER_62_332 ();
 sg13g2_fill_1 FILLER_62_334 ();
 sg13g2_fill_2 FILLER_62_344 ();
 sg13g2_decap_8 FILLER_62_380 ();
 sg13g2_decap_8 FILLER_62_387 ();
 sg13g2_decap_8 FILLER_62_394 ();
 sg13g2_decap_8 FILLER_62_401 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_4 FILLER_63_63 ();
 sg13g2_fill_2 FILLER_63_67 ();
 sg13g2_fill_2 FILLER_63_119 ();
 sg13g2_fill_1 FILLER_63_121 ();
 sg13g2_fill_1 FILLER_63_137 ();
 sg13g2_fill_2 FILLER_63_146 ();
 sg13g2_fill_1 FILLER_63_148 ();
 sg13g2_fill_1 FILLER_63_153 ();
 sg13g2_fill_2 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_182 ();
 sg13g2_fill_2 FILLER_63_207 ();
 sg13g2_fill_1 FILLER_63_209 ();
 sg13g2_fill_2 FILLER_63_229 ();
 sg13g2_fill_1 FILLER_63_231 ();
 sg13g2_fill_1 FILLER_63_252 ();
 sg13g2_fill_2 FILLER_63_266 ();
 sg13g2_fill_1 FILLER_63_274 ();
 sg13g2_fill_1 FILLER_63_283 ();
 sg13g2_fill_2 FILLER_63_326 ();
 sg13g2_fill_1 FILLER_63_328 ();
 sg13g2_fill_2 FILLER_63_340 ();
 sg13g2_decap_8 FILLER_63_377 ();
 sg13g2_decap_8 FILLER_63_384 ();
 sg13g2_decap_8 FILLER_63_391 ();
 sg13g2_decap_8 FILLER_63_398 ();
 sg13g2_decap_4 FILLER_63_405 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_4 FILLER_64_56 ();
 sg13g2_fill_2 FILLER_64_60 ();
 sg13g2_fill_2 FILLER_64_135 ();
 sg13g2_fill_1 FILLER_64_163 ();
 sg13g2_fill_2 FILLER_64_179 ();
 sg13g2_fill_2 FILLER_64_195 ();
 sg13g2_fill_2 FILLER_64_224 ();
 sg13g2_fill_1 FILLER_64_226 ();
 sg13g2_fill_2 FILLER_64_272 ();
 sg13g2_decap_8 FILLER_64_299 ();
 sg13g2_decap_8 FILLER_64_374 ();
 sg13g2_decap_8 FILLER_64_381 ();
 sg13g2_decap_8 FILLER_64_388 ();
 sg13g2_decap_8 FILLER_64_395 ();
 sg13g2_decap_8 FILLER_64_402 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_fill_2 FILLER_65_134 ();
 sg13g2_fill_2 FILLER_65_162 ();
 sg13g2_fill_1 FILLER_65_164 ();
 sg13g2_decap_8 FILLER_65_205 ();
 sg13g2_decap_4 FILLER_65_212 ();
 sg13g2_fill_1 FILLER_65_216 ();
 sg13g2_decap_8 FILLER_65_225 ();
 sg13g2_fill_2 FILLER_65_232 ();
 sg13g2_fill_1 FILLER_65_234 ();
 sg13g2_fill_2 FILLER_65_291 ();
 sg13g2_fill_1 FILLER_65_293 ();
 sg13g2_fill_2 FILLER_65_299 ();
 sg13g2_fill_1 FILLER_65_301 ();
 sg13g2_fill_2 FILLER_65_315 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_fill_1 FILLER_66_63 ();
 sg13g2_fill_1 FILLER_66_82 ();
 sg13g2_fill_2 FILLER_66_99 ();
 sg13g2_fill_1 FILLER_66_101 ();
 sg13g2_fill_2 FILLER_66_111 ();
 sg13g2_decap_8 FILLER_66_132 ();
 sg13g2_fill_2 FILLER_66_139 ();
 sg13g2_fill_1 FILLER_66_141 ();
 sg13g2_fill_1 FILLER_66_146 ();
 sg13g2_fill_2 FILLER_66_169 ();
 sg13g2_fill_1 FILLER_66_171 ();
 sg13g2_fill_2 FILLER_66_186 ();
 sg13g2_fill_1 FILLER_66_207 ();
 sg13g2_fill_2 FILLER_66_218 ();
 sg13g2_fill_1 FILLER_66_220 ();
 sg13g2_fill_1 FILLER_66_227 ();
 sg13g2_decap_8 FILLER_66_254 ();
 sg13g2_decap_4 FILLER_66_261 ();
 sg13g2_fill_1 FILLER_66_265 ();
 sg13g2_decap_8 FILLER_66_270 ();
 sg13g2_fill_2 FILLER_66_277 ();
 sg13g2_fill_2 FILLER_66_295 ();
 sg13g2_fill_1 FILLER_66_297 ();
 sg13g2_fill_2 FILLER_66_306 ();
 sg13g2_fill_1 FILLER_66_308 ();
 sg13g2_fill_2 FILLER_66_317 ();
 sg13g2_decap_8 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_371 ();
 sg13g2_decap_8 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_385 ();
 sg13g2_decap_8 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_66_399 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_4 FILLER_67_140 ();
 sg13g2_fill_1 FILLER_67_144 ();
 sg13g2_decap_4 FILLER_67_171 ();
 sg13g2_fill_1 FILLER_67_175 ();
 sg13g2_fill_2 FILLER_67_192 ();
 sg13g2_fill_1 FILLER_67_240 ();
 sg13g2_fill_2 FILLER_67_254 ();
 sg13g2_fill_1 FILLER_67_256 ();
 sg13g2_fill_2 FILLER_67_272 ();
 sg13g2_fill_1 FILLER_67_274 ();
 sg13g2_fill_1 FILLER_67_311 ();
 sg13g2_fill_2 FILLER_67_360 ();
 sg13g2_fill_1 FILLER_67_362 ();
 sg13g2_decap_8 FILLER_67_389 ();
 sg13g2_decap_8 FILLER_67_396 ();
 sg13g2_decap_4 FILLER_67_403 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_fill_1 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_118 ();
 sg13g2_decap_8 FILLER_68_125 ();
 sg13g2_decap_8 FILLER_68_132 ();
 sg13g2_decap_8 FILLER_68_139 ();
 sg13g2_fill_1 FILLER_68_146 ();
 sg13g2_fill_2 FILLER_68_161 ();
 sg13g2_fill_1 FILLER_68_163 ();
 sg13g2_fill_1 FILLER_68_184 ();
 sg13g2_fill_2 FILLER_68_201 ();
 sg13g2_fill_1 FILLER_68_203 ();
 sg13g2_fill_2 FILLER_68_218 ();
 sg13g2_fill_1 FILLER_68_220 ();
 sg13g2_fill_1 FILLER_68_227 ();
 sg13g2_decap_8 FILLER_68_276 ();
 sg13g2_decap_4 FILLER_68_283 ();
 sg13g2_fill_2 FILLER_68_287 ();
 sg13g2_decap_4 FILLER_68_293 ();
 sg13g2_fill_1 FILLER_68_297 ();
 sg13g2_fill_2 FILLER_68_321 ();
 sg13g2_fill_1 FILLER_68_323 ();
 sg13g2_fill_2 FILLER_68_351 ();
 sg13g2_decap_8 FILLER_68_392 ();
 sg13g2_decap_8 FILLER_68_399 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_4 FILLER_69_84 ();
 sg13g2_fill_1 FILLER_69_88 ();
 sg13g2_decap_8 FILLER_69_93 ();
 sg13g2_decap_8 FILLER_69_122 ();
 sg13g2_decap_4 FILLER_69_129 ();
 sg13g2_fill_1 FILLER_69_164 ();
 sg13g2_fill_2 FILLER_69_189 ();
 sg13g2_fill_1 FILLER_69_191 ();
 sg13g2_fill_1 FILLER_69_207 ();
 sg13g2_fill_2 FILLER_69_217 ();
 sg13g2_decap_4 FILLER_69_228 ();
 sg13g2_decap_8 FILLER_69_244 ();
 sg13g2_fill_1 FILLER_69_251 ();
 sg13g2_decap_8 FILLER_69_261 ();
 sg13g2_fill_2 FILLER_69_268 ();
 sg13g2_decap_8 FILLER_69_284 ();
 sg13g2_fill_1 FILLER_69_324 ();
 sg13g2_fill_2 FILLER_69_347 ();
 sg13g2_fill_2 FILLER_69_367 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_fill_2 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_fill_2 FILLER_70_77 ();
 sg13g2_fill_1 FILLER_70_79 ();
 sg13g2_fill_2 FILLER_70_191 ();
 sg13g2_fill_2 FILLER_70_210 ();
 sg13g2_decap_8 FILLER_70_223 ();
 sg13g2_fill_2 FILLER_70_230 ();
 sg13g2_fill_1 FILLER_70_232 ();
 sg13g2_fill_1 FILLER_70_275 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_fill_2 FILLER_70_307 ();
 sg13g2_fill_2 FILLER_70_376 ();
 sg13g2_fill_1 FILLER_70_378 ();
 sg13g2_fill_2 FILLER_70_406 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_fill_1 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_101 ();
 sg13g2_decap_8 FILLER_71_108 ();
 sg13g2_decap_8 FILLER_71_115 ();
 sg13g2_decap_8 FILLER_71_122 ();
 sg13g2_fill_1 FILLER_71_129 ();
 sg13g2_decap_8 FILLER_71_134 ();
 sg13g2_decap_8 FILLER_71_141 ();
 sg13g2_fill_2 FILLER_71_165 ();
 sg13g2_fill_1 FILLER_71_177 ();
 sg13g2_fill_1 FILLER_71_184 ();
 sg13g2_fill_2 FILLER_71_204 ();
 sg13g2_fill_2 FILLER_71_211 ();
 sg13g2_fill_1 FILLER_71_213 ();
 sg13g2_fill_1 FILLER_71_241 ();
 sg13g2_fill_1 FILLER_71_311 ();
 sg13g2_fill_2 FILLER_71_339 ();
 sg13g2_decap_8 FILLER_71_400 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_fill_1 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_110 ();
 sg13g2_decap_8 FILLER_72_117 ();
 sg13g2_decap_8 FILLER_72_124 ();
 sg13g2_decap_8 FILLER_72_131 ();
 sg13g2_decap_4 FILLER_72_138 ();
 sg13g2_fill_2 FILLER_72_142 ();
 sg13g2_fill_2 FILLER_72_170 ();
 sg13g2_fill_2 FILLER_72_191 ();
 sg13g2_fill_1 FILLER_72_193 ();
 sg13g2_fill_1 FILLER_72_257 ();
 sg13g2_fill_2 FILLER_72_277 ();
 sg13g2_fill_1 FILLER_72_284 ();
 sg13g2_fill_2 FILLER_72_367 ();
 sg13g2_fill_1 FILLER_72_384 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_fill_2 FILLER_73_96 ();
 sg13g2_fill_2 FILLER_73_112 ();
 sg13g2_fill_1 FILLER_73_114 ();
 sg13g2_fill_1 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_124 ();
 sg13g2_decap_8 FILLER_73_131 ();
 sg13g2_decap_8 FILLER_73_138 ();
 sg13g2_fill_2 FILLER_73_145 ();
 sg13g2_fill_2 FILLER_73_206 ();
 sg13g2_fill_1 FILLER_73_208 ();
 sg13g2_fill_2 FILLER_73_260 ();
 sg13g2_fill_1 FILLER_73_262 ();
 sg13g2_fill_2 FILLER_73_268 ();
 sg13g2_fill_1 FILLER_73_270 ();
 sg13g2_fill_2 FILLER_73_291 ();
 sg13g2_fill_1 FILLER_73_293 ();
 sg13g2_fill_2 FILLER_73_315 ();
 sg13g2_fill_1 FILLER_73_317 ();
 sg13g2_fill_1 FILLER_73_329 ();
 sg13g2_fill_1 FILLER_73_348 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_fill_2 FILLER_74_70 ();
 sg13g2_fill_1 FILLER_74_72 ();
 sg13g2_fill_2 FILLER_74_106 ();
 sg13g2_fill_1 FILLER_74_108 ();
 sg13g2_decap_8 FILLER_74_135 ();
 sg13g2_decap_8 FILLER_74_142 ();
 sg13g2_fill_2 FILLER_74_149 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_fill_2 FILLER_74_237 ();
 sg13g2_fill_2 FILLER_74_260 ();
 sg13g2_fill_1 FILLER_74_262 ();
 sg13g2_fill_2 FILLER_74_318 ();
 sg13g2_fill_1 FILLER_74_320 ();
 sg13g2_fill_1 FILLER_74_341 ();
 sg13g2_fill_2 FILLER_74_347 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_4 FILLER_75_70 ();
 sg13g2_fill_2 FILLER_75_74 ();
 sg13g2_fill_2 FILLER_75_102 ();
 sg13g2_fill_1 FILLER_75_109 ();
 sg13g2_decap_8 FILLER_75_148 ();
 sg13g2_fill_2 FILLER_75_185 ();
 sg13g2_decap_4 FILLER_75_200 ();
 sg13g2_fill_2 FILLER_75_204 ();
 sg13g2_fill_1 FILLER_75_210 ();
 sg13g2_fill_2 FILLER_75_225 ();
 sg13g2_fill_1 FILLER_75_240 ();
 sg13g2_fill_1 FILLER_75_285 ();
 sg13g2_fill_2 FILLER_75_295 ();
 sg13g2_fill_1 FILLER_75_297 ();
 sg13g2_fill_2 FILLER_75_321 ();
 sg13g2_fill_1 FILLER_75_323 ();
 sg13g2_fill_2 FILLER_75_381 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_4 FILLER_76_70 ();
 sg13g2_fill_1 FILLER_76_74 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_fill_2 FILLER_76_187 ();
 sg13g2_fill_1 FILLER_76_189 ();
 sg13g2_fill_2 FILLER_76_203 ();
 sg13g2_fill_1 FILLER_76_213 ();
 sg13g2_fill_2 FILLER_76_253 ();
 sg13g2_fill_2 FILLER_76_261 ();
 sg13g2_fill_1 FILLER_76_295 ();
 sg13g2_decap_8 FILLER_76_393 ();
 sg13g2_decap_8 FILLER_76_400 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_fill_2 FILLER_77_70 ();
 sg13g2_fill_1 FILLER_77_72 ();
 sg13g2_fill_2 FILLER_77_95 ();
 sg13g2_fill_1 FILLER_77_106 ();
 sg13g2_decap_8 FILLER_77_139 ();
 sg13g2_decap_8 FILLER_77_146 ();
 sg13g2_decap_8 FILLER_77_153 ();
 sg13g2_decap_8 FILLER_77_160 ();
 sg13g2_fill_1 FILLER_77_167 ();
 sg13g2_decap_4 FILLER_77_194 ();
 sg13g2_fill_1 FILLER_77_198 ();
 sg13g2_fill_2 FILLER_77_237 ();
 sg13g2_fill_1 FILLER_77_362 ();
 sg13g2_fill_2 FILLER_77_374 ();
 sg13g2_decap_4 FILLER_77_403 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_137 ();
 sg13g2_decap_8 FILLER_78_144 ();
 sg13g2_decap_8 FILLER_78_151 ();
 sg13g2_decap_4 FILLER_78_158 ();
 sg13g2_fill_2 FILLER_78_162 ();
 sg13g2_fill_2 FILLER_78_273 ();
 sg13g2_fill_1 FILLER_78_275 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_4 FILLER_78_403 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_fill_2 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_136 ();
 sg13g2_decap_8 FILLER_79_143 ();
 sg13g2_decap_8 FILLER_79_150 ();
 sg13g2_decap_8 FILLER_79_157 ();
 sg13g2_decap_8 FILLER_79_164 ();
 sg13g2_fill_2 FILLER_79_171 ();
 sg13g2_fill_1 FILLER_79_173 ();
 sg13g2_decap_4 FILLER_79_200 ();
 sg13g2_fill_2 FILLER_79_208 ();
 sg13g2_decap_8 FILLER_79_214 ();
 sg13g2_fill_2 FILLER_79_221 ();
 sg13g2_fill_2 FILLER_79_249 ();
 sg13g2_fill_1 FILLER_79_277 ();
 sg13g2_fill_2 FILLER_79_287 ();
 sg13g2_fill_2 FILLER_79_301 ();
 sg13g2_fill_2 FILLER_79_307 ();
 sg13g2_fill_2 FILLER_79_313 ();
 sg13g2_fill_1 FILLER_79_315 ();
 sg13g2_fill_2 FILLER_79_346 ();
 sg13g2_fill_1 FILLER_79_348 ();
 sg13g2_decap_8 FILLER_79_393 ();
 sg13g2_decap_8 FILLER_79_400 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_fill_1 FILLER_80_92 ();
 sg13g2_fill_1 FILLER_80_105 ();
 sg13g2_fill_1 FILLER_80_115 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_fill_2 FILLER_80_172 ();
 sg13g2_fill_2 FILLER_80_182 ();
 sg13g2_decap_4 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_204 ();
 sg13g2_decap_4 FILLER_80_212 ();
 sg13g2_decap_4 FILLER_80_220 ();
 sg13g2_fill_1 FILLER_80_224 ();
 sg13g2_decap_4 FILLER_80_245 ();
 sg13g2_fill_2 FILLER_80_249 ();
 sg13g2_fill_2 FILLER_80_259 ();
 sg13g2_fill_2 FILLER_80_265 ();
 sg13g2_fill_1 FILLER_80_267 ();
 sg13g2_fill_2 FILLER_80_272 ();
 sg13g2_decap_4 FILLER_80_298 ();
 sg13g2_fill_2 FILLER_80_302 ();
 sg13g2_decap_8 FILLER_80_308 ();
 sg13g2_decap_4 FILLER_80_315 ();
 sg13g2_fill_1 FILLER_80_323 ();
 sg13g2_decap_4 FILLER_80_337 ();
 sg13g2_fill_1 FILLER_80_341 ();
 sg13g2_fill_2 FILLER_80_346 ();
 sg13g2_fill_1 FILLER_80_348 ();
 sg13g2_fill_1 FILLER_80_353 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[2] = net18;
 assign uo_out[3] = net19;
 assign uo_out[4] = net20;
 assign uo_out[5] = net21;
 assign uo_out[6] = net22;
 assign uo_out[7] = net23;
endmodule

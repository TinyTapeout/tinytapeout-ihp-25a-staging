module tt_um_wokwi_group_10 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire \proj_10.net10 ;
 wire \proj_10.net11 ;
 wire \proj_10.net12 ;
 wire \proj_12.net10 ;
 wire \proj_12.net15 ;
 wire \proj_12.net16 ;
 wire \proj_12.net17 ;
 wire \proj_12.net18 ;
 wire \proj_12.net20 ;
 wire \proj_12.net3 ;
 wire \proj_12.net4 ;
 wire \proj_12.net5 ;
 wire \proj_12.net6 ;
 wire \proj_12.net7 ;
 wire \proj_12.net8 ;
 wire \proj_12.net9 ;
 wire \proj_13.net10 ;
 wire \proj_13.net11 ;
 wire \proj_13.net12 ;
 wire \proj_13.net18 ;
 wire \proj_13.net19 ;
 wire \proj_13.net9 ;
 wire \proj_14.net7 ;
 wire \proj__0.net12 ;
 wire \proj__0.net13 ;
 wire \proj__0.net14 ;
 wire \proj__0.net15 ;
 wire \proj__0.net16 ;
 wire \proj__0.net17 ;
 wire \proj__0.net18 ;
 wire \proj__0.net19 ;
 wire \proj__0.net20 ;
 wire \proj__0.net6 ;
 wire \proj__0.net7 ;
 wire \proj__1.net10 ;
 wire \proj__1.net11 ;
 wire \proj__1.net12 ;
 wire \proj__1.net13 ;
 wire \proj__1.net14 ;
 wire \proj__1.net15 ;
 wire \proj__1.net16 ;
 wire \proj__1.net17 ;
 wire \proj__1.net18 ;
 wire \proj__1.net19 ;
 wire \proj__1.net20 ;
 wire \proj__1.net21 ;
 wire \proj__1.net22 ;
 wire \proj__1.net23 ;
 wire \proj__1.net24 ;
 wire \proj__1.net25 ;
 wire \proj__1.net26 ;
 wire \proj__1.net27 ;
 wire \proj__1.net28 ;
 wire \proj__1.net29 ;
 wire \proj__1.net30 ;
 wire \proj__1.net31 ;
 wire \proj__1.net32 ;
 wire \proj__1.net6 ;
 wire \proj__1.net7 ;
 wire \proj__1.net8 ;
 wire \proj__2.net10 ;
 wire \proj__2.net11 ;
 wire \proj__2.net12 ;
 wire \proj__2.net9 ;
 wire \proj__3.net12 ;
 wire \proj__3.net13 ;
 wire \proj__3.net6 ;
 wire \proj__4.net10 ;
 wire \proj__4.net11 ;
 wire \proj__4.net12 ;
 wire \proj__4.net18 ;
 wire \proj__4.net9 ;
 wire \proj__5.net10 ;
 wire \proj__5.net11 ;
 wire \proj__5.net12 ;
 wire \proj__5.net13 ;
 wire \proj__5.net14 ;
 wire \proj__5.net9 ;
 wire \proj__6.net10 ;
 wire \proj__6.net11 ;
 wire \proj__6.net8 ;
 wire \proj__6.net9 ;
 wire \proj__7.net10 ;
 wire \proj__7.net9 ;
 wire \proj__8.net15 ;
 wire \proj__8.net16 ;
 wire \proj__8.net17 ;
 wire \proj__8.net18 ;
 wire \proj__8.net19 ;
 wire \proj__8.net2 ;
 wire \proj__8.net20 ;
 wire \proj__8.net21 ;
 wire \proj__8.net22 ;
 wire \proj__8.net23 ;
 wire \proj__8.net24 ;
 wire \proj__8.net25 ;
 wire \proj__8.net26 ;
 wire \proj__8.net27 ;
 wire \proj__8.net28 ;
 wire \proj__8.net29 ;
 wire \proj__8.net3 ;
 wire \proj__8.net30 ;
 wire \proj__8.net31 ;
 wire \proj__8.net32 ;
 wire \proj__8.net33 ;
 wire \proj__8.net34 ;
 wire \proj__8.net35 ;
 wire \proj__8.net36 ;
 wire \proj__8.net37 ;
 wire \proj__8.net38 ;
 wire \proj__8.net39 ;
 wire \proj__8.net4 ;
 wire \proj__8.net40 ;
 wire \proj__8.net41 ;
 wire \proj__8.net42 ;
 wire \proj__8.net43 ;
 wire \proj__8.net44 ;
 wire \proj__8.net45 ;
 wire \proj__8.net46 ;
 wire \proj__8.net47 ;
 wire \proj__8.net48 ;
 wire \proj__8.net5 ;
 wire \proj__8.net6 ;
 wire \proj__8.net7 ;
 wire \proj__8.net8 ;
 wire \proj__8.net9 ;
 wire \proj__9.net10 ;
 wire \proj__9.net11 ;
 wire \proj__9.net12 ;
 wire \proj__9.net4 ;
 wire \proj__9.net5 ;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire \proj_12.flop1/notq ;
 wire net50;
 wire \proj_12.flop2/notq ;
 wire net51;
 wire \proj_12.flop3/notq ;
 wire net52;
 wire \proj_12.flop4/notq ;
 wire net53;
 wire \proj_12.flop5/notq ;
 wire net54;
 wire \proj_12.flop6/notq ;
 wire net55;
 wire \proj_12.flop7/notq ;
 wire net56;
 wire \proj_12.flop8/notq ;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire \proj__8.flop1/notq ;
 wire net66;
 wire \proj__8.flop10/notq ;
 wire net67;
 wire \proj__8.flop11/notq ;
 wire net68;
 wire \proj__8.flop12/notq ;
 wire net69;
 wire \proj__8.flop13/notq ;
 wire net70;
 wire \proj__8.flop14/notq ;
 wire net71;
 wire \proj__8.flop15/notq ;
 wire net72;
 wire net73;
 wire \proj__8.flop17/notq ;
 wire net74;
 wire \proj__8.flop18/notq ;
 wire net75;
 wire \proj__8.flop19/notq ;
 wire net76;
 wire \proj__8.flop2/notq ;
 wire net77;
 wire \proj__8.flop20/notq ;
 wire net78;
 wire net79;
 wire \proj__8.flop3/notq ;
 wire net80;
 wire \proj__8.flop4/notq ;
 wire net81;
 wire \proj__8.flop5/notq ;
 wire net82;
 wire \proj__8.flop6/notq ;
 wire net83;
 wire \proj__8.flop7/notq ;
 wire net84;
 wire \proj__8.flop8/notq ;
 wire \proj__8.flop9/notq ;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;

 sg13g2_inv_1 _087_ (.Y(_044_),
    .A(net25));
 sg13g2_nor2_2 _088_ (.A(net6),
    .B(net7),
    .Y(_045_));
 sg13g2_nor2_2 _089_ (.A(net9),
    .B(net8),
    .Y(_046_));
 sg13g2_nand2_1 _090_ (.Y(_047_),
    .A(_045_),
    .B(_046_));
 sg13g2_nor2_1 _091_ (.A(\proj__0.net6 ),
    .B(_047_),
    .Y(_048_));
 sg13g2_nand2_1 _092_ (.Y(_049_),
    .A(net25),
    .B(net8));
 sg13g2_nor3_2 _093_ (.A(net6),
    .B(net7),
    .C(_049_),
    .Y(_050_));
 sg13g2_nor2b_2 _094_ (.A(net8),
    .B_N(net25),
    .Y(_051_));
 sg13g2_and2_2 _095_ (.A(_045_),
    .B(_051_),
    .X(_052_));
 sg13g2_nor2b_2 _096_ (.A(net7),
    .B_N(net6),
    .Y(_053_));
 sg13g2_nand3_1 _097_ (.B(_051_),
    .C(_053_),
    .A(\proj__9.net4 ),
    .Y(_054_));
 sg13g2_nor2b_2 _098_ (.A(_049_),
    .B_N(_053_),
    .Y(_055_));
 sg13g2_nand3_1 _099_ (.B(_046_),
    .C(_053_),
    .A(\proj__1.net6 ),
    .Y(_056_));
 sg13g2_nor2b_2 _100_ (.A(net25),
    .B_N(net8),
    .Y(_057_));
 sg13g2_nand2b_1 _101_ (.Y(_058_),
    .B(net8),
    .A_N(net25));
 sg13g2_nor2b_2 _102_ (.A(net6),
    .B_N(net7),
    .Y(_059_));
 sg13g2_and2_1 _103_ (.A(_057_),
    .B(_059_),
    .X(_060_));
 sg13g2_nand3_1 _104_ (.B(_057_),
    .C(_059_),
    .A(\proj__6.net8 ),
    .Y(_061_));
 sg13g2_and2_1 _105_ (.A(_046_),
    .B(_059_),
    .X(_062_));
 sg13g2_nand3_1 _106_ (.B(_046_),
    .C(_059_),
    .A(\proj__2.net9 ),
    .Y(_063_));
 sg13g2_nand2_1 _107_ (.Y(_064_),
    .A(net6),
    .B(net7));
 sg13g2_nor2_2 _108_ (.A(_058_),
    .B(_064_),
    .Y(_065_));
 sg13g2_and2_1 _109_ (.A(\proj__7.net9 ),
    .B(_065_),
    .X(_066_));
 sg13g2_and2_2 _110_ (.A(_053_),
    .B(_057_),
    .X(_067_));
 sg13g2_nand3_1 _111_ (.B(_053_),
    .C(_057_),
    .A(\proj__5.net9 ),
    .Y(_068_));
 sg13g2_nand4_1 _112_ (.B(net8),
    .C(\proj_14.net7 ),
    .A(net25),
    .Y(_069_),
    .D(_059_));
 sg13g2_and2_1 _113_ (.A(_051_),
    .B(_059_),
    .X(_070_));
 sg13g2_nand3_1 _114_ (.B(_051_),
    .C(_059_),
    .A(\proj_10.net10 ),
    .Y(_071_));
 sg13g2_nor3_1 _115_ (.A(net25),
    .B(net8),
    .C(_064_),
    .Y(_072_));
 sg13g2_and2_1 _116_ (.A(\proj__3.net6 ),
    .B(_072_),
    .X(_000_));
 sg13g2_nand4_1 _117_ (.B(_063_),
    .C(_068_),
    .A(_061_),
    .Y(_001_),
    .D(_069_));
 sg13g2_a22oi_1 _118_ (.Y(_002_),
    .B1(_052_),
    .B2(\proj__8.net2 ),
    .A2(_050_),
    .A1(\proj_12.net3 ));
 sg13g2_and2_2 _119_ (.A(_045_),
    .B(_057_),
    .X(_003_));
 sg13g2_a22oi_1 _120_ (.Y(_004_),
    .B1(_003_),
    .B2(\proj__4.net9 ),
    .A2(_055_),
    .A1(\proj_13.net9 ));
 sg13g2_and4_1 _121_ (.A(_047_),
    .B(_056_),
    .C(_002_),
    .D(_004_),
    .X(_005_));
 sg13g2_nand2_1 _122_ (.Y(_006_),
    .A(_054_),
    .B(_071_));
 sg13g2_nor4_1 _123_ (.A(_066_),
    .B(_000_),
    .C(_001_),
    .D(_006_),
    .Y(_007_));
 sg13g2_a21oi_2 _124_ (.B1(_048_),
    .Y(uo_out[0]),
    .A2(_007_),
    .A1(_005_));
 sg13g2_nor2_1 _125_ (.A(\proj__0.net7 ),
    .B(_047_),
    .Y(_008_));
 sg13g2_and3_1 _126_ (.X(_009_),
    .A(\proj__9.net5 ),
    .B(_051_),
    .C(_053_));
 sg13g2_and2_1 _127_ (.A(\proj_10.net11 ),
    .B(_070_),
    .X(_010_));
 sg13g2_and3_1 _128_ (.X(_011_),
    .A(\proj__1.net7 ),
    .B(_046_),
    .C(_053_));
 sg13g2_a221oi_1 _129_ (.B2(\proj__4.net10 ),
    .C1(_010_),
    .B1(_003_),
    .A1(net29),
    .Y(_012_),
    .A2(_072_));
 sg13g2_a22oi_1 _130_ (.Y(_013_),
    .B1(_067_),
    .B2(\proj__5.net10 ),
    .A2(_060_),
    .A1(\proj__6.net9 ));
 sg13g2_a22oi_1 _131_ (.Y(_014_),
    .B1(_052_),
    .B2(\proj__8.net3 ),
    .A2(_046_),
    .A1(_045_));
 sg13g2_a221oi_1 _132_ (.B2(\proj_13.net10 ),
    .C1(_009_),
    .B1(_055_),
    .A1(\proj_12.net4 ),
    .Y(_015_),
    .A2(_050_));
 sg13g2_a221oi_1 _133_ (.B2(\proj__7.net9 ),
    .C1(_011_),
    .B1(_065_),
    .A1(\proj__2.net10 ),
    .Y(_016_),
    .A2(_062_));
 sg13g2_and4_1 _134_ (.A(_013_),
    .B(_014_),
    .C(_015_),
    .D(_016_),
    .X(_017_));
 sg13g2_a21oi_2 _135_ (.B1(_008_),
    .Y(uo_out[1]),
    .A2(_017_),
    .A1(_012_));
 sg13g2_nor2_1 _136_ (.A(net25),
    .B(_064_),
    .Y(_018_));
 sg13g2_a22oi_1 _137_ (.Y(_019_),
    .B1(_070_),
    .B2(\proj_10.net12 ),
    .A2(_060_),
    .A1(\proj__6.net10 ));
 sg13g2_a22oi_1 _138_ (.Y(_020_),
    .B1(_067_),
    .B2(\proj__5.net11 ),
    .A2(_055_),
    .A1(\proj_13.net11 ));
 sg13g2_a22oi_1 _139_ (.Y(_021_),
    .B1(_018_),
    .B2(net26),
    .A2(_050_),
    .A1(\proj_12.net5 ));
 sg13g2_a22oi_1 _140_ (.Y(_022_),
    .B1(_003_),
    .B2(\proj__4.net11 ),
    .A2(_062_),
    .A1(\proj__2.net11 ));
 sg13g2_nand4_1 _141_ (.B(_020_),
    .C(_021_),
    .A(_019_),
    .Y(_023_),
    .D(_022_));
 sg13g2_a21o_1 _142_ (.A2(_052_),
    .A1(\proj__8.net4 ),
    .B1(_023_),
    .X(uo_out[2]));
 sg13g2_a21oi_1 _143_ (.A1(\proj_13.net11 ),
    .A2(_055_),
    .Y(_024_),
    .B1(_000_));
 sg13g2_o21ai_1 _144_ (.B1(net1),
    .Y(_025_),
    .A1(_065_),
    .A2(_070_));
 sg13g2_a22oi_1 _145_ (.Y(_026_),
    .B1(_060_),
    .B2(\proj__6.net11 ),
    .A2(_052_),
    .A1(\proj__8.net5 ));
 sg13g2_a22oi_1 _146_ (.Y(_027_),
    .B1(_003_),
    .B2(\proj__4.net12 ),
    .A2(_062_),
    .A1(\proj__2.net12 ));
 sg13g2_a22oi_1 _147_ (.Y(_028_),
    .B1(_067_),
    .B2(\proj__5.net12 ),
    .A2(_050_),
    .A1(\proj_12.net6 ));
 sg13g2_and3_1 _148_ (.X(_029_),
    .A(_025_),
    .B(_026_),
    .C(_028_));
 sg13g2_nand3_1 _149_ (.B(_027_),
    .C(_029_),
    .A(_024_),
    .Y(uo_out[3]));
 sg13g2_a22oi_1 _150_ (.Y(_030_),
    .B1(_058_),
    .B2(_059_),
    .A2(_045_),
    .A1(_044_));
 sg13g2_nand2b_1 _151_ (.Y(_031_),
    .B(_030_),
    .A_N(_065_));
 sg13g2_nand2b_1 _152_ (.Y(_032_),
    .B(_030_),
    .A_N(_067_));
 sg13g2_o21ai_1 _153_ (.B1(net2),
    .Y(_033_),
    .A1(_067_),
    .A2(_031_));
 sg13g2_a22oi_1 _154_ (.Y(_034_),
    .B1(_052_),
    .B2(\proj__8.net6 ),
    .A2(_050_),
    .A1(\proj_12.net7 ));
 sg13g2_nand3_1 _155_ (.B(_033_),
    .C(_034_),
    .A(_024_),
    .Y(uo_out[4]));
 sg13g2_nand2_1 _156_ (.Y(_035_),
    .A(\proj__5.net13 ),
    .B(_067_));
 sg13g2_a22oi_1 _157_ (.Y(_036_),
    .B1(_055_),
    .B2(\proj_13.net12 ),
    .A2(_052_),
    .A1(\proj__8.net7 ));
 sg13g2_a221oi_1 _158_ (.B2(net3),
    .C1(_000_),
    .B1(_031_),
    .A1(\proj_12.net8 ),
    .Y(_037_),
    .A2(_050_));
 sg13g2_nand3_1 _159_ (.B(_036_),
    .C(_037_),
    .A(_035_),
    .Y(uo_out[5]));
 sg13g2_nand2_1 _160_ (.Y(_038_),
    .A(\proj__7.net10 ),
    .B(_065_));
 sg13g2_a22oi_1 _161_ (.Y(_039_),
    .B1(_052_),
    .B2(\proj__8.net8 ),
    .A2(_050_),
    .A1(\proj_12.net9 ));
 sg13g2_a221oi_1 _162_ (.B2(net4),
    .C1(_000_),
    .B1(_032_),
    .A1(net5),
    .Y(_040_),
    .A2(_055_));
 sg13g2_nand3_1 _163_ (.B(_039_),
    .C(_040_),
    .A(_038_),
    .Y(uo_out[6]));
 sg13g2_nand2b_1 _164_ (.Y(_041_),
    .B(net5),
    .A_N(_030_));
 sg13g2_a22oi_1 _165_ (.Y(_042_),
    .B1(_067_),
    .B2(\proj__5.net14 ),
    .A2(_055_),
    .A1(net5));
 sg13g2_a22oi_1 _166_ (.Y(_043_),
    .B1(_052_),
    .B2(\proj__8.net9 ),
    .A2(_050_),
    .A1(\proj_12.net10 ));
 sg13g2_nand3_1 _167_ (.B(_042_),
    .C(_043_),
    .A(_041_),
    .Y(uo_out[7]));
 sg13g2_tielo \proj_12.flop1/_1__11  (.L_LO(net11));
 sg13g2_tielo \proj_12.flop2/_1__12  (.L_LO(net12));
 sg13g2_tielo \proj_12.flop3/_1__13  (.L_LO(net13));
 sg13g2_tielo \proj_12.flop4/_1__14  (.L_LO(net14));
 sg13g2_tielo \proj_12.flop5/_1__15  (.L_LO(net15));
 sg13g2_tielo \proj_12.flop6/_1__16  (.L_LO(net16));
 sg13g2_tielo \proj_12.flop7/_1__17  (.L_LO(net17));
 sg13g2_tielo \proj_12.flop8/_1__18  (.L_LO(net18));
 sg13g2_tielo \proj_12.not1/_0__19  (.L_LO(net19));
 sg13g2_tielo \proj__0.flop1/_1__20  (.L_LO(net20));
 sg13g2_tielo \proj__3.and2/_0__21  (.L_LO(net21));
 sg13g2_tielo \proj__3.and3/_0__22  (.L_LO(net22));
 sg13g2_tielo \proj__8.flop11/_1__23  (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_group_10_24 (.L_LO(net24));
 sg13g2_tielo tt_um_wokwi_group_10_25 (.L_LO(net33));
 sg13g2_tielo tt_um_wokwi_group_10_26 (.L_LO(net34));
 sg13g2_tielo tt_um_wokwi_group_10_27 (.L_LO(net35));
 sg13g2_tielo tt_um_wokwi_group_10_28 (.L_LO(net36));
 sg13g2_tielo tt_um_wokwi_group_10_29 (.L_LO(net37));
 sg13g2_tielo tt_um_wokwi_group_10_30 (.L_LO(net38));
 sg13g2_tielo tt_um_wokwi_group_10_31 (.L_LO(net39));
 sg13g2_tielo tt_um_wokwi_group_10_32 (.L_LO(net40));
 sg13g2_tielo tt_um_wokwi_group_10_33 (.L_LO(net41));
 sg13g2_tielo tt_um_wokwi_group_10_34 (.L_LO(net42));
 sg13g2_tielo tt_um_wokwi_group_10_35 (.L_LO(net43));
 sg13g2_tielo tt_um_wokwi_group_10_36 (.L_LO(net44));
 sg13g2_tielo tt_um_wokwi_group_10_37 (.L_LO(net45));
 sg13g2_tielo tt_um_wokwi_group_10_38 (.L_LO(net46));
 sg13g2_tielo tt_um_wokwi_group_10_39 (.L_LO(net47));
 sg13g2_tiehi \proj_12.flop1/_1__40  (.L_HI(net48));
 sg13g2_and2_1 \proj_10.and1/_0_  (.A(net29),
    .B(net31),
    .X(\proj_10.net11 ));
 sg13g2_nand2_1 \proj_10.nand1/_0_  (.Y(\proj_10.net12 ),
    .A(net26),
    .B(net10));
 sg13g2_or2_1 \proj_10.or1/_0_  (.X(\proj_10.net10 ),
    .B(net32),
    .A(net28));
 sg13g2_dfrbp_1 \proj_12.flop1/_1_  (.CLK(net11),
    .RESET_B(net48),
    .D(\proj_12.net17 ),
    .Q_N(\proj_12.flop1/notq ),
    .Q(\proj_12.net3 ));
 sg13g2_tiehi \proj_12.flop2/_1__41  (.L_HI(net49));
 sg13g2_dfrbp_1 \proj_12.flop2/_1_  (.CLK(net12),
    .RESET_B(net49),
    .D(\proj_12.net3 ),
    .Q_N(\proj_12.flop2/notq ),
    .Q(\proj_12.net4 ));
 sg13g2_tiehi \proj_12.flop3/_1__42  (.L_HI(net50));
 sg13g2_dfrbp_1 \proj_12.flop3/_1_  (.CLK(net13),
    .RESET_B(net50),
    .D(\proj_12.net4 ),
    .Q_N(\proj_12.flop3/notq ),
    .Q(\proj_12.net5 ));
 sg13g2_tiehi \proj_12.flop4/_1__43  (.L_HI(net51));
 sg13g2_dfrbp_1 \proj_12.flop4/_1_  (.CLK(net14),
    .RESET_B(net51),
    .D(\proj_12.net7 ),
    .Q_N(\proj_12.flop4/notq ),
    .Q(\proj_12.net8 ));
 sg13g2_tiehi \proj_12.flop5/_1__44  (.L_HI(net52));
 sg13g2_dfrbp_1 \proj_12.flop5/_1_  (.CLK(net15),
    .RESET_B(net52),
    .D(\proj_12.net6 ),
    .Q_N(\proj_12.flop5/notq ),
    .Q(\proj_12.net7 ));
 sg13g2_tiehi \proj_12.flop6/_1__45  (.L_HI(net53));
 sg13g2_dfrbp_1 \proj_12.flop6/_1_  (.CLK(net16),
    .RESET_B(net53),
    .D(\proj_12.net8 ),
    .Q_N(\proj_12.flop6/notq ),
    .Q(\proj_12.net9 ));
 sg13g2_tiehi \proj_12.flop7/_1__46  (.L_HI(net54));
 sg13g2_dfrbp_1 \proj_12.flop7/_1_  (.CLK(net17),
    .RESET_B(net54),
    .D(\proj_12.net9 ),
    .Q_N(\proj_12.flop7/notq ),
    .Q(\proj_12.net10 ));
 sg13g2_tiehi \proj_12.flop8/_1__47  (.L_HI(net55));
 sg13g2_dfrbp_1 \proj_12.flop8/_1_  (.CLK(net18),
    .RESET_B(net55),
    .D(\proj_12.net5 ),
    .Q_N(\proj_12.flop8/notq ),
    .Q(\proj_12.net6 ));
 sg13g2_tiehi \proj__0.flop1/_1__48  (.L_HI(net56));
 sg13g2_inv_1 \proj_12.not1/_0_  (.Y(\proj_12.net20 ),
    .A(net19));
 sg13g2_or2_1 \proj_12.or1/_0_  (.X(\proj_12.net17 ),
    .B(\proj_12.net16 ),
    .A(\proj_12.net20 ));
 sg13g2_xor2_1 \proj_12.xor1/_0_  (.B(\proj_12.net10 ),
    .A(\proj_12.net15 ),
    .X(\proj_12.net16 ));
 sg13g2_xor2_1 \proj_12.xor2/_0_  (.B(\proj_12.net8 ),
    .A(\proj_12.net18 ),
    .X(\proj_12.net15 ));
 sg13g2_xor2_1 \proj_12.xor3/_0_  (.B(\proj_12.net7 ),
    .A(\proj_12.net6 ),
    .X(\proj_12.net18 ));
 sg13g2_and2_1 \proj_13.and1/_0_  (.A(net28),
    .B(net31),
    .X(\proj_13.net18 ));
 sg13g2_nand2_1 \proj_13.nand1/_0_  (.Y(\proj_13.net12 ),
    .A(net3),
    .B(net2));
 sg13g2_inv_1 \proj_13.not1/_0_  (.Y(\proj_13.net11 ),
    .A(net4));
 sg13g2_or2_1 \proj_13.or1/_0_  (.X(\proj_13.net19 ),
    .B(net27),
    .A(net1));
 sg13g2_or2_1 \proj_13.or2/_0_  (.X(\proj_13.net10 ),
    .B(\proj_13.net19 ),
    .A(\proj_13.net18 ));
 sg13g2_xor2_1 \proj_13.xor1/_0_  (.B(\proj_13.net18 ),
    .A(\proj_13.net19 ),
    .X(\proj_13.net9 ));
 sg13g2_nand2_1 \proj_14.nand1/_0_  (.Y(\proj_14.net7 ),
    .A(net28),
    .B(net32));
 sg13g2_dfrbp_1 \proj__0.flop1/_1_  (.CLK(net20),
    .RESET_B(net56),
    .D(\proj__0.net20 ),
    .Q_N(\proj__0.net7 ),
    .Q(\proj__0.net6 ));
 sg13g2_tiehi \proj__1.flop1/_1__49  (.L_HI(net57));
 sg13g2_inv_1 \proj__0.not1/_0_  (.Y(\proj__0.net13 ),
    .A(\proj__0.net12 ));
 sg13g2_inv_1 \proj__0.not2/_0_  (.Y(\proj__0.net14 ),
    .A(\proj__0.net13 ));
 sg13g2_inv_1 \proj__0.not3/_0_  (.Y(\proj__0.net12 ),
    .A(\proj__0.net14 ));
 sg13g2_inv_1 \proj__0.not4/_0_  (.Y(\proj__0.net16 ),
    .A(\proj__0.net15 ));
 sg13g2_inv_1 \proj__0.not5/_0_  (.Y(\proj__0.net17 ),
    .A(\proj__0.net16 ));
 sg13g2_inv_1 \proj__0.not6/_0_  (.Y(\proj__0.net18 ),
    .A(\proj__0.net17 ));
 sg13g2_inv_1 \proj__0.not7/_0_  (.Y(\proj__0.net19 ),
    .A(\proj__0.net18 ));
 sg13g2_inv_1 \proj__0.not8/_0_  (.Y(\proj__0.net15 ),
    .A(\proj__0.net19 ));
 sg13g2_xor2_1 \proj__0.xor1/_0_  (.B(\proj__0.net15 ),
    .A(\proj__0.net12 ),
    .X(\proj__0.net20 ));
 sg13g2_dfrbp_1 \proj__1.flop1/_1_  (.CLK(\proj__1.net14 ),
    .RESET_B(net57),
    .D(\proj__1.net13 ),
    .Q_N(\proj__1.net13 ),
    .Q(\proj__1.net15 ));
 sg13g2_tiehi \proj__1.flop2/_1__50  (.L_HI(net58));
 sg13g2_dfrbp_1 \proj__1.flop2/_1_  (.CLK(net2),
    .RESET_B(net58),
    .D(\proj__1.net16 ),
    .Q_N(\proj__1.net16 ),
    .Q(\proj__1.net14 ));
 sg13g2_tiehi \proj__1.flop3/_1__51  (.L_HI(net59));
 sg13g2_dfrbp_1 \proj__1.flop3/_1_  (.CLK(\proj__1.net15 ),
    .RESET_B(net59),
    .D(\proj__1.net17 ),
    .Q_N(\proj__1.net17 ),
    .Q(\proj__1.net18 ));
 sg13g2_tiehi \proj__1.flop4/_1__52  (.L_HI(net60));
 sg13g2_dfrbp_1 \proj__1.flop4/_1_  (.CLK(\proj__1.net21 ),
    .RESET_B(net60),
    .D(\proj__1.net20 ),
    .Q_N(\proj__1.net20 ),
    .Q(\proj__1.net22 ));
 sg13g2_tiehi \proj__1.flop5/_1__53  (.L_HI(net61));
 sg13g2_dfrbp_1 \proj__1.flop5/_1_  (.CLK(\proj__1.net18 ),
    .RESET_B(net61),
    .D(\proj__1.net23 ),
    .Q_N(\proj__1.net23 ),
    .Q(\proj__1.net21 ));
 sg13g2_tiehi \proj__1.flop6/_1__54  (.L_HI(net62));
 sg13g2_dfrbp_1 \proj__1.flop6/_1_  (.CLK(\proj__1.net22 ),
    .RESET_B(net62),
    .D(\proj__1.net24 ),
    .Q_N(\proj__1.net24 ),
    .Q(\proj__1.net25 ));
 sg13g2_tiehi \proj__1.flop7/_1__55  (.L_HI(net63));
 sg13g2_dfrbp_1 \proj__1.flop7/_1_  (.CLK(\proj__1.net25 ),
    .RESET_B(net63),
    .D(\proj__1.net28 ),
    .Q_N(\proj__1.net28 ),
    .Q(\proj__1.net29 ));
 sg13g2_tiehi \proj__8.flop1/_1__56  (.L_HI(net64));
 sg13g2_mux2_1 \proj__1.mux1/_0_  (.A0(\proj__1.net14 ),
    .A1(\proj__1.net6 ),
    .S(net28),
    .X(\proj__1.net19 ));
 sg13g2_mux2_1 \proj__1.mux2/_0_  (.A0(\proj__1.net18 ),
    .A1(\proj__1.net15 ),
    .S(net30),
    .X(\proj__1.net26 ));
 sg13g2_mux2_1 \proj__1.mux3/_0_  (.A0(\proj__1.net22 ),
    .A1(\proj__1.net21 ),
    .S(net30),
    .X(\proj__1.net27 ));
 sg13g2_mux2_1 \proj__1.mux4/_0_  (.A0(\proj__1.net29 ),
    .A1(\proj__1.net25 ),
    .S(net30),
    .X(\proj__1.net30 ));
 sg13g2_mux2_1 \proj__1.mux5/_0_  (.A0(\proj__1.net30 ),
    .A1(\proj__1.net27 ),
    .S(net27),
    .X(\proj__1.net31 ));
 sg13g2_mux2_1 \proj__1.mux6/_0_  (.A0(\proj__1.net26 ),
    .A1(\proj__1.net19 ),
    .S(net27),
    .X(\proj__1.net32 ));
 sg13g2_mux2_1 \proj__1.mux7/_0_  (.A0(\proj__1.net31 ),
    .A1(\proj__1.net32 ),
    .S(net1),
    .X(\proj__1.net7 ));
 sg13g2_inv_1 \proj__1.not5/_0_  (.Y(\proj__1.net8 ),
    .A(net32));
 sg13g2_inv_1 \proj__1.not6/_0_  (.Y(\proj__1.net10 ),
    .A(\proj__1.net8 ));
 sg13g2_inv_1 \proj__1.not7/_0_  (.Y(\proj__1.net11 ),
    .A(\proj__1.net10 ));
 sg13g2_inv_1 \proj__1.not8/_0_  (.Y(\proj__1.net12 ),
    .A(\proj__1.net11 ));
 sg13g2_inv_1 \proj__1.not9/_0_  (.Y(\proj__1.net6 ),
    .A(\proj__1.net12 ));
 sg13g2_inv_1 \proj__2.not1/_0_  (.Y(\proj__2.net9 ),
    .A(net31));
 sg13g2_inv_1 \proj__2.not2/_0_  (.Y(\proj__2.net10 ),
    .A(net29));
 sg13g2_inv_1 \proj__2.not3/_0_  (.Y(\proj__2.net11 ),
    .A(net26));
 sg13g2_inv_1 \proj__2.not4/_0_  (.Y(\proj__2.net12 ),
    .A(net1));
 sg13g2_and2_1 \proj__3.and1/_0_  (.A(\proj__3.net13 ),
    .B(\proj__3.net12 ),
    .X(\proj__3.net6 ));
 sg13g2_and2_1 \proj__3.and2/_0_  (.A(net21),
    .B(net4),
    .X(\proj__3.net13 ));
 sg13g2_and2_1 \proj__3.and3/_0_  (.A(net22),
    .B(net32),
    .X(\proj__3.net12 ));
 sg13g2_and2_1 \proj__4.and1/_0_  (.A(net3),
    .B(net26),
    .X(\proj__4.net11 ));
 sg13g2_nand2_1 \proj__4.nand1/_0_  (.Y(\proj__4.net9 ),
    .A(net28),
    .B(\proj__4.net18 ));
 sg13g2_inv_1 \proj__4.not1/_0_  (.Y(\proj__4.net12 ),
    .A(net1));
 sg13g2_or2_1 \proj__4.or1/_0_  (.X(\proj__4.net10 ),
    .B(net31),
    .A(net26));
 sg13g2_xor2_1 \proj__4.xor1/_0_  (.B(net31),
    .A(net28),
    .X(\proj__4.net18 ));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net1),
    .B(net26),
    .X(\proj__5.net12 ));
 sg13g2_nand2_1 \proj__5.nand1/_0_  (.Y(\proj__5.net11 ),
    .A(net26),
    .B(net1));
 sg13g2_inv_1 \proj__5.not1/_0_  (.Y(\proj__5.net14 ),
    .A(net5));
 sg13g2_inv_1 \proj__5.not2/_0_  (.Y(\proj__5.net13 ),
    .A(net3));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net10 ),
    .B(net31),
    .A(net29));
 sg13g2_xor2_1 \proj__5.xor1/_0_  (.B(net32),
    .A(net28),
    .X(\proj__5.net9 ));
 sg13g2_and2_1 \proj__6.and1/_0_  (.A(net26),
    .B(net28),
    .X(\proj__6.net9 ));
 sg13g2_inv_1 \proj__6.not1/_0_  (.Y(\proj__6.net8 ),
    .A(net31));
 sg13g2_or2_1 \proj__6.or1/_0_  (.X(\proj__6.net10 ),
    .B(net1),
    .A(net2));
 sg13g2_xor2_1 \proj__6.xor1/_0_  (.B(net3),
    .A(net4),
    .X(\proj__6.net11 ));
 sg13g2_and2_1 \proj__7.and1/_0_  (.A(net29),
    .B(net31),
    .X(\proj__7.net9 ));
 sg13g2_xor2_1 \proj__7.xor1/_0_  (.B(net4),
    .A(net5),
    .X(\proj__7.net10 ));
 sg13g2_dfrbp_1 \proj__8.flop1/_1_  (.CLK(\proj__8.net15 ),
    .RESET_B(net64),
    .D(\proj__8.net2 ),
    .Q_N(\proj__8.flop1/notq ),
    .Q(\proj__8.net3 ));
 sg13g2_tiehi \proj__8.flop10/_1__57  (.L_HI(net65));
 sg13g2_dfrbp_1 \proj__8.flop10/_1_  (.CLK(\proj__8.net26 ),
    .RESET_B(net65),
    .D(\proj__8.net25 ),
    .Q_N(\proj__8.flop10/notq ),
    .Q(\proj__8.net23 ));
 sg13g2_tiehi \proj__8.flop11/_1__58  (.L_HI(net66));
 sg13g2_dfrbp_1 \proj__8.flop11/_1_  (.CLK(net23),
    .RESET_B(net66),
    .D(\proj__8.net27 ),
    .Q_N(\proj__8.flop11/notq ),
    .Q(\proj__8.net26 ));
 sg13g2_tiehi \proj__8.flop12/_1__59  (.L_HI(net67));
 sg13g2_dfrbp_1 \proj__8.flop12/_1_  (.CLK(\proj__8.net24 ),
    .RESET_B(net67),
    .D(\proj__8.net28 ),
    .Q_N(\proj__8.flop12/notq ),
    .Q(\proj__8.net29 ));
 sg13g2_tiehi \proj__8.flop13/_1__60  (.L_HI(net68));
 sg13g2_dfrbp_1 \proj__8.flop13/_1_  (.CLK(\proj__8.net31 ),
    .RESET_B(net68),
    .D(\proj__8.net30 ),
    .Q_N(\proj__8.flop13/notq ),
    .Q(\proj__8.net32 ));
 sg13g2_tiehi \proj__8.flop14/_1__61  (.L_HI(net69));
 sg13g2_dfrbp_1 \proj__8.flop14/_1_  (.CLK(\proj__8.net34 ),
    .RESET_B(net69),
    .D(\proj__8.net33 ),
    .Q_N(\proj__8.flop14/notq ),
    .Q(\proj__8.net31 ));
 sg13g2_tiehi \proj__8.flop15/_1__62  (.L_HI(net70));
 sg13g2_dfrbp_1 \proj__8.flop15/_1_  (.CLK(\proj__8.net29 ),
    .RESET_B(net70),
    .D(\proj__8.net35 ),
    .Q_N(\proj__8.flop15/notq ),
    .Q(\proj__8.net34 ));
 sg13g2_tiehi \proj__8.flop16/_1__63  (.L_HI(net71));
 sg13g2_dfrbp_1 \proj__8.flop16/_1_  (.CLK(\proj__8.net32 ),
    .RESET_B(net71),
    .D(\proj__8.net36 ),
    .Q_N(\proj__8.net38 ),
    .Q(\proj__8.net37 ));
 sg13g2_tiehi \proj__8.flop17/_1__64  (.L_HI(net72));
 sg13g2_dfrbp_1 \proj__8.flop17/_1_  (.CLK(\proj__8.net40 ),
    .RESET_B(net72),
    .D(\proj__8.net39 ),
    .Q_N(\proj__8.flop17/notq ),
    .Q(\proj__8.net41 ));
 sg13g2_tiehi \proj__8.flop18/_1__65  (.L_HI(net73));
 sg13g2_dfrbp_1 \proj__8.flop18/_1_  (.CLK(\proj__8.net43 ),
    .RESET_B(net73),
    .D(\proj__8.net42 ),
    .Q_N(\proj__8.flop18/notq ),
    .Q(\proj__8.net40 ));
 sg13g2_tiehi \proj__8.flop19/_1__66  (.L_HI(net74));
 sg13g2_dfrbp_1 \proj__8.flop19/_1_  (.CLK(\proj__8.net38 ),
    .RESET_B(net74),
    .D(\proj__8.net44 ),
    .Q_N(\proj__8.flop19/notq ),
    .Q(\proj__8.net43 ));
 sg13g2_tiehi \proj__8.flop2/_1__67  (.L_HI(net75));
 sg13g2_dfrbp_1 \proj__8.flop2/_1_  (.CLK(\proj__8.net15 ),
    .RESET_B(net75),
    .D(\proj__8.net3 ),
    .Q_N(\proj__8.flop2/notq ),
    .Q(\proj__8.net4 ));
 sg13g2_tiehi \proj__8.flop20/_1__68  (.L_HI(net76));
 sg13g2_dfrbp_1 \proj__8.flop20/_1_  (.CLK(\proj__8.net41 ),
    .RESET_B(net76),
    .D(\proj__8.net45 ),
    .Q_N(\proj__8.flop20/notq ),
    .Q(\proj__8.net46 ));
 sg13g2_tiehi \proj__8.flop21/_1__69  (.L_HI(net77));
 sg13g2_dfrbp_1 \proj__8.flop21/_1_  (.CLK(\proj__8.net46 ),
    .RESET_B(net77),
    .D(\proj__8.net47 ),
    .Q_N(\proj__8.net15 ),
    .Q(\proj__8.net48 ));
 sg13g2_tiehi \proj__8.flop3/_1__70  (.L_HI(net78));
 sg13g2_dfrbp_1 \proj__8.flop3/_1_  (.CLK(\proj__8.net15 ),
    .RESET_B(net78),
    .D(\proj__8.net4 ),
    .Q_N(\proj__8.flop3/notq ),
    .Q(\proj__8.net5 ));
 sg13g2_tiehi \proj__8.flop4/_1__71  (.L_HI(net79));
 sg13g2_dfrbp_1 \proj__8.flop4/_1_  (.CLK(\proj__8.net15 ),
    .RESET_B(net79),
    .D(\proj__8.net5 ),
    .Q_N(\proj__8.flop4/notq ),
    .Q(\proj__8.net6 ));
 sg13g2_tiehi \proj__8.flop5/_1__72  (.L_HI(net80));
 sg13g2_dfrbp_1 \proj__8.flop5/_1_  (.CLK(\proj__8.net15 ),
    .RESET_B(net80),
    .D(\proj__8.net16 ),
    .Q_N(\proj__8.flop5/notq ),
    .Q(\proj__8.net2 ));
 sg13g2_tiehi \proj__8.flop6/_1__73  (.L_HI(net81));
 sg13g2_dfrbp_1 \proj__8.flop6/_1_  (.CLK(\proj__8.net15 ),
    .RESET_B(net81),
    .D(\proj__8.net6 ),
    .Q_N(\proj__8.flop6/notq ),
    .Q(\proj__8.net7 ));
 sg13g2_tiehi \proj__8.flop7/_1__74  (.L_HI(net82));
 sg13g2_dfrbp_1 \proj__8.flop7/_1_  (.CLK(\proj__8.net15 ),
    .RESET_B(net82),
    .D(\proj__8.net7 ),
    .Q_N(\proj__8.flop7/notq ),
    .Q(\proj__8.net8 ));
 sg13g2_tiehi \proj__8.flop8/_1__75  (.L_HI(net83));
 sg13g2_dfrbp_1 \proj__8.flop8/_1_  (.CLK(\proj__8.net15 ),
    .RESET_B(net83),
    .D(\proj__8.net8 ),
    .Q_N(\proj__8.flop8/notq ),
    .Q(\proj__8.net9 ));
 sg13g2_tiehi \proj__8.flop9/_1__76  (.L_HI(net84));
 sg13g2_dfrbp_1 \proj__8.flop9/_1_  (.CLK(\proj__8.net23 ),
    .RESET_B(net84),
    .D(\proj__8.net22 ),
    .Q_N(\proj__8.flop9/notq ),
    .Q(\proj__8.net24 ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_inv_1 \proj__8.not1/_0_  (.Y(\proj__8.net16 ),
    .A(\proj__8.net17 ));
 sg13g2_inv_1 \proj__8.not10/_0_  (.Y(\proj__8.net35 ),
    .A(\proj__8.net34 ));
 sg13g2_inv_1 \proj__8.not11/_0_  (.Y(\proj__8.net36 ),
    .A(\proj__8.net37 ));
 sg13g2_inv_1 \proj__8.not12/_0_  (.Y(\proj__8.net39 ),
    .A(\proj__8.net41 ));
 sg13g2_inv_1 \proj__8.not13/_0_  (.Y(\proj__8.net42 ),
    .A(\proj__8.net40 ));
 sg13g2_inv_1 \proj__8.not14/_0_  (.Y(\proj__8.net44 ),
    .A(\proj__8.net43 ));
 sg13g2_inv_1 \proj__8.not15/_0_  (.Y(\proj__8.net45 ),
    .A(\proj__8.net46 ));
 sg13g2_inv_1 \proj__8.not16/_0_  (.Y(\proj__8.net47 ),
    .A(\proj__8.net48 ));
 sg13g2_inv_1 \proj__8.not2/_0_  (.Y(\proj__8.net18 ),
    .A(\proj__8.net19 ));
 sg13g2_inv_1 \proj__8.not3/_0_  (.Y(\proj__8.net20 ),
    .A(\proj__8.net21 ));
 sg13g2_inv_1 \proj__8.not4/_0_  (.Y(\proj__8.net22 ),
    .A(\proj__8.net24 ));
 sg13g2_inv_1 \proj__8.not5/_0_  (.Y(\proj__8.net25 ),
    .A(\proj__8.net23 ));
 sg13g2_inv_1 \proj__8.not6/_0_  (.Y(\proj__8.net27 ),
    .A(\proj__8.net26 ));
 sg13g2_inv_1 \proj__8.not7/_0_  (.Y(\proj__8.net28 ),
    .A(\proj__8.net29 ));
 sg13g2_inv_1 \proj__8.not8/_0_  (.Y(\proj__8.net30 ),
    .A(\proj__8.net32 ));
 sg13g2_inv_1 \proj__8.not9/_0_  (.Y(\proj__8.net33 ),
    .A(\proj__8.net31 ));
 sg13g2_xor2_1 \proj__8.xor1/_0_  (.B(\proj__8.net18 ),
    .A(\proj__8.net5 ),
    .X(\proj__8.net17 ));
 sg13g2_xor2_1 \proj__8.xor2/_0_  (.B(\proj__8.net20 ),
    .A(\proj__8.net6 ),
    .X(\proj__8.net19 ));
 sg13g2_xor2_1 \proj__8.xor3/_0_  (.B(\proj__8.net9 ),
    .A(\proj__8.net7 ),
    .X(\proj__8.net21 ));
 sg13g2_and2_1 \proj__9.and1/_0_  (.A(net30),
    .B(net32),
    .X(\proj__9.net11 ));
 sg13g2_and2_1 \proj__9.and2/_0_  (.A(net27),
    .B(\proj__9.net10 ),
    .X(\proj__9.net12 ));
 sg13g2_or2_1 \proj__9.or1/_0_  (.X(\proj__9.net5 ),
    .B(\proj__9.net11 ),
    .A(\proj__9.net12 ));
 sg13g2_xor2_1 \proj__9.xor1/_0_  (.B(net32),
    .A(net30),
    .X(\proj__9.net10 ));
 sg13g2_xor2_1 \proj__9.xor2/_0_  (.B(\proj__9.net10 ),
    .A(net27),
    .X(\proj__9.net4 ));
 sg13g2_buf_2 fanout25 (.A(net9),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(net27),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(ui_in[2]),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(net30),
    .X(net28));
 sg13g2_buf_1 fanout29 (.A(net30),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(ui_in[1]),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(net32),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(ui_in[0]),
    .X(net32));
 sg13g2_buf_2 input1 (.A(ui_in[3]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[4]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[6]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_tielo \proj_10.nand1/_0__10  (.L_LO(net10));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_4 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_4 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_decap_8 FILLER_27_246 ();
 sg13g2_decap_8 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_decap_4 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_339 ();
 sg13g2_decap_4 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_fill_1 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_4 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_decap_4 FILLER_29_246 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_4 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_decap_4 FILLER_29_323 ();
 sg13g2_fill_1 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_decap_8 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_29_352 ();
 sg13g2_fill_2 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_4 FILLER_29_377 ();
 sg13g2_fill_2 FILLER_29_391 ();
 sg13g2_fill_1 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_4 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_177 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_fill_2 FILLER_30_184 ();
 sg13g2_fill_1 FILLER_30_190 ();
 sg13g2_fill_2 FILLER_30_195 ();
 sg13g2_decap_4 FILLER_30_201 ();
 sg13g2_fill_2 FILLER_30_205 ();
 sg13g2_decap_8 FILLER_30_237 ();
 sg13g2_decap_4 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_265 ();
 sg13g2_decap_8 FILLER_30_272 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_2 FILLER_30_299 ();
 sg13g2_fill_1 FILLER_30_306 ();
 sg13g2_decap_4 FILLER_30_315 ();
 sg13g2_fill_2 FILLER_30_319 ();
 sg13g2_fill_2 FILLER_30_381 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_160 ();
 sg13g2_decap_8 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_decap_8 FILLER_31_208 ();
 sg13g2_decap_4 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_225 ();
 sg13g2_decap_4 FILLER_31_235 ();
 sg13g2_fill_2 FILLER_31_239 ();
 sg13g2_fill_2 FILLER_31_291 ();
 sg13g2_decap_8 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_decap_4 FILLER_31_329 ();
 sg13g2_fill_2 FILLER_31_333 ();
 sg13g2_fill_2 FILLER_31_349 ();
 sg13g2_fill_1 FILLER_31_354 ();
 sg13g2_fill_2 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_fill_2 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_4 FILLER_32_208 ();
 sg13g2_fill_2 FILLER_32_212 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_decap_4 FILLER_32_225 ();
 sg13g2_fill_2 FILLER_32_235 ();
 sg13g2_fill_1 FILLER_32_237 ();
 sg13g2_decap_4 FILLER_32_243 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_decap_4 FILLER_32_260 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_2 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_decap_4 FILLER_32_334 ();
 sg13g2_fill_1 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_fill_2 FILLER_32_361 ();
 sg13g2_fill_1 FILLER_32_363 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_30 ();
 sg13g2_decap_8 FILLER_33_37 ();
 sg13g2_decap_8 FILLER_33_44 ();
 sg13g2_decap_8 FILLER_33_51 ();
 sg13g2_decap_8 FILLER_33_58 ();
 sg13g2_decap_8 FILLER_33_65 ();
 sg13g2_decap_8 FILLER_33_72 ();
 sg13g2_decap_8 FILLER_33_79 ();
 sg13g2_decap_8 FILLER_33_86 ();
 sg13g2_decap_8 FILLER_33_93 ();
 sg13g2_decap_8 FILLER_33_100 ();
 sg13g2_decap_8 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_114 ();
 sg13g2_decap_8 FILLER_33_121 ();
 sg13g2_decap_8 FILLER_33_128 ();
 sg13g2_decap_8 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_142 ();
 sg13g2_decap_8 FILLER_33_149 ();
 sg13g2_decap_8 FILLER_33_156 ();
 sg13g2_decap_8 FILLER_33_163 ();
 sg13g2_fill_2 FILLER_33_200 ();
 sg13g2_fill_1 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_decap_8 FILLER_33_267 ();
 sg13g2_decap_4 FILLER_33_274 ();
 sg13g2_fill_2 FILLER_33_283 ();
 sg13g2_decap_8 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_317 ();
 sg13g2_fill_2 FILLER_33_329 ();
 sg13g2_decap_4 FILLER_33_337 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_fill_1 FILLER_33_351 ();
 sg13g2_fill_2 FILLER_33_367 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_2 FILLER_33_391 ();
 sg13g2_fill_1 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_4 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_179 ();
 sg13g2_decap_8 FILLER_34_185 ();
 sg13g2_decap_8 FILLER_34_192 ();
 sg13g2_decap_8 FILLER_34_199 ();
 sg13g2_decap_8 FILLER_34_206 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_4 FILLER_34_238 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_decap_4 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_306 ();
 sg13g2_decap_8 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_320 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_decap_4 FILLER_34_340 ();
 sg13g2_decap_4 FILLER_34_360 ();
 sg13g2_fill_2 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_370 ();
 sg13g2_fill_2 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_decap_4 FILLER_35_11 ();
 sg13g2_fill_1 FILLER_35_19 ();
 sg13g2_decap_8 FILLER_35_24 ();
 sg13g2_decap_8 FILLER_35_31 ();
 sg13g2_decap_8 FILLER_35_38 ();
 sg13g2_decap_8 FILLER_35_48 ();
 sg13g2_decap_8 FILLER_35_55 ();
 sg13g2_decap_8 FILLER_35_62 ();
 sg13g2_decap_8 FILLER_35_69 ();
 sg13g2_fill_2 FILLER_35_76 ();
 sg13g2_fill_2 FILLER_35_81 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_145 ();
 sg13g2_decap_8 FILLER_35_152 ();
 sg13g2_decap_8 FILLER_35_159 ();
 sg13g2_decap_8 FILLER_35_166 ();
 sg13g2_decap_8 FILLER_35_173 ();
 sg13g2_decap_8 FILLER_35_180 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_253 ();
 sg13g2_decap_8 FILLER_35_264 ();
 sg13g2_decap_4 FILLER_35_280 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_fill_1 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_30 ();
 sg13g2_fill_1 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_88 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_fill_1 FILLER_36_99 ();
 sg13g2_decap_8 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_decap_8 FILLER_36_202 ();
 sg13g2_fill_2 FILLER_36_209 ();
 sg13g2_decap_8 FILLER_36_222 ();
 sg13g2_fill_2 FILLER_36_229 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_2 FILLER_36_269 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_decap_8 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_2 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_19 ();
 sg13g2_decap_4 FILLER_37_47 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_76 ();
 sg13g2_decap_8 FILLER_37_83 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_decap_8 FILLER_37_97 ();
 sg13g2_decap_8 FILLER_37_104 ();
 sg13g2_decap_8 FILLER_37_111 ();
 sg13g2_decap_8 FILLER_37_118 ();
 sg13g2_decap_8 FILLER_37_125 ();
 sg13g2_decap_4 FILLER_37_132 ();
 sg13g2_fill_1 FILLER_37_136 ();
 sg13g2_decap_4 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_145 ();
 sg13g2_decap_4 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_234 ();
 sg13g2_decap_8 FILLER_37_241 ();
 sg13g2_decap_4 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_304 ();
 sg13g2_fill_1 FILLER_37_323 ();
 sg13g2_fill_2 FILLER_37_333 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_341 ();
 sg13g2_fill_1 FILLER_37_347 ();
 sg13g2_decap_8 FILLER_37_360 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_374 ();
 sg13g2_decap_8 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_31 ();
 sg13g2_decap_8 FILLER_38_38 ();
 sg13g2_decap_8 FILLER_38_45 ();
 sg13g2_decap_4 FILLER_38_52 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_176 ();
 sg13g2_decap_8 FILLER_38_185 ();
 sg13g2_decap_4 FILLER_38_192 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_207 ();
 sg13g2_fill_2 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_248 ();
 sg13g2_decap_4 FILLER_38_255 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_decap_8 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_277 ();
 sg13g2_fill_2 FILLER_38_286 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_decap_8 FILLER_38_363 ();
 sg13g2_decap_8 FILLER_38_370 ();
 sg13g2_decap_8 FILLER_38_377 ();
 sg13g2_decap_8 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net24;
 assign uio_oe[1] = net33;
 assign uio_oe[2] = net34;
 assign uio_oe[3] = net35;
 assign uio_oe[4] = net36;
 assign uio_oe[5] = net37;
 assign uio_oe[6] = net38;
 assign uio_oe[7] = net39;
 assign uio_out[0] = net40;
 assign uio_out[1] = net41;
 assign uio_out[2] = net42;
 assign uio_out[3] = net43;
 assign uio_out[4] = net44;
 assign uio_out[5] = net45;
 assign uio_out[6] = net46;
 assign uio_out[7] = net47;
endmodule

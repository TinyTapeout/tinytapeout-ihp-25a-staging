module tt_um_ece298a_8_bit_cpu_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire CF;
 wire Cp;
 wire HF;
 wire Lp;
 wire ZF;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire clk_regs;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire \accumulator_object.bus[0] ;
 wire \accumulator_object.bus[1] ;
 wire \accumulator_object.bus[2] ;
 wire \accumulator_object.bus[3] ;
 wire \accumulator_object.bus[4] ;
 wire \accumulator_object.bus[5] ;
 wire \accumulator_object.bus[6] ;
 wire \accumulator_object.bus[7] ;
 wire \accumulator_object.load ;
 wire \alu_object.addsub.genblk1[0].fa.a ;
 wire \alu_object.addsub.genblk1[0].fa.cin ;
 wire \alu_object.addsub.genblk1[0].fa.sum ;
 wire \alu_object.addsub.genblk1[1].fa.a ;
 wire \alu_object.addsub.genblk1[1].fa.sum ;
 wire \alu_object.addsub.genblk1[2].fa.a ;
 wire \alu_object.addsub.genblk1[2].fa.sum ;
 wire \alu_object.addsub.genblk1[3].fa.a ;
 wire \alu_object.addsub.genblk1[3].fa.sum ;
 wire \alu_object.addsub.genblk1[4].fa.a ;
 wire \alu_object.addsub.genblk1[4].fa.sum ;
 wire \alu_object.addsub.genblk1[5].fa.a ;
 wire \alu_object.addsub.genblk1[5].fa.sum ;
 wire \alu_object.addsub.genblk1[6].fa.a ;
 wire \alu_object.addsub.genblk1[6].fa.sum ;
 wire \alu_object.addsub.genblk1[7].fa.a ;
 wire \alu_object.addsub.genblk1[7].fa.sum ;
 wire \alu_object.addsub.op_b[0] ;
 wire \alu_object.addsub.op_b[1] ;
 wire \alu_object.addsub.op_b[2] ;
 wire \alu_object.addsub.op_b[3] ;
 wire \alu_object.addsub.op_b[4] ;
 wire \alu_object.addsub.op_b[5] ;
 wire \alu_object.addsub.op_b[6] ;
 wire \alu_object.addsub.op_b[7] ;
 wire \b_register.n_load ;
 wire \cb.control_signals[0] ;
 wire \cb.control_signals[10] ;
 wire \cb.control_signals[11] ;
 wire \cb.control_signals[13] ;
 wire \cb.control_signals[2] ;
 wire \cb.control_signals[4] ;
 wire \cb.control_signals[6] ;
 wire \cb.control_signals[7] ;
 wire \cb.control_signals[8] ;
 wire \cb.control_signals[9] ;
 wire \cb.done_load ;
 wire \cb.read_ui_in ;
 wire \cb.stage[0] ;
 wire \cb.stage[1] ;
 wire \cb.stage[2] ;
 wire \input_mar_register.addr[0] ;
 wire \input_mar_register.addr[1] ;
 wire \input_mar_register.addr[2] ;
 wire \input_mar_register.addr[3] ;
 wire \input_mar_register.data[0] ;
 wire \input_mar_register.data[1] ;
 wire \input_mar_register.data[2] ;
 wire \input_mar_register.data[3] ;
 wire \input_mar_register.data[4] ;
 wire \input_mar_register.data[5] ;
 wire \input_mar_register.data[6] ;
 wire \input_mar_register.data[7] ;
 wire \instruction_register.instruction[0] ;
 wire \instruction_register.instruction[1] ;
 wire \instruction_register.instruction[2] ;
 wire \instruction_register.instruction[3] ;
 wire \instruction_register.instruction[4] ;
 wire \instruction_register.instruction[5] ;
 wire \instruction_register.instruction[6] ;
 wire \instruction_register.instruction[7] ;
 wire \pc.set_bit_0.S ;
 wire \pc.set_bit_1.S ;
 wire \pc.set_bit_2.S ;
 wire \pc.set_bit_3.S ;
 wire \ram.RAM[0][0] ;
 wire \ram.RAM[0][1] ;
 wire \ram.RAM[0][2] ;
 wire \ram.RAM[0][3] ;
 wire \ram.RAM[0][4] ;
 wire \ram.RAM[0][5] ;
 wire \ram.RAM[0][6] ;
 wire \ram.RAM[0][7] ;
 wire \ram.RAM[10][0] ;
 wire \ram.RAM[10][1] ;
 wire \ram.RAM[10][2] ;
 wire \ram.RAM[10][3] ;
 wire \ram.RAM[10][4] ;
 wire \ram.RAM[10][5] ;
 wire \ram.RAM[10][6] ;
 wire \ram.RAM[10][7] ;
 wire \ram.RAM[11][0] ;
 wire \ram.RAM[11][1] ;
 wire \ram.RAM[11][2] ;
 wire \ram.RAM[11][3] ;
 wire \ram.RAM[11][4] ;
 wire \ram.RAM[11][5] ;
 wire \ram.RAM[11][6] ;
 wire \ram.RAM[11][7] ;
 wire \ram.RAM[12][0] ;
 wire \ram.RAM[12][1] ;
 wire \ram.RAM[12][2] ;
 wire \ram.RAM[12][3] ;
 wire \ram.RAM[12][4] ;
 wire \ram.RAM[12][5] ;
 wire \ram.RAM[12][6] ;
 wire \ram.RAM[12][7] ;
 wire \ram.RAM[13][0] ;
 wire \ram.RAM[13][1] ;
 wire \ram.RAM[13][2] ;
 wire \ram.RAM[13][3] ;
 wire \ram.RAM[13][4] ;
 wire \ram.RAM[13][5] ;
 wire \ram.RAM[13][6] ;
 wire \ram.RAM[13][7] ;
 wire \ram.RAM[14][0] ;
 wire \ram.RAM[14][1] ;
 wire \ram.RAM[14][2] ;
 wire \ram.RAM[14][3] ;
 wire \ram.RAM[14][4] ;
 wire \ram.RAM[14][5] ;
 wire \ram.RAM[14][6] ;
 wire \ram.RAM[14][7] ;
 wire \ram.RAM[15][0] ;
 wire \ram.RAM[15][1] ;
 wire \ram.RAM[15][2] ;
 wire \ram.RAM[15][3] ;
 wire \ram.RAM[15][4] ;
 wire \ram.RAM[15][5] ;
 wire \ram.RAM[15][6] ;
 wire \ram.RAM[15][7] ;
 wire \ram.RAM[1][0] ;
 wire \ram.RAM[1][1] ;
 wire \ram.RAM[1][2] ;
 wire \ram.RAM[1][3] ;
 wire \ram.RAM[1][4] ;
 wire \ram.RAM[1][5] ;
 wire \ram.RAM[1][6] ;
 wire \ram.RAM[1][7] ;
 wire \ram.RAM[2][0] ;
 wire \ram.RAM[2][1] ;
 wire \ram.RAM[2][2] ;
 wire \ram.RAM[2][3] ;
 wire \ram.RAM[2][4] ;
 wire \ram.RAM[2][5] ;
 wire \ram.RAM[2][6] ;
 wire \ram.RAM[2][7] ;
 wire \ram.RAM[3][0] ;
 wire \ram.RAM[3][1] ;
 wire \ram.RAM[3][2] ;
 wire \ram.RAM[3][3] ;
 wire \ram.RAM[3][4] ;
 wire \ram.RAM[3][5] ;
 wire \ram.RAM[3][6] ;
 wire \ram.RAM[3][7] ;
 wire \ram.RAM[4][0] ;
 wire \ram.RAM[4][1] ;
 wire \ram.RAM[4][2] ;
 wire \ram.RAM[4][3] ;
 wire \ram.RAM[4][4] ;
 wire \ram.RAM[4][5] ;
 wire \ram.RAM[4][6] ;
 wire \ram.RAM[4][7] ;
 wire \ram.RAM[5][0] ;
 wire \ram.RAM[5][1] ;
 wire \ram.RAM[5][2] ;
 wire \ram.RAM[5][3] ;
 wire \ram.RAM[5][4] ;
 wire \ram.RAM[5][5] ;
 wire \ram.RAM[5][6] ;
 wire \ram.RAM[5][7] ;
 wire \ram.RAM[6][0] ;
 wire \ram.RAM[6][1] ;
 wire \ram.RAM[6][2] ;
 wire \ram.RAM[6][3] ;
 wire \ram.RAM[6][4] ;
 wire \ram.RAM[6][5] ;
 wire \ram.RAM[6][6] ;
 wire \ram.RAM[6][7] ;
 wire \ram.RAM[7][0] ;
 wire \ram.RAM[7][1] ;
 wire \ram.RAM[7][2] ;
 wire \ram.RAM[7][3] ;
 wire \ram.RAM[7][4] ;
 wire \ram.RAM[7][5] ;
 wire \ram.RAM[7][6] ;
 wire \ram.RAM[7][7] ;
 wire \ram.RAM[8][0] ;
 wire \ram.RAM[8][1] ;
 wire \ram.RAM[8][2] ;
 wire \ram.RAM[8][3] ;
 wire \ram.RAM[8][4] ;
 wire \ram.RAM[8][5] ;
 wire \ram.RAM[8][6] ;
 wire \ram.RAM[8][7] ;
 wire \ram.RAM[9][0] ;
 wire \ram.RAM[9][1] ;
 wire \ram.RAM[9][2] ;
 wire \ram.RAM[9][3] ;
 wire \ram.RAM[9][4] ;
 wire \ram.RAM[9][5] ;
 wire \ram.RAM[9][6] ;
 wire \ram.RAM[9][7] ;
 wire net19;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire delaynet_0_clk;
 wire delaynet_1_clk;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;

 sg13g2_inv_1 _1016_ (.Y(_0254_),
    .A(net580));
 sg13g2_inv_1 _1017_ (.Y(_0255_),
    .A(net582));
 sg13g2_inv_1 _1018_ (.Y(_0256_),
    .A(net586));
 sg13g2_inv_2 _1019_ (.Y(_0257_),
    .A(\accumulator_object.bus[4] ));
 sg13g2_inv_1 _1020_ (.Y(_0258_),
    .A(net542));
 sg13g2_inv_1 _1021_ (.Y(_0259_),
    .A(net538));
 sg13g2_inv_4 _1022_ (.A(\accumulator_object.bus[1] ),
    .Y(_0260_));
 sg13g2_inv_1 _1023_ (.Y(_0261_),
    .A(net490));
 sg13g2_inv_1 _1024_ (.Y(_0262_),
    .A(net549));
 sg13g2_inv_1 _1025_ (.Y(_0263_),
    .A(net563));
 sg13g2_inv_1 _1026_ (.Y(_0264_),
    .A(net572));
 sg13g2_inv_1 _1027_ (.Y(_0265_),
    .A(net569));
 sg13g2_inv_1 _1028_ (.Y(_0266_),
    .A(net584));
 sg13g2_inv_1 _1029_ (.Y(_0267_),
    .A(net564));
 sg13g2_inv_1 _1030_ (.Y(_0268_),
    .A(net583));
 sg13g2_inv_1 _1031_ (.Y(_0269_),
    .A(net521));
 sg13g2_inv_1 _1032_ (.Y(_0270_),
    .A(net576));
 sg13g2_inv_2 _1033_ (.Y(_0271_),
    .A(net305));
 sg13g2_inv_1 _1034_ (.Y(_0272_),
    .A(_0019_));
 sg13g2_inv_1 _1035_ (.Y(_0273_),
    .A(Lp));
 sg13g2_inv_1 _1036_ (.Y(_0274_),
    .A(\ram.RAM[7][0] ));
 sg13g2_inv_1 _1037_ (.Y(_0275_),
    .A(net550));
 sg13g2_inv_1 _1038_ (.Y(_0276_),
    .A(net514));
 sg13g2_inv_1 _1039_ (.Y(_0277_),
    .A(net547));
 sg13g2_inv_1 _1040_ (.Y(_0278_),
    .A(net553));
 sg13g2_inv_1 _1041_ (.Y(_0279_),
    .A(net511));
 sg13g2_inv_1 _1042_ (.Y(_0280_),
    .A(net467));
 sg13g2_inv_1 _1601__2 (.Y(net233),
    .A(clknet_2_1__leaf_clk));
 sg13g2_nor2_2 _1044_ (.A(\cb.stage[1] ),
    .B(\cb.stage[0] ),
    .Y(_0281_));
 sg13g2_nor2b_1 _1045_ (.A(\cb.stage[1] ),
    .B_N(\cb.stage[2] ),
    .Y(_0282_));
 sg13g2_nand2_2 _1046_ (.Y(_0283_),
    .A(\cb.stage[2] ),
    .B(_0281_));
 sg13g2_nand2_2 _1047_ (.Y(_0284_),
    .A(\cb.stage[1] ),
    .B(\cb.stage[0] ));
 sg13g2_nor2_1 _1048_ (.A(\cb.stage[2] ),
    .B(_0284_),
    .Y(_0285_));
 sg13g2_or2_2 _1049_ (.X(_0286_),
    .B(_0284_),
    .A(\cb.stage[2] ));
 sg13g2_nand2_1 _1050_ (.Y(_0287_),
    .A(_0283_),
    .B(_0286_));
 sg13g2_nand3_1 _1051_ (.B(\instruction_register.instruction[6] ),
    .C(\instruction_register.instruction[4] ),
    .A(_0254_),
    .Y(_0288_));
 sg13g2_nor3_1 _1052_ (.A(net304),
    .B(_0286_),
    .C(_0288_),
    .Y(_0289_));
 sg13g2_nand2_1 _1053_ (.Y(_0065_),
    .A(_0256_),
    .B(_0289_));
 sg13g2_nor3_1 _1054_ (.A(\instruction_register.instruction[7] ),
    .B(_0255_),
    .C(\instruction_register.instruction[4] ),
    .Y(_0290_));
 sg13g2_and2_1 _1055_ (.A(\instruction_register.instruction[5] ),
    .B(_0290_),
    .X(_0291_));
 sg13g2_nor2b_1 _1056_ (.A(net304),
    .B_N(_0291_),
    .Y(_0292_));
 sg13g2_nand2b_1 _1057_ (.Y(_0293_),
    .B(_0292_),
    .A_N(\cb.stage[1] ));
 sg13g2_a22oi_1 _1058_ (.Y(_0223_),
    .B1(_0065_),
    .B2(_0293_),
    .A2(_0286_),
    .A1(_0283_));
 sg13g2_and2_1 _1059_ (.A(\cb.stage[0] ),
    .B(_0282_),
    .X(_0294_));
 sg13g2_nand2_1 _1060_ (.Y(_0295_),
    .A(\cb.stage[0] ),
    .B(_0282_));
 sg13g2_nand3_1 _1061_ (.B(_0255_),
    .C(\instruction_register.instruction[5] ),
    .A(_0254_),
    .Y(_0296_));
 sg13g2_nor3_1 _1062_ (.A(net304),
    .B(_0295_),
    .C(_0296_),
    .Y(_0087_));
 sg13g2_and2_1 _1063_ (.A(_0256_),
    .B(_0290_),
    .X(_0297_));
 sg13g2_nor2_1 _1064_ (.A(net304),
    .B(_0283_),
    .Y(_0298_));
 sg13g2_a21oi_1 _1065_ (.A1(_0297_),
    .A2(_0298_),
    .Y(_0222_),
    .B1(_0087_));
 sg13g2_and3_1 _1066_ (.X(_0086_),
    .A(net304),
    .B(\cb.stage[2] ),
    .C(_0281_));
 sg13g2_a21oi_1 _1067_ (.A1(_0292_),
    .A2(_0294_),
    .Y(_0221_),
    .B1(_0086_));
 sg13g2_nor2b_1 _1068_ (.A(\cb.stage[0] ),
    .B_N(\cb.stage[1] ),
    .Y(_0299_));
 sg13g2_nand2_1 _1069_ (.Y(_0300_),
    .A(_0018_),
    .B(_0299_));
 sg13g2_or2_1 _1070_ (.X(_0055_),
    .B(_0300_),
    .A(net304));
 sg13g2_nor2_1 _1071_ (.A(_0283_),
    .B(_0297_),
    .Y(_0301_));
 sg13g2_a221oi_1 _1072_ (.B2(_0296_),
    .C1(net9),
    .B1(_0301_),
    .A1(_0283_),
    .Y(_0302_),
    .A2(_0300_));
 sg13g2_inv_1 _1073_ (.Y(_0220_),
    .A(_0302_));
 sg13g2_and2_1 _1074_ (.A(net9),
    .B(_0285_),
    .X(_0085_));
 sg13g2_a21oi_1 _1075_ (.A1(_0291_),
    .A2(_0298_),
    .Y(_0219_),
    .B1(_0085_));
 sg13g2_nor2b_1 _1076_ (.A(_0290_),
    .B_N(_0296_),
    .Y(_0303_));
 sg13g2_nor3_1 _1077_ (.A(net304),
    .B(_0286_),
    .C(_0303_),
    .Y(_0304_));
 sg13g2_and2_1 _1078_ (.A(_0018_),
    .B(_0281_),
    .X(_0235_));
 sg13g2_nor2_1 _1079_ (.A(_0304_),
    .B(_0235_),
    .Y(_0218_));
 sg13g2_and2_1 _1080_ (.A(\instruction_register.instruction[4] ),
    .B(_0087_),
    .X(_0088_));
 sg13g2_and2_1 _1081_ (.A(\instruction_register.instruction[5] ),
    .B(_0289_),
    .X(_0067_));
 sg13g2_nor2_1 _1082_ (.A(_0304_),
    .B(_0067_),
    .Y(_0066_));
 sg13g2_or3_1 _1083_ (.A(net304),
    .B(_0283_),
    .C(_0296_),
    .X(_0056_));
 sg13g2_nand2b_2 _1084_ (.Y(_0581_),
    .B(net309),
    .A_N(\cb.control_signals[9] ));
 sg13g2_nand2b_2 _1085_ (.Y(_0577_),
    .B(net308),
    .A_N(\cb.control_signals[6] ));
 sg13g2_nand2_2 _1086_ (.Y(_0569_),
    .A(net309),
    .B(\cb.control_signals[4] ));
 sg13g2_nand2_2 _1087_ (.Y(_0561_),
    .A(net312),
    .B(net249));
 sg13g2_nand2_2 _1088_ (.Y(_0590_),
    .A(net311),
    .B(net251));
 sg13g2_nand2_2 _1089_ (.Y(_0557_),
    .A(net305),
    .B(\cb.control_signals[13] ));
 sg13g2_and4_2 _1090_ (.A(_0577_),
    .B(_0569_),
    .C(_0561_),
    .D(_0557_),
    .X(_0305_));
 sg13g2_nand3b_1 _1091_ (.B(net244),
    .C(_0305_),
    .Y(_0598_),
    .A_N(net250));
 sg13g2_xor2_1 _1092_ (.B(\alu_object.addsub.op_b[0] ),
    .A(\alu_object.addsub.genblk1[0].fa.a ),
    .X(\alu_object.addsub.genblk1[0].fa.sum ));
 sg13g2_mux2_1 _1093_ (.A0(\alu_object.addsub.genblk1[0].fa.cin ),
    .A1(\alu_object.addsub.genblk1[0].fa.a ),
    .S(\alu_object.addsub.op_b[0] ),
    .X(_0306_));
 sg13g2_xor2_1 _1094_ (.B(\alu_object.addsub.op_b[1] ),
    .A(\alu_object.addsub.genblk1[0].fa.cin ),
    .X(_0307_));
 sg13g2_nand2_1 _1095_ (.Y(_0308_),
    .A(_0272_),
    .B(_0307_));
 sg13g2_xnor2_1 _1096_ (.Y(_0309_),
    .A(_0272_),
    .B(_0307_));
 sg13g2_xnor2_1 _1097_ (.Y(\alu_object.addsub.genblk1[1].fa.sum ),
    .A(_0306_),
    .B(_0309_));
 sg13g2_xor2_1 _1098_ (.B(\alu_object.addsub.op_b[2] ),
    .A(\alu_object.addsub.genblk1[0].fa.cin ),
    .X(_0310_));
 sg13g2_nor2_1 _1099_ (.A(\alu_object.addsub.genblk1[2].fa.a ),
    .B(_0310_),
    .Y(_0311_));
 sg13g2_xnor2_1 _1100_ (.Y(_0312_),
    .A(\alu_object.addsub.genblk1[2].fa.a ),
    .B(_0310_));
 sg13g2_o21ai_1 _1101_ (.B1(_0306_),
    .Y(_0313_),
    .A1(_0272_),
    .A2(_0307_));
 sg13g2_nand2_1 _1102_ (.Y(_0314_),
    .A(_0308_),
    .B(_0313_));
 sg13g2_xnor2_1 _1103_ (.Y(\alu_object.addsub.genblk1[2].fa.sum ),
    .A(_0312_),
    .B(_0314_));
 sg13g2_xor2_1 _1104_ (.B(\alu_object.addsub.op_b[3] ),
    .A(\alu_object.addsub.genblk1[0].fa.cin ),
    .X(_0315_));
 sg13g2_and2_1 _1105_ (.A(\alu_object.addsub.genblk1[3].fa.a ),
    .B(_0315_),
    .X(_0316_));
 sg13g2_or2_1 _1106_ (.X(_0317_),
    .B(_0315_),
    .A(\alu_object.addsub.genblk1[3].fa.a ));
 sg13g2_nand2b_1 _1107_ (.Y(_0318_),
    .B(_0317_),
    .A_N(_0316_));
 sg13g2_a21oi_1 _1108_ (.A1(_0308_),
    .A2(_0313_),
    .Y(_0319_),
    .B1(_0311_));
 sg13g2_a21o_1 _1109_ (.A2(_0310_),
    .A1(\alu_object.addsub.genblk1[2].fa.a ),
    .B1(_0319_),
    .X(_0320_));
 sg13g2_xnor2_1 _1110_ (.Y(\alu_object.addsub.genblk1[3].fa.sum ),
    .A(_0318_),
    .B(_0320_));
 sg13g2_xor2_1 _1111_ (.B(\alu_object.addsub.op_b[4] ),
    .A(\alu_object.addsub.genblk1[0].fa.cin ),
    .X(_0321_));
 sg13g2_nor2_1 _1112_ (.A(\alu_object.addsub.genblk1[4].fa.a ),
    .B(_0321_),
    .Y(_0322_));
 sg13g2_xnor2_1 _1113_ (.Y(_0323_),
    .A(_0266_),
    .B(_0321_));
 sg13g2_a21oi_1 _1114_ (.A1(_0317_),
    .A2(_0320_),
    .Y(_0324_),
    .B1(_0316_));
 sg13g2_xnor2_1 _1115_ (.Y(\alu_object.addsub.genblk1[4].fa.sum ),
    .A(_0323_),
    .B(_0324_));
 sg13g2_xor2_1 _1116_ (.B(\alu_object.addsub.op_b[5] ),
    .A(\alu_object.addsub.genblk1[0].fa.cin ),
    .X(_0325_));
 sg13g2_nor2_1 _1117_ (.A(\alu_object.addsub.genblk1[5].fa.a ),
    .B(_0325_),
    .Y(_0326_));
 sg13g2_nand2_1 _1118_ (.Y(_0327_),
    .A(\alu_object.addsub.genblk1[5].fa.a ),
    .B(_0325_));
 sg13g2_nand2b_1 _1119_ (.Y(_0328_),
    .B(_0327_),
    .A_N(_0326_));
 sg13g2_a221oi_1 _1120_ (.B2(\alu_object.addsub.genblk1[4].fa.a ),
    .C1(_0316_),
    .B1(_0321_),
    .A1(_0317_),
    .Y(_0329_),
    .A2(_0320_));
 sg13g2_nor2_1 _1121_ (.A(_0322_),
    .B(_0329_),
    .Y(_0330_));
 sg13g2_xnor2_1 _1122_ (.Y(\alu_object.addsub.genblk1[5].fa.sum ),
    .A(_0328_),
    .B(_0330_));
 sg13g2_xor2_1 _1123_ (.B(\alu_object.addsub.op_b[6] ),
    .A(\alu_object.addsub.genblk1[0].fa.cin ),
    .X(_0331_));
 sg13g2_or2_1 _1124_ (.X(_0332_),
    .B(_0331_),
    .A(\alu_object.addsub.genblk1[6].fa.a ));
 sg13g2_nand2_1 _1125_ (.Y(_0333_),
    .A(\alu_object.addsub.genblk1[6].fa.a ),
    .B(_0331_));
 sg13g2_nand2_1 _1126_ (.Y(_0334_),
    .A(_0332_),
    .B(_0333_));
 sg13g2_or3_1 _1127_ (.A(_0322_),
    .B(_0326_),
    .C(_0329_),
    .X(_0335_));
 sg13g2_and2_1 _1128_ (.A(_0327_),
    .B(_0335_),
    .X(_0336_));
 sg13g2_xnor2_1 _1129_ (.Y(_0337_),
    .A(_0334_),
    .B(_0336_));
 sg13g2_inv_1 _1130_ (.Y(\alu_object.addsub.genblk1[6].fa.sum ),
    .A(_0337_));
 sg13g2_xor2_1 _1131_ (.B(\alu_object.addsub.op_b[7] ),
    .A(\alu_object.addsub.genblk1[0].fa.cin ),
    .X(_0338_));
 sg13g2_nor2_1 _1132_ (.A(\alu_object.addsub.genblk1[7].fa.a ),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_and2_1 _1133_ (.A(\alu_object.addsub.genblk1[7].fa.a ),
    .B(_0338_),
    .X(_0340_));
 sg13g2_or2_1 _1134_ (.X(_0341_),
    .B(_0340_),
    .A(_0339_));
 sg13g2_nand3_1 _1135_ (.B(_0333_),
    .C(_0335_),
    .A(_0327_),
    .Y(_0342_));
 sg13g2_and2_1 _1136_ (.A(_0332_),
    .B(_0342_),
    .X(_0343_));
 sg13g2_nand3_1 _1137_ (.B(_0341_),
    .C(_0342_),
    .A(_0332_),
    .Y(_0344_));
 sg13g2_a21o_1 _1138_ (.A2(_0342_),
    .A1(_0332_),
    .B1(_0341_),
    .X(_0345_));
 sg13g2_nand2_1 _1139_ (.Y(\alu_object.addsub.genblk1[7].fa.sum ),
    .A(_0344_),
    .B(_0345_));
 sg13g2_nand2_1 _1140_ (.Y(_0346_),
    .A(\cb.stage[0] ),
    .B(_0018_));
 sg13g2_nor2_1 _1141_ (.A(\cb.stage[1] ),
    .B(_0346_),
    .Y(_0008_));
 sg13g2_mux2_1 _1142_ (.A0(\ram.RAM[14][0] ),
    .A1(\ram.RAM[15][0] ),
    .S(net301),
    .X(_0347_));
 sg13g2_nor2b_1 _1143_ (.A(net299),
    .B_N(\ram.RAM[12][0] ),
    .Y(_0348_));
 sg13g2_a21oi_1 _1144_ (.A1(net298),
    .A2(\ram.RAM[13][0] ),
    .Y(_0349_),
    .B1(_0348_));
 sg13g2_o21ai_1 _1145_ (.B1(net281),
    .Y(_0350_),
    .A1(net287),
    .A2(_0349_));
 sg13g2_a21oi_1 _1146_ (.A1(net288),
    .A2(_0347_),
    .Y(_0351_),
    .B1(_0350_));
 sg13g2_mux4_1 _1147_ (.S0(net293),
    .A0(\ram.RAM[8][0] ),
    .A1(\ram.RAM[9][0] ),
    .A2(\ram.RAM[10][0] ),
    .A3(\ram.RAM[11][0] ),
    .S1(net284),
    .X(_0352_));
 sg13g2_o21ai_1 _1148_ (.B1(net274),
    .Y(_0353_),
    .A1(net279),
    .A2(_0352_));
 sg13g2_or2_1 _1149_ (.X(_0354_),
    .B(_0353_),
    .A(_0351_));
 sg13g2_mux2_1 _1150_ (.A0(\ram.RAM[2][0] ),
    .A1(\ram.RAM[3][0] ),
    .S(net290),
    .X(_0355_));
 sg13g2_nor2b_1 _1151_ (.A(net290),
    .B_N(\ram.RAM[0][0] ),
    .Y(_0356_));
 sg13g2_a21oi_1 _1152_ (.A1(\ram.RAM[1][0] ),
    .A2(net290),
    .Y(_0357_),
    .B1(_0356_));
 sg13g2_a21oi_1 _1153_ (.A1(net282),
    .A2(_0355_),
    .Y(_0358_),
    .B1(net277));
 sg13g2_o21ai_1 _1154_ (.B1(_0358_),
    .Y(_0359_),
    .A1(net282),
    .A2(_0357_));
 sg13g2_o21ai_1 _1155_ (.B1(net286),
    .Y(_0360_),
    .A1(net295),
    .A2(\ram.RAM[6][0] ));
 sg13g2_a21oi_1 _1156_ (.A1(net297),
    .A2(_0274_),
    .Y(_0361_),
    .B1(_0360_));
 sg13g2_nor2b_1 _1157_ (.A(net297),
    .B_N(\ram.RAM[4][0] ),
    .Y(_0362_));
 sg13g2_a21oi_1 _1158_ (.A1(net298),
    .A2(\ram.RAM[5][0] ),
    .Y(_0363_),
    .B1(_0362_));
 sg13g2_o21ai_1 _1159_ (.B1(net280),
    .Y(_0364_),
    .A1(net286),
    .A2(_0363_));
 sg13g2_o21ai_1 _1160_ (.B1(_0359_),
    .Y(_0365_),
    .A1(_0361_),
    .A2(_0364_));
 sg13g2_o21ai_1 _1161_ (.B1(_0354_),
    .Y(_0010_),
    .A1(net275),
    .A2(_0365_));
 sg13g2_mux4_1 _1162_ (.S0(net293),
    .A0(\ram.RAM[8][1] ),
    .A1(\ram.RAM[9][1] ),
    .A2(\ram.RAM[10][1] ),
    .A3(\ram.RAM[11][1] ),
    .S1(net284),
    .X(_0366_));
 sg13g2_nor2_1 _1163_ (.A(net278),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_nor2b_1 _1164_ (.A(net300),
    .B_N(\ram.RAM[12][1] ),
    .Y(_0368_));
 sg13g2_a21oi_1 _1165_ (.A1(net300),
    .A2(\ram.RAM[13][1] ),
    .Y(_0369_),
    .B1(_0368_));
 sg13g2_o21ai_1 _1166_ (.B1(net289),
    .Y(_0370_),
    .A1(net300),
    .A2(\ram.RAM[14][1] ));
 sg13g2_a21oi_1 _1167_ (.A1(net300),
    .A2(_0275_),
    .Y(_0371_),
    .B1(_0370_));
 sg13g2_o21ai_1 _1168_ (.B1(net278),
    .Y(_0372_),
    .A1(net289),
    .A2(_0369_));
 sg13g2_o21ai_1 _1169_ (.B1(net274),
    .Y(_0373_),
    .A1(_0371_),
    .A2(_0372_));
 sg13g2_nor2b_1 _1170_ (.A(net296),
    .B_N(\ram.RAM[4][1] ),
    .Y(_0374_));
 sg13g2_a21oi_1 _1171_ (.A1(net296),
    .A2(\ram.RAM[5][1] ),
    .Y(_0375_),
    .B1(_0374_));
 sg13g2_mux2_1 _1172_ (.A0(\ram.RAM[6][1] ),
    .A1(\ram.RAM[7][1] ),
    .S(net296),
    .X(_0376_));
 sg13g2_o21ai_1 _1173_ (.B1(net280),
    .Y(_0377_),
    .A1(net287),
    .A2(_0375_));
 sg13g2_a21oi_1 _1174_ (.A1(net287),
    .A2(_0376_),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_mux4_1 _1175_ (.S0(net291),
    .A0(\ram.RAM[0][1] ),
    .A1(\ram.RAM[1][1] ),
    .A2(\ram.RAM[2][1] ),
    .A3(\ram.RAM[3][1] ),
    .S1(net283),
    .X(_0379_));
 sg13g2_nor2_1 _1176_ (.A(net276),
    .B(_0378_),
    .Y(_0380_));
 sg13g2_o21ai_1 _1177_ (.B1(_0380_),
    .Y(_0381_),
    .A1(net277),
    .A2(_0379_));
 sg13g2_o21ai_1 _1178_ (.B1(_0381_),
    .Y(_0011_),
    .A1(_0367_),
    .A2(_0373_));
 sg13g2_mux4_1 _1179_ (.S0(net293),
    .A0(\ram.RAM[8][2] ),
    .A1(\ram.RAM[9][2] ),
    .A2(\ram.RAM[10][2] ),
    .A3(\ram.RAM[11][2] ),
    .S1(net284),
    .X(_0382_));
 sg13g2_nor2_1 _1180_ (.A(net279),
    .B(_0382_),
    .Y(_0383_));
 sg13g2_nor2b_1 _1181_ (.A(net298),
    .B_N(\ram.RAM[12][2] ),
    .Y(_0384_));
 sg13g2_a21oi_1 _1182_ (.A1(net301),
    .A2(\ram.RAM[13][2] ),
    .Y(_0385_),
    .B1(_0384_));
 sg13g2_o21ai_1 _1183_ (.B1(net288),
    .Y(_0386_),
    .A1(net301),
    .A2(\ram.RAM[14][2] ));
 sg13g2_a21oi_1 _1184_ (.A1(net301),
    .A2(_0276_),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_o21ai_1 _1185_ (.B1(net279),
    .Y(_0388_),
    .A1(net288),
    .A2(_0385_));
 sg13g2_o21ai_1 _1186_ (.B1(net275),
    .Y(_0389_),
    .A1(_0387_),
    .A2(_0388_));
 sg13g2_nor2b_1 _1187_ (.A(net297),
    .B_N(\ram.RAM[4][2] ),
    .Y(_0390_));
 sg13g2_a21oi_1 _1188_ (.A1(net297),
    .A2(\ram.RAM[5][2] ),
    .Y(_0391_),
    .B1(_0390_));
 sg13g2_mux2_1 _1189_ (.A0(\ram.RAM[6][2] ),
    .A1(\ram.RAM[7][2] ),
    .S(net297),
    .X(_0392_));
 sg13g2_o21ai_1 _1190_ (.B1(net280),
    .Y(_0393_),
    .A1(net286),
    .A2(_0391_));
 sg13g2_a21oi_1 _1191_ (.A1(net286),
    .A2(_0392_),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_mux4_1 _1192_ (.S0(net291),
    .A0(\ram.RAM[0][2] ),
    .A1(\ram.RAM[1][2] ),
    .A2(\ram.RAM[2][2] ),
    .A3(\ram.RAM[3][2] ),
    .S1(net283),
    .X(_0395_));
 sg13g2_nor2_1 _1193_ (.A(net276),
    .B(_0394_),
    .Y(_0396_));
 sg13g2_o21ai_1 _1194_ (.B1(_0396_),
    .Y(_0397_),
    .A1(net280),
    .A2(_0395_));
 sg13g2_o21ai_1 _1195_ (.B1(_0397_),
    .Y(_0012_),
    .A1(_0383_),
    .A2(_0389_));
 sg13g2_mux4_1 _1196_ (.S0(net293),
    .A0(\ram.RAM[8][3] ),
    .A1(\ram.RAM[9][3] ),
    .A2(\ram.RAM[10][3] ),
    .A3(\ram.RAM[11][3] ),
    .S1(net284),
    .X(_0398_));
 sg13g2_nor2_1 _1197_ (.A(net278),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_nor2b_1 _1198_ (.A(net300),
    .B_N(\ram.RAM[12][3] ),
    .Y(_0400_));
 sg13g2_a21oi_1 _1199_ (.A1(net300),
    .A2(\ram.RAM[13][3] ),
    .Y(_0401_),
    .B1(_0400_));
 sg13g2_o21ai_1 _1200_ (.B1(net284),
    .Y(_0402_),
    .A1(net294),
    .A2(\ram.RAM[14][3] ));
 sg13g2_a21oi_1 _1201_ (.A1(net294),
    .A2(_0277_),
    .Y(_0403_),
    .B1(_0402_));
 sg13g2_o21ai_1 _1202_ (.B1(net278),
    .Y(_0404_),
    .A1(net284),
    .A2(_0401_));
 sg13g2_o21ai_1 _1203_ (.B1(net274),
    .Y(_0405_),
    .A1(_0403_),
    .A2(_0404_));
 sg13g2_mux4_1 _1204_ (.S0(net291),
    .A0(\ram.RAM[0][3] ),
    .A1(\ram.RAM[1][3] ),
    .A2(\ram.RAM[2][3] ),
    .A3(\ram.RAM[3][3] ),
    .S1(net283),
    .X(_0406_));
 sg13g2_mux2_1 _1205_ (.A0(\ram.RAM[6][3] ),
    .A1(\ram.RAM[7][3] ),
    .S(net295),
    .X(_0407_));
 sg13g2_nor2b_1 _1206_ (.A(net295),
    .B_N(\ram.RAM[4][3] ),
    .Y(_0408_));
 sg13g2_a21oi_1 _1207_ (.A1(net295),
    .A2(\ram.RAM[5][3] ),
    .Y(_0409_),
    .B1(_0408_));
 sg13g2_o21ai_1 _1208_ (.B1(net277),
    .Y(_0410_),
    .A1(net287),
    .A2(_0409_));
 sg13g2_a21oi_1 _1209_ (.A1(net287),
    .A2(_0407_),
    .Y(_0411_),
    .B1(_0410_));
 sg13g2_nor2_1 _1210_ (.A(net276),
    .B(_0411_),
    .Y(_0412_));
 sg13g2_o21ai_1 _1211_ (.B1(_0412_),
    .Y(_0413_),
    .A1(net277),
    .A2(_0406_));
 sg13g2_o21ai_1 _1212_ (.B1(_0413_),
    .Y(_0013_),
    .A1(_0399_),
    .A2(_0405_));
 sg13g2_mux4_1 _1213_ (.S0(net293),
    .A0(\ram.RAM[8][4] ),
    .A1(\ram.RAM[9][4] ),
    .A2(\ram.RAM[10][4] ),
    .A3(\ram.RAM[11][4] ),
    .S1(net284),
    .X(_0414_));
 sg13g2_nor2b_1 _1214_ (.A(net300),
    .B_N(\ram.RAM[12][4] ),
    .Y(_0415_));
 sg13g2_a21oi_1 _1215_ (.A1(net300),
    .A2(\ram.RAM[13][4] ),
    .Y(_0416_),
    .B1(_0415_));
 sg13g2_mux2_1 _1216_ (.A0(\ram.RAM[14][4] ),
    .A1(\ram.RAM[15][4] ),
    .S(net303),
    .X(_0417_));
 sg13g2_o21ai_1 _1217_ (.B1(net279),
    .Y(_0418_),
    .A1(net289),
    .A2(_0416_));
 sg13g2_a21oi_1 _1218_ (.A1(net289),
    .A2(_0417_),
    .Y(_0419_),
    .B1(_0418_));
 sg13g2_nor2b_1 _1219_ (.A(_0419_),
    .B_N(net274),
    .Y(_0420_));
 sg13g2_o21ai_1 _1220_ (.B1(_0420_),
    .Y(_0421_),
    .A1(net278),
    .A2(_0414_));
 sg13g2_nor2b_1 _1221_ (.A(net296),
    .B_N(\ram.RAM[4][4] ),
    .Y(_0422_));
 sg13g2_a21oi_1 _1222_ (.A1(net296),
    .A2(\ram.RAM[5][4] ),
    .Y(_0423_),
    .B1(_0422_));
 sg13g2_nor2b_1 _1223_ (.A(net296),
    .B_N(\ram.RAM[6][4] ),
    .Y(_0424_));
 sg13g2_a21oi_1 _1224_ (.A1(net296),
    .A2(\ram.RAM[7][4] ),
    .Y(_0425_),
    .B1(_0424_));
 sg13g2_nor2b_1 _1225_ (.A(net292),
    .B_N(\ram.RAM[2][4] ),
    .Y(_0426_));
 sg13g2_a21oi_1 _1226_ (.A1(net292),
    .A2(\ram.RAM[3][4] ),
    .Y(_0427_),
    .B1(_0426_));
 sg13g2_nor2b_1 _1227_ (.A(net291),
    .B_N(\ram.RAM[0][4] ),
    .Y(_0428_));
 sg13g2_a21oi_1 _1228_ (.A1(net291),
    .A2(\ram.RAM[1][4] ),
    .Y(_0429_),
    .B1(_0428_));
 sg13g2_mux4_1 _1229_ (.S0(net282),
    .A0(_0429_),
    .A1(_0427_),
    .A2(_0423_),
    .A3(_0425_),
    .S1(net277),
    .X(_0430_));
 sg13g2_o21ai_1 _1230_ (.B1(_0421_),
    .Y(_0014_),
    .A1(net274),
    .A2(_0430_));
 sg13g2_mux4_1 _1231_ (.S0(net293),
    .A0(\ram.RAM[8][5] ),
    .A1(\ram.RAM[9][5] ),
    .A2(\ram.RAM[10][5] ),
    .A3(\ram.RAM[11][5] ),
    .S1(net285),
    .X(_0431_));
 sg13g2_nor2b_1 _1232_ (.A(net301),
    .B_N(\ram.RAM[12][5] ),
    .Y(_0432_));
 sg13g2_a21oi_1 _1233_ (.A1(net301),
    .A2(\ram.RAM[13][5] ),
    .Y(_0433_),
    .B1(_0432_));
 sg13g2_mux2_1 _1234_ (.A0(\ram.RAM[14][5] ),
    .A1(\ram.RAM[15][5] ),
    .S(net302),
    .X(_0434_));
 sg13g2_o21ai_1 _1235_ (.B1(net281),
    .Y(_0435_),
    .A1(net288),
    .A2(_0433_));
 sg13g2_a21oi_1 _1236_ (.A1(net289),
    .A2(_0434_),
    .Y(_0436_),
    .B1(_0435_));
 sg13g2_nor2b_1 _1237_ (.A(_0436_),
    .B_N(net275),
    .Y(_0437_));
 sg13g2_o21ai_1 _1238_ (.B1(_0437_),
    .Y(_0438_),
    .A1(net279),
    .A2(_0431_));
 sg13g2_mux2_1 _1239_ (.A0(\ram.RAM[2][5] ),
    .A1(\ram.RAM[3][5] ),
    .S(net290),
    .X(_0439_));
 sg13g2_nor2b_1 _1240_ (.A(net290),
    .B_N(\ram.RAM[0][5] ),
    .Y(_0440_));
 sg13g2_a21oi_1 _1241_ (.A1(net290),
    .A2(\ram.RAM[1][5] ),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_a21oi_1 _1242_ (.A1(net282),
    .A2(_0439_),
    .Y(_0442_),
    .B1(net277));
 sg13g2_o21ai_1 _1243_ (.B1(_0442_),
    .Y(_0443_),
    .A1(net282),
    .A2(_0441_));
 sg13g2_o21ai_1 _1244_ (.B1(net287),
    .Y(_0444_),
    .A1(net295),
    .A2(\ram.RAM[6][5] ));
 sg13g2_a21oi_1 _1245_ (.A1(net295),
    .A2(_0278_),
    .Y(_0445_),
    .B1(_0444_));
 sg13g2_nor2b_1 _1246_ (.A(net297),
    .B_N(\ram.RAM[4][5] ),
    .Y(_0446_));
 sg13g2_a21oi_1 _1247_ (.A1(net298),
    .A2(\ram.RAM[5][5] ),
    .Y(_0447_),
    .B1(_0446_));
 sg13g2_o21ai_1 _1248_ (.B1(net280),
    .Y(_0448_),
    .A1(net286),
    .A2(_0447_));
 sg13g2_o21ai_1 _1249_ (.B1(_0443_),
    .Y(_0449_),
    .A1(_0445_),
    .A2(_0448_));
 sg13g2_o21ai_1 _1250_ (.B1(_0438_),
    .Y(_0015_),
    .A1(net275),
    .A2(_0449_));
 sg13g2_mux4_1 _1251_ (.S0(net293),
    .A0(\ram.RAM[8][6] ),
    .A1(\ram.RAM[9][6] ),
    .A2(\ram.RAM[10][6] ),
    .A3(\ram.RAM[11][6] ),
    .S1(net285),
    .X(_0450_));
 sg13g2_nor2b_1 _1252_ (.A(net301),
    .B_N(\ram.RAM[12][6] ),
    .Y(_0451_));
 sg13g2_a21oi_1 _1253_ (.A1(net302),
    .A2(\ram.RAM[13][6] ),
    .Y(_0452_),
    .B1(_0451_));
 sg13g2_mux2_1 _1254_ (.A0(\ram.RAM[14][6] ),
    .A1(\ram.RAM[15][6] ),
    .S(net302),
    .X(_0453_));
 sg13g2_o21ai_1 _1255_ (.B1(net279),
    .Y(_0454_),
    .A1(net288),
    .A2(_0452_));
 sg13g2_a21oi_1 _1256_ (.A1(net288),
    .A2(_0453_),
    .Y(_0455_),
    .B1(_0454_));
 sg13g2_nor2b_1 _1257_ (.A(_0455_),
    .B_N(net275),
    .Y(_0456_));
 sg13g2_o21ai_1 _1258_ (.B1(_0456_),
    .Y(_0457_),
    .A1(net279),
    .A2(_0450_));
 sg13g2_mux2_1 _1259_ (.A0(\ram.RAM[2][6] ),
    .A1(\ram.RAM[3][6] ),
    .S(net292),
    .X(_0458_));
 sg13g2_nor2b_1 _1260_ (.A(net290),
    .B_N(\ram.RAM[0][6] ),
    .Y(_0459_));
 sg13g2_a21oi_1 _1261_ (.A1(net290),
    .A2(\ram.RAM[1][6] ),
    .Y(_0460_),
    .B1(_0459_));
 sg13g2_a21oi_1 _1262_ (.A1(net282),
    .A2(_0458_),
    .Y(_0461_),
    .B1(net277));
 sg13g2_o21ai_1 _1263_ (.B1(_0461_),
    .Y(_0462_),
    .A1(net283),
    .A2(_0460_));
 sg13g2_o21ai_1 _1264_ (.B1(net286),
    .Y(_0463_),
    .A1(net299),
    .A2(\ram.RAM[6][6] ));
 sg13g2_a21oi_1 _1265_ (.A1(net298),
    .A2(_0279_),
    .Y(_0464_),
    .B1(_0463_));
 sg13g2_nor2b_1 _1266_ (.A(net298),
    .B_N(\ram.RAM[4][6] ),
    .Y(_0465_));
 sg13g2_a21oi_1 _1267_ (.A1(net298),
    .A2(\ram.RAM[5][6] ),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_o21ai_1 _1268_ (.B1(net280),
    .Y(_0467_),
    .A1(net286),
    .A2(_0466_));
 sg13g2_o21ai_1 _1269_ (.B1(_0462_),
    .Y(_0468_),
    .A1(_0464_),
    .A2(_0467_));
 sg13g2_o21ai_1 _1270_ (.B1(_0457_),
    .Y(_0016_),
    .A1(net274),
    .A2(_0468_));
 sg13g2_mux4_1 _1271_ (.S0(net293),
    .A0(\ram.RAM[8][7] ),
    .A1(\ram.RAM[9][7] ),
    .A2(\ram.RAM[10][7] ),
    .A3(\ram.RAM[11][7] ),
    .S1(net284),
    .X(_0469_));
 sg13g2_nor2b_1 _1272_ (.A(net302),
    .B_N(\ram.RAM[12][7] ),
    .Y(_0470_));
 sg13g2_a21oi_1 _1273_ (.A1(net301),
    .A2(\ram.RAM[13][7] ),
    .Y(_0471_),
    .B1(_0470_));
 sg13g2_mux2_1 _1274_ (.A0(\ram.RAM[14][7] ),
    .A1(\ram.RAM[15][7] ),
    .S(net302),
    .X(_0472_));
 sg13g2_o21ai_1 _1275_ (.B1(net279),
    .Y(_0473_),
    .A1(net288),
    .A2(_0471_));
 sg13g2_a21oi_1 _1276_ (.A1(net288),
    .A2(_0472_),
    .Y(_0474_),
    .B1(_0473_));
 sg13g2_nor2b_1 _1277_ (.A(_0474_),
    .B_N(net274),
    .Y(_0475_));
 sg13g2_o21ai_1 _1278_ (.B1(_0475_),
    .Y(_0476_),
    .A1(net278),
    .A2(_0469_));
 sg13g2_mux2_1 _1279_ (.A0(\ram.RAM[2][7] ),
    .A1(\ram.RAM[3][7] ),
    .S(net291),
    .X(_0477_));
 sg13g2_nor2b_1 _1280_ (.A(net291),
    .B_N(\ram.RAM[0][7] ),
    .Y(_0478_));
 sg13g2_a21oi_1 _1281_ (.A1(net291),
    .A2(\ram.RAM[1][7] ),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_a21oi_1 _1282_ (.A1(net282),
    .A2(_0477_),
    .Y(_0480_),
    .B1(net277));
 sg13g2_o21ai_1 _1283_ (.B1(_0480_),
    .Y(_0481_),
    .A1(net282),
    .A2(_0479_));
 sg13g2_o21ai_1 _1284_ (.B1(net287),
    .Y(_0482_),
    .A1(net295),
    .A2(\ram.RAM[6][7] ));
 sg13g2_a21oi_1 _1285_ (.A1(net295),
    .A2(_0280_),
    .Y(_0483_),
    .B1(_0482_));
 sg13g2_nor2b_1 _1286_ (.A(net297),
    .B_N(\ram.RAM[4][7] ),
    .Y(_0484_));
 sg13g2_a21oi_1 _1287_ (.A1(net297),
    .A2(\ram.RAM[5][7] ),
    .Y(_0485_),
    .B1(_0484_));
 sg13g2_o21ai_1 _1288_ (.B1(net280),
    .Y(_0486_),
    .A1(net286),
    .A2(_0485_));
 sg13g2_o21ai_1 _1289_ (.B1(_0481_),
    .Y(_0487_),
    .A1(_0483_),
    .A2(_0486_));
 sg13g2_o21ai_1 _1290_ (.B1(_0476_),
    .Y(_0017_),
    .A1(net274),
    .A2(_0487_));
 sg13g2_nor4_2 _1291_ (.A(\instruction_register.instruction[7] ),
    .B(\instruction_register.instruction[6] ),
    .C(\instruction_register.instruction[5] ),
    .Y(_0488_),
    .D(\instruction_register.instruction[4] ));
 sg13g2_a22oi_1 _1292_ (.Y(_0489_),
    .B1(_0285_),
    .B2(_0488_),
    .A2(net306),
    .A1(net557));
 sg13g2_inv_1 _1293_ (.Y(_0009_),
    .A(_0489_));
 sg13g2_mux2_1 _1294_ (.A0(\accumulator_object.bus[0] ),
    .A1(net579),
    .S(\cb.control_signals[11] ),
    .X(_0004_));
 sg13g2_nand2_1 _1295_ (.Y(_0490_),
    .A(net248),
    .B(net581));
 sg13g2_o21ai_1 _1296_ (.B1(_0490_),
    .Y(_0005_),
    .A1(_0260_),
    .A2(net248));
 sg13g2_mux2_1 _1297_ (.A0(net241),
    .A1(net556),
    .S(net248),
    .X(_0006_));
 sg13g2_mux2_1 _1298_ (.A0(net240),
    .A1(net555),
    .S(net248),
    .X(_0007_));
 sg13g2_nor2b_1 _1299_ (.A(\input_mar_register.addr[0] ),
    .B_N(_0020_),
    .Y(_0491_));
 sg13g2_nand2b_2 _1300_ (.Y(_0492_),
    .B(_0491_),
    .A_N(\input_mar_register.addr[1] ));
 sg13g2_nand2b_2 _1301_ (.Y(_0493_),
    .B(net257),
    .A_N(net256));
 sg13g2_nor2_2 _1302_ (.A(_0492_),
    .B(_0493_),
    .Y(_0494_));
 sg13g2_mux2_1 _1303_ (.A0(net344),
    .A1(net272),
    .S(_0494_),
    .X(_0039_));
 sg13g2_mux2_1 _1304_ (.A0(net363),
    .A1(net270),
    .S(_0494_),
    .X(_0040_));
 sg13g2_mux2_1 _1305_ (.A0(net360),
    .A1(net268),
    .S(_0494_),
    .X(_0041_));
 sg13g2_mux2_1 _1306_ (.A0(net402),
    .A1(net266),
    .S(_0494_),
    .X(_0042_));
 sg13g2_mux2_1 _1307_ (.A0(net367),
    .A1(net264),
    .S(_0494_),
    .X(_0043_));
 sg13g2_mux2_1 _1308_ (.A0(net387),
    .A1(net262),
    .S(_0494_),
    .X(_0044_));
 sg13g2_mux2_1 _1309_ (.A0(net343),
    .A1(net260),
    .S(_0494_),
    .X(_0045_));
 sg13g2_mux2_1 _1310_ (.A0(net371),
    .A1(net258),
    .S(_0494_),
    .X(_0046_));
 sg13g2_mux2_1 _1311_ (.A0(\accumulator_object.bus[0] ),
    .A1(net573),
    .S(net252),
    .X(_0047_));
 sg13g2_nand2_1 _1312_ (.Y(_0495_),
    .A(\cb.control_signals[0] ),
    .B(net552));
 sg13g2_o21ai_1 _1313_ (.B1(_0495_),
    .Y(_0048_),
    .A1(_0260_),
    .A2(net252));
 sg13g2_mux2_1 _1314_ (.A0(\accumulator_object.bus[2] ),
    .A1(net567),
    .S(net252),
    .X(_0049_));
 sg13g2_mux2_1 _1315_ (.A0(\accumulator_object.bus[3] ),
    .A1(net562),
    .S(net252),
    .X(_0050_));
 sg13g2_nand2_1 _1316_ (.Y(_0496_),
    .A(net252),
    .B(net544));
 sg13g2_o21ai_1 _1317_ (.B1(_0496_),
    .Y(_0051_),
    .A1(_0257_),
    .A2(\cb.control_signals[0] ));
 sg13g2_mux2_1 _1318_ (.A0(\accumulator_object.bus[5] ),
    .A1(net574),
    .S(net252),
    .X(_0052_));
 sg13g2_mux2_1 _1319_ (.A0(\accumulator_object.bus[6] ),
    .A1(net575),
    .S(net252),
    .X(_0053_));
 sg13g2_mux2_1 _1320_ (.A0(\accumulator_object.bus[7] ),
    .A1(net577),
    .S(net252),
    .X(_0054_));
 sg13g2_nand3b_1 _1321_ (.B(_0020_),
    .C(\input_mar_register.addr[0] ),
    .Y(_0497_),
    .A_N(\input_mar_register.addr[1] ));
 sg13g2_nor3_2 _1322_ (.A(net257),
    .B(net256),
    .C(_0497_),
    .Y(_0498_));
 sg13g2_mux2_1 _1323_ (.A0(net375),
    .A1(net273),
    .S(_0498_),
    .X(_0057_));
 sg13g2_mux2_1 _1324_ (.A0(net451),
    .A1(net271),
    .S(_0498_),
    .X(_0058_));
 sg13g2_mux2_1 _1325_ (.A0(net472),
    .A1(net269),
    .S(_0498_),
    .X(_0059_));
 sg13g2_mux2_1 _1326_ (.A0(net444),
    .A1(net267),
    .S(_0498_),
    .X(_0060_));
 sg13g2_mux2_1 _1327_ (.A0(net480),
    .A1(net265),
    .S(_0498_),
    .X(_0061_));
 sg13g2_mux2_1 _1328_ (.A0(net483),
    .A1(net263),
    .S(_0498_),
    .X(_0062_));
 sg13g2_mux2_1 _1329_ (.A0(net491),
    .A1(net261),
    .S(_0498_),
    .X(_0063_));
 sg13g2_mux2_1 _1330_ (.A0(net394),
    .A1(net259),
    .S(_0498_),
    .X(_0064_));
 sg13g2_a21oi_1 _1331_ (.A1(net593),
    .A2(_0284_),
    .Y(_0499_),
    .B1(_0287_));
 sg13g2_nand2_1 _1332_ (.Y(_0500_),
    .A(net590),
    .B(_0299_));
 sg13g2_nor3_1 _1333_ (.A(\cb.stage[0] ),
    .B(_0271_),
    .C(_0499_),
    .Y(_0501_));
 sg13g2_a21o_1 _1334_ (.A2(net594),
    .A1(_0500_),
    .B1(HF),
    .X(_0068_));
 sg13g2_nand2_2 _1335_ (.Y(_0502_),
    .A(\input_mar_register.addr[1] ),
    .B(_0491_));
 sg13g2_nand2_2 _1336_ (.Y(_0503_),
    .A(net257),
    .B(net256));
 sg13g2_nor2_2 _1337_ (.A(_0502_),
    .B(_0503_),
    .Y(_0504_));
 sg13g2_mux2_1 _1338_ (.A0(net330),
    .A1(net272),
    .S(_0504_),
    .X(_0069_));
 sg13g2_mux2_1 _1339_ (.A0(net530),
    .A1(\input_mar_register.data[1] ),
    .S(_0504_),
    .X(_0070_));
 sg13g2_mux2_1 _1340_ (.A0(net482),
    .A1(net268),
    .S(_0504_),
    .X(_0071_));
 sg13g2_mux2_1 _1341_ (.A0(net437),
    .A1(net266),
    .S(_0504_),
    .X(_0072_));
 sg13g2_mux2_1 _1342_ (.A0(net383),
    .A1(\input_mar_register.data[4] ),
    .S(_0504_),
    .X(_0073_));
 sg13g2_mux2_1 _1343_ (.A0(net332),
    .A1(net262),
    .S(_0504_),
    .X(_0074_));
 sg13g2_mux2_1 _1344_ (.A0(net352),
    .A1(net260),
    .S(_0504_),
    .X(_0075_));
 sg13g2_mux2_1 _1345_ (.A0(net340),
    .A1(net258),
    .S(_0504_),
    .X(_0076_));
 sg13g2_nand3_1 _1346_ (.B(\input_mar_register.addr[1] ),
    .C(_0020_),
    .A(\input_mar_register.addr[0] ),
    .Y(_0505_));
 sg13g2_nor2_2 _1347_ (.A(_0503_),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_mux2_1 _1348_ (.A0(net545),
    .A1(net272),
    .S(net243),
    .X(_0077_));
 sg13g2_nand2_1 _1349_ (.Y(_0507_),
    .A(net270),
    .B(net243));
 sg13g2_o21ai_1 _1350_ (.B1(_0507_),
    .Y(_0078_),
    .A1(_0275_),
    .A2(net243));
 sg13g2_nand2_1 _1351_ (.Y(_0508_),
    .A(net268),
    .B(_0506_));
 sg13g2_o21ai_1 _1352_ (.B1(_0508_),
    .Y(_0079_),
    .A1(_0276_),
    .A2(_0506_));
 sg13g2_nand2_1 _1353_ (.Y(_0509_),
    .A(net266),
    .B(net243));
 sg13g2_o21ai_1 _1354_ (.B1(_0509_),
    .Y(_0080_),
    .A1(_0277_),
    .A2(net243));
 sg13g2_mux2_1 _1355_ (.A0(net516),
    .A1(net264),
    .S(net243),
    .X(_0081_));
 sg13g2_mux2_1 _1356_ (.A0(net522),
    .A1(net262),
    .S(net243),
    .X(_0082_));
 sg13g2_mux2_1 _1357_ (.A0(net520),
    .A1(net260),
    .S(_0506_),
    .X(_0083_));
 sg13g2_mux2_1 _1358_ (.A0(net498),
    .A1(net258),
    .S(net243),
    .X(_0084_));
 sg13g2_mux2_1 _1359_ (.A0(\accumulator_object.bus[0] ),
    .A1(net578),
    .S(net253),
    .X(_0089_));
 sg13g2_nand2_1 _1360_ (.Y(_0510_),
    .A(net417),
    .B(net253));
 sg13g2_o21ai_1 _1361_ (.B1(_0510_),
    .Y(_0090_),
    .A1(_0260_),
    .A2(net253));
 sg13g2_mux2_1 _1362_ (.A0(net241),
    .A1(net558),
    .S(\b_register.n_load ),
    .X(_0091_));
 sg13g2_mux2_1 _1363_ (.A0(net240),
    .A1(net559),
    .S(\b_register.n_load ),
    .X(_0092_));
 sg13g2_nand2_1 _1364_ (.Y(_0511_),
    .A(net342),
    .B(net253));
 sg13g2_o21ai_1 _1365_ (.B1(_0511_),
    .Y(_0093_),
    .A1(_0257_),
    .A2(net253));
 sg13g2_mux2_1 _1366_ (.A0(\accumulator_object.bus[5] ),
    .A1(net561),
    .S(net253),
    .X(_0094_));
 sg13g2_mux2_1 _1367_ (.A0(\accumulator_object.bus[6] ),
    .A1(net568),
    .S(net253),
    .X(_0095_));
 sg13g2_mux2_1 _1368_ (.A0(\accumulator_object.bus[7] ),
    .A1(net560),
    .S(net253),
    .X(_0096_));
 sg13g2_nand2b_2 _1369_ (.Y(_0512_),
    .B(net256),
    .A_N(net257));
 sg13g2_nor2_2 _1370_ (.A(_0492_),
    .B(_0512_),
    .Y(_0513_));
 sg13g2_mux2_1 _1371_ (.A0(net504),
    .A1(net273),
    .S(_0513_),
    .X(_0097_));
 sg13g2_mux2_1 _1372_ (.A0(net420),
    .A1(net271),
    .S(_0513_),
    .X(_0098_));
 sg13g2_mux2_1 _1373_ (.A0(net510),
    .A1(net269),
    .S(_0513_),
    .X(_0099_));
 sg13g2_mux2_1 _1374_ (.A0(net365),
    .A1(net267),
    .S(_0513_),
    .X(_0100_));
 sg13g2_mux2_1 _1375_ (.A0(net412),
    .A1(net265),
    .S(_0513_),
    .X(_0101_));
 sg13g2_mux2_1 _1376_ (.A0(net460),
    .A1(net263),
    .S(_0513_),
    .X(_0102_));
 sg13g2_mux2_1 _1377_ (.A0(net533),
    .A1(net261),
    .S(_0513_),
    .X(_0103_));
 sg13g2_mux2_1 _1378_ (.A0(net453),
    .A1(net259),
    .S(_0513_),
    .X(_0104_));
 sg13g2_nor2_2 _1379_ (.A(_0497_),
    .B(_0512_),
    .Y(_0514_));
 sg13g2_mux2_1 _1380_ (.A0(net532),
    .A1(net273),
    .S(_0514_),
    .X(_0105_));
 sg13g2_mux2_1 _1381_ (.A0(net540),
    .A1(net271),
    .S(_0514_),
    .X(_0106_));
 sg13g2_mux2_1 _1382_ (.A0(net374),
    .A1(net269),
    .S(_0514_),
    .X(_0107_));
 sg13g2_mux2_1 _1383_ (.A0(net518),
    .A1(net267),
    .S(_0514_),
    .X(_0108_));
 sg13g2_mux2_1 _1384_ (.A0(net536),
    .A1(net265),
    .S(_0514_),
    .X(_0109_));
 sg13g2_mux2_1 _1385_ (.A0(net376),
    .A1(net263),
    .S(_0514_),
    .X(_0110_));
 sg13g2_mux2_1 _1386_ (.A0(net478),
    .A1(net261),
    .S(_0514_),
    .X(_0111_));
 sg13g2_mux2_1 _1387_ (.A0(net433),
    .A1(net259),
    .S(_0514_),
    .X(_0112_));
 sg13g2_nor2_2 _1388_ (.A(_0493_),
    .B(_0505_),
    .Y(_0515_));
 sg13g2_mux2_1 _1389_ (.A0(net429),
    .A1(net272),
    .S(net242),
    .X(_0113_));
 sg13g2_mux2_1 _1390_ (.A0(net502),
    .A1(net270),
    .S(_0515_),
    .X(_0114_));
 sg13g2_mux2_1 _1391_ (.A0(net439),
    .A1(net268),
    .S(_0515_),
    .X(_0115_));
 sg13g2_mux2_1 _1392_ (.A0(net500),
    .A1(net266),
    .S(net242),
    .X(_0116_));
 sg13g2_mux2_1 _1393_ (.A0(net492),
    .A1(net264),
    .S(net242),
    .X(_0117_));
 sg13g2_nand2_1 _1394_ (.Y(_0516_),
    .A(net262),
    .B(net242));
 sg13g2_o21ai_1 _1395_ (.B1(_0516_),
    .Y(_0118_),
    .A1(_0278_),
    .A2(net242));
 sg13g2_nand2_1 _1396_ (.Y(_0517_),
    .A(net260),
    .B(net242));
 sg13g2_o21ai_1 _1397_ (.B1(_0517_),
    .Y(_0119_),
    .A1(_0279_),
    .A2(net242));
 sg13g2_nand2_1 _1398_ (.Y(_0518_),
    .A(net258),
    .B(_0515_));
 sg13g2_o21ai_1 _1399_ (.B1(_0518_),
    .Y(_0120_),
    .A1(_0280_),
    .A2(net242));
 sg13g2_nor2_2 _1400_ (.A(_0493_),
    .B(_0502_),
    .Y(_0519_));
 sg13g2_mux2_1 _1401_ (.A0(net534),
    .A1(net272),
    .S(_0519_),
    .X(_0121_));
 sg13g2_mux2_1 _1402_ (.A0(net328),
    .A1(net270),
    .S(_0519_),
    .X(_0122_));
 sg13g2_mux2_1 _1403_ (.A0(net334),
    .A1(net268),
    .S(_0519_),
    .X(_0123_));
 sg13g2_mux2_1 _1404_ (.A0(net335),
    .A1(net266),
    .S(_0519_),
    .X(_0124_));
 sg13g2_mux2_1 _1405_ (.A0(net350),
    .A1(net264),
    .S(_0519_),
    .X(_0125_));
 sg13g2_mux2_1 _1406_ (.A0(net427),
    .A1(net262),
    .S(_0519_),
    .X(_0126_));
 sg13g2_mux2_1 _1407_ (.A0(net414),
    .A1(net260),
    .S(_0519_),
    .X(_0127_));
 sg13g2_mux2_1 _1408_ (.A0(net404),
    .A1(net258),
    .S(_0519_),
    .X(_0128_));
 sg13g2_nand2b_1 _1409_ (.Y(_0520_),
    .B(net380),
    .A_N(net249));
 sg13g2_or4_1 _1410_ (.A(_0561_),
    .B(\alu_object.addsub.genblk1[0].fa.sum ),
    .C(\alu_object.addsub.genblk1[1].fa.sum ),
    .D(\alu_object.addsub.genblk1[2].fa.sum ),
    .X(_0521_));
 sg13g2_nor4_1 _1411_ (.A(\alu_object.addsub.genblk1[3].fa.sum ),
    .B(\alu_object.addsub.genblk1[4].fa.sum ),
    .C(\alu_object.addsub.genblk1[5].fa.sum ),
    .D(_0521_),
    .Y(_0522_));
 sg13g2_nand4_1 _1412_ (.B(_0344_),
    .C(_0345_),
    .A(_0337_),
    .Y(_0523_),
    .D(_0522_));
 sg13g2_a21oi_1 _1413_ (.A1(_0520_),
    .A2(_0523_),
    .Y(_0129_),
    .B1(_0271_));
 sg13g2_nand2b_1 _1414_ (.Y(_0524_),
    .B(net381),
    .A_N(net249));
 sg13g2_nor2_1 _1415_ (.A(_0561_),
    .B(_0339_),
    .Y(_0525_));
 sg13g2_o21ai_1 _1416_ (.B1(_0525_),
    .Y(_0526_),
    .A1(_0340_),
    .A2(_0343_));
 sg13g2_a21oi_1 _1417_ (.A1(_0524_),
    .A2(_0526_),
    .Y(_0130_),
    .B1(_0271_));
 sg13g2_o21ai_1 _1418_ (.B1(net309),
    .Y(_0527_),
    .A1(\accumulator_object.bus[0] ),
    .A2(net246));
 sg13g2_a21oi_1 _1419_ (.A1(net246),
    .A2(_0270_),
    .Y(_0131_),
    .B1(_0527_));
 sg13g2_o21ai_1 _1420_ (.B1(net313),
    .Y(_0528_),
    .A1(\accumulator_object.bus[1] ),
    .A2(net246));
 sg13g2_a21oi_1 _1421_ (.A1(net245),
    .A2(_0269_),
    .Y(_0132_),
    .B1(_0528_));
 sg13g2_o21ai_1 _1422_ (.B1(net313),
    .Y(_0529_),
    .A1(net241),
    .A2(net245));
 sg13g2_a21oi_1 _1423_ (.A1(net245),
    .A2(_0268_),
    .Y(_0133_),
    .B1(_0529_));
 sg13g2_o21ai_1 _1424_ (.B1(net313),
    .Y(_0530_),
    .A1(net240),
    .A2(net245));
 sg13g2_a21oi_1 _1425_ (.A1(net245),
    .A2(_0267_),
    .Y(_0134_),
    .B1(_0530_));
 sg13g2_o21ai_1 _1426_ (.B1(net311),
    .Y(_0531_),
    .A1(\accumulator_object.bus[4] ),
    .A2(net246));
 sg13g2_a21oi_1 _1427_ (.A1(net246),
    .A2(_0266_),
    .Y(_0135_),
    .B1(_0531_));
 sg13g2_o21ai_1 _1428_ (.B1(net310),
    .Y(_0532_),
    .A1(\accumulator_object.bus[5] ),
    .A2(\accumulator_object.load ));
 sg13g2_a21oi_1 _1429_ (.A1(net245),
    .A2(_0265_),
    .Y(_0136_),
    .B1(_0532_));
 sg13g2_o21ai_1 _1430_ (.B1(net310),
    .Y(_0533_),
    .A1(\accumulator_object.bus[6] ),
    .A2(net245));
 sg13g2_a21oi_1 _1431_ (.A1(net245),
    .A2(_0264_),
    .Y(_0137_),
    .B1(_0533_));
 sg13g2_o21ai_1 _1432_ (.B1(net314),
    .Y(_0534_),
    .A1(\accumulator_object.bus[7] ),
    .A2(net246));
 sg13g2_a21oi_1 _1433_ (.A1(_0263_),
    .A2(net246),
    .Y(_0138_),
    .B1(_0534_));
 sg13g2_mux2_1 _1434_ (.A0(\accumulator_object.bus[0] ),
    .A1(net272),
    .S(net247),
    .X(_0139_));
 sg13g2_nand2_1 _1435_ (.Y(_0535_),
    .A(net270),
    .B(net247));
 sg13g2_o21ai_1 _1436_ (.B1(_0535_),
    .Y(_0140_),
    .A1(_0260_),
    .A2(net247));
 sg13g2_mux2_1 _1437_ (.A0(net241),
    .A1(net268),
    .S(\cb.control_signals[10] ),
    .X(_0141_));
 sg13g2_mux2_1 _1438_ (.A0(net240),
    .A1(net266),
    .S(net247),
    .X(_0142_));
 sg13g2_nand2_1 _1439_ (.Y(_0536_),
    .A(net264),
    .B(net247));
 sg13g2_o21ai_1 _1440_ (.B1(_0536_),
    .Y(_0143_),
    .A1(_0257_),
    .A2(net247));
 sg13g2_mux2_1 _1441_ (.A0(\accumulator_object.bus[5] ),
    .A1(net262),
    .S(\cb.control_signals[10] ),
    .X(_0144_));
 sg13g2_mux2_1 _1442_ (.A0(\accumulator_object.bus[6] ),
    .A1(net260),
    .S(net247),
    .X(_0145_));
 sg13g2_mux2_1 _1443_ (.A0(\accumulator_object.bus[7] ),
    .A1(net258),
    .S(net247),
    .X(_0146_));
 sg13g2_nand2b_1 _1444_ (.Y(_0537_),
    .B(net306),
    .A_N(HF));
 sg13g2_nor2_1 _1445_ (.A(HF),
    .B(_0499_),
    .Y(_0538_));
 sg13g2_nand2b_1 _1446_ (.Y(_0539_),
    .B(_0284_),
    .A_N(_0281_));
 sg13g2_a22oi_1 _1447_ (.Y(_0540_),
    .B1(_0538_),
    .B2(_0539_),
    .A2(_0299_),
    .A1(net590));
 sg13g2_or2_1 _1448_ (.X(_0147_),
    .B(_0540_),
    .A(_0537_));
 sg13g2_nand2_1 _1449_ (.Y(_0541_),
    .A(\cb.stage[2] ),
    .B(_0284_));
 sg13g2_nand3_1 _1450_ (.B(_0538_),
    .C(_0541_),
    .A(_0286_),
    .Y(_0542_));
 sg13g2_a21o_1 _1451_ (.A2(_0542_),
    .A1(_0500_),
    .B1(_0537_),
    .X(_0148_));
 sg13g2_o21ai_1 _1452_ (.B1(net308),
    .Y(_0543_),
    .A1(net254),
    .A2(\accumulator_object.bus[0] ));
 sg13g2_a21oi_1 _1453_ (.A1(net254),
    .A2(_0262_),
    .Y(_0149_),
    .B1(_0543_));
 sg13g2_o21ai_1 _1454_ (.B1(net307),
    .Y(_0544_),
    .A1(net255),
    .A2(\accumulator_object.bus[1] ));
 sg13g2_a21oi_1 _1455_ (.A1(net255),
    .A2(_0261_),
    .Y(_0150_),
    .B1(_0544_));
 sg13g2_o21ai_1 _1456_ (.B1(net307),
    .Y(_0545_),
    .A1(net255),
    .A2(net241));
 sg13g2_a21oi_1 _1457_ (.A1(net255),
    .A2(_0259_),
    .Y(_0151_),
    .B1(_0545_));
 sg13g2_o21ai_1 _1458_ (.B1(net307),
    .Y(_0546_),
    .A1(net255),
    .A2(net240));
 sg13g2_a21oi_1 _1459_ (.A1(net255),
    .A2(_0258_),
    .Y(_0152_),
    .B1(_0546_));
 sg13g2_a21oi_1 _1460_ (.A1(net255),
    .A2(net588),
    .Y(_0547_),
    .B1(_0271_));
 sg13g2_o21ai_1 _1461_ (.B1(_0547_),
    .Y(_0153_),
    .A1(\cb.control_signals[7] ),
    .A2(_0257_));
 sg13g2_o21ai_1 _1462_ (.B1(net308),
    .Y(_0548_),
    .A1(net254),
    .A2(\accumulator_object.bus[5] ));
 sg13g2_a21oi_1 _1463_ (.A1(net254),
    .A2(_0256_),
    .Y(_0154_),
    .B1(_0548_));
 sg13g2_o21ai_1 _1464_ (.B1(net308),
    .Y(_0549_),
    .A1(net254),
    .A2(\accumulator_object.bus[6] ));
 sg13g2_a21oi_1 _1465_ (.A1(net254),
    .A2(_0255_),
    .Y(_0155_),
    .B1(_0549_));
 sg13g2_o21ai_1 _1466_ (.B1(net308),
    .Y(_0550_),
    .A1(\accumulator_object.bus[7] ),
    .A2(net254));
 sg13g2_a21oi_1 _1467_ (.A1(_0254_),
    .A2(net254),
    .Y(_0156_),
    .B1(_0550_));
 sg13g2_nor3_2 _1468_ (.A(net257),
    .B(net256),
    .C(_0505_),
    .Y(_0551_));
 sg13g2_mux2_1 _1469_ (.A0(net543),
    .A1(net273),
    .S(_0551_),
    .X(_0161_));
 sg13g2_mux2_1 _1470_ (.A0(net415),
    .A1(net271),
    .S(_0551_),
    .X(_0162_));
 sg13g2_mux2_1 _1471_ (.A0(net509),
    .A1(net269),
    .S(_0551_),
    .X(_0163_));
 sg13g2_mux2_1 _1472_ (.A0(net455),
    .A1(net267),
    .S(_0551_),
    .X(_0164_));
 sg13g2_mux2_1 _1473_ (.A0(net406),
    .A1(net265),
    .S(_0551_),
    .X(_0165_));
 sg13g2_mux2_1 _1474_ (.A0(net494),
    .A1(net263),
    .S(_0551_),
    .X(_0166_));
 sg13g2_mux2_1 _1475_ (.A0(net473),
    .A1(net261),
    .S(_0551_),
    .X(_0167_));
 sg13g2_mux2_1 _1476_ (.A0(net507),
    .A1(net259),
    .S(_0551_),
    .X(_0168_));
 sg13g2_nor3_2 _1477_ (.A(net257),
    .B(net256),
    .C(_0492_),
    .Y(_0552_));
 sg13g2_mux2_1 _1478_ (.A0(net353),
    .A1(net273),
    .S(_0552_),
    .X(_0169_));
 sg13g2_mux2_1 _1479_ (.A0(net526),
    .A1(net271),
    .S(_0552_),
    .X(_0170_));
 sg13g2_mux2_1 _1480_ (.A0(net513),
    .A1(net269),
    .S(_0552_),
    .X(_0171_));
 sg13g2_mux2_1 _1481_ (.A0(net524),
    .A1(net267),
    .S(_0552_),
    .X(_0172_));
 sg13g2_mux2_1 _1482_ (.A0(net369),
    .A1(net265),
    .S(_0552_),
    .X(_0173_));
 sg13g2_mux2_1 _1483_ (.A0(net354),
    .A1(net263),
    .S(_0552_),
    .X(_0174_));
 sg13g2_mux2_1 _1484_ (.A0(net349),
    .A1(net261),
    .S(_0552_),
    .X(_0175_));
 sg13g2_mux2_1 _1485_ (.A0(net356),
    .A1(net259),
    .S(_0552_),
    .X(_0176_));
 sg13g2_nor2_2 _1486_ (.A(_0502_),
    .B(_0512_),
    .Y(_0553_));
 sg13g2_mux2_1 _1487_ (.A0(net400),
    .A1(net273),
    .S(_0553_),
    .X(_0177_));
 sg13g2_mux2_1 _1488_ (.A0(net463),
    .A1(net271),
    .S(_0553_),
    .X(_0178_));
 sg13g2_mux2_1 _1489_ (.A0(net479),
    .A1(net269),
    .S(_0553_),
    .X(_0179_));
 sg13g2_mux2_1 _1490_ (.A0(net442),
    .A1(net267),
    .S(_0553_),
    .X(_0180_));
 sg13g2_mux2_1 _1491_ (.A0(net474),
    .A1(net265),
    .S(_0553_),
    .X(_0181_));
 sg13g2_mux2_1 _1492_ (.A0(net457),
    .A1(net263),
    .S(_0553_),
    .X(_0182_));
 sg13g2_mux2_1 _1493_ (.A0(net448),
    .A1(net261),
    .S(_0553_),
    .X(_0183_));
 sg13g2_mux2_1 _1494_ (.A0(net496),
    .A1(net259),
    .S(_0553_),
    .X(_0184_));
 sg13g2_nor2_2 _1495_ (.A(_0505_),
    .B(_0512_),
    .Y(_0554_));
 sg13g2_mux2_1 _1496_ (.A0(net462),
    .A1(net273),
    .S(_0554_),
    .X(_0185_));
 sg13g2_mux2_1 _1497_ (.A0(net465),
    .A1(net271),
    .S(_0554_),
    .X(_0186_));
 sg13g2_mux2_1 _1498_ (.A0(net401),
    .A1(net269),
    .S(_0554_),
    .X(_0187_));
 sg13g2_mux2_1 _1499_ (.A0(net396),
    .A1(net267),
    .S(_0554_),
    .X(_0188_));
 sg13g2_mux2_1 _1500_ (.A0(net435),
    .A1(net265),
    .S(_0554_),
    .X(_0189_));
 sg13g2_mux2_1 _1501_ (.A0(net422),
    .A1(net263),
    .S(_0554_),
    .X(_0190_));
 sg13g2_mux2_1 _1502_ (.A0(net471),
    .A1(net261),
    .S(_0554_),
    .X(_0191_));
 sg13g2_mux2_1 _1503_ (.A0(net446),
    .A1(net259),
    .S(_0554_),
    .X(_0192_));
 sg13g2_nor2_2 _1504_ (.A(_0492_),
    .B(_0503_),
    .Y(_0555_));
 sg13g2_mux2_1 _1505_ (.A0(net373),
    .A1(net272),
    .S(_0555_),
    .X(_0193_));
 sg13g2_mux2_1 _1506_ (.A0(net431),
    .A1(net270),
    .S(_0555_),
    .X(_0194_));
 sg13g2_mux2_1 _1507_ (.A0(net358),
    .A1(\input_mar_register.data[2] ),
    .S(_0555_),
    .X(_0195_));
 sg13g2_mux2_1 _1508_ (.A0(net440),
    .A1(\input_mar_register.data[3] ),
    .S(_0555_),
    .X(_0196_));
 sg13g2_mux2_1 _1509_ (.A0(net408),
    .A1(net264),
    .S(_0555_),
    .X(_0197_));
 sg13g2_mux2_1 _1510_ (.A0(net418),
    .A1(net262),
    .S(_0555_),
    .X(_0198_));
 sg13g2_mux2_1 _1511_ (.A0(net346),
    .A1(net260),
    .S(_0555_),
    .X(_0199_));
 sg13g2_mux2_1 _1512_ (.A0(net528),
    .A1(net258),
    .S(_0555_),
    .X(_0200_));
 sg13g2_nor2_2 _1513_ (.A(_0497_),
    .B(_0503_),
    .Y(_0556_));
 sg13g2_mux2_1 _1514_ (.A0(net347),
    .A1(\input_mar_register.data[0] ),
    .S(_0556_),
    .X(_0201_));
 sg13g2_mux2_1 _1515_ (.A0(net449),
    .A1(net270),
    .S(_0556_),
    .X(_0202_));
 sg13g2_mux2_1 _1516_ (.A0(net424),
    .A1(net268),
    .S(_0556_),
    .X(_0203_));
 sg13g2_mux2_1 _1517_ (.A0(net410),
    .A1(net266),
    .S(_0556_),
    .X(_0204_));
 sg13g2_mux2_1 _1518_ (.A0(net398),
    .A1(net264),
    .S(_0556_),
    .X(_0205_));
 sg13g2_mux2_1 _1519_ (.A0(net361),
    .A1(\input_mar_register.data[5] ),
    .S(_0556_),
    .X(_0206_));
 sg13g2_mux2_1 _1520_ (.A0(net489),
    .A1(net260),
    .S(_0556_),
    .X(_0207_));
 sg13g2_mux2_1 _1521_ (.A0(net487),
    .A1(net258),
    .S(_0556_),
    .X(_0208_));
 sg13g2_nor2_2 _1522_ (.A(_0493_),
    .B(_0497_),
    .Y(_0236_));
 sg13g2_mux2_1 _1523_ (.A0(net459),
    .A1(net272),
    .S(_0236_),
    .X(_0209_));
 sg13g2_mux2_1 _1524_ (.A0(net385),
    .A1(net270),
    .S(_0236_),
    .X(_0210_));
 sg13g2_mux2_1 _1525_ (.A0(net393),
    .A1(net268),
    .S(_0236_),
    .X(_0211_));
 sg13g2_mux2_1 _1526_ (.A0(net425),
    .A1(net266),
    .S(_0236_),
    .X(_0212_));
 sg13g2_mux2_1 _1527_ (.A0(net391),
    .A1(net264),
    .S(_0236_),
    .X(_0213_));
 sg13g2_mux2_1 _1528_ (.A0(net505),
    .A1(net262),
    .S(_0236_),
    .X(_0214_));
 sg13g2_mux2_1 _1529_ (.A0(net476),
    .A1(\input_mar_register.data[6] ),
    .S(_0236_),
    .X(_0215_));
 sg13g2_mux2_1 _1530_ (.A0(net485),
    .A1(\input_mar_register.data[7] ),
    .S(_0236_),
    .X(_0216_));
 sg13g2_nand2_1 _1531_ (.Y(_0237_),
    .A(Cp),
    .B(net587));
 sg13g2_nor2_1 _1532_ (.A(Lp),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_nand3_1 _1533_ (.B(net585),
    .C(_0238_),
    .A(net565),
    .Y(_0239_));
 sg13g2_inv_1 _1534_ (.Y(_0240_),
    .A(_0239_));
 sg13g2_o21ai_1 _1535_ (.B1(net305),
    .Y(_0241_),
    .A1(net241),
    .A2(_0273_));
 sg13g2_and2_1 _1536_ (.A(net585),
    .B(_0241_),
    .X(_0242_));
 sg13g2_a221oi_1 _1537_ (.B2(_0238_),
    .C1(net585),
    .B1(net565),
    .A1(net241),
    .Y(_0243_),
    .A2(Lp));
 sg13g2_nor4_1 _1538_ (.A(_0271_),
    .B(_0240_),
    .C(_0242_),
    .D(_0243_),
    .Y(_0217_));
 sg13g2_o21ai_1 _1539_ (.B1(net305),
    .Y(_0244_),
    .A1(Lp),
    .A2(_0237_));
 sg13g2_nand2_1 _1540_ (.Y(_0245_),
    .A(\accumulator_object.bus[0] ),
    .B(Lp));
 sg13g2_o21ai_1 _1541_ (.B1(_0273_),
    .Y(_0246_),
    .A1(Cp),
    .A2(net587));
 sg13g2_a21oi_1 _1542_ (.A1(_0245_),
    .A2(_0246_),
    .Y(_0224_),
    .B1(_0244_));
 sg13g2_nand2b_1 _1543_ (.Y(_0247_),
    .B(Lp),
    .A_N(net240));
 sg13g2_nand4_1 _1544_ (.B(net570),
    .C(_0239_),
    .A(net305),
    .Y(_0248_),
    .D(_0247_));
 sg13g2_a21oi_1 _1545_ (.A1(net240),
    .A2(Lp),
    .Y(_0249_),
    .B1(_0240_));
 sg13g2_nand2b_1 _1546_ (.Y(_0250_),
    .B(net306),
    .A_N(net570));
 sg13g2_o21ai_1 _1547_ (.B1(_0248_),
    .Y(_0225_),
    .A1(_0249_),
    .A2(_0250_));
 sg13g2_nand2_1 _1548_ (.Y(_0251_),
    .A(_0273_),
    .B(_0237_));
 sg13g2_a21oi_1 _1549_ (.A1(net305),
    .A2(_0251_),
    .Y(_0252_),
    .B1(net565));
 sg13g2_a221oi_1 _1550_ (.B2(_0244_),
    .C1(net566),
    .B1(net565),
    .A1(_0260_),
    .Y(_0226_),
    .A2(Lp));
 sg13g2_nor3_2 _1551_ (.A(net257),
    .B(net256),
    .C(_0502_),
    .Y(_0253_));
 sg13g2_mux2_1 _1552_ (.A0(net339),
    .A1(net273),
    .S(_0253_),
    .X(_0227_));
 sg13g2_mux2_1 _1553_ (.A0(net469),
    .A1(net271),
    .S(_0253_),
    .X(_0228_));
 sg13g2_mux2_1 _1554_ (.A0(net539),
    .A1(net269),
    .S(_0253_),
    .X(_0229_));
 sg13g2_mux2_1 _1555_ (.A0(net389),
    .A1(net267),
    .S(_0253_),
    .X(_0230_));
 sg13g2_mux2_1 _1556_ (.A0(net378),
    .A1(net265),
    .S(_0253_),
    .X(_0231_));
 sg13g2_mux2_1 _1557_ (.A0(net326),
    .A1(net263),
    .S(_0253_),
    .X(_0232_));
 sg13g2_mux2_1 _1558_ (.A0(net325),
    .A1(net261),
    .S(_0253_),
    .X(_0233_));
 sg13g2_mux2_1 _1559_ (.A0(net337),
    .A1(net259),
    .S(_0253_),
    .X(_0234_));
 sg13g2_nand2_2 _1560_ (.Y(_0591_),
    .A(net314),
    .B(net251));
 sg13g2_nand2_2 _1561_ (.Y(_0592_),
    .A(net312),
    .B(net251));
 sg13g2_nand2_2 _1562_ (.Y(_0593_),
    .A(net311),
    .B(net251));
 sg13g2_nand2_2 _1563_ (.Y(_0594_),
    .A(net311),
    .B(net251));
 sg13g2_nand2_2 _1564_ (.Y(_0595_),
    .A(net312),
    .B(net251));
 sg13g2_nand2_2 _1565_ (.Y(_0596_),
    .A(net312),
    .B(net251));
 sg13g2_nand3b_1 _1566_ (.B(net244),
    .C(_0305_),
    .Y(_0599_),
    .A_N(net250));
 sg13g2_nand3b_1 _1567_ (.B(net244),
    .C(_0305_),
    .Y(_0600_),
    .A_N(net250));
 sg13g2_nand3b_1 _1568_ (.B(net244),
    .C(_0305_),
    .Y(_0601_),
    .A_N(net250));
 sg13g2_nand3b_1 _1569_ (.B(net244),
    .C(_0305_),
    .Y(_0602_),
    .A_N(net250));
 sg13g2_nand3b_1 _1570_ (.B(net244),
    .C(_0305_),
    .Y(_0603_),
    .A_N(net250));
 sg13g2_nand3b_1 _1571_ (.B(net244),
    .C(_0305_),
    .Y(_0604_),
    .A_N(net250));
 sg13g2_nand2_2 _1572_ (.Y(_0558_),
    .A(net305),
    .B(\cb.control_signals[13] ));
 sg13g2_nand2_2 _1573_ (.Y(_0562_),
    .A(net312),
    .B(\cb.control_signals[2] ));
 sg13g2_nand2_2 _1574_ (.Y(_0563_),
    .A(net310),
    .B(\cb.control_signals[2] ));
 sg13g2_nand2_2 _1575_ (.Y(_0564_),
    .A(net310),
    .B(net249));
 sg13g2_nand2_2 _1576_ (.Y(_0565_),
    .A(net310),
    .B(net249));
 sg13g2_nand2_2 _1577_ (.Y(_0566_),
    .A(net310),
    .B(net249));
 sg13g2_nand2_2 _1578_ (.Y(_0567_),
    .A(net311),
    .B(net249));
 sg13g2_nand2_2 _1579_ (.Y(_0568_),
    .A(net312),
    .B(net249));
 sg13g2_nand2_2 _1580_ (.Y(_0570_),
    .A(net313),
    .B(\cb.control_signals[4] ));
 sg13g2_nand2_2 _1581_ (.Y(_0571_),
    .A(net313),
    .B(\cb.control_signals[4] ));
 sg13g2_nand2_2 _1582_ (.Y(_0572_),
    .A(net313),
    .B(\cb.control_signals[4] ));
 sg13g2_nand2_2 _1583_ (.Y(_0573_),
    .A(net311),
    .B(\cb.control_signals[4] ));
 sg13g2_nand2_2 _1584_ (.Y(_0574_),
    .A(net310),
    .B(\cb.control_signals[4] ));
 sg13g2_nand2_2 _1585_ (.Y(_0575_),
    .A(net310),
    .B(\cb.control_signals[4] ));
 sg13g2_nand2_2 _1586_ (.Y(_0576_),
    .A(net312),
    .B(\cb.control_signals[4] ));
 sg13g2_nand2_2 _1587_ (.Y(_0559_),
    .A(net305),
    .B(\cb.control_signals[13] ));
 sg13g2_nand2_2 _1588_ (.Y(_0560_),
    .A(net306),
    .B(\cb.control_signals[13] ));
 sg13g2_nand2b_2 _1589_ (.Y(_0578_),
    .B(net308),
    .A_N(\cb.control_signals[6] ));
 sg13g2_nand2b_2 _1590_ (.Y(_0582_),
    .B(net309),
    .A_N(\cb.control_signals[9] ));
 sg13g2_nand2b_2 _1591_ (.Y(_0583_),
    .B(net309),
    .A_N(\cb.control_signals[9] ));
 sg13g2_nand2b_2 _1592_ (.Y(_0584_),
    .B(net309),
    .A_N(\cb.control_signals[9] ));
 sg13g2_nand2b_2 _1593_ (.Y(_0585_),
    .B(net309),
    .A_N(\cb.control_signals[9] ));
 sg13g2_nand2b_2 _1594_ (.Y(_0586_),
    .B(net314),
    .A_N(\cb.control_signals[9] ));
 sg13g2_nand2b_2 _1595_ (.Y(_0587_),
    .B(net313),
    .A_N(\cb.control_signals[9] ));
 sg13g2_nand2b_2 _1596_ (.Y(_0588_),
    .B(net309),
    .A_N(\cb.control_signals[9] ));
 sg13g2_nand2b_2 _1597_ (.Y(_0579_),
    .B(net307),
    .A_N(\cb.control_signals[6] ));
 sg13g2_nand2b_2 _1598_ (.Y(_0580_),
    .B(net307),
    .A_N(\cb.control_signals[6] ));
 sg13g2_nand3b_1 _1599_ (.B(net244),
    .C(_0305_),
    .Y(_0597_),
    .A_N(net250));
 sg13g2_nand2_2 _1600_ (.Y(_0589_),
    .A(net311),
    .B(net251));
 sg13g2_inv_1 _1602__3 (.Y(net234),
    .A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 _1603__4 (.Y(net235),
    .A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 _1604__5 (.Y(net236),
    .A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 _1605__6 (.Y(net237),
    .A(clknet_2_0__leaf_clk));
 sg13g2_inv_1 _1606__7 (.Y(net238),
    .A(clknet_2_0__leaf_clk));
 sg13g2_inv_1 _1607__8 (.Y(net239),
    .A(clknet_2_3__leaf_clk));
 sg13g2_inv_1 _1608__9 (.Y(net315),
    .A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 _1609__10 (.Y(net316),
    .A(clknet_2_3__leaf_clk));
 sg13g2_inv_1 _1610__11 (.Y(net317),
    .A(clknet_2_3__leaf_clk));
 sg13g2_inv_1 _1611__12 (.Y(net318),
    .A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 _1616__13 (.Y(net319),
    .A(clknet_2_0__leaf_clk));
 sg13g2_mux2_1 _1612_ (.A0(\accumulator_object.bus[0] ),
    .A1(net579),
    .S(net248),
    .X(_0157_));
 sg13g2_o21ai_1 _1613_ (.B1(_0490_),
    .Y(_0158_),
    .A1(_0260_),
    .A2(net248));
 sg13g2_mux2_1 _1614_ (.A0(net241),
    .A1(net257),
    .S(net248),
    .X(_0159_));
 sg13g2_mux2_1 _1615_ (.A0(net240),
    .A1(net256),
    .S(net248),
    .X(_0160_));
 sg13g2_inv_1 _1617__14 (.Y(net320),
    .A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 _1618__15 (.Y(net321),
    .A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 _1619__16 (.Y(net322),
    .A(clknet_2_0__leaf_clk));
 sg13g2_inv_1 _1620__17 (.Y(net323),
    .A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 _1621__18 (.Y(net324),
    .A(clknet_2_3__leaf_clk));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbp_1 _1622_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net64),
    .D(net345),
    .Q_N(_0800_),
    .Q(\ram.RAM[4][0] ));
 sg13g2_dfrbp_1 _1623_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net189),
    .D(net364),
    .Q_N(_0799_),
    .Q(\ram.RAM[4][1] ));
 sg13g2_dfrbp_1 _1624_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net188),
    .D(_0041_),
    .Q_N(_0798_),
    .Q(\ram.RAM[4][2] ));
 sg13g2_dfrbp_1 _1625_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net187),
    .D(net403),
    .Q_N(_0797_),
    .Q(\ram.RAM[4][3] ));
 sg13g2_dfrbp_1 _1626_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net186),
    .D(net368),
    .Q_N(_0796_),
    .Q(\ram.RAM[4][4] ));
 sg13g2_dfrbp_1 _1627_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net185),
    .D(net388),
    .Q_N(_0795_),
    .Q(\ram.RAM[4][5] ));
 sg13g2_dfrbp_1 _1628_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net184),
    .D(_0045_),
    .Q_N(_0794_),
    .Q(\ram.RAM[4][6] ));
 sg13g2_dfrbp_1 _1629_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net183),
    .D(net372),
    .Q_N(_0793_),
    .Q(\ram.RAM[4][7] ));
 sg13g2_dfrbp_1 _1630_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net182),
    .D(_0047_),
    .Q_N(_0792_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1631_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net181),
    .D(_0048_),
    .Q_N(_0791_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1632_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net180),
    .D(_0049_),
    .Q_N(_0790_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1633_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net179),
    .D(_0050_),
    .Q_N(_0789_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1634_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net178),
    .D(_0051_),
    .Q_N(_0788_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1635_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net177),
    .D(_0052_),
    .Q_N(_0787_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1636_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net176),
    .D(_0053_),
    .Q_N(_0786_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1637_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net175),
    .D(_0054_),
    .Q_N(_0785_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _1638_ (.CLK(net232),
    .RESET_B(net174),
    .D(_0235_),
    .Q_N(_0784_),
    .Q(\cb.control_signals[13] ));
 sg13g2_dfrbp_1 _1639_ (.CLK(net233),
    .RESET_B(net173),
    .D(_0008_),
    .Q_N(_0783_),
    .Q(Cp));
 sg13g2_dfrbp_1 _1640_ (.CLK(net234),
    .RESET_B(net172),
    .D(_0055_),
    .Q_N(_0782_),
    .Q(\cb.control_signals[7] ));
 sg13g2_dfrbp_1 _1641_ (.CLK(net235),
    .RESET_B(net170),
    .D(_0056_),
    .Q_N(_0781_),
    .Q(\b_register.n_load ));
 sg13g2_dfrbp_1 _1642_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net168),
    .D(_0057_),
    .Q_N(_0780_),
    .Q(\ram.RAM[1][0] ));
 sg13g2_dfrbp_1 _1643_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net167),
    .D(net452),
    .Q_N(_0779_),
    .Q(\ram.RAM[1][1] ));
 sg13g2_dfrbp_1 _1644_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net166),
    .D(_0059_),
    .Q_N(_0778_),
    .Q(\ram.RAM[1][2] ));
 sg13g2_dfrbp_1 _1645_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net165),
    .D(net445),
    .Q_N(_0777_),
    .Q(\ram.RAM[1][3] ));
 sg13g2_dfrbp_1 _1646_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net164),
    .D(net481),
    .Q_N(_0776_),
    .Q(\ram.RAM[1][4] ));
 sg13g2_dfrbp_1 _1647_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net163),
    .D(net484),
    .Q_N(_0775_),
    .Q(\ram.RAM[1][5] ));
 sg13g2_dfrbp_1 _1648_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net162),
    .D(_0063_),
    .Q_N(_0774_),
    .Q(\ram.RAM[1][6] ));
 sg13g2_dfrbp_1 _1649_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net161),
    .D(net395),
    .Q_N(_0773_),
    .Q(\ram.RAM[1][7] ));
 sg13g2_dfrbp_1 _1650_ (.CLK(net236),
    .RESET_B(net160),
    .D(_0065_),
    .Q_N(_0772_),
    .Q(\cb.control_signals[0] ));
 sg13g2_dfrbp_1 _1651_ (.CLK(net237),
    .RESET_B(net158),
    .D(_0066_),
    .Q_N(_0771_),
    .Q(\cb.control_signals[6] ));
 sg13g2_dfrbp_1 _1652_ (.CLK(net238),
    .RESET_B(net156),
    .D(_0067_),
    .Q_N(_0770_),
    .Q(Lp));
 sg13g2_dfrbp_1 _1653_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net154),
    .D(_0068_),
    .Q_N(_0769_),
    .Q(\cb.stage[0] ));
 sg13g2_dfrbp_1 _1654_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net153),
    .D(net331),
    .Q_N(_0768_),
    .Q(\ram.RAM[14][0] ));
 sg13g2_dfrbp_1 _1655_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net152),
    .D(net531),
    .Q_N(_0767_),
    .Q(\ram.RAM[14][1] ));
 sg13g2_dfrbp_1 _1656_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net151),
    .D(_0071_),
    .Q_N(_0766_),
    .Q(\ram.RAM[14][2] ));
 sg13g2_dfrbp_1 _1657_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net150),
    .D(net438),
    .Q_N(_0765_),
    .Q(\ram.RAM[14][3] ));
 sg13g2_dfrbp_1 _1658_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net149),
    .D(net384),
    .Q_N(_0764_),
    .Q(\ram.RAM[14][4] ));
 sg13g2_dfrbp_1 _1659_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net148),
    .D(net333),
    .Q_N(_0763_),
    .Q(\ram.RAM[14][5] ));
 sg13g2_dfrbp_1 _1660_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net147),
    .D(_0075_),
    .Q_N(_0762_),
    .Q(\ram.RAM[14][6] ));
 sg13g2_dfrbp_1 _1661_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net65),
    .D(net341),
    .Q_N(_0801_),
    .Q(\ram.RAM[14][7] ));
 sg13g2_dfrbp_1 _1662_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net66),
    .D(_0004_),
    .Q_N(_0802_),
    .Q(_0000_));
 sg13g2_dfrbp_1 _1663_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net67),
    .D(_0005_),
    .Q_N(_0803_),
    .Q(_0001_));
 sg13g2_dfrbp_1 _1664_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net87),
    .D(_0006_),
    .Q_N(_0804_),
    .Q(_0002_));
 sg13g2_dfrbp_1 _1665_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net146),
    .D(_0007_),
    .Q_N(_0761_),
    .Q(_0003_));
 sg13g2_dfrbp_1 _1666_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net145),
    .D(net546),
    .Q_N(_0760_),
    .Q(\ram.RAM[15][0] ));
 sg13g2_dfrbp_1 _1667_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net144),
    .D(net551),
    .Q_N(_0759_),
    .Q(\ram.RAM[15][1] ));
 sg13g2_dfrbp_1 _1668_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net143),
    .D(net515),
    .Q_N(_0758_),
    .Q(\ram.RAM[15][2] ));
 sg13g2_dfrbp_1 _1669_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net142),
    .D(net548),
    .Q_N(_0757_),
    .Q(\ram.RAM[15][3] ));
 sg13g2_dfrbp_1 _1670_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net141),
    .D(net517),
    .Q_N(_0756_),
    .Q(\ram.RAM[15][4] ));
 sg13g2_dfrbp_1 _1671_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net140),
    .D(net523),
    .Q_N(_0755_),
    .Q(\ram.RAM[15][5] ));
 sg13g2_dfrbp_1 _1672_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net139),
    .D(_0083_),
    .Q_N(_0754_),
    .Q(\ram.RAM[15][6] ));
 sg13g2_dfrbp_1 _1673_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net138),
    .D(net499),
    .Q_N(_0753_),
    .Q(\ram.RAM[15][7] ));
 sg13g2_dfrbp_1 _1674_ (.CLK(net239),
    .RESET_B(net137),
    .D(_0085_),
    .Q_N(_0752_),
    .Q(\cb.read_ui_in ));
 sg13g2_dfrbp_1 _1675_ (.CLK(net315),
    .RESET_B(net135),
    .D(_0086_),
    .Q_N(_0751_),
    .Q(\cb.done_load ));
 sg13g2_dfrbp_1 _1676_ (.CLK(net316),
    .RESET_B(net133),
    .D(_0087_),
    .Q_N(_0750_),
    .Q(\cb.control_signals[2] ));
 sg13g2_dfrbp_1 _1677_ (.CLK(net317),
    .RESET_B(net131),
    .D(_0088_),
    .Q_N(_0749_),
    .Q(\alu_object.addsub.genblk1[0].fa.cin ));
 sg13g2_dfrbp_1 _1678_ (.CLK(net318),
    .RESET_B(net129),
    .D(_0009_),
    .Q_N(_0748_),
    .Q(HF));
 sg13g2_dfrbp_1 _1679_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net128),
    .D(_0089_),
    .Q_N(_0747_),
    .Q(\alu_object.addsub.op_b[0] ));
 sg13g2_dfrbp_1 _1680_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net127),
    .D(_0090_),
    .Q_N(_0746_),
    .Q(\alu_object.addsub.op_b[1] ));
 sg13g2_dfrbp_1 _1681_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net126),
    .D(_0091_),
    .Q_N(_0745_),
    .Q(\alu_object.addsub.op_b[2] ));
 sg13g2_dfrbp_1 _1682_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net125),
    .D(_0092_),
    .Q_N(_0744_),
    .Q(\alu_object.addsub.op_b[3] ));
 sg13g2_dfrbp_1 _1683_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net124),
    .D(_0093_),
    .Q_N(_0743_),
    .Q(\alu_object.addsub.op_b[4] ));
 sg13g2_dfrbp_1 _1684_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net123),
    .D(_0094_),
    .Q_N(_0742_),
    .Q(\alu_object.addsub.op_b[5] ));
 sg13g2_dfrbp_1 _1685_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net122),
    .D(_0095_),
    .Q_N(_0741_),
    .Q(\alu_object.addsub.op_b[6] ));
 sg13g2_dfrbp_1 _1686_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net121),
    .D(_0096_),
    .Q_N(_0740_),
    .Q(\alu_object.addsub.op_b[7] ));
 sg13g2_dfrbp_1 _1687_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net120),
    .D(_0097_),
    .Q_N(_0739_),
    .Q(\ram.RAM[8][0] ));
 sg13g2_dfrbp_1 _1688_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net119),
    .D(net421),
    .Q_N(_0738_),
    .Q(\ram.RAM[8][1] ));
 sg13g2_dfrbp_1 _1689_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net118),
    .D(_0099_),
    .Q_N(_0737_),
    .Q(\ram.RAM[8][2] ));
 sg13g2_dfrbp_1 _1690_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net117),
    .D(net366),
    .Q_N(_0736_),
    .Q(\ram.RAM[8][3] ));
 sg13g2_dfrbp_1 _1691_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net116),
    .D(net413),
    .Q_N(_0735_),
    .Q(\ram.RAM[8][4] ));
 sg13g2_dfrbp_1 _1692_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net115),
    .D(net461),
    .Q_N(_0734_),
    .Q(\ram.RAM[8][5] ));
 sg13g2_dfrbp_1 _1693_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net114),
    .D(_0103_),
    .Q_N(_0733_),
    .Q(\ram.RAM[8][6] ));
 sg13g2_dfrbp_1 _1694_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net113),
    .D(net454),
    .Q_N(_0732_),
    .Q(\ram.RAM[8][7] ));
 sg13g2_dfrbp_1 _1695_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net112),
    .D(_0105_),
    .Q_N(_0731_),
    .Q(\ram.RAM[9][0] ));
 sg13g2_dfrbp_1 _1696_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net111),
    .D(net541),
    .Q_N(_0730_),
    .Q(\ram.RAM[9][1] ));
 sg13g2_dfrbp_1 _1697_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net110),
    .D(_0107_),
    .Q_N(_0729_),
    .Q(\ram.RAM[9][2] ));
 sg13g2_dfrbp_1 _1698_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net109),
    .D(net519),
    .Q_N(_0728_),
    .Q(\ram.RAM[9][3] ));
 sg13g2_dfrbp_1 _1699_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net108),
    .D(net537),
    .Q_N(_0727_),
    .Q(\ram.RAM[9][4] ));
 sg13g2_dfrbp_1 _1700_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net107),
    .D(net377),
    .Q_N(_0726_),
    .Q(\ram.RAM[9][5] ));
 sg13g2_dfrbp_1 _1701_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net106),
    .D(_0111_),
    .Q_N(_0725_),
    .Q(\ram.RAM[9][6] ));
 sg13g2_dfrbp_1 _1702_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net105),
    .D(net434),
    .Q_N(_0724_),
    .Q(\ram.RAM[9][7] ));
 sg13g2_dfrbp_1 _1703_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net104),
    .D(net430),
    .Q_N(_0723_),
    .Q(\ram.RAM[7][0] ));
 sg13g2_dfrbp_1 _1704_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net103),
    .D(net503),
    .Q_N(_0722_),
    .Q(\ram.RAM[7][1] ));
 sg13g2_dfrbp_1 _1705_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net102),
    .D(_0115_),
    .Q_N(_0721_),
    .Q(\ram.RAM[7][2] ));
 sg13g2_dfrbp_1 _1706_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net101),
    .D(net501),
    .Q_N(_0720_),
    .Q(\ram.RAM[7][3] ));
 sg13g2_dfrbp_1 _1707_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net100),
    .D(net493),
    .Q_N(_0719_),
    .Q(\ram.RAM[7][4] ));
 sg13g2_dfrbp_1 _1708_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net99),
    .D(net554),
    .Q_N(_0718_),
    .Q(\ram.RAM[7][5] ));
 sg13g2_dfrbp_1 _1709_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net98),
    .D(net512),
    .Q_N(_0717_),
    .Q(\ram.RAM[7][6] ));
 sg13g2_dfrbp_1 _1710_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net97),
    .D(net468),
    .Q_N(_0716_),
    .Q(\ram.RAM[7][7] ));
 sg13g2_dfrbp_1 _1711_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net96),
    .D(net535),
    .Q_N(_0715_),
    .Q(\ram.RAM[6][0] ));
 sg13g2_dfrbp_1 _1712_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net95),
    .D(net329),
    .Q_N(_0714_),
    .Q(\ram.RAM[6][1] ));
 sg13g2_dfrbp_1 _1713_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net94),
    .D(_0123_),
    .Q_N(_0713_),
    .Q(\ram.RAM[6][2] ));
 sg13g2_dfrbp_1 _1714_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net93),
    .D(net336),
    .Q_N(_0712_),
    .Q(\ram.RAM[6][3] ));
 sg13g2_dfrbp_1 _1715_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net92),
    .D(net351),
    .Q_N(_0711_),
    .Q(\ram.RAM[6][4] ));
 sg13g2_dfrbp_1 _1716_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net91),
    .D(net428),
    .Q_N(_0710_),
    .Q(\ram.RAM[6][5] ));
 sg13g2_dfrbp_1 _1717_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net90),
    .D(_0127_),
    .Q_N(_0709_),
    .Q(\ram.RAM[6][6] ));
 sg13g2_dfrbp_1 _1718_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net89),
    .D(net405),
    .Q_N(_0708_),
    .Q(\ram.RAM[6][7] ));
 sg13g2_dfrbp_1 _1719_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net88),
    .D(_0129_),
    .Q_N(_0707_),
    .Q(ZF));
 sg13g2_dfrbp_1 _1720_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net86),
    .D(net382),
    .Q_N(_0706_),
    .Q(CF));
 sg13g2_dfrbp_1 _1721_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net84),
    .D(_0131_),
    .Q_N(_0705_),
    .Q(\alu_object.addsub.genblk1[0].fa.a ));
 sg13g2_dfrbp_1 _1722_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net82),
    .D(_0132_),
    .Q_N(_0019_),
    .Q(\alu_object.addsub.genblk1[1].fa.a ));
 sg13g2_dfrbp_1 _1723_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net80),
    .D(_0133_),
    .Q_N(_0704_),
    .Q(\alu_object.addsub.genblk1[2].fa.a ));
 sg13g2_dfrbp_1 _1724_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net78),
    .D(_0134_),
    .Q_N(_0703_),
    .Q(\alu_object.addsub.genblk1[3].fa.a ));
 sg13g2_dfrbp_1 _1725_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net76),
    .D(_0135_),
    .Q_N(_0702_),
    .Q(\alu_object.addsub.genblk1[4].fa.a ));
 sg13g2_dfrbp_1 _1726_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net74),
    .D(_0136_),
    .Q_N(_0701_),
    .Q(\alu_object.addsub.genblk1[5].fa.a ));
 sg13g2_dfrbp_1 _1727_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net72),
    .D(_0137_),
    .Q_N(_0700_),
    .Q(\alu_object.addsub.genblk1[6].fa.a ));
 sg13g2_dfrbp_1 _1728_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net70),
    .D(_0138_),
    .Q_N(_0699_),
    .Q(\alu_object.addsub.genblk1[7].fa.a ));
 sg13g2_dfrbp_1 _1729_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net68),
    .D(_0139_),
    .Q_N(_0698_),
    .Q(\input_mar_register.data[0] ));
 sg13g2_dfrbp_1 _1730_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net63),
    .D(_0140_),
    .Q_N(_0697_),
    .Q(\input_mar_register.data[1] ));
 sg13g2_dfrbp_1 _1731_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net62),
    .D(_0141_),
    .Q_N(_0696_),
    .Q(\input_mar_register.data[2] ));
 sg13g2_dfrbp_1 _1732_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net61),
    .D(_0142_),
    .Q_N(_0695_),
    .Q(\input_mar_register.data[3] ));
 sg13g2_dfrbp_1 _1733_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net60),
    .D(_0143_),
    .Q_N(_0694_),
    .Q(\input_mar_register.data[4] ));
 sg13g2_dfrbp_1 _1734_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net59),
    .D(_0144_),
    .Q_N(_0693_),
    .Q(\input_mar_register.data[5] ));
 sg13g2_dfrbp_1 _1735_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net58),
    .D(_0145_),
    .Q_N(_0692_),
    .Q(\input_mar_register.data[6] ));
 sg13g2_dfrbp_1 _1736_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net57),
    .D(_0146_),
    .Q_N(_0691_),
    .Q(\input_mar_register.data[7] ));
 sg13g2_dfrbp_1 _1737_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net56),
    .D(_0147_),
    .Q_N(_0690_),
    .Q(\cb.stage[1] ));
 sg13g2_dfrbp_1 _1738_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net55),
    .D(_0148_),
    .Q_N(_0018_),
    .Q(\cb.stage[2] ));
 sg13g2_dfrbp_1 _1739_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net54),
    .D(_0149_),
    .Q_N(_0689_),
    .Q(\instruction_register.instruction[0] ));
 sg13g2_dfrbp_1 _1740_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net52),
    .D(_0150_),
    .Q_N(_0688_),
    .Q(\instruction_register.instruction[1] ));
 sg13g2_dfrbp_1 _1741_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net50),
    .D(_0151_),
    .Q_N(_0687_),
    .Q(\instruction_register.instruction[2] ));
 sg13g2_dfrbp_1 _1742_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net48),
    .D(_0152_),
    .Q_N(_0686_),
    .Q(\instruction_register.instruction[3] ));
 sg13g2_dfrbp_1 _1743_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net46),
    .D(_0153_),
    .Q_N(_0685_),
    .Q(\instruction_register.instruction[4] ));
 sg13g2_dfrbp_1 _1744_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net44),
    .D(_0154_),
    .Q_N(_0684_),
    .Q(\instruction_register.instruction[5] ));
 sg13g2_dfrbp_1 _1745_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net42),
    .D(_0155_),
    .Q_N(_0683_),
    .Q(\instruction_register.instruction[6] ));
 sg13g2_dfrbp_1 _1746_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net40),
    .D(_0156_),
    .Q_N(_0682_),
    .Q(\instruction_register.instruction[7] ));
 sg13g2_dfrbp_1 _1747_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net38),
    .D(_0157_),
    .Q_N(_0681_),
    .Q(\input_mar_register.addr[0] ));
 sg13g2_dfrbp_1 _1748_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net37),
    .D(_0158_),
    .Q_N(_0680_),
    .Q(\input_mar_register.addr[1] ));
 sg13g2_dfrbp_1 _1749_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net36),
    .D(_0159_),
    .Q_N(_0679_),
    .Q(\input_mar_register.addr[2] ));
 sg13g2_dfrbp_1 _1750_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net35),
    .D(_0160_),
    .Q_N(_0678_),
    .Q(\input_mar_register.addr[3] ));
 sg13g2_dfrbp_1 _1751_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net34),
    .D(_0161_),
    .Q_N(_0677_),
    .Q(\ram.RAM[3][0] ));
 sg13g2_dfrbp_1 _1752_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net33),
    .D(net416),
    .Q_N(_0676_),
    .Q(\ram.RAM[3][1] ));
 sg13g2_dfrbp_1 _1753_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net32),
    .D(_0163_),
    .Q_N(_0675_),
    .Q(\ram.RAM[3][2] ));
 sg13g2_dfrbp_1 _1754_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net31),
    .D(net456),
    .Q_N(_0674_),
    .Q(\ram.RAM[3][3] ));
 sg13g2_dfrbp_1 _1755_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net30),
    .D(net407),
    .Q_N(_0673_),
    .Q(\ram.RAM[3][4] ));
 sg13g2_dfrbp_1 _1756_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net29),
    .D(net495),
    .Q_N(_0672_),
    .Q(\ram.RAM[3][5] ));
 sg13g2_dfrbp_1 _1757_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net28),
    .D(_0167_),
    .Q_N(_0671_),
    .Q(\ram.RAM[3][6] ));
 sg13g2_dfrbp_1 _1758_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net27),
    .D(net508),
    .Q_N(_0670_),
    .Q(\ram.RAM[3][7] ));
 sg13g2_dfrbp_1 _1759_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net26),
    .D(_0169_),
    .Q_N(_0669_),
    .Q(\ram.RAM[0][0] ));
 sg13g2_dfrbp_1 _1760_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net25),
    .D(net527),
    .Q_N(_0668_),
    .Q(\ram.RAM[0][1] ));
 sg13g2_dfrbp_1 _1761_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net24),
    .D(_0171_),
    .Q_N(_0667_),
    .Q(\ram.RAM[0][2] ));
 sg13g2_dfrbp_1 _1762_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net226),
    .D(net525),
    .Q_N(_0666_),
    .Q(\ram.RAM[0][3] ));
 sg13g2_dfrbp_1 _1763_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net225),
    .D(net370),
    .Q_N(_0665_),
    .Q(\ram.RAM[0][4] ));
 sg13g2_dfrbp_1 _1764_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net224),
    .D(net355),
    .Q_N(_0664_),
    .Q(\ram.RAM[0][5] ));
 sg13g2_dfrbp_1 _1765_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net223),
    .D(_0175_),
    .Q_N(_0663_),
    .Q(\ram.RAM[0][6] ));
 sg13g2_dfrbp_1 _1766_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net222),
    .D(net357),
    .Q_N(_0662_),
    .Q(\ram.RAM[0][7] ));
 sg13g2_dfrbp_1 _1767_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net221),
    .D(_0177_),
    .Q_N(_0661_),
    .Q(\ram.RAM[10][0] ));
 sg13g2_dfrbp_1 _1768_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net220),
    .D(net464),
    .Q_N(_0660_),
    .Q(\ram.RAM[10][1] ));
 sg13g2_dfrbp_1 _1769_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net219),
    .D(_0179_),
    .Q_N(_0659_),
    .Q(\ram.RAM[10][2] ));
 sg13g2_dfrbp_1 _1770_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net218),
    .D(net443),
    .Q_N(_0658_),
    .Q(\ram.RAM[10][3] ));
 sg13g2_dfrbp_1 _1771_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net217),
    .D(net475),
    .Q_N(_0657_),
    .Q(\ram.RAM[10][4] ));
 sg13g2_dfrbp_1 _1772_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net216),
    .D(net458),
    .Q_N(_0656_),
    .Q(\ram.RAM[10][5] ));
 sg13g2_dfrbp_1 _1773_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net215),
    .D(_0183_),
    .Q_N(_0655_),
    .Q(\ram.RAM[10][6] ));
 sg13g2_dfrbp_1 _1774_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net214),
    .D(net497),
    .Q_N(_0654_),
    .Q(\ram.RAM[10][7] ));
 sg13g2_dfrbp_1 _1775_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net213),
    .D(_0185_),
    .Q_N(_0653_),
    .Q(\ram.RAM[11][0] ));
 sg13g2_dfrbp_1 _1776_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net212),
    .D(net466),
    .Q_N(_0652_),
    .Q(\ram.RAM[11][1] ));
 sg13g2_dfrbp_1 _1777_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net211),
    .D(_0187_),
    .Q_N(_0651_),
    .Q(\ram.RAM[11][2] ));
 sg13g2_dfrbp_1 _1778_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net210),
    .D(net397),
    .Q_N(_0650_),
    .Q(\ram.RAM[11][3] ));
 sg13g2_dfrbp_1 _1779_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net209),
    .D(net436),
    .Q_N(_0649_),
    .Q(\ram.RAM[11][4] ));
 sg13g2_dfrbp_1 _1780_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net208),
    .D(net423),
    .Q_N(_0648_),
    .Q(\ram.RAM[11][5] ));
 sg13g2_dfrbp_1 _1781_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net207),
    .D(_0191_),
    .Q_N(_0647_),
    .Q(\ram.RAM[11][6] ));
 sg13g2_dfrbp_1 _1782_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net206),
    .D(net447),
    .Q_N(_0646_),
    .Q(\ram.RAM[11][7] ));
 sg13g2_dfrbp_1 _1783_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net205),
    .D(_0193_),
    .Q_N(_0645_),
    .Q(\ram.RAM[12][0] ));
 sg13g2_dfrbp_1 _1784_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net204),
    .D(net432),
    .Q_N(_0644_),
    .Q(\ram.RAM[12][1] ));
 sg13g2_dfrbp_1 _1785_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net203),
    .D(net359),
    .Q_N(_0643_),
    .Q(\ram.RAM[12][2] ));
 sg13g2_dfrbp_1 _1786_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net202),
    .D(net441),
    .Q_N(_0642_),
    .Q(\ram.RAM[12][3] ));
 sg13g2_dfrbp_1 _1787_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net201),
    .D(net409),
    .Q_N(_0641_),
    .Q(\ram.RAM[12][4] ));
 sg13g2_dfrbp_1 _1788_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net200),
    .D(net419),
    .Q_N(_0640_),
    .Q(\ram.RAM[12][5] ));
 sg13g2_dfrbp_1 _1789_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net199),
    .D(_0199_),
    .Q_N(_0639_),
    .Q(\ram.RAM[12][6] ));
 sg13g2_dfrbp_1 _1790_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net198),
    .D(net529),
    .Q_N(_0638_),
    .Q(\ram.RAM[12][7] ));
 sg13g2_dfrbp_1 _1791_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net197),
    .D(net348),
    .Q_N(_0637_),
    .Q(\ram.RAM[13][0] ));
 sg13g2_dfrbp_1 _1792_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net196),
    .D(net450),
    .Q_N(_0636_),
    .Q(\ram.RAM[13][1] ));
 sg13g2_dfrbp_1 _1793_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net195),
    .D(_0203_),
    .Q_N(_0635_),
    .Q(\ram.RAM[13][2] ));
 sg13g2_dfrbp_1 _1794_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net194),
    .D(net411),
    .Q_N(_0634_),
    .Q(\ram.RAM[13][3] ));
 sg13g2_dfrbp_1 _1795_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net193),
    .D(net399),
    .Q_N(_0633_),
    .Q(\ram.RAM[13][4] ));
 sg13g2_dfrbp_1 _1796_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net192),
    .D(net362),
    .Q_N(_0632_),
    .Q(\ram.RAM[13][5] ));
 sg13g2_dfrbp_1 _1797_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net191),
    .D(_0207_),
    .Q_N(_0631_),
    .Q(\ram.RAM[13][6] ));
 sg13g2_dfrbp_1 _1798_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net190),
    .D(net488),
    .Q_N(_0630_),
    .Q(\ram.RAM[13][7] ));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net171),
    .D(_0209_),
    .Q_N(_0629_),
    .Q(\ram.RAM[5][0] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net169),
    .D(net386),
    .Q_N(_0628_),
    .Q(\ram.RAM[5][1] ));
 sg13g2_dfrbp_1 _1801_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net159),
    .D(_0211_),
    .Q_N(_0627_),
    .Q(\ram.RAM[5][2] ));
 sg13g2_dfrbp_1 _1802_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net157),
    .D(net426),
    .Q_N(_0626_),
    .Q(\ram.RAM[5][3] ));
 sg13g2_dfrbp_1 _1803_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net155),
    .D(net392),
    .Q_N(_0625_),
    .Q(\ram.RAM[5][4] ));
 sg13g2_dfrbp_1 _1804_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net136),
    .D(net506),
    .Q_N(_0624_),
    .Q(\ram.RAM[5][5] ));
 sg13g2_dfrbp_1 _1805_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net134),
    .D(net477),
    .Q_N(_0623_),
    .Q(\ram.RAM[5][6] ));
 sg13g2_dfrbp_1 _1806_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net132),
    .D(net486),
    .Q_N(_0622_),
    .Q(\ram.RAM[5][7] ));
 sg13g2_dfrbp_1 _1807_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net130),
    .D(_0217_),
    .Q_N(_0621_),
    .Q(\pc.set_bit_2.S ));
 sg13g2_dfrbp_1 _1808_ (.CLK(net319),
    .RESET_B(net85),
    .D(_0218_),
    .Q_N(_0620_),
    .Q(\cb.control_signals[11] ));
 sg13g2_dfrbp_1 _1809_ (.CLK(net320),
    .RESET_B(net81),
    .D(_0219_),
    .Q_N(_0619_),
    .Q(\cb.control_signals[10] ));
 sg13g2_dfrbp_1 _1810_ (.CLK(net321),
    .RESET_B(net77),
    .D(_0220_),
    .Q_N(_0618_),
    .Q(\cb.control_signals[9] ));
 sg13g2_dfrbp_1 _1811_ (.CLK(net322),
    .RESET_B(net73),
    .D(_0221_),
    .Q_N(_0020_),
    .Q(\cb.control_signals[8] ));
 sg13g2_dfrbp_1 _1812_ (.CLK(net323),
    .RESET_B(net69),
    .D(_0222_),
    .Q_N(_0617_),
    .Q(\accumulator_object.load ));
 sg13g2_dfrbp_1 _1813_ (.CLK(net324),
    .RESET_B(net51),
    .D(_0223_),
    .Q_N(_0616_),
    .Q(\cb.control_signals[4] ));
 sg13g2_dfrbp_1 _1814_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net47),
    .D(_0224_),
    .Q_N(_0615_),
    .Q(\pc.set_bit_0.S ));
 sg13g2_dfrbp_1 _1815_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net43),
    .D(net571),
    .Q_N(_0614_),
    .Q(\pc.set_bit_3.S ));
 sg13g2_dfrbp_1 _1816_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net39),
    .D(_0226_),
    .Q_N(_0613_),
    .Q(\pc.set_bit_1.S ));
 sg13g2_dfrbp_1 _1817_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net83),
    .D(_0227_),
    .Q_N(_0612_),
    .Q(\ram.RAM[2][0] ));
 sg13g2_dfrbp_1 _1818_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net79),
    .D(net470),
    .Q_N(_0611_),
    .Q(\ram.RAM[2][1] ));
 sg13g2_dfrbp_1 _1819_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net75),
    .D(_0229_),
    .Q_N(_0610_),
    .Q(\ram.RAM[2][2] ));
 sg13g2_dfrbp_1 _1820_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net71),
    .D(net390),
    .Q_N(_0609_),
    .Q(\ram.RAM[2][3] ));
 sg13g2_dfrbp_1 _1821_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net53),
    .D(net379),
    .Q_N(_0608_),
    .Q(\ram.RAM[2][4] ));
 sg13g2_dfrbp_1 _1822_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net49),
    .D(net327),
    .Q_N(_0607_),
    .Q(\ram.RAM[2][5] ));
 sg13g2_dfrbp_1 _1823_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net45),
    .D(_0233_),
    .Q_N(_0606_),
    .Q(\ram.RAM[2][6] ));
 sg13g2_dfrbp_1 _1824_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net41),
    .D(net338),
    .Q_N(_0605_),
    .Q(\ram.RAM[2][7] ));
 sg13g2_tiehi _1760__25 (.L_HI(net25));
 sg13g2_tiehi _1759__26 (.L_HI(net26));
 sg13g2_tiehi _1758__27 (.L_HI(net27));
 sg13g2_tiehi _1757__28 (.L_HI(net28));
 sg13g2_tiehi _1756__29 (.L_HI(net29));
 sg13g2_tiehi _1755__30 (.L_HI(net30));
 sg13g2_tiehi _1754__31 (.L_HI(net31));
 sg13g2_tiehi _1753__32 (.L_HI(net32));
 sg13g2_tiehi _1752__33 (.L_HI(net33));
 sg13g2_tiehi _1751__34 (.L_HI(net34));
 sg13g2_tiehi _1750__35 (.L_HI(net35));
 sg13g2_tiehi _1749__36 (.L_HI(net36));
 sg13g2_tiehi _1748__37 (.L_HI(net37));
 sg13g2_tiehi _1747__38 (.L_HI(net38));
 sg13g2_tiehi _1816__39 (.L_HI(net39));
 sg13g2_tiehi _1746__40 (.L_HI(net40));
 sg13g2_tiehi _1824__41 (.L_HI(net41));
 sg13g2_tiehi _1745__42 (.L_HI(net42));
 sg13g2_tiehi _1815__43 (.L_HI(net43));
 sg13g2_tiehi _1744__44 (.L_HI(net44));
 sg13g2_tiehi _1823__45 (.L_HI(net45));
 sg13g2_tiehi _1743__46 (.L_HI(net46));
 sg13g2_tiehi _1814__47 (.L_HI(net47));
 sg13g2_tiehi _1742__48 (.L_HI(net48));
 sg13g2_tiehi _1822__49 (.L_HI(net49));
 sg13g2_tiehi _1741__50 (.L_HI(net50));
 sg13g2_tiehi _1813__51 (.L_HI(net51));
 sg13g2_tiehi _1740__52 (.L_HI(net52));
 sg13g2_tiehi _1821__53 (.L_HI(net53));
 sg13g2_tiehi _1739__54 (.L_HI(net54));
 sg13g2_tiehi _1738__55 (.L_HI(net55));
 sg13g2_tiehi _1737__56 (.L_HI(net56));
 sg13g2_tiehi _1736__57 (.L_HI(net57));
 sg13g2_tiehi _1735__58 (.L_HI(net58));
 sg13g2_tiehi _1734__59 (.L_HI(net59));
 sg13g2_tiehi _1733__60 (.L_HI(net60));
 sg13g2_tiehi _1732__61 (.L_HI(net61));
 sg13g2_tiehi _1731__62 (.L_HI(net62));
 sg13g2_tiehi _1730__63 (.L_HI(net63));
 sg13g2_tiehi _1622__64 (.L_HI(net64));
 sg13g2_tiehi _1661__65 (.L_HI(net65));
 sg13g2_tiehi _1662__66 (.L_HI(net66));
 sg13g2_tiehi _1663__67 (.L_HI(net67));
 sg13g2_tiehi _1729__68 (.L_HI(net68));
 sg13g2_tiehi _1812__69 (.L_HI(net69));
 sg13g2_tiehi _1728__70 (.L_HI(net70));
 sg13g2_tiehi _1820__71 (.L_HI(net71));
 sg13g2_tiehi _1727__72 (.L_HI(net72));
 sg13g2_tiehi _1811__73 (.L_HI(net73));
 sg13g2_tiehi _1726__74 (.L_HI(net74));
 sg13g2_tiehi _1819__75 (.L_HI(net75));
 sg13g2_tiehi _1725__76 (.L_HI(net76));
 sg13g2_tiehi _1810__77 (.L_HI(net77));
 sg13g2_tiehi _1724__78 (.L_HI(net78));
 sg13g2_tiehi _1818__79 (.L_HI(net79));
 sg13g2_tiehi _1723__80 (.L_HI(net80));
 sg13g2_tiehi _1809__81 (.L_HI(net81));
 sg13g2_tiehi _1722__82 (.L_HI(net82));
 sg13g2_tiehi _1817__83 (.L_HI(net83));
 sg13g2_tiehi _1721__84 (.L_HI(net84));
 sg13g2_tiehi _1808__85 (.L_HI(net85));
 sg13g2_tiehi _1720__86 (.L_HI(net86));
 sg13g2_tiehi _1664__87 (.L_HI(net87));
 sg13g2_tiehi _1719__88 (.L_HI(net88));
 sg13g2_tiehi _1718__89 (.L_HI(net89));
 sg13g2_tiehi _1717__90 (.L_HI(net90));
 sg13g2_tiehi _1716__91 (.L_HI(net91));
 sg13g2_tiehi _1715__92 (.L_HI(net92));
 sg13g2_tiehi _1714__93 (.L_HI(net93));
 sg13g2_tiehi _1713__94 (.L_HI(net94));
 sg13g2_tiehi _1712__95 (.L_HI(net95));
 sg13g2_tiehi _1711__96 (.L_HI(net96));
 sg13g2_tiehi _1710__97 (.L_HI(net97));
 sg13g2_tiehi _1709__98 (.L_HI(net98));
 sg13g2_tiehi _1708__99 (.L_HI(net99));
 sg13g2_tiehi _1707__100 (.L_HI(net100));
 sg13g2_tiehi _1706__101 (.L_HI(net101));
 sg13g2_tiehi _1705__102 (.L_HI(net102));
 sg13g2_tiehi _1704__103 (.L_HI(net103));
 sg13g2_tiehi _1703__104 (.L_HI(net104));
 sg13g2_tiehi _1702__105 (.L_HI(net105));
 sg13g2_tiehi _1701__106 (.L_HI(net106));
 sg13g2_tiehi _1700__107 (.L_HI(net107));
 sg13g2_tiehi _1699__108 (.L_HI(net108));
 sg13g2_tiehi _1698__109 (.L_HI(net109));
 sg13g2_tiehi _1697__110 (.L_HI(net110));
 sg13g2_tiehi _1696__111 (.L_HI(net111));
 sg13g2_tiehi _1695__112 (.L_HI(net112));
 sg13g2_tiehi _1694__113 (.L_HI(net113));
 sg13g2_tiehi _1693__114 (.L_HI(net114));
 sg13g2_tiehi _1692__115 (.L_HI(net115));
 sg13g2_tiehi _1691__116 (.L_HI(net116));
 sg13g2_tiehi _1690__117 (.L_HI(net117));
 sg13g2_tiehi _1689__118 (.L_HI(net118));
 sg13g2_tiehi _1688__119 (.L_HI(net119));
 sg13g2_tiehi _1687__120 (.L_HI(net120));
 sg13g2_tiehi _1686__121 (.L_HI(net121));
 sg13g2_tiehi _1685__122 (.L_HI(net122));
 sg13g2_tiehi _1684__123 (.L_HI(net123));
 sg13g2_tiehi _1683__124 (.L_HI(net124));
 sg13g2_tiehi _1682__125 (.L_HI(net125));
 sg13g2_tiehi _1681__126 (.L_HI(net126));
 sg13g2_tiehi _1680__127 (.L_HI(net127));
 sg13g2_tiehi _1679__128 (.L_HI(net128));
 sg13g2_tiehi _1678__129 (.L_HI(net129));
 sg13g2_tiehi _1807__130 (.L_HI(net130));
 sg13g2_tiehi _1677__131 (.L_HI(net131));
 sg13g2_tiehi _1806__132 (.L_HI(net132));
 sg13g2_tiehi _1676__133 (.L_HI(net133));
 sg13g2_tiehi _1805__134 (.L_HI(net134));
 sg13g2_tiehi _1675__135 (.L_HI(net135));
 sg13g2_tiehi _1804__136 (.L_HI(net136));
 sg13g2_tiehi _1674__137 (.L_HI(net137));
 sg13g2_tiehi _1673__138 (.L_HI(net138));
 sg13g2_tiehi _1672__139 (.L_HI(net139));
 sg13g2_tiehi _1671__140 (.L_HI(net140));
 sg13g2_tiehi _1670__141 (.L_HI(net141));
 sg13g2_tiehi _1669__142 (.L_HI(net142));
 sg13g2_tiehi _1668__143 (.L_HI(net143));
 sg13g2_tiehi _1667__144 (.L_HI(net144));
 sg13g2_tiehi _1666__145 (.L_HI(net145));
 sg13g2_tiehi _1665__146 (.L_HI(net146));
 sg13g2_tiehi _1660__147 (.L_HI(net147));
 sg13g2_tiehi _1659__148 (.L_HI(net148));
 sg13g2_tiehi _1658__149 (.L_HI(net149));
 sg13g2_tiehi _1657__150 (.L_HI(net150));
 sg13g2_tiehi _1656__151 (.L_HI(net151));
 sg13g2_tiehi _1655__152 (.L_HI(net152));
 sg13g2_tiehi _1654__153 (.L_HI(net153));
 sg13g2_tiehi _1653__154 (.L_HI(net154));
 sg13g2_tiehi _1803__155 (.L_HI(net155));
 sg13g2_tiehi _1652__156 (.L_HI(net156));
 sg13g2_tiehi _1802__157 (.L_HI(net157));
 sg13g2_tiehi _1651__158 (.L_HI(net158));
 sg13g2_tiehi _1801__159 (.L_HI(net159));
 sg13g2_tiehi _1650__160 (.L_HI(net160));
 sg13g2_tiehi _1649__161 (.L_HI(net161));
 sg13g2_tiehi _1648__162 (.L_HI(net162));
 sg13g2_tiehi _1647__163 (.L_HI(net163));
 sg13g2_tiehi _1646__164 (.L_HI(net164));
 sg13g2_tiehi _1645__165 (.L_HI(net165));
 sg13g2_tiehi _1644__166 (.L_HI(net166));
 sg13g2_tiehi _1643__167 (.L_HI(net167));
 sg13g2_tiehi _1642__168 (.L_HI(net168));
 sg13g2_tiehi _1800__169 (.L_HI(net169));
 sg13g2_tiehi _1641__170 (.L_HI(net170));
 sg13g2_tiehi _1799__171 (.L_HI(net171));
 sg13g2_tiehi _1640__172 (.L_HI(net172));
 sg13g2_tiehi _1639__173 (.L_HI(net173));
 sg13g2_tiehi _1638__174 (.L_HI(net174));
 sg13g2_tiehi _1637__175 (.L_HI(net175));
 sg13g2_tiehi _1636__176 (.L_HI(net176));
 sg13g2_tiehi _1635__177 (.L_HI(net177));
 sg13g2_tiehi _1634__178 (.L_HI(net178));
 sg13g2_tiehi _1633__179 (.L_HI(net179));
 sg13g2_tiehi _1632__180 (.L_HI(net180));
 sg13g2_tiehi _1631__181 (.L_HI(net181));
 sg13g2_tiehi _1630__182 (.L_HI(net182));
 sg13g2_tiehi _1629__183 (.L_HI(net183));
 sg13g2_tiehi _1628__184 (.L_HI(net184));
 sg13g2_tiehi _1627__185 (.L_HI(net185));
 sg13g2_tiehi _1626__186 (.L_HI(net186));
 sg13g2_tiehi _1625__187 (.L_HI(net187));
 sg13g2_tiehi _1624__188 (.L_HI(net188));
 sg13g2_tiehi _1623__189 (.L_HI(net189));
 sg13g2_tiehi _1798__190 (.L_HI(net190));
 sg13g2_tiehi _1797__191 (.L_HI(net191));
 sg13g2_tiehi _1796__192 (.L_HI(net192));
 sg13g2_tiehi _1795__193 (.L_HI(net193));
 sg13g2_tiehi _1794__194 (.L_HI(net194));
 sg13g2_tiehi _1793__195 (.L_HI(net195));
 sg13g2_tiehi _1792__196 (.L_HI(net196));
 sg13g2_tiehi _1791__197 (.L_HI(net197));
 sg13g2_tiehi _1790__198 (.L_HI(net198));
 sg13g2_tiehi _1789__199 (.L_HI(net199));
 sg13g2_tiehi _1788__200 (.L_HI(net200));
 sg13g2_tiehi _1787__201 (.L_HI(net201));
 sg13g2_tiehi _1786__202 (.L_HI(net202));
 sg13g2_tiehi _1785__203 (.L_HI(net203));
 sg13g2_tiehi _1784__204 (.L_HI(net204));
 sg13g2_tiehi _1783__205 (.L_HI(net205));
 sg13g2_tiehi _1782__206 (.L_HI(net206));
 sg13g2_tiehi _1781__207 (.L_HI(net207));
 sg13g2_tiehi _1780__208 (.L_HI(net208));
 sg13g2_tiehi _1779__209 (.L_HI(net209));
 sg13g2_tiehi _1778__210 (.L_HI(net210));
 sg13g2_tiehi _1777__211 (.L_HI(net211));
 sg13g2_tiehi _1776__212 (.L_HI(net212));
 sg13g2_tiehi _1775__213 (.L_HI(net213));
 sg13g2_tiehi _1774__214 (.L_HI(net214));
 sg13g2_tiehi _1773__215 (.L_HI(net215));
 sg13g2_tiehi _1772__216 (.L_HI(net216));
 sg13g2_tiehi _1771__217 (.L_HI(net217));
 sg13g2_tiehi _1770__218 (.L_HI(net218));
 sg13g2_tiehi _1769__219 (.L_HI(net219));
 sg13g2_tiehi _1768__220 (.L_HI(net220));
 sg13g2_tiehi _1767__221 (.L_HI(net221));
 sg13g2_tiehi _1766__222 (.L_HI(net222));
 sg13g2_tiehi _1765__223 (.L_HI(net223));
 sg13g2_tiehi _1764__224 (.L_HI(net224));
 sg13g2_tiehi _1763__225 (.L_HI(net225));
 sg13g2_tiehi _1762__226 (.L_HI(net226));
 sg13g2_tiehi tt_um_ece298a_8_bit_cpu_top_227 (.L_HI(net227));
 sg13g2_tiehi tt_um_ece298a_8_bit_cpu_top_228 (.L_HI(net228));
 sg13g2_tiehi tt_um_ece298a_8_bit_cpu_top_229 (.L_HI(net229));
 sg13g2_tiehi tt_um_ece298a_8_bit_cpu_top_230 (.L_HI(net230));
 sg13g2_tiehi tt_um_ece298a_8_bit_cpu_top_231 (.L_HI(net231));
 sg13g2_inv_1 _1043__1 (.Y(net232),
    .A(clknet_2_0__leaf_clk));
 sg13g2_tielo _2093__11 (.L_LO(net11));
 sg13g2_tielo _2094__12 (.L_LO(net12));
 sg13g2_tielo _2095__13 (.L_LO(net13));
 sg13g2_tielo _2096__14 (.L_LO(net14));
 sg13g2_tielo _2097__15 (.L_LO(net15));
 sg13g2_tielo _2098__16 (.L_LO(net16));
 sg13g2_tielo _2099__17 (.L_LO(net17));
 sg13g2_tielo tt_um_ece298a_8_bit_cpu_top_18 (.L_LO(net18));
 sg13g2_tielo tt_um_ece298a_8_bit_cpu_top_19 (.L_LO(net19));
 sg13g2_tielo tt_um_ece298a_8_bit_cpu_top_20 (.L_LO(net20));
 sg13g2_tielo tt_um_ece298a_8_bit_cpu_top_21 (.L_LO(net21));
 sg13g2_tielo tt_um_ece298a_8_bit_cpu_top_22 (.L_LO(net22));
 sg13g2_tielo tt_um_ece298a_8_bit_cpu_top_23 (.L_LO(net23));
 sg13g2_tiehi _1761__24 (.L_HI(net24));
 sg13g2_buf_1 _2047_ (.A(\cb.control_signals[13] ),
    .X(uio_out[1]));
 sg13g2_buf_1 _2048_ (.A(\cb.done_load ),
    .X(uio_out[2]));
 sg13g2_buf_1 _2049_ (.A(CF),
    .X(uio_out[3]));
 sg13g2_buf_1 _2050_ (.A(ZF),
    .X(uio_out[4]));
 sg13g2_buf_1 _2051_ (.A(HF),
    .X(uio_out[5]));
 sg13g2_ebufn_8 _2052_ (.Z(\accumulator_object.bus[0] ),
    .A(\pc.set_bit_0.S ),
    .TE_B(_0557_));
 sg13g2_ebufn_8 _2053_ (.Z(\accumulator_object.bus[1] ),
    .A(\pc.set_bit_1.S ),
    .TE_B(_0558_));
 sg13g2_ebufn_8 _2054_ (.Z(\accumulator_object.bus[2] ),
    .A(\pc.set_bit_2.S ),
    .TE_B(_0559_));
 sg13g2_ebufn_8 _2055_ (.Z(\accumulator_object.bus[3] ),
    .A(\pc.set_bit_3.S ),
    .TE_B(_0560_));
 sg13g2_ebufn_8 _2056_ (.Z(\accumulator_object.bus[0] ),
    .A(\alu_object.addsub.genblk1[0].fa.sum ),
    .TE_B(_0561_));
 sg13g2_ebufn_8 _2057_ (.Z(\accumulator_object.bus[1] ),
    .A(\alu_object.addsub.genblk1[1].fa.sum ),
    .TE_B(_0562_));
 sg13g2_ebufn_8 _2058_ (.Z(\accumulator_object.bus[2] ),
    .A(\alu_object.addsub.genblk1[2].fa.sum ),
    .TE_B(_0563_));
 sg13g2_ebufn_8 _2059_ (.Z(\accumulator_object.bus[3] ),
    .A(\alu_object.addsub.genblk1[3].fa.sum ),
    .TE_B(_0564_));
 sg13g2_ebufn_8 _2060_ (.Z(\accumulator_object.bus[4] ),
    .A(\alu_object.addsub.genblk1[4].fa.sum ),
    .TE_B(_0565_));
 sg13g2_ebufn_8 _2061_ (.Z(\accumulator_object.bus[5] ),
    .A(\alu_object.addsub.genblk1[5].fa.sum ),
    .TE_B(_0566_));
 sg13g2_ebufn_8 _2062_ (.Z(\accumulator_object.bus[6] ),
    .A(\alu_object.addsub.genblk1[6].fa.sum ),
    .TE_B(_0567_));
 sg13g2_ebufn_8 _2063_ (.Z(\accumulator_object.bus[7] ),
    .A(\alu_object.addsub.genblk1[7].fa.sum ),
    .TE_B(_0568_));
 sg13g2_ebufn_8 _2064_ (.Z(\accumulator_object.bus[0] ),
    .A(\alu_object.addsub.genblk1[0].fa.a ),
    .TE_B(_0569_));
 sg13g2_ebufn_8 _2065_ (.Z(\accumulator_object.bus[1] ),
    .A(\alu_object.addsub.genblk1[1].fa.a ),
    .TE_B(_0570_));
 sg13g2_ebufn_8 _2066_ (.Z(\accumulator_object.bus[2] ),
    .A(\alu_object.addsub.genblk1[2].fa.a ),
    .TE_B(_0571_));
 sg13g2_ebufn_8 _2067_ (.Z(\accumulator_object.bus[3] ),
    .A(\alu_object.addsub.genblk1[3].fa.a ),
    .TE_B(_0572_));
 sg13g2_ebufn_8 _2068_ (.Z(\accumulator_object.bus[4] ),
    .A(\alu_object.addsub.genblk1[4].fa.a ),
    .TE_B(_0573_));
 sg13g2_ebufn_8 _2069_ (.Z(\accumulator_object.bus[5] ),
    .A(\alu_object.addsub.genblk1[5].fa.a ),
    .TE_B(_0574_));
 sg13g2_ebufn_8 _2070_ (.Z(\accumulator_object.bus[6] ),
    .A(\alu_object.addsub.genblk1[6].fa.a ),
    .TE_B(_0575_));
 sg13g2_ebufn_8 _2071_ (.Z(\accumulator_object.bus[7] ),
    .A(\alu_object.addsub.genblk1[7].fa.a ),
    .TE_B(_0576_));
 sg13g2_ebufn_8 _2072_ (.Z(\accumulator_object.bus[0] ),
    .A(\instruction_register.instruction[0] ),
    .TE_B(_0577_));
 sg13g2_ebufn_8 _2073_ (.Z(\accumulator_object.bus[1] ),
    .A(\instruction_register.instruction[1] ),
    .TE_B(_0578_));
 sg13g2_ebufn_8 _2074_ (.Z(\accumulator_object.bus[2] ),
    .A(\instruction_register.instruction[2] ),
    .TE_B(_0579_));
 sg13g2_ebufn_8 _2075_ (.Z(\accumulator_object.bus[3] ),
    .A(\instruction_register.instruction[3] ),
    .TE_B(_0580_));
 sg13g2_ebufn_8 _2076_ (.Z(\accumulator_object.bus[0] ),
    .A(_0010_),
    .TE_B(_0581_));
 sg13g2_ebufn_8 _2077_ (.Z(\accumulator_object.bus[1] ),
    .A(_0011_),
    .TE_B(_0582_));
 sg13g2_ebufn_8 _2078_ (.Z(\accumulator_object.bus[2] ),
    .A(_0012_),
    .TE_B(_0583_));
 sg13g2_ebufn_8 _2079_ (.Z(\accumulator_object.bus[3] ),
    .A(_0013_),
    .TE_B(_0584_));
 sg13g2_ebufn_8 _2080_ (.Z(\accumulator_object.bus[4] ),
    .A(_0014_),
    .TE_B(_0585_));
 sg13g2_ebufn_8 _2081_ (.Z(\accumulator_object.bus[5] ),
    .A(_0015_),
    .TE_B(_0586_));
 sg13g2_ebufn_8 _2082_ (.Z(\accumulator_object.bus[6] ),
    .A(_0016_),
    .TE_B(_0587_));
 sg13g2_ebufn_8 _2083_ (.Z(\accumulator_object.bus[7] ),
    .A(_0017_),
    .TE_B(_0588_));
 sg13g2_ebufn_8 _2084_ (.Z(\accumulator_object.bus[0] ),
    .A(net1),
    .TE_B(_0589_));
 sg13g2_ebufn_8 _2085_ (.Z(\accumulator_object.bus[1] ),
    .A(net2),
    .TE_B(_0590_));
 sg13g2_ebufn_8 _2086_ (.Z(\accumulator_object.bus[2] ),
    .A(net3),
    .TE_B(_0591_));
 sg13g2_ebufn_8 _2087_ (.Z(\accumulator_object.bus[3] ),
    .A(net4),
    .TE_B(_0592_));
 sg13g2_ebufn_8 _2088_ (.Z(\accumulator_object.bus[4] ),
    .A(net5),
    .TE_B(_0593_));
 sg13g2_ebufn_8 _2089_ (.Z(\accumulator_object.bus[5] ),
    .A(net6),
    .TE_B(_0594_));
 sg13g2_ebufn_8 _2090_ (.Z(\accumulator_object.bus[6] ),
    .A(net7),
    .TE_B(_0595_));
 sg13g2_ebufn_8 _2091_ (.Z(\accumulator_object.bus[7] ),
    .A(net8),
    .TE_B(_0596_));
 sg13g2_ebufn_8 _2092_ (.Z(\accumulator_object.bus[0] ),
    .A(net10),
    .TE_B(_0597_));
 sg13g2_ebufn_8 _2093_ (.Z(\accumulator_object.bus[1] ),
    .A(net11),
    .TE_B(_0598_));
 sg13g2_ebufn_8 _2094_ (.Z(\accumulator_object.bus[2] ),
    .A(net12),
    .TE_B(_0599_));
 sg13g2_ebufn_8 _2095_ (.Z(\accumulator_object.bus[3] ),
    .A(net13),
    .TE_B(_0600_));
 sg13g2_ebufn_8 _2096_ (.Z(\accumulator_object.bus[4] ),
    .A(net14),
    .TE_B(_0601_));
 sg13g2_ebufn_8 _2097_ (.Z(\accumulator_object.bus[5] ),
    .A(net15),
    .TE_B(_0602_));
 sg13g2_ebufn_8 _2098_ (.Z(\accumulator_object.bus[6] ),
    .A(net16),
    .TE_B(_0603_));
 sg13g2_ebufn_8 _2099_ (.Z(\accumulator_object.bus[7] ),
    .A(net17),
    .TE_B(_0604_));
 sg13g2_buf_4 fanout240 (.X(net240),
    .A(\accumulator_object.bus[3] ));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(\accumulator_object.bus[2] ));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(_0515_));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(_0506_));
 sg13g2_buf_2 fanout244 (.A(_0581_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(net246),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(\accumulator_object.load ),
    .X(net246));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(\cb.control_signals[10] ));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(\cb.control_signals[11] ));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(\cb.control_signals[2] ));
 sg13g2_buf_2 fanout250 (.A(\cb.read_ui_in ),
    .X(net250));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(\cb.read_ui_in ));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(\cb.control_signals[0] ));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(\b_register.n_load ));
 sg13g2_buf_2 fanout254 (.A(net255),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(\cb.control_signals[7] ),
    .X(net255));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(net555));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(net556));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(net595));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(\input_mar_register.data[7] ));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(\input_mar_register.data[6] ));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(\input_mar_register.data[6] ));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(net591));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(\input_mar_register.data[5] ));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(net589));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(\input_mar_register.data[4] ));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(net596));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(\input_mar_register.data[3] ));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(\input_mar_register.data[2] ));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(\input_mar_register.data[2] ));
 sg13g2_buf_2 fanout270 (.A(net592),
    .X(net270));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(\input_mar_register.data[1] ));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(net597));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(net598));
 sg13g2_buf_2 fanout274 (.A(net276),
    .X(net274));
 sg13g2_buf_1 fanout275 (.A(net276),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_0003_),
    .X(net276));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(net281));
 sg13g2_buf_2 fanout278 (.A(net281),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_0002_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(net283),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(net285),
    .X(net283));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(net285));
 sg13g2_buf_2 fanout285 (.A(_0001_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(net287),
    .X(net286));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(_0001_));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_0001_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(net292),
    .X(net290));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(net294));
 sg13g2_buf_1 fanout292 (.A(net294),
    .X(net292));
 sg13g2_buf_8 fanout293 (.A(net294),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_0000_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(net299),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(net299),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(net298),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(net299),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(net303),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(net303),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(net302),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(net303),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_0000_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(net9),
    .X(net304));
 sg13g2_buf_4 fanout305 (.X(net305),
    .A(net306));
 sg13g2_buf_2 fanout306 (.A(net307),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(net308),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(rst_n),
    .X(net308));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(net314));
 sg13g2_buf_4 fanout310 (.X(net310),
    .A(net311));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(net312));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(net313));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(net314));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_tielo _2092__10 (.L_LO(net10));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(delaynet_1_clk));
 sg13g2_buf_2 delaybuf_1_clk (.A(delaynet_1_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ram.RAM[2][6] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ram.RAM[2][5] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0232_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold4 (.A(\ram.RAM[6][1] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0122_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold6 (.A(\ram.RAM[14][0] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0069_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold8 (.A(\ram.RAM[14][5] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0074_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold10 (.A(\ram.RAM[6][2] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold11 (.A(\ram.RAM[6][3] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0124_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold13 (.A(\ram.RAM[2][7] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0234_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold15 (.A(\ram.RAM[2][0] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold16 (.A(\ram.RAM[14][7] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0076_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold18 (.A(\alu_object.addsub.op_b[4] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold19 (.A(\ram.RAM[4][6] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold20 (.A(\ram.RAM[4][0] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0039_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold22 (.A(\ram.RAM[12][6] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold23 (.A(\ram.RAM[13][0] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0201_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold25 (.A(\ram.RAM[0][6] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ram.RAM[6][4] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0125_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold28 (.A(\ram.RAM[14][6] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold29 (.A(\ram.RAM[0][0] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold30 (.A(\ram.RAM[0][5] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0174_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold32 (.A(\ram.RAM[0][7] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0176_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ram.RAM[12][2] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0195_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold36 (.A(\ram.RAM[4][2] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold37 (.A(\ram.RAM[13][5] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0206_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold39 (.A(\ram.RAM[4][1] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0040_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold41 (.A(\ram.RAM[8][3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0100_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold43 (.A(\ram.RAM[4][4] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0043_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold45 (.A(\ram.RAM[0][4] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0173_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold47 (.A(\ram.RAM[4][7] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0046_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold49 (.A(\ram.RAM[12][0] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold50 (.A(\ram.RAM[9][2] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold51 (.A(\ram.RAM[1][0] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ram.RAM[9][5] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0110_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ram.RAM[2][4] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0231_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold56 (.A(ZF),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold57 (.A(CF),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0130_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold59 (.A(\ram.RAM[14][4] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0073_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold61 (.A(\ram.RAM[5][1] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0210_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold63 (.A(\ram.RAM[4][5] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0044_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold65 (.A(\ram.RAM[2][3] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0230_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold67 (.A(\ram.RAM[5][4] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0213_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold69 (.A(\ram.RAM[5][2] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold70 (.A(\ram.RAM[1][7] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0064_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold72 (.A(\ram.RAM[11][3] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0188_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold74 (.A(\ram.RAM[13][4] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0205_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold76 (.A(\ram.RAM[10][0] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold77 (.A(\ram.RAM[11][2] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold78 (.A(\ram.RAM[4][3] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0042_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold80 (.A(\ram.RAM[6][7] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0128_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold82 (.A(\ram.RAM[3][4] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0165_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold84 (.A(\ram.RAM[12][4] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0197_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold86 (.A(\ram.RAM[13][3] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0204_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold88 (.A(\ram.RAM[8][4] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0101_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold90 (.A(\ram.RAM[6][6] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold91 (.A(\ram.RAM[3][1] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0162_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold93 (.A(\alu_object.addsub.op_b[1] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold94 (.A(\ram.RAM[12][5] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0198_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold96 (.A(\ram.RAM[8][1] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0098_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold98 (.A(\ram.RAM[11][5] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0190_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold100 (.A(\ram.RAM[13][2] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold101 (.A(\ram.RAM[5][3] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0212_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold103 (.A(\ram.RAM[6][5] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0126_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold105 (.A(\ram.RAM[7][0] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0113_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold107 (.A(\ram.RAM[12][1] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0194_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold109 (.A(\ram.RAM[9][7] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0112_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold111 (.A(\ram.RAM[11][4] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0189_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold113 (.A(\ram.RAM[14][3] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0072_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold115 (.A(\ram.RAM[7][2] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold116 (.A(\ram.RAM[12][3] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0196_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold118 (.A(\ram.RAM[10][3] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0180_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold120 (.A(\ram.RAM[1][3] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0060_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold122 (.A(\ram.RAM[11][7] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0192_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold124 (.A(\ram.RAM[10][6] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold125 (.A(\ram.RAM[13][1] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0202_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold127 (.A(\ram.RAM[1][1] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0058_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold129 (.A(\ram.RAM[8][7] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0104_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold131 (.A(\ram.RAM[3][3] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0164_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold133 (.A(\ram.RAM[10][5] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0182_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold135 (.A(\ram.RAM[5][0] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold136 (.A(\ram.RAM[8][5] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0102_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold138 (.A(\ram.RAM[11][0] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold139 (.A(\ram.RAM[10][1] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0178_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold141 (.A(\ram.RAM[11][1] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0186_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold143 (.A(\ram.RAM[7][7] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0120_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold145 (.A(\ram.RAM[2][1] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0228_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold147 (.A(\ram.RAM[11][6] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold148 (.A(\ram.RAM[1][2] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold149 (.A(\ram.RAM[3][6] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold150 (.A(\ram.RAM[10][4] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0181_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold152 (.A(\ram.RAM[5][6] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0215_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold154 (.A(\ram.RAM[9][6] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold155 (.A(\ram.RAM[10][2] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold156 (.A(\ram.RAM[1][4] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0061_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold158 (.A(\ram.RAM[14][2] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold159 (.A(\ram.RAM[1][5] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0062_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold161 (.A(\ram.RAM[5][7] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0216_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold163 (.A(\ram.RAM[13][7] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0208_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold165 (.A(\ram.RAM[13][6] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold166 (.A(\instruction_register.instruction[1] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold167 (.A(\ram.RAM[1][6] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold168 (.A(\ram.RAM[7][4] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0117_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold170 (.A(\ram.RAM[3][5] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0166_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold172 (.A(\ram.RAM[10][7] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0184_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold174 (.A(\ram.RAM[15][7] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0084_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold176 (.A(\ram.RAM[7][3] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0116_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold178 (.A(\ram.RAM[7][1] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0114_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold180 (.A(\ram.RAM[8][0] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold181 (.A(\ram.RAM[5][5] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0214_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold183 (.A(\ram.RAM[3][7] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0168_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold185 (.A(\ram.RAM[3][2] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold186 (.A(\ram.RAM[8][2] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold187 (.A(\ram.RAM[7][6] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0119_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold189 (.A(\ram.RAM[0][2] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold190 (.A(\ram.RAM[15][2] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0079_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold192 (.A(\ram.RAM[15][4] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0081_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold194 (.A(\ram.RAM[9][3] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0108_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold196 (.A(\ram.RAM[15][6] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold197 (.A(\alu_object.addsub.genblk1[1].fa.a ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold198 (.A(\ram.RAM[15][5] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0082_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold200 (.A(\ram.RAM[0][3] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0172_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold202 (.A(\ram.RAM[0][1] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0170_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold204 (.A(\ram.RAM[12][7] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0200_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold206 (.A(\ram.RAM[14][1] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0070_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold208 (.A(\ram.RAM[9][0] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold209 (.A(\ram.RAM[8][6] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold210 (.A(\ram.RAM[6][0] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0121_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold212 (.A(\ram.RAM[9][4] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0109_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold214 (.A(\instruction_register.instruction[2] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold215 (.A(\ram.RAM[2][2] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold216 (.A(\ram.RAM[9][1] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0106_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold218 (.A(\instruction_register.instruction[3] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold219 (.A(\ram.RAM[3][0] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold220 (.A(uo_out[4]),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold221 (.A(\ram.RAM[15][0] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0077_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold223 (.A(\ram.RAM[15][3] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0080_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold225 (.A(\instruction_register.instruction[0] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold226 (.A(\ram.RAM[15][1] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0078_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold228 (.A(uo_out[1]),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold229 (.A(\ram.RAM[7][5] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0118_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold231 (.A(\input_mar_register.addr[3] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold232 (.A(\input_mar_register.addr[2] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold233 (.A(HF),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold234 (.A(\alu_object.addsub.op_b[2] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold235 (.A(\alu_object.addsub.op_b[3] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold236 (.A(\alu_object.addsub.op_b[7] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold237 (.A(\alu_object.addsub.op_b[5] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold238 (.A(uo_out[3]),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold239 (.A(\alu_object.addsub.genblk1[7].fa.a ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold240 (.A(\alu_object.addsub.genblk1[3].fa.a ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold241 (.A(\pc.set_bit_1.S ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0252_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold243 (.A(uo_out[2]),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold244 (.A(\alu_object.addsub.op_b[6] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold245 (.A(\alu_object.addsub.genblk1[5].fa.a ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold246 (.A(\pc.set_bit_3.S ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0225_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold248 (.A(\alu_object.addsub.genblk1[6].fa.a ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold249 (.A(uo_out[0]),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold250 (.A(uo_out[5]),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold251 (.A(uo_out[6]),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold252 (.A(\alu_object.addsub.genblk1[0].fa.a ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold253 (.A(uo_out[7]),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold254 (.A(\alu_object.addsub.op_b[0] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold255 (.A(\input_mar_register.addr[0] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold256 (.A(\instruction_register.instruction[7] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold257 (.A(\input_mar_register.addr[1] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold258 (.A(\instruction_register.instruction[6] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold259 (.A(\alu_object.addsub.genblk1[2].fa.a ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold260 (.A(\alu_object.addsub.genblk1[4].fa.a ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold261 (.A(\pc.set_bit_2.S ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold262 (.A(\instruction_register.instruction[5] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold263 (.A(\pc.set_bit_0.S ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold264 (.A(\instruction_register.instruction[4] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold265 (.A(\input_mar_register.data[4] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold266 (.A(\cb.stage[2] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold267 (.A(\input_mar_register.data[5] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold268 (.A(\input_mar_register.data[1] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0018_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0501_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold271 (.A(\input_mar_register.data[7] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold272 (.A(\input_mar_register.data[3] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold273 (.A(\input_mar_register.data[0] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold274 (.A(\input_mar_register.data[0] ),
    .X(net598));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_fill_1 FILLER_0_56 ();
 sg13g2_fill_1 FILLER_0_102 ();
 sg13g2_fill_2 FILLER_0_183 ();
 sg13g2_fill_2 FILLER_0_220 ();
 sg13g2_fill_1 FILLER_0_222 ();
 sg13g2_fill_1 FILLER_0_343 ();
 sg13g2_fill_2 FILLER_0_354 ();
 sg13g2_fill_2 FILLER_0_361 ();
 sg13g2_fill_1 FILLER_0_363 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_4 FILLER_1_35 ();
 sg13g2_fill_2 FILLER_1_39 ();
 sg13g2_fill_2 FILLER_1_45 ();
 sg13g2_fill_1 FILLER_1_47 ();
 sg13g2_fill_2 FILLER_1_69 ();
 sg13g2_fill_1 FILLER_1_71 ();
 sg13g2_fill_2 FILLER_1_103 ();
 sg13g2_fill_2 FILLER_1_151 ();
 sg13g2_fill_2 FILLER_1_227 ();
 sg13g2_fill_2 FILLER_1_244 ();
 sg13g2_fill_1 FILLER_1_246 ();
 sg13g2_fill_1 FILLER_1_278 ();
 sg13g2_fill_2 FILLER_1_314 ();
 sg13g2_fill_1 FILLER_1_316 ();
 sg13g2_fill_1 FILLER_1_353 ();
 sg13g2_fill_1 FILLER_1_368 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_4 FILLER_2_28 ();
 sg13g2_fill_1 FILLER_2_32 ();
 sg13g2_fill_2 FILLER_2_42 ();
 sg13g2_fill_2 FILLER_2_67 ();
 sg13g2_fill_1 FILLER_2_79 ();
 sg13g2_fill_2 FILLER_2_119 ();
 sg13g2_fill_1 FILLER_2_296 ();
 sg13g2_fill_2 FILLER_2_347 ();
 sg13g2_fill_2 FILLER_2_390 ();
 sg13g2_fill_1 FILLER_2_392 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_14 ();
 sg13g2_decap_4 FILLER_3_22 ();
 sg13g2_fill_2 FILLER_3_128 ();
 sg13g2_fill_1 FILLER_3_130 ();
 sg13g2_fill_2 FILLER_3_146 ();
 sg13g2_fill_1 FILLER_3_202 ();
 sg13g2_fill_2 FILLER_3_212 ();
 sg13g2_fill_1 FILLER_3_214 ();
 sg13g2_fill_2 FILLER_3_225 ();
 sg13g2_fill_1 FILLER_3_264 ();
 sg13g2_fill_2 FILLER_3_372 ();
 sg13g2_fill_1 FILLER_3_374 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_17 ();
 sg13g2_fill_1 FILLER_4_29 ();
 sg13g2_fill_2 FILLER_4_58 ();
 sg13g2_fill_2 FILLER_4_166 ();
 sg13g2_fill_1 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_135 ();
 sg13g2_fill_1 FILLER_5_137 ();
 sg13g2_fill_2 FILLER_5_156 ();
 sg13g2_fill_2 FILLER_5_192 ();
 sg13g2_fill_1 FILLER_5_194 ();
 sg13g2_fill_1 FILLER_5_259 ();
 sg13g2_fill_2 FILLER_5_381 ();
 sg13g2_fill_2 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_30 ();
 sg13g2_fill_1 FILLER_6_41 ();
 sg13g2_fill_2 FILLER_6_83 ();
 sg13g2_fill_1 FILLER_6_126 ();
 sg13g2_fill_2 FILLER_6_199 ();
 sg13g2_fill_1 FILLER_6_201 ();
 sg13g2_fill_1 FILLER_6_228 ();
 sg13g2_fill_2 FILLER_6_270 ();
 sg13g2_fill_1 FILLER_6_349 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_fill_2 FILLER_7_26 ();
 sg13g2_fill_2 FILLER_7_54 ();
 sg13g2_fill_1 FILLER_7_103 ();
 sg13g2_fill_2 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_156 ();
 sg13g2_fill_1 FILLER_7_158 ();
 sg13g2_fill_2 FILLER_7_198 ();
 sg13g2_fill_1 FILLER_7_200 ();
 sg13g2_fill_2 FILLER_7_210 ();
 sg13g2_fill_1 FILLER_7_212 ();
 sg13g2_fill_1 FILLER_7_217 ();
 sg13g2_fill_1 FILLER_7_257 ();
 sg13g2_fill_1 FILLER_7_267 ();
 sg13g2_fill_1 FILLER_7_297 ();
 sg13g2_fill_1 FILLER_7_317 ();
 sg13g2_fill_2 FILLER_7_353 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_82 ();
 sg13g2_fill_1 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_192 ();
 sg13g2_fill_1 FILLER_8_230 ();
 sg13g2_fill_2 FILLER_8_320 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_fill_1 FILLER_9_26 ();
 sg13g2_fill_2 FILLER_9_82 ();
 sg13g2_fill_1 FILLER_9_98 ();
 sg13g2_fill_2 FILLER_9_241 ();
 sg13g2_fill_1 FILLER_9_243 ();
 sg13g2_fill_2 FILLER_9_292 ();
 sg13g2_fill_1 FILLER_9_294 ();
 sg13g2_fill_1 FILLER_9_304 ();
 sg13g2_fill_2 FILLER_9_314 ();
 sg13g2_fill_1 FILLER_9_357 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_fill_2 FILLER_10_28 ();
 sg13g2_fill_2 FILLER_10_40 ();
 sg13g2_fill_1 FILLER_10_42 ();
 sg13g2_fill_1 FILLER_10_69 ();
 sg13g2_fill_1 FILLER_10_106 ();
 sg13g2_fill_2 FILLER_10_122 ();
 sg13g2_fill_1 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_153 ();
 sg13g2_fill_2 FILLER_10_283 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_106 ();
 sg13g2_fill_1 FILLER_11_108 ();
 sg13g2_fill_2 FILLER_11_135 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_fill_2 FILLER_11_201 ();
 sg13g2_fill_2 FILLER_11_229 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_fill_1 FILLER_11_253 ();
 sg13g2_fill_1 FILLER_11_305 ();
 sg13g2_fill_2 FILLER_11_342 ();
 sg13g2_fill_2 FILLER_11_370 ();
 sg13g2_fill_1 FILLER_11_382 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_50 ();
 sg13g2_fill_2 FILLER_12_135 ();
 sg13g2_fill_1 FILLER_12_156 ();
 sg13g2_fill_1 FILLER_12_224 ();
 sg13g2_fill_2 FILLER_12_234 ();
 sg13g2_fill_2 FILLER_12_312 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_2 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_73 ();
 sg13g2_fill_2 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_197 ();
 sg13g2_fill_1 FILLER_13_199 ();
 sg13g2_fill_2 FILLER_13_256 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_115 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_180 ();
 sg13g2_fill_1 FILLER_14_212 ();
 sg13g2_fill_1 FILLER_14_279 ();
 sg13g2_fill_2 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_358 ();
 sg13g2_fill_2 FILLER_14_368 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_74 ();
 sg13g2_fill_1 FILLER_15_124 ();
 sg13g2_fill_2 FILLER_15_162 ();
 sg13g2_fill_1 FILLER_15_214 ();
 sg13g2_fill_1 FILLER_15_234 ();
 sg13g2_fill_1 FILLER_15_273 ();
 sg13g2_fill_2 FILLER_15_298 ();
 sg13g2_fill_2 FILLER_15_319 ();
 sg13g2_fill_1 FILLER_15_331 ();
 sg13g2_fill_2 FILLER_15_358 ();
 sg13g2_fill_1 FILLER_15_379 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_1 FILLER_16_87 ();
 sg13g2_fill_2 FILLER_16_140 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_251 ();
 sg13g2_fill_1 FILLER_16_253 ();
 sg13g2_fill_1 FILLER_16_295 ();
 sg13g2_fill_1 FILLER_16_340 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_1 FILLER_17_52 ();
 sg13g2_fill_2 FILLER_17_76 ();
 sg13g2_fill_2 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_fill_2 FILLER_17_175 ();
 sg13g2_fill_1 FILLER_17_177 ();
 sg13g2_fill_2 FILLER_17_273 ();
 sg13g2_fill_1 FILLER_17_295 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_40 ();
 sg13g2_fill_1 FILLER_18_63 ();
 sg13g2_fill_2 FILLER_18_135 ();
 sg13g2_fill_1 FILLER_18_178 ();
 sg13g2_fill_2 FILLER_18_269 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_fill_2 FILLER_18_314 ();
 sg13g2_fill_1 FILLER_18_316 ();
 sg13g2_fill_1 FILLER_18_347 ();
 sg13g2_fill_2 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_18_392 ();
 sg13g2_fill_1 FILLER_18_394 ();
 sg13g2_fill_2 FILLER_19_36 ();
 sg13g2_fill_1 FILLER_19_38 ();
 sg13g2_fill_1 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_99 ();
 sg13g2_fill_1 FILLER_19_104 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_170 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_fill_1 FILLER_19_265 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_fill_2 FILLER_19_312 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_20_40 ();
 sg13g2_fill_1 FILLER_20_67 ();
 sg13g2_fill_1 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_141 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_fill_2 FILLER_20_381 ();
 sg13g2_fill_2 FILLER_21_68 ();
 sg13g2_fill_1 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_fill_1 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_198 ();
 sg13g2_decap_4 FILLER_21_209 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_fill_2 FILLER_21_224 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_292 ();
 sg13g2_fill_1 FILLER_21_305 ();
 sg13g2_fill_1 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_104 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_218 ();
 sg13g2_fill_2 FILLER_22_229 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_242 ();
 sg13g2_fill_1 FILLER_22_298 ();
 sg13g2_fill_1 FILLER_22_335 ();
 sg13g2_fill_2 FILLER_22_371 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_47 ();
 sg13g2_fill_2 FILLER_23_59 ();
 sg13g2_fill_1 FILLER_23_61 ();
 sg13g2_fill_2 FILLER_23_109 ();
 sg13g2_fill_1 FILLER_23_111 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_decap_8 FILLER_23_186 ();
 sg13g2_fill_1 FILLER_23_193 ();
 sg13g2_fill_1 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_310 ();
 sg13g2_fill_1 FILLER_23_312 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_27 ();
 sg13g2_fill_2 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_115 ();
 sg13g2_fill_1 FILLER_24_117 ();
 sg13g2_fill_2 FILLER_24_132 ();
 sg13g2_fill_1 FILLER_24_134 ();
 sg13g2_decap_4 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_169 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_213 ();
 sg13g2_decap_8 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_232 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_fill_2 FILLER_24_239 ();
 sg13g2_fill_1 FILLER_24_241 ();
 sg13g2_fill_1 FILLER_24_271 ();
 sg13g2_fill_2 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_1 FILLER_25_51 ();
 sg13g2_fill_1 FILLER_25_124 ();
 sg13g2_decap_8 FILLER_25_162 ();
 sg13g2_decap_4 FILLER_25_169 ();
 sg13g2_decap_4 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_23 ();
 sg13g2_fill_1 FILLER_26_34 ();
 sg13g2_fill_2 FILLER_26_41 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_fill_1 FILLER_26_86 ();
 sg13g2_fill_1 FILLER_26_104 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_4 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_decap_4 FILLER_26_202 ();
 sg13g2_fill_1 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_fill_1 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_285 ();
 sg13g2_fill_1 FILLER_26_311 ();
 sg13g2_fill_2 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_27_26 ();
 sg13g2_fill_2 FILLER_27_33 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_178 ();
 sg13g2_decap_4 FILLER_27_212 ();
 sg13g2_decap_4 FILLER_27_256 ();
 sg13g2_decap_4 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_323 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_fill_1 FILLER_28_72 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_decap_4 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_202 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_240 ();
 sg13g2_decap_4 FILLER_28_274 ();
 sg13g2_fill_1 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_44 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_fill_1 FILLER_29_99 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_decap_4 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_184 ();
 sg13g2_fill_1 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_205 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_240 ();
 sg13g2_decap_4 FILLER_29_266 ();
 sg13g2_fill_2 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_4 ();
 sg13g2_decap_8 FILLER_30_9 ();
 sg13g2_decap_4 FILLER_30_16 ();
 sg13g2_fill_1 FILLER_30_20 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_115 ();
 sg13g2_decap_4 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_202 ();
 sg13g2_decap_4 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_fill_1 FILLER_30_310 ();
 sg13g2_fill_2 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_31_26 ();
 sg13g2_fill_1 FILLER_31_52 ();
 sg13g2_fill_2 FILLER_31_65 ();
 sg13g2_fill_1 FILLER_31_83 ();
 sg13g2_fill_1 FILLER_31_116 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_decap_4 FILLER_31_225 ();
 sg13g2_decap_8 FILLER_31_233 ();
 sg13g2_fill_2 FILLER_31_240 ();
 sg13g2_decap_4 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_fill_2 FILLER_31_283 ();
 sg13g2_fill_1 FILLER_31_285 ();
 sg13g2_fill_2 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_44 ();
 sg13g2_fill_1 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_117 ();
 sg13g2_fill_1 FILLER_32_124 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_decap_4 FILLER_32_232 ();
 sg13g2_fill_2 FILLER_32_236 ();
 sg13g2_decap_4 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_288 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_fill_2 FILLER_32_310 ();
 sg13g2_fill_2 FILLER_32_347 ();
 sg13g2_fill_1 FILLER_33_53 ();
 sg13g2_fill_2 FILLER_33_64 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_decap_4 FILLER_33_148 ();
 sg13g2_fill_1 FILLER_33_152 ();
 sg13g2_fill_1 FILLER_33_195 ();
 sg13g2_fill_2 FILLER_33_199 ();
 sg13g2_fill_1 FILLER_33_201 ();
 sg13g2_decap_4 FILLER_33_206 ();
 sg13g2_fill_1 FILLER_33_210 ();
 sg13g2_decap_4 FILLER_33_214 ();
 sg13g2_fill_2 FILLER_33_218 ();
 sg13g2_decap_8 FILLER_33_230 ();
 sg13g2_fill_2 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_389 ();
 sg13g2_fill_1 FILLER_33_398 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_fill_1 FILLER_34_39 ();
 sg13g2_fill_1 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_115 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_fill_2 FILLER_34_170 ();
 sg13g2_fill_2 FILLER_34_198 ();
 sg13g2_decap_8 FILLER_34_204 ();
 sg13g2_decap_4 FILLER_34_211 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_252 ();
 sg13g2_fill_1 FILLER_34_254 ();
 sg13g2_fill_2 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_300 ();
 sg13g2_fill_2 FILLER_34_367 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_1 FILLER_35_178 ();
 sg13g2_decap_4 FILLER_35_215 ();
 sg13g2_fill_1 FILLER_35_225 ();
 sg13g2_fill_2 FILLER_35_270 ();
 sg13g2_fill_1 FILLER_35_272 ();
 sg13g2_fill_1 FILLER_35_285 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_316 ();
 sg13g2_fill_2 FILLER_35_332 ();
 sg13g2_fill_2 FILLER_35_363 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_11 ();
 sg13g2_fill_2 FILLER_36_23 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_decap_4 FILLER_36_176 ();
 sg13g2_fill_2 FILLER_36_188 ();
 sg13g2_decap_4 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_212 ();
 sg13g2_fill_1 FILLER_36_238 ();
 sg13g2_fill_2 FILLER_36_360 ();
 sg13g2_fill_2 FILLER_36_398 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_89 ();
 sg13g2_fill_2 FILLER_37_177 ();
 sg13g2_fill_1 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_fill_2 FILLER_37_257 ();
 sg13g2_fill_2 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_314 ();
 sg13g2_fill_1 FILLER_37_316 ();
 sg13g2_fill_2 FILLER_37_353 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_37 ();
 sg13g2_fill_2 FILLER_38_141 ();
 sg13g2_fill_2 FILLER_38_205 ();
 sg13g2_fill_1 FILLER_38_207 ();
 sg13g2_fill_1 FILLER_38_283 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_fill_1 FILLER_38_332 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_377 ();
 assign uio_oe[0] = net18;
 assign uio_oe[1] = net227;
 assign uio_oe[2] = net228;
 assign uio_oe[3] = net229;
 assign uio_oe[4] = net230;
 assign uio_oe[5] = net231;
 assign uio_oe[6] = net19;
 assign uio_oe[7] = net20;
 assign uio_out[0] = net21;
 assign uio_out[6] = net22;
 assign uio_out[7] = net23;
endmodule

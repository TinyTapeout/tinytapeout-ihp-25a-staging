module tt_um_algofoogle_tt09_ring_osc2 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire \c0[0] ;
 wire \c0[1] ;
 wire \c0[2] ;
 wire \c0[3] ;
 wire c0clock;
 wire \c1[0] ;
 wire \c1[1] ;
 wire \c1[2] ;
 wire \c1[3] ;
 wire c1clock;
 wire \c2[0] ;
 wire \c2[1] ;
 wire \c2[2] ;
 wire \c2[3] ;
 wire \c2[4] ;
 wire \c2[5] ;
 wire dummy;
 wire fast_osc;
 wire \ring_1001.inv_in[0] ;
 wire \ring_1001.inv_in[1000] ;
 wire \ring_1001.inv_in[100] ;
 wire \ring_1001.inv_in[101] ;
 wire \ring_1001.inv_in[102] ;
 wire \ring_1001.inv_in[103] ;
 wire \ring_1001.inv_in[104] ;
 wire \ring_1001.inv_in[105] ;
 wire \ring_1001.inv_in[106] ;
 wire \ring_1001.inv_in[107] ;
 wire \ring_1001.inv_in[108] ;
 wire \ring_1001.inv_in[109] ;
 wire \ring_1001.inv_in[10] ;
 wire \ring_1001.inv_in[110] ;
 wire \ring_1001.inv_in[111] ;
 wire \ring_1001.inv_in[112] ;
 wire \ring_1001.inv_in[113] ;
 wire \ring_1001.inv_in[114] ;
 wire \ring_1001.inv_in[115] ;
 wire \ring_1001.inv_in[116] ;
 wire \ring_1001.inv_in[117] ;
 wire \ring_1001.inv_in[118] ;
 wire \ring_1001.inv_in[119] ;
 wire \ring_1001.inv_in[11] ;
 wire \ring_1001.inv_in[120] ;
 wire \ring_1001.inv_in[121] ;
 wire \ring_1001.inv_in[122] ;
 wire \ring_1001.inv_in[123] ;
 wire \ring_1001.inv_in[124] ;
 wire \ring_1001.inv_in[125] ;
 wire \ring_1001.inv_in[126] ;
 wire \ring_1001.inv_in[127] ;
 wire \ring_1001.inv_in[128] ;
 wire \ring_1001.inv_in[129] ;
 wire \ring_1001.inv_in[12] ;
 wire \ring_1001.inv_in[130] ;
 wire \ring_1001.inv_in[131] ;
 wire \ring_1001.inv_in[132] ;
 wire \ring_1001.inv_in[133] ;
 wire \ring_1001.inv_in[134] ;
 wire \ring_1001.inv_in[135] ;
 wire \ring_1001.inv_in[136] ;
 wire \ring_1001.inv_in[137] ;
 wire \ring_1001.inv_in[138] ;
 wire \ring_1001.inv_in[139] ;
 wire \ring_1001.inv_in[13] ;
 wire \ring_1001.inv_in[140] ;
 wire \ring_1001.inv_in[141] ;
 wire \ring_1001.inv_in[142] ;
 wire \ring_1001.inv_in[143] ;
 wire \ring_1001.inv_in[144] ;
 wire \ring_1001.inv_in[145] ;
 wire \ring_1001.inv_in[146] ;
 wire \ring_1001.inv_in[147] ;
 wire \ring_1001.inv_in[148] ;
 wire \ring_1001.inv_in[149] ;
 wire \ring_1001.inv_in[14] ;
 wire \ring_1001.inv_in[150] ;
 wire \ring_1001.inv_in[151] ;
 wire \ring_1001.inv_in[152] ;
 wire \ring_1001.inv_in[153] ;
 wire \ring_1001.inv_in[154] ;
 wire \ring_1001.inv_in[155] ;
 wire \ring_1001.inv_in[156] ;
 wire \ring_1001.inv_in[157] ;
 wire \ring_1001.inv_in[158] ;
 wire \ring_1001.inv_in[159] ;
 wire \ring_1001.inv_in[15] ;
 wire \ring_1001.inv_in[160] ;
 wire \ring_1001.inv_in[161] ;
 wire \ring_1001.inv_in[162] ;
 wire \ring_1001.inv_in[163] ;
 wire \ring_1001.inv_in[164] ;
 wire \ring_1001.inv_in[165] ;
 wire \ring_1001.inv_in[166] ;
 wire \ring_1001.inv_in[167] ;
 wire \ring_1001.inv_in[168] ;
 wire \ring_1001.inv_in[169] ;
 wire \ring_1001.inv_in[16] ;
 wire \ring_1001.inv_in[170] ;
 wire \ring_1001.inv_in[171] ;
 wire \ring_1001.inv_in[172] ;
 wire \ring_1001.inv_in[173] ;
 wire \ring_1001.inv_in[174] ;
 wire \ring_1001.inv_in[175] ;
 wire \ring_1001.inv_in[176] ;
 wire \ring_1001.inv_in[177] ;
 wire \ring_1001.inv_in[178] ;
 wire \ring_1001.inv_in[179] ;
 wire \ring_1001.inv_in[17] ;
 wire \ring_1001.inv_in[180] ;
 wire \ring_1001.inv_in[181] ;
 wire \ring_1001.inv_in[182] ;
 wire \ring_1001.inv_in[183] ;
 wire \ring_1001.inv_in[184] ;
 wire \ring_1001.inv_in[185] ;
 wire \ring_1001.inv_in[186] ;
 wire \ring_1001.inv_in[187] ;
 wire \ring_1001.inv_in[188] ;
 wire \ring_1001.inv_in[189] ;
 wire \ring_1001.inv_in[18] ;
 wire \ring_1001.inv_in[190] ;
 wire \ring_1001.inv_in[191] ;
 wire \ring_1001.inv_in[192] ;
 wire \ring_1001.inv_in[193] ;
 wire \ring_1001.inv_in[194] ;
 wire \ring_1001.inv_in[195] ;
 wire \ring_1001.inv_in[196] ;
 wire \ring_1001.inv_in[197] ;
 wire \ring_1001.inv_in[198] ;
 wire \ring_1001.inv_in[199] ;
 wire \ring_1001.inv_in[19] ;
 wire \ring_1001.inv_in[1] ;
 wire \ring_1001.inv_in[200] ;
 wire \ring_1001.inv_in[201] ;
 wire \ring_1001.inv_in[202] ;
 wire \ring_1001.inv_in[203] ;
 wire \ring_1001.inv_in[204] ;
 wire \ring_1001.inv_in[205] ;
 wire \ring_1001.inv_in[206] ;
 wire \ring_1001.inv_in[207] ;
 wire \ring_1001.inv_in[208] ;
 wire \ring_1001.inv_in[209] ;
 wire \ring_1001.inv_in[20] ;
 wire \ring_1001.inv_in[210] ;
 wire \ring_1001.inv_in[211] ;
 wire \ring_1001.inv_in[212] ;
 wire \ring_1001.inv_in[213] ;
 wire \ring_1001.inv_in[214] ;
 wire \ring_1001.inv_in[215] ;
 wire \ring_1001.inv_in[216] ;
 wire \ring_1001.inv_in[217] ;
 wire \ring_1001.inv_in[218] ;
 wire \ring_1001.inv_in[219] ;
 wire \ring_1001.inv_in[21] ;
 wire \ring_1001.inv_in[220] ;
 wire \ring_1001.inv_in[221] ;
 wire \ring_1001.inv_in[222] ;
 wire \ring_1001.inv_in[223] ;
 wire \ring_1001.inv_in[224] ;
 wire \ring_1001.inv_in[225] ;
 wire \ring_1001.inv_in[226] ;
 wire \ring_1001.inv_in[227] ;
 wire \ring_1001.inv_in[228] ;
 wire \ring_1001.inv_in[229] ;
 wire \ring_1001.inv_in[22] ;
 wire \ring_1001.inv_in[230] ;
 wire \ring_1001.inv_in[231] ;
 wire \ring_1001.inv_in[232] ;
 wire \ring_1001.inv_in[233] ;
 wire \ring_1001.inv_in[234] ;
 wire \ring_1001.inv_in[235] ;
 wire \ring_1001.inv_in[236] ;
 wire \ring_1001.inv_in[237] ;
 wire \ring_1001.inv_in[238] ;
 wire \ring_1001.inv_in[239] ;
 wire \ring_1001.inv_in[23] ;
 wire \ring_1001.inv_in[240] ;
 wire \ring_1001.inv_in[241] ;
 wire \ring_1001.inv_in[242] ;
 wire \ring_1001.inv_in[243] ;
 wire \ring_1001.inv_in[244] ;
 wire \ring_1001.inv_in[245] ;
 wire \ring_1001.inv_in[246] ;
 wire \ring_1001.inv_in[247] ;
 wire \ring_1001.inv_in[248] ;
 wire \ring_1001.inv_in[249] ;
 wire \ring_1001.inv_in[24] ;
 wire \ring_1001.inv_in[250] ;
 wire \ring_1001.inv_in[251] ;
 wire \ring_1001.inv_in[252] ;
 wire \ring_1001.inv_in[253] ;
 wire \ring_1001.inv_in[254] ;
 wire \ring_1001.inv_in[255] ;
 wire \ring_1001.inv_in[256] ;
 wire \ring_1001.inv_in[257] ;
 wire \ring_1001.inv_in[258] ;
 wire \ring_1001.inv_in[259] ;
 wire \ring_1001.inv_in[25] ;
 wire \ring_1001.inv_in[260] ;
 wire \ring_1001.inv_in[261] ;
 wire \ring_1001.inv_in[262] ;
 wire \ring_1001.inv_in[263] ;
 wire \ring_1001.inv_in[264] ;
 wire \ring_1001.inv_in[265] ;
 wire \ring_1001.inv_in[266] ;
 wire \ring_1001.inv_in[267] ;
 wire \ring_1001.inv_in[268] ;
 wire \ring_1001.inv_in[269] ;
 wire \ring_1001.inv_in[26] ;
 wire \ring_1001.inv_in[270] ;
 wire \ring_1001.inv_in[271] ;
 wire \ring_1001.inv_in[272] ;
 wire \ring_1001.inv_in[273] ;
 wire \ring_1001.inv_in[274] ;
 wire \ring_1001.inv_in[275] ;
 wire \ring_1001.inv_in[276] ;
 wire \ring_1001.inv_in[277] ;
 wire \ring_1001.inv_in[278] ;
 wire \ring_1001.inv_in[279] ;
 wire \ring_1001.inv_in[27] ;
 wire \ring_1001.inv_in[280] ;
 wire \ring_1001.inv_in[281] ;
 wire \ring_1001.inv_in[282] ;
 wire \ring_1001.inv_in[283] ;
 wire \ring_1001.inv_in[284] ;
 wire \ring_1001.inv_in[285] ;
 wire \ring_1001.inv_in[286] ;
 wire \ring_1001.inv_in[287] ;
 wire \ring_1001.inv_in[288] ;
 wire \ring_1001.inv_in[289] ;
 wire \ring_1001.inv_in[28] ;
 wire \ring_1001.inv_in[290] ;
 wire \ring_1001.inv_in[291] ;
 wire \ring_1001.inv_in[292] ;
 wire \ring_1001.inv_in[293] ;
 wire \ring_1001.inv_in[294] ;
 wire \ring_1001.inv_in[295] ;
 wire \ring_1001.inv_in[296] ;
 wire \ring_1001.inv_in[297] ;
 wire \ring_1001.inv_in[298] ;
 wire \ring_1001.inv_in[299] ;
 wire \ring_1001.inv_in[29] ;
 wire \ring_1001.inv_in[2] ;
 wire \ring_1001.inv_in[300] ;
 wire \ring_1001.inv_in[301] ;
 wire \ring_1001.inv_in[302] ;
 wire \ring_1001.inv_in[303] ;
 wire \ring_1001.inv_in[304] ;
 wire \ring_1001.inv_in[305] ;
 wire \ring_1001.inv_in[306] ;
 wire \ring_1001.inv_in[307] ;
 wire \ring_1001.inv_in[308] ;
 wire \ring_1001.inv_in[309] ;
 wire \ring_1001.inv_in[30] ;
 wire \ring_1001.inv_in[310] ;
 wire \ring_1001.inv_in[311] ;
 wire \ring_1001.inv_in[312] ;
 wire \ring_1001.inv_in[313] ;
 wire \ring_1001.inv_in[314] ;
 wire \ring_1001.inv_in[315] ;
 wire \ring_1001.inv_in[316] ;
 wire \ring_1001.inv_in[317] ;
 wire \ring_1001.inv_in[318] ;
 wire \ring_1001.inv_in[319] ;
 wire \ring_1001.inv_in[31] ;
 wire \ring_1001.inv_in[320] ;
 wire \ring_1001.inv_in[321] ;
 wire \ring_1001.inv_in[322] ;
 wire \ring_1001.inv_in[323] ;
 wire \ring_1001.inv_in[324] ;
 wire \ring_1001.inv_in[325] ;
 wire \ring_1001.inv_in[326] ;
 wire \ring_1001.inv_in[327] ;
 wire \ring_1001.inv_in[328] ;
 wire \ring_1001.inv_in[329] ;
 wire \ring_1001.inv_in[32] ;
 wire \ring_1001.inv_in[330] ;
 wire \ring_1001.inv_in[331] ;
 wire \ring_1001.inv_in[332] ;
 wire \ring_1001.inv_in[333] ;
 wire \ring_1001.inv_in[334] ;
 wire \ring_1001.inv_in[335] ;
 wire \ring_1001.inv_in[336] ;
 wire \ring_1001.inv_in[337] ;
 wire \ring_1001.inv_in[338] ;
 wire \ring_1001.inv_in[339] ;
 wire \ring_1001.inv_in[33] ;
 wire \ring_1001.inv_in[340] ;
 wire \ring_1001.inv_in[341] ;
 wire \ring_1001.inv_in[342] ;
 wire \ring_1001.inv_in[343] ;
 wire \ring_1001.inv_in[344] ;
 wire \ring_1001.inv_in[345] ;
 wire \ring_1001.inv_in[346] ;
 wire \ring_1001.inv_in[347] ;
 wire \ring_1001.inv_in[348] ;
 wire \ring_1001.inv_in[349] ;
 wire \ring_1001.inv_in[34] ;
 wire \ring_1001.inv_in[350] ;
 wire \ring_1001.inv_in[351] ;
 wire \ring_1001.inv_in[352] ;
 wire \ring_1001.inv_in[353] ;
 wire \ring_1001.inv_in[354] ;
 wire \ring_1001.inv_in[355] ;
 wire \ring_1001.inv_in[356] ;
 wire \ring_1001.inv_in[357] ;
 wire \ring_1001.inv_in[358] ;
 wire \ring_1001.inv_in[359] ;
 wire \ring_1001.inv_in[35] ;
 wire \ring_1001.inv_in[360] ;
 wire \ring_1001.inv_in[361] ;
 wire \ring_1001.inv_in[362] ;
 wire \ring_1001.inv_in[363] ;
 wire \ring_1001.inv_in[364] ;
 wire \ring_1001.inv_in[365] ;
 wire \ring_1001.inv_in[366] ;
 wire \ring_1001.inv_in[367] ;
 wire \ring_1001.inv_in[368] ;
 wire \ring_1001.inv_in[369] ;
 wire \ring_1001.inv_in[36] ;
 wire \ring_1001.inv_in[370] ;
 wire \ring_1001.inv_in[371] ;
 wire \ring_1001.inv_in[372] ;
 wire \ring_1001.inv_in[373] ;
 wire \ring_1001.inv_in[374] ;
 wire \ring_1001.inv_in[375] ;
 wire \ring_1001.inv_in[376] ;
 wire \ring_1001.inv_in[377] ;
 wire \ring_1001.inv_in[378] ;
 wire \ring_1001.inv_in[379] ;
 wire \ring_1001.inv_in[37] ;
 wire \ring_1001.inv_in[380] ;
 wire \ring_1001.inv_in[381] ;
 wire \ring_1001.inv_in[382] ;
 wire \ring_1001.inv_in[383] ;
 wire \ring_1001.inv_in[384] ;
 wire \ring_1001.inv_in[385] ;
 wire \ring_1001.inv_in[386] ;
 wire \ring_1001.inv_in[387] ;
 wire \ring_1001.inv_in[388] ;
 wire \ring_1001.inv_in[389] ;
 wire \ring_1001.inv_in[38] ;
 wire \ring_1001.inv_in[390] ;
 wire \ring_1001.inv_in[391] ;
 wire \ring_1001.inv_in[392] ;
 wire \ring_1001.inv_in[393] ;
 wire \ring_1001.inv_in[394] ;
 wire \ring_1001.inv_in[395] ;
 wire \ring_1001.inv_in[396] ;
 wire \ring_1001.inv_in[397] ;
 wire \ring_1001.inv_in[398] ;
 wire \ring_1001.inv_in[399] ;
 wire \ring_1001.inv_in[39] ;
 wire \ring_1001.inv_in[3] ;
 wire \ring_1001.inv_in[400] ;
 wire \ring_1001.inv_in[401] ;
 wire \ring_1001.inv_in[402] ;
 wire \ring_1001.inv_in[403] ;
 wire \ring_1001.inv_in[404] ;
 wire \ring_1001.inv_in[405] ;
 wire \ring_1001.inv_in[406] ;
 wire \ring_1001.inv_in[407] ;
 wire \ring_1001.inv_in[408] ;
 wire \ring_1001.inv_in[409] ;
 wire \ring_1001.inv_in[40] ;
 wire \ring_1001.inv_in[410] ;
 wire \ring_1001.inv_in[411] ;
 wire \ring_1001.inv_in[412] ;
 wire \ring_1001.inv_in[413] ;
 wire \ring_1001.inv_in[414] ;
 wire \ring_1001.inv_in[415] ;
 wire \ring_1001.inv_in[416] ;
 wire \ring_1001.inv_in[417] ;
 wire \ring_1001.inv_in[418] ;
 wire \ring_1001.inv_in[419] ;
 wire \ring_1001.inv_in[41] ;
 wire \ring_1001.inv_in[420] ;
 wire \ring_1001.inv_in[421] ;
 wire \ring_1001.inv_in[422] ;
 wire \ring_1001.inv_in[423] ;
 wire \ring_1001.inv_in[424] ;
 wire \ring_1001.inv_in[425] ;
 wire \ring_1001.inv_in[426] ;
 wire \ring_1001.inv_in[427] ;
 wire \ring_1001.inv_in[428] ;
 wire \ring_1001.inv_in[429] ;
 wire \ring_1001.inv_in[42] ;
 wire \ring_1001.inv_in[430] ;
 wire \ring_1001.inv_in[431] ;
 wire \ring_1001.inv_in[432] ;
 wire \ring_1001.inv_in[433] ;
 wire \ring_1001.inv_in[434] ;
 wire \ring_1001.inv_in[435] ;
 wire \ring_1001.inv_in[436] ;
 wire \ring_1001.inv_in[437] ;
 wire \ring_1001.inv_in[438] ;
 wire \ring_1001.inv_in[439] ;
 wire \ring_1001.inv_in[43] ;
 wire \ring_1001.inv_in[440] ;
 wire \ring_1001.inv_in[441] ;
 wire \ring_1001.inv_in[442] ;
 wire \ring_1001.inv_in[443] ;
 wire \ring_1001.inv_in[444] ;
 wire \ring_1001.inv_in[445] ;
 wire \ring_1001.inv_in[446] ;
 wire \ring_1001.inv_in[447] ;
 wire \ring_1001.inv_in[448] ;
 wire \ring_1001.inv_in[449] ;
 wire \ring_1001.inv_in[44] ;
 wire \ring_1001.inv_in[450] ;
 wire \ring_1001.inv_in[451] ;
 wire \ring_1001.inv_in[452] ;
 wire \ring_1001.inv_in[453] ;
 wire \ring_1001.inv_in[454] ;
 wire \ring_1001.inv_in[455] ;
 wire \ring_1001.inv_in[456] ;
 wire \ring_1001.inv_in[457] ;
 wire \ring_1001.inv_in[458] ;
 wire \ring_1001.inv_in[459] ;
 wire \ring_1001.inv_in[45] ;
 wire \ring_1001.inv_in[460] ;
 wire \ring_1001.inv_in[461] ;
 wire \ring_1001.inv_in[462] ;
 wire \ring_1001.inv_in[463] ;
 wire \ring_1001.inv_in[464] ;
 wire \ring_1001.inv_in[465] ;
 wire \ring_1001.inv_in[466] ;
 wire \ring_1001.inv_in[467] ;
 wire \ring_1001.inv_in[468] ;
 wire \ring_1001.inv_in[469] ;
 wire \ring_1001.inv_in[46] ;
 wire \ring_1001.inv_in[470] ;
 wire \ring_1001.inv_in[471] ;
 wire \ring_1001.inv_in[472] ;
 wire \ring_1001.inv_in[473] ;
 wire \ring_1001.inv_in[474] ;
 wire \ring_1001.inv_in[475] ;
 wire \ring_1001.inv_in[476] ;
 wire \ring_1001.inv_in[477] ;
 wire \ring_1001.inv_in[478] ;
 wire \ring_1001.inv_in[479] ;
 wire \ring_1001.inv_in[47] ;
 wire \ring_1001.inv_in[480] ;
 wire \ring_1001.inv_in[481] ;
 wire \ring_1001.inv_in[482] ;
 wire \ring_1001.inv_in[483] ;
 wire \ring_1001.inv_in[484] ;
 wire \ring_1001.inv_in[485] ;
 wire \ring_1001.inv_in[486] ;
 wire \ring_1001.inv_in[487] ;
 wire \ring_1001.inv_in[488] ;
 wire \ring_1001.inv_in[489] ;
 wire \ring_1001.inv_in[48] ;
 wire \ring_1001.inv_in[490] ;
 wire \ring_1001.inv_in[491] ;
 wire \ring_1001.inv_in[492] ;
 wire \ring_1001.inv_in[493] ;
 wire \ring_1001.inv_in[494] ;
 wire \ring_1001.inv_in[495] ;
 wire \ring_1001.inv_in[496] ;
 wire \ring_1001.inv_in[497] ;
 wire \ring_1001.inv_in[498] ;
 wire \ring_1001.inv_in[499] ;
 wire \ring_1001.inv_in[49] ;
 wire \ring_1001.inv_in[4] ;
 wire \ring_1001.inv_in[500] ;
 wire \ring_1001.inv_in[501] ;
 wire \ring_1001.inv_in[502] ;
 wire \ring_1001.inv_in[503] ;
 wire \ring_1001.inv_in[504] ;
 wire \ring_1001.inv_in[505] ;
 wire \ring_1001.inv_in[506] ;
 wire \ring_1001.inv_in[507] ;
 wire \ring_1001.inv_in[508] ;
 wire \ring_1001.inv_in[509] ;
 wire \ring_1001.inv_in[50] ;
 wire \ring_1001.inv_in[510] ;
 wire \ring_1001.inv_in[511] ;
 wire \ring_1001.inv_in[512] ;
 wire \ring_1001.inv_in[513] ;
 wire \ring_1001.inv_in[514] ;
 wire \ring_1001.inv_in[515] ;
 wire \ring_1001.inv_in[516] ;
 wire \ring_1001.inv_in[517] ;
 wire \ring_1001.inv_in[518] ;
 wire \ring_1001.inv_in[519] ;
 wire \ring_1001.inv_in[51] ;
 wire \ring_1001.inv_in[520] ;
 wire \ring_1001.inv_in[521] ;
 wire \ring_1001.inv_in[522] ;
 wire \ring_1001.inv_in[523] ;
 wire \ring_1001.inv_in[524] ;
 wire \ring_1001.inv_in[525] ;
 wire \ring_1001.inv_in[526] ;
 wire \ring_1001.inv_in[527] ;
 wire \ring_1001.inv_in[528] ;
 wire \ring_1001.inv_in[529] ;
 wire \ring_1001.inv_in[52] ;
 wire \ring_1001.inv_in[530] ;
 wire \ring_1001.inv_in[531] ;
 wire \ring_1001.inv_in[532] ;
 wire \ring_1001.inv_in[533] ;
 wire \ring_1001.inv_in[534] ;
 wire \ring_1001.inv_in[535] ;
 wire \ring_1001.inv_in[536] ;
 wire \ring_1001.inv_in[537] ;
 wire \ring_1001.inv_in[538] ;
 wire \ring_1001.inv_in[539] ;
 wire \ring_1001.inv_in[53] ;
 wire \ring_1001.inv_in[540] ;
 wire \ring_1001.inv_in[541] ;
 wire \ring_1001.inv_in[542] ;
 wire \ring_1001.inv_in[543] ;
 wire \ring_1001.inv_in[544] ;
 wire \ring_1001.inv_in[545] ;
 wire \ring_1001.inv_in[546] ;
 wire \ring_1001.inv_in[547] ;
 wire \ring_1001.inv_in[548] ;
 wire \ring_1001.inv_in[549] ;
 wire \ring_1001.inv_in[54] ;
 wire \ring_1001.inv_in[550] ;
 wire \ring_1001.inv_in[551] ;
 wire \ring_1001.inv_in[552] ;
 wire \ring_1001.inv_in[553] ;
 wire \ring_1001.inv_in[554] ;
 wire \ring_1001.inv_in[555] ;
 wire \ring_1001.inv_in[556] ;
 wire \ring_1001.inv_in[557] ;
 wire \ring_1001.inv_in[558] ;
 wire \ring_1001.inv_in[559] ;
 wire \ring_1001.inv_in[55] ;
 wire \ring_1001.inv_in[560] ;
 wire \ring_1001.inv_in[561] ;
 wire \ring_1001.inv_in[562] ;
 wire \ring_1001.inv_in[563] ;
 wire \ring_1001.inv_in[564] ;
 wire \ring_1001.inv_in[565] ;
 wire \ring_1001.inv_in[566] ;
 wire \ring_1001.inv_in[567] ;
 wire \ring_1001.inv_in[568] ;
 wire \ring_1001.inv_in[569] ;
 wire \ring_1001.inv_in[56] ;
 wire \ring_1001.inv_in[570] ;
 wire \ring_1001.inv_in[571] ;
 wire \ring_1001.inv_in[572] ;
 wire \ring_1001.inv_in[573] ;
 wire \ring_1001.inv_in[574] ;
 wire \ring_1001.inv_in[575] ;
 wire \ring_1001.inv_in[576] ;
 wire \ring_1001.inv_in[577] ;
 wire \ring_1001.inv_in[578] ;
 wire \ring_1001.inv_in[579] ;
 wire \ring_1001.inv_in[57] ;
 wire \ring_1001.inv_in[580] ;
 wire \ring_1001.inv_in[581] ;
 wire \ring_1001.inv_in[582] ;
 wire \ring_1001.inv_in[583] ;
 wire \ring_1001.inv_in[584] ;
 wire \ring_1001.inv_in[585] ;
 wire \ring_1001.inv_in[586] ;
 wire \ring_1001.inv_in[587] ;
 wire \ring_1001.inv_in[588] ;
 wire \ring_1001.inv_in[589] ;
 wire \ring_1001.inv_in[58] ;
 wire \ring_1001.inv_in[590] ;
 wire \ring_1001.inv_in[591] ;
 wire \ring_1001.inv_in[592] ;
 wire \ring_1001.inv_in[593] ;
 wire \ring_1001.inv_in[594] ;
 wire \ring_1001.inv_in[595] ;
 wire \ring_1001.inv_in[596] ;
 wire \ring_1001.inv_in[597] ;
 wire \ring_1001.inv_in[598] ;
 wire \ring_1001.inv_in[599] ;
 wire \ring_1001.inv_in[59] ;
 wire \ring_1001.inv_in[5] ;
 wire \ring_1001.inv_in[600] ;
 wire \ring_1001.inv_in[601] ;
 wire \ring_1001.inv_in[602] ;
 wire \ring_1001.inv_in[603] ;
 wire \ring_1001.inv_in[604] ;
 wire \ring_1001.inv_in[605] ;
 wire \ring_1001.inv_in[606] ;
 wire \ring_1001.inv_in[607] ;
 wire \ring_1001.inv_in[608] ;
 wire \ring_1001.inv_in[609] ;
 wire \ring_1001.inv_in[60] ;
 wire \ring_1001.inv_in[610] ;
 wire \ring_1001.inv_in[611] ;
 wire \ring_1001.inv_in[612] ;
 wire \ring_1001.inv_in[613] ;
 wire \ring_1001.inv_in[614] ;
 wire \ring_1001.inv_in[615] ;
 wire \ring_1001.inv_in[616] ;
 wire \ring_1001.inv_in[617] ;
 wire \ring_1001.inv_in[618] ;
 wire \ring_1001.inv_in[619] ;
 wire \ring_1001.inv_in[61] ;
 wire \ring_1001.inv_in[620] ;
 wire \ring_1001.inv_in[621] ;
 wire \ring_1001.inv_in[622] ;
 wire \ring_1001.inv_in[623] ;
 wire \ring_1001.inv_in[624] ;
 wire \ring_1001.inv_in[625] ;
 wire \ring_1001.inv_in[626] ;
 wire \ring_1001.inv_in[627] ;
 wire \ring_1001.inv_in[628] ;
 wire \ring_1001.inv_in[629] ;
 wire \ring_1001.inv_in[62] ;
 wire \ring_1001.inv_in[630] ;
 wire \ring_1001.inv_in[631] ;
 wire \ring_1001.inv_in[632] ;
 wire \ring_1001.inv_in[633] ;
 wire \ring_1001.inv_in[634] ;
 wire \ring_1001.inv_in[635] ;
 wire \ring_1001.inv_in[636] ;
 wire \ring_1001.inv_in[637] ;
 wire \ring_1001.inv_in[638] ;
 wire \ring_1001.inv_in[639] ;
 wire \ring_1001.inv_in[63] ;
 wire \ring_1001.inv_in[640] ;
 wire \ring_1001.inv_in[641] ;
 wire \ring_1001.inv_in[642] ;
 wire \ring_1001.inv_in[643] ;
 wire \ring_1001.inv_in[644] ;
 wire \ring_1001.inv_in[645] ;
 wire \ring_1001.inv_in[646] ;
 wire \ring_1001.inv_in[647] ;
 wire \ring_1001.inv_in[648] ;
 wire \ring_1001.inv_in[649] ;
 wire \ring_1001.inv_in[64] ;
 wire \ring_1001.inv_in[650] ;
 wire \ring_1001.inv_in[651] ;
 wire \ring_1001.inv_in[652] ;
 wire \ring_1001.inv_in[653] ;
 wire \ring_1001.inv_in[654] ;
 wire \ring_1001.inv_in[655] ;
 wire \ring_1001.inv_in[656] ;
 wire \ring_1001.inv_in[657] ;
 wire \ring_1001.inv_in[658] ;
 wire \ring_1001.inv_in[659] ;
 wire \ring_1001.inv_in[65] ;
 wire \ring_1001.inv_in[660] ;
 wire \ring_1001.inv_in[661] ;
 wire \ring_1001.inv_in[662] ;
 wire \ring_1001.inv_in[663] ;
 wire \ring_1001.inv_in[664] ;
 wire \ring_1001.inv_in[665] ;
 wire \ring_1001.inv_in[666] ;
 wire \ring_1001.inv_in[667] ;
 wire \ring_1001.inv_in[668] ;
 wire \ring_1001.inv_in[669] ;
 wire \ring_1001.inv_in[66] ;
 wire \ring_1001.inv_in[670] ;
 wire \ring_1001.inv_in[671] ;
 wire \ring_1001.inv_in[672] ;
 wire \ring_1001.inv_in[673] ;
 wire \ring_1001.inv_in[674] ;
 wire \ring_1001.inv_in[675] ;
 wire \ring_1001.inv_in[676] ;
 wire \ring_1001.inv_in[677] ;
 wire \ring_1001.inv_in[678] ;
 wire \ring_1001.inv_in[679] ;
 wire \ring_1001.inv_in[67] ;
 wire \ring_1001.inv_in[680] ;
 wire \ring_1001.inv_in[681] ;
 wire \ring_1001.inv_in[682] ;
 wire \ring_1001.inv_in[683] ;
 wire \ring_1001.inv_in[684] ;
 wire \ring_1001.inv_in[685] ;
 wire \ring_1001.inv_in[686] ;
 wire \ring_1001.inv_in[687] ;
 wire \ring_1001.inv_in[688] ;
 wire \ring_1001.inv_in[689] ;
 wire \ring_1001.inv_in[68] ;
 wire \ring_1001.inv_in[690] ;
 wire \ring_1001.inv_in[691] ;
 wire \ring_1001.inv_in[692] ;
 wire \ring_1001.inv_in[693] ;
 wire \ring_1001.inv_in[694] ;
 wire \ring_1001.inv_in[695] ;
 wire \ring_1001.inv_in[696] ;
 wire \ring_1001.inv_in[697] ;
 wire \ring_1001.inv_in[698] ;
 wire \ring_1001.inv_in[699] ;
 wire \ring_1001.inv_in[69] ;
 wire \ring_1001.inv_in[6] ;
 wire \ring_1001.inv_in[700] ;
 wire \ring_1001.inv_in[701] ;
 wire \ring_1001.inv_in[702] ;
 wire \ring_1001.inv_in[703] ;
 wire \ring_1001.inv_in[704] ;
 wire \ring_1001.inv_in[705] ;
 wire \ring_1001.inv_in[706] ;
 wire \ring_1001.inv_in[707] ;
 wire \ring_1001.inv_in[708] ;
 wire \ring_1001.inv_in[709] ;
 wire \ring_1001.inv_in[70] ;
 wire \ring_1001.inv_in[710] ;
 wire \ring_1001.inv_in[711] ;
 wire \ring_1001.inv_in[712] ;
 wire \ring_1001.inv_in[713] ;
 wire \ring_1001.inv_in[714] ;
 wire \ring_1001.inv_in[715] ;
 wire \ring_1001.inv_in[716] ;
 wire \ring_1001.inv_in[717] ;
 wire \ring_1001.inv_in[718] ;
 wire \ring_1001.inv_in[719] ;
 wire \ring_1001.inv_in[71] ;
 wire \ring_1001.inv_in[720] ;
 wire \ring_1001.inv_in[721] ;
 wire \ring_1001.inv_in[722] ;
 wire \ring_1001.inv_in[723] ;
 wire \ring_1001.inv_in[724] ;
 wire \ring_1001.inv_in[725] ;
 wire \ring_1001.inv_in[726] ;
 wire \ring_1001.inv_in[727] ;
 wire \ring_1001.inv_in[728] ;
 wire \ring_1001.inv_in[729] ;
 wire \ring_1001.inv_in[72] ;
 wire \ring_1001.inv_in[730] ;
 wire \ring_1001.inv_in[731] ;
 wire \ring_1001.inv_in[732] ;
 wire \ring_1001.inv_in[733] ;
 wire \ring_1001.inv_in[734] ;
 wire \ring_1001.inv_in[735] ;
 wire \ring_1001.inv_in[736] ;
 wire \ring_1001.inv_in[737] ;
 wire \ring_1001.inv_in[738] ;
 wire \ring_1001.inv_in[739] ;
 wire \ring_1001.inv_in[73] ;
 wire \ring_1001.inv_in[740] ;
 wire \ring_1001.inv_in[741] ;
 wire \ring_1001.inv_in[742] ;
 wire \ring_1001.inv_in[743] ;
 wire \ring_1001.inv_in[744] ;
 wire \ring_1001.inv_in[745] ;
 wire \ring_1001.inv_in[746] ;
 wire \ring_1001.inv_in[747] ;
 wire \ring_1001.inv_in[748] ;
 wire \ring_1001.inv_in[749] ;
 wire \ring_1001.inv_in[74] ;
 wire \ring_1001.inv_in[750] ;
 wire \ring_1001.inv_in[751] ;
 wire \ring_1001.inv_in[752] ;
 wire \ring_1001.inv_in[753] ;
 wire \ring_1001.inv_in[754] ;
 wire \ring_1001.inv_in[755] ;
 wire \ring_1001.inv_in[756] ;
 wire \ring_1001.inv_in[757] ;
 wire \ring_1001.inv_in[758] ;
 wire \ring_1001.inv_in[759] ;
 wire \ring_1001.inv_in[75] ;
 wire \ring_1001.inv_in[760] ;
 wire \ring_1001.inv_in[761] ;
 wire \ring_1001.inv_in[762] ;
 wire \ring_1001.inv_in[763] ;
 wire \ring_1001.inv_in[764] ;
 wire \ring_1001.inv_in[765] ;
 wire \ring_1001.inv_in[766] ;
 wire \ring_1001.inv_in[767] ;
 wire \ring_1001.inv_in[768] ;
 wire \ring_1001.inv_in[769] ;
 wire \ring_1001.inv_in[76] ;
 wire \ring_1001.inv_in[770] ;
 wire \ring_1001.inv_in[771] ;
 wire \ring_1001.inv_in[772] ;
 wire \ring_1001.inv_in[773] ;
 wire \ring_1001.inv_in[774] ;
 wire \ring_1001.inv_in[775] ;
 wire \ring_1001.inv_in[776] ;
 wire \ring_1001.inv_in[777] ;
 wire \ring_1001.inv_in[778] ;
 wire \ring_1001.inv_in[779] ;
 wire \ring_1001.inv_in[77] ;
 wire \ring_1001.inv_in[780] ;
 wire \ring_1001.inv_in[781] ;
 wire \ring_1001.inv_in[782] ;
 wire \ring_1001.inv_in[783] ;
 wire \ring_1001.inv_in[784] ;
 wire \ring_1001.inv_in[785] ;
 wire \ring_1001.inv_in[786] ;
 wire \ring_1001.inv_in[787] ;
 wire \ring_1001.inv_in[788] ;
 wire \ring_1001.inv_in[789] ;
 wire \ring_1001.inv_in[78] ;
 wire \ring_1001.inv_in[790] ;
 wire \ring_1001.inv_in[791] ;
 wire \ring_1001.inv_in[792] ;
 wire \ring_1001.inv_in[793] ;
 wire \ring_1001.inv_in[794] ;
 wire \ring_1001.inv_in[795] ;
 wire \ring_1001.inv_in[796] ;
 wire \ring_1001.inv_in[797] ;
 wire \ring_1001.inv_in[798] ;
 wire \ring_1001.inv_in[799] ;
 wire \ring_1001.inv_in[79] ;
 wire \ring_1001.inv_in[7] ;
 wire \ring_1001.inv_in[800] ;
 wire \ring_1001.inv_in[801] ;
 wire \ring_1001.inv_in[802] ;
 wire \ring_1001.inv_in[803] ;
 wire \ring_1001.inv_in[804] ;
 wire \ring_1001.inv_in[805] ;
 wire \ring_1001.inv_in[806] ;
 wire \ring_1001.inv_in[807] ;
 wire \ring_1001.inv_in[808] ;
 wire \ring_1001.inv_in[809] ;
 wire \ring_1001.inv_in[80] ;
 wire \ring_1001.inv_in[810] ;
 wire \ring_1001.inv_in[811] ;
 wire \ring_1001.inv_in[812] ;
 wire \ring_1001.inv_in[813] ;
 wire \ring_1001.inv_in[814] ;
 wire \ring_1001.inv_in[815] ;
 wire \ring_1001.inv_in[816] ;
 wire \ring_1001.inv_in[817] ;
 wire \ring_1001.inv_in[818] ;
 wire \ring_1001.inv_in[819] ;
 wire \ring_1001.inv_in[81] ;
 wire \ring_1001.inv_in[820] ;
 wire \ring_1001.inv_in[821] ;
 wire \ring_1001.inv_in[822] ;
 wire \ring_1001.inv_in[823] ;
 wire \ring_1001.inv_in[824] ;
 wire \ring_1001.inv_in[825] ;
 wire \ring_1001.inv_in[826] ;
 wire \ring_1001.inv_in[827] ;
 wire \ring_1001.inv_in[828] ;
 wire \ring_1001.inv_in[829] ;
 wire \ring_1001.inv_in[82] ;
 wire \ring_1001.inv_in[830] ;
 wire \ring_1001.inv_in[831] ;
 wire \ring_1001.inv_in[832] ;
 wire \ring_1001.inv_in[833] ;
 wire \ring_1001.inv_in[834] ;
 wire \ring_1001.inv_in[835] ;
 wire \ring_1001.inv_in[836] ;
 wire \ring_1001.inv_in[837] ;
 wire \ring_1001.inv_in[838] ;
 wire \ring_1001.inv_in[839] ;
 wire \ring_1001.inv_in[83] ;
 wire \ring_1001.inv_in[840] ;
 wire \ring_1001.inv_in[841] ;
 wire \ring_1001.inv_in[842] ;
 wire \ring_1001.inv_in[843] ;
 wire \ring_1001.inv_in[844] ;
 wire \ring_1001.inv_in[845] ;
 wire \ring_1001.inv_in[846] ;
 wire \ring_1001.inv_in[847] ;
 wire \ring_1001.inv_in[848] ;
 wire \ring_1001.inv_in[849] ;
 wire \ring_1001.inv_in[84] ;
 wire \ring_1001.inv_in[850] ;
 wire \ring_1001.inv_in[851] ;
 wire \ring_1001.inv_in[852] ;
 wire \ring_1001.inv_in[853] ;
 wire \ring_1001.inv_in[854] ;
 wire \ring_1001.inv_in[855] ;
 wire \ring_1001.inv_in[856] ;
 wire \ring_1001.inv_in[857] ;
 wire \ring_1001.inv_in[858] ;
 wire \ring_1001.inv_in[859] ;
 wire \ring_1001.inv_in[85] ;
 wire \ring_1001.inv_in[860] ;
 wire \ring_1001.inv_in[861] ;
 wire \ring_1001.inv_in[862] ;
 wire \ring_1001.inv_in[863] ;
 wire \ring_1001.inv_in[864] ;
 wire \ring_1001.inv_in[865] ;
 wire \ring_1001.inv_in[866] ;
 wire \ring_1001.inv_in[867] ;
 wire \ring_1001.inv_in[868] ;
 wire \ring_1001.inv_in[869] ;
 wire \ring_1001.inv_in[86] ;
 wire \ring_1001.inv_in[870] ;
 wire \ring_1001.inv_in[871] ;
 wire \ring_1001.inv_in[872] ;
 wire \ring_1001.inv_in[873] ;
 wire \ring_1001.inv_in[874] ;
 wire \ring_1001.inv_in[875] ;
 wire \ring_1001.inv_in[876] ;
 wire \ring_1001.inv_in[877] ;
 wire \ring_1001.inv_in[878] ;
 wire \ring_1001.inv_in[879] ;
 wire \ring_1001.inv_in[87] ;
 wire \ring_1001.inv_in[880] ;
 wire \ring_1001.inv_in[881] ;
 wire \ring_1001.inv_in[882] ;
 wire \ring_1001.inv_in[883] ;
 wire \ring_1001.inv_in[884] ;
 wire \ring_1001.inv_in[885] ;
 wire \ring_1001.inv_in[886] ;
 wire \ring_1001.inv_in[887] ;
 wire \ring_1001.inv_in[888] ;
 wire \ring_1001.inv_in[889] ;
 wire \ring_1001.inv_in[88] ;
 wire \ring_1001.inv_in[890] ;
 wire \ring_1001.inv_in[891] ;
 wire \ring_1001.inv_in[892] ;
 wire \ring_1001.inv_in[893] ;
 wire \ring_1001.inv_in[894] ;
 wire \ring_1001.inv_in[895] ;
 wire \ring_1001.inv_in[896] ;
 wire \ring_1001.inv_in[897] ;
 wire \ring_1001.inv_in[898] ;
 wire \ring_1001.inv_in[899] ;
 wire \ring_1001.inv_in[89] ;
 wire \ring_1001.inv_in[8] ;
 wire \ring_1001.inv_in[900] ;
 wire \ring_1001.inv_in[901] ;
 wire \ring_1001.inv_in[902] ;
 wire \ring_1001.inv_in[903] ;
 wire \ring_1001.inv_in[904] ;
 wire \ring_1001.inv_in[905] ;
 wire \ring_1001.inv_in[906] ;
 wire \ring_1001.inv_in[907] ;
 wire \ring_1001.inv_in[908] ;
 wire \ring_1001.inv_in[909] ;
 wire \ring_1001.inv_in[90] ;
 wire \ring_1001.inv_in[910] ;
 wire \ring_1001.inv_in[911] ;
 wire \ring_1001.inv_in[912] ;
 wire \ring_1001.inv_in[913] ;
 wire \ring_1001.inv_in[914] ;
 wire \ring_1001.inv_in[915] ;
 wire \ring_1001.inv_in[916] ;
 wire \ring_1001.inv_in[917] ;
 wire \ring_1001.inv_in[918] ;
 wire \ring_1001.inv_in[919] ;
 wire \ring_1001.inv_in[91] ;
 wire \ring_1001.inv_in[920] ;
 wire \ring_1001.inv_in[921] ;
 wire \ring_1001.inv_in[922] ;
 wire \ring_1001.inv_in[923] ;
 wire \ring_1001.inv_in[924] ;
 wire \ring_1001.inv_in[925] ;
 wire \ring_1001.inv_in[926] ;
 wire \ring_1001.inv_in[927] ;
 wire \ring_1001.inv_in[928] ;
 wire \ring_1001.inv_in[929] ;
 wire \ring_1001.inv_in[92] ;
 wire \ring_1001.inv_in[930] ;
 wire \ring_1001.inv_in[931] ;
 wire \ring_1001.inv_in[932] ;
 wire \ring_1001.inv_in[933] ;
 wire \ring_1001.inv_in[934] ;
 wire \ring_1001.inv_in[935] ;
 wire \ring_1001.inv_in[936] ;
 wire \ring_1001.inv_in[937] ;
 wire \ring_1001.inv_in[938] ;
 wire \ring_1001.inv_in[939] ;
 wire \ring_1001.inv_in[93] ;
 wire \ring_1001.inv_in[940] ;
 wire \ring_1001.inv_in[941] ;
 wire \ring_1001.inv_in[942] ;
 wire \ring_1001.inv_in[943] ;
 wire \ring_1001.inv_in[944] ;
 wire \ring_1001.inv_in[945] ;
 wire \ring_1001.inv_in[946] ;
 wire \ring_1001.inv_in[947] ;
 wire \ring_1001.inv_in[948] ;
 wire \ring_1001.inv_in[949] ;
 wire \ring_1001.inv_in[94] ;
 wire \ring_1001.inv_in[950] ;
 wire \ring_1001.inv_in[951] ;
 wire \ring_1001.inv_in[952] ;
 wire \ring_1001.inv_in[953] ;
 wire \ring_1001.inv_in[954] ;
 wire \ring_1001.inv_in[955] ;
 wire \ring_1001.inv_in[956] ;
 wire \ring_1001.inv_in[957] ;
 wire \ring_1001.inv_in[958] ;
 wire \ring_1001.inv_in[959] ;
 wire \ring_1001.inv_in[95] ;
 wire \ring_1001.inv_in[960] ;
 wire \ring_1001.inv_in[961] ;
 wire \ring_1001.inv_in[962] ;
 wire \ring_1001.inv_in[963] ;
 wire \ring_1001.inv_in[964] ;
 wire \ring_1001.inv_in[965] ;
 wire \ring_1001.inv_in[966] ;
 wire \ring_1001.inv_in[967] ;
 wire \ring_1001.inv_in[968] ;
 wire \ring_1001.inv_in[969] ;
 wire \ring_1001.inv_in[96] ;
 wire \ring_1001.inv_in[970] ;
 wire \ring_1001.inv_in[971] ;
 wire \ring_1001.inv_in[972] ;
 wire \ring_1001.inv_in[973] ;
 wire \ring_1001.inv_in[974] ;
 wire \ring_1001.inv_in[975] ;
 wire \ring_1001.inv_in[976] ;
 wire \ring_1001.inv_in[977] ;
 wire \ring_1001.inv_in[978] ;
 wire \ring_1001.inv_in[979] ;
 wire \ring_1001.inv_in[97] ;
 wire \ring_1001.inv_in[980] ;
 wire \ring_1001.inv_in[981] ;
 wire \ring_1001.inv_in[982] ;
 wire \ring_1001.inv_in[983] ;
 wire \ring_1001.inv_in[984] ;
 wire \ring_1001.inv_in[985] ;
 wire \ring_1001.inv_in[986] ;
 wire \ring_1001.inv_in[987] ;
 wire \ring_1001.inv_in[988] ;
 wire \ring_1001.inv_in[989] ;
 wire \ring_1001.inv_in[98] ;
 wire \ring_1001.inv_in[990] ;
 wire \ring_1001.inv_in[991] ;
 wire \ring_1001.inv_in[992] ;
 wire \ring_1001.inv_in[993] ;
 wire \ring_1001.inv_in[994] ;
 wire \ring_1001.inv_in[995] ;
 wire \ring_1001.inv_in[996] ;
 wire \ring_1001.inv_in[997] ;
 wire \ring_1001.inv_in[998] ;
 wire \ring_1001.inv_in[999] ;
 wire \ring_1001.inv_in[99] ;
 wire \ring_1001.inv_in[9] ;
 wire \ring_1001.inv_out[1000] ;
 wire \ring_125.inv_in[100] ;
 wire \ring_125.inv_in[101] ;
 wire \ring_125.inv_in[102] ;
 wire \ring_125.inv_in[103] ;
 wire \ring_125.inv_in[104] ;
 wire \ring_125.inv_in[105] ;
 wire \ring_125.inv_in[106] ;
 wire \ring_125.inv_in[107] ;
 wire \ring_125.inv_in[108] ;
 wire \ring_125.inv_in[109] ;
 wire \ring_125.inv_in[10] ;
 wire \ring_125.inv_in[110] ;
 wire \ring_125.inv_in[111] ;
 wire \ring_125.inv_in[112] ;
 wire \ring_125.inv_in[113] ;
 wire \ring_125.inv_in[114] ;
 wire \ring_125.inv_in[115] ;
 wire \ring_125.inv_in[116] ;
 wire \ring_125.inv_in[117] ;
 wire \ring_125.inv_in[118] ;
 wire \ring_125.inv_in[119] ;
 wire \ring_125.inv_in[11] ;
 wire \ring_125.inv_in[120] ;
 wire \ring_125.inv_in[121] ;
 wire \ring_125.inv_in[122] ;
 wire \ring_125.inv_in[123] ;
 wire \ring_125.inv_in[124] ;
 wire \ring_125.inv_in[12] ;
 wire \ring_125.inv_in[13] ;
 wire \ring_125.inv_in[14] ;
 wire \ring_125.inv_in[15] ;
 wire \ring_125.inv_in[16] ;
 wire \ring_125.inv_in[17] ;
 wire \ring_125.inv_in[18] ;
 wire \ring_125.inv_in[19] ;
 wire \ring_125.inv_in[1] ;
 wire \ring_125.inv_in[20] ;
 wire \ring_125.inv_in[21] ;
 wire \ring_125.inv_in[22] ;
 wire \ring_125.inv_in[23] ;
 wire \ring_125.inv_in[24] ;
 wire \ring_125.inv_in[25] ;
 wire \ring_125.inv_in[26] ;
 wire \ring_125.inv_in[27] ;
 wire \ring_125.inv_in[28] ;
 wire \ring_125.inv_in[29] ;
 wire \ring_125.inv_in[2] ;
 wire \ring_125.inv_in[30] ;
 wire \ring_125.inv_in[31] ;
 wire \ring_125.inv_in[32] ;
 wire \ring_125.inv_in[33] ;
 wire \ring_125.inv_in[34] ;
 wire \ring_125.inv_in[35] ;
 wire \ring_125.inv_in[36] ;
 wire \ring_125.inv_in[37] ;
 wire \ring_125.inv_in[38] ;
 wire \ring_125.inv_in[39] ;
 wire \ring_125.inv_in[3] ;
 wire \ring_125.inv_in[40] ;
 wire \ring_125.inv_in[41] ;
 wire \ring_125.inv_in[42] ;
 wire \ring_125.inv_in[43] ;
 wire \ring_125.inv_in[44] ;
 wire \ring_125.inv_in[45] ;
 wire \ring_125.inv_in[46] ;
 wire \ring_125.inv_in[47] ;
 wire \ring_125.inv_in[48] ;
 wire \ring_125.inv_in[49] ;
 wire \ring_125.inv_in[4] ;
 wire \ring_125.inv_in[50] ;
 wire \ring_125.inv_in[51] ;
 wire \ring_125.inv_in[52] ;
 wire \ring_125.inv_in[53] ;
 wire \ring_125.inv_in[54] ;
 wire \ring_125.inv_in[55] ;
 wire \ring_125.inv_in[56] ;
 wire \ring_125.inv_in[57] ;
 wire \ring_125.inv_in[58] ;
 wire \ring_125.inv_in[59] ;
 wire \ring_125.inv_in[5] ;
 wire \ring_125.inv_in[60] ;
 wire \ring_125.inv_in[61] ;
 wire \ring_125.inv_in[62] ;
 wire \ring_125.inv_in[63] ;
 wire \ring_125.inv_in[64] ;
 wire \ring_125.inv_in[65] ;
 wire \ring_125.inv_in[66] ;
 wire \ring_125.inv_in[67] ;
 wire \ring_125.inv_in[68] ;
 wire \ring_125.inv_in[69] ;
 wire \ring_125.inv_in[6] ;
 wire \ring_125.inv_in[70] ;
 wire \ring_125.inv_in[71] ;
 wire \ring_125.inv_in[72] ;
 wire \ring_125.inv_in[73] ;
 wire \ring_125.inv_in[74] ;
 wire \ring_125.inv_in[75] ;
 wire \ring_125.inv_in[76] ;
 wire \ring_125.inv_in[77] ;
 wire \ring_125.inv_in[78] ;
 wire \ring_125.inv_in[79] ;
 wire \ring_125.inv_in[7] ;
 wire \ring_125.inv_in[80] ;
 wire \ring_125.inv_in[81] ;
 wire \ring_125.inv_in[82] ;
 wire \ring_125.inv_in[83] ;
 wire \ring_125.inv_in[84] ;
 wire \ring_125.inv_in[85] ;
 wire \ring_125.inv_in[86] ;
 wire \ring_125.inv_in[87] ;
 wire \ring_125.inv_in[88] ;
 wire \ring_125.inv_in[89] ;
 wire \ring_125.inv_in[8] ;
 wire \ring_125.inv_in[90] ;
 wire \ring_125.inv_in[91] ;
 wire \ring_125.inv_in[92] ;
 wire \ring_125.inv_in[93] ;
 wire \ring_125.inv_in[94] ;
 wire \ring_125.inv_in[95] ;
 wire \ring_125.inv_in[96] ;
 wire \ring_125.inv_in[97] ;
 wire \ring_125.inv_in[98] ;
 wire \ring_125.inv_in[99] ;
 wire \ring_125.inv_in[9] ;
 wire \ring_125.inv_out[124] ;
 wire \ring_25.inv_in[10] ;
 wire \ring_25.inv_in[11] ;
 wire \ring_25.inv_in[12] ;
 wire \ring_25.inv_in[13] ;
 wire \ring_25.inv_in[14] ;
 wire \ring_25.inv_in[15] ;
 wire \ring_25.inv_in[16] ;
 wire \ring_25.inv_in[17] ;
 wire \ring_25.inv_in[18] ;
 wire \ring_25.inv_in[19] ;
 wire \ring_25.inv_in[1] ;
 wire \ring_25.inv_in[20] ;
 wire \ring_25.inv_in[21] ;
 wire \ring_25.inv_in[22] ;
 wire \ring_25.inv_in[23] ;
 wire \ring_25.inv_in[24] ;
 wire \ring_25.inv_in[2] ;
 wire \ring_25.inv_in[3] ;
 wire \ring_25.inv_in[4] ;
 wire \ring_25.inv_in[5] ;
 wire \ring_25.inv_in[6] ;
 wire \ring_25.inv_in[7] ;
 wire \ring_25.inv_in[8] ;
 wire \ring_25.inv_in[9] ;
 wire \ring_25.inv_out[24] ;
 wire \ring_251.inv_in[0] ;
 wire \ring_251.inv_in[100] ;
 wire \ring_251.inv_in[101] ;
 wire \ring_251.inv_in[102] ;
 wire \ring_251.inv_in[103] ;
 wire \ring_251.inv_in[104] ;
 wire \ring_251.inv_in[105] ;
 wire \ring_251.inv_in[106] ;
 wire \ring_251.inv_in[107] ;
 wire \ring_251.inv_in[108] ;
 wire \ring_251.inv_in[109] ;
 wire \ring_251.inv_in[10] ;
 wire \ring_251.inv_in[110] ;
 wire \ring_251.inv_in[111] ;
 wire \ring_251.inv_in[112] ;
 wire \ring_251.inv_in[113] ;
 wire \ring_251.inv_in[114] ;
 wire \ring_251.inv_in[115] ;
 wire \ring_251.inv_in[116] ;
 wire \ring_251.inv_in[117] ;
 wire \ring_251.inv_in[118] ;
 wire \ring_251.inv_in[119] ;
 wire \ring_251.inv_in[11] ;
 wire \ring_251.inv_in[120] ;
 wire \ring_251.inv_in[121] ;
 wire \ring_251.inv_in[122] ;
 wire \ring_251.inv_in[123] ;
 wire \ring_251.inv_in[124] ;
 wire \ring_251.inv_in[125] ;
 wire \ring_251.inv_in[126] ;
 wire \ring_251.inv_in[127] ;
 wire \ring_251.inv_in[128] ;
 wire \ring_251.inv_in[129] ;
 wire \ring_251.inv_in[12] ;
 wire \ring_251.inv_in[130] ;
 wire \ring_251.inv_in[131] ;
 wire \ring_251.inv_in[132] ;
 wire \ring_251.inv_in[133] ;
 wire \ring_251.inv_in[134] ;
 wire \ring_251.inv_in[135] ;
 wire \ring_251.inv_in[136] ;
 wire \ring_251.inv_in[137] ;
 wire \ring_251.inv_in[138] ;
 wire \ring_251.inv_in[139] ;
 wire \ring_251.inv_in[13] ;
 wire \ring_251.inv_in[140] ;
 wire \ring_251.inv_in[141] ;
 wire \ring_251.inv_in[142] ;
 wire \ring_251.inv_in[143] ;
 wire \ring_251.inv_in[144] ;
 wire \ring_251.inv_in[145] ;
 wire \ring_251.inv_in[146] ;
 wire \ring_251.inv_in[147] ;
 wire \ring_251.inv_in[148] ;
 wire \ring_251.inv_in[149] ;
 wire \ring_251.inv_in[14] ;
 wire \ring_251.inv_in[150] ;
 wire \ring_251.inv_in[151] ;
 wire \ring_251.inv_in[152] ;
 wire \ring_251.inv_in[153] ;
 wire \ring_251.inv_in[154] ;
 wire \ring_251.inv_in[155] ;
 wire \ring_251.inv_in[156] ;
 wire \ring_251.inv_in[157] ;
 wire \ring_251.inv_in[158] ;
 wire \ring_251.inv_in[159] ;
 wire \ring_251.inv_in[15] ;
 wire \ring_251.inv_in[160] ;
 wire \ring_251.inv_in[161] ;
 wire \ring_251.inv_in[162] ;
 wire \ring_251.inv_in[163] ;
 wire \ring_251.inv_in[164] ;
 wire \ring_251.inv_in[165] ;
 wire \ring_251.inv_in[166] ;
 wire \ring_251.inv_in[167] ;
 wire \ring_251.inv_in[168] ;
 wire \ring_251.inv_in[169] ;
 wire \ring_251.inv_in[16] ;
 wire \ring_251.inv_in[170] ;
 wire \ring_251.inv_in[171] ;
 wire \ring_251.inv_in[172] ;
 wire \ring_251.inv_in[173] ;
 wire \ring_251.inv_in[174] ;
 wire \ring_251.inv_in[175] ;
 wire \ring_251.inv_in[176] ;
 wire \ring_251.inv_in[177] ;
 wire \ring_251.inv_in[178] ;
 wire \ring_251.inv_in[179] ;
 wire \ring_251.inv_in[17] ;
 wire \ring_251.inv_in[180] ;
 wire \ring_251.inv_in[181] ;
 wire \ring_251.inv_in[182] ;
 wire \ring_251.inv_in[183] ;
 wire \ring_251.inv_in[184] ;
 wire \ring_251.inv_in[185] ;
 wire \ring_251.inv_in[186] ;
 wire \ring_251.inv_in[187] ;
 wire \ring_251.inv_in[188] ;
 wire \ring_251.inv_in[189] ;
 wire \ring_251.inv_in[18] ;
 wire \ring_251.inv_in[190] ;
 wire \ring_251.inv_in[191] ;
 wire \ring_251.inv_in[192] ;
 wire \ring_251.inv_in[193] ;
 wire \ring_251.inv_in[194] ;
 wire \ring_251.inv_in[195] ;
 wire \ring_251.inv_in[196] ;
 wire \ring_251.inv_in[197] ;
 wire \ring_251.inv_in[198] ;
 wire \ring_251.inv_in[199] ;
 wire \ring_251.inv_in[19] ;
 wire \ring_251.inv_in[1] ;
 wire \ring_251.inv_in[200] ;
 wire \ring_251.inv_in[201] ;
 wire \ring_251.inv_in[202] ;
 wire \ring_251.inv_in[203] ;
 wire \ring_251.inv_in[204] ;
 wire \ring_251.inv_in[205] ;
 wire \ring_251.inv_in[206] ;
 wire \ring_251.inv_in[207] ;
 wire \ring_251.inv_in[208] ;
 wire \ring_251.inv_in[209] ;
 wire \ring_251.inv_in[20] ;
 wire \ring_251.inv_in[210] ;
 wire \ring_251.inv_in[211] ;
 wire \ring_251.inv_in[212] ;
 wire \ring_251.inv_in[213] ;
 wire \ring_251.inv_in[214] ;
 wire \ring_251.inv_in[215] ;
 wire \ring_251.inv_in[216] ;
 wire \ring_251.inv_in[217] ;
 wire \ring_251.inv_in[218] ;
 wire \ring_251.inv_in[219] ;
 wire \ring_251.inv_in[21] ;
 wire \ring_251.inv_in[220] ;
 wire \ring_251.inv_in[221] ;
 wire \ring_251.inv_in[222] ;
 wire \ring_251.inv_in[223] ;
 wire \ring_251.inv_in[224] ;
 wire \ring_251.inv_in[225] ;
 wire \ring_251.inv_in[226] ;
 wire \ring_251.inv_in[227] ;
 wire \ring_251.inv_in[228] ;
 wire \ring_251.inv_in[229] ;
 wire \ring_251.inv_in[22] ;
 wire \ring_251.inv_in[230] ;
 wire \ring_251.inv_in[231] ;
 wire \ring_251.inv_in[232] ;
 wire \ring_251.inv_in[233] ;
 wire \ring_251.inv_in[234] ;
 wire \ring_251.inv_in[235] ;
 wire \ring_251.inv_in[236] ;
 wire \ring_251.inv_in[237] ;
 wire \ring_251.inv_in[238] ;
 wire \ring_251.inv_in[239] ;
 wire \ring_251.inv_in[23] ;
 wire \ring_251.inv_in[240] ;
 wire \ring_251.inv_in[241] ;
 wire \ring_251.inv_in[242] ;
 wire \ring_251.inv_in[243] ;
 wire \ring_251.inv_in[244] ;
 wire \ring_251.inv_in[245] ;
 wire \ring_251.inv_in[246] ;
 wire \ring_251.inv_in[247] ;
 wire \ring_251.inv_in[248] ;
 wire \ring_251.inv_in[249] ;
 wire \ring_251.inv_in[24] ;
 wire \ring_251.inv_in[250] ;
 wire \ring_251.inv_in[25] ;
 wire \ring_251.inv_in[26] ;
 wire \ring_251.inv_in[27] ;
 wire \ring_251.inv_in[28] ;
 wire \ring_251.inv_in[29] ;
 wire \ring_251.inv_in[2] ;
 wire \ring_251.inv_in[30] ;
 wire \ring_251.inv_in[31] ;
 wire \ring_251.inv_in[32] ;
 wire \ring_251.inv_in[33] ;
 wire \ring_251.inv_in[34] ;
 wire \ring_251.inv_in[35] ;
 wire \ring_251.inv_in[36] ;
 wire \ring_251.inv_in[37] ;
 wire \ring_251.inv_in[38] ;
 wire \ring_251.inv_in[39] ;
 wire \ring_251.inv_in[3] ;
 wire \ring_251.inv_in[40] ;
 wire \ring_251.inv_in[41] ;
 wire \ring_251.inv_in[42] ;
 wire \ring_251.inv_in[43] ;
 wire \ring_251.inv_in[44] ;
 wire \ring_251.inv_in[45] ;
 wire \ring_251.inv_in[46] ;
 wire \ring_251.inv_in[47] ;
 wire \ring_251.inv_in[48] ;
 wire \ring_251.inv_in[49] ;
 wire \ring_251.inv_in[4] ;
 wire \ring_251.inv_in[50] ;
 wire \ring_251.inv_in[51] ;
 wire \ring_251.inv_in[52] ;
 wire \ring_251.inv_in[53] ;
 wire \ring_251.inv_in[54] ;
 wire \ring_251.inv_in[55] ;
 wire \ring_251.inv_in[56] ;
 wire \ring_251.inv_in[57] ;
 wire \ring_251.inv_in[58] ;
 wire \ring_251.inv_in[59] ;
 wire \ring_251.inv_in[5] ;
 wire \ring_251.inv_in[60] ;
 wire \ring_251.inv_in[61] ;
 wire \ring_251.inv_in[62] ;
 wire \ring_251.inv_in[63] ;
 wire \ring_251.inv_in[64] ;
 wire \ring_251.inv_in[65] ;
 wire \ring_251.inv_in[66] ;
 wire \ring_251.inv_in[67] ;
 wire \ring_251.inv_in[68] ;
 wire \ring_251.inv_in[69] ;
 wire \ring_251.inv_in[6] ;
 wire \ring_251.inv_in[70] ;
 wire \ring_251.inv_in[71] ;
 wire \ring_251.inv_in[72] ;
 wire \ring_251.inv_in[73] ;
 wire \ring_251.inv_in[74] ;
 wire \ring_251.inv_in[75] ;
 wire \ring_251.inv_in[76] ;
 wire \ring_251.inv_in[77] ;
 wire \ring_251.inv_in[78] ;
 wire \ring_251.inv_in[79] ;
 wire \ring_251.inv_in[7] ;
 wire \ring_251.inv_in[80] ;
 wire \ring_251.inv_in[81] ;
 wire \ring_251.inv_in[82] ;
 wire \ring_251.inv_in[83] ;
 wire \ring_251.inv_in[84] ;
 wire \ring_251.inv_in[85] ;
 wire \ring_251.inv_in[86] ;
 wire \ring_251.inv_in[87] ;
 wire \ring_251.inv_in[88] ;
 wire \ring_251.inv_in[89] ;
 wire \ring_251.inv_in[8] ;
 wire \ring_251.inv_in[90] ;
 wire \ring_251.inv_in[91] ;
 wire \ring_251.inv_in[92] ;
 wire \ring_251.inv_in[93] ;
 wire \ring_251.inv_in[94] ;
 wire \ring_251.inv_in[95] ;
 wire \ring_251.inv_in[96] ;
 wire \ring_251.inv_in[97] ;
 wire \ring_251.inv_in[98] ;
 wire \ring_251.inv_in[99] ;
 wire \ring_251.inv_in[9] ;
 wire \ring_251.inv_out[250] ;
 wire \ring_501.inv_in[100] ;
 wire \ring_501.inv_in[101] ;
 wire \ring_501.inv_in[102] ;
 wire \ring_501.inv_in[103] ;
 wire \ring_501.inv_in[104] ;
 wire \ring_501.inv_in[105] ;
 wire \ring_501.inv_in[106] ;
 wire \ring_501.inv_in[107] ;
 wire \ring_501.inv_in[108] ;
 wire \ring_501.inv_in[109] ;
 wire \ring_501.inv_in[10] ;
 wire \ring_501.inv_in[110] ;
 wire \ring_501.inv_in[111] ;
 wire \ring_501.inv_in[112] ;
 wire \ring_501.inv_in[113] ;
 wire \ring_501.inv_in[114] ;
 wire \ring_501.inv_in[115] ;
 wire \ring_501.inv_in[116] ;
 wire \ring_501.inv_in[117] ;
 wire \ring_501.inv_in[118] ;
 wire \ring_501.inv_in[119] ;
 wire \ring_501.inv_in[11] ;
 wire \ring_501.inv_in[120] ;
 wire \ring_501.inv_in[121] ;
 wire \ring_501.inv_in[122] ;
 wire \ring_501.inv_in[123] ;
 wire \ring_501.inv_in[124] ;
 wire \ring_501.inv_in[125] ;
 wire \ring_501.inv_in[126] ;
 wire \ring_501.inv_in[127] ;
 wire \ring_501.inv_in[128] ;
 wire \ring_501.inv_in[129] ;
 wire \ring_501.inv_in[12] ;
 wire \ring_501.inv_in[130] ;
 wire \ring_501.inv_in[131] ;
 wire \ring_501.inv_in[132] ;
 wire \ring_501.inv_in[133] ;
 wire \ring_501.inv_in[134] ;
 wire \ring_501.inv_in[135] ;
 wire \ring_501.inv_in[136] ;
 wire \ring_501.inv_in[137] ;
 wire \ring_501.inv_in[138] ;
 wire \ring_501.inv_in[139] ;
 wire \ring_501.inv_in[13] ;
 wire \ring_501.inv_in[140] ;
 wire \ring_501.inv_in[141] ;
 wire \ring_501.inv_in[142] ;
 wire \ring_501.inv_in[143] ;
 wire \ring_501.inv_in[144] ;
 wire \ring_501.inv_in[145] ;
 wire \ring_501.inv_in[146] ;
 wire \ring_501.inv_in[147] ;
 wire \ring_501.inv_in[148] ;
 wire \ring_501.inv_in[149] ;
 wire \ring_501.inv_in[14] ;
 wire \ring_501.inv_in[150] ;
 wire \ring_501.inv_in[151] ;
 wire \ring_501.inv_in[152] ;
 wire \ring_501.inv_in[153] ;
 wire \ring_501.inv_in[154] ;
 wire \ring_501.inv_in[155] ;
 wire \ring_501.inv_in[156] ;
 wire \ring_501.inv_in[157] ;
 wire \ring_501.inv_in[158] ;
 wire \ring_501.inv_in[159] ;
 wire \ring_501.inv_in[15] ;
 wire \ring_501.inv_in[160] ;
 wire \ring_501.inv_in[161] ;
 wire \ring_501.inv_in[162] ;
 wire \ring_501.inv_in[163] ;
 wire \ring_501.inv_in[164] ;
 wire \ring_501.inv_in[165] ;
 wire \ring_501.inv_in[166] ;
 wire \ring_501.inv_in[167] ;
 wire \ring_501.inv_in[168] ;
 wire \ring_501.inv_in[169] ;
 wire \ring_501.inv_in[16] ;
 wire \ring_501.inv_in[170] ;
 wire \ring_501.inv_in[171] ;
 wire \ring_501.inv_in[172] ;
 wire \ring_501.inv_in[173] ;
 wire \ring_501.inv_in[174] ;
 wire \ring_501.inv_in[175] ;
 wire \ring_501.inv_in[176] ;
 wire \ring_501.inv_in[177] ;
 wire \ring_501.inv_in[178] ;
 wire \ring_501.inv_in[179] ;
 wire \ring_501.inv_in[17] ;
 wire \ring_501.inv_in[180] ;
 wire \ring_501.inv_in[181] ;
 wire \ring_501.inv_in[182] ;
 wire \ring_501.inv_in[183] ;
 wire \ring_501.inv_in[184] ;
 wire \ring_501.inv_in[185] ;
 wire \ring_501.inv_in[186] ;
 wire \ring_501.inv_in[187] ;
 wire \ring_501.inv_in[188] ;
 wire \ring_501.inv_in[189] ;
 wire \ring_501.inv_in[18] ;
 wire \ring_501.inv_in[190] ;
 wire \ring_501.inv_in[191] ;
 wire \ring_501.inv_in[192] ;
 wire \ring_501.inv_in[193] ;
 wire \ring_501.inv_in[194] ;
 wire \ring_501.inv_in[195] ;
 wire \ring_501.inv_in[196] ;
 wire \ring_501.inv_in[197] ;
 wire \ring_501.inv_in[198] ;
 wire \ring_501.inv_in[199] ;
 wire \ring_501.inv_in[19] ;
 wire \ring_501.inv_in[1] ;
 wire \ring_501.inv_in[200] ;
 wire \ring_501.inv_in[201] ;
 wire \ring_501.inv_in[202] ;
 wire \ring_501.inv_in[203] ;
 wire \ring_501.inv_in[204] ;
 wire \ring_501.inv_in[205] ;
 wire \ring_501.inv_in[206] ;
 wire \ring_501.inv_in[207] ;
 wire \ring_501.inv_in[208] ;
 wire \ring_501.inv_in[209] ;
 wire \ring_501.inv_in[20] ;
 wire \ring_501.inv_in[210] ;
 wire \ring_501.inv_in[211] ;
 wire \ring_501.inv_in[212] ;
 wire \ring_501.inv_in[213] ;
 wire \ring_501.inv_in[214] ;
 wire \ring_501.inv_in[215] ;
 wire \ring_501.inv_in[216] ;
 wire \ring_501.inv_in[217] ;
 wire \ring_501.inv_in[218] ;
 wire \ring_501.inv_in[219] ;
 wire \ring_501.inv_in[21] ;
 wire \ring_501.inv_in[220] ;
 wire \ring_501.inv_in[221] ;
 wire \ring_501.inv_in[222] ;
 wire \ring_501.inv_in[223] ;
 wire \ring_501.inv_in[224] ;
 wire \ring_501.inv_in[225] ;
 wire \ring_501.inv_in[226] ;
 wire \ring_501.inv_in[227] ;
 wire \ring_501.inv_in[228] ;
 wire \ring_501.inv_in[229] ;
 wire \ring_501.inv_in[22] ;
 wire \ring_501.inv_in[230] ;
 wire \ring_501.inv_in[231] ;
 wire \ring_501.inv_in[232] ;
 wire \ring_501.inv_in[233] ;
 wire \ring_501.inv_in[234] ;
 wire \ring_501.inv_in[235] ;
 wire \ring_501.inv_in[236] ;
 wire \ring_501.inv_in[237] ;
 wire \ring_501.inv_in[238] ;
 wire \ring_501.inv_in[239] ;
 wire \ring_501.inv_in[23] ;
 wire \ring_501.inv_in[240] ;
 wire \ring_501.inv_in[241] ;
 wire \ring_501.inv_in[242] ;
 wire \ring_501.inv_in[243] ;
 wire \ring_501.inv_in[244] ;
 wire \ring_501.inv_in[245] ;
 wire \ring_501.inv_in[246] ;
 wire \ring_501.inv_in[247] ;
 wire \ring_501.inv_in[248] ;
 wire \ring_501.inv_in[249] ;
 wire \ring_501.inv_in[24] ;
 wire \ring_501.inv_in[250] ;
 wire \ring_501.inv_in[251] ;
 wire \ring_501.inv_in[252] ;
 wire \ring_501.inv_in[253] ;
 wire \ring_501.inv_in[254] ;
 wire \ring_501.inv_in[255] ;
 wire \ring_501.inv_in[256] ;
 wire \ring_501.inv_in[257] ;
 wire \ring_501.inv_in[258] ;
 wire \ring_501.inv_in[259] ;
 wire \ring_501.inv_in[25] ;
 wire \ring_501.inv_in[260] ;
 wire \ring_501.inv_in[261] ;
 wire \ring_501.inv_in[262] ;
 wire \ring_501.inv_in[263] ;
 wire \ring_501.inv_in[264] ;
 wire \ring_501.inv_in[265] ;
 wire \ring_501.inv_in[266] ;
 wire \ring_501.inv_in[267] ;
 wire \ring_501.inv_in[268] ;
 wire \ring_501.inv_in[269] ;
 wire \ring_501.inv_in[26] ;
 wire \ring_501.inv_in[270] ;
 wire \ring_501.inv_in[271] ;
 wire \ring_501.inv_in[272] ;
 wire \ring_501.inv_in[273] ;
 wire \ring_501.inv_in[274] ;
 wire \ring_501.inv_in[275] ;
 wire \ring_501.inv_in[276] ;
 wire \ring_501.inv_in[277] ;
 wire \ring_501.inv_in[278] ;
 wire \ring_501.inv_in[279] ;
 wire \ring_501.inv_in[27] ;
 wire \ring_501.inv_in[280] ;
 wire \ring_501.inv_in[281] ;
 wire \ring_501.inv_in[282] ;
 wire \ring_501.inv_in[283] ;
 wire \ring_501.inv_in[284] ;
 wire \ring_501.inv_in[285] ;
 wire \ring_501.inv_in[286] ;
 wire \ring_501.inv_in[287] ;
 wire \ring_501.inv_in[288] ;
 wire \ring_501.inv_in[289] ;
 wire \ring_501.inv_in[28] ;
 wire \ring_501.inv_in[290] ;
 wire \ring_501.inv_in[291] ;
 wire \ring_501.inv_in[292] ;
 wire \ring_501.inv_in[293] ;
 wire \ring_501.inv_in[294] ;
 wire \ring_501.inv_in[295] ;
 wire \ring_501.inv_in[296] ;
 wire \ring_501.inv_in[297] ;
 wire \ring_501.inv_in[298] ;
 wire \ring_501.inv_in[299] ;
 wire \ring_501.inv_in[29] ;
 wire \ring_501.inv_in[2] ;
 wire \ring_501.inv_in[300] ;
 wire \ring_501.inv_in[301] ;
 wire \ring_501.inv_in[302] ;
 wire \ring_501.inv_in[303] ;
 wire \ring_501.inv_in[304] ;
 wire \ring_501.inv_in[305] ;
 wire \ring_501.inv_in[306] ;
 wire \ring_501.inv_in[307] ;
 wire \ring_501.inv_in[308] ;
 wire \ring_501.inv_in[309] ;
 wire \ring_501.inv_in[30] ;
 wire \ring_501.inv_in[310] ;
 wire \ring_501.inv_in[311] ;
 wire \ring_501.inv_in[312] ;
 wire \ring_501.inv_in[313] ;
 wire \ring_501.inv_in[314] ;
 wire \ring_501.inv_in[315] ;
 wire \ring_501.inv_in[316] ;
 wire \ring_501.inv_in[317] ;
 wire \ring_501.inv_in[318] ;
 wire \ring_501.inv_in[319] ;
 wire \ring_501.inv_in[31] ;
 wire \ring_501.inv_in[320] ;
 wire \ring_501.inv_in[321] ;
 wire \ring_501.inv_in[322] ;
 wire \ring_501.inv_in[323] ;
 wire \ring_501.inv_in[324] ;
 wire \ring_501.inv_in[325] ;
 wire \ring_501.inv_in[326] ;
 wire \ring_501.inv_in[327] ;
 wire \ring_501.inv_in[328] ;
 wire \ring_501.inv_in[329] ;
 wire \ring_501.inv_in[32] ;
 wire \ring_501.inv_in[330] ;
 wire \ring_501.inv_in[331] ;
 wire \ring_501.inv_in[332] ;
 wire \ring_501.inv_in[333] ;
 wire \ring_501.inv_in[334] ;
 wire \ring_501.inv_in[335] ;
 wire \ring_501.inv_in[336] ;
 wire \ring_501.inv_in[337] ;
 wire \ring_501.inv_in[338] ;
 wire \ring_501.inv_in[339] ;
 wire \ring_501.inv_in[33] ;
 wire \ring_501.inv_in[340] ;
 wire \ring_501.inv_in[341] ;
 wire \ring_501.inv_in[342] ;
 wire \ring_501.inv_in[343] ;
 wire \ring_501.inv_in[344] ;
 wire \ring_501.inv_in[345] ;
 wire \ring_501.inv_in[346] ;
 wire \ring_501.inv_in[347] ;
 wire \ring_501.inv_in[348] ;
 wire \ring_501.inv_in[349] ;
 wire \ring_501.inv_in[34] ;
 wire \ring_501.inv_in[350] ;
 wire \ring_501.inv_in[351] ;
 wire \ring_501.inv_in[352] ;
 wire \ring_501.inv_in[353] ;
 wire \ring_501.inv_in[354] ;
 wire \ring_501.inv_in[355] ;
 wire \ring_501.inv_in[356] ;
 wire \ring_501.inv_in[357] ;
 wire \ring_501.inv_in[358] ;
 wire \ring_501.inv_in[359] ;
 wire \ring_501.inv_in[35] ;
 wire \ring_501.inv_in[360] ;
 wire \ring_501.inv_in[361] ;
 wire \ring_501.inv_in[362] ;
 wire \ring_501.inv_in[363] ;
 wire \ring_501.inv_in[364] ;
 wire \ring_501.inv_in[365] ;
 wire \ring_501.inv_in[366] ;
 wire \ring_501.inv_in[367] ;
 wire \ring_501.inv_in[368] ;
 wire \ring_501.inv_in[369] ;
 wire \ring_501.inv_in[36] ;
 wire \ring_501.inv_in[370] ;
 wire \ring_501.inv_in[371] ;
 wire \ring_501.inv_in[372] ;
 wire \ring_501.inv_in[373] ;
 wire \ring_501.inv_in[374] ;
 wire \ring_501.inv_in[375] ;
 wire \ring_501.inv_in[376] ;
 wire \ring_501.inv_in[377] ;
 wire \ring_501.inv_in[378] ;
 wire \ring_501.inv_in[379] ;
 wire \ring_501.inv_in[37] ;
 wire \ring_501.inv_in[380] ;
 wire \ring_501.inv_in[381] ;
 wire \ring_501.inv_in[382] ;
 wire \ring_501.inv_in[383] ;
 wire \ring_501.inv_in[384] ;
 wire \ring_501.inv_in[385] ;
 wire \ring_501.inv_in[386] ;
 wire \ring_501.inv_in[387] ;
 wire \ring_501.inv_in[388] ;
 wire \ring_501.inv_in[389] ;
 wire \ring_501.inv_in[38] ;
 wire \ring_501.inv_in[390] ;
 wire \ring_501.inv_in[391] ;
 wire \ring_501.inv_in[392] ;
 wire \ring_501.inv_in[393] ;
 wire \ring_501.inv_in[394] ;
 wire \ring_501.inv_in[395] ;
 wire \ring_501.inv_in[396] ;
 wire \ring_501.inv_in[397] ;
 wire \ring_501.inv_in[398] ;
 wire \ring_501.inv_in[399] ;
 wire \ring_501.inv_in[39] ;
 wire \ring_501.inv_in[3] ;
 wire \ring_501.inv_in[400] ;
 wire \ring_501.inv_in[401] ;
 wire \ring_501.inv_in[402] ;
 wire \ring_501.inv_in[403] ;
 wire \ring_501.inv_in[404] ;
 wire \ring_501.inv_in[405] ;
 wire \ring_501.inv_in[406] ;
 wire \ring_501.inv_in[407] ;
 wire \ring_501.inv_in[408] ;
 wire \ring_501.inv_in[409] ;
 wire \ring_501.inv_in[40] ;
 wire \ring_501.inv_in[410] ;
 wire \ring_501.inv_in[411] ;
 wire \ring_501.inv_in[412] ;
 wire \ring_501.inv_in[413] ;
 wire \ring_501.inv_in[414] ;
 wire \ring_501.inv_in[415] ;
 wire \ring_501.inv_in[416] ;
 wire \ring_501.inv_in[417] ;
 wire \ring_501.inv_in[418] ;
 wire \ring_501.inv_in[419] ;
 wire \ring_501.inv_in[41] ;
 wire \ring_501.inv_in[420] ;
 wire \ring_501.inv_in[421] ;
 wire \ring_501.inv_in[422] ;
 wire \ring_501.inv_in[423] ;
 wire \ring_501.inv_in[424] ;
 wire \ring_501.inv_in[425] ;
 wire \ring_501.inv_in[426] ;
 wire \ring_501.inv_in[427] ;
 wire \ring_501.inv_in[428] ;
 wire \ring_501.inv_in[429] ;
 wire \ring_501.inv_in[42] ;
 wire \ring_501.inv_in[430] ;
 wire \ring_501.inv_in[431] ;
 wire \ring_501.inv_in[432] ;
 wire \ring_501.inv_in[433] ;
 wire \ring_501.inv_in[434] ;
 wire \ring_501.inv_in[435] ;
 wire \ring_501.inv_in[436] ;
 wire \ring_501.inv_in[437] ;
 wire \ring_501.inv_in[438] ;
 wire \ring_501.inv_in[439] ;
 wire \ring_501.inv_in[43] ;
 wire \ring_501.inv_in[440] ;
 wire \ring_501.inv_in[441] ;
 wire \ring_501.inv_in[442] ;
 wire \ring_501.inv_in[443] ;
 wire \ring_501.inv_in[444] ;
 wire \ring_501.inv_in[445] ;
 wire \ring_501.inv_in[446] ;
 wire \ring_501.inv_in[447] ;
 wire \ring_501.inv_in[448] ;
 wire \ring_501.inv_in[449] ;
 wire \ring_501.inv_in[44] ;
 wire \ring_501.inv_in[450] ;
 wire \ring_501.inv_in[451] ;
 wire \ring_501.inv_in[452] ;
 wire \ring_501.inv_in[453] ;
 wire \ring_501.inv_in[454] ;
 wire \ring_501.inv_in[455] ;
 wire \ring_501.inv_in[456] ;
 wire \ring_501.inv_in[457] ;
 wire \ring_501.inv_in[458] ;
 wire \ring_501.inv_in[459] ;
 wire \ring_501.inv_in[45] ;
 wire \ring_501.inv_in[460] ;
 wire \ring_501.inv_in[461] ;
 wire \ring_501.inv_in[462] ;
 wire \ring_501.inv_in[463] ;
 wire \ring_501.inv_in[464] ;
 wire \ring_501.inv_in[465] ;
 wire \ring_501.inv_in[466] ;
 wire \ring_501.inv_in[467] ;
 wire \ring_501.inv_in[468] ;
 wire \ring_501.inv_in[469] ;
 wire \ring_501.inv_in[46] ;
 wire \ring_501.inv_in[470] ;
 wire \ring_501.inv_in[471] ;
 wire \ring_501.inv_in[472] ;
 wire \ring_501.inv_in[473] ;
 wire \ring_501.inv_in[474] ;
 wire \ring_501.inv_in[475] ;
 wire \ring_501.inv_in[476] ;
 wire \ring_501.inv_in[477] ;
 wire \ring_501.inv_in[478] ;
 wire \ring_501.inv_in[479] ;
 wire \ring_501.inv_in[47] ;
 wire \ring_501.inv_in[480] ;
 wire \ring_501.inv_in[481] ;
 wire \ring_501.inv_in[482] ;
 wire \ring_501.inv_in[483] ;
 wire \ring_501.inv_in[484] ;
 wire \ring_501.inv_in[485] ;
 wire \ring_501.inv_in[486] ;
 wire \ring_501.inv_in[487] ;
 wire \ring_501.inv_in[488] ;
 wire \ring_501.inv_in[489] ;
 wire \ring_501.inv_in[48] ;
 wire \ring_501.inv_in[490] ;
 wire \ring_501.inv_in[491] ;
 wire \ring_501.inv_in[492] ;
 wire \ring_501.inv_in[493] ;
 wire \ring_501.inv_in[494] ;
 wire \ring_501.inv_in[495] ;
 wire \ring_501.inv_in[496] ;
 wire \ring_501.inv_in[497] ;
 wire \ring_501.inv_in[498] ;
 wire \ring_501.inv_in[499] ;
 wire \ring_501.inv_in[49] ;
 wire \ring_501.inv_in[4] ;
 wire \ring_501.inv_in[500] ;
 wire \ring_501.inv_in[50] ;
 wire \ring_501.inv_in[51] ;
 wire \ring_501.inv_in[52] ;
 wire \ring_501.inv_in[53] ;
 wire \ring_501.inv_in[54] ;
 wire \ring_501.inv_in[55] ;
 wire \ring_501.inv_in[56] ;
 wire \ring_501.inv_in[57] ;
 wire \ring_501.inv_in[58] ;
 wire \ring_501.inv_in[59] ;
 wire \ring_501.inv_in[5] ;
 wire \ring_501.inv_in[60] ;
 wire \ring_501.inv_in[61] ;
 wire \ring_501.inv_in[62] ;
 wire \ring_501.inv_in[63] ;
 wire \ring_501.inv_in[64] ;
 wire \ring_501.inv_in[65] ;
 wire \ring_501.inv_in[66] ;
 wire \ring_501.inv_in[67] ;
 wire \ring_501.inv_in[68] ;
 wire \ring_501.inv_in[69] ;
 wire \ring_501.inv_in[6] ;
 wire \ring_501.inv_in[70] ;
 wire \ring_501.inv_in[71] ;
 wire \ring_501.inv_in[72] ;
 wire \ring_501.inv_in[73] ;
 wire \ring_501.inv_in[74] ;
 wire \ring_501.inv_in[75] ;
 wire \ring_501.inv_in[76] ;
 wire \ring_501.inv_in[77] ;
 wire \ring_501.inv_in[78] ;
 wire \ring_501.inv_in[79] ;
 wire \ring_501.inv_in[7] ;
 wire \ring_501.inv_in[80] ;
 wire \ring_501.inv_in[81] ;
 wire \ring_501.inv_in[82] ;
 wire \ring_501.inv_in[83] ;
 wire \ring_501.inv_in[84] ;
 wire \ring_501.inv_in[85] ;
 wire \ring_501.inv_in[86] ;
 wire \ring_501.inv_in[87] ;
 wire \ring_501.inv_in[88] ;
 wire \ring_501.inv_in[89] ;
 wire \ring_501.inv_in[8] ;
 wire \ring_501.inv_in[90] ;
 wire \ring_501.inv_in[91] ;
 wire \ring_501.inv_in[92] ;
 wire \ring_501.inv_in[93] ;
 wire \ring_501.inv_in[94] ;
 wire \ring_501.inv_in[95] ;
 wire \ring_501.inv_in[96] ;
 wire \ring_501.inv_in[97] ;
 wire \ring_501.inv_in[98] ;
 wire \ring_501.inv_in[99] ;
 wire \ring_501.inv_in[9] ;
 wire \ring_501.inv_out[500] ;
 wire net43;
 wire net44;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net45;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;

 sg13g2_inv_1 _056_ (.Y(_011_),
    .A(\c2[4] ));
 sg13g2_and4_1 _057_ (.A(net6),
    .B(net5),
    .C(net8),
    .D(net7),
    .X(_012_));
 sg13g2_nand3_1 _058_ (.B(net3),
    .C(_012_),
    .A(net4),
    .Y(_013_));
 sg13g2_nand4_1 _059_ (.B(net17),
    .C(net2),
    .A(net18),
    .Y(_014_),
    .D(net1));
 sg13g2_nand4_1 _060_ (.B(net13),
    .C(net16),
    .A(net14),
    .Y(_015_),
    .D(net15));
 sg13g2_nand4_1 _061_ (.B(net9),
    .C(net12),
    .A(net10),
    .Y(_016_),
    .D(net11));
 sg13g2_nor4_1 _062_ (.A(_013_),
    .B(_014_),
    .C(_015_),
    .D(_016_),
    .Y(dummy));
 sg13g2_or3_2 _063_ (.A(net8),
    .B(net10),
    .C(net9),
    .X(uio_out[1]));
 sg13g2_nand2b_1 _064_ (.Y(_017_),
    .B(net4),
    .A_N(\c2[1] ));
 sg13g2_nor2b_1 _065_ (.A(net4),
    .B_N(\c2[1] ),
    .Y(_018_));
 sg13g2_nand2b_1 _066_ (.Y(_019_),
    .B(net3),
    .A_N(\c2[0] ));
 sg13g2_o21ai_1 _067_ (.B1(_017_),
    .Y(uio_out[6]),
    .A1(_018_),
    .A2(_019_));
 sg13g2_or2_2 _068_ (.X(uio_out[7]),
    .B(net5),
    .A(net6));
 sg13g2_and2_2 _069_ (.A(net1),
    .B(\ring_125.inv_out[124] ),
    .X(c1clock));
 sg13g2_and2_1 _070_ (.A(net1),
    .B(\ring_251.inv_out[250] ),
    .X(\ring_251.inv_in[0] ));
 sg13g2_and2_1 _071_ (.A(net1),
    .B(\ring_1001.inv_out[1000] ),
    .X(\ring_1001.inv_in[0] ));
 sg13g2_and2_2 _072_ (.A(net1),
    .B(\ring_25.inv_out[24] ),
    .X(fast_osc));
 sg13g2_and2_2 _073_ (.A(net1),
    .B(\ring_501.inv_out[500] ),
    .X(c0clock));
 sg13g2_xor2_1 _074_ (.B(\c0[1] ),
    .A(\c0[0] ),
    .X(_000_));
 sg13g2_nand3_1 _075_ (.B(\c0[1] ),
    .C(\c0[2] ),
    .A(\c0[0] ),
    .Y(_020_));
 sg13g2_a21o_1 _076_ (.A2(\c0[1] ),
    .A1(\c0[0] ),
    .B1(\c0[2] ),
    .X(_021_));
 sg13g2_and2_1 _077_ (.A(_020_),
    .B(_021_),
    .X(_001_));
 sg13g2_xnor2_1 _078_ (.Y(_002_),
    .A(\c0[3] ),
    .B(_020_));
 sg13g2_xor2_1 _079_ (.B(\c2[0] ),
    .A(\c2[1] ),
    .X(_006_));
 sg13g2_nand3_1 _080_ (.B(\c2[0] ),
    .C(\c2[2] ),
    .A(\c2[1] ),
    .Y(_022_));
 sg13g2_a21o_1 _081_ (.A2(\c2[0] ),
    .A1(\c2[1] ),
    .B1(\c2[2] ),
    .X(_023_));
 sg13g2_and2_1 _082_ (.A(_022_),
    .B(_023_),
    .X(_007_));
 sg13g2_nand4_1 _083_ (.B(\c2[0] ),
    .C(\c2[2] ),
    .A(\c2[1] ),
    .Y(_024_),
    .D(\c2[3] ));
 sg13g2_xnor2_1 _084_ (.Y(_008_),
    .A(\c2[3] ),
    .B(_022_));
 sg13g2_nor2_1 _085_ (.A(_011_),
    .B(_024_),
    .Y(_025_));
 sg13g2_xnor2_1 _086_ (.Y(_009_),
    .A(\c2[4] ),
    .B(_024_));
 sg13g2_xor2_1 _087_ (.B(_025_),
    .A(\c2[5] ),
    .X(_010_));
 sg13g2_xor2_1 _088_ (.B(\c1[1] ),
    .A(\c1[0] ),
    .X(_003_));
 sg13g2_nand3_1 _089_ (.B(\c1[1] ),
    .C(\c1[2] ),
    .A(\c1[0] ),
    .Y(_026_));
 sg13g2_a21o_1 _090_ (.A2(\c1[1] ),
    .A1(\c1[0] ),
    .B1(\c1[2] ),
    .X(_027_));
 sg13g2_and2_1 _091_ (.A(_026_),
    .B(_027_),
    .X(_004_));
 sg13g2_xnor2_1 _092_ (.Y(_005_),
    .A(\c1[3] ),
    .B(_026_));
 sg13g2_dfrbp_1 _093_ (.CLK(fast_osc),
    .RESET_B(net30),
    .D(_028_),
    .Q_N(_028_),
    .Q(\c2[0] ));
 sg13g2_dfrbp_1 _094_ (.CLK(fast_osc),
    .RESET_B(net31),
    .D(_006_),
    .Q_N(_032_),
    .Q(\c2[1] ));
 sg13g2_dfrbp_1 _095_ (.CLK(fast_osc),
    .RESET_B(net32),
    .D(_007_),
    .Q_N(_033_),
    .Q(\c2[2] ));
 sg13g2_dfrbp_1 _096_ (.CLK(fast_osc),
    .RESET_B(net33),
    .D(_008_),
    .Q_N(_034_),
    .Q(\c2[3] ));
 sg13g2_dfrbp_1 _097_ (.CLK(fast_osc),
    .RESET_B(net34),
    .D(_009_),
    .Q_N(_035_),
    .Q(\c2[4] ));
 sg13g2_dfrbp_1 _098_ (.CLK(fast_osc),
    .RESET_B(net35),
    .D(_010_),
    .Q_N(_036_),
    .Q(\c2[5] ));
 sg13g2_dfrbp_1 _099_ (.CLK(c1clock),
    .RESET_B(net36),
    .D(_030_),
    .Q_N(_030_),
    .Q(\c1[0] ));
 sg13g2_dfrbp_1 _100_ (.CLK(c1clock),
    .RESET_B(net37),
    .D(_003_),
    .Q_N(_037_),
    .Q(\c1[1] ));
 sg13g2_dfrbp_1 _101_ (.CLK(c1clock),
    .RESET_B(net38),
    .D(_004_),
    .Q_N(_038_),
    .Q(\c1[2] ));
 sg13g2_dfrbp_1 _102_ (.CLK(c1clock),
    .RESET_B(net39),
    .D(_005_),
    .Q_N(_039_),
    .Q(\c1[3] ));
 sg13g2_dfrbp_1 _103_ (.CLK(c0clock),
    .RESET_B(net40),
    .D(_029_),
    .Q_N(_029_),
    .Q(\c0[0] ));
 sg13g2_dfrbp_1 _104_ (.CLK(c0clock),
    .RESET_B(net41),
    .D(_000_),
    .Q_N(_040_),
    .Q(\c0[1] ));
 sg13g2_dfrbp_1 _105_ (.CLK(c0clock),
    .RESET_B(net28),
    .D(_001_),
    .Q_N(_041_),
    .Q(\c0[2] ));
 sg13g2_dfrbp_1 _106_ (.CLK(c0clock),
    .RESET_B(net29),
    .D(_002_),
    .Q_N(_031_),
    .Q(\c0[3] ));
 sg13g2_tiehi _106__29 (.L_HI(net29));
 sg13g2_tiehi _093__30 (.L_HI(net30));
 sg13g2_tiehi _094__31 (.L_HI(net31));
 sg13g2_tiehi _095__32 (.L_HI(net32));
 sg13g2_tiehi _096__33 (.L_HI(net33));
 sg13g2_tiehi _097__34 (.L_HI(net34));
 sg13g2_tiehi _098__35 (.L_HI(net35));
 sg13g2_tiehi _099__36 (.L_HI(net36));
 sg13g2_tiehi _100__37 (.L_HI(net37));
 sg13g2_tiehi _101__38 (.L_HI(net38));
 sg13g2_tiehi _102__39 (.L_HI(net39));
 sg13g2_tiehi _103__40 (.L_HI(net40));
 sg13g2_tiehi _104__41 (.L_HI(net41));
 sg13g2_tiehi tt_um_algofoogle_tt09_ring_osc2_42 (.L_HI(net42));
 sg13g2_tiehi tt_um_algofoogle_tt09_ring_osc2_43 (.L_HI(net43));
 sg13g2_tiehi tt_um_algofoogle_tt09_ring_osc2_44 (.L_HI(net44));
 sg13g2_tiehi tt_um_algofoogle_tt09_ring_osc2_45 (.L_HI(net45));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc2_20 (.L_LO(net20));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc2_21 (.L_LO(net21));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc2_22 (.L_LO(net22));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc2_23 (.L_LO(net23));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc2_24 (.L_LO(net24));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc2_25 (.L_LO(net25));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc2_26 (.L_LO(net26));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc2_27 (.L_LO(net27));
 sg13g2_tiehi _105__28 (.L_HI(net28));
 sg13g2_buf_1 _134_ (.A(dummy),
    .X(uio_out[0]));
 sg13g2_buf_1 _135_ (.A(c1clock),
    .X(uo_out[0]));
 sg13g2_buf_1 _136_ (.A(\ring_251.inv_in[0] ),
    .X(uo_out[1]));
 sg13g2_buf_1 _137_ (.A(c0clock),
    .X(uo_out[2]));
 sg13g2_buf_1 _138_ (.A(\ring_1001.inv_in[0] ),
    .X(uo_out[3]));
 sg13g2_buf_1 _139_ (.A(\c0[3] ),
    .X(uo_out[4]));
 sg13g2_buf_1 _140_ (.A(\c1[3] ),
    .X(uo_out[5]));
 sg13g2_buf_1 _141_ (.A(\c2[5] ),
    .X(uo_out[6]));
 sg13g2_inv_1 \ring_1001.inv_array[0]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[1] ),
    .A(\ring_1001.inv_in[0] ));
 sg13g2_inv_1 \ring_1001.inv_array[1000]/sky_inverter/_0_  (.Y(\ring_1001.inv_out[1000] ),
    .A(\ring_1001.inv_in[1000] ));
 sg13g2_inv_1 \ring_1001.inv_array[100]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[101] ),
    .A(\ring_1001.inv_in[100] ));
 sg13g2_inv_1 \ring_1001.inv_array[101]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[102] ),
    .A(\ring_1001.inv_in[101] ));
 sg13g2_inv_1 \ring_1001.inv_array[102]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[103] ),
    .A(\ring_1001.inv_in[102] ));
 sg13g2_inv_1 \ring_1001.inv_array[103]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[104] ),
    .A(\ring_1001.inv_in[103] ));
 sg13g2_inv_1 \ring_1001.inv_array[104]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[105] ),
    .A(\ring_1001.inv_in[104] ));
 sg13g2_inv_1 \ring_1001.inv_array[105]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[106] ),
    .A(\ring_1001.inv_in[105] ));
 sg13g2_inv_1 \ring_1001.inv_array[106]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[107] ),
    .A(\ring_1001.inv_in[106] ));
 sg13g2_inv_1 \ring_1001.inv_array[107]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[108] ),
    .A(\ring_1001.inv_in[107] ));
 sg13g2_inv_1 \ring_1001.inv_array[108]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[109] ),
    .A(\ring_1001.inv_in[108] ));
 sg13g2_inv_1 \ring_1001.inv_array[109]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[110] ),
    .A(\ring_1001.inv_in[109] ));
 sg13g2_inv_1 \ring_1001.inv_array[10]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[11] ),
    .A(\ring_1001.inv_in[10] ));
 sg13g2_inv_1 \ring_1001.inv_array[110]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[111] ),
    .A(\ring_1001.inv_in[110] ));
 sg13g2_inv_1 \ring_1001.inv_array[111]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[112] ),
    .A(\ring_1001.inv_in[111] ));
 sg13g2_inv_1 \ring_1001.inv_array[112]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[113] ),
    .A(\ring_1001.inv_in[112] ));
 sg13g2_inv_1 \ring_1001.inv_array[113]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[114] ),
    .A(\ring_1001.inv_in[113] ));
 sg13g2_inv_1 \ring_1001.inv_array[114]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[115] ),
    .A(\ring_1001.inv_in[114] ));
 sg13g2_inv_1 \ring_1001.inv_array[115]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[116] ),
    .A(\ring_1001.inv_in[115] ));
 sg13g2_inv_1 \ring_1001.inv_array[116]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[117] ),
    .A(\ring_1001.inv_in[116] ));
 sg13g2_inv_1 \ring_1001.inv_array[117]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[118] ),
    .A(\ring_1001.inv_in[117] ));
 sg13g2_inv_1 \ring_1001.inv_array[118]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[119] ),
    .A(\ring_1001.inv_in[118] ));
 sg13g2_inv_1 \ring_1001.inv_array[119]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[120] ),
    .A(\ring_1001.inv_in[119] ));
 sg13g2_inv_1 \ring_1001.inv_array[11]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[12] ),
    .A(\ring_1001.inv_in[11] ));
 sg13g2_inv_1 \ring_1001.inv_array[120]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[121] ),
    .A(\ring_1001.inv_in[120] ));
 sg13g2_inv_1 \ring_1001.inv_array[121]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[122] ),
    .A(\ring_1001.inv_in[121] ));
 sg13g2_inv_1 \ring_1001.inv_array[122]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[123] ),
    .A(\ring_1001.inv_in[122] ));
 sg13g2_inv_1 \ring_1001.inv_array[123]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[124] ),
    .A(\ring_1001.inv_in[123] ));
 sg13g2_inv_1 \ring_1001.inv_array[124]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[125] ),
    .A(\ring_1001.inv_in[124] ));
 sg13g2_inv_1 \ring_1001.inv_array[125]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[126] ),
    .A(\ring_1001.inv_in[125] ));
 sg13g2_inv_1 \ring_1001.inv_array[126]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[127] ),
    .A(\ring_1001.inv_in[126] ));
 sg13g2_inv_1 \ring_1001.inv_array[127]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[128] ),
    .A(\ring_1001.inv_in[127] ));
 sg13g2_inv_1 \ring_1001.inv_array[128]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[129] ),
    .A(\ring_1001.inv_in[128] ));
 sg13g2_inv_1 \ring_1001.inv_array[129]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[130] ),
    .A(\ring_1001.inv_in[129] ));
 sg13g2_inv_1 \ring_1001.inv_array[12]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[13] ),
    .A(\ring_1001.inv_in[12] ));
 sg13g2_inv_1 \ring_1001.inv_array[130]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[131] ),
    .A(\ring_1001.inv_in[130] ));
 sg13g2_inv_1 \ring_1001.inv_array[131]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[132] ),
    .A(\ring_1001.inv_in[131] ));
 sg13g2_inv_1 \ring_1001.inv_array[132]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[133] ),
    .A(\ring_1001.inv_in[132] ));
 sg13g2_inv_1 \ring_1001.inv_array[133]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[134] ),
    .A(\ring_1001.inv_in[133] ));
 sg13g2_inv_1 \ring_1001.inv_array[134]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[135] ),
    .A(\ring_1001.inv_in[134] ));
 sg13g2_inv_1 \ring_1001.inv_array[135]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[136] ),
    .A(\ring_1001.inv_in[135] ));
 sg13g2_inv_1 \ring_1001.inv_array[136]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[137] ),
    .A(\ring_1001.inv_in[136] ));
 sg13g2_inv_1 \ring_1001.inv_array[137]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[138] ),
    .A(\ring_1001.inv_in[137] ));
 sg13g2_inv_1 \ring_1001.inv_array[138]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[139] ),
    .A(\ring_1001.inv_in[138] ));
 sg13g2_inv_1 \ring_1001.inv_array[139]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[140] ),
    .A(\ring_1001.inv_in[139] ));
 sg13g2_inv_1 \ring_1001.inv_array[13]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[14] ),
    .A(\ring_1001.inv_in[13] ));
 sg13g2_inv_1 \ring_1001.inv_array[140]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[141] ),
    .A(\ring_1001.inv_in[140] ));
 sg13g2_inv_1 \ring_1001.inv_array[141]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[142] ),
    .A(\ring_1001.inv_in[141] ));
 sg13g2_inv_1 \ring_1001.inv_array[142]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[143] ),
    .A(\ring_1001.inv_in[142] ));
 sg13g2_inv_1 \ring_1001.inv_array[143]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[144] ),
    .A(\ring_1001.inv_in[143] ));
 sg13g2_inv_1 \ring_1001.inv_array[144]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[145] ),
    .A(\ring_1001.inv_in[144] ));
 sg13g2_inv_1 \ring_1001.inv_array[145]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[146] ),
    .A(\ring_1001.inv_in[145] ));
 sg13g2_inv_1 \ring_1001.inv_array[146]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[147] ),
    .A(\ring_1001.inv_in[146] ));
 sg13g2_inv_1 \ring_1001.inv_array[147]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[148] ),
    .A(\ring_1001.inv_in[147] ));
 sg13g2_inv_1 \ring_1001.inv_array[148]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[149] ),
    .A(\ring_1001.inv_in[148] ));
 sg13g2_inv_1 \ring_1001.inv_array[149]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[150] ),
    .A(\ring_1001.inv_in[149] ));
 sg13g2_inv_1 \ring_1001.inv_array[14]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[15] ),
    .A(\ring_1001.inv_in[14] ));
 sg13g2_inv_1 \ring_1001.inv_array[150]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[151] ),
    .A(\ring_1001.inv_in[150] ));
 sg13g2_inv_1 \ring_1001.inv_array[151]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[152] ),
    .A(\ring_1001.inv_in[151] ));
 sg13g2_inv_1 \ring_1001.inv_array[152]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[153] ),
    .A(\ring_1001.inv_in[152] ));
 sg13g2_inv_1 \ring_1001.inv_array[153]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[154] ),
    .A(\ring_1001.inv_in[153] ));
 sg13g2_inv_1 \ring_1001.inv_array[154]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[155] ),
    .A(\ring_1001.inv_in[154] ));
 sg13g2_inv_1 \ring_1001.inv_array[155]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[156] ),
    .A(\ring_1001.inv_in[155] ));
 sg13g2_inv_1 \ring_1001.inv_array[156]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[157] ),
    .A(\ring_1001.inv_in[156] ));
 sg13g2_inv_1 \ring_1001.inv_array[157]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[158] ),
    .A(\ring_1001.inv_in[157] ));
 sg13g2_inv_1 \ring_1001.inv_array[158]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[159] ),
    .A(\ring_1001.inv_in[158] ));
 sg13g2_inv_1 \ring_1001.inv_array[159]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[160] ),
    .A(\ring_1001.inv_in[159] ));
 sg13g2_inv_1 \ring_1001.inv_array[15]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[16] ),
    .A(\ring_1001.inv_in[15] ));
 sg13g2_inv_1 \ring_1001.inv_array[160]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[161] ),
    .A(\ring_1001.inv_in[160] ));
 sg13g2_inv_1 \ring_1001.inv_array[161]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[162] ),
    .A(\ring_1001.inv_in[161] ));
 sg13g2_inv_1 \ring_1001.inv_array[162]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[163] ),
    .A(\ring_1001.inv_in[162] ));
 sg13g2_inv_1 \ring_1001.inv_array[163]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[164] ),
    .A(\ring_1001.inv_in[163] ));
 sg13g2_inv_1 \ring_1001.inv_array[164]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[165] ),
    .A(\ring_1001.inv_in[164] ));
 sg13g2_inv_1 \ring_1001.inv_array[165]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[166] ),
    .A(\ring_1001.inv_in[165] ));
 sg13g2_inv_1 \ring_1001.inv_array[166]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[167] ),
    .A(\ring_1001.inv_in[166] ));
 sg13g2_inv_1 \ring_1001.inv_array[167]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[168] ),
    .A(\ring_1001.inv_in[167] ));
 sg13g2_inv_1 \ring_1001.inv_array[168]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[169] ),
    .A(\ring_1001.inv_in[168] ));
 sg13g2_inv_1 \ring_1001.inv_array[169]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[170] ),
    .A(\ring_1001.inv_in[169] ));
 sg13g2_inv_1 \ring_1001.inv_array[16]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[17] ),
    .A(\ring_1001.inv_in[16] ));
 sg13g2_inv_1 \ring_1001.inv_array[170]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[171] ),
    .A(\ring_1001.inv_in[170] ));
 sg13g2_inv_1 \ring_1001.inv_array[171]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[172] ),
    .A(\ring_1001.inv_in[171] ));
 sg13g2_inv_1 \ring_1001.inv_array[172]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[173] ),
    .A(\ring_1001.inv_in[172] ));
 sg13g2_inv_1 \ring_1001.inv_array[173]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[174] ),
    .A(\ring_1001.inv_in[173] ));
 sg13g2_inv_1 \ring_1001.inv_array[174]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[175] ),
    .A(\ring_1001.inv_in[174] ));
 sg13g2_inv_1 \ring_1001.inv_array[175]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[176] ),
    .A(\ring_1001.inv_in[175] ));
 sg13g2_inv_1 \ring_1001.inv_array[176]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[177] ),
    .A(\ring_1001.inv_in[176] ));
 sg13g2_inv_1 \ring_1001.inv_array[177]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[178] ),
    .A(\ring_1001.inv_in[177] ));
 sg13g2_inv_1 \ring_1001.inv_array[178]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[179] ),
    .A(\ring_1001.inv_in[178] ));
 sg13g2_inv_1 \ring_1001.inv_array[179]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[180] ),
    .A(\ring_1001.inv_in[179] ));
 sg13g2_inv_1 \ring_1001.inv_array[17]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[18] ),
    .A(\ring_1001.inv_in[17] ));
 sg13g2_inv_1 \ring_1001.inv_array[180]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[181] ),
    .A(\ring_1001.inv_in[180] ));
 sg13g2_inv_1 \ring_1001.inv_array[181]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[182] ),
    .A(\ring_1001.inv_in[181] ));
 sg13g2_inv_1 \ring_1001.inv_array[182]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[183] ),
    .A(\ring_1001.inv_in[182] ));
 sg13g2_inv_1 \ring_1001.inv_array[183]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[184] ),
    .A(\ring_1001.inv_in[183] ));
 sg13g2_inv_1 \ring_1001.inv_array[184]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[185] ),
    .A(\ring_1001.inv_in[184] ));
 sg13g2_inv_1 \ring_1001.inv_array[185]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[186] ),
    .A(\ring_1001.inv_in[185] ));
 sg13g2_inv_1 \ring_1001.inv_array[186]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[187] ),
    .A(\ring_1001.inv_in[186] ));
 sg13g2_inv_1 \ring_1001.inv_array[187]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[188] ),
    .A(\ring_1001.inv_in[187] ));
 sg13g2_inv_1 \ring_1001.inv_array[188]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[189] ),
    .A(\ring_1001.inv_in[188] ));
 sg13g2_inv_1 \ring_1001.inv_array[189]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[190] ),
    .A(\ring_1001.inv_in[189] ));
 sg13g2_inv_1 \ring_1001.inv_array[18]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[19] ),
    .A(\ring_1001.inv_in[18] ));
 sg13g2_inv_1 \ring_1001.inv_array[190]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[191] ),
    .A(\ring_1001.inv_in[190] ));
 sg13g2_inv_1 \ring_1001.inv_array[191]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[192] ),
    .A(\ring_1001.inv_in[191] ));
 sg13g2_inv_1 \ring_1001.inv_array[192]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[193] ),
    .A(\ring_1001.inv_in[192] ));
 sg13g2_inv_1 \ring_1001.inv_array[193]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[194] ),
    .A(\ring_1001.inv_in[193] ));
 sg13g2_inv_1 \ring_1001.inv_array[194]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[195] ),
    .A(\ring_1001.inv_in[194] ));
 sg13g2_inv_1 \ring_1001.inv_array[195]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[196] ),
    .A(\ring_1001.inv_in[195] ));
 sg13g2_inv_1 \ring_1001.inv_array[196]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[197] ),
    .A(\ring_1001.inv_in[196] ));
 sg13g2_inv_1 \ring_1001.inv_array[197]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[198] ),
    .A(\ring_1001.inv_in[197] ));
 sg13g2_inv_1 \ring_1001.inv_array[198]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[199] ),
    .A(\ring_1001.inv_in[198] ));
 sg13g2_inv_1 \ring_1001.inv_array[199]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[200] ),
    .A(\ring_1001.inv_in[199] ));
 sg13g2_inv_1 \ring_1001.inv_array[19]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[20] ),
    .A(\ring_1001.inv_in[19] ));
 sg13g2_inv_1 \ring_1001.inv_array[1]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[2] ),
    .A(\ring_1001.inv_in[1] ));
 sg13g2_inv_1 \ring_1001.inv_array[200]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[201] ),
    .A(\ring_1001.inv_in[200] ));
 sg13g2_inv_1 \ring_1001.inv_array[201]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[202] ),
    .A(\ring_1001.inv_in[201] ));
 sg13g2_inv_1 \ring_1001.inv_array[202]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[203] ),
    .A(\ring_1001.inv_in[202] ));
 sg13g2_inv_1 \ring_1001.inv_array[203]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[204] ),
    .A(\ring_1001.inv_in[203] ));
 sg13g2_inv_1 \ring_1001.inv_array[204]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[205] ),
    .A(\ring_1001.inv_in[204] ));
 sg13g2_inv_1 \ring_1001.inv_array[205]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[206] ),
    .A(\ring_1001.inv_in[205] ));
 sg13g2_inv_1 \ring_1001.inv_array[206]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[207] ),
    .A(\ring_1001.inv_in[206] ));
 sg13g2_inv_1 \ring_1001.inv_array[207]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[208] ),
    .A(\ring_1001.inv_in[207] ));
 sg13g2_inv_1 \ring_1001.inv_array[208]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[209] ),
    .A(\ring_1001.inv_in[208] ));
 sg13g2_inv_1 \ring_1001.inv_array[209]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[210] ),
    .A(\ring_1001.inv_in[209] ));
 sg13g2_inv_1 \ring_1001.inv_array[20]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[21] ),
    .A(\ring_1001.inv_in[20] ));
 sg13g2_inv_1 \ring_1001.inv_array[210]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[211] ),
    .A(\ring_1001.inv_in[210] ));
 sg13g2_inv_1 \ring_1001.inv_array[211]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[212] ),
    .A(\ring_1001.inv_in[211] ));
 sg13g2_inv_1 \ring_1001.inv_array[212]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[213] ),
    .A(\ring_1001.inv_in[212] ));
 sg13g2_inv_1 \ring_1001.inv_array[213]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[214] ),
    .A(\ring_1001.inv_in[213] ));
 sg13g2_inv_1 \ring_1001.inv_array[214]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[215] ),
    .A(\ring_1001.inv_in[214] ));
 sg13g2_inv_1 \ring_1001.inv_array[215]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[216] ),
    .A(\ring_1001.inv_in[215] ));
 sg13g2_inv_1 \ring_1001.inv_array[216]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[217] ),
    .A(\ring_1001.inv_in[216] ));
 sg13g2_inv_1 \ring_1001.inv_array[217]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[218] ),
    .A(\ring_1001.inv_in[217] ));
 sg13g2_inv_1 \ring_1001.inv_array[218]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[219] ),
    .A(\ring_1001.inv_in[218] ));
 sg13g2_inv_1 \ring_1001.inv_array[219]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[220] ),
    .A(\ring_1001.inv_in[219] ));
 sg13g2_inv_1 \ring_1001.inv_array[21]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[22] ),
    .A(\ring_1001.inv_in[21] ));
 sg13g2_inv_1 \ring_1001.inv_array[220]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[221] ),
    .A(\ring_1001.inv_in[220] ));
 sg13g2_inv_1 \ring_1001.inv_array[221]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[222] ),
    .A(\ring_1001.inv_in[221] ));
 sg13g2_inv_1 \ring_1001.inv_array[222]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[223] ),
    .A(\ring_1001.inv_in[222] ));
 sg13g2_inv_1 \ring_1001.inv_array[223]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[224] ),
    .A(\ring_1001.inv_in[223] ));
 sg13g2_inv_1 \ring_1001.inv_array[224]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[225] ),
    .A(\ring_1001.inv_in[224] ));
 sg13g2_inv_1 \ring_1001.inv_array[225]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[226] ),
    .A(\ring_1001.inv_in[225] ));
 sg13g2_inv_1 \ring_1001.inv_array[226]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[227] ),
    .A(\ring_1001.inv_in[226] ));
 sg13g2_inv_1 \ring_1001.inv_array[227]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[228] ),
    .A(\ring_1001.inv_in[227] ));
 sg13g2_inv_1 \ring_1001.inv_array[228]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[229] ),
    .A(\ring_1001.inv_in[228] ));
 sg13g2_inv_1 \ring_1001.inv_array[229]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[230] ),
    .A(\ring_1001.inv_in[229] ));
 sg13g2_inv_1 \ring_1001.inv_array[22]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[23] ),
    .A(\ring_1001.inv_in[22] ));
 sg13g2_inv_1 \ring_1001.inv_array[230]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[231] ),
    .A(\ring_1001.inv_in[230] ));
 sg13g2_inv_1 \ring_1001.inv_array[231]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[232] ),
    .A(\ring_1001.inv_in[231] ));
 sg13g2_inv_1 \ring_1001.inv_array[232]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[233] ),
    .A(\ring_1001.inv_in[232] ));
 sg13g2_inv_1 \ring_1001.inv_array[233]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[234] ),
    .A(\ring_1001.inv_in[233] ));
 sg13g2_inv_1 \ring_1001.inv_array[234]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[235] ),
    .A(\ring_1001.inv_in[234] ));
 sg13g2_inv_1 \ring_1001.inv_array[235]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[236] ),
    .A(\ring_1001.inv_in[235] ));
 sg13g2_inv_1 \ring_1001.inv_array[236]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[237] ),
    .A(\ring_1001.inv_in[236] ));
 sg13g2_inv_1 \ring_1001.inv_array[237]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[238] ),
    .A(\ring_1001.inv_in[237] ));
 sg13g2_inv_1 \ring_1001.inv_array[238]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[239] ),
    .A(\ring_1001.inv_in[238] ));
 sg13g2_inv_1 \ring_1001.inv_array[239]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[240] ),
    .A(\ring_1001.inv_in[239] ));
 sg13g2_inv_1 \ring_1001.inv_array[23]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[24] ),
    .A(\ring_1001.inv_in[23] ));
 sg13g2_inv_1 \ring_1001.inv_array[240]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[241] ),
    .A(\ring_1001.inv_in[240] ));
 sg13g2_inv_1 \ring_1001.inv_array[241]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[242] ),
    .A(\ring_1001.inv_in[241] ));
 sg13g2_inv_1 \ring_1001.inv_array[242]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[243] ),
    .A(\ring_1001.inv_in[242] ));
 sg13g2_inv_1 \ring_1001.inv_array[243]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[244] ),
    .A(\ring_1001.inv_in[243] ));
 sg13g2_inv_1 \ring_1001.inv_array[244]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[245] ),
    .A(\ring_1001.inv_in[244] ));
 sg13g2_inv_1 \ring_1001.inv_array[245]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[246] ),
    .A(\ring_1001.inv_in[245] ));
 sg13g2_inv_1 \ring_1001.inv_array[246]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[247] ),
    .A(\ring_1001.inv_in[246] ));
 sg13g2_inv_1 \ring_1001.inv_array[247]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[248] ),
    .A(\ring_1001.inv_in[247] ));
 sg13g2_inv_1 \ring_1001.inv_array[248]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[249] ),
    .A(\ring_1001.inv_in[248] ));
 sg13g2_inv_1 \ring_1001.inv_array[249]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[250] ),
    .A(\ring_1001.inv_in[249] ));
 sg13g2_inv_1 \ring_1001.inv_array[24]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[25] ),
    .A(\ring_1001.inv_in[24] ));
 sg13g2_inv_1 \ring_1001.inv_array[250]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[251] ),
    .A(\ring_1001.inv_in[250] ));
 sg13g2_inv_1 \ring_1001.inv_array[251]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[252] ),
    .A(\ring_1001.inv_in[251] ));
 sg13g2_inv_1 \ring_1001.inv_array[252]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[253] ),
    .A(\ring_1001.inv_in[252] ));
 sg13g2_inv_1 \ring_1001.inv_array[253]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[254] ),
    .A(\ring_1001.inv_in[253] ));
 sg13g2_inv_1 \ring_1001.inv_array[254]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[255] ),
    .A(\ring_1001.inv_in[254] ));
 sg13g2_inv_1 \ring_1001.inv_array[255]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[256] ),
    .A(\ring_1001.inv_in[255] ));
 sg13g2_inv_1 \ring_1001.inv_array[256]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[257] ),
    .A(\ring_1001.inv_in[256] ));
 sg13g2_inv_1 \ring_1001.inv_array[257]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[258] ),
    .A(\ring_1001.inv_in[257] ));
 sg13g2_inv_1 \ring_1001.inv_array[258]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[259] ),
    .A(\ring_1001.inv_in[258] ));
 sg13g2_inv_1 \ring_1001.inv_array[259]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[260] ),
    .A(\ring_1001.inv_in[259] ));
 sg13g2_inv_1 \ring_1001.inv_array[25]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[26] ),
    .A(\ring_1001.inv_in[25] ));
 sg13g2_inv_1 \ring_1001.inv_array[260]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[261] ),
    .A(\ring_1001.inv_in[260] ));
 sg13g2_inv_1 \ring_1001.inv_array[261]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[262] ),
    .A(\ring_1001.inv_in[261] ));
 sg13g2_inv_1 \ring_1001.inv_array[262]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[263] ),
    .A(\ring_1001.inv_in[262] ));
 sg13g2_inv_1 \ring_1001.inv_array[263]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[264] ),
    .A(\ring_1001.inv_in[263] ));
 sg13g2_inv_1 \ring_1001.inv_array[264]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[265] ),
    .A(\ring_1001.inv_in[264] ));
 sg13g2_inv_1 \ring_1001.inv_array[265]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[266] ),
    .A(\ring_1001.inv_in[265] ));
 sg13g2_inv_1 \ring_1001.inv_array[266]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[267] ),
    .A(\ring_1001.inv_in[266] ));
 sg13g2_inv_1 \ring_1001.inv_array[267]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[268] ),
    .A(\ring_1001.inv_in[267] ));
 sg13g2_inv_1 \ring_1001.inv_array[268]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[269] ),
    .A(\ring_1001.inv_in[268] ));
 sg13g2_inv_1 \ring_1001.inv_array[269]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[270] ),
    .A(\ring_1001.inv_in[269] ));
 sg13g2_inv_1 \ring_1001.inv_array[26]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[27] ),
    .A(\ring_1001.inv_in[26] ));
 sg13g2_inv_1 \ring_1001.inv_array[270]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[271] ),
    .A(\ring_1001.inv_in[270] ));
 sg13g2_inv_1 \ring_1001.inv_array[271]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[272] ),
    .A(\ring_1001.inv_in[271] ));
 sg13g2_inv_1 \ring_1001.inv_array[272]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[273] ),
    .A(\ring_1001.inv_in[272] ));
 sg13g2_inv_1 \ring_1001.inv_array[273]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[274] ),
    .A(\ring_1001.inv_in[273] ));
 sg13g2_inv_1 \ring_1001.inv_array[274]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[275] ),
    .A(\ring_1001.inv_in[274] ));
 sg13g2_inv_1 \ring_1001.inv_array[275]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[276] ),
    .A(\ring_1001.inv_in[275] ));
 sg13g2_inv_1 \ring_1001.inv_array[276]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[277] ),
    .A(\ring_1001.inv_in[276] ));
 sg13g2_inv_1 \ring_1001.inv_array[277]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[278] ),
    .A(\ring_1001.inv_in[277] ));
 sg13g2_inv_1 \ring_1001.inv_array[278]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[279] ),
    .A(\ring_1001.inv_in[278] ));
 sg13g2_inv_1 \ring_1001.inv_array[279]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[280] ),
    .A(\ring_1001.inv_in[279] ));
 sg13g2_inv_1 \ring_1001.inv_array[27]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[28] ),
    .A(\ring_1001.inv_in[27] ));
 sg13g2_inv_1 \ring_1001.inv_array[280]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[281] ),
    .A(\ring_1001.inv_in[280] ));
 sg13g2_inv_1 \ring_1001.inv_array[281]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[282] ),
    .A(\ring_1001.inv_in[281] ));
 sg13g2_inv_1 \ring_1001.inv_array[282]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[283] ),
    .A(\ring_1001.inv_in[282] ));
 sg13g2_inv_1 \ring_1001.inv_array[283]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[284] ),
    .A(\ring_1001.inv_in[283] ));
 sg13g2_inv_1 \ring_1001.inv_array[284]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[285] ),
    .A(\ring_1001.inv_in[284] ));
 sg13g2_inv_1 \ring_1001.inv_array[285]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[286] ),
    .A(\ring_1001.inv_in[285] ));
 sg13g2_inv_1 \ring_1001.inv_array[286]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[287] ),
    .A(\ring_1001.inv_in[286] ));
 sg13g2_inv_1 \ring_1001.inv_array[287]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[288] ),
    .A(\ring_1001.inv_in[287] ));
 sg13g2_inv_1 \ring_1001.inv_array[288]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[289] ),
    .A(\ring_1001.inv_in[288] ));
 sg13g2_inv_1 \ring_1001.inv_array[289]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[290] ),
    .A(\ring_1001.inv_in[289] ));
 sg13g2_inv_1 \ring_1001.inv_array[28]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[29] ),
    .A(\ring_1001.inv_in[28] ));
 sg13g2_inv_1 \ring_1001.inv_array[290]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[291] ),
    .A(\ring_1001.inv_in[290] ));
 sg13g2_inv_1 \ring_1001.inv_array[291]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[292] ),
    .A(\ring_1001.inv_in[291] ));
 sg13g2_inv_1 \ring_1001.inv_array[292]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[293] ),
    .A(\ring_1001.inv_in[292] ));
 sg13g2_inv_1 \ring_1001.inv_array[293]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[294] ),
    .A(\ring_1001.inv_in[293] ));
 sg13g2_inv_1 \ring_1001.inv_array[294]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[295] ),
    .A(\ring_1001.inv_in[294] ));
 sg13g2_inv_1 \ring_1001.inv_array[295]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[296] ),
    .A(\ring_1001.inv_in[295] ));
 sg13g2_inv_1 \ring_1001.inv_array[296]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[297] ),
    .A(\ring_1001.inv_in[296] ));
 sg13g2_inv_1 \ring_1001.inv_array[297]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[298] ),
    .A(\ring_1001.inv_in[297] ));
 sg13g2_inv_1 \ring_1001.inv_array[298]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[299] ),
    .A(\ring_1001.inv_in[298] ));
 sg13g2_inv_1 \ring_1001.inv_array[299]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[300] ),
    .A(\ring_1001.inv_in[299] ));
 sg13g2_inv_1 \ring_1001.inv_array[29]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[30] ),
    .A(\ring_1001.inv_in[29] ));
 sg13g2_inv_1 \ring_1001.inv_array[2]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[3] ),
    .A(\ring_1001.inv_in[2] ));
 sg13g2_inv_1 \ring_1001.inv_array[300]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[301] ),
    .A(\ring_1001.inv_in[300] ));
 sg13g2_inv_1 \ring_1001.inv_array[301]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[302] ),
    .A(\ring_1001.inv_in[301] ));
 sg13g2_inv_1 \ring_1001.inv_array[302]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[303] ),
    .A(\ring_1001.inv_in[302] ));
 sg13g2_inv_1 \ring_1001.inv_array[303]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[304] ),
    .A(\ring_1001.inv_in[303] ));
 sg13g2_inv_1 \ring_1001.inv_array[304]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[305] ),
    .A(\ring_1001.inv_in[304] ));
 sg13g2_inv_1 \ring_1001.inv_array[305]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[306] ),
    .A(\ring_1001.inv_in[305] ));
 sg13g2_inv_1 \ring_1001.inv_array[306]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[307] ),
    .A(\ring_1001.inv_in[306] ));
 sg13g2_inv_1 \ring_1001.inv_array[307]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[308] ),
    .A(\ring_1001.inv_in[307] ));
 sg13g2_inv_1 \ring_1001.inv_array[308]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[309] ),
    .A(\ring_1001.inv_in[308] ));
 sg13g2_inv_1 \ring_1001.inv_array[309]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[310] ),
    .A(\ring_1001.inv_in[309] ));
 sg13g2_inv_1 \ring_1001.inv_array[30]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[31] ),
    .A(\ring_1001.inv_in[30] ));
 sg13g2_inv_1 \ring_1001.inv_array[310]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[311] ),
    .A(\ring_1001.inv_in[310] ));
 sg13g2_inv_1 \ring_1001.inv_array[311]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[312] ),
    .A(\ring_1001.inv_in[311] ));
 sg13g2_inv_1 \ring_1001.inv_array[312]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[313] ),
    .A(\ring_1001.inv_in[312] ));
 sg13g2_inv_1 \ring_1001.inv_array[313]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[314] ),
    .A(\ring_1001.inv_in[313] ));
 sg13g2_inv_1 \ring_1001.inv_array[314]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[315] ),
    .A(\ring_1001.inv_in[314] ));
 sg13g2_inv_1 \ring_1001.inv_array[315]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[316] ),
    .A(\ring_1001.inv_in[315] ));
 sg13g2_inv_1 \ring_1001.inv_array[316]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[317] ),
    .A(\ring_1001.inv_in[316] ));
 sg13g2_inv_1 \ring_1001.inv_array[317]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[318] ),
    .A(\ring_1001.inv_in[317] ));
 sg13g2_inv_1 \ring_1001.inv_array[318]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[319] ),
    .A(\ring_1001.inv_in[318] ));
 sg13g2_inv_1 \ring_1001.inv_array[319]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[320] ),
    .A(\ring_1001.inv_in[319] ));
 sg13g2_inv_1 \ring_1001.inv_array[31]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[32] ),
    .A(\ring_1001.inv_in[31] ));
 sg13g2_inv_1 \ring_1001.inv_array[320]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[321] ),
    .A(\ring_1001.inv_in[320] ));
 sg13g2_inv_1 \ring_1001.inv_array[321]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[322] ),
    .A(\ring_1001.inv_in[321] ));
 sg13g2_inv_1 \ring_1001.inv_array[322]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[323] ),
    .A(\ring_1001.inv_in[322] ));
 sg13g2_inv_1 \ring_1001.inv_array[323]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[324] ),
    .A(\ring_1001.inv_in[323] ));
 sg13g2_inv_1 \ring_1001.inv_array[324]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[325] ),
    .A(\ring_1001.inv_in[324] ));
 sg13g2_inv_1 \ring_1001.inv_array[325]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[326] ),
    .A(\ring_1001.inv_in[325] ));
 sg13g2_inv_1 \ring_1001.inv_array[326]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[327] ),
    .A(\ring_1001.inv_in[326] ));
 sg13g2_inv_1 \ring_1001.inv_array[327]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[328] ),
    .A(\ring_1001.inv_in[327] ));
 sg13g2_inv_1 \ring_1001.inv_array[328]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[329] ),
    .A(\ring_1001.inv_in[328] ));
 sg13g2_inv_1 \ring_1001.inv_array[329]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[330] ),
    .A(\ring_1001.inv_in[329] ));
 sg13g2_inv_1 \ring_1001.inv_array[32]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[33] ),
    .A(\ring_1001.inv_in[32] ));
 sg13g2_inv_1 \ring_1001.inv_array[330]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[331] ),
    .A(\ring_1001.inv_in[330] ));
 sg13g2_inv_1 \ring_1001.inv_array[331]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[332] ),
    .A(\ring_1001.inv_in[331] ));
 sg13g2_inv_1 \ring_1001.inv_array[332]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[333] ),
    .A(\ring_1001.inv_in[332] ));
 sg13g2_inv_1 \ring_1001.inv_array[333]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[334] ),
    .A(\ring_1001.inv_in[333] ));
 sg13g2_inv_1 \ring_1001.inv_array[334]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[335] ),
    .A(\ring_1001.inv_in[334] ));
 sg13g2_inv_1 \ring_1001.inv_array[335]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[336] ),
    .A(\ring_1001.inv_in[335] ));
 sg13g2_inv_1 \ring_1001.inv_array[336]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[337] ),
    .A(\ring_1001.inv_in[336] ));
 sg13g2_inv_1 \ring_1001.inv_array[337]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[338] ),
    .A(\ring_1001.inv_in[337] ));
 sg13g2_inv_1 \ring_1001.inv_array[338]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[339] ),
    .A(\ring_1001.inv_in[338] ));
 sg13g2_inv_1 \ring_1001.inv_array[339]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[340] ),
    .A(\ring_1001.inv_in[339] ));
 sg13g2_inv_1 \ring_1001.inv_array[33]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[34] ),
    .A(\ring_1001.inv_in[33] ));
 sg13g2_inv_1 \ring_1001.inv_array[340]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[341] ),
    .A(\ring_1001.inv_in[340] ));
 sg13g2_inv_1 \ring_1001.inv_array[341]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[342] ),
    .A(\ring_1001.inv_in[341] ));
 sg13g2_inv_1 \ring_1001.inv_array[342]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[343] ),
    .A(\ring_1001.inv_in[342] ));
 sg13g2_inv_1 \ring_1001.inv_array[343]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[344] ),
    .A(\ring_1001.inv_in[343] ));
 sg13g2_inv_1 \ring_1001.inv_array[344]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[345] ),
    .A(\ring_1001.inv_in[344] ));
 sg13g2_inv_1 \ring_1001.inv_array[345]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[346] ),
    .A(\ring_1001.inv_in[345] ));
 sg13g2_inv_1 \ring_1001.inv_array[346]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[347] ),
    .A(\ring_1001.inv_in[346] ));
 sg13g2_inv_1 \ring_1001.inv_array[347]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[348] ),
    .A(\ring_1001.inv_in[347] ));
 sg13g2_inv_1 \ring_1001.inv_array[348]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[349] ),
    .A(\ring_1001.inv_in[348] ));
 sg13g2_inv_1 \ring_1001.inv_array[349]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[350] ),
    .A(\ring_1001.inv_in[349] ));
 sg13g2_inv_1 \ring_1001.inv_array[34]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[35] ),
    .A(\ring_1001.inv_in[34] ));
 sg13g2_inv_1 \ring_1001.inv_array[350]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[351] ),
    .A(\ring_1001.inv_in[350] ));
 sg13g2_inv_1 \ring_1001.inv_array[351]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[352] ),
    .A(\ring_1001.inv_in[351] ));
 sg13g2_inv_1 \ring_1001.inv_array[352]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[353] ),
    .A(\ring_1001.inv_in[352] ));
 sg13g2_inv_1 \ring_1001.inv_array[353]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[354] ),
    .A(\ring_1001.inv_in[353] ));
 sg13g2_inv_1 \ring_1001.inv_array[354]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[355] ),
    .A(\ring_1001.inv_in[354] ));
 sg13g2_inv_1 \ring_1001.inv_array[355]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[356] ),
    .A(\ring_1001.inv_in[355] ));
 sg13g2_inv_1 \ring_1001.inv_array[356]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[357] ),
    .A(\ring_1001.inv_in[356] ));
 sg13g2_inv_1 \ring_1001.inv_array[357]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[358] ),
    .A(\ring_1001.inv_in[357] ));
 sg13g2_inv_1 \ring_1001.inv_array[358]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[359] ),
    .A(\ring_1001.inv_in[358] ));
 sg13g2_inv_1 \ring_1001.inv_array[359]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[360] ),
    .A(\ring_1001.inv_in[359] ));
 sg13g2_inv_1 \ring_1001.inv_array[35]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[36] ),
    .A(\ring_1001.inv_in[35] ));
 sg13g2_inv_1 \ring_1001.inv_array[360]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[361] ),
    .A(\ring_1001.inv_in[360] ));
 sg13g2_inv_1 \ring_1001.inv_array[361]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[362] ),
    .A(\ring_1001.inv_in[361] ));
 sg13g2_inv_1 \ring_1001.inv_array[362]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[363] ),
    .A(\ring_1001.inv_in[362] ));
 sg13g2_inv_1 \ring_1001.inv_array[363]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[364] ),
    .A(\ring_1001.inv_in[363] ));
 sg13g2_inv_1 \ring_1001.inv_array[364]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[365] ),
    .A(\ring_1001.inv_in[364] ));
 sg13g2_inv_1 \ring_1001.inv_array[365]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[366] ),
    .A(\ring_1001.inv_in[365] ));
 sg13g2_inv_1 \ring_1001.inv_array[366]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[367] ),
    .A(\ring_1001.inv_in[366] ));
 sg13g2_inv_1 \ring_1001.inv_array[367]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[368] ),
    .A(\ring_1001.inv_in[367] ));
 sg13g2_inv_1 \ring_1001.inv_array[368]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[369] ),
    .A(\ring_1001.inv_in[368] ));
 sg13g2_inv_1 \ring_1001.inv_array[369]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[370] ),
    .A(\ring_1001.inv_in[369] ));
 sg13g2_inv_1 \ring_1001.inv_array[36]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[37] ),
    .A(\ring_1001.inv_in[36] ));
 sg13g2_inv_1 \ring_1001.inv_array[370]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[371] ),
    .A(\ring_1001.inv_in[370] ));
 sg13g2_inv_1 \ring_1001.inv_array[371]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[372] ),
    .A(\ring_1001.inv_in[371] ));
 sg13g2_inv_1 \ring_1001.inv_array[372]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[373] ),
    .A(\ring_1001.inv_in[372] ));
 sg13g2_inv_1 \ring_1001.inv_array[373]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[374] ),
    .A(\ring_1001.inv_in[373] ));
 sg13g2_inv_1 \ring_1001.inv_array[374]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[375] ),
    .A(\ring_1001.inv_in[374] ));
 sg13g2_inv_1 \ring_1001.inv_array[375]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[376] ),
    .A(\ring_1001.inv_in[375] ));
 sg13g2_inv_1 \ring_1001.inv_array[376]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[377] ),
    .A(\ring_1001.inv_in[376] ));
 sg13g2_inv_1 \ring_1001.inv_array[377]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[378] ),
    .A(\ring_1001.inv_in[377] ));
 sg13g2_inv_1 \ring_1001.inv_array[378]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[379] ),
    .A(\ring_1001.inv_in[378] ));
 sg13g2_inv_1 \ring_1001.inv_array[379]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[380] ),
    .A(\ring_1001.inv_in[379] ));
 sg13g2_inv_1 \ring_1001.inv_array[37]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[38] ),
    .A(\ring_1001.inv_in[37] ));
 sg13g2_inv_1 \ring_1001.inv_array[380]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[381] ),
    .A(\ring_1001.inv_in[380] ));
 sg13g2_inv_1 \ring_1001.inv_array[381]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[382] ),
    .A(\ring_1001.inv_in[381] ));
 sg13g2_inv_1 \ring_1001.inv_array[382]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[383] ),
    .A(\ring_1001.inv_in[382] ));
 sg13g2_inv_1 \ring_1001.inv_array[383]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[384] ),
    .A(\ring_1001.inv_in[383] ));
 sg13g2_inv_1 \ring_1001.inv_array[384]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[385] ),
    .A(\ring_1001.inv_in[384] ));
 sg13g2_inv_1 \ring_1001.inv_array[385]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[386] ),
    .A(\ring_1001.inv_in[385] ));
 sg13g2_inv_1 \ring_1001.inv_array[386]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[387] ),
    .A(\ring_1001.inv_in[386] ));
 sg13g2_inv_1 \ring_1001.inv_array[387]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[388] ),
    .A(\ring_1001.inv_in[387] ));
 sg13g2_inv_1 \ring_1001.inv_array[388]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[389] ),
    .A(\ring_1001.inv_in[388] ));
 sg13g2_inv_1 \ring_1001.inv_array[389]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[390] ),
    .A(\ring_1001.inv_in[389] ));
 sg13g2_inv_1 \ring_1001.inv_array[38]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[39] ),
    .A(\ring_1001.inv_in[38] ));
 sg13g2_inv_1 \ring_1001.inv_array[390]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[391] ),
    .A(\ring_1001.inv_in[390] ));
 sg13g2_inv_1 \ring_1001.inv_array[391]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[392] ),
    .A(\ring_1001.inv_in[391] ));
 sg13g2_inv_1 \ring_1001.inv_array[392]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[393] ),
    .A(\ring_1001.inv_in[392] ));
 sg13g2_inv_1 \ring_1001.inv_array[393]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[394] ),
    .A(\ring_1001.inv_in[393] ));
 sg13g2_inv_1 \ring_1001.inv_array[394]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[395] ),
    .A(\ring_1001.inv_in[394] ));
 sg13g2_inv_1 \ring_1001.inv_array[395]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[396] ),
    .A(\ring_1001.inv_in[395] ));
 sg13g2_inv_1 \ring_1001.inv_array[396]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[397] ),
    .A(\ring_1001.inv_in[396] ));
 sg13g2_inv_1 \ring_1001.inv_array[397]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[398] ),
    .A(\ring_1001.inv_in[397] ));
 sg13g2_inv_1 \ring_1001.inv_array[398]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[399] ),
    .A(\ring_1001.inv_in[398] ));
 sg13g2_inv_1 \ring_1001.inv_array[399]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[400] ),
    .A(\ring_1001.inv_in[399] ));
 sg13g2_inv_1 \ring_1001.inv_array[39]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[40] ),
    .A(\ring_1001.inv_in[39] ));
 sg13g2_inv_1 \ring_1001.inv_array[3]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[4] ),
    .A(\ring_1001.inv_in[3] ));
 sg13g2_inv_1 \ring_1001.inv_array[400]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[401] ),
    .A(\ring_1001.inv_in[400] ));
 sg13g2_inv_1 \ring_1001.inv_array[401]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[402] ),
    .A(\ring_1001.inv_in[401] ));
 sg13g2_inv_1 \ring_1001.inv_array[402]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[403] ),
    .A(\ring_1001.inv_in[402] ));
 sg13g2_inv_1 \ring_1001.inv_array[403]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[404] ),
    .A(\ring_1001.inv_in[403] ));
 sg13g2_inv_1 \ring_1001.inv_array[404]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[405] ),
    .A(\ring_1001.inv_in[404] ));
 sg13g2_inv_1 \ring_1001.inv_array[405]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[406] ),
    .A(\ring_1001.inv_in[405] ));
 sg13g2_inv_1 \ring_1001.inv_array[406]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[407] ),
    .A(\ring_1001.inv_in[406] ));
 sg13g2_inv_1 \ring_1001.inv_array[407]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[408] ),
    .A(\ring_1001.inv_in[407] ));
 sg13g2_inv_1 \ring_1001.inv_array[408]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[409] ),
    .A(\ring_1001.inv_in[408] ));
 sg13g2_inv_1 \ring_1001.inv_array[409]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[410] ),
    .A(\ring_1001.inv_in[409] ));
 sg13g2_inv_1 \ring_1001.inv_array[40]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[41] ),
    .A(\ring_1001.inv_in[40] ));
 sg13g2_inv_1 \ring_1001.inv_array[410]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[411] ),
    .A(\ring_1001.inv_in[410] ));
 sg13g2_inv_1 \ring_1001.inv_array[411]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[412] ),
    .A(\ring_1001.inv_in[411] ));
 sg13g2_inv_1 \ring_1001.inv_array[412]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[413] ),
    .A(\ring_1001.inv_in[412] ));
 sg13g2_inv_1 \ring_1001.inv_array[413]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[414] ),
    .A(\ring_1001.inv_in[413] ));
 sg13g2_inv_1 \ring_1001.inv_array[414]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[415] ),
    .A(\ring_1001.inv_in[414] ));
 sg13g2_inv_1 \ring_1001.inv_array[415]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[416] ),
    .A(\ring_1001.inv_in[415] ));
 sg13g2_inv_1 \ring_1001.inv_array[416]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[417] ),
    .A(\ring_1001.inv_in[416] ));
 sg13g2_inv_1 \ring_1001.inv_array[417]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[418] ),
    .A(\ring_1001.inv_in[417] ));
 sg13g2_inv_1 \ring_1001.inv_array[418]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[419] ),
    .A(\ring_1001.inv_in[418] ));
 sg13g2_inv_1 \ring_1001.inv_array[419]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[420] ),
    .A(\ring_1001.inv_in[419] ));
 sg13g2_inv_1 \ring_1001.inv_array[41]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[42] ),
    .A(\ring_1001.inv_in[41] ));
 sg13g2_inv_1 \ring_1001.inv_array[420]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[421] ),
    .A(\ring_1001.inv_in[420] ));
 sg13g2_inv_1 \ring_1001.inv_array[421]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[422] ),
    .A(\ring_1001.inv_in[421] ));
 sg13g2_inv_1 \ring_1001.inv_array[422]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[423] ),
    .A(\ring_1001.inv_in[422] ));
 sg13g2_inv_1 \ring_1001.inv_array[423]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[424] ),
    .A(\ring_1001.inv_in[423] ));
 sg13g2_inv_1 \ring_1001.inv_array[424]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[425] ),
    .A(\ring_1001.inv_in[424] ));
 sg13g2_inv_1 \ring_1001.inv_array[425]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[426] ),
    .A(\ring_1001.inv_in[425] ));
 sg13g2_inv_1 \ring_1001.inv_array[426]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[427] ),
    .A(\ring_1001.inv_in[426] ));
 sg13g2_inv_1 \ring_1001.inv_array[427]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[428] ),
    .A(\ring_1001.inv_in[427] ));
 sg13g2_inv_1 \ring_1001.inv_array[428]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[429] ),
    .A(\ring_1001.inv_in[428] ));
 sg13g2_inv_1 \ring_1001.inv_array[429]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[430] ),
    .A(\ring_1001.inv_in[429] ));
 sg13g2_inv_1 \ring_1001.inv_array[42]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[43] ),
    .A(\ring_1001.inv_in[42] ));
 sg13g2_inv_1 \ring_1001.inv_array[430]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[431] ),
    .A(\ring_1001.inv_in[430] ));
 sg13g2_inv_1 \ring_1001.inv_array[431]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[432] ),
    .A(\ring_1001.inv_in[431] ));
 sg13g2_inv_1 \ring_1001.inv_array[432]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[433] ),
    .A(\ring_1001.inv_in[432] ));
 sg13g2_inv_1 \ring_1001.inv_array[433]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[434] ),
    .A(\ring_1001.inv_in[433] ));
 sg13g2_inv_1 \ring_1001.inv_array[434]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[435] ),
    .A(\ring_1001.inv_in[434] ));
 sg13g2_inv_1 \ring_1001.inv_array[435]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[436] ),
    .A(\ring_1001.inv_in[435] ));
 sg13g2_inv_1 \ring_1001.inv_array[436]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[437] ),
    .A(\ring_1001.inv_in[436] ));
 sg13g2_inv_1 \ring_1001.inv_array[437]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[438] ),
    .A(\ring_1001.inv_in[437] ));
 sg13g2_inv_1 \ring_1001.inv_array[438]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[439] ),
    .A(\ring_1001.inv_in[438] ));
 sg13g2_inv_1 \ring_1001.inv_array[439]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[440] ),
    .A(\ring_1001.inv_in[439] ));
 sg13g2_inv_1 \ring_1001.inv_array[43]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[44] ),
    .A(\ring_1001.inv_in[43] ));
 sg13g2_inv_1 \ring_1001.inv_array[440]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[441] ),
    .A(\ring_1001.inv_in[440] ));
 sg13g2_inv_1 \ring_1001.inv_array[441]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[442] ),
    .A(\ring_1001.inv_in[441] ));
 sg13g2_inv_1 \ring_1001.inv_array[442]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[443] ),
    .A(\ring_1001.inv_in[442] ));
 sg13g2_inv_1 \ring_1001.inv_array[443]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[444] ),
    .A(\ring_1001.inv_in[443] ));
 sg13g2_inv_1 \ring_1001.inv_array[444]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[445] ),
    .A(\ring_1001.inv_in[444] ));
 sg13g2_inv_1 \ring_1001.inv_array[445]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[446] ),
    .A(\ring_1001.inv_in[445] ));
 sg13g2_inv_1 \ring_1001.inv_array[446]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[447] ),
    .A(\ring_1001.inv_in[446] ));
 sg13g2_inv_1 \ring_1001.inv_array[447]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[448] ),
    .A(\ring_1001.inv_in[447] ));
 sg13g2_inv_1 \ring_1001.inv_array[448]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[449] ),
    .A(\ring_1001.inv_in[448] ));
 sg13g2_inv_1 \ring_1001.inv_array[449]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[450] ),
    .A(\ring_1001.inv_in[449] ));
 sg13g2_inv_1 \ring_1001.inv_array[44]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[45] ),
    .A(\ring_1001.inv_in[44] ));
 sg13g2_inv_1 \ring_1001.inv_array[450]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[451] ),
    .A(\ring_1001.inv_in[450] ));
 sg13g2_inv_1 \ring_1001.inv_array[451]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[452] ),
    .A(\ring_1001.inv_in[451] ));
 sg13g2_inv_1 \ring_1001.inv_array[452]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[453] ),
    .A(\ring_1001.inv_in[452] ));
 sg13g2_inv_1 \ring_1001.inv_array[453]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[454] ),
    .A(\ring_1001.inv_in[453] ));
 sg13g2_inv_1 \ring_1001.inv_array[454]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[455] ),
    .A(\ring_1001.inv_in[454] ));
 sg13g2_inv_1 \ring_1001.inv_array[455]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[456] ),
    .A(\ring_1001.inv_in[455] ));
 sg13g2_inv_1 \ring_1001.inv_array[456]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[457] ),
    .A(\ring_1001.inv_in[456] ));
 sg13g2_inv_1 \ring_1001.inv_array[457]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[458] ),
    .A(\ring_1001.inv_in[457] ));
 sg13g2_inv_1 \ring_1001.inv_array[458]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[459] ),
    .A(\ring_1001.inv_in[458] ));
 sg13g2_inv_1 \ring_1001.inv_array[459]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[460] ),
    .A(\ring_1001.inv_in[459] ));
 sg13g2_inv_1 \ring_1001.inv_array[45]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[46] ),
    .A(\ring_1001.inv_in[45] ));
 sg13g2_inv_1 \ring_1001.inv_array[460]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[461] ),
    .A(\ring_1001.inv_in[460] ));
 sg13g2_inv_1 \ring_1001.inv_array[461]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[462] ),
    .A(\ring_1001.inv_in[461] ));
 sg13g2_inv_1 \ring_1001.inv_array[462]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[463] ),
    .A(\ring_1001.inv_in[462] ));
 sg13g2_inv_1 \ring_1001.inv_array[463]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[464] ),
    .A(\ring_1001.inv_in[463] ));
 sg13g2_inv_1 \ring_1001.inv_array[464]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[465] ),
    .A(\ring_1001.inv_in[464] ));
 sg13g2_inv_1 \ring_1001.inv_array[465]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[466] ),
    .A(\ring_1001.inv_in[465] ));
 sg13g2_inv_1 \ring_1001.inv_array[466]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[467] ),
    .A(\ring_1001.inv_in[466] ));
 sg13g2_inv_1 \ring_1001.inv_array[467]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[468] ),
    .A(\ring_1001.inv_in[467] ));
 sg13g2_inv_1 \ring_1001.inv_array[468]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[469] ),
    .A(\ring_1001.inv_in[468] ));
 sg13g2_inv_1 \ring_1001.inv_array[469]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[470] ),
    .A(\ring_1001.inv_in[469] ));
 sg13g2_inv_1 \ring_1001.inv_array[46]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[47] ),
    .A(\ring_1001.inv_in[46] ));
 sg13g2_inv_1 \ring_1001.inv_array[470]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[471] ),
    .A(\ring_1001.inv_in[470] ));
 sg13g2_inv_1 \ring_1001.inv_array[471]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[472] ),
    .A(\ring_1001.inv_in[471] ));
 sg13g2_inv_1 \ring_1001.inv_array[472]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[473] ),
    .A(\ring_1001.inv_in[472] ));
 sg13g2_inv_1 \ring_1001.inv_array[473]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[474] ),
    .A(\ring_1001.inv_in[473] ));
 sg13g2_inv_1 \ring_1001.inv_array[474]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[475] ),
    .A(\ring_1001.inv_in[474] ));
 sg13g2_inv_1 \ring_1001.inv_array[475]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[476] ),
    .A(\ring_1001.inv_in[475] ));
 sg13g2_inv_1 \ring_1001.inv_array[476]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[477] ),
    .A(\ring_1001.inv_in[476] ));
 sg13g2_inv_1 \ring_1001.inv_array[477]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[478] ),
    .A(\ring_1001.inv_in[477] ));
 sg13g2_inv_1 \ring_1001.inv_array[478]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[479] ),
    .A(\ring_1001.inv_in[478] ));
 sg13g2_inv_1 \ring_1001.inv_array[479]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[480] ),
    .A(\ring_1001.inv_in[479] ));
 sg13g2_inv_1 \ring_1001.inv_array[47]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[48] ),
    .A(\ring_1001.inv_in[47] ));
 sg13g2_inv_1 \ring_1001.inv_array[480]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[481] ),
    .A(\ring_1001.inv_in[480] ));
 sg13g2_inv_1 \ring_1001.inv_array[481]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[482] ),
    .A(\ring_1001.inv_in[481] ));
 sg13g2_inv_1 \ring_1001.inv_array[482]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[483] ),
    .A(\ring_1001.inv_in[482] ));
 sg13g2_inv_1 \ring_1001.inv_array[483]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[484] ),
    .A(\ring_1001.inv_in[483] ));
 sg13g2_inv_1 \ring_1001.inv_array[484]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[485] ),
    .A(\ring_1001.inv_in[484] ));
 sg13g2_inv_1 \ring_1001.inv_array[485]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[486] ),
    .A(\ring_1001.inv_in[485] ));
 sg13g2_inv_1 \ring_1001.inv_array[486]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[487] ),
    .A(\ring_1001.inv_in[486] ));
 sg13g2_inv_1 \ring_1001.inv_array[487]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[488] ),
    .A(\ring_1001.inv_in[487] ));
 sg13g2_inv_1 \ring_1001.inv_array[488]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[489] ),
    .A(\ring_1001.inv_in[488] ));
 sg13g2_inv_1 \ring_1001.inv_array[489]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[490] ),
    .A(\ring_1001.inv_in[489] ));
 sg13g2_inv_1 \ring_1001.inv_array[48]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[49] ),
    .A(\ring_1001.inv_in[48] ));
 sg13g2_inv_1 \ring_1001.inv_array[490]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[491] ),
    .A(\ring_1001.inv_in[490] ));
 sg13g2_inv_1 \ring_1001.inv_array[491]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[492] ),
    .A(\ring_1001.inv_in[491] ));
 sg13g2_inv_1 \ring_1001.inv_array[492]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[493] ),
    .A(\ring_1001.inv_in[492] ));
 sg13g2_inv_1 \ring_1001.inv_array[493]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[494] ),
    .A(\ring_1001.inv_in[493] ));
 sg13g2_inv_1 \ring_1001.inv_array[494]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[495] ),
    .A(\ring_1001.inv_in[494] ));
 sg13g2_inv_1 \ring_1001.inv_array[495]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[496] ),
    .A(\ring_1001.inv_in[495] ));
 sg13g2_inv_1 \ring_1001.inv_array[496]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[497] ),
    .A(\ring_1001.inv_in[496] ));
 sg13g2_inv_1 \ring_1001.inv_array[497]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[498] ),
    .A(\ring_1001.inv_in[497] ));
 sg13g2_inv_1 \ring_1001.inv_array[498]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[499] ),
    .A(\ring_1001.inv_in[498] ));
 sg13g2_inv_1 \ring_1001.inv_array[499]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[500] ),
    .A(\ring_1001.inv_in[499] ));
 sg13g2_inv_1 \ring_1001.inv_array[49]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[50] ),
    .A(\ring_1001.inv_in[49] ));
 sg13g2_inv_1 \ring_1001.inv_array[4]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[5] ),
    .A(\ring_1001.inv_in[4] ));
 sg13g2_inv_1 \ring_1001.inv_array[500]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[501] ),
    .A(\ring_1001.inv_in[500] ));
 sg13g2_inv_1 \ring_1001.inv_array[501]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[502] ),
    .A(\ring_1001.inv_in[501] ));
 sg13g2_inv_1 \ring_1001.inv_array[502]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[503] ),
    .A(\ring_1001.inv_in[502] ));
 sg13g2_inv_1 \ring_1001.inv_array[503]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[504] ),
    .A(\ring_1001.inv_in[503] ));
 sg13g2_inv_1 \ring_1001.inv_array[504]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[505] ),
    .A(\ring_1001.inv_in[504] ));
 sg13g2_inv_1 \ring_1001.inv_array[505]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[506] ),
    .A(\ring_1001.inv_in[505] ));
 sg13g2_inv_1 \ring_1001.inv_array[506]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[507] ),
    .A(\ring_1001.inv_in[506] ));
 sg13g2_inv_1 \ring_1001.inv_array[507]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[508] ),
    .A(\ring_1001.inv_in[507] ));
 sg13g2_inv_1 \ring_1001.inv_array[508]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[509] ),
    .A(\ring_1001.inv_in[508] ));
 sg13g2_inv_1 \ring_1001.inv_array[509]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[510] ),
    .A(\ring_1001.inv_in[509] ));
 sg13g2_inv_1 \ring_1001.inv_array[50]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[51] ),
    .A(\ring_1001.inv_in[50] ));
 sg13g2_inv_1 \ring_1001.inv_array[510]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[511] ),
    .A(\ring_1001.inv_in[510] ));
 sg13g2_inv_1 \ring_1001.inv_array[511]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[512] ),
    .A(\ring_1001.inv_in[511] ));
 sg13g2_inv_1 \ring_1001.inv_array[512]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[513] ),
    .A(\ring_1001.inv_in[512] ));
 sg13g2_inv_1 \ring_1001.inv_array[513]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[514] ),
    .A(\ring_1001.inv_in[513] ));
 sg13g2_inv_1 \ring_1001.inv_array[514]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[515] ),
    .A(\ring_1001.inv_in[514] ));
 sg13g2_inv_1 \ring_1001.inv_array[515]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[516] ),
    .A(\ring_1001.inv_in[515] ));
 sg13g2_inv_1 \ring_1001.inv_array[516]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[517] ),
    .A(\ring_1001.inv_in[516] ));
 sg13g2_inv_1 \ring_1001.inv_array[517]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[518] ),
    .A(\ring_1001.inv_in[517] ));
 sg13g2_inv_1 \ring_1001.inv_array[518]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[519] ),
    .A(\ring_1001.inv_in[518] ));
 sg13g2_inv_1 \ring_1001.inv_array[519]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[520] ),
    .A(\ring_1001.inv_in[519] ));
 sg13g2_inv_1 \ring_1001.inv_array[51]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[52] ),
    .A(\ring_1001.inv_in[51] ));
 sg13g2_inv_1 \ring_1001.inv_array[520]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[521] ),
    .A(\ring_1001.inv_in[520] ));
 sg13g2_inv_1 \ring_1001.inv_array[521]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[522] ),
    .A(\ring_1001.inv_in[521] ));
 sg13g2_inv_1 \ring_1001.inv_array[522]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[523] ),
    .A(\ring_1001.inv_in[522] ));
 sg13g2_inv_1 \ring_1001.inv_array[523]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[524] ),
    .A(\ring_1001.inv_in[523] ));
 sg13g2_inv_1 \ring_1001.inv_array[524]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[525] ),
    .A(\ring_1001.inv_in[524] ));
 sg13g2_inv_1 \ring_1001.inv_array[525]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[526] ),
    .A(\ring_1001.inv_in[525] ));
 sg13g2_inv_1 \ring_1001.inv_array[526]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[527] ),
    .A(\ring_1001.inv_in[526] ));
 sg13g2_inv_1 \ring_1001.inv_array[527]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[528] ),
    .A(\ring_1001.inv_in[527] ));
 sg13g2_inv_1 \ring_1001.inv_array[528]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[529] ),
    .A(\ring_1001.inv_in[528] ));
 sg13g2_inv_1 \ring_1001.inv_array[529]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[530] ),
    .A(\ring_1001.inv_in[529] ));
 sg13g2_inv_1 \ring_1001.inv_array[52]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[53] ),
    .A(\ring_1001.inv_in[52] ));
 sg13g2_inv_1 \ring_1001.inv_array[530]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[531] ),
    .A(\ring_1001.inv_in[530] ));
 sg13g2_inv_1 \ring_1001.inv_array[531]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[532] ),
    .A(\ring_1001.inv_in[531] ));
 sg13g2_inv_1 \ring_1001.inv_array[532]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[533] ),
    .A(\ring_1001.inv_in[532] ));
 sg13g2_inv_1 \ring_1001.inv_array[533]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[534] ),
    .A(\ring_1001.inv_in[533] ));
 sg13g2_inv_1 \ring_1001.inv_array[534]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[535] ),
    .A(\ring_1001.inv_in[534] ));
 sg13g2_inv_1 \ring_1001.inv_array[535]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[536] ),
    .A(\ring_1001.inv_in[535] ));
 sg13g2_inv_1 \ring_1001.inv_array[536]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[537] ),
    .A(\ring_1001.inv_in[536] ));
 sg13g2_inv_1 \ring_1001.inv_array[537]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[538] ),
    .A(\ring_1001.inv_in[537] ));
 sg13g2_inv_1 \ring_1001.inv_array[538]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[539] ),
    .A(\ring_1001.inv_in[538] ));
 sg13g2_inv_1 \ring_1001.inv_array[539]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[540] ),
    .A(\ring_1001.inv_in[539] ));
 sg13g2_inv_1 \ring_1001.inv_array[53]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[54] ),
    .A(\ring_1001.inv_in[53] ));
 sg13g2_inv_1 \ring_1001.inv_array[540]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[541] ),
    .A(\ring_1001.inv_in[540] ));
 sg13g2_inv_1 \ring_1001.inv_array[541]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[542] ),
    .A(\ring_1001.inv_in[541] ));
 sg13g2_inv_1 \ring_1001.inv_array[542]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[543] ),
    .A(\ring_1001.inv_in[542] ));
 sg13g2_inv_1 \ring_1001.inv_array[543]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[544] ),
    .A(\ring_1001.inv_in[543] ));
 sg13g2_inv_1 \ring_1001.inv_array[544]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[545] ),
    .A(\ring_1001.inv_in[544] ));
 sg13g2_inv_1 \ring_1001.inv_array[545]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[546] ),
    .A(\ring_1001.inv_in[545] ));
 sg13g2_inv_1 \ring_1001.inv_array[546]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[547] ),
    .A(\ring_1001.inv_in[546] ));
 sg13g2_inv_1 \ring_1001.inv_array[547]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[548] ),
    .A(\ring_1001.inv_in[547] ));
 sg13g2_inv_1 \ring_1001.inv_array[548]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[549] ),
    .A(\ring_1001.inv_in[548] ));
 sg13g2_inv_1 \ring_1001.inv_array[549]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[550] ),
    .A(\ring_1001.inv_in[549] ));
 sg13g2_inv_1 \ring_1001.inv_array[54]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[55] ),
    .A(\ring_1001.inv_in[54] ));
 sg13g2_inv_1 \ring_1001.inv_array[550]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[551] ),
    .A(\ring_1001.inv_in[550] ));
 sg13g2_inv_1 \ring_1001.inv_array[551]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[552] ),
    .A(\ring_1001.inv_in[551] ));
 sg13g2_inv_1 \ring_1001.inv_array[552]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[553] ),
    .A(\ring_1001.inv_in[552] ));
 sg13g2_inv_1 \ring_1001.inv_array[553]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[554] ),
    .A(\ring_1001.inv_in[553] ));
 sg13g2_inv_1 \ring_1001.inv_array[554]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[555] ),
    .A(\ring_1001.inv_in[554] ));
 sg13g2_inv_1 \ring_1001.inv_array[555]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[556] ),
    .A(\ring_1001.inv_in[555] ));
 sg13g2_inv_1 \ring_1001.inv_array[556]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[557] ),
    .A(\ring_1001.inv_in[556] ));
 sg13g2_inv_1 \ring_1001.inv_array[557]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[558] ),
    .A(\ring_1001.inv_in[557] ));
 sg13g2_inv_1 \ring_1001.inv_array[558]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[559] ),
    .A(\ring_1001.inv_in[558] ));
 sg13g2_inv_1 \ring_1001.inv_array[559]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[560] ),
    .A(\ring_1001.inv_in[559] ));
 sg13g2_inv_1 \ring_1001.inv_array[55]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[56] ),
    .A(\ring_1001.inv_in[55] ));
 sg13g2_inv_1 \ring_1001.inv_array[560]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[561] ),
    .A(\ring_1001.inv_in[560] ));
 sg13g2_inv_1 \ring_1001.inv_array[561]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[562] ),
    .A(\ring_1001.inv_in[561] ));
 sg13g2_inv_1 \ring_1001.inv_array[562]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[563] ),
    .A(\ring_1001.inv_in[562] ));
 sg13g2_inv_1 \ring_1001.inv_array[563]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[564] ),
    .A(\ring_1001.inv_in[563] ));
 sg13g2_inv_1 \ring_1001.inv_array[564]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[565] ),
    .A(\ring_1001.inv_in[564] ));
 sg13g2_inv_1 \ring_1001.inv_array[565]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[566] ),
    .A(\ring_1001.inv_in[565] ));
 sg13g2_inv_1 \ring_1001.inv_array[566]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[567] ),
    .A(\ring_1001.inv_in[566] ));
 sg13g2_inv_1 \ring_1001.inv_array[567]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[568] ),
    .A(\ring_1001.inv_in[567] ));
 sg13g2_inv_1 \ring_1001.inv_array[568]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[569] ),
    .A(\ring_1001.inv_in[568] ));
 sg13g2_inv_1 \ring_1001.inv_array[569]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[570] ),
    .A(\ring_1001.inv_in[569] ));
 sg13g2_inv_1 \ring_1001.inv_array[56]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[57] ),
    .A(\ring_1001.inv_in[56] ));
 sg13g2_inv_1 \ring_1001.inv_array[570]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[571] ),
    .A(\ring_1001.inv_in[570] ));
 sg13g2_inv_1 \ring_1001.inv_array[571]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[572] ),
    .A(\ring_1001.inv_in[571] ));
 sg13g2_inv_1 \ring_1001.inv_array[572]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[573] ),
    .A(\ring_1001.inv_in[572] ));
 sg13g2_inv_1 \ring_1001.inv_array[573]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[574] ),
    .A(\ring_1001.inv_in[573] ));
 sg13g2_inv_1 \ring_1001.inv_array[574]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[575] ),
    .A(\ring_1001.inv_in[574] ));
 sg13g2_inv_1 \ring_1001.inv_array[575]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[576] ),
    .A(\ring_1001.inv_in[575] ));
 sg13g2_inv_1 \ring_1001.inv_array[576]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[577] ),
    .A(\ring_1001.inv_in[576] ));
 sg13g2_inv_1 \ring_1001.inv_array[577]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[578] ),
    .A(\ring_1001.inv_in[577] ));
 sg13g2_inv_1 \ring_1001.inv_array[578]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[579] ),
    .A(\ring_1001.inv_in[578] ));
 sg13g2_inv_1 \ring_1001.inv_array[579]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[580] ),
    .A(\ring_1001.inv_in[579] ));
 sg13g2_inv_1 \ring_1001.inv_array[57]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[58] ),
    .A(\ring_1001.inv_in[57] ));
 sg13g2_inv_1 \ring_1001.inv_array[580]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[581] ),
    .A(\ring_1001.inv_in[580] ));
 sg13g2_inv_1 \ring_1001.inv_array[581]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[582] ),
    .A(\ring_1001.inv_in[581] ));
 sg13g2_inv_1 \ring_1001.inv_array[582]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[583] ),
    .A(\ring_1001.inv_in[582] ));
 sg13g2_inv_1 \ring_1001.inv_array[583]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[584] ),
    .A(\ring_1001.inv_in[583] ));
 sg13g2_inv_1 \ring_1001.inv_array[584]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[585] ),
    .A(\ring_1001.inv_in[584] ));
 sg13g2_inv_1 \ring_1001.inv_array[585]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[586] ),
    .A(\ring_1001.inv_in[585] ));
 sg13g2_inv_1 \ring_1001.inv_array[586]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[587] ),
    .A(\ring_1001.inv_in[586] ));
 sg13g2_inv_1 \ring_1001.inv_array[587]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[588] ),
    .A(\ring_1001.inv_in[587] ));
 sg13g2_inv_1 \ring_1001.inv_array[588]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[589] ),
    .A(\ring_1001.inv_in[588] ));
 sg13g2_inv_1 \ring_1001.inv_array[589]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[590] ),
    .A(\ring_1001.inv_in[589] ));
 sg13g2_inv_1 \ring_1001.inv_array[58]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[59] ),
    .A(\ring_1001.inv_in[58] ));
 sg13g2_inv_1 \ring_1001.inv_array[590]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[591] ),
    .A(\ring_1001.inv_in[590] ));
 sg13g2_inv_1 \ring_1001.inv_array[591]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[592] ),
    .A(\ring_1001.inv_in[591] ));
 sg13g2_inv_1 \ring_1001.inv_array[592]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[593] ),
    .A(\ring_1001.inv_in[592] ));
 sg13g2_inv_1 \ring_1001.inv_array[593]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[594] ),
    .A(\ring_1001.inv_in[593] ));
 sg13g2_inv_1 \ring_1001.inv_array[594]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[595] ),
    .A(\ring_1001.inv_in[594] ));
 sg13g2_inv_1 \ring_1001.inv_array[595]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[596] ),
    .A(\ring_1001.inv_in[595] ));
 sg13g2_inv_1 \ring_1001.inv_array[596]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[597] ),
    .A(\ring_1001.inv_in[596] ));
 sg13g2_inv_1 \ring_1001.inv_array[597]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[598] ),
    .A(\ring_1001.inv_in[597] ));
 sg13g2_inv_1 \ring_1001.inv_array[598]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[599] ),
    .A(\ring_1001.inv_in[598] ));
 sg13g2_inv_1 \ring_1001.inv_array[599]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[600] ),
    .A(\ring_1001.inv_in[599] ));
 sg13g2_inv_1 \ring_1001.inv_array[59]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[60] ),
    .A(\ring_1001.inv_in[59] ));
 sg13g2_inv_1 \ring_1001.inv_array[5]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[6] ),
    .A(\ring_1001.inv_in[5] ));
 sg13g2_inv_1 \ring_1001.inv_array[600]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[601] ),
    .A(\ring_1001.inv_in[600] ));
 sg13g2_inv_1 \ring_1001.inv_array[601]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[602] ),
    .A(\ring_1001.inv_in[601] ));
 sg13g2_inv_1 \ring_1001.inv_array[602]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[603] ),
    .A(\ring_1001.inv_in[602] ));
 sg13g2_inv_1 \ring_1001.inv_array[603]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[604] ),
    .A(\ring_1001.inv_in[603] ));
 sg13g2_inv_1 \ring_1001.inv_array[604]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[605] ),
    .A(\ring_1001.inv_in[604] ));
 sg13g2_inv_1 \ring_1001.inv_array[605]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[606] ),
    .A(\ring_1001.inv_in[605] ));
 sg13g2_inv_1 \ring_1001.inv_array[606]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[607] ),
    .A(\ring_1001.inv_in[606] ));
 sg13g2_inv_1 \ring_1001.inv_array[607]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[608] ),
    .A(\ring_1001.inv_in[607] ));
 sg13g2_inv_1 \ring_1001.inv_array[608]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[609] ),
    .A(\ring_1001.inv_in[608] ));
 sg13g2_inv_1 \ring_1001.inv_array[609]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[610] ),
    .A(\ring_1001.inv_in[609] ));
 sg13g2_inv_1 \ring_1001.inv_array[60]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[61] ),
    .A(\ring_1001.inv_in[60] ));
 sg13g2_inv_1 \ring_1001.inv_array[610]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[611] ),
    .A(\ring_1001.inv_in[610] ));
 sg13g2_inv_1 \ring_1001.inv_array[611]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[612] ),
    .A(\ring_1001.inv_in[611] ));
 sg13g2_inv_1 \ring_1001.inv_array[612]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[613] ),
    .A(\ring_1001.inv_in[612] ));
 sg13g2_inv_1 \ring_1001.inv_array[613]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[614] ),
    .A(\ring_1001.inv_in[613] ));
 sg13g2_inv_1 \ring_1001.inv_array[614]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[615] ),
    .A(\ring_1001.inv_in[614] ));
 sg13g2_inv_1 \ring_1001.inv_array[615]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[616] ),
    .A(\ring_1001.inv_in[615] ));
 sg13g2_inv_1 \ring_1001.inv_array[616]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[617] ),
    .A(\ring_1001.inv_in[616] ));
 sg13g2_inv_1 \ring_1001.inv_array[617]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[618] ),
    .A(\ring_1001.inv_in[617] ));
 sg13g2_inv_1 \ring_1001.inv_array[618]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[619] ),
    .A(\ring_1001.inv_in[618] ));
 sg13g2_inv_1 \ring_1001.inv_array[619]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[620] ),
    .A(\ring_1001.inv_in[619] ));
 sg13g2_inv_1 \ring_1001.inv_array[61]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[62] ),
    .A(\ring_1001.inv_in[61] ));
 sg13g2_inv_1 \ring_1001.inv_array[620]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[621] ),
    .A(\ring_1001.inv_in[620] ));
 sg13g2_inv_1 \ring_1001.inv_array[621]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[622] ),
    .A(\ring_1001.inv_in[621] ));
 sg13g2_inv_1 \ring_1001.inv_array[622]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[623] ),
    .A(\ring_1001.inv_in[622] ));
 sg13g2_inv_1 \ring_1001.inv_array[623]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[624] ),
    .A(\ring_1001.inv_in[623] ));
 sg13g2_inv_1 \ring_1001.inv_array[624]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[625] ),
    .A(\ring_1001.inv_in[624] ));
 sg13g2_inv_1 \ring_1001.inv_array[625]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[626] ),
    .A(\ring_1001.inv_in[625] ));
 sg13g2_inv_1 \ring_1001.inv_array[626]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[627] ),
    .A(\ring_1001.inv_in[626] ));
 sg13g2_inv_1 \ring_1001.inv_array[627]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[628] ),
    .A(\ring_1001.inv_in[627] ));
 sg13g2_inv_1 \ring_1001.inv_array[628]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[629] ),
    .A(\ring_1001.inv_in[628] ));
 sg13g2_inv_1 \ring_1001.inv_array[629]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[630] ),
    .A(\ring_1001.inv_in[629] ));
 sg13g2_inv_1 \ring_1001.inv_array[62]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[63] ),
    .A(\ring_1001.inv_in[62] ));
 sg13g2_inv_1 \ring_1001.inv_array[630]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[631] ),
    .A(\ring_1001.inv_in[630] ));
 sg13g2_inv_1 \ring_1001.inv_array[631]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[632] ),
    .A(\ring_1001.inv_in[631] ));
 sg13g2_inv_1 \ring_1001.inv_array[632]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[633] ),
    .A(\ring_1001.inv_in[632] ));
 sg13g2_inv_1 \ring_1001.inv_array[633]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[634] ),
    .A(\ring_1001.inv_in[633] ));
 sg13g2_inv_1 \ring_1001.inv_array[634]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[635] ),
    .A(\ring_1001.inv_in[634] ));
 sg13g2_inv_1 \ring_1001.inv_array[635]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[636] ),
    .A(\ring_1001.inv_in[635] ));
 sg13g2_inv_1 \ring_1001.inv_array[636]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[637] ),
    .A(\ring_1001.inv_in[636] ));
 sg13g2_inv_1 \ring_1001.inv_array[637]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[638] ),
    .A(\ring_1001.inv_in[637] ));
 sg13g2_inv_1 \ring_1001.inv_array[638]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[639] ),
    .A(\ring_1001.inv_in[638] ));
 sg13g2_inv_1 \ring_1001.inv_array[639]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[640] ),
    .A(\ring_1001.inv_in[639] ));
 sg13g2_inv_1 \ring_1001.inv_array[63]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[64] ),
    .A(\ring_1001.inv_in[63] ));
 sg13g2_inv_1 \ring_1001.inv_array[640]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[641] ),
    .A(\ring_1001.inv_in[640] ));
 sg13g2_inv_1 \ring_1001.inv_array[641]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[642] ),
    .A(\ring_1001.inv_in[641] ));
 sg13g2_inv_1 \ring_1001.inv_array[642]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[643] ),
    .A(\ring_1001.inv_in[642] ));
 sg13g2_inv_1 \ring_1001.inv_array[643]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[644] ),
    .A(\ring_1001.inv_in[643] ));
 sg13g2_inv_1 \ring_1001.inv_array[644]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[645] ),
    .A(\ring_1001.inv_in[644] ));
 sg13g2_inv_1 \ring_1001.inv_array[645]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[646] ),
    .A(\ring_1001.inv_in[645] ));
 sg13g2_inv_1 \ring_1001.inv_array[646]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[647] ),
    .A(\ring_1001.inv_in[646] ));
 sg13g2_inv_1 \ring_1001.inv_array[647]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[648] ),
    .A(\ring_1001.inv_in[647] ));
 sg13g2_inv_1 \ring_1001.inv_array[648]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[649] ),
    .A(\ring_1001.inv_in[648] ));
 sg13g2_inv_1 \ring_1001.inv_array[649]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[650] ),
    .A(\ring_1001.inv_in[649] ));
 sg13g2_inv_1 \ring_1001.inv_array[64]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[65] ),
    .A(\ring_1001.inv_in[64] ));
 sg13g2_inv_1 \ring_1001.inv_array[650]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[651] ),
    .A(\ring_1001.inv_in[650] ));
 sg13g2_inv_1 \ring_1001.inv_array[651]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[652] ),
    .A(\ring_1001.inv_in[651] ));
 sg13g2_inv_1 \ring_1001.inv_array[652]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[653] ),
    .A(\ring_1001.inv_in[652] ));
 sg13g2_inv_1 \ring_1001.inv_array[653]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[654] ),
    .A(\ring_1001.inv_in[653] ));
 sg13g2_inv_1 \ring_1001.inv_array[654]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[655] ),
    .A(\ring_1001.inv_in[654] ));
 sg13g2_inv_1 \ring_1001.inv_array[655]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[656] ),
    .A(\ring_1001.inv_in[655] ));
 sg13g2_inv_1 \ring_1001.inv_array[656]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[657] ),
    .A(\ring_1001.inv_in[656] ));
 sg13g2_inv_1 \ring_1001.inv_array[657]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[658] ),
    .A(\ring_1001.inv_in[657] ));
 sg13g2_inv_1 \ring_1001.inv_array[658]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[659] ),
    .A(\ring_1001.inv_in[658] ));
 sg13g2_inv_1 \ring_1001.inv_array[659]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[660] ),
    .A(\ring_1001.inv_in[659] ));
 sg13g2_inv_1 \ring_1001.inv_array[65]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[66] ),
    .A(\ring_1001.inv_in[65] ));
 sg13g2_inv_1 \ring_1001.inv_array[660]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[661] ),
    .A(\ring_1001.inv_in[660] ));
 sg13g2_inv_1 \ring_1001.inv_array[661]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[662] ),
    .A(\ring_1001.inv_in[661] ));
 sg13g2_inv_1 \ring_1001.inv_array[662]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[663] ),
    .A(\ring_1001.inv_in[662] ));
 sg13g2_inv_1 \ring_1001.inv_array[663]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[664] ),
    .A(\ring_1001.inv_in[663] ));
 sg13g2_inv_1 \ring_1001.inv_array[664]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[665] ),
    .A(\ring_1001.inv_in[664] ));
 sg13g2_inv_1 \ring_1001.inv_array[665]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[666] ),
    .A(\ring_1001.inv_in[665] ));
 sg13g2_inv_1 \ring_1001.inv_array[666]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[667] ),
    .A(\ring_1001.inv_in[666] ));
 sg13g2_inv_1 \ring_1001.inv_array[667]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[668] ),
    .A(\ring_1001.inv_in[667] ));
 sg13g2_inv_1 \ring_1001.inv_array[668]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[669] ),
    .A(\ring_1001.inv_in[668] ));
 sg13g2_inv_1 \ring_1001.inv_array[669]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[670] ),
    .A(\ring_1001.inv_in[669] ));
 sg13g2_inv_1 \ring_1001.inv_array[66]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[67] ),
    .A(\ring_1001.inv_in[66] ));
 sg13g2_inv_1 \ring_1001.inv_array[670]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[671] ),
    .A(\ring_1001.inv_in[670] ));
 sg13g2_inv_1 \ring_1001.inv_array[671]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[672] ),
    .A(\ring_1001.inv_in[671] ));
 sg13g2_inv_1 \ring_1001.inv_array[672]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[673] ),
    .A(\ring_1001.inv_in[672] ));
 sg13g2_inv_1 \ring_1001.inv_array[673]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[674] ),
    .A(\ring_1001.inv_in[673] ));
 sg13g2_inv_1 \ring_1001.inv_array[674]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[675] ),
    .A(\ring_1001.inv_in[674] ));
 sg13g2_inv_1 \ring_1001.inv_array[675]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[676] ),
    .A(\ring_1001.inv_in[675] ));
 sg13g2_inv_1 \ring_1001.inv_array[676]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[677] ),
    .A(\ring_1001.inv_in[676] ));
 sg13g2_inv_1 \ring_1001.inv_array[677]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[678] ),
    .A(\ring_1001.inv_in[677] ));
 sg13g2_inv_1 \ring_1001.inv_array[678]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[679] ),
    .A(\ring_1001.inv_in[678] ));
 sg13g2_inv_1 \ring_1001.inv_array[679]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[680] ),
    .A(\ring_1001.inv_in[679] ));
 sg13g2_inv_1 \ring_1001.inv_array[67]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[68] ),
    .A(\ring_1001.inv_in[67] ));
 sg13g2_inv_1 \ring_1001.inv_array[680]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[681] ),
    .A(\ring_1001.inv_in[680] ));
 sg13g2_inv_1 \ring_1001.inv_array[681]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[682] ),
    .A(\ring_1001.inv_in[681] ));
 sg13g2_inv_1 \ring_1001.inv_array[682]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[683] ),
    .A(\ring_1001.inv_in[682] ));
 sg13g2_inv_1 \ring_1001.inv_array[683]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[684] ),
    .A(\ring_1001.inv_in[683] ));
 sg13g2_inv_1 \ring_1001.inv_array[684]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[685] ),
    .A(\ring_1001.inv_in[684] ));
 sg13g2_inv_1 \ring_1001.inv_array[685]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[686] ),
    .A(\ring_1001.inv_in[685] ));
 sg13g2_inv_1 \ring_1001.inv_array[686]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[687] ),
    .A(\ring_1001.inv_in[686] ));
 sg13g2_inv_1 \ring_1001.inv_array[687]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[688] ),
    .A(\ring_1001.inv_in[687] ));
 sg13g2_inv_1 \ring_1001.inv_array[688]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[689] ),
    .A(\ring_1001.inv_in[688] ));
 sg13g2_inv_1 \ring_1001.inv_array[689]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[690] ),
    .A(\ring_1001.inv_in[689] ));
 sg13g2_inv_1 \ring_1001.inv_array[68]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[69] ),
    .A(\ring_1001.inv_in[68] ));
 sg13g2_inv_1 \ring_1001.inv_array[690]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[691] ),
    .A(\ring_1001.inv_in[690] ));
 sg13g2_inv_1 \ring_1001.inv_array[691]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[692] ),
    .A(\ring_1001.inv_in[691] ));
 sg13g2_inv_1 \ring_1001.inv_array[692]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[693] ),
    .A(\ring_1001.inv_in[692] ));
 sg13g2_inv_1 \ring_1001.inv_array[693]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[694] ),
    .A(\ring_1001.inv_in[693] ));
 sg13g2_inv_1 \ring_1001.inv_array[694]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[695] ),
    .A(\ring_1001.inv_in[694] ));
 sg13g2_inv_1 \ring_1001.inv_array[695]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[696] ),
    .A(\ring_1001.inv_in[695] ));
 sg13g2_inv_1 \ring_1001.inv_array[696]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[697] ),
    .A(\ring_1001.inv_in[696] ));
 sg13g2_inv_1 \ring_1001.inv_array[697]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[698] ),
    .A(\ring_1001.inv_in[697] ));
 sg13g2_inv_1 \ring_1001.inv_array[698]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[699] ),
    .A(\ring_1001.inv_in[698] ));
 sg13g2_inv_1 \ring_1001.inv_array[699]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[700] ),
    .A(\ring_1001.inv_in[699] ));
 sg13g2_inv_1 \ring_1001.inv_array[69]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[70] ),
    .A(\ring_1001.inv_in[69] ));
 sg13g2_inv_1 \ring_1001.inv_array[6]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[7] ),
    .A(\ring_1001.inv_in[6] ));
 sg13g2_inv_1 \ring_1001.inv_array[700]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[701] ),
    .A(\ring_1001.inv_in[700] ));
 sg13g2_inv_1 \ring_1001.inv_array[701]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[702] ),
    .A(\ring_1001.inv_in[701] ));
 sg13g2_inv_1 \ring_1001.inv_array[702]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[703] ),
    .A(\ring_1001.inv_in[702] ));
 sg13g2_inv_1 \ring_1001.inv_array[703]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[704] ),
    .A(\ring_1001.inv_in[703] ));
 sg13g2_inv_1 \ring_1001.inv_array[704]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[705] ),
    .A(\ring_1001.inv_in[704] ));
 sg13g2_inv_1 \ring_1001.inv_array[705]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[706] ),
    .A(\ring_1001.inv_in[705] ));
 sg13g2_inv_1 \ring_1001.inv_array[706]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[707] ),
    .A(\ring_1001.inv_in[706] ));
 sg13g2_inv_1 \ring_1001.inv_array[707]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[708] ),
    .A(\ring_1001.inv_in[707] ));
 sg13g2_inv_1 \ring_1001.inv_array[708]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[709] ),
    .A(\ring_1001.inv_in[708] ));
 sg13g2_inv_1 \ring_1001.inv_array[709]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[710] ),
    .A(\ring_1001.inv_in[709] ));
 sg13g2_inv_1 \ring_1001.inv_array[70]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[71] ),
    .A(\ring_1001.inv_in[70] ));
 sg13g2_inv_1 \ring_1001.inv_array[710]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[711] ),
    .A(\ring_1001.inv_in[710] ));
 sg13g2_inv_1 \ring_1001.inv_array[711]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[712] ),
    .A(\ring_1001.inv_in[711] ));
 sg13g2_inv_1 \ring_1001.inv_array[712]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[713] ),
    .A(\ring_1001.inv_in[712] ));
 sg13g2_inv_1 \ring_1001.inv_array[713]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[714] ),
    .A(\ring_1001.inv_in[713] ));
 sg13g2_inv_1 \ring_1001.inv_array[714]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[715] ),
    .A(\ring_1001.inv_in[714] ));
 sg13g2_inv_1 \ring_1001.inv_array[715]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[716] ),
    .A(\ring_1001.inv_in[715] ));
 sg13g2_inv_1 \ring_1001.inv_array[716]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[717] ),
    .A(\ring_1001.inv_in[716] ));
 sg13g2_inv_1 \ring_1001.inv_array[717]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[718] ),
    .A(\ring_1001.inv_in[717] ));
 sg13g2_inv_1 \ring_1001.inv_array[718]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[719] ),
    .A(\ring_1001.inv_in[718] ));
 sg13g2_inv_1 \ring_1001.inv_array[719]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[720] ),
    .A(\ring_1001.inv_in[719] ));
 sg13g2_inv_1 \ring_1001.inv_array[71]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[72] ),
    .A(\ring_1001.inv_in[71] ));
 sg13g2_inv_1 \ring_1001.inv_array[720]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[721] ),
    .A(\ring_1001.inv_in[720] ));
 sg13g2_inv_1 \ring_1001.inv_array[721]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[722] ),
    .A(\ring_1001.inv_in[721] ));
 sg13g2_inv_1 \ring_1001.inv_array[722]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[723] ),
    .A(\ring_1001.inv_in[722] ));
 sg13g2_inv_1 \ring_1001.inv_array[723]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[724] ),
    .A(\ring_1001.inv_in[723] ));
 sg13g2_inv_1 \ring_1001.inv_array[724]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[725] ),
    .A(\ring_1001.inv_in[724] ));
 sg13g2_inv_1 \ring_1001.inv_array[725]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[726] ),
    .A(\ring_1001.inv_in[725] ));
 sg13g2_inv_1 \ring_1001.inv_array[726]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[727] ),
    .A(\ring_1001.inv_in[726] ));
 sg13g2_inv_1 \ring_1001.inv_array[727]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[728] ),
    .A(\ring_1001.inv_in[727] ));
 sg13g2_inv_1 \ring_1001.inv_array[728]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[729] ),
    .A(\ring_1001.inv_in[728] ));
 sg13g2_inv_1 \ring_1001.inv_array[729]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[730] ),
    .A(\ring_1001.inv_in[729] ));
 sg13g2_inv_1 \ring_1001.inv_array[72]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[73] ),
    .A(\ring_1001.inv_in[72] ));
 sg13g2_inv_1 \ring_1001.inv_array[730]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[731] ),
    .A(\ring_1001.inv_in[730] ));
 sg13g2_inv_1 \ring_1001.inv_array[731]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[732] ),
    .A(\ring_1001.inv_in[731] ));
 sg13g2_inv_1 \ring_1001.inv_array[732]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[733] ),
    .A(\ring_1001.inv_in[732] ));
 sg13g2_inv_1 \ring_1001.inv_array[733]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[734] ),
    .A(\ring_1001.inv_in[733] ));
 sg13g2_inv_1 \ring_1001.inv_array[734]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[735] ),
    .A(\ring_1001.inv_in[734] ));
 sg13g2_inv_1 \ring_1001.inv_array[735]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[736] ),
    .A(\ring_1001.inv_in[735] ));
 sg13g2_inv_1 \ring_1001.inv_array[736]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[737] ),
    .A(\ring_1001.inv_in[736] ));
 sg13g2_inv_1 \ring_1001.inv_array[737]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[738] ),
    .A(\ring_1001.inv_in[737] ));
 sg13g2_inv_1 \ring_1001.inv_array[738]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[739] ),
    .A(\ring_1001.inv_in[738] ));
 sg13g2_inv_1 \ring_1001.inv_array[739]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[740] ),
    .A(\ring_1001.inv_in[739] ));
 sg13g2_inv_1 \ring_1001.inv_array[73]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[74] ),
    .A(\ring_1001.inv_in[73] ));
 sg13g2_inv_1 \ring_1001.inv_array[740]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[741] ),
    .A(\ring_1001.inv_in[740] ));
 sg13g2_inv_1 \ring_1001.inv_array[741]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[742] ),
    .A(\ring_1001.inv_in[741] ));
 sg13g2_inv_1 \ring_1001.inv_array[742]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[743] ),
    .A(\ring_1001.inv_in[742] ));
 sg13g2_inv_1 \ring_1001.inv_array[743]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[744] ),
    .A(\ring_1001.inv_in[743] ));
 sg13g2_inv_1 \ring_1001.inv_array[744]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[745] ),
    .A(\ring_1001.inv_in[744] ));
 sg13g2_inv_1 \ring_1001.inv_array[745]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[746] ),
    .A(\ring_1001.inv_in[745] ));
 sg13g2_inv_1 \ring_1001.inv_array[746]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[747] ),
    .A(\ring_1001.inv_in[746] ));
 sg13g2_inv_1 \ring_1001.inv_array[747]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[748] ),
    .A(\ring_1001.inv_in[747] ));
 sg13g2_inv_1 \ring_1001.inv_array[748]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[749] ),
    .A(\ring_1001.inv_in[748] ));
 sg13g2_inv_1 \ring_1001.inv_array[749]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[750] ),
    .A(\ring_1001.inv_in[749] ));
 sg13g2_inv_1 \ring_1001.inv_array[74]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[75] ),
    .A(\ring_1001.inv_in[74] ));
 sg13g2_inv_1 \ring_1001.inv_array[750]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[751] ),
    .A(\ring_1001.inv_in[750] ));
 sg13g2_inv_1 \ring_1001.inv_array[751]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[752] ),
    .A(\ring_1001.inv_in[751] ));
 sg13g2_inv_1 \ring_1001.inv_array[752]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[753] ),
    .A(\ring_1001.inv_in[752] ));
 sg13g2_inv_1 \ring_1001.inv_array[753]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[754] ),
    .A(\ring_1001.inv_in[753] ));
 sg13g2_inv_1 \ring_1001.inv_array[754]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[755] ),
    .A(\ring_1001.inv_in[754] ));
 sg13g2_inv_1 \ring_1001.inv_array[755]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[756] ),
    .A(\ring_1001.inv_in[755] ));
 sg13g2_inv_1 \ring_1001.inv_array[756]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[757] ),
    .A(\ring_1001.inv_in[756] ));
 sg13g2_inv_1 \ring_1001.inv_array[757]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[758] ),
    .A(\ring_1001.inv_in[757] ));
 sg13g2_inv_1 \ring_1001.inv_array[758]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[759] ),
    .A(\ring_1001.inv_in[758] ));
 sg13g2_inv_1 \ring_1001.inv_array[759]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[760] ),
    .A(\ring_1001.inv_in[759] ));
 sg13g2_inv_1 \ring_1001.inv_array[75]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[76] ),
    .A(\ring_1001.inv_in[75] ));
 sg13g2_inv_1 \ring_1001.inv_array[760]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[761] ),
    .A(\ring_1001.inv_in[760] ));
 sg13g2_inv_1 \ring_1001.inv_array[761]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[762] ),
    .A(\ring_1001.inv_in[761] ));
 sg13g2_inv_1 \ring_1001.inv_array[762]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[763] ),
    .A(\ring_1001.inv_in[762] ));
 sg13g2_inv_1 \ring_1001.inv_array[763]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[764] ),
    .A(\ring_1001.inv_in[763] ));
 sg13g2_inv_1 \ring_1001.inv_array[764]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[765] ),
    .A(\ring_1001.inv_in[764] ));
 sg13g2_inv_1 \ring_1001.inv_array[765]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[766] ),
    .A(\ring_1001.inv_in[765] ));
 sg13g2_inv_1 \ring_1001.inv_array[766]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[767] ),
    .A(\ring_1001.inv_in[766] ));
 sg13g2_inv_1 \ring_1001.inv_array[767]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[768] ),
    .A(\ring_1001.inv_in[767] ));
 sg13g2_inv_1 \ring_1001.inv_array[768]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[769] ),
    .A(\ring_1001.inv_in[768] ));
 sg13g2_inv_1 \ring_1001.inv_array[769]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[770] ),
    .A(\ring_1001.inv_in[769] ));
 sg13g2_inv_1 \ring_1001.inv_array[76]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[77] ),
    .A(\ring_1001.inv_in[76] ));
 sg13g2_inv_1 \ring_1001.inv_array[770]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[771] ),
    .A(\ring_1001.inv_in[770] ));
 sg13g2_inv_1 \ring_1001.inv_array[771]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[772] ),
    .A(\ring_1001.inv_in[771] ));
 sg13g2_inv_1 \ring_1001.inv_array[772]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[773] ),
    .A(\ring_1001.inv_in[772] ));
 sg13g2_inv_1 \ring_1001.inv_array[773]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[774] ),
    .A(\ring_1001.inv_in[773] ));
 sg13g2_inv_1 \ring_1001.inv_array[774]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[775] ),
    .A(\ring_1001.inv_in[774] ));
 sg13g2_inv_1 \ring_1001.inv_array[775]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[776] ),
    .A(\ring_1001.inv_in[775] ));
 sg13g2_inv_1 \ring_1001.inv_array[776]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[777] ),
    .A(\ring_1001.inv_in[776] ));
 sg13g2_inv_1 \ring_1001.inv_array[777]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[778] ),
    .A(\ring_1001.inv_in[777] ));
 sg13g2_inv_1 \ring_1001.inv_array[778]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[779] ),
    .A(\ring_1001.inv_in[778] ));
 sg13g2_inv_1 \ring_1001.inv_array[779]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[780] ),
    .A(\ring_1001.inv_in[779] ));
 sg13g2_inv_1 \ring_1001.inv_array[77]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[78] ),
    .A(\ring_1001.inv_in[77] ));
 sg13g2_inv_1 \ring_1001.inv_array[780]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[781] ),
    .A(\ring_1001.inv_in[780] ));
 sg13g2_inv_1 \ring_1001.inv_array[781]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[782] ),
    .A(\ring_1001.inv_in[781] ));
 sg13g2_inv_1 \ring_1001.inv_array[782]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[783] ),
    .A(\ring_1001.inv_in[782] ));
 sg13g2_inv_1 \ring_1001.inv_array[783]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[784] ),
    .A(\ring_1001.inv_in[783] ));
 sg13g2_inv_1 \ring_1001.inv_array[784]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[785] ),
    .A(\ring_1001.inv_in[784] ));
 sg13g2_inv_1 \ring_1001.inv_array[785]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[786] ),
    .A(\ring_1001.inv_in[785] ));
 sg13g2_inv_1 \ring_1001.inv_array[786]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[787] ),
    .A(\ring_1001.inv_in[786] ));
 sg13g2_inv_1 \ring_1001.inv_array[787]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[788] ),
    .A(\ring_1001.inv_in[787] ));
 sg13g2_inv_1 \ring_1001.inv_array[788]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[789] ),
    .A(\ring_1001.inv_in[788] ));
 sg13g2_inv_1 \ring_1001.inv_array[789]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[790] ),
    .A(\ring_1001.inv_in[789] ));
 sg13g2_inv_1 \ring_1001.inv_array[78]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[79] ),
    .A(\ring_1001.inv_in[78] ));
 sg13g2_inv_1 \ring_1001.inv_array[790]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[791] ),
    .A(\ring_1001.inv_in[790] ));
 sg13g2_inv_1 \ring_1001.inv_array[791]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[792] ),
    .A(\ring_1001.inv_in[791] ));
 sg13g2_inv_1 \ring_1001.inv_array[792]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[793] ),
    .A(\ring_1001.inv_in[792] ));
 sg13g2_inv_1 \ring_1001.inv_array[793]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[794] ),
    .A(\ring_1001.inv_in[793] ));
 sg13g2_inv_1 \ring_1001.inv_array[794]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[795] ),
    .A(\ring_1001.inv_in[794] ));
 sg13g2_inv_1 \ring_1001.inv_array[795]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[796] ),
    .A(\ring_1001.inv_in[795] ));
 sg13g2_inv_1 \ring_1001.inv_array[796]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[797] ),
    .A(\ring_1001.inv_in[796] ));
 sg13g2_inv_1 \ring_1001.inv_array[797]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[798] ),
    .A(\ring_1001.inv_in[797] ));
 sg13g2_inv_1 \ring_1001.inv_array[798]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[799] ),
    .A(\ring_1001.inv_in[798] ));
 sg13g2_inv_1 \ring_1001.inv_array[799]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[800] ),
    .A(\ring_1001.inv_in[799] ));
 sg13g2_inv_1 \ring_1001.inv_array[79]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[80] ),
    .A(\ring_1001.inv_in[79] ));
 sg13g2_inv_1 \ring_1001.inv_array[7]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[8] ),
    .A(\ring_1001.inv_in[7] ));
 sg13g2_inv_1 \ring_1001.inv_array[800]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[801] ),
    .A(\ring_1001.inv_in[800] ));
 sg13g2_inv_1 \ring_1001.inv_array[801]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[802] ),
    .A(\ring_1001.inv_in[801] ));
 sg13g2_inv_1 \ring_1001.inv_array[802]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[803] ),
    .A(\ring_1001.inv_in[802] ));
 sg13g2_inv_1 \ring_1001.inv_array[803]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[804] ),
    .A(\ring_1001.inv_in[803] ));
 sg13g2_inv_1 \ring_1001.inv_array[804]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[805] ),
    .A(\ring_1001.inv_in[804] ));
 sg13g2_inv_1 \ring_1001.inv_array[805]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[806] ),
    .A(\ring_1001.inv_in[805] ));
 sg13g2_inv_1 \ring_1001.inv_array[806]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[807] ),
    .A(\ring_1001.inv_in[806] ));
 sg13g2_inv_1 \ring_1001.inv_array[807]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[808] ),
    .A(\ring_1001.inv_in[807] ));
 sg13g2_inv_1 \ring_1001.inv_array[808]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[809] ),
    .A(\ring_1001.inv_in[808] ));
 sg13g2_inv_1 \ring_1001.inv_array[809]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[810] ),
    .A(\ring_1001.inv_in[809] ));
 sg13g2_inv_1 \ring_1001.inv_array[80]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[81] ),
    .A(\ring_1001.inv_in[80] ));
 sg13g2_inv_1 \ring_1001.inv_array[810]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[811] ),
    .A(\ring_1001.inv_in[810] ));
 sg13g2_inv_1 \ring_1001.inv_array[811]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[812] ),
    .A(\ring_1001.inv_in[811] ));
 sg13g2_inv_1 \ring_1001.inv_array[812]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[813] ),
    .A(\ring_1001.inv_in[812] ));
 sg13g2_inv_1 \ring_1001.inv_array[813]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[814] ),
    .A(\ring_1001.inv_in[813] ));
 sg13g2_inv_1 \ring_1001.inv_array[814]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[815] ),
    .A(\ring_1001.inv_in[814] ));
 sg13g2_inv_1 \ring_1001.inv_array[815]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[816] ),
    .A(\ring_1001.inv_in[815] ));
 sg13g2_inv_1 \ring_1001.inv_array[816]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[817] ),
    .A(\ring_1001.inv_in[816] ));
 sg13g2_inv_1 \ring_1001.inv_array[817]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[818] ),
    .A(\ring_1001.inv_in[817] ));
 sg13g2_inv_1 \ring_1001.inv_array[818]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[819] ),
    .A(\ring_1001.inv_in[818] ));
 sg13g2_inv_1 \ring_1001.inv_array[819]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[820] ),
    .A(\ring_1001.inv_in[819] ));
 sg13g2_inv_1 \ring_1001.inv_array[81]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[82] ),
    .A(\ring_1001.inv_in[81] ));
 sg13g2_inv_1 \ring_1001.inv_array[820]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[821] ),
    .A(\ring_1001.inv_in[820] ));
 sg13g2_inv_1 \ring_1001.inv_array[821]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[822] ),
    .A(\ring_1001.inv_in[821] ));
 sg13g2_inv_1 \ring_1001.inv_array[822]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[823] ),
    .A(\ring_1001.inv_in[822] ));
 sg13g2_inv_1 \ring_1001.inv_array[823]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[824] ),
    .A(\ring_1001.inv_in[823] ));
 sg13g2_inv_1 \ring_1001.inv_array[824]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[825] ),
    .A(\ring_1001.inv_in[824] ));
 sg13g2_inv_1 \ring_1001.inv_array[825]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[826] ),
    .A(\ring_1001.inv_in[825] ));
 sg13g2_inv_1 \ring_1001.inv_array[826]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[827] ),
    .A(\ring_1001.inv_in[826] ));
 sg13g2_inv_1 \ring_1001.inv_array[827]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[828] ),
    .A(\ring_1001.inv_in[827] ));
 sg13g2_inv_1 \ring_1001.inv_array[828]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[829] ),
    .A(\ring_1001.inv_in[828] ));
 sg13g2_inv_1 \ring_1001.inv_array[829]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[830] ),
    .A(\ring_1001.inv_in[829] ));
 sg13g2_inv_1 \ring_1001.inv_array[82]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[83] ),
    .A(\ring_1001.inv_in[82] ));
 sg13g2_inv_1 \ring_1001.inv_array[830]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[831] ),
    .A(\ring_1001.inv_in[830] ));
 sg13g2_inv_1 \ring_1001.inv_array[831]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[832] ),
    .A(\ring_1001.inv_in[831] ));
 sg13g2_inv_1 \ring_1001.inv_array[832]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[833] ),
    .A(\ring_1001.inv_in[832] ));
 sg13g2_inv_1 \ring_1001.inv_array[833]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[834] ),
    .A(\ring_1001.inv_in[833] ));
 sg13g2_inv_1 \ring_1001.inv_array[834]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[835] ),
    .A(\ring_1001.inv_in[834] ));
 sg13g2_inv_1 \ring_1001.inv_array[835]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[836] ),
    .A(\ring_1001.inv_in[835] ));
 sg13g2_inv_1 \ring_1001.inv_array[836]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[837] ),
    .A(\ring_1001.inv_in[836] ));
 sg13g2_inv_1 \ring_1001.inv_array[837]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[838] ),
    .A(\ring_1001.inv_in[837] ));
 sg13g2_inv_1 \ring_1001.inv_array[838]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[839] ),
    .A(\ring_1001.inv_in[838] ));
 sg13g2_inv_1 \ring_1001.inv_array[839]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[840] ),
    .A(\ring_1001.inv_in[839] ));
 sg13g2_inv_1 \ring_1001.inv_array[83]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[84] ),
    .A(\ring_1001.inv_in[83] ));
 sg13g2_inv_1 \ring_1001.inv_array[840]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[841] ),
    .A(\ring_1001.inv_in[840] ));
 sg13g2_inv_1 \ring_1001.inv_array[841]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[842] ),
    .A(\ring_1001.inv_in[841] ));
 sg13g2_inv_1 \ring_1001.inv_array[842]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[843] ),
    .A(\ring_1001.inv_in[842] ));
 sg13g2_inv_1 \ring_1001.inv_array[843]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[844] ),
    .A(\ring_1001.inv_in[843] ));
 sg13g2_inv_1 \ring_1001.inv_array[844]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[845] ),
    .A(\ring_1001.inv_in[844] ));
 sg13g2_inv_1 \ring_1001.inv_array[845]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[846] ),
    .A(\ring_1001.inv_in[845] ));
 sg13g2_inv_1 \ring_1001.inv_array[846]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[847] ),
    .A(\ring_1001.inv_in[846] ));
 sg13g2_inv_1 \ring_1001.inv_array[847]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[848] ),
    .A(\ring_1001.inv_in[847] ));
 sg13g2_inv_1 \ring_1001.inv_array[848]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[849] ),
    .A(\ring_1001.inv_in[848] ));
 sg13g2_inv_1 \ring_1001.inv_array[849]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[850] ),
    .A(\ring_1001.inv_in[849] ));
 sg13g2_inv_1 \ring_1001.inv_array[84]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[85] ),
    .A(\ring_1001.inv_in[84] ));
 sg13g2_inv_1 \ring_1001.inv_array[850]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[851] ),
    .A(\ring_1001.inv_in[850] ));
 sg13g2_inv_1 \ring_1001.inv_array[851]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[852] ),
    .A(\ring_1001.inv_in[851] ));
 sg13g2_inv_1 \ring_1001.inv_array[852]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[853] ),
    .A(\ring_1001.inv_in[852] ));
 sg13g2_inv_1 \ring_1001.inv_array[853]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[854] ),
    .A(\ring_1001.inv_in[853] ));
 sg13g2_inv_1 \ring_1001.inv_array[854]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[855] ),
    .A(\ring_1001.inv_in[854] ));
 sg13g2_inv_1 \ring_1001.inv_array[855]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[856] ),
    .A(\ring_1001.inv_in[855] ));
 sg13g2_inv_1 \ring_1001.inv_array[856]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[857] ),
    .A(\ring_1001.inv_in[856] ));
 sg13g2_inv_1 \ring_1001.inv_array[857]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[858] ),
    .A(\ring_1001.inv_in[857] ));
 sg13g2_inv_1 \ring_1001.inv_array[858]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[859] ),
    .A(\ring_1001.inv_in[858] ));
 sg13g2_inv_1 \ring_1001.inv_array[859]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[860] ),
    .A(\ring_1001.inv_in[859] ));
 sg13g2_inv_1 \ring_1001.inv_array[85]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[86] ),
    .A(\ring_1001.inv_in[85] ));
 sg13g2_inv_1 \ring_1001.inv_array[860]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[861] ),
    .A(\ring_1001.inv_in[860] ));
 sg13g2_inv_1 \ring_1001.inv_array[861]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[862] ),
    .A(\ring_1001.inv_in[861] ));
 sg13g2_inv_1 \ring_1001.inv_array[862]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[863] ),
    .A(\ring_1001.inv_in[862] ));
 sg13g2_inv_1 \ring_1001.inv_array[863]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[864] ),
    .A(\ring_1001.inv_in[863] ));
 sg13g2_inv_1 \ring_1001.inv_array[864]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[865] ),
    .A(\ring_1001.inv_in[864] ));
 sg13g2_inv_1 \ring_1001.inv_array[865]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[866] ),
    .A(\ring_1001.inv_in[865] ));
 sg13g2_inv_1 \ring_1001.inv_array[866]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[867] ),
    .A(\ring_1001.inv_in[866] ));
 sg13g2_inv_1 \ring_1001.inv_array[867]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[868] ),
    .A(\ring_1001.inv_in[867] ));
 sg13g2_inv_1 \ring_1001.inv_array[868]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[869] ),
    .A(\ring_1001.inv_in[868] ));
 sg13g2_inv_1 \ring_1001.inv_array[869]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[870] ),
    .A(\ring_1001.inv_in[869] ));
 sg13g2_inv_1 \ring_1001.inv_array[86]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[87] ),
    .A(\ring_1001.inv_in[86] ));
 sg13g2_inv_1 \ring_1001.inv_array[870]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[871] ),
    .A(\ring_1001.inv_in[870] ));
 sg13g2_inv_1 \ring_1001.inv_array[871]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[872] ),
    .A(\ring_1001.inv_in[871] ));
 sg13g2_inv_1 \ring_1001.inv_array[872]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[873] ),
    .A(\ring_1001.inv_in[872] ));
 sg13g2_inv_1 \ring_1001.inv_array[873]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[874] ),
    .A(\ring_1001.inv_in[873] ));
 sg13g2_inv_1 \ring_1001.inv_array[874]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[875] ),
    .A(\ring_1001.inv_in[874] ));
 sg13g2_inv_1 \ring_1001.inv_array[875]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[876] ),
    .A(\ring_1001.inv_in[875] ));
 sg13g2_inv_1 \ring_1001.inv_array[876]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[877] ),
    .A(\ring_1001.inv_in[876] ));
 sg13g2_inv_1 \ring_1001.inv_array[877]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[878] ),
    .A(\ring_1001.inv_in[877] ));
 sg13g2_inv_1 \ring_1001.inv_array[878]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[879] ),
    .A(\ring_1001.inv_in[878] ));
 sg13g2_inv_1 \ring_1001.inv_array[879]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[880] ),
    .A(\ring_1001.inv_in[879] ));
 sg13g2_inv_1 \ring_1001.inv_array[87]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[88] ),
    .A(\ring_1001.inv_in[87] ));
 sg13g2_inv_1 \ring_1001.inv_array[880]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[881] ),
    .A(\ring_1001.inv_in[880] ));
 sg13g2_inv_1 \ring_1001.inv_array[881]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[882] ),
    .A(\ring_1001.inv_in[881] ));
 sg13g2_inv_1 \ring_1001.inv_array[882]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[883] ),
    .A(\ring_1001.inv_in[882] ));
 sg13g2_inv_1 \ring_1001.inv_array[883]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[884] ),
    .A(\ring_1001.inv_in[883] ));
 sg13g2_inv_1 \ring_1001.inv_array[884]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[885] ),
    .A(\ring_1001.inv_in[884] ));
 sg13g2_inv_1 \ring_1001.inv_array[885]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[886] ),
    .A(\ring_1001.inv_in[885] ));
 sg13g2_inv_1 \ring_1001.inv_array[886]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[887] ),
    .A(\ring_1001.inv_in[886] ));
 sg13g2_inv_1 \ring_1001.inv_array[887]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[888] ),
    .A(\ring_1001.inv_in[887] ));
 sg13g2_inv_1 \ring_1001.inv_array[888]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[889] ),
    .A(\ring_1001.inv_in[888] ));
 sg13g2_inv_1 \ring_1001.inv_array[889]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[890] ),
    .A(\ring_1001.inv_in[889] ));
 sg13g2_inv_1 \ring_1001.inv_array[88]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[89] ),
    .A(\ring_1001.inv_in[88] ));
 sg13g2_inv_1 \ring_1001.inv_array[890]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[891] ),
    .A(\ring_1001.inv_in[890] ));
 sg13g2_inv_1 \ring_1001.inv_array[891]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[892] ),
    .A(\ring_1001.inv_in[891] ));
 sg13g2_inv_1 \ring_1001.inv_array[892]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[893] ),
    .A(\ring_1001.inv_in[892] ));
 sg13g2_inv_1 \ring_1001.inv_array[893]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[894] ),
    .A(\ring_1001.inv_in[893] ));
 sg13g2_inv_1 \ring_1001.inv_array[894]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[895] ),
    .A(\ring_1001.inv_in[894] ));
 sg13g2_inv_1 \ring_1001.inv_array[895]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[896] ),
    .A(\ring_1001.inv_in[895] ));
 sg13g2_inv_1 \ring_1001.inv_array[896]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[897] ),
    .A(\ring_1001.inv_in[896] ));
 sg13g2_inv_1 \ring_1001.inv_array[897]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[898] ),
    .A(\ring_1001.inv_in[897] ));
 sg13g2_inv_1 \ring_1001.inv_array[898]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[899] ),
    .A(\ring_1001.inv_in[898] ));
 sg13g2_inv_1 \ring_1001.inv_array[899]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[900] ),
    .A(\ring_1001.inv_in[899] ));
 sg13g2_inv_1 \ring_1001.inv_array[89]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[90] ),
    .A(\ring_1001.inv_in[89] ));
 sg13g2_inv_1 \ring_1001.inv_array[8]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[9] ),
    .A(\ring_1001.inv_in[8] ));
 sg13g2_inv_1 \ring_1001.inv_array[900]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[901] ),
    .A(\ring_1001.inv_in[900] ));
 sg13g2_inv_1 \ring_1001.inv_array[901]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[902] ),
    .A(\ring_1001.inv_in[901] ));
 sg13g2_inv_1 \ring_1001.inv_array[902]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[903] ),
    .A(\ring_1001.inv_in[902] ));
 sg13g2_inv_1 \ring_1001.inv_array[903]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[904] ),
    .A(\ring_1001.inv_in[903] ));
 sg13g2_inv_1 \ring_1001.inv_array[904]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[905] ),
    .A(\ring_1001.inv_in[904] ));
 sg13g2_inv_1 \ring_1001.inv_array[905]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[906] ),
    .A(\ring_1001.inv_in[905] ));
 sg13g2_inv_1 \ring_1001.inv_array[906]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[907] ),
    .A(\ring_1001.inv_in[906] ));
 sg13g2_inv_1 \ring_1001.inv_array[907]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[908] ),
    .A(\ring_1001.inv_in[907] ));
 sg13g2_inv_1 \ring_1001.inv_array[908]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[909] ),
    .A(\ring_1001.inv_in[908] ));
 sg13g2_inv_1 \ring_1001.inv_array[909]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[910] ),
    .A(\ring_1001.inv_in[909] ));
 sg13g2_inv_1 \ring_1001.inv_array[90]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[91] ),
    .A(\ring_1001.inv_in[90] ));
 sg13g2_inv_1 \ring_1001.inv_array[910]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[911] ),
    .A(\ring_1001.inv_in[910] ));
 sg13g2_inv_1 \ring_1001.inv_array[911]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[912] ),
    .A(\ring_1001.inv_in[911] ));
 sg13g2_inv_1 \ring_1001.inv_array[912]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[913] ),
    .A(\ring_1001.inv_in[912] ));
 sg13g2_inv_1 \ring_1001.inv_array[913]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[914] ),
    .A(\ring_1001.inv_in[913] ));
 sg13g2_inv_1 \ring_1001.inv_array[914]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[915] ),
    .A(\ring_1001.inv_in[914] ));
 sg13g2_inv_1 \ring_1001.inv_array[915]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[916] ),
    .A(\ring_1001.inv_in[915] ));
 sg13g2_inv_1 \ring_1001.inv_array[916]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[917] ),
    .A(\ring_1001.inv_in[916] ));
 sg13g2_inv_1 \ring_1001.inv_array[917]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[918] ),
    .A(\ring_1001.inv_in[917] ));
 sg13g2_inv_1 \ring_1001.inv_array[918]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[919] ),
    .A(\ring_1001.inv_in[918] ));
 sg13g2_inv_1 \ring_1001.inv_array[919]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[920] ),
    .A(\ring_1001.inv_in[919] ));
 sg13g2_inv_1 \ring_1001.inv_array[91]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[92] ),
    .A(\ring_1001.inv_in[91] ));
 sg13g2_inv_1 \ring_1001.inv_array[920]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[921] ),
    .A(\ring_1001.inv_in[920] ));
 sg13g2_inv_1 \ring_1001.inv_array[921]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[922] ),
    .A(\ring_1001.inv_in[921] ));
 sg13g2_inv_1 \ring_1001.inv_array[922]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[923] ),
    .A(\ring_1001.inv_in[922] ));
 sg13g2_inv_1 \ring_1001.inv_array[923]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[924] ),
    .A(\ring_1001.inv_in[923] ));
 sg13g2_inv_1 \ring_1001.inv_array[924]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[925] ),
    .A(\ring_1001.inv_in[924] ));
 sg13g2_inv_1 \ring_1001.inv_array[925]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[926] ),
    .A(\ring_1001.inv_in[925] ));
 sg13g2_inv_1 \ring_1001.inv_array[926]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[927] ),
    .A(\ring_1001.inv_in[926] ));
 sg13g2_inv_1 \ring_1001.inv_array[927]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[928] ),
    .A(\ring_1001.inv_in[927] ));
 sg13g2_inv_1 \ring_1001.inv_array[928]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[929] ),
    .A(\ring_1001.inv_in[928] ));
 sg13g2_inv_1 \ring_1001.inv_array[929]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[930] ),
    .A(\ring_1001.inv_in[929] ));
 sg13g2_inv_1 \ring_1001.inv_array[92]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[93] ),
    .A(\ring_1001.inv_in[92] ));
 sg13g2_inv_1 \ring_1001.inv_array[930]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[931] ),
    .A(\ring_1001.inv_in[930] ));
 sg13g2_inv_1 \ring_1001.inv_array[931]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[932] ),
    .A(\ring_1001.inv_in[931] ));
 sg13g2_inv_1 \ring_1001.inv_array[932]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[933] ),
    .A(\ring_1001.inv_in[932] ));
 sg13g2_inv_1 \ring_1001.inv_array[933]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[934] ),
    .A(\ring_1001.inv_in[933] ));
 sg13g2_inv_1 \ring_1001.inv_array[934]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[935] ),
    .A(\ring_1001.inv_in[934] ));
 sg13g2_inv_1 \ring_1001.inv_array[935]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[936] ),
    .A(\ring_1001.inv_in[935] ));
 sg13g2_inv_1 \ring_1001.inv_array[936]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[937] ),
    .A(\ring_1001.inv_in[936] ));
 sg13g2_inv_1 \ring_1001.inv_array[937]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[938] ),
    .A(\ring_1001.inv_in[937] ));
 sg13g2_inv_1 \ring_1001.inv_array[938]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[939] ),
    .A(\ring_1001.inv_in[938] ));
 sg13g2_inv_1 \ring_1001.inv_array[939]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[940] ),
    .A(\ring_1001.inv_in[939] ));
 sg13g2_inv_1 \ring_1001.inv_array[93]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[94] ),
    .A(\ring_1001.inv_in[93] ));
 sg13g2_inv_1 \ring_1001.inv_array[940]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[941] ),
    .A(\ring_1001.inv_in[940] ));
 sg13g2_inv_1 \ring_1001.inv_array[941]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[942] ),
    .A(\ring_1001.inv_in[941] ));
 sg13g2_inv_1 \ring_1001.inv_array[942]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[943] ),
    .A(\ring_1001.inv_in[942] ));
 sg13g2_inv_1 \ring_1001.inv_array[943]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[944] ),
    .A(\ring_1001.inv_in[943] ));
 sg13g2_inv_1 \ring_1001.inv_array[944]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[945] ),
    .A(\ring_1001.inv_in[944] ));
 sg13g2_inv_1 \ring_1001.inv_array[945]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[946] ),
    .A(\ring_1001.inv_in[945] ));
 sg13g2_inv_1 \ring_1001.inv_array[946]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[947] ),
    .A(\ring_1001.inv_in[946] ));
 sg13g2_inv_1 \ring_1001.inv_array[947]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[948] ),
    .A(\ring_1001.inv_in[947] ));
 sg13g2_inv_1 \ring_1001.inv_array[948]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[949] ),
    .A(\ring_1001.inv_in[948] ));
 sg13g2_inv_1 \ring_1001.inv_array[949]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[950] ),
    .A(\ring_1001.inv_in[949] ));
 sg13g2_inv_1 \ring_1001.inv_array[94]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[95] ),
    .A(\ring_1001.inv_in[94] ));
 sg13g2_inv_1 \ring_1001.inv_array[950]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[951] ),
    .A(\ring_1001.inv_in[950] ));
 sg13g2_inv_1 \ring_1001.inv_array[951]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[952] ),
    .A(\ring_1001.inv_in[951] ));
 sg13g2_inv_1 \ring_1001.inv_array[952]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[953] ),
    .A(\ring_1001.inv_in[952] ));
 sg13g2_inv_1 \ring_1001.inv_array[953]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[954] ),
    .A(\ring_1001.inv_in[953] ));
 sg13g2_inv_1 \ring_1001.inv_array[954]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[955] ),
    .A(\ring_1001.inv_in[954] ));
 sg13g2_inv_1 \ring_1001.inv_array[955]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[956] ),
    .A(\ring_1001.inv_in[955] ));
 sg13g2_inv_1 \ring_1001.inv_array[956]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[957] ),
    .A(\ring_1001.inv_in[956] ));
 sg13g2_inv_1 \ring_1001.inv_array[957]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[958] ),
    .A(\ring_1001.inv_in[957] ));
 sg13g2_inv_1 \ring_1001.inv_array[958]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[959] ),
    .A(\ring_1001.inv_in[958] ));
 sg13g2_inv_1 \ring_1001.inv_array[959]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[960] ),
    .A(\ring_1001.inv_in[959] ));
 sg13g2_inv_1 \ring_1001.inv_array[95]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[96] ),
    .A(\ring_1001.inv_in[95] ));
 sg13g2_inv_1 \ring_1001.inv_array[960]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[961] ),
    .A(\ring_1001.inv_in[960] ));
 sg13g2_inv_1 \ring_1001.inv_array[961]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[962] ),
    .A(\ring_1001.inv_in[961] ));
 sg13g2_inv_1 \ring_1001.inv_array[962]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[963] ),
    .A(\ring_1001.inv_in[962] ));
 sg13g2_inv_1 \ring_1001.inv_array[963]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[964] ),
    .A(\ring_1001.inv_in[963] ));
 sg13g2_inv_1 \ring_1001.inv_array[964]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[965] ),
    .A(\ring_1001.inv_in[964] ));
 sg13g2_inv_1 \ring_1001.inv_array[965]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[966] ),
    .A(\ring_1001.inv_in[965] ));
 sg13g2_inv_1 \ring_1001.inv_array[966]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[967] ),
    .A(\ring_1001.inv_in[966] ));
 sg13g2_inv_1 \ring_1001.inv_array[967]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[968] ),
    .A(\ring_1001.inv_in[967] ));
 sg13g2_inv_1 \ring_1001.inv_array[968]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[969] ),
    .A(\ring_1001.inv_in[968] ));
 sg13g2_inv_1 \ring_1001.inv_array[969]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[970] ),
    .A(\ring_1001.inv_in[969] ));
 sg13g2_inv_1 \ring_1001.inv_array[96]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[97] ),
    .A(\ring_1001.inv_in[96] ));
 sg13g2_inv_1 \ring_1001.inv_array[970]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[971] ),
    .A(\ring_1001.inv_in[970] ));
 sg13g2_inv_1 \ring_1001.inv_array[971]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[972] ),
    .A(\ring_1001.inv_in[971] ));
 sg13g2_inv_1 \ring_1001.inv_array[972]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[973] ),
    .A(\ring_1001.inv_in[972] ));
 sg13g2_inv_1 \ring_1001.inv_array[973]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[974] ),
    .A(\ring_1001.inv_in[973] ));
 sg13g2_inv_1 \ring_1001.inv_array[974]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[975] ),
    .A(\ring_1001.inv_in[974] ));
 sg13g2_inv_1 \ring_1001.inv_array[975]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[976] ),
    .A(\ring_1001.inv_in[975] ));
 sg13g2_inv_1 \ring_1001.inv_array[976]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[977] ),
    .A(\ring_1001.inv_in[976] ));
 sg13g2_inv_1 \ring_1001.inv_array[977]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[978] ),
    .A(\ring_1001.inv_in[977] ));
 sg13g2_inv_1 \ring_1001.inv_array[978]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[979] ),
    .A(\ring_1001.inv_in[978] ));
 sg13g2_inv_1 \ring_1001.inv_array[979]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[980] ),
    .A(\ring_1001.inv_in[979] ));
 sg13g2_inv_1 \ring_1001.inv_array[97]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[98] ),
    .A(\ring_1001.inv_in[97] ));
 sg13g2_inv_1 \ring_1001.inv_array[980]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[981] ),
    .A(\ring_1001.inv_in[980] ));
 sg13g2_inv_1 \ring_1001.inv_array[981]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[982] ),
    .A(\ring_1001.inv_in[981] ));
 sg13g2_inv_1 \ring_1001.inv_array[982]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[983] ),
    .A(\ring_1001.inv_in[982] ));
 sg13g2_inv_1 \ring_1001.inv_array[983]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[984] ),
    .A(\ring_1001.inv_in[983] ));
 sg13g2_inv_1 \ring_1001.inv_array[984]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[985] ),
    .A(\ring_1001.inv_in[984] ));
 sg13g2_inv_1 \ring_1001.inv_array[985]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[986] ),
    .A(\ring_1001.inv_in[985] ));
 sg13g2_inv_1 \ring_1001.inv_array[986]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[987] ),
    .A(\ring_1001.inv_in[986] ));
 sg13g2_inv_1 \ring_1001.inv_array[987]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[988] ),
    .A(\ring_1001.inv_in[987] ));
 sg13g2_inv_1 \ring_1001.inv_array[988]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[989] ),
    .A(\ring_1001.inv_in[988] ));
 sg13g2_inv_1 \ring_1001.inv_array[989]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[990] ),
    .A(\ring_1001.inv_in[989] ));
 sg13g2_inv_1 \ring_1001.inv_array[98]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[99] ),
    .A(\ring_1001.inv_in[98] ));
 sg13g2_inv_1 \ring_1001.inv_array[990]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[991] ),
    .A(\ring_1001.inv_in[990] ));
 sg13g2_inv_1 \ring_1001.inv_array[991]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[992] ),
    .A(\ring_1001.inv_in[991] ));
 sg13g2_inv_1 \ring_1001.inv_array[992]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[993] ),
    .A(\ring_1001.inv_in[992] ));
 sg13g2_inv_1 \ring_1001.inv_array[993]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[994] ),
    .A(\ring_1001.inv_in[993] ));
 sg13g2_inv_1 \ring_1001.inv_array[994]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[995] ),
    .A(\ring_1001.inv_in[994] ));
 sg13g2_inv_1 \ring_1001.inv_array[995]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[996] ),
    .A(\ring_1001.inv_in[995] ));
 sg13g2_inv_1 \ring_1001.inv_array[996]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[997] ),
    .A(\ring_1001.inv_in[996] ));
 sg13g2_inv_1 \ring_1001.inv_array[997]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[998] ),
    .A(\ring_1001.inv_in[997] ));
 sg13g2_inv_1 \ring_1001.inv_array[998]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[999] ),
    .A(\ring_1001.inv_in[998] ));
 sg13g2_inv_1 \ring_1001.inv_array[999]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[1000] ),
    .A(\ring_1001.inv_in[999] ));
 sg13g2_inv_1 \ring_1001.inv_array[99]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[100] ),
    .A(\ring_1001.inv_in[99] ));
 sg13g2_inv_1 \ring_1001.inv_array[9]/sky_inverter/_0_  (.Y(\ring_1001.inv_in[10] ),
    .A(\ring_1001.inv_in[9] ));
 sg13g2_inv_1 \ring_125.inv_array[0]/sky_inverter/_0_  (.Y(\ring_125.inv_in[1] ),
    .A(c1clock));
 sg13g2_inv_1 \ring_125.inv_array[100]/sky_inverter/_0_  (.Y(\ring_125.inv_in[101] ),
    .A(\ring_125.inv_in[100] ));
 sg13g2_inv_1 \ring_125.inv_array[101]/sky_inverter/_0_  (.Y(\ring_125.inv_in[102] ),
    .A(\ring_125.inv_in[101] ));
 sg13g2_inv_1 \ring_125.inv_array[102]/sky_inverter/_0_  (.Y(\ring_125.inv_in[103] ),
    .A(\ring_125.inv_in[102] ));
 sg13g2_inv_1 \ring_125.inv_array[103]/sky_inverter/_0_  (.Y(\ring_125.inv_in[104] ),
    .A(\ring_125.inv_in[103] ));
 sg13g2_inv_1 \ring_125.inv_array[104]/sky_inverter/_0_  (.Y(\ring_125.inv_in[105] ),
    .A(\ring_125.inv_in[104] ));
 sg13g2_inv_1 \ring_125.inv_array[105]/sky_inverter/_0_  (.Y(\ring_125.inv_in[106] ),
    .A(\ring_125.inv_in[105] ));
 sg13g2_inv_1 \ring_125.inv_array[106]/sky_inverter/_0_  (.Y(\ring_125.inv_in[107] ),
    .A(\ring_125.inv_in[106] ));
 sg13g2_inv_1 \ring_125.inv_array[107]/sky_inverter/_0_  (.Y(\ring_125.inv_in[108] ),
    .A(\ring_125.inv_in[107] ));
 sg13g2_inv_1 \ring_125.inv_array[108]/sky_inverter/_0_  (.Y(\ring_125.inv_in[109] ),
    .A(\ring_125.inv_in[108] ));
 sg13g2_inv_1 \ring_125.inv_array[109]/sky_inverter/_0_  (.Y(\ring_125.inv_in[110] ),
    .A(\ring_125.inv_in[109] ));
 sg13g2_inv_1 \ring_125.inv_array[10]/sky_inverter/_0_  (.Y(\ring_125.inv_in[11] ),
    .A(\ring_125.inv_in[10] ));
 sg13g2_inv_1 \ring_125.inv_array[110]/sky_inverter/_0_  (.Y(\ring_125.inv_in[111] ),
    .A(\ring_125.inv_in[110] ));
 sg13g2_inv_1 \ring_125.inv_array[111]/sky_inverter/_0_  (.Y(\ring_125.inv_in[112] ),
    .A(\ring_125.inv_in[111] ));
 sg13g2_inv_1 \ring_125.inv_array[112]/sky_inverter/_0_  (.Y(\ring_125.inv_in[113] ),
    .A(\ring_125.inv_in[112] ));
 sg13g2_inv_1 \ring_125.inv_array[113]/sky_inverter/_0_  (.Y(\ring_125.inv_in[114] ),
    .A(\ring_125.inv_in[113] ));
 sg13g2_inv_1 \ring_125.inv_array[114]/sky_inverter/_0_  (.Y(\ring_125.inv_in[115] ),
    .A(\ring_125.inv_in[114] ));
 sg13g2_inv_1 \ring_125.inv_array[115]/sky_inverter/_0_  (.Y(\ring_125.inv_in[116] ),
    .A(\ring_125.inv_in[115] ));
 sg13g2_inv_1 \ring_125.inv_array[116]/sky_inverter/_0_  (.Y(\ring_125.inv_in[117] ),
    .A(\ring_125.inv_in[116] ));
 sg13g2_inv_1 \ring_125.inv_array[117]/sky_inverter/_0_  (.Y(\ring_125.inv_in[118] ),
    .A(\ring_125.inv_in[117] ));
 sg13g2_inv_1 \ring_125.inv_array[118]/sky_inverter/_0_  (.Y(\ring_125.inv_in[119] ),
    .A(\ring_125.inv_in[118] ));
 sg13g2_inv_1 \ring_125.inv_array[119]/sky_inverter/_0_  (.Y(\ring_125.inv_in[120] ),
    .A(\ring_125.inv_in[119] ));
 sg13g2_inv_1 \ring_125.inv_array[11]/sky_inverter/_0_  (.Y(\ring_125.inv_in[12] ),
    .A(\ring_125.inv_in[11] ));
 sg13g2_inv_1 \ring_125.inv_array[120]/sky_inverter/_0_  (.Y(\ring_125.inv_in[121] ),
    .A(\ring_125.inv_in[120] ));
 sg13g2_inv_1 \ring_125.inv_array[121]/sky_inverter/_0_  (.Y(\ring_125.inv_in[122] ),
    .A(\ring_125.inv_in[121] ));
 sg13g2_inv_1 \ring_125.inv_array[122]/sky_inverter/_0_  (.Y(\ring_125.inv_in[123] ),
    .A(\ring_125.inv_in[122] ));
 sg13g2_inv_1 \ring_125.inv_array[123]/sky_inverter/_0_  (.Y(\ring_125.inv_in[124] ),
    .A(\ring_125.inv_in[123] ));
 sg13g2_inv_1 \ring_125.inv_array[124]/sky_inverter/_0_  (.Y(\ring_125.inv_out[124] ),
    .A(\ring_125.inv_in[124] ));
 sg13g2_inv_1 \ring_125.inv_array[12]/sky_inverter/_0_  (.Y(\ring_125.inv_in[13] ),
    .A(\ring_125.inv_in[12] ));
 sg13g2_inv_1 \ring_125.inv_array[13]/sky_inverter/_0_  (.Y(\ring_125.inv_in[14] ),
    .A(\ring_125.inv_in[13] ));
 sg13g2_inv_1 \ring_125.inv_array[14]/sky_inverter/_0_  (.Y(\ring_125.inv_in[15] ),
    .A(\ring_125.inv_in[14] ));
 sg13g2_inv_1 \ring_125.inv_array[15]/sky_inverter/_0_  (.Y(\ring_125.inv_in[16] ),
    .A(\ring_125.inv_in[15] ));
 sg13g2_inv_1 \ring_125.inv_array[16]/sky_inverter/_0_  (.Y(\ring_125.inv_in[17] ),
    .A(\ring_125.inv_in[16] ));
 sg13g2_inv_1 \ring_125.inv_array[17]/sky_inverter/_0_  (.Y(\ring_125.inv_in[18] ),
    .A(\ring_125.inv_in[17] ));
 sg13g2_inv_1 \ring_125.inv_array[18]/sky_inverter/_0_  (.Y(\ring_125.inv_in[19] ),
    .A(\ring_125.inv_in[18] ));
 sg13g2_inv_1 \ring_125.inv_array[19]/sky_inverter/_0_  (.Y(\ring_125.inv_in[20] ),
    .A(\ring_125.inv_in[19] ));
 sg13g2_inv_1 \ring_125.inv_array[1]/sky_inverter/_0_  (.Y(\ring_125.inv_in[2] ),
    .A(\ring_125.inv_in[1] ));
 sg13g2_inv_1 \ring_125.inv_array[20]/sky_inverter/_0_  (.Y(\ring_125.inv_in[21] ),
    .A(\ring_125.inv_in[20] ));
 sg13g2_inv_1 \ring_125.inv_array[21]/sky_inverter/_0_  (.Y(\ring_125.inv_in[22] ),
    .A(\ring_125.inv_in[21] ));
 sg13g2_inv_1 \ring_125.inv_array[22]/sky_inverter/_0_  (.Y(\ring_125.inv_in[23] ),
    .A(\ring_125.inv_in[22] ));
 sg13g2_inv_1 \ring_125.inv_array[23]/sky_inverter/_0_  (.Y(\ring_125.inv_in[24] ),
    .A(\ring_125.inv_in[23] ));
 sg13g2_inv_1 \ring_125.inv_array[24]/sky_inverter/_0_  (.Y(\ring_125.inv_in[25] ),
    .A(\ring_125.inv_in[24] ));
 sg13g2_inv_1 \ring_125.inv_array[25]/sky_inverter/_0_  (.Y(\ring_125.inv_in[26] ),
    .A(\ring_125.inv_in[25] ));
 sg13g2_inv_1 \ring_125.inv_array[26]/sky_inverter/_0_  (.Y(\ring_125.inv_in[27] ),
    .A(\ring_125.inv_in[26] ));
 sg13g2_inv_1 \ring_125.inv_array[27]/sky_inverter/_0_  (.Y(\ring_125.inv_in[28] ),
    .A(\ring_125.inv_in[27] ));
 sg13g2_inv_1 \ring_125.inv_array[28]/sky_inverter/_0_  (.Y(\ring_125.inv_in[29] ),
    .A(\ring_125.inv_in[28] ));
 sg13g2_inv_1 \ring_125.inv_array[29]/sky_inverter/_0_  (.Y(\ring_125.inv_in[30] ),
    .A(\ring_125.inv_in[29] ));
 sg13g2_inv_1 \ring_125.inv_array[2]/sky_inverter/_0_  (.Y(\ring_125.inv_in[3] ),
    .A(\ring_125.inv_in[2] ));
 sg13g2_inv_1 \ring_125.inv_array[30]/sky_inverter/_0_  (.Y(\ring_125.inv_in[31] ),
    .A(\ring_125.inv_in[30] ));
 sg13g2_inv_1 \ring_125.inv_array[31]/sky_inverter/_0_  (.Y(\ring_125.inv_in[32] ),
    .A(\ring_125.inv_in[31] ));
 sg13g2_inv_1 \ring_125.inv_array[32]/sky_inverter/_0_  (.Y(\ring_125.inv_in[33] ),
    .A(\ring_125.inv_in[32] ));
 sg13g2_inv_1 \ring_125.inv_array[33]/sky_inverter/_0_  (.Y(\ring_125.inv_in[34] ),
    .A(\ring_125.inv_in[33] ));
 sg13g2_inv_1 \ring_125.inv_array[34]/sky_inverter/_0_  (.Y(\ring_125.inv_in[35] ),
    .A(\ring_125.inv_in[34] ));
 sg13g2_inv_1 \ring_125.inv_array[35]/sky_inverter/_0_  (.Y(\ring_125.inv_in[36] ),
    .A(\ring_125.inv_in[35] ));
 sg13g2_inv_1 \ring_125.inv_array[36]/sky_inverter/_0_  (.Y(\ring_125.inv_in[37] ),
    .A(\ring_125.inv_in[36] ));
 sg13g2_inv_1 \ring_125.inv_array[37]/sky_inverter/_0_  (.Y(\ring_125.inv_in[38] ),
    .A(\ring_125.inv_in[37] ));
 sg13g2_inv_1 \ring_125.inv_array[38]/sky_inverter/_0_  (.Y(\ring_125.inv_in[39] ),
    .A(\ring_125.inv_in[38] ));
 sg13g2_inv_1 \ring_125.inv_array[39]/sky_inverter/_0_  (.Y(\ring_125.inv_in[40] ),
    .A(\ring_125.inv_in[39] ));
 sg13g2_inv_1 \ring_125.inv_array[3]/sky_inverter/_0_  (.Y(\ring_125.inv_in[4] ),
    .A(\ring_125.inv_in[3] ));
 sg13g2_inv_1 \ring_125.inv_array[40]/sky_inverter/_0_  (.Y(\ring_125.inv_in[41] ),
    .A(\ring_125.inv_in[40] ));
 sg13g2_inv_1 \ring_125.inv_array[41]/sky_inverter/_0_  (.Y(\ring_125.inv_in[42] ),
    .A(\ring_125.inv_in[41] ));
 sg13g2_inv_1 \ring_125.inv_array[42]/sky_inverter/_0_  (.Y(\ring_125.inv_in[43] ),
    .A(\ring_125.inv_in[42] ));
 sg13g2_inv_1 \ring_125.inv_array[43]/sky_inverter/_0_  (.Y(\ring_125.inv_in[44] ),
    .A(\ring_125.inv_in[43] ));
 sg13g2_inv_1 \ring_125.inv_array[44]/sky_inverter/_0_  (.Y(\ring_125.inv_in[45] ),
    .A(\ring_125.inv_in[44] ));
 sg13g2_inv_1 \ring_125.inv_array[45]/sky_inverter/_0_  (.Y(\ring_125.inv_in[46] ),
    .A(\ring_125.inv_in[45] ));
 sg13g2_inv_1 \ring_125.inv_array[46]/sky_inverter/_0_  (.Y(\ring_125.inv_in[47] ),
    .A(\ring_125.inv_in[46] ));
 sg13g2_inv_1 \ring_125.inv_array[47]/sky_inverter/_0_  (.Y(\ring_125.inv_in[48] ),
    .A(\ring_125.inv_in[47] ));
 sg13g2_inv_1 \ring_125.inv_array[48]/sky_inverter/_0_  (.Y(\ring_125.inv_in[49] ),
    .A(\ring_125.inv_in[48] ));
 sg13g2_inv_1 \ring_125.inv_array[49]/sky_inverter/_0_  (.Y(\ring_125.inv_in[50] ),
    .A(\ring_125.inv_in[49] ));
 sg13g2_inv_1 \ring_125.inv_array[4]/sky_inverter/_0_  (.Y(\ring_125.inv_in[5] ),
    .A(\ring_125.inv_in[4] ));
 sg13g2_inv_1 \ring_125.inv_array[50]/sky_inverter/_0_  (.Y(\ring_125.inv_in[51] ),
    .A(\ring_125.inv_in[50] ));
 sg13g2_inv_1 \ring_125.inv_array[51]/sky_inverter/_0_  (.Y(\ring_125.inv_in[52] ),
    .A(\ring_125.inv_in[51] ));
 sg13g2_inv_1 \ring_125.inv_array[52]/sky_inverter/_0_  (.Y(\ring_125.inv_in[53] ),
    .A(\ring_125.inv_in[52] ));
 sg13g2_inv_1 \ring_125.inv_array[53]/sky_inverter/_0_  (.Y(\ring_125.inv_in[54] ),
    .A(\ring_125.inv_in[53] ));
 sg13g2_inv_1 \ring_125.inv_array[54]/sky_inverter/_0_  (.Y(\ring_125.inv_in[55] ),
    .A(\ring_125.inv_in[54] ));
 sg13g2_inv_1 \ring_125.inv_array[55]/sky_inverter/_0_  (.Y(\ring_125.inv_in[56] ),
    .A(\ring_125.inv_in[55] ));
 sg13g2_inv_1 \ring_125.inv_array[56]/sky_inverter/_0_  (.Y(\ring_125.inv_in[57] ),
    .A(\ring_125.inv_in[56] ));
 sg13g2_inv_1 \ring_125.inv_array[57]/sky_inverter/_0_  (.Y(\ring_125.inv_in[58] ),
    .A(\ring_125.inv_in[57] ));
 sg13g2_inv_1 \ring_125.inv_array[58]/sky_inverter/_0_  (.Y(\ring_125.inv_in[59] ),
    .A(\ring_125.inv_in[58] ));
 sg13g2_inv_1 \ring_125.inv_array[59]/sky_inverter/_0_  (.Y(\ring_125.inv_in[60] ),
    .A(\ring_125.inv_in[59] ));
 sg13g2_inv_1 \ring_125.inv_array[5]/sky_inverter/_0_  (.Y(\ring_125.inv_in[6] ),
    .A(\ring_125.inv_in[5] ));
 sg13g2_inv_1 \ring_125.inv_array[60]/sky_inverter/_0_  (.Y(\ring_125.inv_in[61] ),
    .A(\ring_125.inv_in[60] ));
 sg13g2_inv_1 \ring_125.inv_array[61]/sky_inverter/_0_  (.Y(\ring_125.inv_in[62] ),
    .A(\ring_125.inv_in[61] ));
 sg13g2_inv_1 \ring_125.inv_array[62]/sky_inverter/_0_  (.Y(\ring_125.inv_in[63] ),
    .A(\ring_125.inv_in[62] ));
 sg13g2_inv_1 \ring_125.inv_array[63]/sky_inverter/_0_  (.Y(\ring_125.inv_in[64] ),
    .A(\ring_125.inv_in[63] ));
 sg13g2_inv_1 \ring_125.inv_array[64]/sky_inverter/_0_  (.Y(\ring_125.inv_in[65] ),
    .A(\ring_125.inv_in[64] ));
 sg13g2_inv_1 \ring_125.inv_array[65]/sky_inverter/_0_  (.Y(\ring_125.inv_in[66] ),
    .A(\ring_125.inv_in[65] ));
 sg13g2_inv_1 \ring_125.inv_array[66]/sky_inverter/_0_  (.Y(\ring_125.inv_in[67] ),
    .A(\ring_125.inv_in[66] ));
 sg13g2_inv_1 \ring_125.inv_array[67]/sky_inverter/_0_  (.Y(\ring_125.inv_in[68] ),
    .A(\ring_125.inv_in[67] ));
 sg13g2_inv_1 \ring_125.inv_array[68]/sky_inverter/_0_  (.Y(\ring_125.inv_in[69] ),
    .A(\ring_125.inv_in[68] ));
 sg13g2_inv_1 \ring_125.inv_array[69]/sky_inverter/_0_  (.Y(\ring_125.inv_in[70] ),
    .A(\ring_125.inv_in[69] ));
 sg13g2_inv_1 \ring_125.inv_array[6]/sky_inverter/_0_  (.Y(\ring_125.inv_in[7] ),
    .A(\ring_125.inv_in[6] ));
 sg13g2_inv_1 \ring_125.inv_array[70]/sky_inverter/_0_  (.Y(\ring_125.inv_in[71] ),
    .A(\ring_125.inv_in[70] ));
 sg13g2_inv_1 \ring_125.inv_array[71]/sky_inverter/_0_  (.Y(\ring_125.inv_in[72] ),
    .A(\ring_125.inv_in[71] ));
 sg13g2_inv_1 \ring_125.inv_array[72]/sky_inverter/_0_  (.Y(\ring_125.inv_in[73] ),
    .A(\ring_125.inv_in[72] ));
 sg13g2_inv_1 \ring_125.inv_array[73]/sky_inverter/_0_  (.Y(\ring_125.inv_in[74] ),
    .A(\ring_125.inv_in[73] ));
 sg13g2_inv_1 \ring_125.inv_array[74]/sky_inverter/_0_  (.Y(\ring_125.inv_in[75] ),
    .A(\ring_125.inv_in[74] ));
 sg13g2_inv_1 \ring_125.inv_array[75]/sky_inverter/_0_  (.Y(\ring_125.inv_in[76] ),
    .A(\ring_125.inv_in[75] ));
 sg13g2_inv_1 \ring_125.inv_array[76]/sky_inverter/_0_  (.Y(\ring_125.inv_in[77] ),
    .A(\ring_125.inv_in[76] ));
 sg13g2_inv_1 \ring_125.inv_array[77]/sky_inverter/_0_  (.Y(\ring_125.inv_in[78] ),
    .A(\ring_125.inv_in[77] ));
 sg13g2_inv_1 \ring_125.inv_array[78]/sky_inverter/_0_  (.Y(\ring_125.inv_in[79] ),
    .A(\ring_125.inv_in[78] ));
 sg13g2_inv_1 \ring_125.inv_array[79]/sky_inverter/_0_  (.Y(\ring_125.inv_in[80] ),
    .A(\ring_125.inv_in[79] ));
 sg13g2_inv_1 \ring_125.inv_array[7]/sky_inverter/_0_  (.Y(\ring_125.inv_in[8] ),
    .A(\ring_125.inv_in[7] ));
 sg13g2_inv_1 \ring_125.inv_array[80]/sky_inverter/_0_  (.Y(\ring_125.inv_in[81] ),
    .A(\ring_125.inv_in[80] ));
 sg13g2_inv_1 \ring_125.inv_array[81]/sky_inverter/_0_  (.Y(\ring_125.inv_in[82] ),
    .A(\ring_125.inv_in[81] ));
 sg13g2_inv_1 \ring_125.inv_array[82]/sky_inverter/_0_  (.Y(\ring_125.inv_in[83] ),
    .A(\ring_125.inv_in[82] ));
 sg13g2_inv_1 \ring_125.inv_array[83]/sky_inverter/_0_  (.Y(\ring_125.inv_in[84] ),
    .A(\ring_125.inv_in[83] ));
 sg13g2_inv_1 \ring_125.inv_array[84]/sky_inverter/_0_  (.Y(\ring_125.inv_in[85] ),
    .A(\ring_125.inv_in[84] ));
 sg13g2_inv_1 \ring_125.inv_array[85]/sky_inverter/_0_  (.Y(\ring_125.inv_in[86] ),
    .A(\ring_125.inv_in[85] ));
 sg13g2_inv_1 \ring_125.inv_array[86]/sky_inverter/_0_  (.Y(\ring_125.inv_in[87] ),
    .A(\ring_125.inv_in[86] ));
 sg13g2_inv_1 \ring_125.inv_array[87]/sky_inverter/_0_  (.Y(\ring_125.inv_in[88] ),
    .A(\ring_125.inv_in[87] ));
 sg13g2_inv_1 \ring_125.inv_array[88]/sky_inverter/_0_  (.Y(\ring_125.inv_in[89] ),
    .A(\ring_125.inv_in[88] ));
 sg13g2_inv_1 \ring_125.inv_array[89]/sky_inverter/_0_  (.Y(\ring_125.inv_in[90] ),
    .A(\ring_125.inv_in[89] ));
 sg13g2_inv_1 \ring_125.inv_array[8]/sky_inverter/_0_  (.Y(\ring_125.inv_in[9] ),
    .A(\ring_125.inv_in[8] ));
 sg13g2_inv_1 \ring_125.inv_array[90]/sky_inverter/_0_  (.Y(\ring_125.inv_in[91] ),
    .A(\ring_125.inv_in[90] ));
 sg13g2_inv_1 \ring_125.inv_array[91]/sky_inverter/_0_  (.Y(\ring_125.inv_in[92] ),
    .A(\ring_125.inv_in[91] ));
 sg13g2_inv_1 \ring_125.inv_array[92]/sky_inverter/_0_  (.Y(\ring_125.inv_in[93] ),
    .A(\ring_125.inv_in[92] ));
 sg13g2_inv_1 \ring_125.inv_array[93]/sky_inverter/_0_  (.Y(\ring_125.inv_in[94] ),
    .A(\ring_125.inv_in[93] ));
 sg13g2_inv_1 \ring_125.inv_array[94]/sky_inverter/_0_  (.Y(\ring_125.inv_in[95] ),
    .A(\ring_125.inv_in[94] ));
 sg13g2_inv_1 \ring_125.inv_array[95]/sky_inverter/_0_  (.Y(\ring_125.inv_in[96] ),
    .A(\ring_125.inv_in[95] ));
 sg13g2_inv_1 \ring_125.inv_array[96]/sky_inverter/_0_  (.Y(\ring_125.inv_in[97] ),
    .A(\ring_125.inv_in[96] ));
 sg13g2_inv_1 \ring_125.inv_array[97]/sky_inverter/_0_  (.Y(\ring_125.inv_in[98] ),
    .A(\ring_125.inv_in[97] ));
 sg13g2_inv_1 \ring_125.inv_array[98]/sky_inverter/_0_  (.Y(\ring_125.inv_in[99] ),
    .A(\ring_125.inv_in[98] ));
 sg13g2_inv_1 \ring_125.inv_array[99]/sky_inverter/_0_  (.Y(\ring_125.inv_in[100] ),
    .A(\ring_125.inv_in[99] ));
 sg13g2_inv_1 \ring_125.inv_array[9]/sky_inverter/_0_  (.Y(\ring_125.inv_in[10] ),
    .A(\ring_125.inv_in[9] ));
 sg13g2_inv_1 \ring_25.inv_array[0]/sky_inverter/_0_  (.Y(\ring_25.inv_in[1] ),
    .A(fast_osc));
 sg13g2_inv_1 \ring_25.inv_array[10]/sky_inverter/_0_  (.Y(\ring_25.inv_in[11] ),
    .A(\ring_25.inv_in[10] ));
 sg13g2_inv_1 \ring_25.inv_array[11]/sky_inverter/_0_  (.Y(\ring_25.inv_in[12] ),
    .A(\ring_25.inv_in[11] ));
 sg13g2_inv_1 \ring_25.inv_array[12]/sky_inverter/_0_  (.Y(\ring_25.inv_in[13] ),
    .A(\ring_25.inv_in[12] ));
 sg13g2_inv_1 \ring_25.inv_array[13]/sky_inverter/_0_  (.Y(\ring_25.inv_in[14] ),
    .A(\ring_25.inv_in[13] ));
 sg13g2_inv_1 \ring_25.inv_array[14]/sky_inverter/_0_  (.Y(\ring_25.inv_in[15] ),
    .A(\ring_25.inv_in[14] ));
 sg13g2_inv_1 \ring_25.inv_array[15]/sky_inverter/_0_  (.Y(\ring_25.inv_in[16] ),
    .A(\ring_25.inv_in[15] ));
 sg13g2_inv_1 \ring_25.inv_array[16]/sky_inverter/_0_  (.Y(\ring_25.inv_in[17] ),
    .A(\ring_25.inv_in[16] ));
 sg13g2_inv_1 \ring_25.inv_array[17]/sky_inverter/_0_  (.Y(\ring_25.inv_in[18] ),
    .A(\ring_25.inv_in[17] ));
 sg13g2_inv_1 \ring_25.inv_array[18]/sky_inverter/_0_  (.Y(\ring_25.inv_in[19] ),
    .A(\ring_25.inv_in[18] ));
 sg13g2_inv_1 \ring_25.inv_array[19]/sky_inverter/_0_  (.Y(\ring_25.inv_in[20] ),
    .A(\ring_25.inv_in[19] ));
 sg13g2_inv_1 \ring_25.inv_array[1]/sky_inverter/_0_  (.Y(\ring_25.inv_in[2] ),
    .A(\ring_25.inv_in[1] ));
 sg13g2_inv_1 \ring_25.inv_array[20]/sky_inverter/_0_  (.Y(\ring_25.inv_in[21] ),
    .A(\ring_25.inv_in[20] ));
 sg13g2_inv_1 \ring_25.inv_array[21]/sky_inverter/_0_  (.Y(\ring_25.inv_in[22] ),
    .A(\ring_25.inv_in[21] ));
 sg13g2_inv_1 \ring_25.inv_array[22]/sky_inverter/_0_  (.Y(\ring_25.inv_in[23] ),
    .A(\ring_25.inv_in[22] ));
 sg13g2_inv_1 \ring_25.inv_array[23]/sky_inverter/_0_  (.Y(\ring_25.inv_in[24] ),
    .A(\ring_25.inv_in[23] ));
 sg13g2_inv_1 \ring_25.inv_array[24]/sky_inverter/_0_  (.Y(\ring_25.inv_out[24] ),
    .A(\ring_25.inv_in[24] ));
 sg13g2_inv_1 \ring_25.inv_array[2]/sky_inverter/_0_  (.Y(\ring_25.inv_in[3] ),
    .A(\ring_25.inv_in[2] ));
 sg13g2_inv_1 \ring_25.inv_array[3]/sky_inverter/_0_  (.Y(\ring_25.inv_in[4] ),
    .A(\ring_25.inv_in[3] ));
 sg13g2_inv_1 \ring_25.inv_array[4]/sky_inverter/_0_  (.Y(\ring_25.inv_in[5] ),
    .A(\ring_25.inv_in[4] ));
 sg13g2_inv_1 \ring_25.inv_array[5]/sky_inverter/_0_  (.Y(\ring_25.inv_in[6] ),
    .A(\ring_25.inv_in[5] ));
 sg13g2_inv_1 \ring_25.inv_array[6]/sky_inverter/_0_  (.Y(\ring_25.inv_in[7] ),
    .A(\ring_25.inv_in[6] ));
 sg13g2_inv_1 \ring_25.inv_array[7]/sky_inverter/_0_  (.Y(\ring_25.inv_in[8] ),
    .A(\ring_25.inv_in[7] ));
 sg13g2_inv_1 \ring_25.inv_array[8]/sky_inverter/_0_  (.Y(\ring_25.inv_in[9] ),
    .A(\ring_25.inv_in[8] ));
 sg13g2_inv_1 \ring_25.inv_array[9]/sky_inverter/_0_  (.Y(\ring_25.inv_in[10] ),
    .A(\ring_25.inv_in[9] ));
 sg13g2_inv_1 \ring_251.inv_array[0]/sky_inverter/_0_  (.Y(\ring_251.inv_in[1] ),
    .A(\ring_251.inv_in[0] ));
 sg13g2_inv_1 \ring_251.inv_array[100]/sky_inverter/_0_  (.Y(\ring_251.inv_in[101] ),
    .A(\ring_251.inv_in[100] ));
 sg13g2_inv_1 \ring_251.inv_array[101]/sky_inverter/_0_  (.Y(\ring_251.inv_in[102] ),
    .A(\ring_251.inv_in[101] ));
 sg13g2_inv_1 \ring_251.inv_array[102]/sky_inverter/_0_  (.Y(\ring_251.inv_in[103] ),
    .A(\ring_251.inv_in[102] ));
 sg13g2_inv_1 \ring_251.inv_array[103]/sky_inverter/_0_  (.Y(\ring_251.inv_in[104] ),
    .A(\ring_251.inv_in[103] ));
 sg13g2_inv_1 \ring_251.inv_array[104]/sky_inverter/_0_  (.Y(\ring_251.inv_in[105] ),
    .A(\ring_251.inv_in[104] ));
 sg13g2_inv_1 \ring_251.inv_array[105]/sky_inverter/_0_  (.Y(\ring_251.inv_in[106] ),
    .A(\ring_251.inv_in[105] ));
 sg13g2_inv_1 \ring_251.inv_array[106]/sky_inverter/_0_  (.Y(\ring_251.inv_in[107] ),
    .A(\ring_251.inv_in[106] ));
 sg13g2_inv_1 \ring_251.inv_array[107]/sky_inverter/_0_  (.Y(\ring_251.inv_in[108] ),
    .A(\ring_251.inv_in[107] ));
 sg13g2_inv_1 \ring_251.inv_array[108]/sky_inverter/_0_  (.Y(\ring_251.inv_in[109] ),
    .A(\ring_251.inv_in[108] ));
 sg13g2_inv_1 \ring_251.inv_array[109]/sky_inverter/_0_  (.Y(\ring_251.inv_in[110] ),
    .A(\ring_251.inv_in[109] ));
 sg13g2_inv_1 \ring_251.inv_array[10]/sky_inverter/_0_  (.Y(\ring_251.inv_in[11] ),
    .A(\ring_251.inv_in[10] ));
 sg13g2_inv_1 \ring_251.inv_array[110]/sky_inverter/_0_  (.Y(\ring_251.inv_in[111] ),
    .A(\ring_251.inv_in[110] ));
 sg13g2_inv_1 \ring_251.inv_array[111]/sky_inverter/_0_  (.Y(\ring_251.inv_in[112] ),
    .A(\ring_251.inv_in[111] ));
 sg13g2_inv_1 \ring_251.inv_array[112]/sky_inverter/_0_  (.Y(\ring_251.inv_in[113] ),
    .A(\ring_251.inv_in[112] ));
 sg13g2_inv_1 \ring_251.inv_array[113]/sky_inverter/_0_  (.Y(\ring_251.inv_in[114] ),
    .A(\ring_251.inv_in[113] ));
 sg13g2_inv_1 \ring_251.inv_array[114]/sky_inverter/_0_  (.Y(\ring_251.inv_in[115] ),
    .A(\ring_251.inv_in[114] ));
 sg13g2_inv_1 \ring_251.inv_array[115]/sky_inverter/_0_  (.Y(\ring_251.inv_in[116] ),
    .A(\ring_251.inv_in[115] ));
 sg13g2_inv_1 \ring_251.inv_array[116]/sky_inverter/_0_  (.Y(\ring_251.inv_in[117] ),
    .A(\ring_251.inv_in[116] ));
 sg13g2_inv_1 \ring_251.inv_array[117]/sky_inverter/_0_  (.Y(\ring_251.inv_in[118] ),
    .A(\ring_251.inv_in[117] ));
 sg13g2_inv_1 \ring_251.inv_array[118]/sky_inverter/_0_  (.Y(\ring_251.inv_in[119] ),
    .A(\ring_251.inv_in[118] ));
 sg13g2_inv_1 \ring_251.inv_array[119]/sky_inverter/_0_  (.Y(\ring_251.inv_in[120] ),
    .A(\ring_251.inv_in[119] ));
 sg13g2_inv_1 \ring_251.inv_array[11]/sky_inverter/_0_  (.Y(\ring_251.inv_in[12] ),
    .A(\ring_251.inv_in[11] ));
 sg13g2_inv_1 \ring_251.inv_array[120]/sky_inverter/_0_  (.Y(\ring_251.inv_in[121] ),
    .A(\ring_251.inv_in[120] ));
 sg13g2_inv_1 \ring_251.inv_array[121]/sky_inverter/_0_  (.Y(\ring_251.inv_in[122] ),
    .A(\ring_251.inv_in[121] ));
 sg13g2_inv_1 \ring_251.inv_array[122]/sky_inverter/_0_  (.Y(\ring_251.inv_in[123] ),
    .A(\ring_251.inv_in[122] ));
 sg13g2_inv_1 \ring_251.inv_array[123]/sky_inverter/_0_  (.Y(\ring_251.inv_in[124] ),
    .A(\ring_251.inv_in[123] ));
 sg13g2_inv_1 \ring_251.inv_array[124]/sky_inverter/_0_  (.Y(\ring_251.inv_in[125] ),
    .A(\ring_251.inv_in[124] ));
 sg13g2_inv_1 \ring_251.inv_array[125]/sky_inverter/_0_  (.Y(\ring_251.inv_in[126] ),
    .A(\ring_251.inv_in[125] ));
 sg13g2_inv_1 \ring_251.inv_array[126]/sky_inverter/_0_  (.Y(\ring_251.inv_in[127] ),
    .A(\ring_251.inv_in[126] ));
 sg13g2_inv_1 \ring_251.inv_array[127]/sky_inverter/_0_  (.Y(\ring_251.inv_in[128] ),
    .A(\ring_251.inv_in[127] ));
 sg13g2_inv_1 \ring_251.inv_array[128]/sky_inverter/_0_  (.Y(\ring_251.inv_in[129] ),
    .A(\ring_251.inv_in[128] ));
 sg13g2_inv_1 \ring_251.inv_array[129]/sky_inverter/_0_  (.Y(\ring_251.inv_in[130] ),
    .A(\ring_251.inv_in[129] ));
 sg13g2_inv_1 \ring_251.inv_array[12]/sky_inverter/_0_  (.Y(\ring_251.inv_in[13] ),
    .A(\ring_251.inv_in[12] ));
 sg13g2_inv_1 \ring_251.inv_array[130]/sky_inverter/_0_  (.Y(\ring_251.inv_in[131] ),
    .A(\ring_251.inv_in[130] ));
 sg13g2_inv_1 \ring_251.inv_array[131]/sky_inverter/_0_  (.Y(\ring_251.inv_in[132] ),
    .A(\ring_251.inv_in[131] ));
 sg13g2_inv_1 \ring_251.inv_array[132]/sky_inverter/_0_  (.Y(\ring_251.inv_in[133] ),
    .A(\ring_251.inv_in[132] ));
 sg13g2_inv_1 \ring_251.inv_array[133]/sky_inverter/_0_  (.Y(\ring_251.inv_in[134] ),
    .A(\ring_251.inv_in[133] ));
 sg13g2_inv_1 \ring_251.inv_array[134]/sky_inverter/_0_  (.Y(\ring_251.inv_in[135] ),
    .A(\ring_251.inv_in[134] ));
 sg13g2_inv_1 \ring_251.inv_array[135]/sky_inverter/_0_  (.Y(\ring_251.inv_in[136] ),
    .A(\ring_251.inv_in[135] ));
 sg13g2_inv_1 \ring_251.inv_array[136]/sky_inverter/_0_  (.Y(\ring_251.inv_in[137] ),
    .A(\ring_251.inv_in[136] ));
 sg13g2_inv_1 \ring_251.inv_array[137]/sky_inverter/_0_  (.Y(\ring_251.inv_in[138] ),
    .A(\ring_251.inv_in[137] ));
 sg13g2_inv_1 \ring_251.inv_array[138]/sky_inverter/_0_  (.Y(\ring_251.inv_in[139] ),
    .A(\ring_251.inv_in[138] ));
 sg13g2_inv_1 \ring_251.inv_array[139]/sky_inverter/_0_  (.Y(\ring_251.inv_in[140] ),
    .A(\ring_251.inv_in[139] ));
 sg13g2_inv_1 \ring_251.inv_array[13]/sky_inverter/_0_  (.Y(\ring_251.inv_in[14] ),
    .A(\ring_251.inv_in[13] ));
 sg13g2_inv_1 \ring_251.inv_array[140]/sky_inverter/_0_  (.Y(\ring_251.inv_in[141] ),
    .A(\ring_251.inv_in[140] ));
 sg13g2_inv_1 \ring_251.inv_array[141]/sky_inverter/_0_  (.Y(\ring_251.inv_in[142] ),
    .A(\ring_251.inv_in[141] ));
 sg13g2_inv_1 \ring_251.inv_array[142]/sky_inverter/_0_  (.Y(\ring_251.inv_in[143] ),
    .A(\ring_251.inv_in[142] ));
 sg13g2_inv_1 \ring_251.inv_array[143]/sky_inverter/_0_  (.Y(\ring_251.inv_in[144] ),
    .A(\ring_251.inv_in[143] ));
 sg13g2_inv_1 \ring_251.inv_array[144]/sky_inverter/_0_  (.Y(\ring_251.inv_in[145] ),
    .A(\ring_251.inv_in[144] ));
 sg13g2_inv_1 \ring_251.inv_array[145]/sky_inverter/_0_  (.Y(\ring_251.inv_in[146] ),
    .A(\ring_251.inv_in[145] ));
 sg13g2_inv_1 \ring_251.inv_array[146]/sky_inverter/_0_  (.Y(\ring_251.inv_in[147] ),
    .A(\ring_251.inv_in[146] ));
 sg13g2_inv_1 \ring_251.inv_array[147]/sky_inverter/_0_  (.Y(\ring_251.inv_in[148] ),
    .A(\ring_251.inv_in[147] ));
 sg13g2_inv_1 \ring_251.inv_array[148]/sky_inverter/_0_  (.Y(\ring_251.inv_in[149] ),
    .A(\ring_251.inv_in[148] ));
 sg13g2_inv_1 \ring_251.inv_array[149]/sky_inverter/_0_  (.Y(\ring_251.inv_in[150] ),
    .A(\ring_251.inv_in[149] ));
 sg13g2_inv_1 \ring_251.inv_array[14]/sky_inverter/_0_  (.Y(\ring_251.inv_in[15] ),
    .A(\ring_251.inv_in[14] ));
 sg13g2_inv_1 \ring_251.inv_array[150]/sky_inverter/_0_  (.Y(\ring_251.inv_in[151] ),
    .A(\ring_251.inv_in[150] ));
 sg13g2_inv_1 \ring_251.inv_array[151]/sky_inverter/_0_  (.Y(\ring_251.inv_in[152] ),
    .A(\ring_251.inv_in[151] ));
 sg13g2_inv_1 \ring_251.inv_array[152]/sky_inverter/_0_  (.Y(\ring_251.inv_in[153] ),
    .A(\ring_251.inv_in[152] ));
 sg13g2_inv_1 \ring_251.inv_array[153]/sky_inverter/_0_  (.Y(\ring_251.inv_in[154] ),
    .A(\ring_251.inv_in[153] ));
 sg13g2_inv_1 \ring_251.inv_array[154]/sky_inverter/_0_  (.Y(\ring_251.inv_in[155] ),
    .A(\ring_251.inv_in[154] ));
 sg13g2_inv_1 \ring_251.inv_array[155]/sky_inverter/_0_  (.Y(\ring_251.inv_in[156] ),
    .A(\ring_251.inv_in[155] ));
 sg13g2_inv_1 \ring_251.inv_array[156]/sky_inverter/_0_  (.Y(\ring_251.inv_in[157] ),
    .A(\ring_251.inv_in[156] ));
 sg13g2_inv_1 \ring_251.inv_array[157]/sky_inverter/_0_  (.Y(\ring_251.inv_in[158] ),
    .A(\ring_251.inv_in[157] ));
 sg13g2_inv_1 \ring_251.inv_array[158]/sky_inverter/_0_  (.Y(\ring_251.inv_in[159] ),
    .A(\ring_251.inv_in[158] ));
 sg13g2_inv_1 \ring_251.inv_array[159]/sky_inverter/_0_  (.Y(\ring_251.inv_in[160] ),
    .A(\ring_251.inv_in[159] ));
 sg13g2_inv_1 \ring_251.inv_array[15]/sky_inverter/_0_  (.Y(\ring_251.inv_in[16] ),
    .A(\ring_251.inv_in[15] ));
 sg13g2_inv_1 \ring_251.inv_array[160]/sky_inverter/_0_  (.Y(\ring_251.inv_in[161] ),
    .A(\ring_251.inv_in[160] ));
 sg13g2_inv_1 \ring_251.inv_array[161]/sky_inverter/_0_  (.Y(\ring_251.inv_in[162] ),
    .A(\ring_251.inv_in[161] ));
 sg13g2_inv_1 \ring_251.inv_array[162]/sky_inverter/_0_  (.Y(\ring_251.inv_in[163] ),
    .A(\ring_251.inv_in[162] ));
 sg13g2_inv_1 \ring_251.inv_array[163]/sky_inverter/_0_  (.Y(\ring_251.inv_in[164] ),
    .A(\ring_251.inv_in[163] ));
 sg13g2_inv_1 \ring_251.inv_array[164]/sky_inverter/_0_  (.Y(\ring_251.inv_in[165] ),
    .A(\ring_251.inv_in[164] ));
 sg13g2_inv_1 \ring_251.inv_array[165]/sky_inverter/_0_  (.Y(\ring_251.inv_in[166] ),
    .A(\ring_251.inv_in[165] ));
 sg13g2_inv_1 \ring_251.inv_array[166]/sky_inverter/_0_  (.Y(\ring_251.inv_in[167] ),
    .A(\ring_251.inv_in[166] ));
 sg13g2_inv_1 \ring_251.inv_array[167]/sky_inverter/_0_  (.Y(\ring_251.inv_in[168] ),
    .A(\ring_251.inv_in[167] ));
 sg13g2_inv_1 \ring_251.inv_array[168]/sky_inverter/_0_  (.Y(\ring_251.inv_in[169] ),
    .A(\ring_251.inv_in[168] ));
 sg13g2_inv_1 \ring_251.inv_array[169]/sky_inverter/_0_  (.Y(\ring_251.inv_in[170] ),
    .A(\ring_251.inv_in[169] ));
 sg13g2_inv_1 \ring_251.inv_array[16]/sky_inverter/_0_  (.Y(\ring_251.inv_in[17] ),
    .A(\ring_251.inv_in[16] ));
 sg13g2_inv_1 \ring_251.inv_array[170]/sky_inverter/_0_  (.Y(\ring_251.inv_in[171] ),
    .A(\ring_251.inv_in[170] ));
 sg13g2_inv_1 \ring_251.inv_array[171]/sky_inverter/_0_  (.Y(\ring_251.inv_in[172] ),
    .A(\ring_251.inv_in[171] ));
 sg13g2_inv_1 \ring_251.inv_array[172]/sky_inverter/_0_  (.Y(\ring_251.inv_in[173] ),
    .A(\ring_251.inv_in[172] ));
 sg13g2_inv_1 \ring_251.inv_array[173]/sky_inverter/_0_  (.Y(\ring_251.inv_in[174] ),
    .A(\ring_251.inv_in[173] ));
 sg13g2_inv_1 \ring_251.inv_array[174]/sky_inverter/_0_  (.Y(\ring_251.inv_in[175] ),
    .A(\ring_251.inv_in[174] ));
 sg13g2_inv_1 \ring_251.inv_array[175]/sky_inverter/_0_  (.Y(\ring_251.inv_in[176] ),
    .A(\ring_251.inv_in[175] ));
 sg13g2_inv_1 \ring_251.inv_array[176]/sky_inverter/_0_  (.Y(\ring_251.inv_in[177] ),
    .A(\ring_251.inv_in[176] ));
 sg13g2_inv_1 \ring_251.inv_array[177]/sky_inverter/_0_  (.Y(\ring_251.inv_in[178] ),
    .A(\ring_251.inv_in[177] ));
 sg13g2_inv_1 \ring_251.inv_array[178]/sky_inverter/_0_  (.Y(\ring_251.inv_in[179] ),
    .A(\ring_251.inv_in[178] ));
 sg13g2_inv_1 \ring_251.inv_array[179]/sky_inverter/_0_  (.Y(\ring_251.inv_in[180] ),
    .A(\ring_251.inv_in[179] ));
 sg13g2_inv_1 \ring_251.inv_array[17]/sky_inverter/_0_  (.Y(\ring_251.inv_in[18] ),
    .A(\ring_251.inv_in[17] ));
 sg13g2_inv_1 \ring_251.inv_array[180]/sky_inverter/_0_  (.Y(\ring_251.inv_in[181] ),
    .A(\ring_251.inv_in[180] ));
 sg13g2_inv_1 \ring_251.inv_array[181]/sky_inverter/_0_  (.Y(\ring_251.inv_in[182] ),
    .A(\ring_251.inv_in[181] ));
 sg13g2_inv_1 \ring_251.inv_array[182]/sky_inverter/_0_  (.Y(\ring_251.inv_in[183] ),
    .A(\ring_251.inv_in[182] ));
 sg13g2_inv_1 \ring_251.inv_array[183]/sky_inverter/_0_  (.Y(\ring_251.inv_in[184] ),
    .A(\ring_251.inv_in[183] ));
 sg13g2_inv_1 \ring_251.inv_array[184]/sky_inverter/_0_  (.Y(\ring_251.inv_in[185] ),
    .A(\ring_251.inv_in[184] ));
 sg13g2_inv_1 \ring_251.inv_array[185]/sky_inverter/_0_  (.Y(\ring_251.inv_in[186] ),
    .A(\ring_251.inv_in[185] ));
 sg13g2_inv_1 \ring_251.inv_array[186]/sky_inverter/_0_  (.Y(\ring_251.inv_in[187] ),
    .A(\ring_251.inv_in[186] ));
 sg13g2_inv_1 \ring_251.inv_array[187]/sky_inverter/_0_  (.Y(\ring_251.inv_in[188] ),
    .A(\ring_251.inv_in[187] ));
 sg13g2_inv_1 \ring_251.inv_array[188]/sky_inverter/_0_  (.Y(\ring_251.inv_in[189] ),
    .A(\ring_251.inv_in[188] ));
 sg13g2_inv_1 \ring_251.inv_array[189]/sky_inverter/_0_  (.Y(\ring_251.inv_in[190] ),
    .A(\ring_251.inv_in[189] ));
 sg13g2_inv_1 \ring_251.inv_array[18]/sky_inverter/_0_  (.Y(\ring_251.inv_in[19] ),
    .A(\ring_251.inv_in[18] ));
 sg13g2_inv_1 \ring_251.inv_array[190]/sky_inverter/_0_  (.Y(\ring_251.inv_in[191] ),
    .A(\ring_251.inv_in[190] ));
 sg13g2_inv_1 \ring_251.inv_array[191]/sky_inverter/_0_  (.Y(\ring_251.inv_in[192] ),
    .A(\ring_251.inv_in[191] ));
 sg13g2_inv_1 \ring_251.inv_array[192]/sky_inverter/_0_  (.Y(\ring_251.inv_in[193] ),
    .A(\ring_251.inv_in[192] ));
 sg13g2_inv_1 \ring_251.inv_array[193]/sky_inverter/_0_  (.Y(\ring_251.inv_in[194] ),
    .A(\ring_251.inv_in[193] ));
 sg13g2_inv_1 \ring_251.inv_array[194]/sky_inverter/_0_  (.Y(\ring_251.inv_in[195] ),
    .A(\ring_251.inv_in[194] ));
 sg13g2_inv_1 \ring_251.inv_array[195]/sky_inverter/_0_  (.Y(\ring_251.inv_in[196] ),
    .A(\ring_251.inv_in[195] ));
 sg13g2_inv_1 \ring_251.inv_array[196]/sky_inverter/_0_  (.Y(\ring_251.inv_in[197] ),
    .A(\ring_251.inv_in[196] ));
 sg13g2_inv_1 \ring_251.inv_array[197]/sky_inverter/_0_  (.Y(\ring_251.inv_in[198] ),
    .A(\ring_251.inv_in[197] ));
 sg13g2_inv_1 \ring_251.inv_array[198]/sky_inverter/_0_  (.Y(\ring_251.inv_in[199] ),
    .A(\ring_251.inv_in[198] ));
 sg13g2_inv_1 \ring_251.inv_array[199]/sky_inverter/_0_  (.Y(\ring_251.inv_in[200] ),
    .A(\ring_251.inv_in[199] ));
 sg13g2_inv_1 \ring_251.inv_array[19]/sky_inverter/_0_  (.Y(\ring_251.inv_in[20] ),
    .A(\ring_251.inv_in[19] ));
 sg13g2_inv_1 \ring_251.inv_array[1]/sky_inverter/_0_  (.Y(\ring_251.inv_in[2] ),
    .A(\ring_251.inv_in[1] ));
 sg13g2_inv_1 \ring_251.inv_array[200]/sky_inverter/_0_  (.Y(\ring_251.inv_in[201] ),
    .A(\ring_251.inv_in[200] ));
 sg13g2_inv_1 \ring_251.inv_array[201]/sky_inverter/_0_  (.Y(\ring_251.inv_in[202] ),
    .A(\ring_251.inv_in[201] ));
 sg13g2_inv_1 \ring_251.inv_array[202]/sky_inverter/_0_  (.Y(\ring_251.inv_in[203] ),
    .A(\ring_251.inv_in[202] ));
 sg13g2_inv_1 \ring_251.inv_array[203]/sky_inverter/_0_  (.Y(\ring_251.inv_in[204] ),
    .A(\ring_251.inv_in[203] ));
 sg13g2_inv_1 \ring_251.inv_array[204]/sky_inverter/_0_  (.Y(\ring_251.inv_in[205] ),
    .A(\ring_251.inv_in[204] ));
 sg13g2_inv_1 \ring_251.inv_array[205]/sky_inverter/_0_  (.Y(\ring_251.inv_in[206] ),
    .A(\ring_251.inv_in[205] ));
 sg13g2_inv_1 \ring_251.inv_array[206]/sky_inverter/_0_  (.Y(\ring_251.inv_in[207] ),
    .A(\ring_251.inv_in[206] ));
 sg13g2_inv_1 \ring_251.inv_array[207]/sky_inverter/_0_  (.Y(\ring_251.inv_in[208] ),
    .A(\ring_251.inv_in[207] ));
 sg13g2_inv_1 \ring_251.inv_array[208]/sky_inverter/_0_  (.Y(\ring_251.inv_in[209] ),
    .A(\ring_251.inv_in[208] ));
 sg13g2_inv_1 \ring_251.inv_array[209]/sky_inverter/_0_  (.Y(\ring_251.inv_in[210] ),
    .A(\ring_251.inv_in[209] ));
 sg13g2_inv_1 \ring_251.inv_array[20]/sky_inverter/_0_  (.Y(\ring_251.inv_in[21] ),
    .A(\ring_251.inv_in[20] ));
 sg13g2_inv_1 \ring_251.inv_array[210]/sky_inverter/_0_  (.Y(\ring_251.inv_in[211] ),
    .A(\ring_251.inv_in[210] ));
 sg13g2_inv_1 \ring_251.inv_array[211]/sky_inverter/_0_  (.Y(\ring_251.inv_in[212] ),
    .A(\ring_251.inv_in[211] ));
 sg13g2_inv_1 \ring_251.inv_array[212]/sky_inverter/_0_  (.Y(\ring_251.inv_in[213] ),
    .A(\ring_251.inv_in[212] ));
 sg13g2_inv_1 \ring_251.inv_array[213]/sky_inverter/_0_  (.Y(\ring_251.inv_in[214] ),
    .A(\ring_251.inv_in[213] ));
 sg13g2_inv_1 \ring_251.inv_array[214]/sky_inverter/_0_  (.Y(\ring_251.inv_in[215] ),
    .A(\ring_251.inv_in[214] ));
 sg13g2_inv_1 \ring_251.inv_array[215]/sky_inverter/_0_  (.Y(\ring_251.inv_in[216] ),
    .A(\ring_251.inv_in[215] ));
 sg13g2_inv_1 \ring_251.inv_array[216]/sky_inverter/_0_  (.Y(\ring_251.inv_in[217] ),
    .A(\ring_251.inv_in[216] ));
 sg13g2_inv_1 \ring_251.inv_array[217]/sky_inverter/_0_  (.Y(\ring_251.inv_in[218] ),
    .A(\ring_251.inv_in[217] ));
 sg13g2_inv_1 \ring_251.inv_array[218]/sky_inverter/_0_  (.Y(\ring_251.inv_in[219] ),
    .A(\ring_251.inv_in[218] ));
 sg13g2_inv_1 \ring_251.inv_array[219]/sky_inverter/_0_  (.Y(\ring_251.inv_in[220] ),
    .A(\ring_251.inv_in[219] ));
 sg13g2_inv_1 \ring_251.inv_array[21]/sky_inverter/_0_  (.Y(\ring_251.inv_in[22] ),
    .A(\ring_251.inv_in[21] ));
 sg13g2_inv_1 \ring_251.inv_array[220]/sky_inverter/_0_  (.Y(\ring_251.inv_in[221] ),
    .A(\ring_251.inv_in[220] ));
 sg13g2_inv_1 \ring_251.inv_array[221]/sky_inverter/_0_  (.Y(\ring_251.inv_in[222] ),
    .A(\ring_251.inv_in[221] ));
 sg13g2_inv_1 \ring_251.inv_array[222]/sky_inverter/_0_  (.Y(\ring_251.inv_in[223] ),
    .A(\ring_251.inv_in[222] ));
 sg13g2_inv_1 \ring_251.inv_array[223]/sky_inverter/_0_  (.Y(\ring_251.inv_in[224] ),
    .A(\ring_251.inv_in[223] ));
 sg13g2_inv_1 \ring_251.inv_array[224]/sky_inverter/_0_  (.Y(\ring_251.inv_in[225] ),
    .A(\ring_251.inv_in[224] ));
 sg13g2_inv_1 \ring_251.inv_array[225]/sky_inverter/_0_  (.Y(\ring_251.inv_in[226] ),
    .A(\ring_251.inv_in[225] ));
 sg13g2_inv_1 \ring_251.inv_array[226]/sky_inverter/_0_  (.Y(\ring_251.inv_in[227] ),
    .A(\ring_251.inv_in[226] ));
 sg13g2_inv_1 \ring_251.inv_array[227]/sky_inverter/_0_  (.Y(\ring_251.inv_in[228] ),
    .A(\ring_251.inv_in[227] ));
 sg13g2_inv_1 \ring_251.inv_array[228]/sky_inverter/_0_  (.Y(\ring_251.inv_in[229] ),
    .A(\ring_251.inv_in[228] ));
 sg13g2_inv_1 \ring_251.inv_array[229]/sky_inverter/_0_  (.Y(\ring_251.inv_in[230] ),
    .A(\ring_251.inv_in[229] ));
 sg13g2_inv_1 \ring_251.inv_array[22]/sky_inverter/_0_  (.Y(\ring_251.inv_in[23] ),
    .A(\ring_251.inv_in[22] ));
 sg13g2_inv_1 \ring_251.inv_array[230]/sky_inverter/_0_  (.Y(\ring_251.inv_in[231] ),
    .A(\ring_251.inv_in[230] ));
 sg13g2_inv_1 \ring_251.inv_array[231]/sky_inverter/_0_  (.Y(\ring_251.inv_in[232] ),
    .A(\ring_251.inv_in[231] ));
 sg13g2_inv_1 \ring_251.inv_array[232]/sky_inverter/_0_  (.Y(\ring_251.inv_in[233] ),
    .A(\ring_251.inv_in[232] ));
 sg13g2_inv_1 \ring_251.inv_array[233]/sky_inverter/_0_  (.Y(\ring_251.inv_in[234] ),
    .A(\ring_251.inv_in[233] ));
 sg13g2_inv_1 \ring_251.inv_array[234]/sky_inverter/_0_  (.Y(\ring_251.inv_in[235] ),
    .A(\ring_251.inv_in[234] ));
 sg13g2_inv_1 \ring_251.inv_array[235]/sky_inverter/_0_  (.Y(\ring_251.inv_in[236] ),
    .A(\ring_251.inv_in[235] ));
 sg13g2_inv_1 \ring_251.inv_array[236]/sky_inverter/_0_  (.Y(\ring_251.inv_in[237] ),
    .A(\ring_251.inv_in[236] ));
 sg13g2_inv_1 \ring_251.inv_array[237]/sky_inverter/_0_  (.Y(\ring_251.inv_in[238] ),
    .A(\ring_251.inv_in[237] ));
 sg13g2_inv_1 \ring_251.inv_array[238]/sky_inverter/_0_  (.Y(\ring_251.inv_in[239] ),
    .A(\ring_251.inv_in[238] ));
 sg13g2_inv_1 \ring_251.inv_array[239]/sky_inverter/_0_  (.Y(\ring_251.inv_in[240] ),
    .A(\ring_251.inv_in[239] ));
 sg13g2_inv_1 \ring_251.inv_array[23]/sky_inverter/_0_  (.Y(\ring_251.inv_in[24] ),
    .A(\ring_251.inv_in[23] ));
 sg13g2_inv_1 \ring_251.inv_array[240]/sky_inverter/_0_  (.Y(\ring_251.inv_in[241] ),
    .A(\ring_251.inv_in[240] ));
 sg13g2_inv_1 \ring_251.inv_array[241]/sky_inverter/_0_  (.Y(\ring_251.inv_in[242] ),
    .A(\ring_251.inv_in[241] ));
 sg13g2_inv_1 \ring_251.inv_array[242]/sky_inverter/_0_  (.Y(\ring_251.inv_in[243] ),
    .A(\ring_251.inv_in[242] ));
 sg13g2_inv_1 \ring_251.inv_array[243]/sky_inverter/_0_  (.Y(\ring_251.inv_in[244] ),
    .A(\ring_251.inv_in[243] ));
 sg13g2_inv_1 \ring_251.inv_array[244]/sky_inverter/_0_  (.Y(\ring_251.inv_in[245] ),
    .A(\ring_251.inv_in[244] ));
 sg13g2_inv_1 \ring_251.inv_array[245]/sky_inverter/_0_  (.Y(\ring_251.inv_in[246] ),
    .A(\ring_251.inv_in[245] ));
 sg13g2_inv_1 \ring_251.inv_array[246]/sky_inverter/_0_  (.Y(\ring_251.inv_in[247] ),
    .A(\ring_251.inv_in[246] ));
 sg13g2_inv_1 \ring_251.inv_array[247]/sky_inverter/_0_  (.Y(\ring_251.inv_in[248] ),
    .A(\ring_251.inv_in[247] ));
 sg13g2_inv_1 \ring_251.inv_array[248]/sky_inverter/_0_  (.Y(\ring_251.inv_in[249] ),
    .A(\ring_251.inv_in[248] ));
 sg13g2_inv_1 \ring_251.inv_array[249]/sky_inverter/_0_  (.Y(\ring_251.inv_in[250] ),
    .A(\ring_251.inv_in[249] ));
 sg13g2_inv_1 \ring_251.inv_array[24]/sky_inverter/_0_  (.Y(\ring_251.inv_in[25] ),
    .A(\ring_251.inv_in[24] ));
 sg13g2_inv_1 \ring_251.inv_array[250]/sky_inverter/_0_  (.Y(\ring_251.inv_out[250] ),
    .A(\ring_251.inv_in[250] ));
 sg13g2_inv_1 \ring_251.inv_array[25]/sky_inverter/_0_  (.Y(\ring_251.inv_in[26] ),
    .A(\ring_251.inv_in[25] ));
 sg13g2_inv_1 \ring_251.inv_array[26]/sky_inverter/_0_  (.Y(\ring_251.inv_in[27] ),
    .A(\ring_251.inv_in[26] ));
 sg13g2_inv_1 \ring_251.inv_array[27]/sky_inverter/_0_  (.Y(\ring_251.inv_in[28] ),
    .A(\ring_251.inv_in[27] ));
 sg13g2_inv_1 \ring_251.inv_array[28]/sky_inverter/_0_  (.Y(\ring_251.inv_in[29] ),
    .A(\ring_251.inv_in[28] ));
 sg13g2_inv_1 \ring_251.inv_array[29]/sky_inverter/_0_  (.Y(\ring_251.inv_in[30] ),
    .A(\ring_251.inv_in[29] ));
 sg13g2_inv_1 \ring_251.inv_array[2]/sky_inverter/_0_  (.Y(\ring_251.inv_in[3] ),
    .A(\ring_251.inv_in[2] ));
 sg13g2_inv_1 \ring_251.inv_array[30]/sky_inverter/_0_  (.Y(\ring_251.inv_in[31] ),
    .A(\ring_251.inv_in[30] ));
 sg13g2_inv_1 \ring_251.inv_array[31]/sky_inverter/_0_  (.Y(\ring_251.inv_in[32] ),
    .A(\ring_251.inv_in[31] ));
 sg13g2_inv_1 \ring_251.inv_array[32]/sky_inverter/_0_  (.Y(\ring_251.inv_in[33] ),
    .A(\ring_251.inv_in[32] ));
 sg13g2_inv_1 \ring_251.inv_array[33]/sky_inverter/_0_  (.Y(\ring_251.inv_in[34] ),
    .A(\ring_251.inv_in[33] ));
 sg13g2_inv_1 \ring_251.inv_array[34]/sky_inverter/_0_  (.Y(\ring_251.inv_in[35] ),
    .A(\ring_251.inv_in[34] ));
 sg13g2_inv_1 \ring_251.inv_array[35]/sky_inverter/_0_  (.Y(\ring_251.inv_in[36] ),
    .A(\ring_251.inv_in[35] ));
 sg13g2_inv_1 \ring_251.inv_array[36]/sky_inverter/_0_  (.Y(\ring_251.inv_in[37] ),
    .A(\ring_251.inv_in[36] ));
 sg13g2_inv_1 \ring_251.inv_array[37]/sky_inverter/_0_  (.Y(\ring_251.inv_in[38] ),
    .A(\ring_251.inv_in[37] ));
 sg13g2_inv_1 \ring_251.inv_array[38]/sky_inverter/_0_  (.Y(\ring_251.inv_in[39] ),
    .A(\ring_251.inv_in[38] ));
 sg13g2_inv_1 \ring_251.inv_array[39]/sky_inverter/_0_  (.Y(\ring_251.inv_in[40] ),
    .A(\ring_251.inv_in[39] ));
 sg13g2_inv_1 \ring_251.inv_array[3]/sky_inverter/_0_  (.Y(\ring_251.inv_in[4] ),
    .A(\ring_251.inv_in[3] ));
 sg13g2_inv_1 \ring_251.inv_array[40]/sky_inverter/_0_  (.Y(\ring_251.inv_in[41] ),
    .A(\ring_251.inv_in[40] ));
 sg13g2_inv_1 \ring_251.inv_array[41]/sky_inverter/_0_  (.Y(\ring_251.inv_in[42] ),
    .A(\ring_251.inv_in[41] ));
 sg13g2_inv_1 \ring_251.inv_array[42]/sky_inverter/_0_  (.Y(\ring_251.inv_in[43] ),
    .A(\ring_251.inv_in[42] ));
 sg13g2_inv_1 \ring_251.inv_array[43]/sky_inverter/_0_  (.Y(\ring_251.inv_in[44] ),
    .A(\ring_251.inv_in[43] ));
 sg13g2_inv_1 \ring_251.inv_array[44]/sky_inverter/_0_  (.Y(\ring_251.inv_in[45] ),
    .A(\ring_251.inv_in[44] ));
 sg13g2_inv_1 \ring_251.inv_array[45]/sky_inverter/_0_  (.Y(\ring_251.inv_in[46] ),
    .A(\ring_251.inv_in[45] ));
 sg13g2_inv_1 \ring_251.inv_array[46]/sky_inverter/_0_  (.Y(\ring_251.inv_in[47] ),
    .A(\ring_251.inv_in[46] ));
 sg13g2_inv_1 \ring_251.inv_array[47]/sky_inverter/_0_  (.Y(\ring_251.inv_in[48] ),
    .A(\ring_251.inv_in[47] ));
 sg13g2_inv_1 \ring_251.inv_array[48]/sky_inverter/_0_  (.Y(\ring_251.inv_in[49] ),
    .A(\ring_251.inv_in[48] ));
 sg13g2_inv_1 \ring_251.inv_array[49]/sky_inverter/_0_  (.Y(\ring_251.inv_in[50] ),
    .A(\ring_251.inv_in[49] ));
 sg13g2_inv_1 \ring_251.inv_array[4]/sky_inverter/_0_  (.Y(\ring_251.inv_in[5] ),
    .A(\ring_251.inv_in[4] ));
 sg13g2_inv_1 \ring_251.inv_array[50]/sky_inverter/_0_  (.Y(\ring_251.inv_in[51] ),
    .A(\ring_251.inv_in[50] ));
 sg13g2_inv_1 \ring_251.inv_array[51]/sky_inverter/_0_  (.Y(\ring_251.inv_in[52] ),
    .A(\ring_251.inv_in[51] ));
 sg13g2_inv_1 \ring_251.inv_array[52]/sky_inverter/_0_  (.Y(\ring_251.inv_in[53] ),
    .A(\ring_251.inv_in[52] ));
 sg13g2_inv_1 \ring_251.inv_array[53]/sky_inverter/_0_  (.Y(\ring_251.inv_in[54] ),
    .A(\ring_251.inv_in[53] ));
 sg13g2_inv_1 \ring_251.inv_array[54]/sky_inverter/_0_  (.Y(\ring_251.inv_in[55] ),
    .A(\ring_251.inv_in[54] ));
 sg13g2_inv_1 \ring_251.inv_array[55]/sky_inverter/_0_  (.Y(\ring_251.inv_in[56] ),
    .A(\ring_251.inv_in[55] ));
 sg13g2_inv_1 \ring_251.inv_array[56]/sky_inverter/_0_  (.Y(\ring_251.inv_in[57] ),
    .A(\ring_251.inv_in[56] ));
 sg13g2_inv_1 \ring_251.inv_array[57]/sky_inverter/_0_  (.Y(\ring_251.inv_in[58] ),
    .A(\ring_251.inv_in[57] ));
 sg13g2_inv_1 \ring_251.inv_array[58]/sky_inverter/_0_  (.Y(\ring_251.inv_in[59] ),
    .A(\ring_251.inv_in[58] ));
 sg13g2_inv_1 \ring_251.inv_array[59]/sky_inverter/_0_  (.Y(\ring_251.inv_in[60] ),
    .A(\ring_251.inv_in[59] ));
 sg13g2_inv_1 \ring_251.inv_array[5]/sky_inverter/_0_  (.Y(\ring_251.inv_in[6] ),
    .A(\ring_251.inv_in[5] ));
 sg13g2_inv_1 \ring_251.inv_array[60]/sky_inverter/_0_  (.Y(\ring_251.inv_in[61] ),
    .A(\ring_251.inv_in[60] ));
 sg13g2_inv_1 \ring_251.inv_array[61]/sky_inverter/_0_  (.Y(\ring_251.inv_in[62] ),
    .A(\ring_251.inv_in[61] ));
 sg13g2_inv_1 \ring_251.inv_array[62]/sky_inverter/_0_  (.Y(\ring_251.inv_in[63] ),
    .A(\ring_251.inv_in[62] ));
 sg13g2_inv_1 \ring_251.inv_array[63]/sky_inverter/_0_  (.Y(\ring_251.inv_in[64] ),
    .A(\ring_251.inv_in[63] ));
 sg13g2_inv_1 \ring_251.inv_array[64]/sky_inverter/_0_  (.Y(\ring_251.inv_in[65] ),
    .A(\ring_251.inv_in[64] ));
 sg13g2_inv_1 \ring_251.inv_array[65]/sky_inverter/_0_  (.Y(\ring_251.inv_in[66] ),
    .A(\ring_251.inv_in[65] ));
 sg13g2_inv_1 \ring_251.inv_array[66]/sky_inverter/_0_  (.Y(\ring_251.inv_in[67] ),
    .A(\ring_251.inv_in[66] ));
 sg13g2_inv_1 \ring_251.inv_array[67]/sky_inverter/_0_  (.Y(\ring_251.inv_in[68] ),
    .A(\ring_251.inv_in[67] ));
 sg13g2_inv_1 \ring_251.inv_array[68]/sky_inverter/_0_  (.Y(\ring_251.inv_in[69] ),
    .A(\ring_251.inv_in[68] ));
 sg13g2_inv_1 \ring_251.inv_array[69]/sky_inverter/_0_  (.Y(\ring_251.inv_in[70] ),
    .A(\ring_251.inv_in[69] ));
 sg13g2_inv_1 \ring_251.inv_array[6]/sky_inverter/_0_  (.Y(\ring_251.inv_in[7] ),
    .A(\ring_251.inv_in[6] ));
 sg13g2_inv_1 \ring_251.inv_array[70]/sky_inverter/_0_  (.Y(\ring_251.inv_in[71] ),
    .A(\ring_251.inv_in[70] ));
 sg13g2_inv_1 \ring_251.inv_array[71]/sky_inverter/_0_  (.Y(\ring_251.inv_in[72] ),
    .A(\ring_251.inv_in[71] ));
 sg13g2_inv_1 \ring_251.inv_array[72]/sky_inverter/_0_  (.Y(\ring_251.inv_in[73] ),
    .A(\ring_251.inv_in[72] ));
 sg13g2_inv_1 \ring_251.inv_array[73]/sky_inverter/_0_  (.Y(\ring_251.inv_in[74] ),
    .A(\ring_251.inv_in[73] ));
 sg13g2_inv_1 \ring_251.inv_array[74]/sky_inverter/_0_  (.Y(\ring_251.inv_in[75] ),
    .A(\ring_251.inv_in[74] ));
 sg13g2_inv_1 \ring_251.inv_array[75]/sky_inverter/_0_  (.Y(\ring_251.inv_in[76] ),
    .A(\ring_251.inv_in[75] ));
 sg13g2_inv_1 \ring_251.inv_array[76]/sky_inverter/_0_  (.Y(\ring_251.inv_in[77] ),
    .A(\ring_251.inv_in[76] ));
 sg13g2_inv_1 \ring_251.inv_array[77]/sky_inverter/_0_  (.Y(\ring_251.inv_in[78] ),
    .A(\ring_251.inv_in[77] ));
 sg13g2_inv_1 \ring_251.inv_array[78]/sky_inverter/_0_  (.Y(\ring_251.inv_in[79] ),
    .A(\ring_251.inv_in[78] ));
 sg13g2_inv_1 \ring_251.inv_array[79]/sky_inverter/_0_  (.Y(\ring_251.inv_in[80] ),
    .A(\ring_251.inv_in[79] ));
 sg13g2_inv_1 \ring_251.inv_array[7]/sky_inverter/_0_  (.Y(\ring_251.inv_in[8] ),
    .A(\ring_251.inv_in[7] ));
 sg13g2_inv_1 \ring_251.inv_array[80]/sky_inverter/_0_  (.Y(\ring_251.inv_in[81] ),
    .A(\ring_251.inv_in[80] ));
 sg13g2_inv_1 \ring_251.inv_array[81]/sky_inverter/_0_  (.Y(\ring_251.inv_in[82] ),
    .A(\ring_251.inv_in[81] ));
 sg13g2_inv_1 \ring_251.inv_array[82]/sky_inverter/_0_  (.Y(\ring_251.inv_in[83] ),
    .A(\ring_251.inv_in[82] ));
 sg13g2_inv_1 \ring_251.inv_array[83]/sky_inverter/_0_  (.Y(\ring_251.inv_in[84] ),
    .A(\ring_251.inv_in[83] ));
 sg13g2_inv_1 \ring_251.inv_array[84]/sky_inverter/_0_  (.Y(\ring_251.inv_in[85] ),
    .A(\ring_251.inv_in[84] ));
 sg13g2_inv_1 \ring_251.inv_array[85]/sky_inverter/_0_  (.Y(\ring_251.inv_in[86] ),
    .A(\ring_251.inv_in[85] ));
 sg13g2_inv_1 \ring_251.inv_array[86]/sky_inverter/_0_  (.Y(\ring_251.inv_in[87] ),
    .A(\ring_251.inv_in[86] ));
 sg13g2_inv_1 \ring_251.inv_array[87]/sky_inverter/_0_  (.Y(\ring_251.inv_in[88] ),
    .A(\ring_251.inv_in[87] ));
 sg13g2_inv_1 \ring_251.inv_array[88]/sky_inverter/_0_  (.Y(\ring_251.inv_in[89] ),
    .A(\ring_251.inv_in[88] ));
 sg13g2_inv_1 \ring_251.inv_array[89]/sky_inverter/_0_  (.Y(\ring_251.inv_in[90] ),
    .A(\ring_251.inv_in[89] ));
 sg13g2_inv_1 \ring_251.inv_array[8]/sky_inverter/_0_  (.Y(\ring_251.inv_in[9] ),
    .A(\ring_251.inv_in[8] ));
 sg13g2_inv_1 \ring_251.inv_array[90]/sky_inverter/_0_  (.Y(\ring_251.inv_in[91] ),
    .A(\ring_251.inv_in[90] ));
 sg13g2_inv_1 \ring_251.inv_array[91]/sky_inverter/_0_  (.Y(\ring_251.inv_in[92] ),
    .A(\ring_251.inv_in[91] ));
 sg13g2_inv_1 \ring_251.inv_array[92]/sky_inverter/_0_  (.Y(\ring_251.inv_in[93] ),
    .A(\ring_251.inv_in[92] ));
 sg13g2_inv_1 \ring_251.inv_array[93]/sky_inverter/_0_  (.Y(\ring_251.inv_in[94] ),
    .A(\ring_251.inv_in[93] ));
 sg13g2_inv_1 \ring_251.inv_array[94]/sky_inverter/_0_  (.Y(\ring_251.inv_in[95] ),
    .A(\ring_251.inv_in[94] ));
 sg13g2_inv_1 \ring_251.inv_array[95]/sky_inverter/_0_  (.Y(\ring_251.inv_in[96] ),
    .A(\ring_251.inv_in[95] ));
 sg13g2_inv_1 \ring_251.inv_array[96]/sky_inverter/_0_  (.Y(\ring_251.inv_in[97] ),
    .A(\ring_251.inv_in[96] ));
 sg13g2_inv_1 \ring_251.inv_array[97]/sky_inverter/_0_  (.Y(\ring_251.inv_in[98] ),
    .A(\ring_251.inv_in[97] ));
 sg13g2_inv_1 \ring_251.inv_array[98]/sky_inverter/_0_  (.Y(\ring_251.inv_in[99] ),
    .A(\ring_251.inv_in[98] ));
 sg13g2_inv_1 \ring_251.inv_array[99]/sky_inverter/_0_  (.Y(\ring_251.inv_in[100] ),
    .A(\ring_251.inv_in[99] ));
 sg13g2_inv_1 \ring_251.inv_array[9]/sky_inverter/_0_  (.Y(\ring_251.inv_in[10] ),
    .A(\ring_251.inv_in[9] ));
 sg13g2_inv_1 \ring_501.inv_array[0]/sky_inverter/_0_  (.Y(\ring_501.inv_in[1] ),
    .A(c0clock));
 sg13g2_inv_1 \ring_501.inv_array[100]/sky_inverter/_0_  (.Y(\ring_501.inv_in[101] ),
    .A(\ring_501.inv_in[100] ));
 sg13g2_inv_1 \ring_501.inv_array[101]/sky_inverter/_0_  (.Y(\ring_501.inv_in[102] ),
    .A(\ring_501.inv_in[101] ));
 sg13g2_inv_1 \ring_501.inv_array[102]/sky_inverter/_0_  (.Y(\ring_501.inv_in[103] ),
    .A(\ring_501.inv_in[102] ));
 sg13g2_inv_1 \ring_501.inv_array[103]/sky_inverter/_0_  (.Y(\ring_501.inv_in[104] ),
    .A(\ring_501.inv_in[103] ));
 sg13g2_inv_1 \ring_501.inv_array[104]/sky_inverter/_0_  (.Y(\ring_501.inv_in[105] ),
    .A(\ring_501.inv_in[104] ));
 sg13g2_inv_1 \ring_501.inv_array[105]/sky_inverter/_0_  (.Y(\ring_501.inv_in[106] ),
    .A(\ring_501.inv_in[105] ));
 sg13g2_inv_1 \ring_501.inv_array[106]/sky_inverter/_0_  (.Y(\ring_501.inv_in[107] ),
    .A(\ring_501.inv_in[106] ));
 sg13g2_inv_1 \ring_501.inv_array[107]/sky_inverter/_0_  (.Y(\ring_501.inv_in[108] ),
    .A(\ring_501.inv_in[107] ));
 sg13g2_inv_1 \ring_501.inv_array[108]/sky_inverter/_0_  (.Y(\ring_501.inv_in[109] ),
    .A(\ring_501.inv_in[108] ));
 sg13g2_inv_1 \ring_501.inv_array[109]/sky_inverter/_0_  (.Y(\ring_501.inv_in[110] ),
    .A(\ring_501.inv_in[109] ));
 sg13g2_inv_1 \ring_501.inv_array[10]/sky_inverter/_0_  (.Y(\ring_501.inv_in[11] ),
    .A(\ring_501.inv_in[10] ));
 sg13g2_inv_1 \ring_501.inv_array[110]/sky_inverter/_0_  (.Y(\ring_501.inv_in[111] ),
    .A(\ring_501.inv_in[110] ));
 sg13g2_inv_1 \ring_501.inv_array[111]/sky_inverter/_0_  (.Y(\ring_501.inv_in[112] ),
    .A(\ring_501.inv_in[111] ));
 sg13g2_inv_1 \ring_501.inv_array[112]/sky_inverter/_0_  (.Y(\ring_501.inv_in[113] ),
    .A(\ring_501.inv_in[112] ));
 sg13g2_inv_1 \ring_501.inv_array[113]/sky_inverter/_0_  (.Y(\ring_501.inv_in[114] ),
    .A(\ring_501.inv_in[113] ));
 sg13g2_inv_1 \ring_501.inv_array[114]/sky_inverter/_0_  (.Y(\ring_501.inv_in[115] ),
    .A(\ring_501.inv_in[114] ));
 sg13g2_inv_1 \ring_501.inv_array[115]/sky_inverter/_0_  (.Y(\ring_501.inv_in[116] ),
    .A(\ring_501.inv_in[115] ));
 sg13g2_inv_1 \ring_501.inv_array[116]/sky_inverter/_0_  (.Y(\ring_501.inv_in[117] ),
    .A(\ring_501.inv_in[116] ));
 sg13g2_inv_1 \ring_501.inv_array[117]/sky_inverter/_0_  (.Y(\ring_501.inv_in[118] ),
    .A(\ring_501.inv_in[117] ));
 sg13g2_inv_1 \ring_501.inv_array[118]/sky_inverter/_0_  (.Y(\ring_501.inv_in[119] ),
    .A(\ring_501.inv_in[118] ));
 sg13g2_inv_1 \ring_501.inv_array[119]/sky_inverter/_0_  (.Y(\ring_501.inv_in[120] ),
    .A(\ring_501.inv_in[119] ));
 sg13g2_inv_1 \ring_501.inv_array[11]/sky_inverter/_0_  (.Y(\ring_501.inv_in[12] ),
    .A(\ring_501.inv_in[11] ));
 sg13g2_inv_1 \ring_501.inv_array[120]/sky_inverter/_0_  (.Y(\ring_501.inv_in[121] ),
    .A(\ring_501.inv_in[120] ));
 sg13g2_inv_1 \ring_501.inv_array[121]/sky_inverter/_0_  (.Y(\ring_501.inv_in[122] ),
    .A(\ring_501.inv_in[121] ));
 sg13g2_inv_1 \ring_501.inv_array[122]/sky_inverter/_0_  (.Y(\ring_501.inv_in[123] ),
    .A(\ring_501.inv_in[122] ));
 sg13g2_inv_1 \ring_501.inv_array[123]/sky_inverter/_0_  (.Y(\ring_501.inv_in[124] ),
    .A(\ring_501.inv_in[123] ));
 sg13g2_inv_1 \ring_501.inv_array[124]/sky_inverter/_0_  (.Y(\ring_501.inv_in[125] ),
    .A(\ring_501.inv_in[124] ));
 sg13g2_inv_1 \ring_501.inv_array[125]/sky_inverter/_0_  (.Y(\ring_501.inv_in[126] ),
    .A(\ring_501.inv_in[125] ));
 sg13g2_inv_1 \ring_501.inv_array[126]/sky_inverter/_0_  (.Y(\ring_501.inv_in[127] ),
    .A(\ring_501.inv_in[126] ));
 sg13g2_inv_1 \ring_501.inv_array[127]/sky_inverter/_0_  (.Y(\ring_501.inv_in[128] ),
    .A(\ring_501.inv_in[127] ));
 sg13g2_inv_1 \ring_501.inv_array[128]/sky_inverter/_0_  (.Y(\ring_501.inv_in[129] ),
    .A(\ring_501.inv_in[128] ));
 sg13g2_inv_1 \ring_501.inv_array[129]/sky_inverter/_0_  (.Y(\ring_501.inv_in[130] ),
    .A(\ring_501.inv_in[129] ));
 sg13g2_inv_1 \ring_501.inv_array[12]/sky_inverter/_0_  (.Y(\ring_501.inv_in[13] ),
    .A(\ring_501.inv_in[12] ));
 sg13g2_inv_1 \ring_501.inv_array[130]/sky_inverter/_0_  (.Y(\ring_501.inv_in[131] ),
    .A(\ring_501.inv_in[130] ));
 sg13g2_inv_1 \ring_501.inv_array[131]/sky_inverter/_0_  (.Y(\ring_501.inv_in[132] ),
    .A(\ring_501.inv_in[131] ));
 sg13g2_inv_1 \ring_501.inv_array[132]/sky_inverter/_0_  (.Y(\ring_501.inv_in[133] ),
    .A(\ring_501.inv_in[132] ));
 sg13g2_inv_1 \ring_501.inv_array[133]/sky_inverter/_0_  (.Y(\ring_501.inv_in[134] ),
    .A(\ring_501.inv_in[133] ));
 sg13g2_inv_1 \ring_501.inv_array[134]/sky_inverter/_0_  (.Y(\ring_501.inv_in[135] ),
    .A(\ring_501.inv_in[134] ));
 sg13g2_inv_1 \ring_501.inv_array[135]/sky_inverter/_0_  (.Y(\ring_501.inv_in[136] ),
    .A(\ring_501.inv_in[135] ));
 sg13g2_inv_1 \ring_501.inv_array[136]/sky_inverter/_0_  (.Y(\ring_501.inv_in[137] ),
    .A(\ring_501.inv_in[136] ));
 sg13g2_inv_1 \ring_501.inv_array[137]/sky_inverter/_0_  (.Y(\ring_501.inv_in[138] ),
    .A(\ring_501.inv_in[137] ));
 sg13g2_inv_1 \ring_501.inv_array[138]/sky_inverter/_0_  (.Y(\ring_501.inv_in[139] ),
    .A(\ring_501.inv_in[138] ));
 sg13g2_inv_1 \ring_501.inv_array[139]/sky_inverter/_0_  (.Y(\ring_501.inv_in[140] ),
    .A(\ring_501.inv_in[139] ));
 sg13g2_inv_1 \ring_501.inv_array[13]/sky_inverter/_0_  (.Y(\ring_501.inv_in[14] ),
    .A(\ring_501.inv_in[13] ));
 sg13g2_inv_1 \ring_501.inv_array[140]/sky_inverter/_0_  (.Y(\ring_501.inv_in[141] ),
    .A(\ring_501.inv_in[140] ));
 sg13g2_inv_1 \ring_501.inv_array[141]/sky_inverter/_0_  (.Y(\ring_501.inv_in[142] ),
    .A(\ring_501.inv_in[141] ));
 sg13g2_inv_1 \ring_501.inv_array[142]/sky_inverter/_0_  (.Y(\ring_501.inv_in[143] ),
    .A(\ring_501.inv_in[142] ));
 sg13g2_inv_1 \ring_501.inv_array[143]/sky_inverter/_0_  (.Y(\ring_501.inv_in[144] ),
    .A(\ring_501.inv_in[143] ));
 sg13g2_inv_1 \ring_501.inv_array[144]/sky_inverter/_0_  (.Y(\ring_501.inv_in[145] ),
    .A(\ring_501.inv_in[144] ));
 sg13g2_inv_1 \ring_501.inv_array[145]/sky_inverter/_0_  (.Y(\ring_501.inv_in[146] ),
    .A(\ring_501.inv_in[145] ));
 sg13g2_inv_1 \ring_501.inv_array[146]/sky_inverter/_0_  (.Y(\ring_501.inv_in[147] ),
    .A(\ring_501.inv_in[146] ));
 sg13g2_inv_1 \ring_501.inv_array[147]/sky_inverter/_0_  (.Y(\ring_501.inv_in[148] ),
    .A(\ring_501.inv_in[147] ));
 sg13g2_inv_1 \ring_501.inv_array[148]/sky_inverter/_0_  (.Y(\ring_501.inv_in[149] ),
    .A(\ring_501.inv_in[148] ));
 sg13g2_inv_1 \ring_501.inv_array[149]/sky_inverter/_0_  (.Y(\ring_501.inv_in[150] ),
    .A(\ring_501.inv_in[149] ));
 sg13g2_inv_1 \ring_501.inv_array[14]/sky_inverter/_0_  (.Y(\ring_501.inv_in[15] ),
    .A(\ring_501.inv_in[14] ));
 sg13g2_inv_1 \ring_501.inv_array[150]/sky_inverter/_0_  (.Y(\ring_501.inv_in[151] ),
    .A(\ring_501.inv_in[150] ));
 sg13g2_inv_1 \ring_501.inv_array[151]/sky_inverter/_0_  (.Y(\ring_501.inv_in[152] ),
    .A(\ring_501.inv_in[151] ));
 sg13g2_inv_1 \ring_501.inv_array[152]/sky_inverter/_0_  (.Y(\ring_501.inv_in[153] ),
    .A(\ring_501.inv_in[152] ));
 sg13g2_inv_1 \ring_501.inv_array[153]/sky_inverter/_0_  (.Y(\ring_501.inv_in[154] ),
    .A(\ring_501.inv_in[153] ));
 sg13g2_inv_1 \ring_501.inv_array[154]/sky_inverter/_0_  (.Y(\ring_501.inv_in[155] ),
    .A(\ring_501.inv_in[154] ));
 sg13g2_inv_1 \ring_501.inv_array[155]/sky_inverter/_0_  (.Y(\ring_501.inv_in[156] ),
    .A(\ring_501.inv_in[155] ));
 sg13g2_inv_1 \ring_501.inv_array[156]/sky_inverter/_0_  (.Y(\ring_501.inv_in[157] ),
    .A(\ring_501.inv_in[156] ));
 sg13g2_inv_1 \ring_501.inv_array[157]/sky_inverter/_0_  (.Y(\ring_501.inv_in[158] ),
    .A(\ring_501.inv_in[157] ));
 sg13g2_inv_1 \ring_501.inv_array[158]/sky_inverter/_0_  (.Y(\ring_501.inv_in[159] ),
    .A(\ring_501.inv_in[158] ));
 sg13g2_inv_1 \ring_501.inv_array[159]/sky_inverter/_0_  (.Y(\ring_501.inv_in[160] ),
    .A(\ring_501.inv_in[159] ));
 sg13g2_inv_1 \ring_501.inv_array[15]/sky_inverter/_0_  (.Y(\ring_501.inv_in[16] ),
    .A(\ring_501.inv_in[15] ));
 sg13g2_inv_1 \ring_501.inv_array[160]/sky_inverter/_0_  (.Y(\ring_501.inv_in[161] ),
    .A(\ring_501.inv_in[160] ));
 sg13g2_inv_1 \ring_501.inv_array[161]/sky_inverter/_0_  (.Y(\ring_501.inv_in[162] ),
    .A(\ring_501.inv_in[161] ));
 sg13g2_inv_1 \ring_501.inv_array[162]/sky_inverter/_0_  (.Y(\ring_501.inv_in[163] ),
    .A(\ring_501.inv_in[162] ));
 sg13g2_inv_1 \ring_501.inv_array[163]/sky_inverter/_0_  (.Y(\ring_501.inv_in[164] ),
    .A(\ring_501.inv_in[163] ));
 sg13g2_inv_1 \ring_501.inv_array[164]/sky_inverter/_0_  (.Y(\ring_501.inv_in[165] ),
    .A(\ring_501.inv_in[164] ));
 sg13g2_inv_1 \ring_501.inv_array[165]/sky_inverter/_0_  (.Y(\ring_501.inv_in[166] ),
    .A(\ring_501.inv_in[165] ));
 sg13g2_inv_1 \ring_501.inv_array[166]/sky_inverter/_0_  (.Y(\ring_501.inv_in[167] ),
    .A(\ring_501.inv_in[166] ));
 sg13g2_inv_1 \ring_501.inv_array[167]/sky_inverter/_0_  (.Y(\ring_501.inv_in[168] ),
    .A(\ring_501.inv_in[167] ));
 sg13g2_inv_1 \ring_501.inv_array[168]/sky_inverter/_0_  (.Y(\ring_501.inv_in[169] ),
    .A(\ring_501.inv_in[168] ));
 sg13g2_inv_1 \ring_501.inv_array[169]/sky_inverter/_0_  (.Y(\ring_501.inv_in[170] ),
    .A(\ring_501.inv_in[169] ));
 sg13g2_inv_1 \ring_501.inv_array[16]/sky_inverter/_0_  (.Y(\ring_501.inv_in[17] ),
    .A(\ring_501.inv_in[16] ));
 sg13g2_inv_1 \ring_501.inv_array[170]/sky_inverter/_0_  (.Y(\ring_501.inv_in[171] ),
    .A(\ring_501.inv_in[170] ));
 sg13g2_inv_1 \ring_501.inv_array[171]/sky_inverter/_0_  (.Y(\ring_501.inv_in[172] ),
    .A(\ring_501.inv_in[171] ));
 sg13g2_inv_1 \ring_501.inv_array[172]/sky_inverter/_0_  (.Y(\ring_501.inv_in[173] ),
    .A(\ring_501.inv_in[172] ));
 sg13g2_inv_1 \ring_501.inv_array[173]/sky_inverter/_0_  (.Y(\ring_501.inv_in[174] ),
    .A(\ring_501.inv_in[173] ));
 sg13g2_inv_1 \ring_501.inv_array[174]/sky_inverter/_0_  (.Y(\ring_501.inv_in[175] ),
    .A(\ring_501.inv_in[174] ));
 sg13g2_inv_1 \ring_501.inv_array[175]/sky_inverter/_0_  (.Y(\ring_501.inv_in[176] ),
    .A(\ring_501.inv_in[175] ));
 sg13g2_inv_1 \ring_501.inv_array[176]/sky_inverter/_0_  (.Y(\ring_501.inv_in[177] ),
    .A(\ring_501.inv_in[176] ));
 sg13g2_inv_1 \ring_501.inv_array[177]/sky_inverter/_0_  (.Y(\ring_501.inv_in[178] ),
    .A(\ring_501.inv_in[177] ));
 sg13g2_inv_1 \ring_501.inv_array[178]/sky_inverter/_0_  (.Y(\ring_501.inv_in[179] ),
    .A(\ring_501.inv_in[178] ));
 sg13g2_inv_1 \ring_501.inv_array[179]/sky_inverter/_0_  (.Y(\ring_501.inv_in[180] ),
    .A(\ring_501.inv_in[179] ));
 sg13g2_inv_1 \ring_501.inv_array[17]/sky_inverter/_0_  (.Y(\ring_501.inv_in[18] ),
    .A(\ring_501.inv_in[17] ));
 sg13g2_inv_1 \ring_501.inv_array[180]/sky_inverter/_0_  (.Y(\ring_501.inv_in[181] ),
    .A(\ring_501.inv_in[180] ));
 sg13g2_inv_1 \ring_501.inv_array[181]/sky_inverter/_0_  (.Y(\ring_501.inv_in[182] ),
    .A(\ring_501.inv_in[181] ));
 sg13g2_inv_1 \ring_501.inv_array[182]/sky_inverter/_0_  (.Y(\ring_501.inv_in[183] ),
    .A(\ring_501.inv_in[182] ));
 sg13g2_inv_1 \ring_501.inv_array[183]/sky_inverter/_0_  (.Y(\ring_501.inv_in[184] ),
    .A(\ring_501.inv_in[183] ));
 sg13g2_inv_1 \ring_501.inv_array[184]/sky_inverter/_0_  (.Y(\ring_501.inv_in[185] ),
    .A(\ring_501.inv_in[184] ));
 sg13g2_inv_1 \ring_501.inv_array[185]/sky_inverter/_0_  (.Y(\ring_501.inv_in[186] ),
    .A(\ring_501.inv_in[185] ));
 sg13g2_inv_1 \ring_501.inv_array[186]/sky_inverter/_0_  (.Y(\ring_501.inv_in[187] ),
    .A(\ring_501.inv_in[186] ));
 sg13g2_inv_1 \ring_501.inv_array[187]/sky_inverter/_0_  (.Y(\ring_501.inv_in[188] ),
    .A(\ring_501.inv_in[187] ));
 sg13g2_inv_1 \ring_501.inv_array[188]/sky_inverter/_0_  (.Y(\ring_501.inv_in[189] ),
    .A(\ring_501.inv_in[188] ));
 sg13g2_inv_1 \ring_501.inv_array[189]/sky_inverter/_0_  (.Y(\ring_501.inv_in[190] ),
    .A(\ring_501.inv_in[189] ));
 sg13g2_inv_1 \ring_501.inv_array[18]/sky_inverter/_0_  (.Y(\ring_501.inv_in[19] ),
    .A(\ring_501.inv_in[18] ));
 sg13g2_inv_1 \ring_501.inv_array[190]/sky_inverter/_0_  (.Y(\ring_501.inv_in[191] ),
    .A(\ring_501.inv_in[190] ));
 sg13g2_inv_1 \ring_501.inv_array[191]/sky_inverter/_0_  (.Y(\ring_501.inv_in[192] ),
    .A(\ring_501.inv_in[191] ));
 sg13g2_inv_1 \ring_501.inv_array[192]/sky_inverter/_0_  (.Y(\ring_501.inv_in[193] ),
    .A(\ring_501.inv_in[192] ));
 sg13g2_inv_1 \ring_501.inv_array[193]/sky_inverter/_0_  (.Y(\ring_501.inv_in[194] ),
    .A(\ring_501.inv_in[193] ));
 sg13g2_inv_1 \ring_501.inv_array[194]/sky_inverter/_0_  (.Y(\ring_501.inv_in[195] ),
    .A(\ring_501.inv_in[194] ));
 sg13g2_inv_1 \ring_501.inv_array[195]/sky_inverter/_0_  (.Y(\ring_501.inv_in[196] ),
    .A(\ring_501.inv_in[195] ));
 sg13g2_inv_1 \ring_501.inv_array[196]/sky_inverter/_0_  (.Y(\ring_501.inv_in[197] ),
    .A(\ring_501.inv_in[196] ));
 sg13g2_inv_1 \ring_501.inv_array[197]/sky_inverter/_0_  (.Y(\ring_501.inv_in[198] ),
    .A(\ring_501.inv_in[197] ));
 sg13g2_inv_1 \ring_501.inv_array[198]/sky_inverter/_0_  (.Y(\ring_501.inv_in[199] ),
    .A(\ring_501.inv_in[198] ));
 sg13g2_inv_1 \ring_501.inv_array[199]/sky_inverter/_0_  (.Y(\ring_501.inv_in[200] ),
    .A(\ring_501.inv_in[199] ));
 sg13g2_inv_1 \ring_501.inv_array[19]/sky_inverter/_0_  (.Y(\ring_501.inv_in[20] ),
    .A(\ring_501.inv_in[19] ));
 sg13g2_inv_1 \ring_501.inv_array[1]/sky_inverter/_0_  (.Y(\ring_501.inv_in[2] ),
    .A(\ring_501.inv_in[1] ));
 sg13g2_inv_1 \ring_501.inv_array[200]/sky_inverter/_0_  (.Y(\ring_501.inv_in[201] ),
    .A(\ring_501.inv_in[200] ));
 sg13g2_inv_1 \ring_501.inv_array[201]/sky_inverter/_0_  (.Y(\ring_501.inv_in[202] ),
    .A(\ring_501.inv_in[201] ));
 sg13g2_inv_1 \ring_501.inv_array[202]/sky_inverter/_0_  (.Y(\ring_501.inv_in[203] ),
    .A(\ring_501.inv_in[202] ));
 sg13g2_inv_1 \ring_501.inv_array[203]/sky_inverter/_0_  (.Y(\ring_501.inv_in[204] ),
    .A(\ring_501.inv_in[203] ));
 sg13g2_inv_1 \ring_501.inv_array[204]/sky_inverter/_0_  (.Y(\ring_501.inv_in[205] ),
    .A(\ring_501.inv_in[204] ));
 sg13g2_inv_1 \ring_501.inv_array[205]/sky_inverter/_0_  (.Y(\ring_501.inv_in[206] ),
    .A(\ring_501.inv_in[205] ));
 sg13g2_inv_1 \ring_501.inv_array[206]/sky_inverter/_0_  (.Y(\ring_501.inv_in[207] ),
    .A(\ring_501.inv_in[206] ));
 sg13g2_inv_1 \ring_501.inv_array[207]/sky_inverter/_0_  (.Y(\ring_501.inv_in[208] ),
    .A(\ring_501.inv_in[207] ));
 sg13g2_inv_1 \ring_501.inv_array[208]/sky_inverter/_0_  (.Y(\ring_501.inv_in[209] ),
    .A(\ring_501.inv_in[208] ));
 sg13g2_inv_1 \ring_501.inv_array[209]/sky_inverter/_0_  (.Y(\ring_501.inv_in[210] ),
    .A(\ring_501.inv_in[209] ));
 sg13g2_inv_1 \ring_501.inv_array[20]/sky_inverter/_0_  (.Y(\ring_501.inv_in[21] ),
    .A(\ring_501.inv_in[20] ));
 sg13g2_inv_1 \ring_501.inv_array[210]/sky_inverter/_0_  (.Y(\ring_501.inv_in[211] ),
    .A(\ring_501.inv_in[210] ));
 sg13g2_inv_1 \ring_501.inv_array[211]/sky_inverter/_0_  (.Y(\ring_501.inv_in[212] ),
    .A(\ring_501.inv_in[211] ));
 sg13g2_inv_1 \ring_501.inv_array[212]/sky_inverter/_0_  (.Y(\ring_501.inv_in[213] ),
    .A(\ring_501.inv_in[212] ));
 sg13g2_inv_1 \ring_501.inv_array[213]/sky_inverter/_0_  (.Y(\ring_501.inv_in[214] ),
    .A(\ring_501.inv_in[213] ));
 sg13g2_inv_1 \ring_501.inv_array[214]/sky_inverter/_0_  (.Y(\ring_501.inv_in[215] ),
    .A(\ring_501.inv_in[214] ));
 sg13g2_inv_1 \ring_501.inv_array[215]/sky_inverter/_0_  (.Y(\ring_501.inv_in[216] ),
    .A(\ring_501.inv_in[215] ));
 sg13g2_inv_1 \ring_501.inv_array[216]/sky_inverter/_0_  (.Y(\ring_501.inv_in[217] ),
    .A(\ring_501.inv_in[216] ));
 sg13g2_inv_1 \ring_501.inv_array[217]/sky_inverter/_0_  (.Y(\ring_501.inv_in[218] ),
    .A(\ring_501.inv_in[217] ));
 sg13g2_inv_1 \ring_501.inv_array[218]/sky_inverter/_0_  (.Y(\ring_501.inv_in[219] ),
    .A(\ring_501.inv_in[218] ));
 sg13g2_inv_1 \ring_501.inv_array[219]/sky_inverter/_0_  (.Y(\ring_501.inv_in[220] ),
    .A(\ring_501.inv_in[219] ));
 sg13g2_inv_1 \ring_501.inv_array[21]/sky_inverter/_0_  (.Y(\ring_501.inv_in[22] ),
    .A(\ring_501.inv_in[21] ));
 sg13g2_inv_1 \ring_501.inv_array[220]/sky_inverter/_0_  (.Y(\ring_501.inv_in[221] ),
    .A(\ring_501.inv_in[220] ));
 sg13g2_inv_1 \ring_501.inv_array[221]/sky_inverter/_0_  (.Y(\ring_501.inv_in[222] ),
    .A(\ring_501.inv_in[221] ));
 sg13g2_inv_1 \ring_501.inv_array[222]/sky_inverter/_0_  (.Y(\ring_501.inv_in[223] ),
    .A(\ring_501.inv_in[222] ));
 sg13g2_inv_1 \ring_501.inv_array[223]/sky_inverter/_0_  (.Y(\ring_501.inv_in[224] ),
    .A(\ring_501.inv_in[223] ));
 sg13g2_inv_1 \ring_501.inv_array[224]/sky_inverter/_0_  (.Y(\ring_501.inv_in[225] ),
    .A(\ring_501.inv_in[224] ));
 sg13g2_inv_1 \ring_501.inv_array[225]/sky_inverter/_0_  (.Y(\ring_501.inv_in[226] ),
    .A(\ring_501.inv_in[225] ));
 sg13g2_inv_1 \ring_501.inv_array[226]/sky_inverter/_0_  (.Y(\ring_501.inv_in[227] ),
    .A(\ring_501.inv_in[226] ));
 sg13g2_inv_1 \ring_501.inv_array[227]/sky_inverter/_0_  (.Y(\ring_501.inv_in[228] ),
    .A(\ring_501.inv_in[227] ));
 sg13g2_inv_1 \ring_501.inv_array[228]/sky_inverter/_0_  (.Y(\ring_501.inv_in[229] ),
    .A(\ring_501.inv_in[228] ));
 sg13g2_inv_1 \ring_501.inv_array[229]/sky_inverter/_0_  (.Y(\ring_501.inv_in[230] ),
    .A(\ring_501.inv_in[229] ));
 sg13g2_inv_1 \ring_501.inv_array[22]/sky_inverter/_0_  (.Y(\ring_501.inv_in[23] ),
    .A(\ring_501.inv_in[22] ));
 sg13g2_inv_1 \ring_501.inv_array[230]/sky_inverter/_0_  (.Y(\ring_501.inv_in[231] ),
    .A(\ring_501.inv_in[230] ));
 sg13g2_inv_1 \ring_501.inv_array[231]/sky_inverter/_0_  (.Y(\ring_501.inv_in[232] ),
    .A(\ring_501.inv_in[231] ));
 sg13g2_inv_1 \ring_501.inv_array[232]/sky_inverter/_0_  (.Y(\ring_501.inv_in[233] ),
    .A(\ring_501.inv_in[232] ));
 sg13g2_inv_1 \ring_501.inv_array[233]/sky_inverter/_0_  (.Y(\ring_501.inv_in[234] ),
    .A(\ring_501.inv_in[233] ));
 sg13g2_inv_1 \ring_501.inv_array[234]/sky_inverter/_0_  (.Y(\ring_501.inv_in[235] ),
    .A(\ring_501.inv_in[234] ));
 sg13g2_inv_1 \ring_501.inv_array[235]/sky_inverter/_0_  (.Y(\ring_501.inv_in[236] ),
    .A(\ring_501.inv_in[235] ));
 sg13g2_inv_1 \ring_501.inv_array[236]/sky_inverter/_0_  (.Y(\ring_501.inv_in[237] ),
    .A(\ring_501.inv_in[236] ));
 sg13g2_inv_1 \ring_501.inv_array[237]/sky_inverter/_0_  (.Y(\ring_501.inv_in[238] ),
    .A(\ring_501.inv_in[237] ));
 sg13g2_inv_1 \ring_501.inv_array[238]/sky_inverter/_0_  (.Y(\ring_501.inv_in[239] ),
    .A(\ring_501.inv_in[238] ));
 sg13g2_inv_1 \ring_501.inv_array[239]/sky_inverter/_0_  (.Y(\ring_501.inv_in[240] ),
    .A(\ring_501.inv_in[239] ));
 sg13g2_inv_1 \ring_501.inv_array[23]/sky_inverter/_0_  (.Y(\ring_501.inv_in[24] ),
    .A(\ring_501.inv_in[23] ));
 sg13g2_inv_1 \ring_501.inv_array[240]/sky_inverter/_0_  (.Y(\ring_501.inv_in[241] ),
    .A(\ring_501.inv_in[240] ));
 sg13g2_inv_1 \ring_501.inv_array[241]/sky_inverter/_0_  (.Y(\ring_501.inv_in[242] ),
    .A(\ring_501.inv_in[241] ));
 sg13g2_inv_1 \ring_501.inv_array[242]/sky_inverter/_0_  (.Y(\ring_501.inv_in[243] ),
    .A(\ring_501.inv_in[242] ));
 sg13g2_inv_1 \ring_501.inv_array[243]/sky_inverter/_0_  (.Y(\ring_501.inv_in[244] ),
    .A(\ring_501.inv_in[243] ));
 sg13g2_inv_1 \ring_501.inv_array[244]/sky_inverter/_0_  (.Y(\ring_501.inv_in[245] ),
    .A(\ring_501.inv_in[244] ));
 sg13g2_inv_1 \ring_501.inv_array[245]/sky_inverter/_0_  (.Y(\ring_501.inv_in[246] ),
    .A(\ring_501.inv_in[245] ));
 sg13g2_inv_1 \ring_501.inv_array[246]/sky_inverter/_0_  (.Y(\ring_501.inv_in[247] ),
    .A(\ring_501.inv_in[246] ));
 sg13g2_inv_1 \ring_501.inv_array[247]/sky_inverter/_0_  (.Y(\ring_501.inv_in[248] ),
    .A(\ring_501.inv_in[247] ));
 sg13g2_inv_1 \ring_501.inv_array[248]/sky_inverter/_0_  (.Y(\ring_501.inv_in[249] ),
    .A(\ring_501.inv_in[248] ));
 sg13g2_inv_1 \ring_501.inv_array[249]/sky_inverter/_0_  (.Y(\ring_501.inv_in[250] ),
    .A(\ring_501.inv_in[249] ));
 sg13g2_inv_1 \ring_501.inv_array[24]/sky_inverter/_0_  (.Y(\ring_501.inv_in[25] ),
    .A(\ring_501.inv_in[24] ));
 sg13g2_inv_1 \ring_501.inv_array[250]/sky_inverter/_0_  (.Y(\ring_501.inv_in[251] ),
    .A(\ring_501.inv_in[250] ));
 sg13g2_inv_1 \ring_501.inv_array[251]/sky_inverter/_0_  (.Y(\ring_501.inv_in[252] ),
    .A(\ring_501.inv_in[251] ));
 sg13g2_inv_1 \ring_501.inv_array[252]/sky_inverter/_0_  (.Y(\ring_501.inv_in[253] ),
    .A(\ring_501.inv_in[252] ));
 sg13g2_inv_1 \ring_501.inv_array[253]/sky_inverter/_0_  (.Y(\ring_501.inv_in[254] ),
    .A(\ring_501.inv_in[253] ));
 sg13g2_inv_1 \ring_501.inv_array[254]/sky_inverter/_0_  (.Y(\ring_501.inv_in[255] ),
    .A(\ring_501.inv_in[254] ));
 sg13g2_inv_1 \ring_501.inv_array[255]/sky_inverter/_0_  (.Y(\ring_501.inv_in[256] ),
    .A(\ring_501.inv_in[255] ));
 sg13g2_inv_1 \ring_501.inv_array[256]/sky_inverter/_0_  (.Y(\ring_501.inv_in[257] ),
    .A(\ring_501.inv_in[256] ));
 sg13g2_inv_1 \ring_501.inv_array[257]/sky_inverter/_0_  (.Y(\ring_501.inv_in[258] ),
    .A(\ring_501.inv_in[257] ));
 sg13g2_inv_1 \ring_501.inv_array[258]/sky_inverter/_0_  (.Y(\ring_501.inv_in[259] ),
    .A(\ring_501.inv_in[258] ));
 sg13g2_inv_1 \ring_501.inv_array[259]/sky_inverter/_0_  (.Y(\ring_501.inv_in[260] ),
    .A(\ring_501.inv_in[259] ));
 sg13g2_inv_1 \ring_501.inv_array[25]/sky_inverter/_0_  (.Y(\ring_501.inv_in[26] ),
    .A(\ring_501.inv_in[25] ));
 sg13g2_inv_1 \ring_501.inv_array[260]/sky_inverter/_0_  (.Y(\ring_501.inv_in[261] ),
    .A(\ring_501.inv_in[260] ));
 sg13g2_inv_1 \ring_501.inv_array[261]/sky_inverter/_0_  (.Y(\ring_501.inv_in[262] ),
    .A(\ring_501.inv_in[261] ));
 sg13g2_inv_1 \ring_501.inv_array[262]/sky_inverter/_0_  (.Y(\ring_501.inv_in[263] ),
    .A(\ring_501.inv_in[262] ));
 sg13g2_inv_1 \ring_501.inv_array[263]/sky_inverter/_0_  (.Y(\ring_501.inv_in[264] ),
    .A(\ring_501.inv_in[263] ));
 sg13g2_inv_1 \ring_501.inv_array[264]/sky_inverter/_0_  (.Y(\ring_501.inv_in[265] ),
    .A(\ring_501.inv_in[264] ));
 sg13g2_inv_1 \ring_501.inv_array[265]/sky_inverter/_0_  (.Y(\ring_501.inv_in[266] ),
    .A(\ring_501.inv_in[265] ));
 sg13g2_inv_1 \ring_501.inv_array[266]/sky_inverter/_0_  (.Y(\ring_501.inv_in[267] ),
    .A(\ring_501.inv_in[266] ));
 sg13g2_inv_1 \ring_501.inv_array[267]/sky_inverter/_0_  (.Y(\ring_501.inv_in[268] ),
    .A(\ring_501.inv_in[267] ));
 sg13g2_inv_1 \ring_501.inv_array[268]/sky_inverter/_0_  (.Y(\ring_501.inv_in[269] ),
    .A(\ring_501.inv_in[268] ));
 sg13g2_inv_1 \ring_501.inv_array[269]/sky_inverter/_0_  (.Y(\ring_501.inv_in[270] ),
    .A(\ring_501.inv_in[269] ));
 sg13g2_inv_1 \ring_501.inv_array[26]/sky_inverter/_0_  (.Y(\ring_501.inv_in[27] ),
    .A(\ring_501.inv_in[26] ));
 sg13g2_inv_1 \ring_501.inv_array[270]/sky_inverter/_0_  (.Y(\ring_501.inv_in[271] ),
    .A(\ring_501.inv_in[270] ));
 sg13g2_inv_1 \ring_501.inv_array[271]/sky_inverter/_0_  (.Y(\ring_501.inv_in[272] ),
    .A(\ring_501.inv_in[271] ));
 sg13g2_inv_1 \ring_501.inv_array[272]/sky_inverter/_0_  (.Y(\ring_501.inv_in[273] ),
    .A(\ring_501.inv_in[272] ));
 sg13g2_inv_1 \ring_501.inv_array[273]/sky_inverter/_0_  (.Y(\ring_501.inv_in[274] ),
    .A(\ring_501.inv_in[273] ));
 sg13g2_inv_1 \ring_501.inv_array[274]/sky_inverter/_0_  (.Y(\ring_501.inv_in[275] ),
    .A(\ring_501.inv_in[274] ));
 sg13g2_inv_1 \ring_501.inv_array[275]/sky_inverter/_0_  (.Y(\ring_501.inv_in[276] ),
    .A(\ring_501.inv_in[275] ));
 sg13g2_inv_1 \ring_501.inv_array[276]/sky_inverter/_0_  (.Y(\ring_501.inv_in[277] ),
    .A(\ring_501.inv_in[276] ));
 sg13g2_inv_1 \ring_501.inv_array[277]/sky_inverter/_0_  (.Y(\ring_501.inv_in[278] ),
    .A(\ring_501.inv_in[277] ));
 sg13g2_inv_1 \ring_501.inv_array[278]/sky_inverter/_0_  (.Y(\ring_501.inv_in[279] ),
    .A(\ring_501.inv_in[278] ));
 sg13g2_inv_1 \ring_501.inv_array[279]/sky_inverter/_0_  (.Y(\ring_501.inv_in[280] ),
    .A(\ring_501.inv_in[279] ));
 sg13g2_inv_1 \ring_501.inv_array[27]/sky_inverter/_0_  (.Y(\ring_501.inv_in[28] ),
    .A(\ring_501.inv_in[27] ));
 sg13g2_inv_1 \ring_501.inv_array[280]/sky_inverter/_0_  (.Y(\ring_501.inv_in[281] ),
    .A(\ring_501.inv_in[280] ));
 sg13g2_inv_1 \ring_501.inv_array[281]/sky_inverter/_0_  (.Y(\ring_501.inv_in[282] ),
    .A(\ring_501.inv_in[281] ));
 sg13g2_inv_1 \ring_501.inv_array[282]/sky_inverter/_0_  (.Y(\ring_501.inv_in[283] ),
    .A(\ring_501.inv_in[282] ));
 sg13g2_inv_1 \ring_501.inv_array[283]/sky_inverter/_0_  (.Y(\ring_501.inv_in[284] ),
    .A(\ring_501.inv_in[283] ));
 sg13g2_inv_1 \ring_501.inv_array[284]/sky_inverter/_0_  (.Y(\ring_501.inv_in[285] ),
    .A(\ring_501.inv_in[284] ));
 sg13g2_inv_1 \ring_501.inv_array[285]/sky_inverter/_0_  (.Y(\ring_501.inv_in[286] ),
    .A(\ring_501.inv_in[285] ));
 sg13g2_inv_1 \ring_501.inv_array[286]/sky_inverter/_0_  (.Y(\ring_501.inv_in[287] ),
    .A(\ring_501.inv_in[286] ));
 sg13g2_inv_1 \ring_501.inv_array[287]/sky_inverter/_0_  (.Y(\ring_501.inv_in[288] ),
    .A(\ring_501.inv_in[287] ));
 sg13g2_inv_1 \ring_501.inv_array[288]/sky_inverter/_0_  (.Y(\ring_501.inv_in[289] ),
    .A(\ring_501.inv_in[288] ));
 sg13g2_inv_1 \ring_501.inv_array[289]/sky_inverter/_0_  (.Y(\ring_501.inv_in[290] ),
    .A(\ring_501.inv_in[289] ));
 sg13g2_inv_1 \ring_501.inv_array[28]/sky_inverter/_0_  (.Y(\ring_501.inv_in[29] ),
    .A(\ring_501.inv_in[28] ));
 sg13g2_inv_1 \ring_501.inv_array[290]/sky_inverter/_0_  (.Y(\ring_501.inv_in[291] ),
    .A(\ring_501.inv_in[290] ));
 sg13g2_inv_1 \ring_501.inv_array[291]/sky_inverter/_0_  (.Y(\ring_501.inv_in[292] ),
    .A(\ring_501.inv_in[291] ));
 sg13g2_inv_1 \ring_501.inv_array[292]/sky_inverter/_0_  (.Y(\ring_501.inv_in[293] ),
    .A(\ring_501.inv_in[292] ));
 sg13g2_inv_1 \ring_501.inv_array[293]/sky_inverter/_0_  (.Y(\ring_501.inv_in[294] ),
    .A(\ring_501.inv_in[293] ));
 sg13g2_inv_1 \ring_501.inv_array[294]/sky_inverter/_0_  (.Y(\ring_501.inv_in[295] ),
    .A(\ring_501.inv_in[294] ));
 sg13g2_inv_1 \ring_501.inv_array[295]/sky_inverter/_0_  (.Y(\ring_501.inv_in[296] ),
    .A(\ring_501.inv_in[295] ));
 sg13g2_inv_1 \ring_501.inv_array[296]/sky_inverter/_0_  (.Y(\ring_501.inv_in[297] ),
    .A(\ring_501.inv_in[296] ));
 sg13g2_inv_1 \ring_501.inv_array[297]/sky_inverter/_0_  (.Y(\ring_501.inv_in[298] ),
    .A(\ring_501.inv_in[297] ));
 sg13g2_inv_1 \ring_501.inv_array[298]/sky_inverter/_0_  (.Y(\ring_501.inv_in[299] ),
    .A(\ring_501.inv_in[298] ));
 sg13g2_inv_1 \ring_501.inv_array[299]/sky_inverter/_0_  (.Y(\ring_501.inv_in[300] ),
    .A(\ring_501.inv_in[299] ));
 sg13g2_inv_1 \ring_501.inv_array[29]/sky_inverter/_0_  (.Y(\ring_501.inv_in[30] ),
    .A(\ring_501.inv_in[29] ));
 sg13g2_inv_1 \ring_501.inv_array[2]/sky_inverter/_0_  (.Y(\ring_501.inv_in[3] ),
    .A(\ring_501.inv_in[2] ));
 sg13g2_inv_1 \ring_501.inv_array[300]/sky_inverter/_0_  (.Y(\ring_501.inv_in[301] ),
    .A(\ring_501.inv_in[300] ));
 sg13g2_inv_1 \ring_501.inv_array[301]/sky_inverter/_0_  (.Y(\ring_501.inv_in[302] ),
    .A(\ring_501.inv_in[301] ));
 sg13g2_inv_1 \ring_501.inv_array[302]/sky_inverter/_0_  (.Y(\ring_501.inv_in[303] ),
    .A(\ring_501.inv_in[302] ));
 sg13g2_inv_1 \ring_501.inv_array[303]/sky_inverter/_0_  (.Y(\ring_501.inv_in[304] ),
    .A(\ring_501.inv_in[303] ));
 sg13g2_inv_1 \ring_501.inv_array[304]/sky_inverter/_0_  (.Y(\ring_501.inv_in[305] ),
    .A(\ring_501.inv_in[304] ));
 sg13g2_inv_1 \ring_501.inv_array[305]/sky_inverter/_0_  (.Y(\ring_501.inv_in[306] ),
    .A(\ring_501.inv_in[305] ));
 sg13g2_inv_1 \ring_501.inv_array[306]/sky_inverter/_0_  (.Y(\ring_501.inv_in[307] ),
    .A(\ring_501.inv_in[306] ));
 sg13g2_inv_1 \ring_501.inv_array[307]/sky_inverter/_0_  (.Y(\ring_501.inv_in[308] ),
    .A(\ring_501.inv_in[307] ));
 sg13g2_inv_1 \ring_501.inv_array[308]/sky_inverter/_0_  (.Y(\ring_501.inv_in[309] ),
    .A(\ring_501.inv_in[308] ));
 sg13g2_inv_1 \ring_501.inv_array[309]/sky_inverter/_0_  (.Y(\ring_501.inv_in[310] ),
    .A(\ring_501.inv_in[309] ));
 sg13g2_inv_1 \ring_501.inv_array[30]/sky_inverter/_0_  (.Y(\ring_501.inv_in[31] ),
    .A(\ring_501.inv_in[30] ));
 sg13g2_inv_1 \ring_501.inv_array[310]/sky_inverter/_0_  (.Y(\ring_501.inv_in[311] ),
    .A(\ring_501.inv_in[310] ));
 sg13g2_inv_1 \ring_501.inv_array[311]/sky_inverter/_0_  (.Y(\ring_501.inv_in[312] ),
    .A(\ring_501.inv_in[311] ));
 sg13g2_inv_1 \ring_501.inv_array[312]/sky_inverter/_0_  (.Y(\ring_501.inv_in[313] ),
    .A(\ring_501.inv_in[312] ));
 sg13g2_inv_1 \ring_501.inv_array[313]/sky_inverter/_0_  (.Y(\ring_501.inv_in[314] ),
    .A(\ring_501.inv_in[313] ));
 sg13g2_inv_1 \ring_501.inv_array[314]/sky_inverter/_0_  (.Y(\ring_501.inv_in[315] ),
    .A(\ring_501.inv_in[314] ));
 sg13g2_inv_1 \ring_501.inv_array[315]/sky_inverter/_0_  (.Y(\ring_501.inv_in[316] ),
    .A(\ring_501.inv_in[315] ));
 sg13g2_inv_1 \ring_501.inv_array[316]/sky_inverter/_0_  (.Y(\ring_501.inv_in[317] ),
    .A(\ring_501.inv_in[316] ));
 sg13g2_inv_1 \ring_501.inv_array[317]/sky_inverter/_0_  (.Y(\ring_501.inv_in[318] ),
    .A(\ring_501.inv_in[317] ));
 sg13g2_inv_1 \ring_501.inv_array[318]/sky_inverter/_0_  (.Y(\ring_501.inv_in[319] ),
    .A(\ring_501.inv_in[318] ));
 sg13g2_inv_1 \ring_501.inv_array[319]/sky_inverter/_0_  (.Y(\ring_501.inv_in[320] ),
    .A(\ring_501.inv_in[319] ));
 sg13g2_inv_1 \ring_501.inv_array[31]/sky_inverter/_0_  (.Y(\ring_501.inv_in[32] ),
    .A(\ring_501.inv_in[31] ));
 sg13g2_inv_1 \ring_501.inv_array[320]/sky_inverter/_0_  (.Y(\ring_501.inv_in[321] ),
    .A(\ring_501.inv_in[320] ));
 sg13g2_inv_1 \ring_501.inv_array[321]/sky_inverter/_0_  (.Y(\ring_501.inv_in[322] ),
    .A(\ring_501.inv_in[321] ));
 sg13g2_inv_1 \ring_501.inv_array[322]/sky_inverter/_0_  (.Y(\ring_501.inv_in[323] ),
    .A(\ring_501.inv_in[322] ));
 sg13g2_inv_1 \ring_501.inv_array[323]/sky_inverter/_0_  (.Y(\ring_501.inv_in[324] ),
    .A(\ring_501.inv_in[323] ));
 sg13g2_inv_1 \ring_501.inv_array[324]/sky_inverter/_0_  (.Y(\ring_501.inv_in[325] ),
    .A(\ring_501.inv_in[324] ));
 sg13g2_inv_1 \ring_501.inv_array[325]/sky_inverter/_0_  (.Y(\ring_501.inv_in[326] ),
    .A(\ring_501.inv_in[325] ));
 sg13g2_inv_1 \ring_501.inv_array[326]/sky_inverter/_0_  (.Y(\ring_501.inv_in[327] ),
    .A(\ring_501.inv_in[326] ));
 sg13g2_inv_1 \ring_501.inv_array[327]/sky_inverter/_0_  (.Y(\ring_501.inv_in[328] ),
    .A(\ring_501.inv_in[327] ));
 sg13g2_inv_1 \ring_501.inv_array[328]/sky_inverter/_0_  (.Y(\ring_501.inv_in[329] ),
    .A(\ring_501.inv_in[328] ));
 sg13g2_inv_1 \ring_501.inv_array[329]/sky_inverter/_0_  (.Y(\ring_501.inv_in[330] ),
    .A(\ring_501.inv_in[329] ));
 sg13g2_inv_1 \ring_501.inv_array[32]/sky_inverter/_0_  (.Y(\ring_501.inv_in[33] ),
    .A(\ring_501.inv_in[32] ));
 sg13g2_inv_1 \ring_501.inv_array[330]/sky_inverter/_0_  (.Y(\ring_501.inv_in[331] ),
    .A(\ring_501.inv_in[330] ));
 sg13g2_inv_1 \ring_501.inv_array[331]/sky_inverter/_0_  (.Y(\ring_501.inv_in[332] ),
    .A(\ring_501.inv_in[331] ));
 sg13g2_inv_1 \ring_501.inv_array[332]/sky_inverter/_0_  (.Y(\ring_501.inv_in[333] ),
    .A(\ring_501.inv_in[332] ));
 sg13g2_inv_1 \ring_501.inv_array[333]/sky_inverter/_0_  (.Y(\ring_501.inv_in[334] ),
    .A(\ring_501.inv_in[333] ));
 sg13g2_inv_1 \ring_501.inv_array[334]/sky_inverter/_0_  (.Y(\ring_501.inv_in[335] ),
    .A(\ring_501.inv_in[334] ));
 sg13g2_inv_1 \ring_501.inv_array[335]/sky_inverter/_0_  (.Y(\ring_501.inv_in[336] ),
    .A(\ring_501.inv_in[335] ));
 sg13g2_inv_1 \ring_501.inv_array[336]/sky_inverter/_0_  (.Y(\ring_501.inv_in[337] ),
    .A(\ring_501.inv_in[336] ));
 sg13g2_inv_1 \ring_501.inv_array[337]/sky_inverter/_0_  (.Y(\ring_501.inv_in[338] ),
    .A(\ring_501.inv_in[337] ));
 sg13g2_inv_1 \ring_501.inv_array[338]/sky_inverter/_0_  (.Y(\ring_501.inv_in[339] ),
    .A(\ring_501.inv_in[338] ));
 sg13g2_inv_1 \ring_501.inv_array[339]/sky_inverter/_0_  (.Y(\ring_501.inv_in[340] ),
    .A(\ring_501.inv_in[339] ));
 sg13g2_inv_1 \ring_501.inv_array[33]/sky_inverter/_0_  (.Y(\ring_501.inv_in[34] ),
    .A(\ring_501.inv_in[33] ));
 sg13g2_inv_1 \ring_501.inv_array[340]/sky_inverter/_0_  (.Y(\ring_501.inv_in[341] ),
    .A(\ring_501.inv_in[340] ));
 sg13g2_inv_1 \ring_501.inv_array[341]/sky_inverter/_0_  (.Y(\ring_501.inv_in[342] ),
    .A(\ring_501.inv_in[341] ));
 sg13g2_inv_1 \ring_501.inv_array[342]/sky_inverter/_0_  (.Y(\ring_501.inv_in[343] ),
    .A(\ring_501.inv_in[342] ));
 sg13g2_inv_1 \ring_501.inv_array[343]/sky_inverter/_0_  (.Y(\ring_501.inv_in[344] ),
    .A(\ring_501.inv_in[343] ));
 sg13g2_inv_1 \ring_501.inv_array[344]/sky_inverter/_0_  (.Y(\ring_501.inv_in[345] ),
    .A(\ring_501.inv_in[344] ));
 sg13g2_inv_1 \ring_501.inv_array[345]/sky_inverter/_0_  (.Y(\ring_501.inv_in[346] ),
    .A(\ring_501.inv_in[345] ));
 sg13g2_inv_1 \ring_501.inv_array[346]/sky_inverter/_0_  (.Y(\ring_501.inv_in[347] ),
    .A(\ring_501.inv_in[346] ));
 sg13g2_inv_1 \ring_501.inv_array[347]/sky_inverter/_0_  (.Y(\ring_501.inv_in[348] ),
    .A(\ring_501.inv_in[347] ));
 sg13g2_inv_1 \ring_501.inv_array[348]/sky_inverter/_0_  (.Y(\ring_501.inv_in[349] ),
    .A(\ring_501.inv_in[348] ));
 sg13g2_inv_1 \ring_501.inv_array[349]/sky_inverter/_0_  (.Y(\ring_501.inv_in[350] ),
    .A(\ring_501.inv_in[349] ));
 sg13g2_inv_1 \ring_501.inv_array[34]/sky_inverter/_0_  (.Y(\ring_501.inv_in[35] ),
    .A(\ring_501.inv_in[34] ));
 sg13g2_inv_1 \ring_501.inv_array[350]/sky_inverter/_0_  (.Y(\ring_501.inv_in[351] ),
    .A(\ring_501.inv_in[350] ));
 sg13g2_inv_1 \ring_501.inv_array[351]/sky_inverter/_0_  (.Y(\ring_501.inv_in[352] ),
    .A(\ring_501.inv_in[351] ));
 sg13g2_inv_1 \ring_501.inv_array[352]/sky_inverter/_0_  (.Y(\ring_501.inv_in[353] ),
    .A(\ring_501.inv_in[352] ));
 sg13g2_inv_1 \ring_501.inv_array[353]/sky_inverter/_0_  (.Y(\ring_501.inv_in[354] ),
    .A(\ring_501.inv_in[353] ));
 sg13g2_inv_1 \ring_501.inv_array[354]/sky_inverter/_0_  (.Y(\ring_501.inv_in[355] ),
    .A(\ring_501.inv_in[354] ));
 sg13g2_inv_1 \ring_501.inv_array[355]/sky_inverter/_0_  (.Y(\ring_501.inv_in[356] ),
    .A(\ring_501.inv_in[355] ));
 sg13g2_inv_1 \ring_501.inv_array[356]/sky_inverter/_0_  (.Y(\ring_501.inv_in[357] ),
    .A(\ring_501.inv_in[356] ));
 sg13g2_inv_1 \ring_501.inv_array[357]/sky_inverter/_0_  (.Y(\ring_501.inv_in[358] ),
    .A(\ring_501.inv_in[357] ));
 sg13g2_inv_1 \ring_501.inv_array[358]/sky_inverter/_0_  (.Y(\ring_501.inv_in[359] ),
    .A(\ring_501.inv_in[358] ));
 sg13g2_inv_1 \ring_501.inv_array[359]/sky_inverter/_0_  (.Y(\ring_501.inv_in[360] ),
    .A(\ring_501.inv_in[359] ));
 sg13g2_inv_1 \ring_501.inv_array[35]/sky_inverter/_0_  (.Y(\ring_501.inv_in[36] ),
    .A(\ring_501.inv_in[35] ));
 sg13g2_inv_1 \ring_501.inv_array[360]/sky_inverter/_0_  (.Y(\ring_501.inv_in[361] ),
    .A(\ring_501.inv_in[360] ));
 sg13g2_inv_1 \ring_501.inv_array[361]/sky_inverter/_0_  (.Y(\ring_501.inv_in[362] ),
    .A(\ring_501.inv_in[361] ));
 sg13g2_inv_1 \ring_501.inv_array[362]/sky_inverter/_0_  (.Y(\ring_501.inv_in[363] ),
    .A(\ring_501.inv_in[362] ));
 sg13g2_inv_1 \ring_501.inv_array[363]/sky_inverter/_0_  (.Y(\ring_501.inv_in[364] ),
    .A(\ring_501.inv_in[363] ));
 sg13g2_inv_1 \ring_501.inv_array[364]/sky_inverter/_0_  (.Y(\ring_501.inv_in[365] ),
    .A(\ring_501.inv_in[364] ));
 sg13g2_inv_1 \ring_501.inv_array[365]/sky_inverter/_0_  (.Y(\ring_501.inv_in[366] ),
    .A(\ring_501.inv_in[365] ));
 sg13g2_inv_1 \ring_501.inv_array[366]/sky_inverter/_0_  (.Y(\ring_501.inv_in[367] ),
    .A(\ring_501.inv_in[366] ));
 sg13g2_inv_1 \ring_501.inv_array[367]/sky_inverter/_0_  (.Y(\ring_501.inv_in[368] ),
    .A(\ring_501.inv_in[367] ));
 sg13g2_inv_1 \ring_501.inv_array[368]/sky_inverter/_0_  (.Y(\ring_501.inv_in[369] ),
    .A(\ring_501.inv_in[368] ));
 sg13g2_inv_1 \ring_501.inv_array[369]/sky_inverter/_0_  (.Y(\ring_501.inv_in[370] ),
    .A(\ring_501.inv_in[369] ));
 sg13g2_inv_1 \ring_501.inv_array[36]/sky_inverter/_0_  (.Y(\ring_501.inv_in[37] ),
    .A(\ring_501.inv_in[36] ));
 sg13g2_inv_1 \ring_501.inv_array[370]/sky_inverter/_0_  (.Y(\ring_501.inv_in[371] ),
    .A(\ring_501.inv_in[370] ));
 sg13g2_inv_1 \ring_501.inv_array[371]/sky_inverter/_0_  (.Y(\ring_501.inv_in[372] ),
    .A(\ring_501.inv_in[371] ));
 sg13g2_inv_1 \ring_501.inv_array[372]/sky_inverter/_0_  (.Y(\ring_501.inv_in[373] ),
    .A(\ring_501.inv_in[372] ));
 sg13g2_inv_1 \ring_501.inv_array[373]/sky_inverter/_0_  (.Y(\ring_501.inv_in[374] ),
    .A(\ring_501.inv_in[373] ));
 sg13g2_inv_1 \ring_501.inv_array[374]/sky_inverter/_0_  (.Y(\ring_501.inv_in[375] ),
    .A(\ring_501.inv_in[374] ));
 sg13g2_inv_1 \ring_501.inv_array[375]/sky_inverter/_0_  (.Y(\ring_501.inv_in[376] ),
    .A(\ring_501.inv_in[375] ));
 sg13g2_inv_1 \ring_501.inv_array[376]/sky_inverter/_0_  (.Y(\ring_501.inv_in[377] ),
    .A(\ring_501.inv_in[376] ));
 sg13g2_inv_1 \ring_501.inv_array[377]/sky_inverter/_0_  (.Y(\ring_501.inv_in[378] ),
    .A(\ring_501.inv_in[377] ));
 sg13g2_inv_1 \ring_501.inv_array[378]/sky_inverter/_0_  (.Y(\ring_501.inv_in[379] ),
    .A(\ring_501.inv_in[378] ));
 sg13g2_inv_1 \ring_501.inv_array[379]/sky_inverter/_0_  (.Y(\ring_501.inv_in[380] ),
    .A(\ring_501.inv_in[379] ));
 sg13g2_inv_1 \ring_501.inv_array[37]/sky_inverter/_0_  (.Y(\ring_501.inv_in[38] ),
    .A(\ring_501.inv_in[37] ));
 sg13g2_inv_1 \ring_501.inv_array[380]/sky_inverter/_0_  (.Y(\ring_501.inv_in[381] ),
    .A(\ring_501.inv_in[380] ));
 sg13g2_inv_1 \ring_501.inv_array[381]/sky_inverter/_0_  (.Y(\ring_501.inv_in[382] ),
    .A(\ring_501.inv_in[381] ));
 sg13g2_inv_1 \ring_501.inv_array[382]/sky_inverter/_0_  (.Y(\ring_501.inv_in[383] ),
    .A(\ring_501.inv_in[382] ));
 sg13g2_inv_1 \ring_501.inv_array[383]/sky_inverter/_0_  (.Y(\ring_501.inv_in[384] ),
    .A(\ring_501.inv_in[383] ));
 sg13g2_inv_1 \ring_501.inv_array[384]/sky_inverter/_0_  (.Y(\ring_501.inv_in[385] ),
    .A(\ring_501.inv_in[384] ));
 sg13g2_inv_1 \ring_501.inv_array[385]/sky_inverter/_0_  (.Y(\ring_501.inv_in[386] ),
    .A(\ring_501.inv_in[385] ));
 sg13g2_inv_1 \ring_501.inv_array[386]/sky_inverter/_0_  (.Y(\ring_501.inv_in[387] ),
    .A(\ring_501.inv_in[386] ));
 sg13g2_inv_1 \ring_501.inv_array[387]/sky_inverter/_0_  (.Y(\ring_501.inv_in[388] ),
    .A(\ring_501.inv_in[387] ));
 sg13g2_inv_1 \ring_501.inv_array[388]/sky_inverter/_0_  (.Y(\ring_501.inv_in[389] ),
    .A(\ring_501.inv_in[388] ));
 sg13g2_inv_1 \ring_501.inv_array[389]/sky_inverter/_0_  (.Y(\ring_501.inv_in[390] ),
    .A(\ring_501.inv_in[389] ));
 sg13g2_inv_1 \ring_501.inv_array[38]/sky_inverter/_0_  (.Y(\ring_501.inv_in[39] ),
    .A(\ring_501.inv_in[38] ));
 sg13g2_inv_1 \ring_501.inv_array[390]/sky_inverter/_0_  (.Y(\ring_501.inv_in[391] ),
    .A(\ring_501.inv_in[390] ));
 sg13g2_inv_1 \ring_501.inv_array[391]/sky_inverter/_0_  (.Y(\ring_501.inv_in[392] ),
    .A(\ring_501.inv_in[391] ));
 sg13g2_inv_1 \ring_501.inv_array[392]/sky_inverter/_0_  (.Y(\ring_501.inv_in[393] ),
    .A(\ring_501.inv_in[392] ));
 sg13g2_inv_1 \ring_501.inv_array[393]/sky_inverter/_0_  (.Y(\ring_501.inv_in[394] ),
    .A(\ring_501.inv_in[393] ));
 sg13g2_inv_1 \ring_501.inv_array[394]/sky_inverter/_0_  (.Y(\ring_501.inv_in[395] ),
    .A(\ring_501.inv_in[394] ));
 sg13g2_inv_1 \ring_501.inv_array[395]/sky_inverter/_0_  (.Y(\ring_501.inv_in[396] ),
    .A(\ring_501.inv_in[395] ));
 sg13g2_inv_1 \ring_501.inv_array[396]/sky_inverter/_0_  (.Y(\ring_501.inv_in[397] ),
    .A(\ring_501.inv_in[396] ));
 sg13g2_inv_1 \ring_501.inv_array[397]/sky_inverter/_0_  (.Y(\ring_501.inv_in[398] ),
    .A(\ring_501.inv_in[397] ));
 sg13g2_inv_1 \ring_501.inv_array[398]/sky_inverter/_0_  (.Y(\ring_501.inv_in[399] ),
    .A(\ring_501.inv_in[398] ));
 sg13g2_inv_1 \ring_501.inv_array[399]/sky_inverter/_0_  (.Y(\ring_501.inv_in[400] ),
    .A(\ring_501.inv_in[399] ));
 sg13g2_inv_1 \ring_501.inv_array[39]/sky_inverter/_0_  (.Y(\ring_501.inv_in[40] ),
    .A(\ring_501.inv_in[39] ));
 sg13g2_inv_1 \ring_501.inv_array[3]/sky_inverter/_0_  (.Y(\ring_501.inv_in[4] ),
    .A(\ring_501.inv_in[3] ));
 sg13g2_inv_1 \ring_501.inv_array[400]/sky_inverter/_0_  (.Y(\ring_501.inv_in[401] ),
    .A(\ring_501.inv_in[400] ));
 sg13g2_inv_1 \ring_501.inv_array[401]/sky_inverter/_0_  (.Y(\ring_501.inv_in[402] ),
    .A(\ring_501.inv_in[401] ));
 sg13g2_inv_1 \ring_501.inv_array[402]/sky_inverter/_0_  (.Y(\ring_501.inv_in[403] ),
    .A(\ring_501.inv_in[402] ));
 sg13g2_inv_1 \ring_501.inv_array[403]/sky_inverter/_0_  (.Y(\ring_501.inv_in[404] ),
    .A(\ring_501.inv_in[403] ));
 sg13g2_inv_1 \ring_501.inv_array[404]/sky_inverter/_0_  (.Y(\ring_501.inv_in[405] ),
    .A(\ring_501.inv_in[404] ));
 sg13g2_inv_1 \ring_501.inv_array[405]/sky_inverter/_0_  (.Y(\ring_501.inv_in[406] ),
    .A(\ring_501.inv_in[405] ));
 sg13g2_inv_1 \ring_501.inv_array[406]/sky_inverter/_0_  (.Y(\ring_501.inv_in[407] ),
    .A(\ring_501.inv_in[406] ));
 sg13g2_inv_1 \ring_501.inv_array[407]/sky_inverter/_0_  (.Y(\ring_501.inv_in[408] ),
    .A(\ring_501.inv_in[407] ));
 sg13g2_inv_1 \ring_501.inv_array[408]/sky_inverter/_0_  (.Y(\ring_501.inv_in[409] ),
    .A(\ring_501.inv_in[408] ));
 sg13g2_inv_1 \ring_501.inv_array[409]/sky_inverter/_0_  (.Y(\ring_501.inv_in[410] ),
    .A(\ring_501.inv_in[409] ));
 sg13g2_inv_1 \ring_501.inv_array[40]/sky_inverter/_0_  (.Y(\ring_501.inv_in[41] ),
    .A(\ring_501.inv_in[40] ));
 sg13g2_inv_1 \ring_501.inv_array[410]/sky_inverter/_0_  (.Y(\ring_501.inv_in[411] ),
    .A(\ring_501.inv_in[410] ));
 sg13g2_inv_1 \ring_501.inv_array[411]/sky_inverter/_0_  (.Y(\ring_501.inv_in[412] ),
    .A(\ring_501.inv_in[411] ));
 sg13g2_inv_1 \ring_501.inv_array[412]/sky_inverter/_0_  (.Y(\ring_501.inv_in[413] ),
    .A(\ring_501.inv_in[412] ));
 sg13g2_inv_1 \ring_501.inv_array[413]/sky_inverter/_0_  (.Y(\ring_501.inv_in[414] ),
    .A(\ring_501.inv_in[413] ));
 sg13g2_inv_1 \ring_501.inv_array[414]/sky_inverter/_0_  (.Y(\ring_501.inv_in[415] ),
    .A(\ring_501.inv_in[414] ));
 sg13g2_inv_1 \ring_501.inv_array[415]/sky_inverter/_0_  (.Y(\ring_501.inv_in[416] ),
    .A(\ring_501.inv_in[415] ));
 sg13g2_inv_1 \ring_501.inv_array[416]/sky_inverter/_0_  (.Y(\ring_501.inv_in[417] ),
    .A(\ring_501.inv_in[416] ));
 sg13g2_inv_1 \ring_501.inv_array[417]/sky_inverter/_0_  (.Y(\ring_501.inv_in[418] ),
    .A(\ring_501.inv_in[417] ));
 sg13g2_inv_1 \ring_501.inv_array[418]/sky_inverter/_0_  (.Y(\ring_501.inv_in[419] ),
    .A(\ring_501.inv_in[418] ));
 sg13g2_inv_1 \ring_501.inv_array[419]/sky_inverter/_0_  (.Y(\ring_501.inv_in[420] ),
    .A(\ring_501.inv_in[419] ));
 sg13g2_inv_1 \ring_501.inv_array[41]/sky_inverter/_0_  (.Y(\ring_501.inv_in[42] ),
    .A(\ring_501.inv_in[41] ));
 sg13g2_inv_1 \ring_501.inv_array[420]/sky_inverter/_0_  (.Y(\ring_501.inv_in[421] ),
    .A(\ring_501.inv_in[420] ));
 sg13g2_inv_1 \ring_501.inv_array[421]/sky_inverter/_0_  (.Y(\ring_501.inv_in[422] ),
    .A(\ring_501.inv_in[421] ));
 sg13g2_inv_1 \ring_501.inv_array[422]/sky_inverter/_0_  (.Y(\ring_501.inv_in[423] ),
    .A(\ring_501.inv_in[422] ));
 sg13g2_inv_1 \ring_501.inv_array[423]/sky_inverter/_0_  (.Y(\ring_501.inv_in[424] ),
    .A(\ring_501.inv_in[423] ));
 sg13g2_inv_1 \ring_501.inv_array[424]/sky_inverter/_0_  (.Y(\ring_501.inv_in[425] ),
    .A(\ring_501.inv_in[424] ));
 sg13g2_inv_1 \ring_501.inv_array[425]/sky_inverter/_0_  (.Y(\ring_501.inv_in[426] ),
    .A(\ring_501.inv_in[425] ));
 sg13g2_inv_1 \ring_501.inv_array[426]/sky_inverter/_0_  (.Y(\ring_501.inv_in[427] ),
    .A(\ring_501.inv_in[426] ));
 sg13g2_inv_1 \ring_501.inv_array[427]/sky_inverter/_0_  (.Y(\ring_501.inv_in[428] ),
    .A(\ring_501.inv_in[427] ));
 sg13g2_inv_1 \ring_501.inv_array[428]/sky_inverter/_0_  (.Y(\ring_501.inv_in[429] ),
    .A(\ring_501.inv_in[428] ));
 sg13g2_inv_1 \ring_501.inv_array[429]/sky_inverter/_0_  (.Y(\ring_501.inv_in[430] ),
    .A(\ring_501.inv_in[429] ));
 sg13g2_inv_1 \ring_501.inv_array[42]/sky_inverter/_0_  (.Y(\ring_501.inv_in[43] ),
    .A(\ring_501.inv_in[42] ));
 sg13g2_inv_1 \ring_501.inv_array[430]/sky_inverter/_0_  (.Y(\ring_501.inv_in[431] ),
    .A(\ring_501.inv_in[430] ));
 sg13g2_inv_1 \ring_501.inv_array[431]/sky_inverter/_0_  (.Y(\ring_501.inv_in[432] ),
    .A(\ring_501.inv_in[431] ));
 sg13g2_inv_1 \ring_501.inv_array[432]/sky_inverter/_0_  (.Y(\ring_501.inv_in[433] ),
    .A(\ring_501.inv_in[432] ));
 sg13g2_inv_1 \ring_501.inv_array[433]/sky_inverter/_0_  (.Y(\ring_501.inv_in[434] ),
    .A(\ring_501.inv_in[433] ));
 sg13g2_inv_1 \ring_501.inv_array[434]/sky_inverter/_0_  (.Y(\ring_501.inv_in[435] ),
    .A(\ring_501.inv_in[434] ));
 sg13g2_inv_1 \ring_501.inv_array[435]/sky_inverter/_0_  (.Y(\ring_501.inv_in[436] ),
    .A(\ring_501.inv_in[435] ));
 sg13g2_inv_1 \ring_501.inv_array[436]/sky_inverter/_0_  (.Y(\ring_501.inv_in[437] ),
    .A(\ring_501.inv_in[436] ));
 sg13g2_inv_1 \ring_501.inv_array[437]/sky_inverter/_0_  (.Y(\ring_501.inv_in[438] ),
    .A(\ring_501.inv_in[437] ));
 sg13g2_inv_1 \ring_501.inv_array[438]/sky_inverter/_0_  (.Y(\ring_501.inv_in[439] ),
    .A(\ring_501.inv_in[438] ));
 sg13g2_inv_1 \ring_501.inv_array[439]/sky_inverter/_0_  (.Y(\ring_501.inv_in[440] ),
    .A(\ring_501.inv_in[439] ));
 sg13g2_inv_1 \ring_501.inv_array[43]/sky_inverter/_0_  (.Y(\ring_501.inv_in[44] ),
    .A(\ring_501.inv_in[43] ));
 sg13g2_inv_1 \ring_501.inv_array[440]/sky_inverter/_0_  (.Y(\ring_501.inv_in[441] ),
    .A(\ring_501.inv_in[440] ));
 sg13g2_inv_1 \ring_501.inv_array[441]/sky_inverter/_0_  (.Y(\ring_501.inv_in[442] ),
    .A(\ring_501.inv_in[441] ));
 sg13g2_inv_1 \ring_501.inv_array[442]/sky_inverter/_0_  (.Y(\ring_501.inv_in[443] ),
    .A(\ring_501.inv_in[442] ));
 sg13g2_inv_1 \ring_501.inv_array[443]/sky_inverter/_0_  (.Y(\ring_501.inv_in[444] ),
    .A(\ring_501.inv_in[443] ));
 sg13g2_inv_1 \ring_501.inv_array[444]/sky_inverter/_0_  (.Y(\ring_501.inv_in[445] ),
    .A(\ring_501.inv_in[444] ));
 sg13g2_inv_1 \ring_501.inv_array[445]/sky_inverter/_0_  (.Y(\ring_501.inv_in[446] ),
    .A(\ring_501.inv_in[445] ));
 sg13g2_inv_1 \ring_501.inv_array[446]/sky_inverter/_0_  (.Y(\ring_501.inv_in[447] ),
    .A(\ring_501.inv_in[446] ));
 sg13g2_inv_1 \ring_501.inv_array[447]/sky_inverter/_0_  (.Y(\ring_501.inv_in[448] ),
    .A(\ring_501.inv_in[447] ));
 sg13g2_inv_1 \ring_501.inv_array[448]/sky_inverter/_0_  (.Y(\ring_501.inv_in[449] ),
    .A(\ring_501.inv_in[448] ));
 sg13g2_inv_1 \ring_501.inv_array[449]/sky_inverter/_0_  (.Y(\ring_501.inv_in[450] ),
    .A(\ring_501.inv_in[449] ));
 sg13g2_inv_1 \ring_501.inv_array[44]/sky_inverter/_0_  (.Y(\ring_501.inv_in[45] ),
    .A(\ring_501.inv_in[44] ));
 sg13g2_inv_1 \ring_501.inv_array[450]/sky_inverter/_0_  (.Y(\ring_501.inv_in[451] ),
    .A(\ring_501.inv_in[450] ));
 sg13g2_inv_1 \ring_501.inv_array[451]/sky_inverter/_0_  (.Y(\ring_501.inv_in[452] ),
    .A(\ring_501.inv_in[451] ));
 sg13g2_inv_1 \ring_501.inv_array[452]/sky_inverter/_0_  (.Y(\ring_501.inv_in[453] ),
    .A(\ring_501.inv_in[452] ));
 sg13g2_inv_1 \ring_501.inv_array[453]/sky_inverter/_0_  (.Y(\ring_501.inv_in[454] ),
    .A(\ring_501.inv_in[453] ));
 sg13g2_inv_1 \ring_501.inv_array[454]/sky_inverter/_0_  (.Y(\ring_501.inv_in[455] ),
    .A(\ring_501.inv_in[454] ));
 sg13g2_inv_1 \ring_501.inv_array[455]/sky_inverter/_0_  (.Y(\ring_501.inv_in[456] ),
    .A(\ring_501.inv_in[455] ));
 sg13g2_inv_1 \ring_501.inv_array[456]/sky_inverter/_0_  (.Y(\ring_501.inv_in[457] ),
    .A(\ring_501.inv_in[456] ));
 sg13g2_inv_1 \ring_501.inv_array[457]/sky_inverter/_0_  (.Y(\ring_501.inv_in[458] ),
    .A(\ring_501.inv_in[457] ));
 sg13g2_inv_1 \ring_501.inv_array[458]/sky_inverter/_0_  (.Y(\ring_501.inv_in[459] ),
    .A(\ring_501.inv_in[458] ));
 sg13g2_inv_1 \ring_501.inv_array[459]/sky_inverter/_0_  (.Y(\ring_501.inv_in[460] ),
    .A(\ring_501.inv_in[459] ));
 sg13g2_inv_1 \ring_501.inv_array[45]/sky_inverter/_0_  (.Y(\ring_501.inv_in[46] ),
    .A(\ring_501.inv_in[45] ));
 sg13g2_inv_1 \ring_501.inv_array[460]/sky_inverter/_0_  (.Y(\ring_501.inv_in[461] ),
    .A(\ring_501.inv_in[460] ));
 sg13g2_inv_1 \ring_501.inv_array[461]/sky_inverter/_0_  (.Y(\ring_501.inv_in[462] ),
    .A(\ring_501.inv_in[461] ));
 sg13g2_inv_1 \ring_501.inv_array[462]/sky_inverter/_0_  (.Y(\ring_501.inv_in[463] ),
    .A(\ring_501.inv_in[462] ));
 sg13g2_inv_1 \ring_501.inv_array[463]/sky_inverter/_0_  (.Y(\ring_501.inv_in[464] ),
    .A(\ring_501.inv_in[463] ));
 sg13g2_inv_1 \ring_501.inv_array[464]/sky_inverter/_0_  (.Y(\ring_501.inv_in[465] ),
    .A(\ring_501.inv_in[464] ));
 sg13g2_inv_1 \ring_501.inv_array[465]/sky_inverter/_0_  (.Y(\ring_501.inv_in[466] ),
    .A(\ring_501.inv_in[465] ));
 sg13g2_inv_1 \ring_501.inv_array[466]/sky_inverter/_0_  (.Y(\ring_501.inv_in[467] ),
    .A(\ring_501.inv_in[466] ));
 sg13g2_inv_1 \ring_501.inv_array[467]/sky_inverter/_0_  (.Y(\ring_501.inv_in[468] ),
    .A(\ring_501.inv_in[467] ));
 sg13g2_inv_1 \ring_501.inv_array[468]/sky_inverter/_0_  (.Y(\ring_501.inv_in[469] ),
    .A(\ring_501.inv_in[468] ));
 sg13g2_inv_1 \ring_501.inv_array[469]/sky_inverter/_0_  (.Y(\ring_501.inv_in[470] ),
    .A(\ring_501.inv_in[469] ));
 sg13g2_inv_1 \ring_501.inv_array[46]/sky_inverter/_0_  (.Y(\ring_501.inv_in[47] ),
    .A(\ring_501.inv_in[46] ));
 sg13g2_inv_1 \ring_501.inv_array[470]/sky_inverter/_0_  (.Y(\ring_501.inv_in[471] ),
    .A(\ring_501.inv_in[470] ));
 sg13g2_inv_1 \ring_501.inv_array[471]/sky_inverter/_0_  (.Y(\ring_501.inv_in[472] ),
    .A(\ring_501.inv_in[471] ));
 sg13g2_inv_1 \ring_501.inv_array[472]/sky_inverter/_0_  (.Y(\ring_501.inv_in[473] ),
    .A(\ring_501.inv_in[472] ));
 sg13g2_inv_1 \ring_501.inv_array[473]/sky_inverter/_0_  (.Y(\ring_501.inv_in[474] ),
    .A(\ring_501.inv_in[473] ));
 sg13g2_inv_1 \ring_501.inv_array[474]/sky_inverter/_0_  (.Y(\ring_501.inv_in[475] ),
    .A(\ring_501.inv_in[474] ));
 sg13g2_inv_1 \ring_501.inv_array[475]/sky_inverter/_0_  (.Y(\ring_501.inv_in[476] ),
    .A(\ring_501.inv_in[475] ));
 sg13g2_inv_1 \ring_501.inv_array[476]/sky_inverter/_0_  (.Y(\ring_501.inv_in[477] ),
    .A(\ring_501.inv_in[476] ));
 sg13g2_inv_1 \ring_501.inv_array[477]/sky_inverter/_0_  (.Y(\ring_501.inv_in[478] ),
    .A(\ring_501.inv_in[477] ));
 sg13g2_inv_1 \ring_501.inv_array[478]/sky_inverter/_0_  (.Y(\ring_501.inv_in[479] ),
    .A(\ring_501.inv_in[478] ));
 sg13g2_inv_1 \ring_501.inv_array[479]/sky_inverter/_0_  (.Y(\ring_501.inv_in[480] ),
    .A(\ring_501.inv_in[479] ));
 sg13g2_inv_1 \ring_501.inv_array[47]/sky_inverter/_0_  (.Y(\ring_501.inv_in[48] ),
    .A(\ring_501.inv_in[47] ));
 sg13g2_inv_1 \ring_501.inv_array[480]/sky_inverter/_0_  (.Y(\ring_501.inv_in[481] ),
    .A(\ring_501.inv_in[480] ));
 sg13g2_inv_1 \ring_501.inv_array[481]/sky_inverter/_0_  (.Y(\ring_501.inv_in[482] ),
    .A(\ring_501.inv_in[481] ));
 sg13g2_inv_1 \ring_501.inv_array[482]/sky_inverter/_0_  (.Y(\ring_501.inv_in[483] ),
    .A(\ring_501.inv_in[482] ));
 sg13g2_inv_1 \ring_501.inv_array[483]/sky_inverter/_0_  (.Y(\ring_501.inv_in[484] ),
    .A(\ring_501.inv_in[483] ));
 sg13g2_inv_1 \ring_501.inv_array[484]/sky_inverter/_0_  (.Y(\ring_501.inv_in[485] ),
    .A(\ring_501.inv_in[484] ));
 sg13g2_inv_1 \ring_501.inv_array[485]/sky_inverter/_0_  (.Y(\ring_501.inv_in[486] ),
    .A(\ring_501.inv_in[485] ));
 sg13g2_inv_1 \ring_501.inv_array[486]/sky_inverter/_0_  (.Y(\ring_501.inv_in[487] ),
    .A(\ring_501.inv_in[486] ));
 sg13g2_inv_1 \ring_501.inv_array[487]/sky_inverter/_0_  (.Y(\ring_501.inv_in[488] ),
    .A(\ring_501.inv_in[487] ));
 sg13g2_inv_1 \ring_501.inv_array[488]/sky_inverter/_0_  (.Y(\ring_501.inv_in[489] ),
    .A(\ring_501.inv_in[488] ));
 sg13g2_inv_1 \ring_501.inv_array[489]/sky_inverter/_0_  (.Y(\ring_501.inv_in[490] ),
    .A(\ring_501.inv_in[489] ));
 sg13g2_inv_1 \ring_501.inv_array[48]/sky_inverter/_0_  (.Y(\ring_501.inv_in[49] ),
    .A(\ring_501.inv_in[48] ));
 sg13g2_inv_1 \ring_501.inv_array[490]/sky_inverter/_0_  (.Y(\ring_501.inv_in[491] ),
    .A(\ring_501.inv_in[490] ));
 sg13g2_inv_1 \ring_501.inv_array[491]/sky_inverter/_0_  (.Y(\ring_501.inv_in[492] ),
    .A(\ring_501.inv_in[491] ));
 sg13g2_inv_1 \ring_501.inv_array[492]/sky_inverter/_0_  (.Y(\ring_501.inv_in[493] ),
    .A(\ring_501.inv_in[492] ));
 sg13g2_inv_1 \ring_501.inv_array[493]/sky_inverter/_0_  (.Y(\ring_501.inv_in[494] ),
    .A(\ring_501.inv_in[493] ));
 sg13g2_inv_1 \ring_501.inv_array[494]/sky_inverter/_0_  (.Y(\ring_501.inv_in[495] ),
    .A(\ring_501.inv_in[494] ));
 sg13g2_inv_1 \ring_501.inv_array[495]/sky_inverter/_0_  (.Y(\ring_501.inv_in[496] ),
    .A(\ring_501.inv_in[495] ));
 sg13g2_inv_1 \ring_501.inv_array[496]/sky_inverter/_0_  (.Y(\ring_501.inv_in[497] ),
    .A(\ring_501.inv_in[496] ));
 sg13g2_inv_1 \ring_501.inv_array[497]/sky_inverter/_0_  (.Y(\ring_501.inv_in[498] ),
    .A(\ring_501.inv_in[497] ));
 sg13g2_inv_1 \ring_501.inv_array[498]/sky_inverter/_0_  (.Y(\ring_501.inv_in[499] ),
    .A(\ring_501.inv_in[498] ));
 sg13g2_inv_1 \ring_501.inv_array[499]/sky_inverter/_0_  (.Y(\ring_501.inv_in[500] ),
    .A(\ring_501.inv_in[499] ));
 sg13g2_inv_1 \ring_501.inv_array[49]/sky_inverter/_0_  (.Y(\ring_501.inv_in[50] ),
    .A(\ring_501.inv_in[49] ));
 sg13g2_inv_1 \ring_501.inv_array[4]/sky_inverter/_0_  (.Y(\ring_501.inv_in[5] ),
    .A(\ring_501.inv_in[4] ));
 sg13g2_inv_1 \ring_501.inv_array[500]/sky_inverter/_0_  (.Y(\ring_501.inv_out[500] ),
    .A(\ring_501.inv_in[500] ));
 sg13g2_inv_1 \ring_501.inv_array[50]/sky_inverter/_0_  (.Y(\ring_501.inv_in[51] ),
    .A(\ring_501.inv_in[50] ));
 sg13g2_inv_1 \ring_501.inv_array[51]/sky_inverter/_0_  (.Y(\ring_501.inv_in[52] ),
    .A(\ring_501.inv_in[51] ));
 sg13g2_inv_1 \ring_501.inv_array[52]/sky_inverter/_0_  (.Y(\ring_501.inv_in[53] ),
    .A(\ring_501.inv_in[52] ));
 sg13g2_inv_1 \ring_501.inv_array[53]/sky_inverter/_0_  (.Y(\ring_501.inv_in[54] ),
    .A(\ring_501.inv_in[53] ));
 sg13g2_inv_1 \ring_501.inv_array[54]/sky_inverter/_0_  (.Y(\ring_501.inv_in[55] ),
    .A(\ring_501.inv_in[54] ));
 sg13g2_inv_1 \ring_501.inv_array[55]/sky_inverter/_0_  (.Y(\ring_501.inv_in[56] ),
    .A(\ring_501.inv_in[55] ));
 sg13g2_inv_1 \ring_501.inv_array[56]/sky_inverter/_0_  (.Y(\ring_501.inv_in[57] ),
    .A(\ring_501.inv_in[56] ));
 sg13g2_inv_1 \ring_501.inv_array[57]/sky_inverter/_0_  (.Y(\ring_501.inv_in[58] ),
    .A(\ring_501.inv_in[57] ));
 sg13g2_inv_1 \ring_501.inv_array[58]/sky_inverter/_0_  (.Y(\ring_501.inv_in[59] ),
    .A(\ring_501.inv_in[58] ));
 sg13g2_inv_1 \ring_501.inv_array[59]/sky_inverter/_0_  (.Y(\ring_501.inv_in[60] ),
    .A(\ring_501.inv_in[59] ));
 sg13g2_inv_1 \ring_501.inv_array[5]/sky_inverter/_0_  (.Y(\ring_501.inv_in[6] ),
    .A(\ring_501.inv_in[5] ));
 sg13g2_inv_1 \ring_501.inv_array[60]/sky_inverter/_0_  (.Y(\ring_501.inv_in[61] ),
    .A(\ring_501.inv_in[60] ));
 sg13g2_inv_1 \ring_501.inv_array[61]/sky_inverter/_0_  (.Y(\ring_501.inv_in[62] ),
    .A(\ring_501.inv_in[61] ));
 sg13g2_inv_1 \ring_501.inv_array[62]/sky_inverter/_0_  (.Y(\ring_501.inv_in[63] ),
    .A(\ring_501.inv_in[62] ));
 sg13g2_inv_1 \ring_501.inv_array[63]/sky_inverter/_0_  (.Y(\ring_501.inv_in[64] ),
    .A(\ring_501.inv_in[63] ));
 sg13g2_inv_1 \ring_501.inv_array[64]/sky_inverter/_0_  (.Y(\ring_501.inv_in[65] ),
    .A(\ring_501.inv_in[64] ));
 sg13g2_inv_1 \ring_501.inv_array[65]/sky_inverter/_0_  (.Y(\ring_501.inv_in[66] ),
    .A(\ring_501.inv_in[65] ));
 sg13g2_inv_1 \ring_501.inv_array[66]/sky_inverter/_0_  (.Y(\ring_501.inv_in[67] ),
    .A(\ring_501.inv_in[66] ));
 sg13g2_inv_1 \ring_501.inv_array[67]/sky_inverter/_0_  (.Y(\ring_501.inv_in[68] ),
    .A(\ring_501.inv_in[67] ));
 sg13g2_inv_1 \ring_501.inv_array[68]/sky_inverter/_0_  (.Y(\ring_501.inv_in[69] ),
    .A(\ring_501.inv_in[68] ));
 sg13g2_inv_1 \ring_501.inv_array[69]/sky_inverter/_0_  (.Y(\ring_501.inv_in[70] ),
    .A(\ring_501.inv_in[69] ));
 sg13g2_inv_1 \ring_501.inv_array[6]/sky_inverter/_0_  (.Y(\ring_501.inv_in[7] ),
    .A(\ring_501.inv_in[6] ));
 sg13g2_inv_1 \ring_501.inv_array[70]/sky_inverter/_0_  (.Y(\ring_501.inv_in[71] ),
    .A(\ring_501.inv_in[70] ));
 sg13g2_inv_1 \ring_501.inv_array[71]/sky_inverter/_0_  (.Y(\ring_501.inv_in[72] ),
    .A(\ring_501.inv_in[71] ));
 sg13g2_inv_1 \ring_501.inv_array[72]/sky_inverter/_0_  (.Y(\ring_501.inv_in[73] ),
    .A(\ring_501.inv_in[72] ));
 sg13g2_inv_1 \ring_501.inv_array[73]/sky_inverter/_0_  (.Y(\ring_501.inv_in[74] ),
    .A(\ring_501.inv_in[73] ));
 sg13g2_inv_1 \ring_501.inv_array[74]/sky_inverter/_0_  (.Y(\ring_501.inv_in[75] ),
    .A(\ring_501.inv_in[74] ));
 sg13g2_inv_1 \ring_501.inv_array[75]/sky_inverter/_0_  (.Y(\ring_501.inv_in[76] ),
    .A(\ring_501.inv_in[75] ));
 sg13g2_inv_1 \ring_501.inv_array[76]/sky_inverter/_0_  (.Y(\ring_501.inv_in[77] ),
    .A(\ring_501.inv_in[76] ));
 sg13g2_inv_1 \ring_501.inv_array[77]/sky_inverter/_0_  (.Y(\ring_501.inv_in[78] ),
    .A(\ring_501.inv_in[77] ));
 sg13g2_inv_1 \ring_501.inv_array[78]/sky_inverter/_0_  (.Y(\ring_501.inv_in[79] ),
    .A(\ring_501.inv_in[78] ));
 sg13g2_inv_1 \ring_501.inv_array[79]/sky_inverter/_0_  (.Y(\ring_501.inv_in[80] ),
    .A(\ring_501.inv_in[79] ));
 sg13g2_inv_1 \ring_501.inv_array[7]/sky_inverter/_0_  (.Y(\ring_501.inv_in[8] ),
    .A(\ring_501.inv_in[7] ));
 sg13g2_inv_1 \ring_501.inv_array[80]/sky_inverter/_0_  (.Y(\ring_501.inv_in[81] ),
    .A(\ring_501.inv_in[80] ));
 sg13g2_inv_1 \ring_501.inv_array[81]/sky_inverter/_0_  (.Y(\ring_501.inv_in[82] ),
    .A(\ring_501.inv_in[81] ));
 sg13g2_inv_1 \ring_501.inv_array[82]/sky_inverter/_0_  (.Y(\ring_501.inv_in[83] ),
    .A(\ring_501.inv_in[82] ));
 sg13g2_inv_1 \ring_501.inv_array[83]/sky_inverter/_0_  (.Y(\ring_501.inv_in[84] ),
    .A(\ring_501.inv_in[83] ));
 sg13g2_inv_1 \ring_501.inv_array[84]/sky_inverter/_0_  (.Y(\ring_501.inv_in[85] ),
    .A(\ring_501.inv_in[84] ));
 sg13g2_inv_1 \ring_501.inv_array[85]/sky_inverter/_0_  (.Y(\ring_501.inv_in[86] ),
    .A(\ring_501.inv_in[85] ));
 sg13g2_inv_1 \ring_501.inv_array[86]/sky_inverter/_0_  (.Y(\ring_501.inv_in[87] ),
    .A(\ring_501.inv_in[86] ));
 sg13g2_inv_1 \ring_501.inv_array[87]/sky_inverter/_0_  (.Y(\ring_501.inv_in[88] ),
    .A(\ring_501.inv_in[87] ));
 sg13g2_inv_1 \ring_501.inv_array[88]/sky_inverter/_0_  (.Y(\ring_501.inv_in[89] ),
    .A(\ring_501.inv_in[88] ));
 sg13g2_inv_1 \ring_501.inv_array[89]/sky_inverter/_0_  (.Y(\ring_501.inv_in[90] ),
    .A(\ring_501.inv_in[89] ));
 sg13g2_inv_1 \ring_501.inv_array[8]/sky_inverter/_0_  (.Y(\ring_501.inv_in[9] ),
    .A(\ring_501.inv_in[8] ));
 sg13g2_inv_1 \ring_501.inv_array[90]/sky_inverter/_0_  (.Y(\ring_501.inv_in[91] ),
    .A(\ring_501.inv_in[90] ));
 sg13g2_inv_1 \ring_501.inv_array[91]/sky_inverter/_0_  (.Y(\ring_501.inv_in[92] ),
    .A(\ring_501.inv_in[91] ));
 sg13g2_inv_1 \ring_501.inv_array[92]/sky_inverter/_0_  (.Y(\ring_501.inv_in[93] ),
    .A(\ring_501.inv_in[92] ));
 sg13g2_inv_1 \ring_501.inv_array[93]/sky_inverter/_0_  (.Y(\ring_501.inv_in[94] ),
    .A(\ring_501.inv_in[93] ));
 sg13g2_inv_1 \ring_501.inv_array[94]/sky_inverter/_0_  (.Y(\ring_501.inv_in[95] ),
    .A(\ring_501.inv_in[94] ));
 sg13g2_inv_1 \ring_501.inv_array[95]/sky_inverter/_0_  (.Y(\ring_501.inv_in[96] ),
    .A(\ring_501.inv_in[95] ));
 sg13g2_inv_1 \ring_501.inv_array[96]/sky_inverter/_0_  (.Y(\ring_501.inv_in[97] ),
    .A(\ring_501.inv_in[96] ));
 sg13g2_inv_1 \ring_501.inv_array[97]/sky_inverter/_0_  (.Y(\ring_501.inv_in[98] ),
    .A(\ring_501.inv_in[97] ));
 sg13g2_inv_1 \ring_501.inv_array[98]/sky_inverter/_0_  (.Y(\ring_501.inv_in[99] ),
    .A(\ring_501.inv_in[98] ));
 sg13g2_inv_1 \ring_501.inv_array[99]/sky_inverter/_0_  (.Y(\ring_501.inv_in[100] ),
    .A(\ring_501.inv_in[99] ));
 sg13g2_inv_1 \ring_501.inv_array[9]/sky_inverter/_0_  (.Y(\ring_501.inv_in[10] ),
    .A(\ring_501.inv_in[9] ));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[0]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[2]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[3]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[4]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[5]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[6]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(ui_in[7]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[0]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[1]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[2]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[3]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[4]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[5]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(uio_in[6]),
    .X(net17));
 sg13g2_buf_1 input18 (.A(uio_in[7]),
    .X(net18));
 sg13g2_tielo tt_um_algofoogle_tt09_ring_osc2_19 (.L_LO(net19));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_4 FILLER_0_147 ();
 sg13g2_fill_2 FILLER_0_160 ();
 sg13g2_fill_2 FILLER_0_165 ();
 sg13g2_fill_1 FILLER_0_167 ();
 sg13g2_fill_2 FILLER_0_183 ();
 sg13g2_fill_1 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_4 FILLER_0_217 ();
 sg13g2_decap_4 FILLER_0_230 ();
 sg13g2_fill_1 FILLER_0_237 ();
 sg13g2_fill_1 FILLER_0_250 ();
 sg13g2_fill_1 FILLER_0_260 ();
 sg13g2_decap_8 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_293 ();
 sg13g2_decap_8 FILLER_0_300 ();
 sg13g2_decap_8 FILLER_0_307 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_8 FILLER_0_321 ();
 sg13g2_decap_8 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_4 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_fill_2 FILLER_1_140 ();
 sg13g2_fill_2 FILLER_1_205 ();
 sg13g2_fill_1 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_286 ();
 sg13g2_decap_8 FILLER_1_293 ();
 sg13g2_decap_8 FILLER_1_300 ();
 sg13g2_decap_8 FILLER_1_307 ();
 sg13g2_decap_8 FILLER_1_314 ();
 sg13g2_decap_8 FILLER_1_321 ();
 sg13g2_decap_8 FILLER_1_328 ();
 sg13g2_decap_8 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_342 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_162 ();
 sg13g2_decap_8 FILLER_2_169 ();
 sg13g2_fill_2 FILLER_2_176 ();
 sg13g2_fill_1 FILLER_2_178 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_4 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_212 ();
 sg13g2_decap_8 FILLER_2_219 ();
 sg13g2_decap_4 FILLER_2_226 ();
 sg13g2_fill_2 FILLER_2_230 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_fill_2 FILLER_2_259 ();
 sg13g2_fill_1 FILLER_2_261 ();
 sg13g2_fill_2 FILLER_2_265 ();
 sg13g2_fill_1 FILLER_2_267 ();
 sg13g2_fill_2 FILLER_2_271 ();
 sg13g2_decap_8 FILLER_2_285 ();
 sg13g2_decap_8 FILLER_2_292 ();
 sg13g2_decap_8 FILLER_2_299 ();
 sg13g2_decap_8 FILLER_2_306 ();
 sg13g2_decap_8 FILLER_2_313 ();
 sg13g2_decap_8 FILLER_2_320 ();
 sg13g2_decap_8 FILLER_2_327 ();
 sg13g2_decap_8 FILLER_2_334 ();
 sg13g2_decap_8 FILLER_2_341 ();
 sg13g2_decap_8 FILLER_2_348 ();
 sg13g2_decap_8 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_4 FILLER_2_404 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_195 ();
 sg13g2_decap_4 FILLER_3_202 ();
 sg13g2_fill_1 FILLER_3_206 ();
 sg13g2_fill_1 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_247 ();
 sg13g2_fill_2 FILLER_3_254 ();
 sg13g2_fill_1 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_fill_1 FILLER_4_133 ();
 sg13g2_decap_4 FILLER_4_137 ();
 sg13g2_fill_1 FILLER_4_141 ();
 sg13g2_fill_1 FILLER_4_145 ();
 sg13g2_fill_2 FILLER_4_149 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_4 FILLER_4_161 ();
 sg13g2_fill_2 FILLER_4_165 ();
 sg13g2_fill_2 FILLER_4_176 ();
 sg13g2_decap_8 FILLER_4_184 ();
 sg13g2_decap_8 FILLER_4_191 ();
 sg13g2_fill_1 FILLER_4_198 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_fill_2 FILLER_4_231 ();
 sg13g2_fill_1 FILLER_4_233 ();
 sg13g2_decap_8 FILLER_4_243 ();
 sg13g2_fill_2 FILLER_4_250 ();
 sg13g2_decap_8 FILLER_4_267 ();
 sg13g2_decap_8 FILLER_4_274 ();
 sg13g2_decap_8 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_288 ();
 sg13g2_decap_8 FILLER_4_295 ();
 sg13g2_decap_8 FILLER_4_302 ();
 sg13g2_decap_8 FILLER_4_309 ();
 sg13g2_decap_8 FILLER_4_316 ();
 sg13g2_decap_8 FILLER_4_323 ();
 sg13g2_decap_8 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_344 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_fill_2 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_161 ();
 sg13g2_fill_1 FILLER_5_174 ();
 sg13g2_fill_2 FILLER_5_181 ();
 sg13g2_fill_1 FILLER_5_183 ();
 sg13g2_decap_8 FILLER_5_187 ();
 sg13g2_decap_4 FILLER_5_194 ();
 sg13g2_fill_2 FILLER_5_198 ();
 sg13g2_fill_1 FILLER_5_218 ();
 sg13g2_decap_8 FILLER_5_222 ();
 sg13g2_fill_2 FILLER_5_229 ();
 sg13g2_fill_1 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_244 ();
 sg13g2_fill_2 FILLER_5_251 ();
 sg13g2_decap_8 FILLER_5_268 ();
 sg13g2_decap_8 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_282 ();
 sg13g2_decap_8 FILLER_5_289 ();
 sg13g2_decap_8 FILLER_5_296 ();
 sg13g2_decap_8 FILLER_5_303 ();
 sg13g2_decap_8 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_317 ();
 sg13g2_decap_8 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_331 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_fill_1 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_145 ();
 sg13g2_decap_8 FILLER_6_152 ();
 sg13g2_decap_4 FILLER_6_159 ();
 sg13g2_fill_1 FILLER_6_163 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_fill_2 FILLER_6_210 ();
 sg13g2_fill_1 FILLER_6_212 ();
 sg13g2_decap_4 FILLER_6_231 ();
 sg13g2_fill_1 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_4 FILLER_7_119 ();
 sg13g2_fill_1 FILLER_7_123 ();
 sg13g2_decap_8 FILLER_7_142 ();
 sg13g2_decap_8 FILLER_7_149 ();
 sg13g2_decap_8 FILLER_7_156 ();
 sg13g2_fill_2 FILLER_7_163 ();
 sg13g2_decap_8 FILLER_7_180 ();
 sg13g2_fill_1 FILLER_7_187 ();
 sg13g2_decap_8 FILLER_7_209 ();
 sg13g2_decap_4 FILLER_7_216 ();
 sg13g2_fill_1 FILLER_7_220 ();
 sg13g2_decap_8 FILLER_7_236 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_decap_8 FILLER_7_250 ();
 sg13g2_decap_8 FILLER_7_257 ();
 sg13g2_decap_8 FILLER_7_264 ();
 sg13g2_decap_8 FILLER_7_271 ();
 sg13g2_decap_8 FILLER_7_278 ();
 sg13g2_decap_8 FILLER_7_285 ();
 sg13g2_decap_8 FILLER_7_292 ();
 sg13g2_decap_8 FILLER_7_299 ();
 sg13g2_decap_8 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_327 ();
 sg13g2_decap_8 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_341 ();
 sg13g2_decap_8 FILLER_7_348 ();
 sg13g2_decap_8 FILLER_7_355 ();
 sg13g2_decap_8 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_369 ();
 sg13g2_decap_8 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_4 FILLER_8_126 ();
 sg13g2_fill_1 FILLER_8_130 ();
 sg13g2_decap_4 FILLER_8_179 ();
 sg13g2_fill_2 FILLER_8_183 ();
 sg13g2_decap_4 FILLER_8_188 ();
 sg13g2_fill_1 FILLER_8_192 ();
 sg13g2_decap_8 FILLER_8_214 ();
 sg13g2_fill_2 FILLER_8_221 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_fill_2 FILLER_9_145 ();
 sg13g2_fill_1 FILLER_9_147 ();
 sg13g2_decap_4 FILLER_9_151 ();
 sg13g2_fill_1 FILLER_9_155 ();
 sg13g2_fill_2 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_fill_2 FILLER_9_165 ();
 sg13g2_fill_1 FILLER_9_167 ();
 sg13g2_decap_8 FILLER_9_171 ();
 sg13g2_fill_1 FILLER_9_178 ();
 sg13g2_decap_8 FILLER_9_206 ();
 sg13g2_decap_8 FILLER_9_213 ();
 sg13g2_fill_2 FILLER_9_220 ();
 sg13g2_fill_1 FILLER_9_222 ();
 sg13g2_decap_4 FILLER_9_226 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_fill_1 FILLER_9_243 ();
 sg13g2_decap_8 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_254 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_decap_8 FILLER_9_268 ();
 sg13g2_decap_8 FILLER_9_275 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_decap_8 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_303 ();
 sg13g2_decap_8 FILLER_9_310 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_4 FILLER_10_119 ();
 sg13g2_fill_1 FILLER_10_123 ();
 sg13g2_fill_1 FILLER_10_181 ();
 sg13g2_decap_8 FILLER_10_188 ();
 sg13g2_decap_8 FILLER_10_195 ();
 sg13g2_decap_8 FILLER_10_202 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_fill_2 FILLER_10_273 ();
 sg13g2_fill_1 FILLER_10_278 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_296 ();
 sg13g2_decap_8 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_126 ();
 sg13g2_fill_1 FILLER_11_128 ();
 sg13g2_decap_8 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_fill_2 FILLER_11_165 ();
 sg13g2_fill_2 FILLER_11_170 ();
 sg13g2_fill_2 FILLER_11_178 ();
 sg13g2_fill_1 FILLER_11_180 ();
 sg13g2_decap_8 FILLER_11_184 ();
 sg13g2_decap_4 FILLER_11_191 ();
 sg13g2_fill_1 FILLER_11_195 ();
 sg13g2_decap_8 FILLER_11_211 ();
 sg13g2_decap_4 FILLER_11_218 ();
 sg13g2_fill_1 FILLER_11_222 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_fill_2 FILLER_11_249 ();
 sg13g2_fill_1 FILLER_11_254 ();
 sg13g2_fill_1 FILLER_11_258 ();
 sg13g2_fill_2 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_fill_2 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_128 ();
 sg13g2_fill_2 FILLER_12_156 ();
 sg13g2_decap_8 FILLER_12_209 ();
 sg13g2_fill_2 FILLER_12_228 ();
 sg13g2_decap_4 FILLER_12_233 ();
 sg13g2_fill_2 FILLER_12_237 ();
 sg13g2_fill_2 FILLER_12_251 ();
 sg13g2_fill_1 FILLER_12_253 ();
 sg13g2_decap_8 FILLER_12_257 ();
 sg13g2_fill_2 FILLER_12_264 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_fill_1 FILLER_12_282 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_324 ();
 sg13g2_decap_8 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_338 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_4 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_159 ();
 sg13g2_fill_1 FILLER_13_181 ();
 sg13g2_decap_8 FILLER_13_188 ();
 sg13g2_decap_8 FILLER_13_195 ();
 sg13g2_decap_8 FILLER_13_202 ();
 sg13g2_decap_8 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_216 ();
 sg13g2_fill_1 FILLER_13_218 ();
 sg13g2_decap_8 FILLER_13_285 ();
 sg13g2_fill_2 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_318 ();
 sg13g2_decap_8 FILLER_13_325 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_decap_8 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_decap_8 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_4 FILLER_14_133 ();
 sg13g2_fill_2 FILLER_14_137 ();
 sg13g2_decap_4 FILLER_14_160 ();
 sg13g2_decap_8 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_216 ();
 sg13g2_decap_8 FILLER_14_223 ();
 sg13g2_decap_8 FILLER_14_230 ();
 sg13g2_decap_8 FILLER_14_237 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_258 ();
 sg13g2_fill_2 FILLER_14_265 ();
 sg13g2_fill_1 FILLER_14_267 ();
 sg13g2_decap_8 FILLER_14_283 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_fill_1 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_4 FILLER_15_105 ();
 sg13g2_fill_1 FILLER_15_109 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_decap_8 FILLER_15_135 ();
 sg13g2_fill_1 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_4 FILLER_15_189 ();
 sg13g2_fill_2 FILLER_15_193 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_4 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_4 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_292 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_4 FILLER_16_98 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_fill_1 FILLER_16_122 ();
 sg13g2_decap_8 FILLER_16_144 ();
 sg13g2_decap_4 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_decap_8 FILLER_16_177 ();
 sg13g2_decap_4 FILLER_16_184 ();
 sg13g2_fill_2 FILLER_16_188 ();
 sg13g2_decap_8 FILLER_16_208 ();
 sg13g2_decap_8 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_222 ();
 sg13g2_fill_2 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_240 ();
 sg13g2_fill_1 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_306 ();
 sg13g2_decap_8 FILLER_16_313 ();
 sg13g2_decap_8 FILLER_16_320 ();
 sg13g2_decap_8 FILLER_16_327 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_355 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_fill_2 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_118 ();
 sg13g2_fill_2 FILLER_17_125 ();
 sg13g2_fill_1 FILLER_17_127 ();
 sg13g2_decap_4 FILLER_17_146 ();
 sg13g2_decap_8 FILLER_17_153 ();
 sg13g2_fill_2 FILLER_17_160 ();
 sg13g2_decap_4 FILLER_17_180 ();
 sg13g2_fill_2 FILLER_17_184 ();
 sg13g2_decap_8 FILLER_17_204 ();
 sg13g2_fill_2 FILLER_17_211 ();
 sg13g2_fill_1 FILLER_17_213 ();
 sg13g2_decap_8 FILLER_17_274 ();
 sg13g2_decap_8 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_288 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_4 FILLER_18_98 ();
 sg13g2_fill_2 FILLER_18_102 ();
 sg13g2_decap_4 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_decap_4 FILLER_18_175 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_4 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_decap_8 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_decap_4 FILLER_18_251 ();
 sg13g2_fill_2 FILLER_18_255 ();
 sg13g2_decap_8 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_288 ();
 sg13g2_decap_8 FILLER_18_295 ();
 sg13g2_decap_8 FILLER_18_302 ();
 sg13g2_decap_8 FILLER_18_309 ();
 sg13g2_decap_8 FILLER_18_316 ();
 sg13g2_decap_8 FILLER_18_323 ();
 sg13g2_decap_8 FILLER_18_330 ();
 sg13g2_decap_8 FILLER_18_337 ();
 sg13g2_decap_8 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_18_372 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_4 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_122 ();
 sg13g2_decap_4 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_146 ();
 sg13g2_decap_8 FILLER_19_150 ();
 sg13g2_decap_8 FILLER_19_157 ();
 sg13g2_decap_8 FILLER_19_164 ();
 sg13g2_decap_8 FILLER_19_171 ();
 sg13g2_fill_2 FILLER_19_178 ();
 sg13g2_decap_8 FILLER_19_195 ();
 sg13g2_fill_2 FILLER_19_202 ();
 sg13g2_decap_8 FILLER_19_219 ();
 sg13g2_decap_8 FILLER_19_226 ();
 sg13g2_fill_1 FILLER_19_236 ();
 sg13g2_fill_1 FILLER_19_240 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_250 ();
 sg13g2_decap_4 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_4 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_78 ();
 sg13g2_decap_8 FILLER_20_85 ();
 sg13g2_fill_2 FILLER_20_92 ();
 sg13g2_fill_1 FILLER_20_94 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_fill_2 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_122 ();
 sg13g2_fill_1 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_fill_2 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_4 FILLER_20_217 ();
 sg13g2_decap_4 FILLER_20_257 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_decap_8 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_285 ();
 sg13g2_fill_2 FILLER_20_292 ();
 sg13g2_fill_1 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_4 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_63 ();
 sg13g2_decap_4 FILLER_21_115 ();
 sg13g2_fill_1 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_135 ();
 sg13g2_fill_1 FILLER_21_142 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_decap_4 FILLER_21_173 ();
 sg13g2_decap_4 FILLER_21_180 ();
 sg13g2_fill_2 FILLER_21_184 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_decap_4 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_232 ();
 sg13g2_fill_2 FILLER_21_239 ();
 sg13g2_fill_1 FILLER_21_241 ();
 sg13g2_decap_8 FILLER_21_257 ();
 sg13g2_decap_4 FILLER_21_264 ();
 sg13g2_fill_2 FILLER_21_268 ();
 sg13g2_decap_8 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_4 FILLER_21_351 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_63 ();
 sg13g2_decap_4 FILLER_22_79 ();
 sg13g2_fill_1 FILLER_22_83 ();
 sg13g2_fill_1 FILLER_22_87 ();
 sg13g2_fill_1 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_fill_1 FILLER_22_118 ();
 sg13g2_decap_8 FILLER_22_131 ();
 sg13g2_decap_4 FILLER_22_138 ();
 sg13g2_fill_2 FILLER_22_157 ();
 sg13g2_fill_1 FILLER_22_159 ();
 sg13g2_decap_8 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_227 ();
 sg13g2_fill_1 FILLER_22_229 ();
 sg13g2_fill_2 FILLER_22_233 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_4 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_fill_1 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_fill_2 FILLER_22_381 ();
 sg13g2_fill_1 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_4 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_83 ();
 sg13g2_decap_8 FILLER_23_90 ();
 sg13g2_decap_8 FILLER_23_97 ();
 sg13g2_decap_4 FILLER_23_104 ();
 sg13g2_fill_1 FILLER_23_117 ();
 sg13g2_fill_2 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_fill_1 FILLER_23_158 ();
 sg13g2_decap_8 FILLER_23_177 ();
 sg13g2_decap_8 FILLER_23_184 ();
 sg13g2_decap_4 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_195 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_4 FILLER_23_221 ();
 sg13g2_fill_2 FILLER_23_243 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_260 ();
 sg13g2_fill_2 FILLER_23_267 ();
 sg13g2_decap_4 FILLER_23_272 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_281 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_decap_4 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_291 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_decap_4 FILLER_23_380 ();
 sg13g2_fill_2 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_4 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_95 ();
 sg13g2_decap_4 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_124 ();
 sg13g2_fill_2 FILLER_24_131 ();
 sg13g2_fill_1 FILLER_24_133 ();
 sg13g2_decap_4 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_153 ();
 sg13g2_decap_8 FILLER_24_173 ();
 sg13g2_decap_4 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_4 FILLER_24_214 ();
 sg13g2_fill_1 FILLER_24_218 ();
 sg13g2_decap_8 FILLER_24_237 ();
 sg13g2_decap_4 FILLER_24_244 ();
 sg13g2_fill_1 FILLER_24_248 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_decap_4 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_fill_2 FILLER_25_77 ();
 sg13g2_fill_1 FILLER_25_79 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_127 ();
 sg13g2_fill_2 FILLER_25_134 ();
 sg13g2_fill_2 FILLER_25_151 ();
 sg13g2_decap_4 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_169 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_247 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_decap_8 FILLER_25_269 ();
 sg13g2_decap_8 FILLER_25_276 ();
 sg13g2_decap_4 FILLER_25_283 ();
 sg13g2_fill_1 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_291 ();
 sg13g2_fill_1 FILLER_25_298 ();
 sg13g2_decap_4 FILLER_25_305 ();
 sg13g2_decap_4 FILLER_25_336 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_fill_1 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_11 ();
 sg13g2_decap_4 FILLER_26_16 ();
 sg13g2_fill_1 FILLER_26_20 ();
 sg13g2_decap_8 FILLER_26_24 ();
 sg13g2_decap_8 FILLER_26_31 ();
 sg13g2_decap_4 FILLER_26_38 ();
 sg13g2_decap_8 FILLER_26_69 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_78 ();
 sg13g2_decap_8 FILLER_26_100 ();
 sg13g2_decap_4 FILLER_26_107 ();
 sg13g2_decap_8 FILLER_26_129 ();
 sg13g2_decap_4 FILLER_26_136 ();
 sg13g2_fill_1 FILLER_26_140 ();
 sg13g2_fill_1 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_fill_2 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_169 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_4 FILLER_26_195 ();
 sg13g2_fill_2 FILLER_26_199 ();
 sg13g2_decap_4 FILLER_26_219 ();
 sg13g2_fill_1 FILLER_26_223 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_fill_2 FILLER_26_249 ();
 sg13g2_fill_1 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_decap_4 FILLER_26_274 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_4 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_338 ();
 sg13g2_decap_4 FILLER_26_345 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_fill_1 FILLER_26_373 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_40 ();
 sg13g2_decap_4 FILLER_27_50 ();
 sg13g2_fill_2 FILLER_27_54 ();
 sg13g2_fill_2 FILLER_27_74 ();
 sg13g2_fill_1 FILLER_27_76 ();
 sg13g2_decap_8 FILLER_27_95 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_fill_1 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_165 ();
 sg13g2_fill_2 FILLER_27_172 ();
 sg13g2_decap_8 FILLER_27_195 ();
 sg13g2_fill_2 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_decap_4 FILLER_27_220 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_decap_4 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_decap_8 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_274 ();
 sg13g2_fill_2 FILLER_27_291 ();
 sg13g2_fill_1 FILLER_27_293 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_323 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_decap_8 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_59 ();
 sg13g2_decap_8 FILLER_28_66 ();
 sg13g2_decap_4 FILLER_28_73 ();
 sg13g2_decap_8 FILLER_28_95 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_125 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_decap_8 FILLER_28_148 ();
 sg13g2_fill_2 FILLER_28_155 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_fill_1 FILLER_28_176 ();
 sg13g2_decap_8 FILLER_28_192 ();
 sg13g2_decap_8 FILLER_28_199 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_243 ();
 sg13g2_fill_2 FILLER_28_250 ();
 sg13g2_fill_1 FILLER_28_252 ();
 sg13g2_decap_4 FILLER_28_268 ();
 sg13g2_fill_2 FILLER_28_272 ();
 sg13g2_decap_8 FILLER_28_292 ();
 sg13g2_decap_4 FILLER_28_299 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_decap_8 FILLER_28_320 ();
 sg13g2_decap_8 FILLER_28_327 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_fill_2 FILLER_28_361 ();
 sg13g2_fill_1 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_fill_1 FILLER_29_44 ();
 sg13g2_fill_2 FILLER_29_66 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_fill_1 FILLER_29_81 ();
 sg13g2_fill_1 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_4 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_146 ();
 sg13g2_fill_1 FILLER_29_153 ();
 sg13g2_fill_2 FILLER_29_172 ();
 sg13g2_fill_1 FILLER_29_174 ();
 sg13g2_decap_8 FILLER_29_190 ();
 sg13g2_decap_8 FILLER_29_197 ();
 sg13g2_decap_8 FILLER_29_204 ();
 sg13g2_decap_4 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_230 ();
 sg13g2_decap_4 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_288 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_fill_2 FILLER_29_347 ();
 sg13g2_fill_1 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_4 FILLER_29_363 ();
 sg13g2_decap_4 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_31 ();
 sg13g2_decap_8 FILLER_30_41 ();
 sg13g2_decap_4 FILLER_30_48 ();
 sg13g2_fill_1 FILLER_30_52 ();
 sg13g2_decap_4 FILLER_30_62 ();
 sg13g2_fill_1 FILLER_30_66 ();
 sg13g2_fill_2 FILLER_30_85 ();
 sg13g2_decap_8 FILLER_30_90 ();
 sg13g2_decap_8 FILLER_30_97 ();
 sg13g2_decap_8 FILLER_30_104 ();
 sg13g2_decap_8 FILLER_30_111 ();
 sg13g2_decap_8 FILLER_30_118 ();
 sg13g2_decap_8 FILLER_30_143 ();
 sg13g2_decap_8 FILLER_30_150 ();
 sg13g2_decap_4 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_fill_2 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_199 ();
 sg13g2_decap_8 FILLER_30_206 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_fill_2 FILLER_30_223 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_fill_1 FILLER_30_240 ();
 sg13g2_decap_8 FILLER_30_262 ();
 sg13g2_fill_1 FILLER_30_269 ();
 sg13g2_decap_8 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_4 FILLER_30_319 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_decap_8 FILLER_30_363 ();
 sg13g2_decap_4 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_23 ();
 sg13g2_decap_8 FILLER_31_30 ();
 sg13g2_decap_8 FILLER_31_37 ();
 sg13g2_decap_8 FILLER_31_44 ();
 sg13g2_decap_4 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_decap_8 FILLER_31_89 ();
 sg13g2_decap_8 FILLER_31_96 ();
 sg13g2_decap_8 FILLER_31_103 ();
 sg13g2_decap_8 FILLER_31_110 ();
 sg13g2_decap_8 FILLER_31_117 ();
 sg13g2_decap_8 FILLER_31_142 ();
 sg13g2_decap_8 FILLER_31_149 ();
 sg13g2_decap_8 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_163 ();
 sg13g2_decap_8 FILLER_31_185 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_225 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_decap_4 FILLER_31_242 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_fill_2 FILLER_31_273 ();
 sg13g2_fill_1 FILLER_31_290 ();
 sg13g2_decap_8 FILLER_31_297 ();
 sg13g2_decap_4 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_308 ();
 sg13g2_fill_2 FILLER_31_330 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_decap_8 FILLER_31_339 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_1 FILLER_31_368 ();
 sg13g2_decap_4 FILLER_31_372 ();
 sg13g2_fill_2 FILLER_31_376 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_decap_4 FILLER_32_20 ();
 sg13g2_fill_2 FILLER_32_24 ();
 sg13g2_decap_8 FILLER_32_44 ();
 sg13g2_decap_4 FILLER_32_51 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_82 ();
 sg13g2_decap_8 FILLER_32_89 ();
 sg13g2_decap_8 FILLER_32_96 ();
 sg13g2_decap_8 FILLER_32_103 ();
 sg13g2_decap_8 FILLER_32_110 ();
 sg13g2_decap_8 FILLER_32_117 ();
 sg13g2_fill_2 FILLER_32_124 ();
 sg13g2_fill_1 FILLER_32_126 ();
 sg13g2_fill_1 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_4 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_271 ();
 sg13g2_decap_4 FILLER_32_295 ();
 sg13g2_decap_8 FILLER_32_317 ();
 sg13g2_fill_2 FILLER_32_324 ();
 sg13g2_decap_4 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_29 ();
 sg13g2_decap_4 FILLER_33_36 ();
 sg13g2_fill_1 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_110 ();
 sg13g2_fill_2 FILLER_33_114 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_123 ();
 sg13g2_fill_2 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_137 ();
 sg13g2_decap_4 FILLER_33_144 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_decap_8 FILLER_33_165 ();
 sg13g2_fill_2 FILLER_33_172 ();
 sg13g2_fill_1 FILLER_33_174 ();
 sg13g2_decap_8 FILLER_33_178 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_fill_1 FILLER_33_209 ();
 sg13g2_decap_8 FILLER_33_216 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_235 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_decap_4 FILLER_33_254 ();
 sg13g2_decap_4 FILLER_33_270 ();
 sg13g2_fill_2 FILLER_33_274 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_296 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_decap_4 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_363 ();
 sg13g2_decap_8 FILLER_33_370 ();
 sg13g2_decap_4 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_15 ();
 sg13g2_fill_2 FILLER_34_19 ();
 sg13g2_fill_1 FILLER_34_24 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_4 FILLER_34_35 ();
 sg13g2_fill_2 FILLER_34_39 ();
 sg13g2_decap_8 FILLER_34_53 ();
 sg13g2_fill_1 FILLER_34_60 ();
 sg13g2_fill_1 FILLER_34_73 ();
 sg13g2_decap_8 FILLER_34_80 ();
 sg13g2_decap_4 FILLER_34_87 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_decap_4 FILLER_34_159 ();
 sg13g2_decap_8 FILLER_34_169 ();
 sg13g2_decap_4 FILLER_34_176 ();
 sg13g2_fill_2 FILLER_34_180 ();
 sg13g2_decap_8 FILLER_34_188 ();
 sg13g2_decap_8 FILLER_34_199 ();
 sg13g2_decap_4 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_210 ();
 sg13g2_fill_2 FILLER_34_251 ();
 sg13g2_decap_8 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_2 FILLER_35_51 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_86 ();
 sg13g2_decap_8 FILLER_35_93 ();
 sg13g2_fill_1 FILLER_35_100 ();
 sg13g2_decap_8 FILLER_35_110 ();
 sg13g2_decap_8 FILLER_35_117 ();
 sg13g2_decap_8 FILLER_35_124 ();
 sg13g2_decap_8 FILLER_35_131 ();
 sg13g2_decap_8 FILLER_35_138 ();
 sg13g2_decap_8 FILLER_35_145 ();
 sg13g2_decap_4 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_156 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_decap_8 FILLER_35_235 ();
 sg13g2_decap_4 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_decap_8 FILLER_35_251 ();
 sg13g2_decap_8 FILLER_35_258 ();
 sg13g2_decap_8 FILLER_35_269 ();
 sg13g2_fill_1 FILLER_35_276 ();
 sg13g2_decap_8 FILLER_35_286 ();
 sg13g2_decap_8 FILLER_35_293 ();
 sg13g2_decap_8 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_decap_8 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_384 ();
 sg13g2_decap_8 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_20 ();
 sg13g2_fill_1 FILLER_36_22 ();
 sg13g2_decap_4 FILLER_36_26 ();
 sg13g2_fill_2 FILLER_36_30 ();
 sg13g2_fill_2 FILLER_36_38 ();
 sg13g2_fill_1 FILLER_36_40 ();
 sg13g2_fill_2 FILLER_36_44 ();
 sg13g2_fill_1 FILLER_36_46 ();
 sg13g2_decap_8 FILLER_36_74 ();
 sg13g2_decap_4 FILLER_36_81 ();
 sg13g2_fill_2 FILLER_36_85 ();
 sg13g2_decap_4 FILLER_36_108 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_fill_2 FILLER_36_125 ();
 sg13g2_fill_1 FILLER_36_127 ();
 sg13g2_decap_8 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_138 ();
 sg13g2_decap_8 FILLER_36_145 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_179 ();
 sg13g2_decap_8 FILLER_36_186 ();
 sg13g2_decap_4 FILLER_36_193 ();
 sg13g2_fill_2 FILLER_36_197 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_fill_2 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_decap_8 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_4 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_11 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_decap_8 FILLER_37_58 ();
 sg13g2_decap_8 FILLER_37_65 ();
 sg13g2_decap_8 FILLER_37_72 ();
 sg13g2_decap_8 FILLER_37_79 ();
 sg13g2_fill_1 FILLER_37_86 ();
 sg13g2_fill_1 FILLER_37_99 ();
 sg13g2_fill_1 FILLER_37_103 ();
 sg13g2_fill_1 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_150 ();
 sg13g2_fill_1 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_170 ();
 sg13g2_decap_8 FILLER_37_177 ();
 sg13g2_decap_4 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_188 ();
 sg13g2_fill_1 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_37_391 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_4 ();
 sg13g2_fill_1 FILLER_38_12 ();
 sg13g2_fill_1 FILLER_38_16 ();
 sg13g2_fill_1 FILLER_38_20 ();
 sg13g2_decap_8 FILLER_38_24 ();
 sg13g2_decap_8 FILLER_38_31 ();
 sg13g2_decap_8 FILLER_38_38 ();
 sg13g2_decap_8 FILLER_38_45 ();
 sg13g2_decap_4 FILLER_38_52 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_100 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_167 ();
 sg13g2_decap_8 FILLER_38_174 ();
 sg13g2_fill_2 FILLER_38_181 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_decap_8 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_195 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_4 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_245 ();
 sg13g2_fill_1 FILLER_38_247 ();
 sg13g2_decap_4 FILLER_38_252 ();
 sg13g2_decap_4 FILLER_38_268 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_decap_4 FILLER_38_301 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_4 FILLER_38_387 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net42;
 assign uio_oe[1] = net43;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net44;
 assign uio_oe[7] = net45;
 assign uio_out[2] = net23;
 assign uio_out[3] = net24;
 assign uio_out[4] = net25;
 assign uio_out[5] = net26;
 assign uo_out[7] = net27;
endmodule

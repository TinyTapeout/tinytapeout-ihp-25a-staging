module tt_um_wokwi_group_7 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire net11;
 wire net12;
 wire net13;
 wire \proj_10.net4 ;
 wire \proj_10.net5 ;
 wire \proj_10.net6 ;
 wire \proj_10.net7 ;
 wire \proj_11.net10 ;
 wire \proj_11.net11 ;
 wire \proj_11.net17 ;
 wire \proj_11.net18 ;
 wire \proj_11.net19 ;
 wire \proj_11.net20 ;
 wire \proj_11.net21 ;
 wire \proj_11.net6 ;
 wire \proj_11.net7 ;
 wire \proj_11.net8 ;
 wire \proj_11.net9 ;
 wire \proj_12.net14 ;
 wire \proj_12.net4 ;
 wire \proj_12.net5 ;
 wire \proj_12.net6 ;
 wire \proj_12.net7 ;
 wire \proj_12.net8 ;
 wire \proj_13.net11 ;
 wire \proj_13.net12 ;
 wire \proj_13.net13 ;
 wire \proj_13.net4 ;
 wire \proj_13.net5 ;
 wire \proj_14.net6 ;
 wire \proj_14.net7 ;
 wire \proj_14.net8 ;
 wire \proj__0.net10 ;
 wire \proj__0.net11 ;
 wire \proj__0.net12 ;
 wire \proj__0.net13 ;
 wire \proj__0.net19 ;
 wire \proj__0.net20 ;
 wire \proj__0.net21 ;
 wire \proj__0.net22 ;
 wire \proj__0.net23 ;
 wire \proj__0.net24 ;
 wire \proj__0.net25 ;
 wire \proj__0.net26 ;
 wire \proj__0.net27 ;
 wire \proj__0.net28 ;
 wire \proj__0.net29 ;
 wire \proj__0.net30 ;
 wire \proj__0.net31 ;
 wire \proj__0.net32 ;
 wire \proj__0.net33 ;
 wire \proj__0.net34 ;
 wire \proj__0.net35 ;
 wire \proj__0.net36 ;
 wire \proj__0.net9 ;
 wire \proj__1.net7 ;
 wire \proj__2.net10 ;
 wire \proj__2.net11 ;
 wire \proj__2.net17 ;
 wire \proj__2.net18 ;
 wire \proj__2.net19 ;
 wire \proj__2.net20 ;
 wire \proj__2.net21 ;
 wire \proj__2.net22 ;
 wire \proj__2.net23 ;
 wire \proj__2.net24 ;
 wire \proj__2.net25 ;
 wire \proj__2.net26 ;
 wire \proj__2.net27 ;
 wire \proj__2.net28 ;
 wire \proj__2.net29 ;
 wire \proj__2.net30 ;
 wire \proj__2.net31 ;
 wire \proj__2.net32 ;
 wire \proj__2.net33 ;
 wire \proj__2.net34 ;
 wire \proj__2.net35 ;
 wire \proj__2.net36 ;
 wire \proj__2.net37 ;
 wire \proj__2.net38 ;
 wire \proj__2.net39 ;
 wire \proj__2.net40 ;
 wire \proj__2.net41 ;
 wire \proj__2.net42 ;
 wire \proj__2.net43 ;
 wire \proj__2.net44 ;
 wire \proj__2.net45 ;
 wire \proj__2.net46 ;
 wire \proj__2.net47 ;
 wire \proj__2.net48 ;
 wire \proj__2.net49 ;
 wire \proj__2.net5 ;
 wire \proj__2.net50 ;
 wire \proj__2.net51 ;
 wire \proj__2.net52 ;
 wire \proj__2.net53 ;
 wire \proj__2.net54 ;
 wire \proj__2.net55 ;
 wire \proj__2.net56 ;
 wire \proj__2.net57 ;
 wire \proj__2.net58 ;
 wire \proj__2.net59 ;
 wire \proj__2.net6 ;
 wire \proj__2.net60 ;
 wire \proj__2.net61 ;
 wire \proj__2.net62 ;
 wire \proj__2.net63 ;
 wire \proj__2.net64 ;
 wire \proj__2.net65 ;
 wire \proj__2.net66 ;
 wire \proj__2.net67 ;
 wire \proj__2.net68 ;
 wire \proj__2.net69 ;
 wire \proj__2.net7 ;
 wire \proj__2.net70 ;
 wire \proj__2.net71 ;
 wire \proj__2.net72 ;
 wire \proj__2.net73 ;
 wire \proj__2.net74 ;
 wire \proj__2.net75 ;
 wire \proj__2.net76 ;
 wire \proj__2.net77 ;
 wire \proj__2.net78 ;
 wire \proj__2.net79 ;
 wire \proj__2.net8 ;
 wire \proj__2.net80 ;
 wire \proj__2.net81 ;
 wire \proj__2.net82 ;
 wire \proj__2.net83 ;
 wire \proj__2.net84 ;
 wire \proj__2.net85 ;
 wire \proj__2.net86 ;
 wire \proj__2.net87 ;
 wire \proj__2.net9 ;
 wire \proj__3.net10 ;
 wire \proj__3.net11 ;
 wire \proj__3.net12 ;
 wire \proj__3.net18 ;
 wire \proj__3.net19 ;
 wire \proj__3.net20 ;
 wire \proj__3.net21 ;
 wire \proj__3.net9 ;
 wire \proj__4.net10 ;
 wire \proj__4.net11 ;
 wire \proj__4.net12 ;
 wire \proj__4.net9 ;
 wire \proj__5.net7 ;
 wire \proj__5.net8 ;
 wire \proj__5.net9 ;
 wire \proj__6.net10 ;
 wire \proj__6.net9 ;
 wire \proj__7.net10 ;
 wire \proj__7.net11 ;
 wire \proj__7.net12 ;
 wire \proj__7.net13 ;
 wire \proj__7.net14 ;
 wire \proj__7.net15 ;
 wire \proj__7.net21 ;
 wire \proj__7.net22 ;
 wire \proj__7.net23 ;
 wire \proj__7.net24 ;
 wire \proj__7.net25 ;
 wire \proj__7.net26 ;
 wire \proj__7.net27 ;
 wire \proj__7.net28 ;
 wire \proj__7.net9 ;
 wire \proj__8.net10 ;
 wire \proj__8.net11 ;
 wire \proj__8.net12 ;
 wire \proj__8.net4 ;
 wire \proj__8.net5 ;
 wire \proj__9.net10 ;
 wire \proj__9.net11 ;
 wire \proj__9.net12 ;
 wire \proj__9.net9 ;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire \proj_11.flop1/notq ;
 wire net33;
 wire \proj_11.flop2/notq ;
 wire net34;
 wire \proj_11.flop5/notq ;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;

 sg13g2_inv_1 _074_ (.Y(_048_),
    .A(\proj__0.net10 ));
 sg13g2_inv_1 _075_ (.Y(_049_),
    .A(\proj__0.net11 ));
 sg13g2_inv_1 _076_ (.Y(_050_),
    .A(\proj__0.net12 ));
 sg13g2_nor2_2 _077_ (.A(net7),
    .B(net6),
    .Y(_051_));
 sg13g2_nor2b_2 _078_ (.A(net9),
    .B_N(net8),
    .Y(_052_));
 sg13g2_and2_2 _079_ (.A(_051_),
    .B(_052_),
    .X(_053_));
 sg13g2_and2_1 _080_ (.A(net7),
    .B(net6),
    .X(_054_));
 sg13g2_and2_2 _081_ (.A(_052_),
    .B(_054_),
    .X(_055_));
 sg13g2_nor2b_2 _082_ (.A(net6),
    .B_N(net7),
    .Y(_056_));
 sg13g2_nor2_1 _083_ (.A(net9),
    .B(net8),
    .Y(_057_));
 sg13g2_and2_2 _084_ (.A(_056_),
    .B(_057_),
    .X(_058_));
 sg13g2_and3_2 _085_ (.X(_059_),
    .A(net9),
    .B(net8),
    .C(_051_));
 sg13g2_nor2b_1 _086_ (.A(net8),
    .B_N(net9),
    .Y(_060_));
 sg13g2_and2_1 _087_ (.A(_056_),
    .B(_060_),
    .X(_061_));
 sg13g2_and2_1 _088_ (.A(_051_),
    .B(_060_),
    .X(_062_));
 sg13g2_and2_1 _089_ (.A(_052_),
    .B(_056_),
    .X(_063_));
 sg13g2_nor2b_2 _090_ (.A(net7),
    .B_N(net6),
    .Y(_064_));
 sg13g2_and3_1 _091_ (.X(_065_),
    .A(net9),
    .B(net8),
    .C(_064_));
 sg13g2_nand2_1 _092_ (.Y(_066_),
    .A(\proj_13.net4 ),
    .B(_065_));
 sg13g2_and2_2 _093_ (.A(_054_),
    .B(_060_),
    .X(_067_));
 sg13g2_and2_2 _094_ (.A(_060_),
    .B(_064_),
    .X(_068_));
 sg13g2_and2_1 _095_ (.A(_051_),
    .B(_057_),
    .X(_069_));
 sg13g2_nand3_1 _096_ (.B(_057_),
    .C(_064_),
    .A(\proj__1.net7 ),
    .Y(_070_));
 sg13g2_a22oi_1 _097_ (.Y(_000_),
    .B1(net71),
    .B2(\proj__0.net9 ),
    .A2(_063_),
    .A1(\proj__6.net9 ));
 sg13g2_a22oi_1 _098_ (.Y(_001_),
    .B1(_067_),
    .B2(\proj_11.net6 ),
    .A2(_061_),
    .A1(\proj_10.net4 ));
 sg13g2_a22oi_1 _099_ (.Y(_002_),
    .B1(_058_),
    .B2(\proj__2.net5 ),
    .A2(_053_),
    .A1(\proj__4.net9 ));
 sg13g2_a22oi_1 _100_ (.Y(_003_),
    .B1(_062_),
    .B2(\proj__8.net4 ),
    .A2(_059_),
    .A1(\proj_12.net4 ));
 sg13g2_and4_1 _101_ (.A(_000_),
    .B(_001_),
    .C(_002_),
    .D(_003_),
    .X(_004_));
 sg13g2_a22oi_1 _102_ (.Y(_005_),
    .B1(_068_),
    .B2(\proj__9.net9 ),
    .A2(_055_),
    .A1(\proj__7.net9 ));
 sg13g2_nand4_1 _103_ (.B(_070_),
    .C(_004_),
    .A(_066_),
    .Y(uo_out[0]),
    .D(_005_));
 sg13g2_and3_1 _104_ (.X(_006_),
    .A(net9),
    .B(net8),
    .C(_056_));
 sg13g2_a21oi_1 _105_ (.A1(\proj_14.net6 ),
    .A2(_006_),
    .Y(_007_),
    .B1(net71));
 sg13g2_a22oi_1 _106_ (.Y(_008_),
    .B1(_067_),
    .B2(\proj_11.net7 ),
    .A2(_065_),
    .A1(\proj_13.net5 ));
 sg13g2_a22oi_1 _107_ (.Y(_009_),
    .B1(_062_),
    .B2(\proj__8.net5 ),
    .A2(_059_),
    .A1(\proj_12.net5 ));
 sg13g2_and2_1 _108_ (.A(_052_),
    .B(_064_),
    .X(_010_));
 sg13g2_a22oi_1 _109_ (.Y(_011_),
    .B1(_010_),
    .B2(\proj__5.net7 ),
    .A2(_063_),
    .A1(\proj__6.net10 ));
 sg13g2_a22oi_1 _110_ (.Y(_012_),
    .B1(_068_),
    .B2(\proj__9.net10 ),
    .A2(_061_),
    .A1(\proj_10.net5 ));
 sg13g2_a22oi_1 _111_ (.Y(_013_),
    .B1(_055_),
    .B2(\proj__7.net10 ),
    .A2(_053_),
    .A1(\proj__4.net10 ));
 sg13g2_and2_2 _112_ (.A(_054_),
    .B(_057_),
    .X(_014_));
 sg13g2_a22oi_1 _113_ (.Y(_015_),
    .B1(_014_),
    .B2(\proj__3.net9 ),
    .A2(_058_),
    .A1(\proj__2.net6 ));
 sg13g2_and4_1 _114_ (.A(_007_),
    .B(_008_),
    .C(_009_),
    .D(_015_),
    .X(_016_));
 sg13g2_and3_1 _115_ (.X(_017_),
    .A(_011_),
    .B(_012_),
    .C(_013_));
 sg13g2_a22oi_1 _116_ (.Y(uo_out[1]),
    .B1(_016_),
    .B2(_017_),
    .A2(net71),
    .A1(_048_));
 sg13g2_a22oi_1 _117_ (.Y(_018_),
    .B1(_067_),
    .B2(\proj_11.net8 ),
    .A2(_061_),
    .A1(\proj_10.net6 ));
 sg13g2_a22oi_1 _118_ (.Y(_019_),
    .B1(_014_),
    .B2(\proj__3.net10 ),
    .A2(_053_),
    .A1(\proj__4.net11 ));
 sg13g2_a22oi_1 _119_ (.Y(_020_),
    .B1(_068_),
    .B2(\proj__9.net11 ),
    .A2(_059_),
    .A1(\proj_12.net6 ));
 sg13g2_and2_1 _120_ (.A(_019_),
    .B(_020_),
    .X(_021_));
 sg13g2_a22oi_1 _121_ (.Y(_022_),
    .B1(_058_),
    .B2(\proj__2.net7 ),
    .A2(_055_),
    .A1(\proj__7.net11 ));
 sg13g2_and3_1 _122_ (.X(_023_),
    .A(_007_),
    .B(_018_),
    .C(_022_));
 sg13g2_a22oi_1 _123_ (.Y(uo_out[2]),
    .B1(_021_),
    .B2(_023_),
    .A2(net71),
    .A1(_049_));
 sg13g2_nand2_1 _124_ (.Y(_024_),
    .A(\proj_11.net9 ),
    .B(_067_));
 sg13g2_a22oi_1 _125_ (.Y(_025_),
    .B1(_063_),
    .B2(net3),
    .A2(_059_),
    .A1(\proj_12.net7 ));
 sg13g2_nand2_1 _126_ (.Y(_026_),
    .A(\proj_10.net7 ),
    .B(_061_));
 sg13g2_a21o_1 _127_ (.A2(_068_),
    .A1(\proj__9.net12 ),
    .B1(net71),
    .X(_027_));
 sg13g2_a221oi_1 _128_ (.B2(\proj__3.net11 ),
    .C1(_027_),
    .B1(_014_),
    .A1(\proj__2.net8 ),
    .Y(_028_),
    .A2(_058_));
 sg13g2_a22oi_1 _129_ (.Y(_029_),
    .B1(_055_),
    .B2(\proj__7.net12 ),
    .A2(_053_),
    .A1(\proj__4.net12 ));
 sg13g2_and4_1 _130_ (.A(_024_),
    .B(_025_),
    .C(_026_),
    .D(_029_),
    .X(_030_));
 sg13g2_a22oi_1 _131_ (.Y(uo_out[3]),
    .B1(_028_),
    .B2(_030_),
    .A2(net71),
    .A1(_050_));
 sg13g2_nor2b_1 _132_ (.A(net8),
    .B_N(_064_),
    .Y(_031_));
 sg13g2_or3_1 _133_ (.A(_053_),
    .B(_063_),
    .C(_031_),
    .X(_032_));
 sg13g2_nand2_1 _134_ (.Y(_033_),
    .A(net2),
    .B(_032_));
 sg13g2_a22oi_1 _135_ (.Y(_034_),
    .B1(_014_),
    .B2(\proj__3.net12 ),
    .A2(_055_),
    .A1(\proj__7.net13 ));
 sg13g2_a22oi_1 _136_ (.Y(_035_),
    .B1(_059_),
    .B2(net86),
    .A2(_058_),
    .A1(\proj__2.net9 ));
 sg13g2_a22oi_1 _137_ (.Y(_036_),
    .B1(_069_),
    .B2(\proj__0.net13 ),
    .A2(_067_),
    .A1(\proj_11.net10 ));
 sg13g2_nand4_1 _138_ (.B(_034_),
    .C(_035_),
    .A(_033_),
    .Y(uo_out[4]),
    .D(_036_));
 sg13g2_and3_1 _139_ (.X(_037_),
    .A(\proj__5.net8 ),
    .B(_052_),
    .C(_064_));
 sg13g2_a221oi_1 _140_ (.B2(\proj__2.net10 ),
    .C1(_037_),
    .B1(_058_),
    .A1(\proj__7.net14 ),
    .Y(_038_),
    .A2(_055_));
 sg13g2_o21ai_1 _141_ (.B1(net3),
    .Y(_039_),
    .A1(_053_),
    .A2(_031_));
 sg13g2_a22oi_1 _142_ (.Y(_040_),
    .B1(net71),
    .B2(\proj__0.net13 ),
    .A2(_067_),
    .A1(\proj_11.net11 ));
 sg13g2_nand3_1 _143_ (.B(_039_),
    .C(_040_),
    .A(_038_),
    .Y(uo_out[5]));
 sg13g2_nand2_1 _144_ (.Y(_041_),
    .A(net4),
    .B(_032_));
 sg13g2_nand2_1 _145_ (.Y(_042_),
    .A(\proj__2.net11 ),
    .B(_058_));
 sg13g2_a22oi_1 _146_ (.Y(_043_),
    .B1(_059_),
    .B2(\proj_12.net8 ),
    .A2(_055_),
    .A1(\proj__7.net15 ));
 sg13g2_a22oi_1 _147_ (.Y(_044_),
    .B1(_006_),
    .B2(\proj_14.net7 ),
    .A2(net71),
    .A1(\proj__0.net9 ));
 sg13g2_nand4_1 _148_ (.B(_042_),
    .C(_043_),
    .A(_041_),
    .Y(uo_out[6]),
    .D(_044_));
 sg13g2_nand2_1 _149_ (.Y(_045_),
    .A(net5),
    .B(_032_));
 sg13g2_nand2_1 _150_ (.Y(_046_),
    .A(\proj_14.net8 ),
    .B(_006_));
 sg13g2_nand3_1 _151_ (.B(_052_),
    .C(_064_),
    .A(\proj__5.net9 ),
    .Y(_047_));
 sg13g2_nand3_1 _152_ (.B(_046_),
    .C(_047_),
    .A(_045_),
    .Y(uo_out[7]));
 sg13g2_tielo \proj_10.flop2/_1__11  (.L_LO(net11));
 sg13g2_tielo \proj_11.flop1/_1__12  (.L_LO(net12));
 sg13g2_tielo tt_um_wokwi_group_7_13 (.L_LO(net13));
 sg13g2_tielo tt_um_wokwi_group_7_14 (.L_LO(net14));
 sg13g2_tielo tt_um_wokwi_group_7_15 (.L_LO(net15));
 sg13g2_tielo tt_um_wokwi_group_7_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_group_7_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_group_7_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_group_7_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_group_7_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_group_7_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_group_7_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_group_7_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_group_7_24 (.L_LO(net24));
 sg13g2_tielo tt_um_wokwi_group_7_25 (.L_LO(net25));
 sg13g2_tielo tt_um_wokwi_group_7_26 (.L_LO(net26));
 sg13g2_tielo tt_um_wokwi_group_7_27 (.L_LO(net27));
 sg13g2_tielo tt_um_wokwi_group_7_28 (.L_LO(net28));
 sg13g2_tiehi \proj_10.flop1/_1__29  (.L_HI(net29));
 sg13g2_dfrbp_1 \proj_10.flop1/_1_  (.CLK(net10),
    .RESET_B(net29),
    .D(net88),
    .Q_N(\proj_10.net5 ),
    .Q(\proj_10.net4 ));
 sg13g2_tiehi \proj_10.flop2/_1__30  (.L_HI(net30));
 sg13g2_dfrbp_1 \proj_10.flop2/_1_  (.CLK(net11),
    .RESET_B(net30),
    .D(net79),
    .Q_N(\proj_10.net6 ),
    .Q(\proj_10.net7 ));
 sg13g2_tiehi \proj_11.flop1/_1__31  (.L_HI(net31));
 sg13g2_and2_1 \proj_11.and1/_0_  (.A(net78),
    .B(net82),
    .X(\proj_11.net11 ));
 sg13g2_dfrbp_1 \proj_11.flop1/_1_  (.CLK(net12),
    .RESET_B(net31),
    .D(\proj_11.net17 ),
    .Q_N(\proj_11.flop1/notq ),
    .Q(\proj_11.net9 ));
 sg13g2_tiehi \proj_11.flop2/_1__32  (.L_HI(net32));
 sg13g2_dfrbp_1 \proj_11.flop2/_1_  (.CLK(\proj_11.net8 ),
    .RESET_B(net32),
    .D(\proj_11.net19 ),
    .Q_N(\proj_11.flop2/notq ),
    .Q(\proj_11.net7 ));
 sg13g2_tiehi \proj_11.flop3/_1__33  (.L_HI(net33));
 sg13g2_dfrbp_1 \proj_11.flop3/_1_  (.CLK(\proj_11.net7 ),
    .RESET_B(net33),
    .D(\proj_11.net20 ),
    .Q_N(\proj_11.net6 ),
    .Q(\proj_11.net21 ));
 sg13g2_tiehi \proj_11.flop5/_1__34  (.L_HI(net34));
 sg13g2_dfrbp_1 \proj_11.flop5/_1_  (.CLK(\proj_11.net9 ),
    .RESET_B(net34),
    .D(\proj_11.net18 ),
    .Q_N(\proj_11.flop5/notq ),
    .Q(\proj_11.net8 ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_nand2_1 \proj_11.nand1/_0_  (.Y(\proj_11.net10 ),
    .A(net87),
    .B(net90));
 sg13g2_inv_1 \proj_11.not1/_0_  (.Y(\proj_11.net17 ),
    .A(\proj_11.net9 ));
 sg13g2_inv_1 \proj_11.not2/_0_  (.Y(\proj_11.net18 ),
    .A(\proj_11.net8 ));
 sg13g2_inv_1 \proj_11.not3/_0_  (.Y(\proj_11.net19 ),
    .A(\proj_11.net7 ));
 sg13g2_inv_1 \proj_11.not4/_0_  (.Y(\proj_11.net20 ),
    .A(\proj_11.net21 ));
 sg13g2_or2_1 \proj_12.or1/_0_  (.X(\proj_12.net14 ),
    .B(net88),
    .A(net83));
 sg13g2_or2_1 \proj_12.or2/_0_  (.X(\proj_12.net8 ),
    .B(net81),
    .A(net85));
 sg13g2_or2_1 \proj_12.or3/_0_  (.X(\proj_12.net6 ),
    .B(net88),
    .A(net79));
 sg13g2_or2_1 \proj_12.or4/_0_  (.X(\proj_12.net7 ),
    .B(net84),
    .A(net80));
 sg13g2_or2_1 \proj_12.or5/_0_  (.X(\proj_12.net4 ),
    .B(net83),
    .A(net79));
 sg13g2_or2_1 \proj_12.or6/_0_  (.X(\proj_12.net5 ),
    .B(net79),
    .A(\proj_12.net14 ));
 sg13g2_and2_1 \proj_13.and1/_0_  (.A(net84),
    .B(net89),
    .X(\proj_13.net12 ));
 sg13g2_and2_1 \proj_13.and2/_0_  (.A(\proj_13.net11 ),
    .B(net80),
    .X(\proj_13.net13 ));
 sg13g2_or2_1 \proj_13.or1/_0_  (.X(\proj_13.net5 ),
    .B(\proj_13.net13 ),
    .A(\proj_13.net12 ));
 sg13g2_xor2_1 \proj_13.xor1/_0_  (.B(\proj_13.net11 ),
    .A(net80),
    .X(\proj_13.net4 ));
 sg13g2_xor2_1 \proj_13.xor2/_0_  (.B(net89),
    .A(net84),
    .X(\proj_13.net11 ));
 sg13g2_and2_1 \proj_14.and1/_0_  (.A(net83),
    .B(net88),
    .X(\proj_14.net6 ));
 sg13g2_inv_1 \proj_14.not1/_0_  (.Y(\proj_14.net7 ),
    .A(net4));
 sg13g2_xor2_1 \proj_14.xor1/_0_  (.B(net3),
    .A(net5),
    .X(\proj_14.net8 ));
 sg13g2_and2_1 \proj__0.and1/_0_  (.A(net4),
    .B(\proj__0.net21 ),
    .X(\proj__0.net22 ));
 sg13g2_and2_1 \proj__0.and10/_0_  (.A(\proj__0.net19 ),
    .B(net86),
    .X(\proj__0.net31 ));
 sg13g2_and2_1 \proj__0.and11/_0_  (.A(\proj__0.net29 ),
    .B(\proj__0.net30 ),
    .X(\proj__0.net32 ));
 sg13g2_and2_1 \proj__0.and12/_0_  (.A(\proj__0.net28 ),
    .B(\proj__0.net31 ),
    .X(\proj__0.net33 ));
 sg13g2_and2_1 \proj__0.and13/_0_  (.A(\proj__0.net33 ),
    .B(\proj__0.net32 ),
    .X(\proj__0.net34 ));
 sg13g2_and2_1 \proj__0.and14/_0_  (.A(\proj__0.net35 ),
    .B(\proj__0.net34 ),
    .X(\proj__0.net9 ));
 sg13g2_and2_1 \proj__0.and15/_0_  (.A(\proj__0.net13 ),
    .B(\proj__0.net10 ),
    .X(\proj__0.net35 ));
 sg13g2_and2_1 \proj__0.and16/_0_  (.A(\proj__0.net11 ),
    .B(\proj__0.net36 ),
    .X(\proj__0.net12 ));
 sg13g2_and2_1 \proj__0.and2/_0_  (.A(\proj__0.net19 ),
    .B(net4),
    .X(\proj__0.net23 ));
 sg13g2_and2_1 \proj__0.and3/_0_  (.A(net82),
    .B(\proj__0.net20 ),
    .X(\proj__0.net25 ));
 sg13g2_and2_1 \proj__0.and4/_0_  (.A(\proj__0.net24 ),
    .B(net81),
    .X(\proj__0.net26 ));
 sg13g2_and2_1 \proj__0.and5/_0_  (.A(\proj__0.net23 ),
    .B(\proj__0.net22 ),
    .X(\proj__0.net13 ));
 sg13g2_and2_1 \proj__0.and6/_0_  (.A(\proj__0.net26 ),
    .B(\proj__0.net25 ),
    .X(\proj__0.net10 ));
 sg13g2_and2_1 \proj__0.and7/_0_  (.A(\proj__0.net27 ),
    .B(net86),
    .X(\proj__0.net28 ));
 sg13g2_and2_1 \proj__0.and8/_0_  (.A(\proj__0.net21 ),
    .B(net86),
    .X(\proj__0.net29 ));
 sg13g2_and2_1 \proj__0.and9/_0_  (.A(net86),
    .B(\proj__0.net24 ),
    .X(\proj__0.net30 ));
 sg13g2_inv_1 \proj__0.not1/_0_  (.Y(\proj__0.net19 ),
    .A(net5));
 sg13g2_inv_1 \proj__0.not2/_0_  (.Y(\proj__0.net20 ),
    .A(net91));
 sg13g2_inv_1 \proj__0.not3/_0_  (.Y(\proj__0.net21 ),
    .A(net3));
 sg13g2_inv_1 \proj__0.not4/_0_  (.Y(\proj__0.net24 ),
    .A(net78));
 sg13g2_inv_1 \proj__0.not5/_0_  (.Y(\proj__0.net27 ),
    .A(net2));
 sg13g2_inv_1 \proj__0.not6/_0_  (.Y(\proj__0.net11 ),
    .A(\proj__0.net35 ));
 sg13g2_inv_1 \proj__0.not7/_0_  (.Y(\proj__0.net36 ),
    .A(\proj__0.net34 ));
 sg13g2_and2_1 \proj__1.and1/_0_  (.A(net83),
    .B(net89),
    .X(\proj__1.net7 ));
 sg13g2_and2_1 \proj__2.and10/_0_  (.A(net74),
    .B(net75),
    .X(\proj__2.net33 ));
 sg13g2_and2_1 \proj__2.and11/_0_  (.A(net72),
    .B(net74),
    .X(\proj__2.net34 ));
 sg13g2_and2_1 \proj__2.and12/_0_  (.A(net73),
    .B(\proj__2.net17 ),
    .X(\proj__2.net35 ));
 sg13g2_and2_1 \proj__2.and13/_0_  (.A(net72),
    .B(\proj__2.net35 ),
    .X(\proj__2.net36 ));
 sg13g2_and2_1 \proj__2.and14/_0_  (.A(net87),
    .B(\proj__2.net17 ),
    .X(\proj__2.net37 ));
 sg13g2_and2_1 \proj__2.and15/_0_  (.A(net90),
    .B(\proj__2.net37 ),
    .X(\proj__2.net38 ));
 sg13g2_and2_1 \proj__2.and16/_0_  (.A(net73),
    .B(net77),
    .X(\proj__2.net39 ));
 sg13g2_and2_1 \proj__2.and17/_0_  (.A(net90),
    .B(\proj__2.net39 ),
    .X(\proj__2.net40 ));
 sg13g2_and2_1 \proj__2.and18/_0_  (.A(net73),
    .B(net75),
    .X(\proj__2.net44 ));
 sg13g2_and2_1 \proj__2.and19/_0_  (.A(net90),
    .B(net75),
    .X(\proj__2.net45 ));
 sg13g2_and2_1 \proj__2.and2/_0_  (.A(net72),
    .B(net74),
    .X(\proj__2.net21 ));
 sg13g2_and2_1 \proj__2.and20/_0_  (.A(net90),
    .B(net73),
    .X(\proj__2.net46 ));
 sg13g2_and2_1 \proj__2.and21/_0_  (.A(net82),
    .B(net75),
    .X(\proj__2.net47 ));
 sg13g2_and2_1 \proj__2.and22/_0_  (.A(net74),
    .B(net76),
    .X(\proj__2.net48 ));
 sg13g2_and2_1 \proj__2.and23/_0_  (.A(\proj__2.net19 ),
    .B(net77),
    .X(\proj__2.net52 ));
 sg13g2_and2_1 \proj__2.and24/_0_  (.A(net74),
    .B(net75),
    .X(\proj__2.net53 ));
 sg13g2_and2_1 \proj__2.and25/_0_  (.A(net72),
    .B(\proj__2.net53 ),
    .X(\proj__2.net54 ));
 sg13g2_and2_1 \proj__2.and26/_0_  (.A(net87),
    .B(net74),
    .X(\proj__2.net55 ));
 sg13g2_and2_1 \proj__2.and27/_0_  (.A(net91),
    .B(\proj__2.net55 ),
    .X(\proj__2.net56 ));
 sg13g2_and2_1 \proj__2.and28/_0_  (.A(net73),
    .B(net81),
    .X(\proj__2.net57 ));
 sg13g2_and2_1 \proj__2.and29/_0_  (.A(net91),
    .B(\proj__2.net57 ),
    .X(\proj__2.net58 ));
 sg13g2_and2_1 \proj__2.and3/_0_  (.A(net87),
    .B(net75),
    .X(\proj__2.net22 ));
 sg13g2_and2_1 \proj__2.and30/_0_  (.A(net87),
    .B(net82),
    .X(\proj__2.net59 ));
 sg13g2_and2_1 \proj__2.and31/_0_  (.A(net72),
    .B(\proj__2.net59 ),
    .X(\proj__2.net60 ));
 sg13g2_and2_1 \proj__2.and32/_0_  (.A(net72),
    .B(\proj__2.net18 ),
    .X(\proj__2.net64 ));
 sg13g2_and2_1 \proj__2.and33/_0_  (.A(\proj__2.net20 ),
    .B(net85),
    .X(\proj__2.net65 ));
 sg13g2_and2_1 \proj__2.and34/_0_  (.A(net85),
    .B(net77),
    .X(\proj__2.net66 ));
 sg13g2_and2_1 \proj__2.and35/_0_  (.A(net81),
    .B(net78),
    .X(\proj__2.net67 ));
 sg13g2_and2_1 \proj__2.and36/_0_  (.A(net72),
    .B(\proj__2.net19 ),
    .X(\proj__2.net70 ));
 sg13g2_and2_1 \proj__2.and37/_0_  (.A(\proj__2.net20 ),
    .B(net81),
    .X(\proj__2.net71 ));
 sg13g2_and2_1 \proj__2.and38/_0_  (.A(net74),
    .B(net77),
    .X(\proj__2.net72 ));
 sg13g2_and2_1 \proj__2.and39/_0_  (.A(net85),
    .B(net77),
    .X(\proj__2.net73 ));
 sg13g2_and2_1 \proj__2.and4/_0_  (.A(net1),
    .B(net80),
    .X(\proj__2.net23 ));
 sg13g2_and2_1 \proj__2.and40/_0_  (.A(net81),
    .B(net75),
    .X(\proj__2.net74 ));
 sg13g2_and2_1 \proj__2.and41/_0_  (.A(net73),
    .B(\proj__2.net74 ),
    .X(\proj__2.net75 ));
 sg13g2_and2_1 \proj__2.and42/_0_  (.A(net85),
    .B(\proj__2.net18 ),
    .X(\proj__2.net79 ));
 sg13g2_and2_1 \proj__2.and43/_0_  (.A(\proj__2.net20 ),
    .B(net85),
    .X(\proj__2.net80 ));
 sg13g2_and2_1 \proj__2.and44/_0_  (.A(\proj__2.net18 ),
    .B(net77),
    .X(\proj__2.net81 ));
 sg13g2_and2_1 \proj__2.and45/_0_  (.A(net91),
    .B(net77),
    .X(\proj__2.net82 ));
 sg13g2_and2_1 \proj__2.and46/_0_  (.A(net81),
    .B(\proj__2.net17 ),
    .X(\proj__2.net83 ));
 sg13g2_and2_1 \proj__2.and47/_0_  (.A(net73),
    .B(\proj__2.net83 ),
    .X(\proj__2.net84 ));
 sg13g2_and2_1 \proj__2.and5/_0_  (.A(net72),
    .B(net76),
    .X(\proj__2.net24 ));
 sg13g2_and2_1 \proj__2.and6/_0_  (.A(net82),
    .B(net75),
    .X(\proj__2.net25 ));
 sg13g2_and2_1 \proj__2.and7/_0_  (.A(net90),
    .B(\proj__2.net25 ),
    .X(\proj__2.net26 ));
 sg13g2_and2_1 \proj__2.and8/_0_  (.A(net74),
    .B(net76),
    .X(\proj__2.net27 ));
 sg13g2_and2_1 \proj__2.and9/_0_  (.A(net73),
    .B(\proj__2.net27 ),
    .X(\proj__2.net28 ));
 sg13g2_inv_1 \proj__2.not1/_0_  (.Y(\proj__2.net17 ),
    .A(net77));
 sg13g2_inv_1 \proj__2.not3/_0_  (.Y(\proj__2.net18 ),
    .A(net81));
 sg13g2_inv_1 \proj__2.not4/_0_  (.Y(\proj__2.net19 ),
    .A(net85));
 sg13g2_inv_1 \proj__2.not5/_0_  (.Y(\proj__2.net20 ),
    .A(net90));
 sg13g2_or2_1 \proj__2.or10/_0_  (.X(\proj__2.net6 ),
    .B(\proj__2.net43 ),
    .A(\proj__2.net40 ));
 sg13g2_or2_1 \proj__2.or11/_0_  (.X(\proj__2.net7 ),
    .B(\proj__2.net51 ),
    .A(\proj__2.net48 ));
 sg13g2_or2_1 \proj__2.or12/_0_  (.X(\proj__2.net49 ),
    .B(\proj__2.net44 ),
    .A(\proj__2.net45 ));
 sg13g2_or2_1 \proj__2.or13/_0_  (.X(\proj__2.net50 ),
    .B(\proj__2.net46 ),
    .A(\proj__2.net47 ));
 sg13g2_or2_1 \proj__2.or14/_0_  (.X(\proj__2.net51 ),
    .B(\proj__2.net49 ),
    .A(\proj__2.net50 ));
 sg13g2_or2_1 \proj__2.or15/_0_  (.X(\proj__2.net61 ),
    .B(\proj__2.net52 ),
    .A(\proj__2.net54 ));
 sg13g2_or2_1 \proj__2.or16/_0_  (.X(\proj__2.net62 ),
    .B(\proj__2.net56 ),
    .A(\proj__2.net58 ));
 sg13g2_or2_1 \proj__2.or17/_0_  (.X(\proj__2.net63 ),
    .B(\proj__2.net61 ),
    .A(\proj__2.net62 ));
 sg13g2_or2_1 \proj__2.or18/_0_  (.X(\proj__2.net8 ),
    .B(\proj__2.net63 ),
    .A(\proj__2.net60 ));
 sg13g2_or2_1 \proj__2.or19/_0_  (.X(\proj__2.net68 ),
    .B(\proj__2.net64 ),
    .A(\proj__2.net65 ));
 sg13g2_or2_1 \proj__2.or2/_0_  (.X(\proj__2.net41 ),
    .B(\proj__2.net33 ),
    .A(\proj__2.net34 ));
 sg13g2_or2_1 \proj__2.or20/_0_  (.X(\proj__2.net69 ),
    .B(\proj__2.net66 ),
    .A(\proj__2.net67 ));
 sg13g2_or2_1 \proj__2.or21/_0_  (.X(\proj__2.net76 ),
    .B(\proj__2.net70 ),
    .A(\proj__2.net71 ));
 sg13g2_or2_1 \proj__2.or22/_0_  (.X(\proj__2.net9 ),
    .B(\proj__2.net68 ),
    .A(\proj__2.net69 ));
 sg13g2_or2_1 \proj__2.or23/_0_  (.X(\proj__2.net77 ),
    .B(\proj__2.net72 ),
    .A(\proj__2.net73 ));
 sg13g2_or2_1 \proj__2.or24/_0_  (.X(\proj__2.net78 ),
    .B(\proj__2.net76 ),
    .A(\proj__2.net77 ));
 sg13g2_or2_1 \proj__2.or25/_0_  (.X(\proj__2.net85 ),
    .B(\proj__2.net79 ),
    .A(\proj__2.net80 ));
 sg13g2_or2_1 \proj__2.or26/_0_  (.X(\proj__2.net10 ),
    .B(\proj__2.net78 ),
    .A(\proj__2.net75 ));
 sg13g2_or2_1 \proj__2.or27/_0_  (.X(\proj__2.net86 ),
    .B(\proj__2.net81 ),
    .A(\proj__2.net82 ));
 sg13g2_or2_1 \proj__2.or28/_0_  (.X(\proj__2.net87 ),
    .B(\proj__2.net85 ),
    .A(\proj__2.net86 ));
 sg13g2_or2_1 \proj__2.or29/_0_  (.X(\proj__2.net11 ),
    .B(\proj__2.net87 ),
    .A(\proj__2.net84 ));
 sg13g2_or2_1 \proj__2.or3/_0_  (.X(\proj__2.net29 ),
    .B(\proj__2.net21 ),
    .A(\proj__2.net22 ));
 sg13g2_or2_1 \proj__2.or4/_0_  (.X(\proj__2.net30 ),
    .B(\proj__2.net23 ),
    .A(\proj__2.net24 ));
 sg13g2_or2_1 \proj__2.or5/_0_  (.X(\proj__2.net31 ),
    .B(\proj__2.net29 ),
    .A(\proj__2.net30 ));
 sg13g2_or2_1 \proj__2.or6/_0_  (.X(\proj__2.net32 ),
    .B(\proj__2.net26 ),
    .A(\proj__2.net28 ));
 sg13g2_or2_1 \proj__2.or7/_0_  (.X(\proj__2.net5 ),
    .B(\proj__2.net31 ),
    .A(\proj__2.net32 ));
 sg13g2_or2_1 \proj__2.or8/_0_  (.X(\proj__2.net42 ),
    .B(\proj__2.net36 ),
    .A(\proj__2.net38 ));
 sg13g2_or2_1 \proj__2.or9/_0_  (.X(\proj__2.net43 ),
    .B(\proj__2.net41 ),
    .A(\proj__2.net42 ));
 sg13g2_and2_1 \proj__3.and1/_0_  (.A(\proj__3.net20 ),
    .B(net3),
    .X(\proj__3.net12 ));
 sg13g2_and2_1 \proj__3.and2/_0_  (.A(\proj__3.net21 ),
    .B(net2),
    .X(\proj__3.net11 ));
 sg13g2_and2_1 \proj__3.and3/_0_  (.A(\proj__3.net18 ),
    .B(net90),
    .X(\proj__3.net9 ));
 sg13g2_and2_1 \proj__3.and4/_0_  (.A(\proj__3.net19 ),
    .B(net82),
    .X(\proj__3.net10 ));
 sg13g2_inv_1 \proj__3.not1/_0_  (.Y(\proj__3.net18 ),
    .A(net5));
 sg13g2_inv_1 \proj__3.not2/_0_  (.Y(\proj__3.net19 ),
    .A(net4));
 sg13g2_inv_1 \proj__3.not3/_0_  (.Y(\proj__3.net20 ),
    .A(net85));
 sg13g2_inv_1 \proj__3.not4/_0_  (.Y(\proj__3.net21 ),
    .A(net78));
 sg13g2_inv_1 \proj__4.not1/_0_  (.Y(\proj__4.net9 ),
    .A(net89));
 sg13g2_inv_1 \proj__4.not2/_0_  (.Y(\proj__4.net10 ),
    .A(net84));
 sg13g2_inv_1 \proj__4.not3/_0_  (.Y(\proj__4.net11 ),
    .A(net82));
 sg13g2_inv_1 \proj__4.not4/_0_  (.Y(\proj__4.net12 ),
    .A(net76));
 sg13g2_and2_1 \proj__5.and1/_0_  (.A(net80),
    .B(net84),
    .X(\proj__5.net7 ));
 sg13g2_nand2_1 \proj__5.nand1/_0_  (.Y(\proj__5.net9 ),
    .A(net5),
    .B(net4));
 sg13g2_or2_1 \proj__5.or1/_0_  (.X(\proj__5.net8 ),
    .B(net78),
    .A(net2));
 sg13g2_and2_1 \proj__6.and1/_0_  (.A(net84),
    .B(net89),
    .X(\proj__6.net9 ));
 sg13g2_xor2_1 \proj__6.xor1/_0_  (.B(net80),
    .A(net76),
    .X(\proj__6.net10 ));
 sg13g2_and2_1 \proj__7.and1/_0_  (.A(net76),
    .B(net84),
    .X(\proj__7.net21 ));
 sg13g2_and2_1 \proj__7.and2/_0_  (.A(net80),
    .B(net83),
    .X(\proj__7.net22 ));
 sg13g2_and2_1 \proj__7.and3/_0_  (.A(net76),
    .B(net89),
    .X(\proj__7.net23 ));
 sg13g2_and2_1 \proj__7.and4/_0_  (.A(net79),
    .B(net88),
    .X(\proj__7.net9 ));
 sg13g2_and2_1 \proj__7.and5/_0_  (.A(\proj__7.net23 ),
    .B(\proj__7.net22 ),
    .X(\proj__7.net24 ));
 sg13g2_and2_1 \proj__7.and6/_0_  (.A(\proj__7.net21 ),
    .B(\proj__7.net24 ),
    .X(\proj__7.net12 ));
 sg13g2_and2_1 \proj__7.and7/_0_  (.A(net5),
    .B(net3),
    .X(\proj__7.net26 ));
 sg13g2_and2_1 \proj__7.and8/_0_  (.A(net4),
    .B(net2),
    .X(\proj__7.net27 ));
 sg13g2_and2_1 \proj__7.and9/_0_  (.A(\proj__7.net25 ),
    .B(\proj__7.net27 ),
    .X(\proj__7.net28 ));
 sg13g2_or2_1 \proj__7.or1/_0_  (.X(\proj__7.net15 ),
    .B(\proj__7.net28 ),
    .A(\proj__7.net26 ));
 sg13g2_xor2_1 \proj__7.xor1/_0_  (.B(\proj__7.net23 ),
    .A(\proj__7.net22 ),
    .X(\proj__7.net10 ));
 sg13g2_xor2_1 \proj__7.xor2/_0_  (.B(\proj__7.net24 ),
    .A(\proj__7.net21 ),
    .X(\proj__7.net11 ));
 sg13g2_xor2_1 \proj__7.xor3/_0_  (.B(net3),
    .A(net5),
    .X(\proj__7.net25 ));
 sg13g2_xor2_1 \proj__7.xor4/_0_  (.B(net2),
    .A(net4),
    .X(\proj__7.net13 ));
 sg13g2_xor2_1 \proj__7.xor5/_0_  (.B(\proj__7.net27 ),
    .A(\proj__7.net25 ),
    .X(\proj__7.net14 ));
 sg13g2_and2_1 \proj__8.and1/_0_  (.A(net79),
    .B(\proj__8.net10 ),
    .X(\proj__8.net11 ));
 sg13g2_and2_1 \proj__8.and2/_0_  (.A(net83),
    .B(net88),
    .X(\proj__8.net12 ));
 sg13g2_or2_1 \proj__8.or1/_0_  (.X(\proj__8.net5 ),
    .B(\proj__8.net11 ),
    .A(\proj__8.net12 ));
 sg13g2_xor2_1 \proj__8.xor1/_0_  (.B(net88),
    .A(net83),
    .X(\proj__8.net10 ));
 sg13g2_xor2_1 \proj__8.xor2/_0_  (.B(\proj__8.net10 ),
    .A(net79),
    .X(\proj__8.net4 ));
 sg13g2_inv_1 \proj__9.not1/_0_  (.Y(\proj__9.net9 ),
    .A(net88));
 sg13g2_inv_1 \proj__9.not2/_0_  (.Y(\proj__9.net10 ),
    .A(net83));
 sg13g2_inv_1 \proj__9.not3/_0_  (.Y(\proj__9.net11 ),
    .A(net79));
 sg13g2_inv_1 \proj__9.not4/_0_  (.Y(\proj__9.net12 ),
    .A(net76));
 sg13g2_buf_2 fanout71 (.A(_069_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(\proj__2.net20 ),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(\proj__2.net19 ),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(\proj__2.net18 ),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(\proj__2.net17 ),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(net78),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(net78),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(ui_in[3]),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(net80),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(ui_in[2]),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(net82),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(ui_in[2]),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(net84),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(net1),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(net87),
    .X(net85));
 sg13g2_buf_1 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(net1),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(net89),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(ui_in[0]),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(ui_in[0]),
    .X(net90));
 sg13g2_buf_1 fanout91 (.A(ui_in[0]),
    .X(net91));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[4]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[6]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_tielo \proj_10.flop1/_1__10  (.L_LO(net10));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_4 FILLER_26_280 ();
 sg13g2_fill_1 FILLER_26_284 ();
 sg13g2_decap_8 FILLER_26_290 ();
 sg13g2_decap_8 FILLER_26_297 ();
 sg13g2_decap_4 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_318 ();
 sg13g2_decap_8 FILLER_26_325 ();
 sg13g2_fill_1 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_338 ();
 sg13g2_fill_2 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_fill_2 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_4 FILLER_27_245 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_decap_8 FILLER_27_258 ();
 sg13g2_decap_8 FILLER_27_265 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_fill_1 FILLER_27_279 ();
 sg13g2_decap_4 FILLER_27_300 ();
 sg13g2_fill_2 FILLER_27_324 ();
 sg13g2_decap_4 FILLER_27_346 ();
 sg13g2_fill_1 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_8 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_245 ();
 sg13g2_decap_4 FILLER_28_264 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_decap_8 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_282 ();
 sg13g2_decap_4 FILLER_28_289 ();
 sg13g2_decap_4 FILLER_28_313 ();
 sg13g2_decap_4 FILLER_28_322 ();
 sg13g2_decap_4 FILLER_28_346 ();
 sg13g2_fill_2 FILLER_28_350 ();
 sg13g2_decap_4 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_371 ();
 sg13g2_decap_4 FILLER_28_377 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_4 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_fill_1 FILLER_29_247 ();
 sg13g2_decap_4 FILLER_29_263 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_decap_8 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_240 ();
 sg13g2_decap_4 FILLER_30_263 ();
 sg13g2_decap_4 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_294 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_decap_4 FILLER_30_302 ();
 sg13g2_decap_4 FILLER_30_316 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_fill_2 FILLER_30_336 ();
 sg13g2_decap_4 FILLER_30_356 ();
 sg13g2_decap_4 FILLER_30_370 ();
 sg13g2_fill_1 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_4 FILLER_31_182 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_decap_8 FILLER_31_191 ();
 sg13g2_decap_8 FILLER_31_198 ();
 sg13g2_decap_8 FILLER_31_205 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_fill_2 FILLER_31_219 ();
 sg13g2_fill_1 FILLER_31_221 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_decap_8 FILLER_31_237 ();
 sg13g2_fill_1 FILLER_31_250 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_decap_4 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_290 ();
 sg13g2_fill_1 FILLER_31_304 ();
 sg13g2_decap_4 FILLER_31_308 ();
 sg13g2_decap_4 FILLER_31_316 ();
 sg13g2_decap_8 FILLER_31_323 ();
 sg13g2_decap_4 FILLER_31_330 ();
 sg13g2_fill_2 FILLER_31_334 ();
 sg13g2_decap_4 FILLER_31_341 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_fill_2 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_fill_1 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_288 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_319 ();
 sg13g2_fill_2 FILLER_32_333 ();
 sg13g2_fill_2 FILLER_32_346 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_decap_4 FILLER_32_370 ();
 sg13g2_fill_2 FILLER_32_374 ();
 sg13g2_decap_4 FILLER_32_386 ();
 sg13g2_fill_2 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_4 FILLER_33_189 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_decap_8 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_218 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_244 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_269 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_323 ();
 sg13g2_decap_8 FILLER_33_330 ();
 sg13g2_fill_2 FILLER_33_340 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_decap_4 FILLER_33_358 ();
 sg13g2_fill_2 FILLER_33_362 ();
 sg13g2_decap_4 FILLER_33_372 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_fill_2 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_264 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_fill_2 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_decap_4 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_340 ();
 sg13g2_fill_1 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_fill_1 FILLER_35_198 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_222 ();
 sg13g2_decap_8 FILLER_35_228 ();
 sg13g2_fill_2 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_decap_4 FILLER_35_259 ();
 sg13g2_fill_1 FILLER_35_263 ();
 sg13g2_decap_4 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_272 ();
 sg13g2_fill_2 FILLER_35_284 ();
 sg13g2_decap_4 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_decap_4 FILLER_35_330 ();
 sg13g2_fill_2 FILLER_35_355 ();
 sg13g2_decap_8 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_decap_8 FILLER_35_383 ();
 sg13g2_decap_8 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_4 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_200 ();
 sg13g2_decap_4 FILLER_36_235 ();
 sg13g2_fill_2 FILLER_36_239 ();
 sg13g2_fill_2 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_279 ();
 sg13g2_fill_1 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_288 ();
 sg13g2_decap_8 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_302 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_2 FILLER_36_332 ();
 sg13g2_fill_2 FILLER_36_356 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_fill_2 FILLER_37_210 ();
 sg13g2_fill_1 FILLER_37_212 ();
 sg13g2_decap_4 FILLER_37_242 ();
 sg13g2_fill_2 FILLER_37_246 ();
 sg13g2_decap_4 FILLER_37_261 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_290 ();
 sg13g2_fill_2 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_305 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_325 ();
 sg13g2_fill_1 FILLER_37_345 ();
 sg13g2_decap_8 FILLER_37_356 ();
 sg13g2_decap_8 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_370 ();
 sg13g2_decap_8 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_37_384 ();
 sg13g2_decap_8 FILLER_37_391 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_4 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_219 ();
 sg13g2_fill_2 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_4 FILLER_38_245 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_262 ();
 sg13g2_decap_8 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net17;
 assign uio_oe[5] = net18;
 assign uio_oe[6] = net19;
 assign uio_oe[7] = net20;
 assign uio_out[0] = net21;
 assign uio_out[1] = net22;
 assign uio_out[2] = net23;
 assign uio_out[3] = net24;
 assign uio_out[4] = net25;
 assign uio_out[5] = net26;
 assign uio_out[6] = net27;
 assign uio_out[7] = net28;
endmodule

module tt_um_zec_square1 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire \frame_no[0] ;
 wire \frame_no[1] ;
 wire \frame_no[2] ;
 wire \frame_no[3] ;
 wire \frame_no[4] ;
 wire \frame_no[5] ;
 wire \frame_no[6] ;
 wire \frame_no[7] ;
 wire \frame_no[8] ;
 wire \hpos[0] ;
 wire \hpos[1] ;
 wire \hpos[2] ;
 wire \hpos[3] ;
 wire \hpos[4] ;
 wire \hpos[5] ;
 wire \hpos[6] ;
 wire \hpos[7] ;
 wire \hpos[8] ;
 wire \hpos[9] ;
 wire hsync;
 wire prev_vsync;
 wire \project_audio.f_counter[0] ;
 wire \project_audio.f_counter[1] ;
 wire \project_audio.f_counter[2] ;
 wire \project_audio.freq[0][0] ;
 wire \project_audio.freq[0][10] ;
 wire \project_audio.freq[0][11] ;
 wire \project_audio.freq[0][1] ;
 wire \project_audio.freq[0][2] ;
 wire \project_audio.freq[0][3] ;
 wire \project_audio.freq[0][4] ;
 wire \project_audio.freq[0][5] ;
 wire \project_audio.freq[0][6] ;
 wire \project_audio.freq[0][7] ;
 wire \project_audio.freq[0][8] ;
 wire \project_audio.freq[0][9] ;
 wire \project_audio.freq[1][0] ;
 wire \project_audio.freq[1][10] ;
 wire \project_audio.freq[1][11] ;
 wire \project_audio.freq[1][1] ;
 wire \project_audio.freq[1][2] ;
 wire \project_audio.freq[1][3] ;
 wire \project_audio.freq[1][4] ;
 wire \project_audio.freq[1][5] ;
 wire \project_audio.freq[1][6] ;
 wire \project_audio.freq[1][7] ;
 wire \project_audio.freq[1][8] ;
 wire \project_audio.freq[1][9] ;
 wire \project_audio.freq[2][0] ;
 wire \project_audio.freq[2][10] ;
 wire \project_audio.freq[2][11] ;
 wire \project_audio.freq[2][1] ;
 wire \project_audio.freq[2][2] ;
 wire \project_audio.freq[2][3] ;
 wire \project_audio.freq[2][4] ;
 wire \project_audio.freq[2][5] ;
 wire \project_audio.freq[2][6] ;
 wire \project_audio.freq[2][7] ;
 wire \project_audio.freq[2][8] ;
 wire \project_audio.freq[2][9] ;
 wire \project_audio.freq[3][0] ;
 wire \project_audio.freq[3][10] ;
 wire \project_audio.freq[3][11] ;
 wire \project_audio.freq[3][1] ;
 wire \project_audio.freq[3][2] ;
 wire \project_audio.freq[3][3] ;
 wire \project_audio.freq[3][4] ;
 wire \project_audio.freq[3][5] ;
 wire \project_audio.freq[3][6] ;
 wire \project_audio.freq[3][7] ;
 wire \project_audio.freq[3][8] ;
 wire \project_audio.freq[3][9] ;
 wire \project_audio.freq[4][0] ;
 wire \project_audio.freq[4][10] ;
 wire \project_audio.freq[4][11] ;
 wire \project_audio.freq[4][1] ;
 wire \project_audio.freq[4][2] ;
 wire \project_audio.freq[4][3] ;
 wire \project_audio.freq[4][4] ;
 wire \project_audio.freq[4][5] ;
 wire \project_audio.freq[4][6] ;
 wire \project_audio.freq[4][7] ;
 wire \project_audio.freq[4][8] ;
 wire \project_audio.freq[4][9] ;
 wire \project_audio.freq[5][0] ;
 wire \project_audio.freq[5][10] ;
 wire \project_audio.freq[5][11] ;
 wire \project_audio.freq[5][1] ;
 wire \project_audio.freq[5][2] ;
 wire \project_audio.freq[5][3] ;
 wire \project_audio.freq[5][4] ;
 wire \project_audio.freq[5][5] ;
 wire \project_audio.freq[5][6] ;
 wire \project_audio.freq[5][7] ;
 wire \project_audio.freq[5][8] ;
 wire \project_audio.freq[5][9] ;
 wire \project_audio.freq[6][0] ;
 wire \project_audio.freq[6][10] ;
 wire \project_audio.freq[6][11] ;
 wire \project_audio.freq[6][1] ;
 wire \project_audio.freq[6][2] ;
 wire \project_audio.freq[6][3] ;
 wire \project_audio.freq[6][4] ;
 wire \project_audio.freq[6][5] ;
 wire \project_audio.freq[6][6] ;
 wire \project_audio.freq[6][7] ;
 wire \project_audio.freq[6][8] ;
 wire \project_audio.freq[6][9] ;
 wire \project_audio.freq[7][0] ;
 wire \project_audio.freq[7][10] ;
 wire \project_audio.freq[7][11] ;
 wire \project_audio.freq[7][1] ;
 wire \project_audio.freq[7][2] ;
 wire \project_audio.freq[7][3] ;
 wire \project_audio.freq[7][4] ;
 wire \project_audio.freq[7][5] ;
 wire \project_audio.freq[7][6] ;
 wire \project_audio.freq[7][7] ;
 wire \project_audio.freq[7][8] ;
 wire \project_audio.freq[7][9] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[0] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[10] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[11] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[12] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[13] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[14] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[15] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[1] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[2] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[3] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[4] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[5] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[6] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[7] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[8] ;
 wire \project_audio.genblk1[0].n_c_oh_my.phase[9] ;
 wire \project_audio.genblk1[0].n_c_oh_my.snd ;
 wire \project_audio.genblk1[0].n_c_oh_my.step ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[0] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[10] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[11] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[12] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[13] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[14] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[15] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[1] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[2] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[3] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[4] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[5] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[6] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[7] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[8] ;
 wire \project_audio.genblk1[1].n_c_oh_my.phase[9] ;
 wire \project_audio.genblk1[1].n_c_oh_my.snd ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[0] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[10] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[11] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[12] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[13] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[14] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[15] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[1] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[2] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[3] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[4] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[5] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[6] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[7] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[8] ;
 wire \project_audio.genblk1[2].n_c_oh_my.phase[9] ;
 wire \project_audio.genblk1[2].n_c_oh_my.snd ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[0] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[10] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[11] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[12] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[13] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[14] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[15] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[1] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[2] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[3] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[4] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[5] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[6] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[7] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[8] ;
 wire \project_audio.genblk1[3].n_c_oh_my.phase[9] ;
 wire \project_audio.genblk1[3].n_c_oh_my.snd ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[0] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[10] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[11] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[12] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[13] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[14] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[15] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[1] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[2] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[3] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[4] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[5] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[6] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[7] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[8] ;
 wire \project_audio.genblk1[4].n_c_oh_my.phase[9] ;
 wire \project_audio.genblk1[4].n_c_oh_my.snd ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[0] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[10] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[11] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[12] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[13] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[14] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[15] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[1] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[2] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[3] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[4] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[5] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[6] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[7] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[8] ;
 wire \project_audio.genblk1[5].n_c_oh_my.phase[9] ;
 wire \project_audio.genblk1[5].n_c_oh_my.snd ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[0] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[10] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[11] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[12] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[13] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[14] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[15] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[1] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[2] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[3] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[4] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[5] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[6] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[7] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[8] ;
 wire \project_audio.genblk1[6].n_c_oh_my.phase[9] ;
 wire \project_audio.genblk1[6].n_c_oh_my.snd ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[0] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[10] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[11] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[12] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[13] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[14] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[15] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[1] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[2] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[3] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[4] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[5] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[6] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[7] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[8] ;
 wire \project_audio.genblk1[7].n_c_oh_my.phase[9] ;
 wire \project_audio.genblk1[7].n_c_oh_my.snd ;
 wire \project_audio.iter.counter[0] ;
 wire \project_audio.iter.counter[10] ;
 wire \project_audio.iter.counter[11] ;
 wire \project_audio.iter.counter[12] ;
 wire \project_audio.iter.counter[13] ;
 wire \project_audio.iter.counter[1] ;
 wire \project_audio.iter.counter[2] ;
 wire \project_audio.iter.counter[3] ;
 wire \project_audio.iter.counter[4] ;
 wire \project_audio.iter.counter[5] ;
 wire \project_audio.iter.counter[6] ;
 wire \project_audio.iter.counter[7] ;
 wire \project_audio.iter.counter[8] ;
 wire \project_audio.iter.counter[9] ;
 wire \project_audio.iter.mult1_shift[0] ;
 wire \project_audio.iter.mult1_shift[10] ;
 wire \project_audio.iter.mult1_shift[11] ;
 wire \project_audio.iter.mult1_shift[12] ;
 wire \project_audio.iter.mult1_shift[13] ;
 wire \project_audio.iter.mult1_shift[14] ;
 wire \project_audio.iter.mult1_shift[15] ;
 wire \project_audio.iter.mult1_shift[16] ;
 wire \project_audio.iter.mult1_shift[17] ;
 wire \project_audio.iter.mult1_shift[18] ;
 wire \project_audio.iter.mult1_shift[19] ;
 wire \project_audio.iter.mult1_shift[1] ;
 wire \project_audio.iter.mult1_shift[20] ;
 wire \project_audio.iter.mult1_shift[21] ;
 wire \project_audio.iter.mult1_shift[22] ;
 wire \project_audio.iter.mult1_shift[23] ;
 wire \project_audio.iter.mult1_shift[24] ;
 wire \project_audio.iter.mult1_shift[25] ;
 wire \project_audio.iter.mult1_shift[26] ;
 wire \project_audio.iter.mult1_shift[27] ;
 wire \project_audio.iter.mult1_shift[28] ;
 wire \project_audio.iter.mult1_shift[29] ;
 wire \project_audio.iter.mult1_shift[2] ;
 wire \project_audio.iter.mult1_shift[30] ;
 wire \project_audio.iter.mult1_shift[31] ;
 wire \project_audio.iter.mult1_shift[3] ;
 wire \project_audio.iter.mult1_shift[4] ;
 wire \project_audio.iter.mult1_shift[5] ;
 wire \project_audio.iter.mult1_shift[6] ;
 wire \project_audio.iter.mult1_shift[7] ;
 wire \project_audio.iter.mult1_shift[8] ;
 wire \project_audio.iter.mult1_shift[9] ;
 wire \project_audio.iter.mult2_shift[0] ;
 wire \project_audio.iter.mult2_shift[10] ;
 wire \project_audio.iter.mult2_shift[11] ;
 wire \project_audio.iter.mult2_shift[12] ;
 wire \project_audio.iter.mult2_shift[13] ;
 wire \project_audio.iter.mult2_shift[14] ;
 wire \project_audio.iter.mult2_shift[15] ;
 wire \project_audio.iter.mult2_shift[1] ;
 wire \project_audio.iter.mult2_shift[2] ;
 wire \project_audio.iter.mult2_shift[3] ;
 wire \project_audio.iter.mult2_shift[4] ;
 wire \project_audio.iter.mult2_shift[5] ;
 wire \project_audio.iter.mult2_shift[6] ;
 wire \project_audio.iter.mult2_shift[7] ;
 wire \project_audio.iter.mult2_shift[8] ;
 wire \project_audio.iter.mult2_shift[9] ;
 wire \project_audio.iter.mult_accum[0] ;
 wire \project_audio.iter.mult_accum[10] ;
 wire \project_audio.iter.mult_accum[11] ;
 wire \project_audio.iter.mult_accum[12] ;
 wire \project_audio.iter.mult_accum[13] ;
 wire \project_audio.iter.mult_accum[14] ;
 wire \project_audio.iter.mult_accum[15] ;
 wire \project_audio.iter.mult_accum[16] ;
 wire \project_audio.iter.mult_accum[17] ;
 wire \project_audio.iter.mult_accum[18] ;
 wire \project_audio.iter.mult_accum[19] ;
 wire \project_audio.iter.mult_accum[1] ;
 wire \project_audio.iter.mult_accum[20] ;
 wire \project_audio.iter.mult_accum[21] ;
 wire \project_audio.iter.mult_accum[22] ;
 wire \project_audio.iter.mult_accum[23] ;
 wire \project_audio.iter.mult_accum[24] ;
 wire \project_audio.iter.mult_accum[25] ;
 wire \project_audio.iter.mult_accum[26] ;
 wire \project_audio.iter.mult_accum[27] ;
 wire \project_audio.iter.mult_accum[28] ;
 wire \project_audio.iter.mult_accum[29] ;
 wire \project_audio.iter.mult_accum[2] ;
 wire \project_audio.iter.mult_accum[30] ;
 wire \project_audio.iter.mult_accum[31] ;
 wire \project_audio.iter.mult_accum[3] ;
 wire \project_audio.iter.mult_accum[4] ;
 wire \project_audio.iter.mult_accum[5] ;
 wire \project_audio.iter.mult_accum[6] ;
 wire \project_audio.iter.mult_accum[7] ;
 wire \project_audio.iter.mult_accum[8] ;
 wire \project_audio.iter.mult_accum[9] ;
 wire \project_audio.iter.next_ready ;
 wire \project_audio.iter.r[0] ;
 wire \project_audio.iter.r[10] ;
 wire \project_audio.iter.r[11] ;
 wire \project_audio.iter.r[12] ;
 wire \project_audio.iter.r[13] ;
 wire \project_audio.iter.r[14] ;
 wire \project_audio.iter.r[15] ;
 wire \project_audio.iter.r[16] ;
 wire \project_audio.iter.r[17] ;
 wire \project_audio.iter.r[1] ;
 wire \project_audio.iter.r[2] ;
 wire \project_audio.iter.r[3] ;
 wire \project_audio.iter.r[4] ;
 wire \project_audio.iter.r[5] ;
 wire \project_audio.iter.r[6] ;
 wire \project_audio.iter.r[7] ;
 wire \project_audio.iter.r[8] ;
 wire \project_audio.iter.r[9] ;
 wire \project_audio.iter.x[0] ;
 wire \project_audio.iter.x[10] ;
 wire \project_audio.iter.x[11] ;
 wire \project_audio.iter.x[12] ;
 wire \project_audio.iter.x[13] ;
 wire \project_audio.iter.x[14] ;
 wire \project_audio.iter.x[15] ;
 wire \project_audio.iter.x[1] ;
 wire \project_audio.iter.x[2] ;
 wire \project_audio.iter.x[3] ;
 wire \project_audio.iter.x[4] ;
 wire \project_audio.iter.x[5] ;
 wire \project_audio.iter.x[6] ;
 wire \project_audio.iter.x[7] ;
 wire \project_audio.iter.x[8] ;
 wire \project_audio.iter.x[9] ;
 wire \project_audio.mixer.audio_out ;
 wire \project_audio.mixer.counter[0] ;
 wire \project_audio.mixer.counter[1] ;
 wire \project_audio.mixer.counter[2] ;
 wire \project_audio.mixer.counter[3] ;
 wire \project_audio.nco_increment_gen.counter[0] ;
 wire \project_audio.nco_increment_gen.counter[1] ;
 wire \project_audio.nco_increment_gen.counter[2] ;
 wire \project_audio.nco_increment_gen.counter[3] ;
 wire \project_audio.nco_increment_gen.counter[4] ;
 wire \project_audio.nco_increment_gen.counter[5] ;
 wire \project_audio.nco_increment_gen.counter[6] ;
 wire \project_audio.nco_increment_gen.counter[7] ;
 wire \project_audio.nco_increment_gen.counter[8] ;
 wire \project_audio.r_counter ;
 wire \sync_gen.vpos[0] ;
 wire \sync_gen.vpos[1] ;
 wire \sync_gen.vpos[2] ;
 wire \sync_gen.vpos[3] ;
 wire \sync_gen.vpos[4] ;
 wire \sync_gen.vpos[5] ;
 wire \sync_gen.vpos[6] ;
 wire \sync_gen.vpos[7] ;
 wire \sync_gen.vpos[8] ;
 wire \sync_gen.vpos[9] ;
 wire \sync_gen.vsync ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_leaf_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net1;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;

 sg13g2_inv_1 _3362_ (.Y(_2452_),
    .A(net1216));
 sg13g2_inv_2 _3363_ (.Y(_2453_),
    .A(net1198));
 sg13g2_inv_2 _3364_ (.Y(_2454_),
    .A(net626));
 sg13g2_inv_1 _3365_ (.Y(_2455_),
    .A(net627));
 sg13g2_inv_1 _3366_ (.Y(_2456_),
    .A(net629));
 sg13g2_inv_1 _3367_ (.Y(_2457_),
    .A(net1146));
 sg13g2_inv_1 _3368_ (.Y(_2458_),
    .A(net1204));
 sg13g2_inv_1 _3369_ (.Y(_2459_),
    .A(net1200));
 sg13g2_inv_1 _3370_ (.Y(_2460_),
    .A(net1218));
 sg13g2_inv_1 _3371_ (.Y(_2461_),
    .A(net1186));
 sg13g2_inv_1 _3372_ (.Y(_2462_),
    .A(net1158));
 sg13g2_inv_1 _3373_ (.Y(_2463_),
    .A(net1229));
 sg13g2_inv_1 _3374_ (.Y(_2464_),
    .A(net1238));
 sg13g2_inv_2 _3375_ (.Y(_2465_),
    .A(net1234));
 sg13g2_inv_2 _3376_ (.Y(_2466_),
    .A(net858));
 sg13g2_inv_2 _3377_ (.Y(_2467_),
    .A(net1224));
 sg13g2_inv_2 _3378_ (.Y(_2468_),
    .A(net1223));
 sg13g2_inv_1 _3379_ (.Y(_2469_),
    .A(net1219));
 sg13g2_inv_1 _3380_ (.Y(_2470_),
    .A(\project_audio.iter.mult_accum[16] ));
 sg13g2_inv_1 _3381_ (.Y(_2471_),
    .A(net455));
 sg13g2_inv_1 _3382_ (.Y(_2472_),
    .A(net740));
 sg13g2_inv_1 _3383_ (.Y(_2473_),
    .A(net538));
 sg13g2_inv_1 _3384_ (.Y(_2474_),
    .A(net483));
 sg13g2_inv_1 _3385_ (.Y(_2475_),
    .A(net511));
 sg13g2_inv_1 _3386_ (.Y(_2476_),
    .A(net756));
 sg13g2_inv_1 _3387_ (.Y(_2477_),
    .A(net476));
 sg13g2_inv_1 _3388_ (.Y(_2478_),
    .A(net525));
 sg13g2_inv_1 _3389_ (.Y(_2479_),
    .A(net748));
 sg13g2_inv_1 _3390_ (.Y(_2480_),
    .A(net480));
 sg13g2_inv_1 _3391_ (.Y(_2481_),
    .A(net492));
 sg13g2_inv_1 _3392_ (.Y(_2482_),
    .A(net786));
 sg13g2_inv_1 _3393_ (.Y(_2483_),
    .A(net487));
 sg13g2_inv_1 _3394_ (.Y(_2484_),
    .A(net494));
 sg13g2_inv_1 _3395_ (.Y(_2485_),
    .A(net795));
 sg13g2_inv_1 _3396_ (.Y(_2486_),
    .A(net510));
 sg13g2_inv_1 _3397_ (.Y(_2487_),
    .A(net530));
 sg13g2_inv_1 _3398_ (.Y(_2488_),
    .A(net736));
 sg13g2_inv_1 _3399_ (.Y(_2489_),
    .A(net503));
 sg13g2_inv_1 _3400_ (.Y(_2490_),
    .A(net535));
 sg13g2_inv_1 _3401_ (.Y(_2491_),
    .A(net735));
 sg13g2_inv_1 _3402_ (.Y(_2492_),
    .A(net524));
 sg13g2_inv_1 _3403_ (.Y(_2493_),
    .A(net1055));
 sg13g2_inv_1 _3404_ (.Y(_2494_),
    .A(\project_audio.iter.mult1_shift[29] ));
 sg13g2_inv_1 _3405_ (.Y(_2495_),
    .A(net800));
 sg13g2_inv_1 _3406_ (.Y(_2496_),
    .A(\project_audio.iter.mult1_shift[27] ));
 sg13g2_inv_1 _3407_ (.Y(_2497_),
    .A(net867));
 sg13g2_inv_1 _3408_ (.Y(_2498_),
    .A(\project_audio.iter.mult1_shift[25] ));
 sg13g2_inv_1 _3409_ (.Y(_2499_),
    .A(\project_audio.iter.mult1_shift[24] ));
 sg13g2_inv_1 _3410_ (.Y(_2500_),
    .A(net819));
 sg13g2_inv_1 _3411_ (.Y(_2501_),
    .A(net891));
 sg13g2_inv_1 _3412_ (.Y(_2502_),
    .A(net948));
 sg13g2_inv_1 _3413_ (.Y(_2503_),
    .A(\project_audio.iter.mult1_shift[20] ));
 sg13g2_inv_1 _3414_ (.Y(_2504_),
    .A(net887));
 sg13g2_inv_1 _3415_ (.Y(_2505_),
    .A(net1062));
 sg13g2_inv_1 _3416_ (.Y(_2506_),
    .A(\sync_gen.vpos[7] ));
 sg13g2_inv_2 _3417_ (.Y(_2507_),
    .A(net1225));
 sg13g2_inv_1 _3418_ (.Y(_2508_),
    .A(\sync_gen.vpos[5] ));
 sg13g2_inv_1 _3419_ (.Y(_2509_),
    .A(\frame_no[4] ));
 sg13g2_inv_1 _3420_ (.Y(_2510_),
    .A(net439));
 sg13g2_inv_1 _3421_ (.Y(_2511_),
    .A(\project_audio.iter.counter[0] ));
 sg13g2_inv_1 _3422_ (.Y(_2512_),
    .A(_0021_));
 sg13g2_inv_1 _3423_ (.Y(_2513_),
    .A(net693));
 sg13g2_inv_1 _3424_ (.Y(_2514_),
    .A(net827));
 sg13g2_inv_1 _3425_ (.Y(_2515_),
    .A(_0001_));
 sg13g2_inv_1 _3426_ (.Y(_2516_),
    .A(net1189));
 sg13g2_inv_1 _3427_ (.Y(_2517_),
    .A(\project_audio.iter.mult1_shift[9] ));
 sg13g2_inv_1 _3428_ (.Y(_2518_),
    .A(_0017_));
 sg13g2_inv_1 _3429_ (.Y(_2519_),
    .A(net760));
 sg13g2_or4_1 _3430_ (.A(\project_audio.iter.counter[9] ),
    .B(\project_audio.iter.counter[8] ),
    .C(\project_audio.iter.counter[11] ),
    .D(\project_audio.iter.counter[12] ),
    .X(_2520_));
 sg13g2_nor3_2 _3431_ (.A(\project_audio.iter.counter[10] ),
    .B(\project_audio.iter.counter[13] ),
    .C(_2520_),
    .Y(_2521_));
 sg13g2_nor2_1 _3432_ (.A(\project_audio.iter.counter[7] ),
    .B(\project_audio.iter.counter[6] ),
    .Y(_2522_));
 sg13g2_nor3_2 _3433_ (.A(\project_audio.iter.counter[5] ),
    .B(\project_audio.iter.counter[7] ),
    .C(\project_audio.iter.counter[6] ),
    .Y(_2523_));
 sg13g2_nand2_2 _3434_ (.Y(_2524_),
    .A(_2521_),
    .B(_2523_));
 sg13g2_nor3_2 _3435_ (.A(\project_audio.iter.counter[3] ),
    .B(\project_audio.iter.counter[2] ),
    .C(\project_audio.iter.counter[4] ),
    .Y(_2525_));
 sg13g2_nand2_1 _3436_ (.Y(_2526_),
    .A(_2522_),
    .B(_2525_));
 sg13g2_nand2b_1 _3437_ (.Y(_2527_),
    .B(_2521_),
    .A_N(\project_audio.iter.counter[1] ));
 sg13g2_nor3_1 _3438_ (.A(\project_audio.iter.counter[1] ),
    .B(\project_audio.iter.counter[3] ),
    .C(\project_audio.iter.counter[2] ),
    .Y(_2528_));
 sg13g2_o21ai_1 _3439_ (.B1(_2524_),
    .Y(_2529_),
    .A1(_2526_),
    .A2(_2527_));
 sg13g2_inv_1 _3440_ (.Y(_2530_),
    .A(_2529_));
 sg13g2_nand2b_1 _3441_ (.Y(_2531_),
    .B(\project_audio.iter.counter[4] ),
    .A_N(_2528_));
 sg13g2_nor2b_1 _3442_ (.A(\project_audio.iter.counter[8] ),
    .B_N(_2523_),
    .Y(_2532_));
 sg13g2_a21oi_2 _3443_ (.B1(_2530_),
    .Y(_2533_),
    .A2(_2532_),
    .A1(_2531_));
 sg13g2_nand2_1 _3444_ (.Y(_2534_),
    .A(\project_audio.iter.counter[0] ),
    .B(\project_audio.iter.counter[4] ));
 sg13g2_nor2_1 _3445_ (.A(\project_audio.iter.counter[1] ),
    .B(net1211),
    .Y(_2535_));
 sg13g2_and4_1 _3446_ (.A(_2521_),
    .B(_2523_),
    .C(_2531_),
    .D(_2534_),
    .X(_2536_));
 sg13g2_nor2_2 _3447_ (.A(_2533_),
    .B(_2536_),
    .Y(_2537_));
 sg13g2_nor2_1 _3448_ (.A(net682),
    .B(_2530_),
    .Y(_2538_));
 sg13g2_nand2_1 _3449_ (.Y(_2539_),
    .A(net690),
    .B(_2529_));
 sg13g2_nand3b_1 _3450_ (.B(_2537_),
    .C(net567),
    .Y(_2540_),
    .A_N(_0002_));
 sg13g2_nand2_2 _3451_ (.Y(_2541_),
    .A(_2525_),
    .B(_2535_));
 sg13g2_nor2_2 _3452_ (.A(_2524_),
    .B(_2541_),
    .Y(_2542_));
 sg13g2_or2_1 _3453_ (.X(_2543_),
    .B(_2541_),
    .A(_2524_));
 sg13g2_nor2_1 _3454_ (.A(net682),
    .B(_2543_),
    .Y(_2544_));
 sg13g2_a22oi_1 _3455_ (.Y(_2545_),
    .B1(net577),
    .B2(\project_audio.iter.x[0] ),
    .A2(net581),
    .A1(net1119));
 sg13g2_nand2_1 _3456_ (.Y(_0045_),
    .A(_2540_),
    .B(net1120));
 sg13g2_nor2_1 _3457_ (.A(net881),
    .B(net582),
    .Y(_2546_));
 sg13g2_nor2_1 _3458_ (.A(net1045),
    .B(net567),
    .Y(_2547_));
 sg13g2_a21o_1 _3459_ (.A2(net577),
    .A1(_2468_),
    .B1(_2547_),
    .X(_2548_));
 sg13g2_nor2_2 _3460_ (.A(net581),
    .B(_2542_),
    .Y(_2549_));
 sg13g2_nand2_1 _3461_ (.Y(_2550_),
    .A(net567),
    .B(_2543_));
 sg13g2_a21o_1 _3462_ (.A2(_2541_),
    .A1(_2536_),
    .B1(_2533_),
    .X(_2551_));
 sg13g2_a21oi_2 _3463_ (.B1(_2533_),
    .Y(_2552_),
    .A2(_2541_),
    .A1(_2536_));
 sg13g2_nor2_1 _3464_ (.A(net1119),
    .B(_2552_),
    .Y(_2553_));
 sg13g2_a221oi_1 _3465_ (.B2(_2553_),
    .C1(_2548_),
    .B1(_2549_),
    .A1(_2537_),
    .Y(_0046_),
    .A2(_2546_));
 sg13g2_nand2_1 _3466_ (.Y(_2554_),
    .A(_2467_),
    .B(net577));
 sg13g2_o21ai_1 _3467_ (.B1(_2554_),
    .Y(_2555_),
    .A1(net912),
    .A2(net567));
 sg13g2_nand2_1 _3468_ (.Y(_2556_),
    .A(net720),
    .B(net550));
 sg13g2_a21oi_1 _3469_ (.A1(net1045),
    .A2(net555),
    .Y(_2557_),
    .B1(net562));
 sg13g2_a21oi_1 _3470_ (.A1(_2556_),
    .A2(_2557_),
    .Y(_0047_),
    .B1(_2555_));
 sg13g2_nand2_1 _3471_ (.Y(_2558_),
    .A(_2466_),
    .B(net578));
 sg13g2_o21ai_1 _3472_ (.B1(_2558_),
    .Y(_2559_),
    .A1(\project_audio.iter.mult1_shift[3] ),
    .A2(net567));
 sg13g2_nand2_1 _3473_ (.Y(_2560_),
    .A(net485),
    .B(net550));
 sg13g2_a21oi_1 _3474_ (.A1(net912),
    .A2(net555),
    .Y(_2561_),
    .B1(net562));
 sg13g2_a21oi_1 _3475_ (.A1(_2560_),
    .A2(_2561_),
    .Y(_0048_),
    .B1(_2559_));
 sg13g2_nand2_1 _3476_ (.Y(_2562_),
    .A(\project_audio.iter.r[4] ),
    .B(net550));
 sg13g2_a21oi_1 _3477_ (.A1(\project_audio.iter.mult1_shift[3] ),
    .A2(net555),
    .Y(_2563_),
    .B1(_2542_));
 sg13g2_a221oi_1 _3478_ (.B2(_2563_),
    .C1(net581),
    .B1(_2562_),
    .A1(_2465_),
    .Y(_2564_),
    .A2(_2542_));
 sg13g2_a21o_1 _3479_ (.A2(net581),
    .A1(net1080),
    .B1(_2564_),
    .X(_0049_));
 sg13g2_nand2_1 _3480_ (.Y(_2565_),
    .A(\project_audio.iter.r[5] ),
    .B(net550));
 sg13g2_a21oi_1 _3481_ (.A1(net1080),
    .A2(net555),
    .Y(_2566_),
    .B1(_2542_));
 sg13g2_a221oi_1 _3482_ (.B2(_2566_),
    .C1(net581),
    .B1(_2565_),
    .A1(_2464_),
    .Y(_2567_),
    .A2(_2542_));
 sg13g2_a21o_1 _3483_ (.A2(net581),
    .A1(net1142),
    .B1(_2567_),
    .X(_0050_));
 sg13g2_nand2_1 _3484_ (.Y(_2568_),
    .A(_2463_),
    .B(net577));
 sg13g2_o21ai_1 _3485_ (.B1(_2568_),
    .Y(_2569_),
    .A1(\project_audio.iter.mult1_shift[6] ),
    .A2(net567));
 sg13g2_nand2_1 _3486_ (.Y(_2570_),
    .A(net1059),
    .B(net551));
 sg13g2_a21oi_1 _3487_ (.A1(\project_audio.iter.mult1_shift[5] ),
    .A2(net555),
    .Y(_0463_),
    .B1(net562));
 sg13g2_a21oi_1 _3488_ (.A1(_2570_),
    .A2(_0463_),
    .Y(_0051_),
    .B1(_2569_));
 sg13g2_nand2_1 _3489_ (.Y(_0464_),
    .A(_2462_),
    .B(net577));
 sg13g2_o21ai_1 _3490_ (.B1(_0464_),
    .Y(_0465_),
    .A1(net1077),
    .A2(net573));
 sg13g2_nand2_1 _3491_ (.Y(_0466_),
    .A(net1137),
    .B(net550));
 sg13g2_a21oi_1 _3492_ (.A1(\project_audio.iter.mult1_shift[6] ),
    .A2(net556),
    .Y(_0467_),
    .B1(net562));
 sg13g2_a21oi_1 _3493_ (.A1(_0466_),
    .A2(_0467_),
    .Y(_0052_),
    .B1(_0465_));
 sg13g2_nand2_1 _3494_ (.Y(_0468_),
    .A(_2461_),
    .B(net577));
 sg13g2_o21ai_1 _3495_ (.B1(_0468_),
    .Y(_0469_),
    .A1(\project_audio.iter.mult1_shift[8] ),
    .A2(net573));
 sg13g2_nand2_1 _3496_ (.Y(_0470_),
    .A(net904),
    .B(net550));
 sg13g2_a21oi_1 _3497_ (.A1(net1077),
    .A2(net556),
    .Y(_0471_),
    .B1(net562));
 sg13g2_a21oi_1 _3498_ (.A1(_0470_),
    .A2(_0471_),
    .Y(_0053_),
    .B1(_0469_));
 sg13g2_nand2_1 _3499_ (.Y(_0472_),
    .A(net1135),
    .B(net556));
 sg13g2_a21oi_1 _3500_ (.A1(\project_audio.iter.r[9] ),
    .A2(net550),
    .Y(_0473_),
    .B1(net563));
 sg13g2_nor3_1 _3501_ (.A(\project_audio.iter.x[9] ),
    .B(net581),
    .C(_2543_),
    .Y(_0474_));
 sg13g2_a221oi_1 _3502_ (.B2(_0473_),
    .C1(_0474_),
    .B1(_0472_),
    .A1(_2517_),
    .Y(_0054_),
    .A2(net581));
 sg13g2_nand2_1 _3503_ (.Y(_0475_),
    .A(_2459_),
    .B(net580));
 sg13g2_o21ai_1 _3504_ (.B1(_0475_),
    .Y(_0476_),
    .A1(net1167),
    .A2(net573));
 sg13g2_nand2_1 _3505_ (.Y(_0477_),
    .A(net1152),
    .B(net550));
 sg13g2_a21oi_1 _3506_ (.A1(\project_audio.iter.mult1_shift[9] ),
    .A2(net556),
    .Y(_0478_),
    .B1(net563));
 sg13g2_a21oi_1 _3507_ (.A1(_0477_),
    .A2(_0478_),
    .Y(_0055_),
    .B1(_0476_));
 sg13g2_nand2_1 _3508_ (.Y(_0479_),
    .A(_2458_),
    .B(net580));
 sg13g2_o21ai_1 _3509_ (.B1(_0479_),
    .Y(_0480_),
    .A1(net1057),
    .A2(net574));
 sg13g2_nand2_1 _3510_ (.Y(_0481_),
    .A(net1000),
    .B(net551));
 sg13g2_a21oi_1 _3511_ (.A1(\project_audio.iter.mult1_shift[10] ),
    .A2(net556),
    .Y(_0482_),
    .B1(net563));
 sg13g2_a21oi_1 _3512_ (.A1(_0481_),
    .A2(_0482_),
    .Y(_0056_),
    .B1(_0480_));
 sg13g2_nand2_1 _3513_ (.Y(_0483_),
    .A(\project_audio.iter.r[12] ),
    .B(net551));
 sg13g2_a21oi_1 _3514_ (.A1(\project_audio.iter.mult1_shift[11] ),
    .A2(net556),
    .Y(_0484_),
    .B1(_2542_));
 sg13g2_a221oi_1 _3515_ (.B2(_0484_),
    .C1(net582),
    .B1(_0483_),
    .A1(_2456_),
    .Y(_0485_),
    .A2(_2542_));
 sg13g2_a21o_1 _3516_ (.A2(net582),
    .A1(net1147),
    .B1(_0485_),
    .X(_0057_));
 sg13g2_nand2_1 _3517_ (.Y(_0486_),
    .A(_2455_),
    .B(net580));
 sg13g2_o21ai_1 _3518_ (.B1(_0486_),
    .Y(_0487_),
    .A1(net1173),
    .A2(net574));
 sg13g2_nand2_1 _3519_ (.Y(_0488_),
    .A(net1150),
    .B(net551));
 sg13g2_a21oi_1 _3520_ (.A1(net1147),
    .A2(net556),
    .Y(_0489_),
    .B1(net563));
 sg13g2_a21oi_1 _3521_ (.A1(_0488_),
    .A2(_0489_),
    .Y(_0058_),
    .B1(_0487_));
 sg13g2_nand2_1 _3522_ (.Y(_0490_),
    .A(_2454_),
    .B(net577));
 sg13g2_o21ai_1 _3523_ (.B1(_0490_),
    .Y(_0491_),
    .A1(net1190),
    .A2(net574));
 sg13g2_nand2_1 _3524_ (.Y(_0492_),
    .A(\project_audio.iter.r[14] ),
    .B(net552));
 sg13g2_a21oi_1 _3525_ (.A1(net1173),
    .A2(net557),
    .Y(_0493_),
    .B1(net562));
 sg13g2_a21oi_1 _3526_ (.A1(_0492_),
    .A2(_0493_),
    .Y(_0059_),
    .B1(_0491_));
 sg13g2_nand2_1 _3527_ (.Y(_0494_),
    .A(_2453_),
    .B(net577));
 sg13g2_o21ai_1 _3528_ (.B1(_0494_),
    .Y(_0495_),
    .A1(net1170),
    .A2(net574));
 sg13g2_nand2_1 _3529_ (.Y(_0496_),
    .A(net1139),
    .B(net552));
 sg13g2_a21oi_1 _3530_ (.A1(\project_audio.iter.mult1_shift[14] ),
    .A2(net556),
    .Y(_0497_),
    .B1(net562));
 sg13g2_a21oi_1 _3531_ (.A1(_0496_),
    .A2(_0497_),
    .Y(_0060_),
    .B1(_0495_));
 sg13g2_and2_1 _3532_ (.A(\project_audio.iter.next_ready ),
    .B(net688),
    .X(_0498_));
 sg13g2_nand2_2 _3533_ (.Y(_0499_),
    .A(net1182),
    .B(net688));
 sg13g2_nor2_2 _3534_ (.A(_0021_),
    .B(_0499_),
    .Y(_0500_));
 sg13g2_nor2b_2 _3535_ (.A(\project_audio.f_counter[1] ),
    .B_N(\project_audio.f_counter[2] ),
    .Y(_0501_));
 sg13g2_nand2_2 _3536_ (.Y(_0502_),
    .A(_0500_),
    .B(_0501_));
 sg13g2_a21oi_1 _3537_ (.A1(_0500_),
    .A2(_0501_),
    .Y(_0503_),
    .B1(net684));
 sg13g2_nand2_1 _3538_ (.Y(_0504_),
    .A(net474),
    .B(net613));
 sg13g2_nand2_2 _3539_ (.Y(_0505_),
    .A(\project_audio.iter.x[9] ),
    .B(\project_audio.iter.x[8] ));
 sg13g2_nor3_2 _3540_ (.A(_0030_),
    .B(_0031_),
    .C(_0505_),
    .Y(_0506_));
 sg13g2_nand2_2 _3541_ (.Y(_0507_),
    .A(net628),
    .B(\project_audio.iter.x[11] ));
 sg13g2_nor2_1 _3542_ (.A(net627),
    .B(_0507_),
    .Y(_0508_));
 sg13g2_xor2_1 _3543_ (.B(\project_audio.iter.x[8] ),
    .A(\project_audio.iter.x[9] ),
    .X(_0509_));
 sg13g2_nand2_2 _3544_ (.Y(_0510_),
    .A(net627),
    .B(net628));
 sg13g2_xor2_1 _3545_ (.B(net628),
    .A(net627),
    .X(_0511_));
 sg13g2_mux2_1 _3546_ (.A0(net627),
    .A1(_0511_),
    .S(_0507_),
    .X(_0512_));
 sg13g2_a21oi_1 _3547_ (.A1(_0509_),
    .A2(_0512_),
    .Y(_0513_),
    .B1(_0508_));
 sg13g2_nand2_2 _3548_ (.Y(_0514_),
    .A(\project_audio.iter.x[10] ),
    .B(\project_audio.iter.x[9] ));
 sg13g2_xor2_1 _3549_ (.B(\project_audio.iter.x[9] ),
    .A(\project_audio.iter.x[10] ),
    .X(_0515_));
 sg13g2_nor2_1 _3550_ (.A(net625),
    .B(_0510_),
    .Y(_0516_));
 sg13g2_nand2_2 _3551_ (.Y(_0517_),
    .A(net625),
    .B(\project_audio.iter.x[13] ));
 sg13g2_xor2_1 _3552_ (.B(net627),
    .A(net625),
    .X(_0518_));
 sg13g2_mux2_1 _3553_ (.A0(net625),
    .A1(_0518_),
    .S(_0510_),
    .X(_0519_));
 sg13g2_xnor2_1 _3554_ (.Y(_0520_),
    .A(_0515_),
    .B(_0519_));
 sg13g2_nor2_1 _3555_ (.A(_0513_),
    .B(_0520_),
    .Y(_0521_));
 sg13g2_xor2_1 _3556_ (.B(_0505_),
    .A(_0031_),
    .X(_0522_));
 sg13g2_xor2_1 _3557_ (.B(_0520_),
    .A(_0513_),
    .X(_0523_));
 sg13g2_a21oi_1 _3558_ (.A1(_0522_),
    .A2(_0523_),
    .Y(_0524_),
    .B1(_0521_));
 sg13g2_xor2_1 _3559_ (.B(_0514_),
    .A(_0032_),
    .X(_0525_));
 sg13g2_a21oi_1 _3560_ (.A1(_0515_),
    .A2(_0519_),
    .Y(_0526_),
    .B1(_0516_));
 sg13g2_nand2_2 _3561_ (.Y(_0527_),
    .A(\project_audio.iter.x[11] ),
    .B(\project_audio.iter.x[10] ));
 sg13g2_xor2_1 _3562_ (.B(\project_audio.iter.x[10] ),
    .A(\project_audio.iter.x[11] ),
    .X(_0528_));
 sg13g2_nor2_1 _3563_ (.A(_2453_),
    .B(net625),
    .Y(_0529_));
 sg13g2_nand2_1 _3564_ (.Y(_0530_),
    .A(\project_audio.iter.x[15] ),
    .B(\project_audio.iter.x[13] ));
 sg13g2_xor2_1 _3565_ (.B(net627),
    .A(\project_audio.iter.x[15] ),
    .X(_0531_));
 sg13g2_nor2_1 _3566_ (.A(\project_audio.iter.x[15] ),
    .B(net626),
    .Y(_0532_));
 sg13g2_a21oi_1 _3567_ (.A1(net625),
    .A2(_0531_),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_xnor2_1 _3568_ (.Y(_0534_),
    .A(_0528_),
    .B(_0533_));
 sg13g2_nor2_1 _3569_ (.A(_0526_),
    .B(_0534_),
    .Y(_0535_));
 sg13g2_xor2_1 _3570_ (.B(_0534_),
    .A(_0526_),
    .X(_0536_));
 sg13g2_xnor2_1 _3571_ (.Y(_0537_),
    .A(_0525_),
    .B(_0536_));
 sg13g2_nor2_1 _3572_ (.A(_0524_),
    .B(_0537_),
    .Y(_0538_));
 sg13g2_o21ai_1 _3573_ (.B1(_0030_),
    .Y(_0539_),
    .A1(_0031_),
    .A2(_0505_));
 sg13g2_nor2b_1 _3574_ (.A(_0506_),
    .B_N(_0539_),
    .Y(_0540_));
 sg13g2_xor2_1 _3575_ (.B(_0537_),
    .A(_0524_),
    .X(_0541_));
 sg13g2_a21oi_1 _3576_ (.A1(_0540_),
    .A2(_0541_),
    .Y(_0542_),
    .B1(_0538_));
 sg13g2_nor3_2 _3577_ (.A(_0031_),
    .B(_0032_),
    .C(_0514_),
    .Y(_0543_));
 sg13g2_o21ai_1 _3578_ (.B1(_0031_),
    .Y(_0544_),
    .A1(_0032_),
    .A2(_0514_));
 sg13g2_nand2b_1 _3579_ (.Y(_0545_),
    .B(_0544_),
    .A_N(_0543_));
 sg13g2_inv_1 _3580_ (.Y(_0546_),
    .A(_0545_));
 sg13g2_a21oi_1 _3581_ (.A1(_0525_),
    .A2(_0536_),
    .Y(_0547_),
    .B1(_0535_));
 sg13g2_xor2_1 _3582_ (.B(_0527_),
    .A(_0033_),
    .X(_0548_));
 sg13g2_nor2_1 _3583_ (.A(\project_audio.iter.x[15] ),
    .B(_0517_),
    .Y(_0549_));
 sg13g2_a21oi_1 _3584_ (.A1(_0528_),
    .A2(_0533_),
    .Y(_0550_),
    .B1(_0549_));
 sg13g2_xor2_1 _3585_ (.B(\project_audio.iter.x[11] ),
    .A(net628),
    .X(_0551_));
 sg13g2_xnor2_1 _3586_ (.Y(_0552_),
    .A(_0529_),
    .B(_0551_));
 sg13g2_nor2_1 _3587_ (.A(_0550_),
    .B(_0552_),
    .Y(_0553_));
 sg13g2_xor2_1 _3588_ (.B(_0552_),
    .A(_0550_),
    .X(_0554_));
 sg13g2_xnor2_1 _3589_ (.Y(_0555_),
    .A(_0548_),
    .B(_0554_));
 sg13g2_nor2_1 _3590_ (.A(_0547_),
    .B(_0555_),
    .Y(_0556_));
 sg13g2_xor2_1 _3591_ (.B(_0555_),
    .A(_0547_),
    .X(_0557_));
 sg13g2_xnor2_1 _3592_ (.Y(_0558_),
    .A(_0546_),
    .B(_0557_));
 sg13g2_nor2_1 _3593_ (.A(_0542_),
    .B(_0558_),
    .Y(_0559_));
 sg13g2_xor2_1 _3594_ (.B(_0558_),
    .A(_0542_),
    .X(_0560_));
 sg13g2_xnor2_1 _3595_ (.Y(_0561_),
    .A(_0506_),
    .B(_0560_));
 sg13g2_nor2_1 _3596_ (.A(net628),
    .B(_0527_),
    .Y(_0562_));
 sg13g2_nand2_1 _3597_ (.Y(_0563_),
    .A(\project_audio.iter.x[8] ),
    .B(\project_audio.iter.x[7] ));
 sg13g2_xor2_1 _3598_ (.B(net630),
    .A(\project_audio.iter.x[8] ),
    .X(_0564_));
 sg13g2_mux2_1 _3599_ (.A0(net628),
    .A1(_0551_),
    .S(_0527_),
    .X(_0565_));
 sg13g2_a21oi_1 _3600_ (.A1(_0564_),
    .A2(_0565_),
    .Y(_0566_),
    .B1(_0562_));
 sg13g2_xnor2_1 _3601_ (.Y(_0567_),
    .A(_0509_),
    .B(_0512_));
 sg13g2_nor2_1 _3602_ (.A(_0566_),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_xor2_1 _3603_ (.B(_0567_),
    .A(_0566_),
    .X(_0569_));
 sg13g2_xor2_1 _3604_ (.B(_0563_),
    .A(_0030_),
    .X(_0570_));
 sg13g2_a21oi_1 _3605_ (.A1(_0569_),
    .A2(_0570_),
    .Y(_0571_),
    .B1(_0568_));
 sg13g2_xnor2_1 _3606_ (.Y(_0572_),
    .A(_0522_),
    .B(_0523_));
 sg13g2_nor2_1 _3607_ (.A(_0571_),
    .B(_0572_),
    .Y(_0573_));
 sg13g2_nand3_1 _3608_ (.B(net630),
    .C(\project_audio.iter.x[5] ),
    .A(\project_audio.iter.x[8] ),
    .Y(_0574_));
 sg13g2_nor2_1 _3609_ (.A(_0029_),
    .B(_0574_),
    .Y(_0575_));
 sg13g2_xor2_1 _3610_ (.B(_0574_),
    .A(_0029_),
    .X(_0576_));
 sg13g2_xor2_1 _3611_ (.B(_0572_),
    .A(_0571_),
    .X(_0577_));
 sg13g2_a21oi_1 _3612_ (.A1(_0576_),
    .A2(_0577_),
    .Y(_0578_),
    .B1(_0573_));
 sg13g2_xor2_1 _3613_ (.B(_0541_),
    .A(_0540_),
    .X(_0579_));
 sg13g2_nor2b_1 _3614_ (.A(_0578_),
    .B_N(_0579_),
    .Y(_0580_));
 sg13g2_xnor2_1 _3615_ (.Y(_0581_),
    .A(_0578_),
    .B(_0579_));
 sg13g2_a21oi_1 _3616_ (.A1(_0575_),
    .A2(_0581_),
    .Y(_0582_),
    .B1(_0580_));
 sg13g2_nor2_1 _3617_ (.A(_0561_),
    .B(_0582_),
    .Y(_0583_));
 sg13g2_inv_1 _3618_ (.Y(_0584_),
    .A(_0583_));
 sg13g2_xnor2_1 _3619_ (.Y(_0585_),
    .A(_0561_),
    .B(_0582_));
 sg13g2_inv_1 _3620_ (.Y(_0586_),
    .A(_0585_));
 sg13g2_nand2_2 _3621_ (.Y(_0587_),
    .A(\project_audio.iter.x[4] ),
    .B(net631));
 sg13g2_nor3_2 _3622_ (.A(_0025_),
    .B(_0026_),
    .C(_0587_),
    .Y(_0588_));
 sg13g2_inv_1 _3623_ (.Y(_0589_),
    .A(_0588_));
 sg13g2_o21ai_1 _3624_ (.B1(_0025_),
    .Y(_0590_),
    .A1(_0026_),
    .A2(_0587_));
 sg13g2_nand2_1 _3625_ (.Y(_0591_),
    .A(_0589_),
    .B(_0590_));
 sg13g2_nand2_2 _3626_ (.Y(_0592_),
    .A(net630),
    .B(\project_audio.iter.x[6] ));
 sg13g2_nor2_1 _3627_ (.A(\project_audio.iter.x[8] ),
    .B(_0592_),
    .Y(_0593_));
 sg13g2_mux2_1 _3628_ (.A0(\project_audio.iter.x[8] ),
    .A1(_0564_),
    .S(_0592_),
    .X(_0594_));
 sg13g2_xor2_1 _3629_ (.B(net631),
    .A(\project_audio.iter.x[4] ),
    .X(_0595_));
 sg13g2_a21oi_1 _3630_ (.A1(_0594_),
    .A2(_0595_),
    .Y(_0596_),
    .B1(_0593_));
 sg13g2_nand2_2 _3631_ (.Y(_0597_),
    .A(\project_audio.iter.x[5] ),
    .B(\project_audio.iter.x[4] ));
 sg13g2_xnor2_1 _3632_ (.Y(_0598_),
    .A(\project_audio.iter.x[5] ),
    .B(\project_audio.iter.x[4] ));
 sg13g2_inv_1 _3633_ (.Y(_0599_),
    .A(_0598_));
 sg13g2_nor2_1 _3634_ (.A(\project_audio.iter.x[9] ),
    .B(_0563_),
    .Y(_0600_));
 sg13g2_mux2_1 _3635_ (.A0(\project_audio.iter.x[9] ),
    .A1(_0509_),
    .S(_0563_),
    .X(_0601_));
 sg13g2_xnor2_1 _3636_ (.Y(_0602_),
    .A(_0598_),
    .B(_0601_));
 sg13g2_nand2b_1 _3637_ (.Y(_0603_),
    .B(_0602_),
    .A_N(_0596_));
 sg13g2_xor2_1 _3638_ (.B(_0602_),
    .A(_0596_),
    .X(_0604_));
 sg13g2_xnor2_1 _3639_ (.Y(_0605_),
    .A(_2468_),
    .B(_0587_));
 sg13g2_o21ai_1 _3640_ (.B1(_0603_),
    .Y(_0606_),
    .A1(_0604_),
    .A2(_0605_));
 sg13g2_a21oi_1 _3641_ (.A1(_0599_),
    .A2(_0601_),
    .Y(_0607_),
    .B1(_0600_));
 sg13g2_nand2_2 _3642_ (.Y(_0608_),
    .A(\project_audio.iter.x[6] ),
    .B(\project_audio.iter.x[5] ));
 sg13g2_xor2_1 _3643_ (.B(\project_audio.iter.x[5] ),
    .A(\project_audio.iter.x[6] ),
    .X(_0609_));
 sg13g2_nor2_1 _3644_ (.A(\project_audio.iter.x[10] ),
    .B(_0505_),
    .Y(_0610_));
 sg13g2_mux2_1 _3645_ (.A0(\project_audio.iter.x[10] ),
    .A1(_0515_),
    .S(_0505_),
    .X(_0611_));
 sg13g2_xor2_1 _3646_ (.B(_0611_),
    .A(_0609_),
    .X(_0612_));
 sg13g2_nand2b_1 _3647_ (.Y(_0613_),
    .B(_0612_),
    .A_N(_0607_));
 sg13g2_nor2b_1 _3648_ (.A(_0612_),
    .B_N(_0607_),
    .Y(_0614_));
 sg13g2_xnor2_1 _3649_ (.Y(_0615_),
    .A(_0607_),
    .B(_0612_));
 sg13g2_xnor2_1 _3650_ (.Y(_0616_),
    .A(_2467_),
    .B(_0597_));
 sg13g2_xnor2_1 _3651_ (.Y(_0617_),
    .A(_0615_),
    .B(_0616_));
 sg13g2_nand2_1 _3652_ (.Y(_0618_),
    .A(_0606_),
    .B(_0617_));
 sg13g2_xnor2_1 _3653_ (.Y(_0619_),
    .A(_0606_),
    .B(_0617_));
 sg13g2_xor2_1 _3654_ (.B(_0619_),
    .A(_0591_),
    .X(_0620_));
 sg13g2_nor2_1 _3655_ (.A(net630),
    .B(_0608_),
    .Y(_0621_));
 sg13g2_xor2_1 _3656_ (.B(\project_audio.iter.x[6] ),
    .A(net630),
    .X(_0622_));
 sg13g2_mux2_1 _3657_ (.A0(net630),
    .A1(_0622_),
    .S(_0608_),
    .X(_0623_));
 sg13g2_nand2_2 _3658_ (.Y(_0624_),
    .A(net631),
    .B(\project_audio.iter.x[2] ));
 sg13g2_xor2_1 _3659_ (.B(\project_audio.iter.x[2] ),
    .A(net631),
    .X(_0625_));
 sg13g2_a21oi_1 _3660_ (.A1(_0623_),
    .A2(_0625_),
    .Y(_0626_),
    .B1(_0621_));
 sg13g2_xnor2_1 _3661_ (.Y(_0627_),
    .A(_0594_),
    .B(_0595_));
 sg13g2_nor2_1 _3662_ (.A(_0626_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nor2_1 _3663_ (.A(_0025_),
    .B(_0624_),
    .Y(_0629_));
 sg13g2_xor2_1 _3664_ (.B(_0624_),
    .A(_0025_),
    .X(_0630_));
 sg13g2_xor2_1 _3665_ (.B(_0627_),
    .A(_0626_),
    .X(_0631_));
 sg13g2_a21oi_1 _3666_ (.A1(_0630_),
    .A2(_0631_),
    .Y(_0632_),
    .B1(_0628_));
 sg13g2_xnor2_1 _3667_ (.Y(_0633_),
    .A(_0604_),
    .B(_0605_));
 sg13g2_nor2_1 _3668_ (.A(_0632_),
    .B(_0633_),
    .Y(_0634_));
 sg13g2_xor2_1 _3669_ (.B(_0633_),
    .A(_0632_),
    .X(_0635_));
 sg13g2_a21oi_1 _3670_ (.A1(_0629_),
    .A2(_0635_),
    .Y(_0636_),
    .B1(_0634_));
 sg13g2_nor2b_1 _3671_ (.A(_0636_),
    .B_N(_0620_),
    .Y(_0637_));
 sg13g2_o21ai_1 _3672_ (.B1(_0618_),
    .Y(_0638_),
    .A1(_0591_),
    .A2(_0619_));
 sg13g2_nor3_1 _3673_ (.A(_0026_),
    .B(_0027_),
    .C(_0597_),
    .Y(_0639_));
 sg13g2_inv_1 _3674_ (.Y(_0640_),
    .A(_0639_));
 sg13g2_o21ai_1 _3675_ (.B1(_0026_),
    .Y(_0641_),
    .A1(_0027_),
    .A2(_0597_));
 sg13g2_nand2_1 _3676_ (.Y(_0642_),
    .A(_0640_),
    .B(_0641_));
 sg13g2_o21ai_1 _3677_ (.B1(_0613_),
    .Y(_0643_),
    .A1(_0614_),
    .A2(_0616_));
 sg13g2_a21oi_1 _3678_ (.A1(_0609_),
    .A2(_0611_),
    .Y(_0644_),
    .B1(_0610_));
 sg13g2_nor2_1 _3679_ (.A(\project_audio.iter.x[11] ),
    .B(_0514_),
    .Y(_0645_));
 sg13g2_mux2_1 _3680_ (.A0(\project_audio.iter.x[11] ),
    .A1(_0528_),
    .S(_0514_),
    .X(_0646_));
 sg13g2_xor2_1 _3681_ (.B(_0646_),
    .A(_0622_),
    .X(_0647_));
 sg13g2_nand2b_1 _3682_ (.Y(_0648_),
    .B(_0647_),
    .A_N(_0644_));
 sg13g2_nor2b_1 _3683_ (.A(_0647_),
    .B_N(_0644_),
    .Y(_0649_));
 sg13g2_xnor2_1 _3684_ (.Y(_0650_),
    .A(_0644_),
    .B(_0647_));
 sg13g2_xnor2_1 _3685_ (.Y(_0651_),
    .A(_2466_),
    .B(_0608_));
 sg13g2_xnor2_1 _3686_ (.Y(_0652_),
    .A(_0650_),
    .B(_0651_));
 sg13g2_nand2_1 _3687_ (.Y(_0653_),
    .A(_0643_),
    .B(_0652_));
 sg13g2_xnor2_1 _3688_ (.Y(_0654_),
    .A(_0643_),
    .B(_0652_));
 sg13g2_xor2_1 _3689_ (.B(_0654_),
    .A(_0642_),
    .X(_0655_));
 sg13g2_nand2_1 _3690_ (.Y(_0656_),
    .A(_0638_),
    .B(_0655_));
 sg13g2_xnor2_1 _3691_ (.Y(_0657_),
    .A(_0638_),
    .B(_0655_));
 sg13g2_xnor2_1 _3692_ (.Y(_0658_),
    .A(_0588_),
    .B(_0657_));
 sg13g2_nor2_1 _3693_ (.A(_0637_),
    .B(_0658_),
    .Y(_0659_));
 sg13g2_nor2_1 _3694_ (.A(\project_audio.iter.x[5] ),
    .B(_0587_),
    .Y(_0660_));
 sg13g2_nand2_1 _3695_ (.Y(_0661_),
    .A(_0587_),
    .B(_0598_));
 sg13g2_nand2b_1 _3696_ (.Y(_0662_),
    .B(_0661_),
    .A_N(_0660_));
 sg13g2_nand2_2 _3697_ (.Y(_0663_),
    .A(\project_audio.iter.x[1] ),
    .B(\project_audio.iter.x[0] ));
 sg13g2_inv_1 _3698_ (.Y(_0664_),
    .A(_0663_));
 sg13g2_xor2_1 _3699_ (.B(\project_audio.iter.x[0] ),
    .A(\project_audio.iter.x[1] ),
    .X(_0665_));
 sg13g2_a21oi_1 _3700_ (.A1(_0661_),
    .A2(_0665_),
    .Y(_0666_),
    .B1(_0660_));
 sg13g2_nor2_1 _3701_ (.A(\project_audio.iter.x[6] ),
    .B(_0597_),
    .Y(_0667_));
 sg13g2_mux2_1 _3702_ (.A0(\project_audio.iter.x[6] ),
    .A1(_0609_),
    .S(_0597_),
    .X(_0668_));
 sg13g2_nand2_2 _3703_ (.Y(_0669_),
    .A(\project_audio.iter.x[2] ),
    .B(\project_audio.iter.x[1] ));
 sg13g2_inv_1 _3704_ (.Y(_0670_),
    .A(_0669_));
 sg13g2_xor2_1 _3705_ (.B(\project_audio.iter.x[1] ),
    .A(\project_audio.iter.x[2] ),
    .X(_0671_));
 sg13g2_xnor2_1 _3706_ (.Y(_0672_),
    .A(_0668_),
    .B(_0671_));
 sg13g2_nor2_1 _3707_ (.A(_0666_),
    .B(_0672_),
    .Y(_0673_));
 sg13g2_xor2_1 _3708_ (.B(_0672_),
    .A(_0666_),
    .X(_0674_));
 sg13g2_a21oi_2 _3709_ (.B1(_0673_),
    .Y(_0675_),
    .A2(_0674_),
    .A1(_0664_));
 sg13g2_a21oi_1 _3710_ (.A1(_0668_),
    .A2(_0671_),
    .Y(_0676_),
    .B1(_0667_));
 sg13g2_xnor2_1 _3711_ (.Y(_0677_),
    .A(_0623_),
    .B(_0625_));
 sg13g2_nor2_1 _3712_ (.A(_0676_),
    .B(_0677_),
    .Y(_0678_));
 sg13g2_xor2_1 _3713_ (.B(_0677_),
    .A(_0676_),
    .X(_0679_));
 sg13g2_xnor2_1 _3714_ (.Y(_0680_),
    .A(_0670_),
    .B(_0679_));
 sg13g2_nor2_1 _3715_ (.A(_0675_),
    .B(_0680_),
    .Y(_0681_));
 sg13g2_xnor2_1 _3716_ (.Y(_0682_),
    .A(_0630_),
    .B(_0631_));
 sg13g2_a21oi_2 _3717_ (.B1(_0678_),
    .Y(_0683_),
    .A2(_0679_),
    .A1(_0670_));
 sg13g2_nor2_1 _3718_ (.A(_0682_),
    .B(_0683_),
    .Y(_0684_));
 sg13g2_xnor2_1 _3719_ (.Y(_0685_),
    .A(_0682_),
    .B(_0683_));
 sg13g2_or3_1 _3720_ (.A(_0675_),
    .B(_0680_),
    .C(_0685_),
    .X(_0686_));
 sg13g2_xnor2_1 _3721_ (.Y(_0687_),
    .A(_0629_),
    .B(_0635_));
 sg13g2_xor2_1 _3722_ (.B(_0687_),
    .A(_0684_),
    .X(_0688_));
 sg13g2_or2_1 _3723_ (.X(_0689_),
    .B(_0688_),
    .A(_0686_));
 sg13g2_xnor2_1 _3724_ (.Y(_0690_),
    .A(_0686_),
    .B(_0688_));
 sg13g2_xnor2_1 _3725_ (.Y(_0691_),
    .A(_0663_),
    .B(_0674_));
 sg13g2_mux2_1 _3726_ (.A0(_0675_),
    .A1(_0673_),
    .S(_0680_),
    .X(_0692_));
 sg13g2_xor2_1 _3727_ (.B(_0665_),
    .A(_0662_),
    .X(_0693_));
 sg13g2_nor2_1 _3728_ (.A(\project_audio.iter.x[4] ),
    .B(_0624_),
    .Y(_0694_));
 sg13g2_nor2b_1 _3729_ (.A(_0595_),
    .B_N(_0624_),
    .Y(_0695_));
 sg13g2_nor2_1 _3730_ (.A(_0694_),
    .B(_0695_),
    .Y(_0696_));
 sg13g2_a21oi_1 _3731_ (.A1(\project_audio.iter.x[0] ),
    .A2(_0696_),
    .Y(_0697_),
    .B1(_0694_));
 sg13g2_nor2_1 _3732_ (.A(_0693_),
    .B(_0697_),
    .Y(_0698_));
 sg13g2_nand3_1 _3733_ (.B(_0692_),
    .C(_0698_),
    .A(_0691_),
    .Y(_0699_));
 sg13g2_xor2_1 _3734_ (.B(_0685_),
    .A(_0681_),
    .X(_0700_));
 sg13g2_nor2_1 _3735_ (.A(_0699_),
    .B(_0700_),
    .Y(_0701_));
 sg13g2_xnor2_1 _3736_ (.Y(_0702_),
    .A(\project_audio.iter.x[0] ),
    .B(_0696_));
 sg13g2_nor3_1 _3737_ (.A(net631),
    .B(_0669_),
    .C(_0702_),
    .Y(_0703_));
 sg13g2_nand3_1 _3738_ (.B(_0692_),
    .C(_0703_),
    .A(_0691_),
    .Y(_0704_));
 sg13g2_o21ai_1 _3739_ (.B1(_0702_),
    .Y(_0705_),
    .A1(net631),
    .A2(_0669_));
 sg13g2_nor2_1 _3740_ (.A(\project_audio.iter.x[2] ),
    .B(_0663_),
    .Y(_0706_));
 sg13g2_nor4_1 _3741_ (.A(_2466_),
    .B(\project_audio.iter.x[2] ),
    .C(_0663_),
    .D(_0702_),
    .Y(_0707_));
 sg13g2_nand2b_1 _3742_ (.Y(_0708_),
    .B(_0707_),
    .A_N(_0592_));
 sg13g2_xnor2_1 _3743_ (.Y(_0709_),
    .A(_0693_),
    .B(_0697_));
 sg13g2_a21oi_1 _3744_ (.A1(_0704_),
    .A2(_0708_),
    .Y(_0710_),
    .B1(_0709_));
 sg13g2_xor2_1 _3745_ (.B(_0700_),
    .A(_0699_),
    .X(_0711_));
 sg13g2_a21oi_1 _3746_ (.A1(_0710_),
    .A2(_0711_),
    .Y(_0712_),
    .B1(_0701_));
 sg13g2_or2_1 _3747_ (.X(_0713_),
    .B(_0712_),
    .A(_0690_));
 sg13g2_o21ai_1 _3748_ (.B1(_0689_),
    .Y(_0714_),
    .A1(_0690_),
    .A2(_0712_));
 sg13g2_xor2_1 _3749_ (.B(_0636_),
    .A(_0620_),
    .X(_0715_));
 sg13g2_inv_1 _3750_ (.Y(_0716_),
    .A(_0715_));
 sg13g2_nor4_1 _3751_ (.A(_0682_),
    .B(_0683_),
    .C(_0687_),
    .D(_0715_),
    .Y(_0717_));
 sg13g2_a221oi_1 _3752_ (.B2(_0620_),
    .C1(_0717_),
    .B1(_0714_),
    .A1(_0637_),
    .Y(_0718_),
    .A2(_0658_));
 sg13g2_xor2_1 _3753_ (.B(_0658_),
    .A(_0637_),
    .X(_0719_));
 sg13g2_o21ai_1 _3754_ (.B1(_0648_),
    .Y(_0720_),
    .A1(_0649_),
    .A2(_0651_));
 sg13g2_nand3_1 _3755_ (.B(\project_audio.iter.x[6] ),
    .C(\project_audio.iter.x[4] ),
    .A(net630),
    .Y(_0721_));
 sg13g2_xnor2_1 _3756_ (.Y(_0722_),
    .A(_2465_),
    .B(_0592_));
 sg13g2_a21oi_1 _3757_ (.A1(_0622_),
    .A2(_0646_),
    .Y(_0723_),
    .B1(_0645_));
 sg13g2_xor2_1 _3758_ (.B(_0565_),
    .A(_0564_),
    .X(_0724_));
 sg13g2_nand2b_1 _3759_ (.Y(_0725_),
    .B(_0724_),
    .A_N(_0723_));
 sg13g2_nor2b_1 _3760_ (.A(_0724_),
    .B_N(_0723_),
    .Y(_0726_));
 sg13g2_xnor2_1 _3761_ (.Y(_0727_),
    .A(_0723_),
    .B(_0724_));
 sg13g2_xnor2_1 _3762_ (.Y(_0728_),
    .A(_0722_),
    .B(_0727_));
 sg13g2_nand2_1 _3763_ (.Y(_0729_),
    .A(_0720_),
    .B(_0728_));
 sg13g2_nor3_1 _3764_ (.A(_0027_),
    .B(_0028_),
    .C(_0608_),
    .Y(_0730_));
 sg13g2_inv_1 _3765_ (.Y(_0731_),
    .A(_0730_));
 sg13g2_o21ai_1 _3766_ (.B1(_0027_),
    .Y(_0732_),
    .A1(_0028_),
    .A2(_0608_));
 sg13g2_nand2_1 _3767_ (.Y(_0733_),
    .A(_0731_),
    .B(_0732_));
 sg13g2_xnor2_1 _3768_ (.Y(_0734_),
    .A(_0720_),
    .B(_0728_));
 sg13g2_o21ai_1 _3769_ (.B1(_0729_),
    .Y(_0735_),
    .A1(_0733_),
    .A2(_0734_));
 sg13g2_nor2_1 _3770_ (.A(_0028_),
    .B(_0721_),
    .Y(_0736_));
 sg13g2_xor2_1 _3771_ (.B(_0721_),
    .A(_0028_),
    .X(_0737_));
 sg13g2_o21ai_1 _3772_ (.B1(_0725_),
    .Y(_0738_),
    .A1(_0722_),
    .A2(_0726_));
 sg13g2_xor2_1 _3773_ (.B(_0570_),
    .A(_0569_),
    .X(_0739_));
 sg13g2_and2_1 _3774_ (.A(_0738_),
    .B(_0739_),
    .X(_0740_));
 sg13g2_or2_1 _3775_ (.X(_0741_),
    .B(_0739_),
    .A(_0738_));
 sg13g2_xor2_1 _3776_ (.B(_0739_),
    .A(_0738_),
    .X(_0742_));
 sg13g2_xnor2_1 _3777_ (.Y(_0743_),
    .A(_0737_),
    .B(_0742_));
 sg13g2_nand2b_1 _3778_ (.Y(_0744_),
    .B(_0735_),
    .A_N(_0743_));
 sg13g2_xor2_1 _3779_ (.B(_0743_),
    .A(_0735_),
    .X(_0745_));
 sg13g2_or2_1 _3780_ (.X(_0746_),
    .B(_0745_),
    .A(_0731_));
 sg13g2_a21oi_1 _3781_ (.A1(_0737_),
    .A2(_0741_),
    .Y(_0747_),
    .B1(_0740_));
 sg13g2_xnor2_1 _3782_ (.Y(_0748_),
    .A(_0576_),
    .B(_0577_));
 sg13g2_nor2_1 _3783_ (.A(_0747_),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_xor2_1 _3784_ (.B(_0748_),
    .A(_0747_),
    .X(_0750_));
 sg13g2_xnor2_1 _3785_ (.Y(_0751_),
    .A(_0736_),
    .B(_0750_));
 sg13g2_a21oi_1 _3786_ (.A1(_0744_),
    .A2(_0746_),
    .Y(_0752_),
    .B1(_0751_));
 sg13g2_a21o_1 _3787_ (.A2(_0746_),
    .A1(_0744_),
    .B1(_0751_),
    .X(_0753_));
 sg13g2_a21oi_2 _3788_ (.B1(_0749_),
    .Y(_0754_),
    .A2(_0750_),
    .A1(_0736_));
 sg13g2_xnor2_1 _3789_ (.Y(_0755_),
    .A(_0575_),
    .B(_0581_));
 sg13g2_nor2_1 _3790_ (.A(_0754_),
    .B(_0755_),
    .Y(_0756_));
 sg13g2_nand2_1 _3791_ (.Y(_0757_),
    .A(_0754_),
    .B(_0755_));
 sg13g2_xor2_1 _3792_ (.B(_0755_),
    .A(_0754_),
    .X(_0758_));
 sg13g2_nand2b_1 _3793_ (.Y(_0759_),
    .B(_0757_),
    .A_N(_0756_));
 sg13g2_nand3_1 _3794_ (.B(_0746_),
    .C(_0751_),
    .A(_0744_),
    .Y(_0760_));
 sg13g2_nand2_1 _3795_ (.Y(_0761_),
    .A(_0758_),
    .B(_0760_));
 sg13g2_and3_1 _3796_ (.X(_0762_),
    .A(_0753_),
    .B(_0758_),
    .C(_0760_));
 sg13g2_nand3_1 _3797_ (.B(_0758_),
    .C(_0760_),
    .A(_0753_),
    .Y(_0763_));
 sg13g2_o21ai_1 _3798_ (.B1(_0656_),
    .Y(_0764_),
    .A1(_0589_),
    .A2(_0657_));
 sg13g2_o21ai_1 _3799_ (.B1(_0653_),
    .Y(_0765_),
    .A1(_0642_),
    .A2(_0654_));
 sg13g2_xor2_1 _3800_ (.B(_0734_),
    .A(_0733_),
    .X(_0766_));
 sg13g2_nand2_1 _3801_ (.Y(_0767_),
    .A(_0765_),
    .B(_0766_));
 sg13g2_xnor2_1 _3802_ (.Y(_0768_),
    .A(_0765_),
    .B(_0766_));
 sg13g2_xnor2_1 _3803_ (.Y(_0769_),
    .A(_0639_),
    .B(_0768_));
 sg13g2_nand2_1 _3804_ (.Y(_0770_),
    .A(_0764_),
    .B(_0769_));
 sg13g2_nor2_1 _3805_ (.A(_0764_),
    .B(_0769_),
    .Y(_0771_));
 sg13g2_or2_1 _3806_ (.X(_0772_),
    .B(_0769_),
    .A(_0764_));
 sg13g2_xnor2_1 _3807_ (.Y(_0773_),
    .A(_0731_),
    .B(_0745_));
 sg13g2_o21ai_1 _3808_ (.B1(_0767_),
    .Y(_0774_),
    .A1(_0640_),
    .A2(_0768_));
 sg13g2_nor2b_1 _3809_ (.A(_0774_),
    .B_N(_0773_),
    .Y(_0775_));
 sg13g2_nand2b_1 _3810_ (.Y(_0776_),
    .B(_0774_),
    .A_N(_0773_));
 sg13g2_xnor2_1 _3811_ (.Y(_0777_),
    .A(_0773_),
    .B(_0774_));
 sg13g2_nand3_1 _3812_ (.B(_0772_),
    .C(_0777_),
    .A(_0770_),
    .Y(_0778_));
 sg13g2_nor4_2 _3813_ (.A(_0659_),
    .B(_0718_),
    .C(_0763_),
    .Y(_0779_),
    .D(_0778_));
 sg13g2_or4_1 _3814_ (.A(_0659_),
    .B(_0718_),
    .C(_0763_),
    .D(_0778_),
    .X(_0780_));
 sg13g2_a21o_1 _3815_ (.A2(_0776_),
    .A1(_0770_),
    .B1(_0775_),
    .X(_0781_));
 sg13g2_a21oi_1 _3816_ (.A1(_0770_),
    .A2(_0776_),
    .Y(_0782_),
    .B1(_0775_));
 sg13g2_o21ai_1 _3817_ (.B1(_0757_),
    .Y(_0783_),
    .A1(_0752_),
    .A2(_0756_));
 sg13g2_a221oi_1 _3818_ (.B2(_0782_),
    .C1(_0756_),
    .B1(_0762_),
    .A1(_0752_),
    .Y(_0784_),
    .A2(_0757_));
 sg13g2_o21ai_1 _3819_ (.B1(_0783_),
    .Y(_0785_),
    .A1(_0763_),
    .A2(_0781_));
 sg13g2_nor3_1 _3820_ (.A(_0586_),
    .B(_0779_),
    .C(_0785_),
    .Y(_0786_));
 sg13g2_a21oi_1 _3821_ (.A1(_0780_),
    .A2(_0784_),
    .Y(_0787_),
    .B1(_0585_));
 sg13g2_o21ai_1 _3822_ (.B1(_0586_),
    .Y(_0788_),
    .A1(_0779_),
    .A2(_0785_));
 sg13g2_a21o_1 _3823_ (.A2(_0781_),
    .A1(_0753_),
    .B1(_0761_),
    .X(_0789_));
 sg13g2_a21oi_1 _3824_ (.A1(_0620_),
    .A2(_0714_),
    .Y(_0790_),
    .B1(_0717_));
 sg13g2_xnor2_1 _3825_ (.Y(_0791_),
    .A(_0719_),
    .B(_0790_));
 sg13g2_o21ai_1 _3826_ (.B1(_0771_),
    .Y(_0792_),
    .A1(_0659_),
    .A2(_0718_));
 sg13g2_xnor2_1 _3827_ (.Y(_0793_),
    .A(_0710_),
    .B(_0711_));
 sg13g2_nand2_1 _3828_ (.Y(_0794_),
    .A(_0665_),
    .B(_0671_));
 sg13g2_mux2_1 _3829_ (.A0(net631),
    .A1(_0625_),
    .S(_0669_),
    .X(_0795_));
 sg13g2_nor2_1 _3830_ (.A(_0706_),
    .B(_0795_),
    .Y(_0796_));
 sg13g2_a21oi_1 _3831_ (.A1(net631),
    .A2(_0706_),
    .Y(_0797_),
    .B1(_0796_));
 sg13g2_nand3b_1 _3832_ (.B(_0705_),
    .C(_0797_),
    .Y(_0798_),
    .A_N(_0703_));
 sg13g2_o21ai_1 _3833_ (.B1(_0798_),
    .Y(_0799_),
    .A1(_0702_),
    .A2(_0794_));
 sg13g2_nor2_1 _3834_ (.A(net630),
    .B(_0709_),
    .Y(_0800_));
 sg13g2_nand3_1 _3835_ (.B(_0799_),
    .C(_0800_),
    .A(_0691_),
    .Y(_0801_));
 sg13g2_a22oi_1 _3836_ (.Y(_0802_),
    .B1(_0793_),
    .B2(_0801_),
    .A2(_0712_),
    .A1(_0690_));
 sg13g2_nand4_1 _3837_ (.B(_0716_),
    .C(_0777_),
    .A(_0713_),
    .Y(_0803_),
    .D(_0802_));
 sg13g2_a221oi_1 _3838_ (.B2(_0781_),
    .C1(_0803_),
    .B1(_0761_),
    .A1(_0753_),
    .Y(_0804_),
    .A2(_0759_));
 sg13g2_nand4_1 _3839_ (.B(_0791_),
    .C(_0792_),
    .A(_0789_),
    .Y(_0805_),
    .D(_0804_));
 sg13g2_nor3_2 _3840_ (.A(_0786_),
    .B(_0787_),
    .C(_0805_),
    .Y(_0806_));
 sg13g2_o21ai_1 _3841_ (.B1(_0805_),
    .Y(_0807_),
    .A1(_0786_),
    .A2(_0787_));
 sg13g2_nand2b_2 _3842_ (.Y(_0808_),
    .B(_0807_),
    .A_N(_0806_));
 sg13g2_o21ai_1 _3843_ (.B1(_0504_),
    .Y(_0061_),
    .A1(net615),
    .A2(_0808_));
 sg13g2_nand2_1 _3844_ (.Y(_0809_),
    .A(net718),
    .B(net614));
 sg13g2_a21oi_1 _3845_ (.A1(_0546_),
    .A2(_0557_),
    .Y(_0810_),
    .B1(_0556_));
 sg13g2_nor3_2 _3846_ (.A(_0032_),
    .B(_0033_),
    .C(_0527_),
    .Y(_0811_));
 sg13g2_o21ai_1 _3847_ (.B1(_0032_),
    .Y(_0812_),
    .A1(_0033_),
    .A2(_0527_));
 sg13g2_nand2b_1 _3848_ (.Y(_0813_),
    .B(_0812_),
    .A_N(_0811_));
 sg13g2_a21oi_1 _3849_ (.A1(_0548_),
    .A2(_0554_),
    .Y(_0814_),
    .B1(_0553_));
 sg13g2_nand2_1 _3850_ (.Y(_0815_),
    .A(\project_audio.iter.x[15] ),
    .B(net626));
 sg13g2_o21ai_1 _3851_ (.B1(\project_audio.iter.x[15] ),
    .Y(_0816_),
    .A1(net625),
    .A2(_0551_));
 sg13g2_nor2b_1 _3852_ (.A(_0816_),
    .B_N(_0511_),
    .Y(_0817_));
 sg13g2_xnor2_1 _3853_ (.Y(_0818_),
    .A(_0511_),
    .B(_0816_));
 sg13g2_xor2_1 _3854_ (.B(_0507_),
    .A(_0034_),
    .X(_0819_));
 sg13g2_xnor2_1 _3855_ (.Y(_0820_),
    .A(_0818_),
    .B(_0819_));
 sg13g2_nor2_1 _3856_ (.A(_0814_),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_xnor2_1 _3857_ (.Y(_0822_),
    .A(_0814_),
    .B(_0820_));
 sg13g2_nor2_1 _3858_ (.A(_0813_),
    .B(_0822_),
    .Y(_0823_));
 sg13g2_xor2_1 _3859_ (.B(_0822_),
    .A(_0813_),
    .X(_0824_));
 sg13g2_nand2b_1 _3860_ (.Y(_0825_),
    .B(_0824_),
    .A_N(_0810_));
 sg13g2_xnor2_1 _3861_ (.Y(_0826_),
    .A(_0810_),
    .B(_0824_));
 sg13g2_nand2_1 _3862_ (.Y(_0827_),
    .A(_0543_),
    .B(_0826_));
 sg13g2_xnor2_1 _3863_ (.Y(_0828_),
    .A(_0543_),
    .B(_0826_));
 sg13g2_a21oi_2 _3864_ (.B1(_0559_),
    .Y(_0829_),
    .A2(_0560_),
    .A1(_0506_));
 sg13g2_nand2_1 _3865_ (.Y(_0830_),
    .A(_0828_),
    .B(_0829_));
 sg13g2_nor2_1 _3866_ (.A(_0828_),
    .B(_0829_),
    .Y(_0831_));
 sg13g2_xnor2_1 _3867_ (.Y(_0832_),
    .A(_0828_),
    .B(_0829_));
 sg13g2_a21o_1 _3868_ (.A2(_0788_),
    .A1(_0584_),
    .B1(_0832_),
    .X(_0833_));
 sg13g2_nand3_1 _3869_ (.B(_0788_),
    .C(_0832_),
    .A(_0584_),
    .Y(_0834_));
 sg13g2_and2_1 _3870_ (.A(_0833_),
    .B(_0834_),
    .X(_0835_));
 sg13g2_nand3_1 _3871_ (.B(_0833_),
    .C(_0834_),
    .A(_0806_),
    .Y(_0836_));
 sg13g2_xnor2_1 _3872_ (.Y(_0837_),
    .A(_0806_),
    .B(_0835_));
 sg13g2_o21ai_1 _3873_ (.B1(_0809_),
    .Y(_0062_),
    .A1(_0502_),
    .A2(_0837_));
 sg13g2_nand2_1 _3874_ (.Y(_0838_),
    .A(net754),
    .B(net613));
 sg13g2_nor3_2 _3875_ (.A(_0033_),
    .B(_0034_),
    .C(_0507_),
    .Y(_0839_));
 sg13g2_o21ai_1 _3876_ (.B1(_0033_),
    .Y(_0840_),
    .A1(_0034_),
    .A2(_0507_));
 sg13g2_nand2b_1 _3877_ (.Y(_0841_),
    .B(_0840_),
    .A_N(_0839_));
 sg13g2_xor2_1 _3878_ (.B(_0510_),
    .A(_0035_),
    .X(_0842_));
 sg13g2_nand2_1 _3879_ (.Y(_0843_),
    .A(_0518_),
    .B(_0842_));
 sg13g2_xnor2_1 _3880_ (.Y(_0844_),
    .A(_0518_),
    .B(_0842_));
 sg13g2_a21oi_1 _3881_ (.A1(_0818_),
    .A2(_0819_),
    .Y(_0845_),
    .B1(_0817_));
 sg13g2_xor2_1 _3882_ (.B(_0845_),
    .A(_0844_),
    .X(_0846_));
 sg13g2_nand2b_1 _3883_ (.Y(_0847_),
    .B(_0846_),
    .A_N(_0841_));
 sg13g2_xnor2_1 _3884_ (.Y(_0848_),
    .A(_0841_),
    .B(_0846_));
 sg13g2_o21ai_1 _3885_ (.B1(_0848_),
    .Y(_0849_),
    .A1(_0821_),
    .A2(_0823_));
 sg13g2_or3_1 _3886_ (.A(_0821_),
    .B(_0823_),
    .C(_0848_),
    .X(_0850_));
 sg13g2_and2_1 _3887_ (.A(_0849_),
    .B(_0850_),
    .X(_0851_));
 sg13g2_nand2_1 _3888_ (.Y(_0852_),
    .A(_0811_),
    .B(_0851_));
 sg13g2_xnor2_1 _3889_ (.Y(_0853_),
    .A(_0811_),
    .B(_0851_));
 sg13g2_a21oi_1 _3890_ (.A1(_0825_),
    .A2(_0827_),
    .Y(_0854_),
    .B1(_0853_));
 sg13g2_inv_1 _3891_ (.Y(_0855_),
    .A(_0854_));
 sg13g2_nand3_1 _3892_ (.B(_0827_),
    .C(_0853_),
    .A(_0825_),
    .Y(_0856_));
 sg13g2_nor2b_1 _3893_ (.A(_0854_),
    .B_N(_0856_),
    .Y(_0857_));
 sg13g2_or2_1 _3894_ (.X(_0858_),
    .B(_0832_),
    .A(_0585_));
 sg13g2_a21oi_1 _3895_ (.A1(_0780_),
    .A2(_0784_),
    .Y(_0859_),
    .B1(_0858_));
 sg13g2_a21o_1 _3896_ (.A2(_0784_),
    .A1(_0780_),
    .B1(_0858_),
    .X(_0860_));
 sg13g2_o21ai_1 _3897_ (.B1(_0830_),
    .Y(_0861_),
    .A1(_0583_),
    .A2(_0831_));
 sg13g2_inv_1 _3898_ (.Y(_0862_),
    .A(_0861_));
 sg13g2_nor3_1 _3899_ (.A(_0857_),
    .B(_0859_),
    .C(_0862_),
    .Y(_0863_));
 sg13g2_o21ai_1 _3900_ (.B1(_0857_),
    .Y(_0864_),
    .A1(_0859_),
    .A2(_0862_));
 sg13g2_nand2b_2 _3901_ (.Y(_0865_),
    .B(_0864_),
    .A_N(_0863_));
 sg13g2_xnor2_1 _3902_ (.Y(_0866_),
    .A(_0836_),
    .B(_0865_));
 sg13g2_o21ai_1 _3903_ (.B1(_0838_),
    .Y(_0063_),
    .A1(_0502_),
    .A2(_0866_));
 sg13g2_nand2_1 _3904_ (.Y(_0867_),
    .A(net729),
    .B(net613));
 sg13g2_o21ai_1 _3905_ (.B1(_0847_),
    .Y(_0868_),
    .A1(_0844_),
    .A2(_0845_));
 sg13g2_nor3_2 _3906_ (.A(_0034_),
    .B(_0035_),
    .C(_0510_),
    .Y(_0869_));
 sg13g2_o21ai_1 _3907_ (.B1(_0034_),
    .Y(_0870_),
    .A1(_0035_),
    .A2(_0510_));
 sg13g2_nand2b_1 _3908_ (.Y(_0871_),
    .B(_0870_),
    .A_N(_0869_));
 sg13g2_nand2b_1 _3909_ (.Y(_0872_),
    .B(_0815_),
    .A_N(_0532_));
 sg13g2_xor2_1 _3910_ (.B(_0517_),
    .A(_0036_),
    .X(_0873_));
 sg13g2_nand2b_1 _3911_ (.Y(_0874_),
    .B(_0873_),
    .A_N(_0872_));
 sg13g2_xor2_1 _3912_ (.B(_0873_),
    .A(_0872_),
    .X(_0875_));
 sg13g2_xor2_1 _3913_ (.B(_0875_),
    .A(_0843_),
    .X(_0876_));
 sg13g2_nand2b_1 _3914_ (.Y(_0877_),
    .B(_0876_),
    .A_N(_0871_));
 sg13g2_xnor2_1 _3915_ (.Y(_0878_),
    .A(_0871_),
    .B(_0876_));
 sg13g2_nand2_1 _3916_ (.Y(_0879_),
    .A(_0868_),
    .B(_0878_));
 sg13g2_xor2_1 _3917_ (.B(_0878_),
    .A(_0868_),
    .X(_0880_));
 sg13g2_nand2_1 _3918_ (.Y(_0881_),
    .A(_0839_),
    .B(_0880_));
 sg13g2_xnor2_1 _3919_ (.Y(_0882_),
    .A(_0839_),
    .B(_0880_));
 sg13g2_a21o_1 _3920_ (.A2(_0852_),
    .A1(_0849_),
    .B1(_0882_),
    .X(_0883_));
 sg13g2_nand3_1 _3921_ (.B(_0852_),
    .C(_0882_),
    .A(_0849_),
    .Y(_0884_));
 sg13g2_and2_1 _3922_ (.A(_0883_),
    .B(_0884_),
    .X(_0885_));
 sg13g2_inv_1 _3923_ (.Y(_0886_),
    .A(_0885_));
 sg13g2_and3_1 _3924_ (.X(_0887_),
    .A(_0855_),
    .B(_0864_),
    .C(_0886_));
 sg13g2_a21oi_1 _3925_ (.A1(_0855_),
    .A2(_0864_),
    .Y(_0888_),
    .B1(_0886_));
 sg13g2_or2_1 _3926_ (.X(_0889_),
    .B(_0888_),
    .A(_0887_));
 sg13g2_nor4_2 _3927_ (.A(_0836_),
    .B(_0865_),
    .C(_0887_),
    .Y(_0890_),
    .D(_0888_));
 sg13g2_o21ai_1 _3928_ (.B1(_0889_),
    .Y(_0891_),
    .A1(_0836_),
    .A2(_0865_));
 sg13g2_nand2b_2 _3929_ (.Y(_0892_),
    .B(_0891_),
    .A_N(_0890_));
 sg13g2_o21ai_1 _3930_ (.B1(_0867_),
    .Y(_0064_),
    .A1(net615),
    .A2(_0892_));
 sg13g2_nand2_1 _3931_ (.Y(_0893_),
    .A(net517),
    .B(net613));
 sg13g2_o21ai_1 _3932_ (.B1(_0877_),
    .Y(_0894_),
    .A1(_0843_),
    .A2(_0875_));
 sg13g2_nor3_2 _3933_ (.A(_0035_),
    .B(_0036_),
    .C(_0517_),
    .Y(_0895_));
 sg13g2_o21ai_1 _3934_ (.B1(_0035_),
    .Y(_0896_),
    .A1(_0036_),
    .A2(_0517_));
 sg13g2_nor2b_1 _3935_ (.A(_0895_),
    .B_N(_0896_),
    .Y(_0897_));
 sg13g2_nor2_1 _3936_ (.A(_0037_),
    .B(_0815_),
    .Y(_0898_));
 sg13g2_a21oi_1 _3937_ (.A1(_2454_),
    .A2(_0037_),
    .Y(_0899_),
    .B1(_2453_));
 sg13g2_nor2b_1 _3938_ (.A(_0898_),
    .B_N(_0899_),
    .Y(_0900_));
 sg13g2_a21oi_1 _3939_ (.A1(_2453_),
    .A2(_0037_),
    .Y(_0901_),
    .B1(_0900_));
 sg13g2_nor2b_1 _3940_ (.A(_0874_),
    .B_N(_0901_),
    .Y(_0902_));
 sg13g2_xnor2_1 _3941_ (.Y(_0903_),
    .A(_0874_),
    .B(_0901_));
 sg13g2_xor2_1 _3942_ (.B(_0903_),
    .A(_0897_),
    .X(_0904_));
 sg13g2_and2_1 _3943_ (.A(_0894_),
    .B(_0904_),
    .X(_0905_));
 sg13g2_xor2_1 _3944_ (.B(_0904_),
    .A(_0894_),
    .X(_0906_));
 sg13g2_xnor2_1 _3945_ (.Y(_0907_),
    .A(_0869_),
    .B(_0906_));
 sg13g2_a21oi_1 _3946_ (.A1(_0879_),
    .A2(_0881_),
    .Y(_0908_),
    .B1(_0907_));
 sg13g2_nand3_1 _3947_ (.B(_0881_),
    .C(_0907_),
    .A(_0879_),
    .Y(_0909_));
 sg13g2_nand2b_1 _3948_ (.Y(_0910_),
    .B(_0909_),
    .A_N(_0908_));
 sg13g2_inv_1 _3949_ (.Y(_0911_),
    .A(_0910_));
 sg13g2_nand2_1 _3950_ (.Y(_0912_),
    .A(_0854_),
    .B(_0884_));
 sg13g2_and3_1 _3951_ (.X(_0913_),
    .A(_0861_),
    .B(_0883_),
    .C(_0912_));
 sg13g2_nand2_1 _3952_ (.Y(_0914_),
    .A(_0856_),
    .B(_0884_));
 sg13g2_a22oi_1 _3953_ (.Y(_0915_),
    .B1(_0914_),
    .B2(_0883_),
    .A2(_0913_),
    .A1(_0860_));
 sg13g2_xnor2_1 _3954_ (.Y(_0916_),
    .A(_0910_),
    .B(_0915_));
 sg13g2_xnor2_1 _3955_ (.Y(_0917_),
    .A(_0890_),
    .B(_0916_));
 sg13g2_o21ai_1 _3956_ (.B1(_0893_),
    .Y(_0065_),
    .A1(net615),
    .A2(_0917_));
 sg13g2_nand2_1 _3957_ (.Y(_0918_),
    .A(net469),
    .B(net613));
 sg13g2_a21oi_1 _3958_ (.A1(_0911_),
    .A2(_0915_),
    .Y(_0919_),
    .B1(_0908_));
 sg13g2_a21oi_2 _3959_ (.B1(_0905_),
    .Y(_0920_),
    .A2(_0906_),
    .A1(_0869_));
 sg13g2_a21oi_1 _3960_ (.A1(_0897_),
    .A2(_0903_),
    .Y(_0921_),
    .B1(_0902_));
 sg13g2_nor3_1 _3961_ (.A(_0036_),
    .B(_0037_),
    .C(_0815_),
    .Y(_0922_));
 sg13g2_xor2_1 _3962_ (.B(_0898_),
    .A(_0036_),
    .X(_0923_));
 sg13g2_xnor2_1 _3963_ (.Y(_0924_),
    .A(_0038_),
    .B(_0900_));
 sg13g2_nor2b_1 _3964_ (.A(_0923_),
    .B_N(_0924_),
    .Y(_0925_));
 sg13g2_xor2_1 _3965_ (.B(_0924_),
    .A(_0923_),
    .X(_0926_));
 sg13g2_nor2_1 _3966_ (.A(_0921_),
    .B(_0926_),
    .Y(_0927_));
 sg13g2_xor2_1 _3967_ (.B(_0926_),
    .A(_0921_),
    .X(_0928_));
 sg13g2_xnor2_1 _3968_ (.Y(_0929_),
    .A(_0895_),
    .B(_0928_));
 sg13g2_nor2_1 _3969_ (.A(_0920_),
    .B(_0929_),
    .Y(_0930_));
 sg13g2_xor2_1 _3970_ (.B(_0929_),
    .A(_0920_),
    .X(_0931_));
 sg13g2_xnor2_1 _3971_ (.Y(_0932_),
    .A(_0919_),
    .B(_0931_));
 sg13g2_nand3_1 _3972_ (.B(_0916_),
    .C(_0932_),
    .A(_0890_),
    .Y(_0933_));
 sg13g2_a21o_1 _3973_ (.A2(_0916_),
    .A1(_0890_),
    .B1(_0932_),
    .X(_0934_));
 sg13g2_nand2_2 _3974_ (.Y(_0935_),
    .A(_0933_),
    .B(_0934_));
 sg13g2_o21ai_1 _3975_ (.B1(_0918_),
    .Y(_0066_),
    .A1(net615),
    .A2(_0935_));
 sg13g2_nand2_1 _3976_ (.Y(_0936_),
    .A(net527),
    .B(net613));
 sg13g2_xor2_1 _3977_ (.B(net629),
    .A(net626),
    .X(_0937_));
 sg13g2_a21o_1 _3978_ (.A2(_0900_),
    .A1(net627),
    .B1(_0925_),
    .X(_0938_));
 sg13g2_nand2_1 _3979_ (.Y(_0939_),
    .A(_0937_),
    .B(_0938_));
 sg13g2_xor2_1 _3980_ (.B(_0938_),
    .A(_0937_),
    .X(_0940_));
 sg13g2_nand2_1 _3981_ (.Y(_0941_),
    .A(_0922_),
    .B(_0940_));
 sg13g2_xnor2_1 _3982_ (.Y(_0942_),
    .A(_0922_),
    .B(_0940_));
 sg13g2_a21oi_1 _3983_ (.A1(_0895_),
    .A2(_0928_),
    .Y(_0943_),
    .B1(_0927_));
 sg13g2_or2_1 _3984_ (.X(_0944_),
    .B(_0943_),
    .A(_0942_));
 sg13g2_xnor2_1 _3985_ (.Y(_0945_),
    .A(_0942_),
    .B(_0943_));
 sg13g2_nand2_1 _3986_ (.Y(_0946_),
    .A(_0911_),
    .B(_0931_));
 sg13g2_a221oi_1 _3987_ (.B2(_0883_),
    .C1(_0946_),
    .B1(_0914_),
    .A1(_0860_),
    .Y(_0947_),
    .A2(_0913_));
 sg13g2_nor2_1 _3988_ (.A(_0908_),
    .B(_0930_),
    .Y(_0948_));
 sg13g2_a21oi_1 _3989_ (.A1(_0920_),
    .A2(_0929_),
    .Y(_0949_),
    .B1(_0948_));
 sg13g2_nor2_1 _3990_ (.A(_0947_),
    .B(_0949_),
    .Y(_0950_));
 sg13g2_xor2_1 _3991_ (.B(_0950_),
    .A(_0945_),
    .X(_0951_));
 sg13g2_nand4_1 _3992_ (.B(_0916_),
    .C(_0932_),
    .A(_0890_),
    .Y(_0952_),
    .D(_0951_));
 sg13g2_xor2_1 _3993_ (.B(_0951_),
    .A(_0933_),
    .X(_0953_));
 sg13g2_o21ai_1 _3994_ (.B1(_0936_),
    .Y(_0067_),
    .A1(net615),
    .A2(_0953_));
 sg13g2_nand2_1 _3995_ (.Y(_0954_),
    .A(net744),
    .B(net613));
 sg13g2_nand3_1 _3996_ (.B(net628),
    .C(_0531_),
    .A(net626),
    .Y(_0955_));
 sg13g2_a21o_1 _3997_ (.A2(net628),
    .A1(net625),
    .B1(_0531_),
    .X(_0956_));
 sg13g2_nand2_1 _3998_ (.Y(_0957_),
    .A(_0955_),
    .B(_0956_));
 sg13g2_a21oi_1 _3999_ (.A1(_0939_),
    .A2(_0941_),
    .Y(_0958_),
    .B1(_0957_));
 sg13g2_nand3_1 _4000_ (.B(_0941_),
    .C(_0957_),
    .A(_0939_),
    .Y(_0959_));
 sg13g2_nand2b_1 _4001_ (.Y(_0960_),
    .B(_0959_),
    .A_N(_0958_));
 sg13g2_o21ai_1 _4002_ (.B1(_0944_),
    .Y(_0961_),
    .A1(_0945_),
    .A2(_0950_));
 sg13g2_xor2_1 _4003_ (.B(_0961_),
    .A(_0960_),
    .X(_0962_));
 sg13g2_nor2_1 _4004_ (.A(_0952_),
    .B(_0962_),
    .Y(_0963_));
 sg13g2_xnor2_1 _4005_ (.Y(_0964_),
    .A(_0952_),
    .B(_0962_));
 sg13g2_o21ai_1 _4006_ (.B1(_0954_),
    .Y(_0068_),
    .A1(_0502_),
    .A2(_0964_));
 sg13g2_nand2_1 _4007_ (.Y(_0965_),
    .A(net788),
    .B(net613));
 sg13g2_nand2_1 _4008_ (.Y(_0966_),
    .A(_0530_),
    .B(_0955_));
 sg13g2_nor2_1 _4009_ (.A(_0039_),
    .B(_0530_),
    .Y(_0967_));
 sg13g2_nor2_1 _4010_ (.A(_0039_),
    .B(_0955_),
    .Y(_0968_));
 sg13g2_xor2_1 _4011_ (.B(_0966_),
    .A(_0039_),
    .X(_0969_));
 sg13g2_nor2_1 _4012_ (.A(_0945_),
    .B(_0960_),
    .Y(_0970_));
 sg13g2_o21ai_1 _4013_ (.B1(_0970_),
    .Y(_0971_),
    .A1(_0947_),
    .A2(_0949_));
 sg13g2_nor2_1 _4014_ (.A(_0944_),
    .B(_0960_),
    .Y(_0972_));
 sg13g2_nor2_1 _4015_ (.A(_0958_),
    .B(_0972_),
    .Y(_0973_));
 sg13g2_a21oi_1 _4016_ (.A1(_0971_),
    .A2(_0973_),
    .Y(_0974_),
    .B1(_0969_));
 sg13g2_nand3_1 _4017_ (.B(_0971_),
    .C(_0973_),
    .A(_0969_),
    .Y(_0975_));
 sg13g2_nand2b_1 _4018_ (.Y(_0976_),
    .B(_0975_),
    .A_N(_0974_));
 sg13g2_nor3_1 _4019_ (.A(_0952_),
    .B(_0962_),
    .C(_0976_),
    .Y(_0977_));
 sg13g2_xor2_1 _4020_ (.B(_0976_),
    .A(_0963_),
    .X(_0978_));
 sg13g2_o21ai_1 _4021_ (.B1(_0965_),
    .Y(_0069_),
    .A1(net615),
    .A2(_0978_));
 sg13g2_nand2_1 _4022_ (.Y(_0979_),
    .A(net830),
    .B(net614));
 sg13g2_nor2_1 _4023_ (.A(_0968_),
    .B(_0974_),
    .Y(_0980_));
 sg13g2_xnor2_1 _4024_ (.Y(_0981_),
    .A(_2515_),
    .B(_0967_));
 sg13g2_nor2_1 _4025_ (.A(_0980_),
    .B(_0981_),
    .Y(_0982_));
 sg13g2_xor2_1 _4026_ (.B(_0981_),
    .A(_0980_),
    .X(_0983_));
 sg13g2_xnor2_1 _4027_ (.Y(_0984_),
    .A(_0977_),
    .B(_0983_));
 sg13g2_o21ai_1 _4028_ (.B1(_0979_),
    .Y(_0070_),
    .A1(net615),
    .A2(_0984_));
 sg13g2_nand2_1 _4029_ (.Y(_0985_),
    .A(net798),
    .B(net614));
 sg13g2_a221oi_1 _4030_ (.B2(_0983_),
    .C1(_0982_),
    .B1(_0977_),
    .A1(_2515_),
    .Y(_0986_),
    .A2(_0967_));
 sg13g2_o21ai_1 _4031_ (.B1(_0985_),
    .Y(_0071_),
    .A1(net615),
    .A2(_0986_));
 sg13g2_and2_1 _4032_ (.A(net462),
    .B(net614),
    .X(_0072_));
 sg13g2_nor2_2 _4033_ (.A(\project_audio.f_counter[0] ),
    .B(_0499_),
    .Y(_0987_));
 sg13g2_nand3_1 _4034_ (.B(net624),
    .C(_0987_),
    .A(\project_audio.f_counter[2] ),
    .Y(_0988_));
 sg13g2_and2_1 _4035_ (.A(net712),
    .B(net612),
    .X(_0989_));
 sg13g2_nand2_1 _4036_ (.Y(_0990_),
    .A(net749),
    .B(net592));
 sg13g2_o21ai_1 _4037_ (.B1(_0990_),
    .Y(_0073_),
    .A1(_0808_),
    .A2(net611));
 sg13g2_nand2_1 _4038_ (.Y(_0991_),
    .A(net807),
    .B(net592));
 sg13g2_o21ai_1 _4039_ (.B1(_0991_),
    .Y(_0074_),
    .A1(_0837_),
    .A2(net611));
 sg13g2_nand2_1 _4040_ (.Y(_0992_),
    .A(net509),
    .B(net592));
 sg13g2_o21ai_1 _4041_ (.B1(_0992_),
    .Y(_0075_),
    .A1(_0866_),
    .A2(net611));
 sg13g2_nand2_1 _4042_ (.Y(_0993_),
    .A(net792),
    .B(net592));
 sg13g2_o21ai_1 _4043_ (.B1(_0993_),
    .Y(_0076_),
    .A1(_0892_),
    .A2(net611));
 sg13g2_nand2_1 _4044_ (.Y(_0994_),
    .A(net533),
    .B(net592));
 sg13g2_o21ai_1 _4045_ (.B1(_0994_),
    .Y(_0077_),
    .A1(_0917_),
    .A2(net611));
 sg13g2_nand2_1 _4046_ (.Y(_0995_),
    .A(net475),
    .B(net592));
 sg13g2_o21ai_1 _4047_ (.B1(_0995_),
    .Y(_0078_),
    .A1(_0935_),
    .A2(net612));
 sg13g2_nand2_1 _4048_ (.Y(_0996_),
    .A(net772),
    .B(net593));
 sg13g2_o21ai_1 _4049_ (.B1(_0996_),
    .Y(_0079_),
    .A1(_0953_),
    .A2(net612));
 sg13g2_nand2_1 _4050_ (.Y(_0997_),
    .A(net743),
    .B(net592));
 sg13g2_o21ai_1 _4051_ (.B1(_0997_),
    .Y(_0080_),
    .A1(_0964_),
    .A2(net612));
 sg13g2_nand2_1 _4052_ (.Y(_0998_),
    .A(net776),
    .B(net592));
 sg13g2_o21ai_1 _4053_ (.B1(_0998_),
    .Y(_0081_),
    .A1(_0978_),
    .A2(net611));
 sg13g2_nand2_1 _4054_ (.Y(_0999_),
    .A(net812),
    .B(net593));
 sg13g2_o21ai_1 _4055_ (.B1(_0999_),
    .Y(_0082_),
    .A1(_0984_),
    .A2(net611));
 sg13g2_nand2_1 _4056_ (.Y(_1000_),
    .A(net794),
    .B(net593));
 sg13g2_o21ai_1 _4057_ (.B1(_1000_),
    .Y(_0083_),
    .A1(_0986_),
    .A2(net611));
 sg13g2_and2_1 _4058_ (.A(net444),
    .B(net593),
    .X(_0084_));
 sg13g2_nand3_1 _4059_ (.B(net624),
    .C(_0500_),
    .A(\project_audio.f_counter[2] ),
    .Y(_1001_));
 sg13g2_and2_1 _4060_ (.A(net701),
    .B(net609),
    .X(_1002_));
 sg13g2_nand2_1 _4061_ (.Y(_1003_),
    .A(net528),
    .B(net590));
 sg13g2_o21ai_1 _4062_ (.B1(_1003_),
    .Y(_0085_),
    .A1(_0808_),
    .A2(net609));
 sg13g2_nand2_1 _4063_ (.Y(_1004_),
    .A(net777),
    .B(net590));
 sg13g2_o21ai_1 _4064_ (.B1(_1004_),
    .Y(_0086_),
    .A1(_0837_),
    .A2(net609));
 sg13g2_nand2_1 _4065_ (.Y(_1005_),
    .A(net778),
    .B(net590));
 sg13g2_o21ai_1 _4066_ (.B1(_1005_),
    .Y(_0087_),
    .A1(_0866_),
    .A2(net609));
 sg13g2_nand2_1 _4067_ (.Y(_1006_),
    .A(net806),
    .B(net591));
 sg13g2_o21ai_1 _4068_ (.B1(_1006_),
    .Y(_0088_),
    .A1(_0892_),
    .A2(net610));
 sg13g2_nand2_1 _4069_ (.Y(_1007_),
    .A(net499),
    .B(net591));
 sg13g2_o21ai_1 _4070_ (.B1(_1007_),
    .Y(_0089_),
    .A1(_0917_),
    .A2(net610));
 sg13g2_nand2_1 _4071_ (.Y(_1008_),
    .A(net810),
    .B(net591));
 sg13g2_o21ai_1 _4072_ (.B1(_1008_),
    .Y(_0090_),
    .A1(_0935_),
    .A2(net610));
 sg13g2_nand2_1 _4073_ (.Y(_1009_),
    .A(net829),
    .B(net591));
 sg13g2_o21ai_1 _4074_ (.B1(_1009_),
    .Y(_0091_),
    .A1(_0953_),
    .A2(net609));
 sg13g2_nand2_1 _4075_ (.Y(_1010_),
    .A(net727),
    .B(net590));
 sg13g2_o21ai_1 _4076_ (.B1(_1010_),
    .Y(_0092_),
    .A1(_0964_),
    .A2(net610));
 sg13g2_nand2_1 _4077_ (.Y(_1011_),
    .A(net781),
    .B(net590));
 sg13g2_o21ai_1 _4078_ (.B1(_1011_),
    .Y(_0093_),
    .A1(_0978_),
    .A2(net609));
 sg13g2_nand2_1 _4079_ (.Y(_1012_),
    .A(net851),
    .B(net590));
 sg13g2_o21ai_1 _4080_ (.B1(_1012_),
    .Y(_0094_),
    .A1(_0984_),
    .A2(net609));
 sg13g2_nand2_1 _4081_ (.Y(_1013_),
    .A(net717),
    .B(net590));
 sg13g2_o21ai_1 _4082_ (.B1(_1013_),
    .Y(_0095_),
    .A1(_0986_),
    .A2(net609));
 sg13g2_and2_1 _4083_ (.A(net447),
    .B(net590),
    .X(_0096_));
 sg13g2_nor3_1 _4084_ (.A(\hpos[5] ),
    .B(\hpos[7] ),
    .C(\hpos[6] ),
    .Y(_1014_));
 sg13g2_nand2_1 _4085_ (.Y(_1015_),
    .A(\hpos[8] ),
    .B(_1014_));
 sg13g2_nand2_1 _4086_ (.Y(_1016_),
    .A(\hpos[0] ),
    .B(net1208));
 sg13g2_and4_1 _4087_ (.A(\hpos[0] ),
    .B(net813),
    .C(net910),
    .D(\hpos[1] ),
    .X(_1017_));
 sg13g2_and2_1 _4088_ (.A(net920),
    .B(_1017_),
    .X(_1018_));
 sg13g2_o21ai_1 _4089_ (.B1(net929),
    .Y(_1019_),
    .A1(_1015_),
    .A2(_1018_));
 sg13g2_a21oi_2 _4090_ (.B1(_1019_),
    .Y(_1020_),
    .A2(_1015_),
    .A1(_0023_));
 sg13g2_nor2_2 _4091_ (.A(net680),
    .B(_1020_),
    .Y(_1021_));
 sg13g2_nand2b_2 _4092_ (.Y(_1022_),
    .B(net691),
    .A_N(_1020_));
 sg13g2_and2_1 _4093_ (.A(net434),
    .B(_1021_),
    .X(_0097_));
 sg13g2_or2_1 _4094_ (.X(_1023_),
    .B(net1208),
    .A(\hpos[0] ));
 sg13g2_and3_1 _4095_ (.X(_0098_),
    .A(_1016_),
    .B(_1021_),
    .C(net1209));
 sg13g2_xor2_1 _4096_ (.B(_1016_),
    .A(net910),
    .X(_1024_));
 sg13g2_nor2_1 _4097_ (.A(_1022_),
    .B(net911),
    .Y(_0099_));
 sg13g2_nor2_1 _4098_ (.A(_0008_),
    .B(_1016_),
    .Y(_1025_));
 sg13g2_xnor2_1 _4099_ (.Y(_1026_),
    .A(net813),
    .B(_1025_));
 sg13g2_nor2_1 _4100_ (.A(_1022_),
    .B(net814),
    .Y(_0100_));
 sg13g2_nor2_1 _4101_ (.A(net920),
    .B(_1017_),
    .Y(_1027_));
 sg13g2_nor3_1 _4102_ (.A(_1018_),
    .B(_1022_),
    .C(net921),
    .Y(_0101_));
 sg13g2_nor2b_1 _4103_ (.A(net860),
    .B_N(_1017_),
    .Y(_1028_));
 sg13g2_xnor2_1 _4104_ (.Y(_1029_),
    .A(\hpos[5] ),
    .B(_1028_));
 sg13g2_nor2_1 _4105_ (.A(_1022_),
    .B(net861),
    .Y(_0102_));
 sg13g2_and3_1 _4106_ (.X(_1030_),
    .A(\hpos[5] ),
    .B(net1163),
    .C(\hpos[6] ));
 sg13g2_and2_1 _4107_ (.A(\hpos[5] ),
    .B(_1018_),
    .X(_1031_));
 sg13g2_o21ai_1 _4108_ (.B1(_1021_),
    .Y(_1032_),
    .A1(net821),
    .A2(_1031_));
 sg13g2_a21oi_1 _4109_ (.A1(net821),
    .A2(_1031_),
    .Y(_0103_),
    .B1(_1032_));
 sg13g2_nor2b_1 _4110_ (.A(_0012_),
    .B_N(_1031_),
    .Y(_1033_));
 sg13g2_xnor2_1 _4111_ (.Y(_1034_),
    .A(net1051),
    .B(_1033_));
 sg13g2_nor2_1 _4112_ (.A(_1022_),
    .B(net1052),
    .Y(_0104_));
 sg13g2_nand3_1 _4113_ (.B(_1017_),
    .C(_1030_),
    .A(net1051),
    .Y(_1035_));
 sg13g2_xor2_1 _4114_ (.B(_1035_),
    .A(net1067),
    .X(_1036_));
 sg13g2_nor2_1 _4115_ (.A(_1022_),
    .B(_1036_),
    .Y(_0105_));
 sg13g2_nor2_1 _4116_ (.A(_0023_),
    .B(_1035_),
    .Y(_1037_));
 sg13g2_nor2_1 _4117_ (.A(net929),
    .B(_1037_),
    .Y(_1038_));
 sg13g2_nor2_1 _4118_ (.A(_1022_),
    .B(net930),
    .Y(_0106_));
 sg13g2_nor4_1 _4119_ (.A(\sync_gen.vpos[9] ),
    .B(_2508_),
    .C(\sync_gen.vpos[4] ),
    .D(\sync_gen.vpos[2] ),
    .Y(_1039_));
 sg13g2_nand4_1 _4120_ (.B(net1201),
    .C(net1225),
    .A(\sync_gen.vpos[8] ),
    .Y(_1040_),
    .D(_1039_));
 sg13g2_nor4_1 _4121_ (.A(\sync_gen.vpos[3] ),
    .B(\sync_gen.vpos[1] ),
    .C(\sync_gen.vpos[0] ),
    .D(_1040_),
    .Y(_1041_));
 sg13g2_nor3_1 _4122_ (.A(net815),
    .B(net680),
    .C(net929),
    .Y(_1042_));
 sg13g2_nor3_1 _4123_ (.A(_2506_),
    .B(_2507_),
    .C(_0022_),
    .Y(_1043_));
 sg13g2_a21oi_1 _4124_ (.A1(\sync_gen.vpos[8] ),
    .A2(_1043_),
    .Y(_1044_),
    .B1(_1041_));
 sg13g2_nand2_2 _4125_ (.Y(_1045_),
    .A(_1042_),
    .B(_1044_));
 sg13g2_nor2_2 _4126_ (.A(net675),
    .B(net677),
    .Y(_1046_));
 sg13g2_or2_2 _4127_ (.X(_1047_),
    .B(net677),
    .A(net675));
 sg13g2_nor2_2 _4128_ (.A(net677),
    .B(net679),
    .Y(_1048_));
 sg13g2_nor2_2 _4129_ (.A(\frame_no[0] ),
    .B(_1047_),
    .Y(_1049_));
 sg13g2_nand2b_1 _4130_ (.Y(_1050_),
    .B(_1046_),
    .A_N(net679));
 sg13g2_xnor2_1 _4131_ (.Y(_1051_),
    .A(_0013_),
    .B(_0019_));
 sg13g2_xnor2_1 _4132_ (.Y(_1052_),
    .A(\sync_gen.vpos[7] ),
    .B(_1051_));
 sg13g2_nor2_1 _4133_ (.A(\frame_no[4] ),
    .B(net673),
    .Y(_1053_));
 sg13g2_nor2_2 _4134_ (.A(net670),
    .B(\frame_no[4] ),
    .Y(_1054_));
 sg13g2_nand2b_2 _4135_ (.Y(_1055_),
    .B(_1054_),
    .A_N(\frame_no[6] ));
 sg13g2_or2_1 _4136_ (.X(_1056_),
    .B(_1055_),
    .A(net622));
 sg13g2_xnor2_1 _4137_ (.Y(_1057_),
    .A(\sync_gen.vpos[3] ),
    .B(_0009_));
 sg13g2_xor2_1 _4138_ (.B(_1057_),
    .A(_0015_),
    .X(_1058_));
 sg13g2_xnor2_1 _4139_ (.Y(_1059_),
    .A(_0015_),
    .B(_1057_));
 sg13g2_xnor2_1 _4140_ (.Y(_1060_),
    .A(_0012_),
    .B(_0018_));
 sg13g2_xnor2_1 _4141_ (.Y(_1061_),
    .A(_2507_),
    .B(_1060_));
 sg13g2_nand2b_1 _4142_ (.Y(_1062_),
    .B(_1054_),
    .A_N(net672));
 sg13g2_nand2_2 _4143_ (.Y(_1063_),
    .A(_1054_),
    .B(net621));
 sg13g2_nor2_1 _4144_ (.A(net672),
    .B(_1063_),
    .Y(_1064_));
 sg13g2_a21oi_1 _4145_ (.A1(_1056_),
    .A2(_1063_),
    .Y(_1065_),
    .B1(net673));
 sg13g2_xnor2_1 _4146_ (.Y(_1066_),
    .A(_0011_),
    .B(_0016_));
 sg13g2_xnor2_1 _4147_ (.Y(_1067_),
    .A(\sync_gen.vpos[5] ),
    .B(_1066_));
 sg13g2_and2_1 _4148_ (.A(_2518_),
    .B(net619),
    .X(_1068_));
 sg13g2_xor2_1 _4149_ (.B(_0010_),
    .A(\sync_gen.vpos[4] ),
    .X(_1069_));
 sg13g2_xnor2_1 _4150_ (.Y(_1070_),
    .A(\frame_no[4] ),
    .B(_1069_));
 sg13g2_xnor2_1 _4151_ (.Y(_1071_),
    .A(_0023_),
    .B(_0020_));
 sg13g2_xnor2_1 _4152_ (.Y(_1072_),
    .A(\sync_gen.vpos[8] ),
    .B(_1071_));
 sg13g2_or2_2 _4153_ (.X(_1073_),
    .B(_1055_),
    .A(\frame_no[7] ));
 sg13g2_nor2_1 _4154_ (.A(_1072_),
    .B(_1073_),
    .Y(_1074_));
 sg13g2_o21ai_1 _4155_ (.B1(_1070_),
    .Y(_1075_),
    .A1(net618),
    .A2(_1073_));
 sg13g2_nor2_2 _4156_ (.A(net673),
    .B(net676),
    .Y(_1076_));
 sg13g2_nor2_1 _4157_ (.A(net672),
    .B(_1050_),
    .Y(_1077_));
 sg13g2_nand2_1 _4158_ (.Y(_1078_),
    .A(_1048_),
    .B(_1076_));
 sg13g2_o21ai_1 _4159_ (.B1(_1078_),
    .Y(_1079_),
    .A1(net620),
    .A2(_1070_));
 sg13g2_nand2b_1 _4160_ (.Y(_1080_),
    .B(_1062_),
    .A_N(_1061_));
 sg13g2_xnor2_1 _4161_ (.Y(_1081_),
    .A(\sync_gen.vpos[2] ),
    .B(_0008_));
 sg13g2_xnor2_1 _4162_ (.Y(_1082_),
    .A(_0014_),
    .B(_1048_));
 sg13g2_xnor2_1 _4163_ (.Y(_1083_),
    .A(_1081_),
    .B(_1082_));
 sg13g2_nor2_1 _4164_ (.A(_1073_),
    .B(_1078_),
    .Y(_1084_));
 sg13g2_xnor2_1 _4165_ (.Y(_1085_),
    .A(net679),
    .B(\hpos[0] ));
 sg13g2_xnor2_1 _4166_ (.Y(_1086_),
    .A(\sync_gen.vpos[0] ),
    .B(_1085_));
 sg13g2_xnor2_1 _4167_ (.Y(_1087_),
    .A(net677),
    .B(_0007_));
 sg13g2_xnor2_1 _4168_ (.Y(_1088_),
    .A(\sync_gen.vpos[1] ),
    .B(_1087_));
 sg13g2_xnor2_1 _4169_ (.Y(_1089_),
    .A(\frame_no[0] ),
    .B(_1088_));
 sg13g2_inv_1 _4170_ (.Y(_1090_),
    .A(_1089_));
 sg13g2_and2_1 _4171_ (.A(_1086_),
    .B(_1089_),
    .X(_1091_));
 sg13g2_nor2b_2 _4172_ (.A(net622),
    .B_N(net621),
    .Y(_1092_));
 sg13g2_nand2_1 _4173_ (.Y(_1093_),
    .A(_1058_),
    .B(_1092_));
 sg13g2_o21ai_1 _4174_ (.B1(net623),
    .Y(_1094_),
    .A1(net671),
    .A2(_1055_));
 sg13g2_inv_1 _4175_ (.Y(_1095_),
    .A(_1094_));
 sg13g2_o21ai_1 _4176_ (.B1(_1093_),
    .Y(_1096_),
    .A1(_1050_),
    .A2(_1095_));
 sg13g2_xnor2_1 _4177_ (.Y(_1097_),
    .A(_0017_),
    .B(_1069_));
 sg13g2_o21ai_1 _4178_ (.B1(net623),
    .Y(_1098_),
    .A1(\frame_no[7] ),
    .A2(net618));
 sg13g2_nand2b_1 _4179_ (.Y(_1099_),
    .B(_1098_),
    .A_N(_1055_));
 sg13g2_inv_1 _4180_ (.Y(_1100_),
    .A(_1099_));
 sg13g2_nor2_1 _4181_ (.A(_1097_),
    .B(_1100_),
    .Y(_1101_));
 sg13g2_xnor2_1 _4182_ (.Y(_1102_),
    .A(_1053_),
    .B(net620));
 sg13g2_o21ai_1 _4183_ (.B1(_1047_),
    .Y(_1103_),
    .A1(net620),
    .A2(_1093_));
 sg13g2_nor2_1 _4184_ (.A(_1086_),
    .B(_1088_),
    .Y(_1104_));
 sg13g2_xor2_1 _4185_ (.B(_1081_),
    .A(net676),
    .X(_1105_));
 sg13g2_xnor2_1 _4186_ (.Y(_1106_),
    .A(net678),
    .B(_1105_));
 sg13g2_nor2b_1 _4187_ (.A(_1106_),
    .B_N(_1104_),
    .Y(_1107_));
 sg13g2_nand2b_1 _4188_ (.Y(_1108_),
    .B(_1097_),
    .A_N(net618));
 sg13g2_o21ai_1 _4189_ (.B1(_1108_),
    .Y(_1109_),
    .A1(net671),
    .A2(_1047_));
 sg13g2_nand2_2 _4190_ (.Y(_1110_),
    .A(net618),
    .B(_1073_));
 sg13g2_nand4_1 _4191_ (.B(_1094_),
    .C(_1109_),
    .A(_1080_),
    .Y(_1111_),
    .D(_1110_));
 sg13g2_o21ai_1 _4192_ (.B1(_1070_),
    .Y(_1112_),
    .A1(_2518_),
    .A2(net619));
 sg13g2_nand3b_1 _4193_ (.B(_1063_),
    .C(_1099_),
    .Y(_1113_),
    .A_N(_1112_));
 sg13g2_xor2_1 _4194_ (.B(_1105_),
    .A(_1048_),
    .X(_1114_));
 sg13g2_nand2_1 _4195_ (.Y(_1115_),
    .A(_1091_),
    .B(_1114_));
 sg13g2_nor2_1 _4196_ (.A(net619),
    .B(net618),
    .Y(_1116_));
 sg13g2_nand2_1 _4197_ (.Y(_1117_),
    .A(_1061_),
    .B(_1116_));
 sg13g2_nand2_2 _4198_ (.Y(_1118_),
    .A(net674),
    .B(net676));
 sg13g2_o21ai_1 _4199_ (.B1(net675),
    .Y(_1119_),
    .A1(net678),
    .A2(net679));
 sg13g2_and2_1 _4200_ (.A(net672),
    .B(_1070_),
    .X(_1120_));
 sg13g2_nand2_1 _4201_ (.Y(_1121_),
    .A(net671),
    .B(_1070_));
 sg13g2_a21oi_1 _4202_ (.A1(net672),
    .A2(_1117_),
    .Y(_1122_),
    .B1(_1058_));
 sg13g2_a21oi_1 _4203_ (.A1(_1121_),
    .A2(_1122_),
    .Y(_1123_),
    .B1(_1119_));
 sg13g2_nand2_1 _4204_ (.Y(_1124_),
    .A(net669),
    .B(net622));
 sg13g2_nand2_1 _4205_ (.Y(_1125_),
    .A(_1110_),
    .B(_1124_));
 sg13g2_or2_1 _4206_ (.X(_1126_),
    .B(net621),
    .A(_1054_));
 sg13g2_nor2b_1 _4207_ (.A(_1086_),
    .B_N(_1088_),
    .Y(_1127_));
 sg13g2_nand2_1 _4208_ (.Y(_1128_),
    .A(_1105_),
    .B(_1127_));
 sg13g2_xnor2_1 _4209_ (.Y(_1129_),
    .A(net674),
    .B(_1057_));
 sg13g2_xor2_1 _4210_ (.B(_1057_),
    .A(net674),
    .X(_1130_));
 sg13g2_xnor2_1 _4211_ (.Y(_1131_),
    .A(net675),
    .B(_1129_));
 sg13g2_nand2_1 _4212_ (.Y(_1132_),
    .A(_1113_),
    .B(_1118_));
 sg13g2_nor2_1 _4213_ (.A(\frame_no[4] ),
    .B(net619),
    .Y(_1133_));
 sg13g2_nand2_1 _4214_ (.Y(_1134_),
    .A(net622),
    .B(_1055_));
 sg13g2_nor3_2 _4215_ (.A(_1074_),
    .B(_1097_),
    .C(_1133_),
    .Y(_1135_));
 sg13g2_nand3_1 _4216_ (.B(_1134_),
    .C(_1135_),
    .A(_1056_),
    .Y(_1136_));
 sg13g2_nand2_1 _4217_ (.Y(_1137_),
    .A(net675),
    .B(net678));
 sg13g2_nand3_1 _4218_ (.B(net677),
    .C(net679),
    .A(net676),
    .Y(_1138_));
 sg13g2_nand2_2 _4219_ (.Y(_1139_),
    .A(net677),
    .B(net679));
 sg13g2_inv_1 _4220_ (.Y(_1140_),
    .A(_1139_));
 sg13g2_o21ai_1 _4221_ (.B1(_0015_),
    .Y(_1141_),
    .A1(net674),
    .A2(_1138_));
 sg13g2_nand2b_1 _4222_ (.Y(_1142_),
    .B(_1136_),
    .A_N(_1141_));
 sg13g2_nor2_2 _4223_ (.A(net619),
    .B(_1108_),
    .Y(_1143_));
 sg13g2_nand2b_1 _4224_ (.Y(_1144_),
    .B(_1143_),
    .A_N(net622));
 sg13g2_nand2_2 _4225_ (.Y(_1145_),
    .A(_0014_),
    .B(_1139_));
 sg13g2_nand3b_1 _4226_ (.B(_1130_),
    .C(_1145_),
    .Y(_1146_),
    .A_N(_1081_));
 sg13g2_nand2_1 _4227_ (.Y(_1147_),
    .A(\frame_no[4] ),
    .B(net619));
 sg13g2_and2_1 _4228_ (.A(_1110_),
    .B(_1147_),
    .X(_1148_));
 sg13g2_xnor2_1 _4229_ (.Y(_1149_),
    .A(_0014_),
    .B(_1139_));
 sg13g2_nand2_1 _4230_ (.Y(_1150_),
    .A(_1081_),
    .B(_1149_));
 sg13g2_o21ai_1 _4231_ (.B1(_1129_),
    .Y(_1151_),
    .A1(_0014_),
    .A2(_1139_));
 sg13g2_and4_1 _4232_ (.A(_1146_),
    .B(_1148_),
    .C(_1150_),
    .D(_1151_),
    .X(_1152_));
 sg13g2_nor2b_2 _4233_ (.A(net670),
    .B_N(net619),
    .Y(_1153_));
 sg13g2_xor2_1 _4234_ (.B(_1153_),
    .A(net621),
    .X(_1154_));
 sg13g2_nand4_1 _4235_ (.B(_1090_),
    .C(_1152_),
    .A(_1086_),
    .Y(_1155_),
    .D(_1154_));
 sg13g2_a21oi_1 _4236_ (.A1(_1141_),
    .A2(_1144_),
    .Y(_1156_),
    .B1(_1155_));
 sg13g2_nand2b_1 _4237_ (.Y(_1157_),
    .B(_1075_),
    .A_N(net671));
 sg13g2_o21ai_1 _4238_ (.B1(_1080_),
    .Y(_1158_),
    .A1(net671),
    .A2(_1063_));
 sg13g2_nor2b_1 _4239_ (.A(_1105_),
    .B_N(_1127_),
    .Y(_1159_));
 sg13g2_nor2_1 _4240_ (.A(net623),
    .B(net618),
    .Y(_1160_));
 sg13g2_o21ai_1 _4241_ (.B1(net618),
    .Y(_1161_),
    .A1(net672),
    .A2(_1073_));
 sg13g2_nand2_1 _4242_ (.Y(_1162_),
    .A(_1094_),
    .B(_1161_));
 sg13g2_nand2_1 _4243_ (.Y(_1163_),
    .A(_1121_),
    .B(_1130_));
 sg13g2_o21ai_1 _4244_ (.B1(_1102_),
    .Y(_1164_),
    .A1(net671),
    .A2(_1056_));
 sg13g2_nor2_1 _4245_ (.A(_1163_),
    .B(_1164_),
    .Y(_1165_));
 sg13g2_nand3_1 _4246_ (.B(_1159_),
    .C(_1165_),
    .A(_1157_),
    .Y(_1166_));
 sg13g2_nor3_1 _4247_ (.A(_1158_),
    .B(_1162_),
    .C(_1166_),
    .Y(_1167_));
 sg13g2_and2_1 _4248_ (.A(_1063_),
    .B(_1135_),
    .X(_1168_));
 sg13g2_nor2_1 _4249_ (.A(net676),
    .B(_1140_),
    .Y(_1169_));
 sg13g2_o21ai_1 _4250_ (.B1(net673),
    .Y(_1170_),
    .A1(net675),
    .A2(_1140_));
 sg13g2_nor2b_1 _4251_ (.A(_1168_),
    .B_N(_1170_),
    .Y(_1171_));
 sg13g2_nand2_1 _4252_ (.Y(_1172_),
    .A(_1126_),
    .B(_1148_));
 sg13g2_o21ai_1 _4253_ (.B1(net622),
    .Y(_1173_),
    .A1(net669),
    .A2(net621));
 sg13g2_nor3_1 _4254_ (.A(net669),
    .B(net622),
    .C(net621),
    .Y(_1174_));
 sg13g2_xnor2_1 _4255_ (.Y(_1175_),
    .A(_1129_),
    .B(_1145_));
 sg13g2_nor2_1 _4256_ (.A(_1174_),
    .B(_1175_),
    .Y(_1176_));
 sg13g2_nand4_1 _4257_ (.B(_1148_),
    .C(_1173_),
    .A(_1126_),
    .Y(_1177_),
    .D(_1176_));
 sg13g2_xnor2_1 _4258_ (.Y(_1178_),
    .A(_1105_),
    .B(_1139_));
 sg13g2_nand3_1 _4259_ (.B(_1090_),
    .C(_1178_),
    .A(_1086_),
    .Y(_1179_));
 sg13g2_a21oi_1 _4260_ (.A1(net621),
    .A2(_1143_),
    .Y(_1180_),
    .B1(_1170_));
 sg13g2_nor4_1 _4261_ (.A(_1171_),
    .B(_1177_),
    .C(_1179_),
    .D(_1180_),
    .Y(_1181_));
 sg13g2_nand2_1 _4262_ (.Y(_1182_),
    .A(net671),
    .B(_1047_));
 sg13g2_o21ai_1 _4263_ (.B1(_0017_),
    .Y(_1183_),
    .A1(\frame_no[4] ),
    .A2(_1182_));
 sg13g2_nor3_1 _4264_ (.A(net669),
    .B(net670),
    .C(_1183_),
    .Y(_1184_));
 sg13g2_xnor2_1 _4265_ (.Y(_1185_),
    .A(net620),
    .B(_1183_));
 sg13g2_nand2_1 _4266_ (.Y(_1186_),
    .A(_1046_),
    .B(_1130_));
 sg13g2_nor2b_1 _4267_ (.A(_1070_),
    .B_N(_1182_),
    .Y(_1187_));
 sg13g2_o21ai_1 _4268_ (.B1(_1186_),
    .Y(_1188_),
    .A1(_1160_),
    .A2(_1184_));
 sg13g2_a22oi_1 _4269_ (.Y(_1189_),
    .B1(_1184_),
    .B2(_1098_),
    .A2(_1163_),
    .A1(_1047_));
 sg13g2_nand2_1 _4270_ (.Y(_1190_),
    .A(_1107_),
    .B(_1189_));
 sg13g2_nor4_1 _4271_ (.A(_1185_),
    .B(_1187_),
    .C(_1188_),
    .D(_1190_),
    .Y(_1191_));
 sg13g2_nand3_1 _4272_ (.B(net675),
    .C(net678),
    .A(net673),
    .Y(_1192_));
 sg13g2_o21ai_1 _4273_ (.B1(_0017_),
    .Y(_1193_),
    .A1(\frame_no[4] ),
    .A2(_1192_));
 sg13g2_nor3_1 _4274_ (.A(net669),
    .B(net670),
    .C(_1193_),
    .Y(_1194_));
 sg13g2_xor2_1 _4275_ (.B(_1193_),
    .A(net620),
    .X(_1195_));
 sg13g2_nor2_1 _4276_ (.A(_0015_),
    .B(_1137_),
    .Y(_1196_));
 sg13g2_xnor2_1 _4277_ (.Y(_1197_),
    .A(_1070_),
    .B(_1196_));
 sg13g2_xnor2_1 _4278_ (.Y(_1198_),
    .A(_1059_),
    .B(_1137_));
 sg13g2_o21ai_1 _4279_ (.B1(_1195_),
    .Y(_1199_),
    .A1(_1160_),
    .A2(_1194_));
 sg13g2_nor3_1 _4280_ (.A(_1197_),
    .B(_1198_),
    .C(_1199_),
    .Y(_1200_));
 sg13g2_nand2_1 _4281_ (.Y(_1201_),
    .A(_1104_),
    .B(_1106_));
 sg13g2_a21oi_1 _4282_ (.A1(_1098_),
    .A2(_1194_),
    .Y(_1202_),
    .B1(_1201_));
 sg13g2_a21oi_1 _4283_ (.A1(_1200_),
    .A2(_1202_),
    .Y(_1203_),
    .B1(_1191_));
 sg13g2_a21oi_1 _4284_ (.A1(\frame_no[7] ),
    .A2(net618),
    .Y(_1204_),
    .B1(_1203_));
 sg13g2_nand2_1 _4285_ (.Y(_1205_),
    .A(_1154_),
    .B(_1204_));
 sg13g2_nand2_1 _4286_ (.Y(_1206_),
    .A(net672),
    .B(_1050_));
 sg13g2_nand2b_1 _4287_ (.Y(_1207_),
    .B(_1063_),
    .A_N(_1136_));
 sg13g2_nand2_2 _4288_ (.Y(_1208_),
    .A(_1092_),
    .B(_1143_));
 sg13g2_nand2b_1 _4289_ (.Y(_1209_),
    .B(_1208_),
    .A_N(_1206_));
 sg13g2_xnor2_1 _4290_ (.Y(_1210_),
    .A(_1049_),
    .B(_1129_));
 sg13g2_and4_1 _4291_ (.A(_1083_),
    .B(_1126_),
    .C(_1148_),
    .D(_1210_),
    .X(_1211_));
 sg13g2_nand3_1 _4292_ (.B(_1209_),
    .C(_1211_),
    .A(_1091_),
    .Y(_1212_));
 sg13g2_a21oi_1 _4293_ (.A1(_1206_),
    .A2(_1207_),
    .Y(_1213_),
    .B1(_1212_));
 sg13g2_nand4_1 _4294_ (.B(_1080_),
    .C(_1091_),
    .A(_1079_),
    .Y(_1214_),
    .D(_1096_));
 sg13g2_o21ai_1 _4295_ (.B1(_1049_),
    .Y(_1215_),
    .A1(_1058_),
    .A2(_1065_));
 sg13g2_o21ai_1 _4296_ (.B1(_1077_),
    .Y(_1216_),
    .A1(_1068_),
    .A2(_1112_));
 sg13g2_xnor2_1 _4297_ (.Y(_1217_),
    .A(_1072_),
    .B(_1084_));
 sg13g2_nand4_1 _4298_ (.B(_1215_),
    .C(_1216_),
    .A(_1083_),
    .Y(_1218_),
    .D(_1217_));
 sg13g2_nor2_1 _4299_ (.A(_1046_),
    .B(net619),
    .Y(_1219_));
 sg13g2_o21ai_1 _4300_ (.B1(_1046_),
    .Y(_1220_),
    .A1(_1058_),
    .A2(_1064_));
 sg13g2_o21ai_1 _4301_ (.B1(_1107_),
    .Y(_1221_),
    .A1(_1102_),
    .A2(_1219_));
 sg13g2_nor3_1 _4302_ (.A(net671),
    .B(_1047_),
    .C(_1101_),
    .Y(_1222_));
 sg13g2_nor3_1 _4303_ (.A(_1111_),
    .B(_1221_),
    .C(_1222_),
    .Y(_1223_));
 sg13g2_nand3_1 _4304_ (.B(_1220_),
    .C(_1223_),
    .A(_1103_),
    .Y(_1224_));
 sg13g2_o21ai_1 _4305_ (.B1(_1224_),
    .Y(_1225_),
    .A1(_1214_),
    .A2(_1218_));
 sg13g2_nor2_1 _4306_ (.A(_1213_),
    .B(_1225_),
    .Y(_1226_));
 sg13g2_a21oi_1 _4307_ (.A1(_1142_),
    .A2(_1156_),
    .Y(_1227_),
    .B1(_1181_));
 sg13g2_o21ai_1 _4308_ (.B1(_1113_),
    .Y(_1228_),
    .A1(_1048_),
    .A2(_1118_));
 sg13g2_a22oi_1 _4309_ (.Y(_1229_),
    .B1(_1119_),
    .B2(_1059_),
    .A2(net621),
    .A1(net622));
 sg13g2_nand3b_1 _4310_ (.B(_1126_),
    .C(_1229_),
    .Y(_1230_),
    .A_N(_1068_));
 sg13g2_nor4_1 _4311_ (.A(_1115_),
    .B(_1123_),
    .C(_1125_),
    .D(_1230_),
    .Y(_1231_));
 sg13g2_a21oi_1 _4312_ (.A1(_1054_),
    .A2(_1118_),
    .Y(_1232_),
    .B1(_1092_));
 sg13g2_a21oi_1 _4313_ (.A1(_1120_),
    .A2(_1130_),
    .Y(_1233_),
    .B1(_1232_));
 sg13g2_o21ai_1 _4314_ (.B1(_1233_),
    .Y(_1234_),
    .A1(_1116_),
    .A2(_1118_));
 sg13g2_nor4_1 _4315_ (.A(_1068_),
    .B(_1125_),
    .C(_1128_),
    .D(_1131_),
    .Y(_1235_));
 sg13g2_nor2b_1 _4316_ (.A(_1234_),
    .B_N(_1235_),
    .Y(_1236_));
 sg13g2_a221oi_1 _4317_ (.B2(_1132_),
    .C1(_1167_),
    .B1(_1236_),
    .A1(_1228_),
    .Y(_1237_),
    .A2(_1231_));
 sg13g2_nand4_1 _4318_ (.B(_1226_),
    .C(_1227_),
    .A(_1205_),
    .Y(_1238_),
    .D(_1237_));
 sg13g2_inv_1 _4319_ (.Y(_1239_),
    .A(_1238_));
 sg13g2_xnor2_1 _4320_ (.Y(_1240_),
    .A(net669),
    .B(_0012_));
 sg13g2_xnor2_1 _4321_ (.Y(_1241_),
    .A(_2507_),
    .B(_1240_));
 sg13g2_xor2_1 _4322_ (.B(net670),
    .A(\sync_gen.vpos[5] ),
    .X(_1242_));
 sg13g2_xnor2_1 _4323_ (.Y(_1243_),
    .A(_0011_),
    .B(_1242_));
 sg13g2_xor2_1 _4324_ (.B(\frame_no[7] ),
    .A(\sync_gen.vpos[7] ),
    .X(_1244_));
 sg13g2_xnor2_1 _4325_ (.Y(_1245_),
    .A(_0013_),
    .B(_1244_));
 sg13g2_xnor2_1 _4326_ (.Y(_1246_),
    .A(\sync_gen.vpos[8] ),
    .B(\frame_no[8] ));
 sg13g2_xnor2_1 _4327_ (.Y(_1247_),
    .A(_0023_),
    .B(_1246_));
 sg13g2_nor4_1 _4328_ (.A(_1070_),
    .B(_1241_),
    .C(_1243_),
    .D(_1245_),
    .Y(_1248_));
 sg13g2_nand4_1 _4329_ (.B(_1159_),
    .C(_1247_),
    .A(_1129_),
    .Y(_1249_),
    .D(_1248_));
 sg13g2_inv_1 _4330_ (.Y(_1250_),
    .A(_1249_));
 sg13g2_a21oi_2 _4331_ (.B1(_1045_),
    .Y(_0109_),
    .A2(_1249_),
    .A1(_1239_));
 sg13g2_inv_1 _4332_ (.Y(_1251_),
    .A(_0109_));
 sg13g2_o21ai_1 _4333_ (.B1(_0015_),
    .Y(_1252_),
    .A1(net673),
    .A2(_1119_));
 sg13g2_xnor2_1 _4334_ (.Y(_1253_),
    .A(_1119_),
    .B(_1129_));
 sg13g2_mux2_1 _4335_ (.A0(_1207_),
    .A1(_1208_),
    .S(_1252_),
    .X(_1254_));
 sg13g2_nor4_1 _4336_ (.A(_1115_),
    .B(_1172_),
    .C(_1253_),
    .D(_1254_),
    .Y(_1255_));
 sg13g2_a21oi_1 _4337_ (.A1(_1076_),
    .A2(_1139_),
    .Y(_1256_),
    .B1(_1143_));
 sg13g2_nor2_1 _4338_ (.A(_1092_),
    .B(_1153_),
    .Y(_1257_));
 sg13g2_xnor2_1 _4339_ (.Y(_1258_),
    .A(_1058_),
    .B(_1145_));
 sg13g2_nand4_1 _4340_ (.B(_1124_),
    .C(_1147_),
    .A(_1110_),
    .Y(_1259_),
    .D(_1258_));
 sg13g2_nor3_1 _4341_ (.A(_1256_),
    .B(_1257_),
    .C(_1259_),
    .Y(_1260_));
 sg13g2_nand2_1 _4342_ (.Y(_1261_),
    .A(_1056_),
    .B(_1168_));
 sg13g2_nand2_1 _4343_ (.Y(_1262_),
    .A(_1076_),
    .B(_1261_));
 sg13g2_a21oi_1 _4344_ (.A1(_1092_),
    .A2(_1143_),
    .Y(_1263_),
    .B1(_1076_));
 sg13g2_nand2_1 _4345_ (.Y(_1264_),
    .A(_1131_),
    .B(_1134_));
 sg13g2_nor4_1 _4346_ (.A(_1128_),
    .B(_1172_),
    .C(_1263_),
    .D(_1264_),
    .Y(_1265_));
 sg13g2_nor2_1 _4347_ (.A(_1162_),
    .B(_1201_),
    .Y(_1266_));
 sg13g2_nand2_1 _4348_ (.Y(_1267_),
    .A(_1057_),
    .B(_1100_));
 sg13g2_nor2_1 _4349_ (.A(_1135_),
    .B(_1140_),
    .Y(_1268_));
 sg13g2_nand2_1 _4350_ (.Y(_1269_),
    .A(_1102_),
    .B(_1130_));
 sg13g2_xnor2_1 _4351_ (.Y(_1270_),
    .A(_0015_),
    .B(_1097_));
 sg13g2_nor3_1 _4352_ (.A(_1158_),
    .B(_1269_),
    .C(_1270_),
    .Y(_1271_));
 sg13g2_a22oi_1 _4353_ (.Y(_1272_),
    .B1(_1267_),
    .B2(_1271_),
    .A2(net677),
    .A1(net675));
 sg13g2_nor2_1 _4354_ (.A(_1130_),
    .B(_1208_),
    .Y(_1273_));
 sg13g2_a221oi_1 _4355_ (.B2(_1076_),
    .C1(_1179_),
    .B1(_1268_),
    .A1(_1065_),
    .Y(_1274_),
    .A2(_1169_));
 sg13g2_a221oi_1 _4356_ (.B2(_1260_),
    .C1(_1255_),
    .B1(_1274_),
    .A1(_1262_),
    .Y(_1275_),
    .A2(_1265_));
 sg13g2_o21ai_1 _4357_ (.B1(_1266_),
    .Y(_1276_),
    .A1(_1137_),
    .A2(_1273_));
 sg13g2_o21ai_1 _4358_ (.B1(_1275_),
    .Y(_1277_),
    .A1(_1272_),
    .A2(_1276_));
 sg13g2_o21ai_1 _4359_ (.B1(net692),
    .Y(_1278_),
    .A1(_1238_),
    .A2(_1277_));
 sg13g2_and2_1 _4360_ (.A(_0109_),
    .B(_1278_),
    .X(_0107_));
 sg13g2_nor3_1 _4361_ (.A(_1225_),
    .B(_1250_),
    .C(_1277_),
    .Y(_1279_));
 sg13g2_nor2_1 _4362_ (.A(_1045_),
    .B(_1279_),
    .Y(_0110_));
 sg13g2_nor2b_2 _4363_ (.A(net1236),
    .B_N(net793),
    .Y(_1280_));
 sg13g2_o21ai_1 _4364_ (.B1(net691),
    .Y(_1281_),
    .A1(net679),
    .A2(_1280_));
 sg13g2_a21oi_1 _4365_ (.A1(_2510_),
    .A2(_1280_),
    .Y(_0111_),
    .B1(_1281_));
 sg13g2_a21oi_1 _4366_ (.A1(net679),
    .A2(_1280_),
    .Y(_1282_),
    .B1(net677));
 sg13g2_nand2_2 _4367_ (.Y(_1283_),
    .A(_1140_),
    .B(_1280_));
 sg13g2_nand2_1 _4368_ (.Y(_1284_),
    .A(net691),
    .B(_1283_));
 sg13g2_nor2_1 _4369_ (.A(net1222),
    .B(_1284_),
    .Y(_0112_));
 sg13g2_o21ai_1 _4370_ (.B1(net691),
    .Y(_1285_),
    .A1(net676),
    .A2(_1280_));
 sg13g2_a21oi_1 _4371_ (.A1(_1149_),
    .A2(_1280_),
    .Y(_0113_),
    .B1(_1285_));
 sg13g2_nor2_1 _4372_ (.A(_0014_),
    .B(_1283_),
    .Y(_1286_));
 sg13g2_o21ai_1 _4373_ (.B1(net691),
    .Y(_1287_),
    .A1(net674),
    .A2(_1286_));
 sg13g2_a21oi_1 _4374_ (.A1(net674),
    .A2(_1286_),
    .Y(_0114_),
    .B1(_1287_));
 sg13g2_o21ai_1 _4375_ (.B1(_2509_),
    .Y(_1288_),
    .A1(_1118_),
    .A2(_1283_));
 sg13g2_nor3_2 _4376_ (.A(_2509_),
    .B(_1118_),
    .C(_1283_),
    .Y(_1289_));
 sg13g2_nand2_1 _4377_ (.Y(_1290_),
    .A(net691),
    .B(_1288_));
 sg13g2_nor2_1 _4378_ (.A(_1289_),
    .B(_1290_),
    .Y(_0115_));
 sg13g2_nor3_1 _4379_ (.A(_0017_),
    .B(_1118_),
    .C(_1283_),
    .Y(_1291_));
 sg13g2_o21ai_1 _4380_ (.B1(net691),
    .Y(_1292_),
    .A1(net670),
    .A2(_1291_));
 sg13g2_a21oi_1 _4381_ (.A1(net670),
    .A2(_1291_),
    .Y(_0116_),
    .B1(_1292_));
 sg13g2_nand2_1 _4382_ (.Y(_1293_),
    .A(net670),
    .B(_1289_));
 sg13g2_xor2_1 _4383_ (.B(_1293_),
    .A(net669),
    .X(_1294_));
 sg13g2_nor2_1 _4384_ (.A(net680),
    .B(_1294_),
    .Y(_0117_));
 sg13g2_nor2_1 _4385_ (.A(net1122),
    .B(_1293_),
    .Y(_1295_));
 sg13g2_o21ai_1 _4386_ (.B1(net692),
    .Y(_1296_),
    .A1(\frame_no[7] ),
    .A2(_1295_));
 sg13g2_a21oi_1 _4387_ (.A1(\frame_no[7] ),
    .A2(_1295_),
    .Y(_0118_),
    .B1(_1296_));
 sg13g2_and4_1 _4388_ (.A(\frame_no[7] ),
    .B(net669),
    .C(\frame_no[5] ),
    .D(_1289_),
    .X(_1297_));
 sg13g2_o21ai_1 _4389_ (.B1(net692),
    .Y(_1298_),
    .A1(net457),
    .A2(_1297_));
 sg13g2_a21oi_1 _4390_ (.A1(net457),
    .A2(_1297_),
    .Y(_0119_),
    .B1(_1298_));
 sg13g2_nor2_1 _4391_ (.A(_1251_),
    .B(_1278_),
    .Y(_0120_));
 sg13g2_nor2b_1 _4392_ (.A(_1278_),
    .B_N(_0110_),
    .Y(_0121_));
 sg13g2_or3_1 _4393_ (.A(\sync_gen.vpos[6] ),
    .B(\sync_gen.vpos[5] ),
    .C(\sync_gen.vpos[4] ),
    .X(_1299_));
 sg13g2_and2_1 _4394_ (.A(\sync_gen.vpos[3] ),
    .B(\sync_gen.vpos[2] ),
    .X(_1300_));
 sg13g2_nor4_1 _4395_ (.A(\sync_gen.vpos[8] ),
    .B(\sync_gen.vpos[7] ),
    .C(_1299_),
    .D(_1300_),
    .Y(_1301_));
 sg13g2_nand2b_2 _4396_ (.Y(_1302_),
    .B(net815),
    .A_N(_1301_));
 sg13g2_a21oi_1 _4397_ (.A1(_1020_),
    .A2(_1302_),
    .Y(_1303_),
    .B1(net1195));
 sg13g2_and2_1 _4398_ (.A(\sync_gen.vpos[0] ),
    .B(_1020_),
    .X(_1304_));
 sg13g2_nor3_1 _4399_ (.A(net680),
    .B(net1196),
    .C(_1304_),
    .Y(_0122_));
 sg13g2_a21oi_2 _4400_ (.B1(_1021_),
    .Y(_1305_),
    .A2(_1302_),
    .A1(net693));
 sg13g2_xnor2_1 _4401_ (.Y(_1306_),
    .A(net1235),
    .B(_1304_));
 sg13g2_nor2_1 _4402_ (.A(_1305_),
    .B(_1306_),
    .Y(_0123_));
 sg13g2_a21oi_1 _4403_ (.A1(\sync_gen.vpos[1] ),
    .A2(_1304_),
    .Y(_1307_),
    .B1(net1104));
 sg13g2_and3_1 _4404_ (.X(_1308_),
    .A(net1104),
    .B(\sync_gen.vpos[1] ),
    .C(_1304_));
 sg13g2_nor3_1 _4405_ (.A(_1305_),
    .B(net1105),
    .C(_1308_),
    .Y(_0124_));
 sg13g2_xnor2_1 _4406_ (.Y(_1309_),
    .A(net1220),
    .B(_1308_));
 sg13g2_nor2_1 _4407_ (.A(_1305_),
    .B(_1309_),
    .Y(_0125_));
 sg13g2_a21oi_1 _4408_ (.A1(\sync_gen.vpos[3] ),
    .A2(_1308_),
    .Y(_1310_),
    .B1(net917));
 sg13g2_and4_1 _4409_ (.A(\sync_gen.vpos[4] ),
    .B(\sync_gen.vpos[1] ),
    .C(\sync_gen.vpos[0] ),
    .D(_1300_),
    .X(_1311_));
 sg13g2_a21oi_1 _4410_ (.A1(_1022_),
    .A2(_1311_),
    .Y(_1312_),
    .B1(_1305_));
 sg13g2_nor2b_1 _4411_ (.A(net918),
    .B_N(_1312_),
    .Y(_0126_));
 sg13g2_xnor2_1 _4412_ (.Y(_1313_),
    .A(_0022_),
    .B(_1311_));
 sg13g2_and3_1 _4413_ (.X(_1314_),
    .A(_1020_),
    .B(_1302_),
    .C(_1313_));
 sg13g2_a22oi_1 _4414_ (.Y(_1315_),
    .B1(_1314_),
    .B2(net692),
    .A2(_1021_),
    .A1(net1187));
 sg13g2_inv_1 _4415_ (.Y(_0127_),
    .A(net1188));
 sg13g2_nand3_1 _4416_ (.B(_1020_),
    .C(_1311_),
    .A(net1187),
    .Y(_1316_));
 sg13g2_and2_1 _4417_ (.A(_2507_),
    .B(_1316_),
    .X(_1317_));
 sg13g2_nor2_1 _4418_ (.A(_2507_),
    .B(_1316_),
    .Y(_1318_));
 sg13g2_nor3_1 _4419_ (.A(_1305_),
    .B(_1317_),
    .C(_1318_),
    .Y(_0128_));
 sg13g2_a21oi_1 _4420_ (.A1(_1302_),
    .A2(_1318_),
    .Y(_1319_),
    .B1(net1201));
 sg13g2_and2_1 _4421_ (.A(net1201),
    .B(_1318_),
    .X(_1320_));
 sg13g2_nor3_1 _4422_ (.A(_1305_),
    .B(net1202),
    .C(_1320_),
    .Y(_0129_));
 sg13g2_xnor2_1 _4423_ (.Y(_1321_),
    .A(net1228),
    .B(_1320_));
 sg13g2_nor2_1 _4424_ (.A(_1305_),
    .B(_1321_),
    .Y(_0130_));
 sg13g2_a21oi_1 _4425_ (.A1(\sync_gen.vpos[8] ),
    .A2(_1320_),
    .Y(_1322_),
    .B1(net815));
 sg13g2_nor2_1 _4426_ (.A(_1305_),
    .B(net816),
    .Y(_0131_));
 sg13g2_nor3_1 _4427_ (.A(\hpos[5] ),
    .B(net920),
    .C(net821),
    .Y(_1323_));
 sg13g2_nand3_1 _4428_ (.B(net929),
    .C(net1051),
    .A(net691),
    .Y(_1324_));
 sg13g2_or4_1 _4429_ (.A(net1067),
    .B(_1030_),
    .C(_1323_),
    .D(_1324_),
    .X(_0132_));
 sg13g2_nand3_1 _4430_ (.B(\sync_gen.vpos[1] ),
    .C(net692),
    .A(net1220),
    .Y(_1325_));
 sg13g2_o21ai_1 _4431_ (.B1(_1300_),
    .Y(_1326_),
    .A1(\sync_gen.vpos[1] ),
    .A2(\sync_gen.vpos[0] ));
 sg13g2_nor2_1 _4432_ (.A(\sync_gen.vpos[0] ),
    .B(_1043_),
    .Y(_1327_));
 sg13g2_a21oi_1 _4433_ (.A1(_1043_),
    .A2(_1326_),
    .Y(_1328_),
    .B1(_1327_));
 sg13g2_or3_1 _4434_ (.A(net1226),
    .B(_1325_),
    .C(_1328_),
    .X(_0133_));
 sg13g2_and3_1 _4435_ (.X(_1329_),
    .A(\project_audio.nco_increment_gen.counter[0] ),
    .B(net464),
    .C(net497));
 sg13g2_and2_1 _4436_ (.A(net751),
    .B(_1329_),
    .X(_1330_));
 sg13g2_and2_1 _4437_ (.A(net790),
    .B(_1330_),
    .X(_1331_));
 sg13g2_and2_1 _4438_ (.A(net862),
    .B(_1331_),
    .X(_1332_));
 sg13g2_nand3_1 _4439_ (.B(net782),
    .C(_1332_),
    .A(net459),
    .Y(_1333_));
 sg13g2_nand2_1 _4440_ (.Y(_1334_),
    .A(net693),
    .B(_1333_));
 sg13g2_nand2_1 _4441_ (.Y(_1335_),
    .A(net693),
    .B(_0024_));
 sg13g2_o21ai_1 _4442_ (.B1(net693),
    .Y(_1336_),
    .A1(_0024_),
    .A2(_1333_));
 sg13g2_nor2b_1 _4443_ (.A(_1336_),
    .B_N(net435),
    .Y(_0134_));
 sg13g2_xnor2_1 _4444_ (.Y(_1337_),
    .A(net963),
    .B(net497));
 sg13g2_nor2_1 _4445_ (.A(_1336_),
    .B(_1337_),
    .Y(_0135_));
 sg13g2_a21oi_1 _4446_ (.A1(\project_audio.nco_increment_gen.counter[0] ),
    .A2(\project_audio.nco_increment_gen.counter[1] ),
    .Y(_1338_),
    .B1(net464));
 sg13g2_nor3_1 _4447_ (.A(_1329_),
    .B(_1336_),
    .C(net465),
    .Y(_0136_));
 sg13g2_nor2_1 _4448_ (.A(net751),
    .B(_1329_),
    .Y(_1339_));
 sg13g2_nor3_1 _4449_ (.A(_1330_),
    .B(_1336_),
    .C(net752),
    .Y(_0137_));
 sg13g2_nor2_1 _4450_ (.A(net790),
    .B(_1330_),
    .Y(_1340_));
 sg13g2_nor3_1 _4451_ (.A(_1331_),
    .B(_1336_),
    .C(_1340_),
    .Y(_0138_));
 sg13g2_nor2_1 _4452_ (.A(net862),
    .B(_1331_),
    .Y(_1341_));
 sg13g2_nor3_1 _4453_ (.A(net680),
    .B(_1332_),
    .C(_1341_),
    .Y(_0139_));
 sg13g2_o21ai_1 _4454_ (.B1(net693),
    .Y(_1342_),
    .A1(net782),
    .A2(_1332_));
 sg13g2_a21oi_1 _4455_ (.A1(net782),
    .A2(_1332_),
    .Y(_0140_),
    .B1(_1342_));
 sg13g2_a21oi_1 _4456_ (.A1(\project_audio.nco_increment_gen.counter[6] ),
    .A2(_1332_),
    .Y(_1343_),
    .B1(net459));
 sg13g2_nor2_1 _4457_ (.A(_1334_),
    .B(net460),
    .Y(_0141_));
 sg13g2_nand2b_1 _4458_ (.Y(_1344_),
    .B(_2514_),
    .A_N(_1335_));
 sg13g2_a22oi_1 _4459_ (.Y(_0142_),
    .B1(_1334_),
    .B2(_1344_),
    .A2(_1333_),
    .A1(_2514_));
 sg13g2_nand2_2 _4460_ (.Y(_1345_),
    .A(_0501_),
    .B(_0987_));
 sg13g2_a21oi_1 _4461_ (.A1(_0501_),
    .A2(_0987_),
    .Y(_1346_),
    .B1(net684));
 sg13g2_nand2_1 _4462_ (.Y(_1347_),
    .A(net482),
    .B(net607));
 sg13g2_o21ai_1 _4463_ (.B1(_1347_),
    .Y(_0143_),
    .A1(_0808_),
    .A2(net608));
 sg13g2_nand2_1 _4464_ (.Y(_1348_),
    .A(net764),
    .B(net607));
 sg13g2_o21ai_1 _4465_ (.B1(_1348_),
    .Y(_0144_),
    .A1(_0837_),
    .A2(net608));
 sg13g2_nand2_1 _4466_ (.Y(_1349_),
    .A(net518),
    .B(net607));
 sg13g2_o21ai_1 _4467_ (.B1(_1349_),
    .Y(_0145_),
    .A1(_0866_),
    .A2(_1345_));
 sg13g2_nand2_1 _4468_ (.Y(_1350_),
    .A(net796),
    .B(net607));
 sg13g2_o21ai_1 _4469_ (.B1(_1350_),
    .Y(_0146_),
    .A1(_0892_),
    .A2(_1345_));
 sg13g2_nand2_1 _4470_ (.Y(_1351_),
    .A(net520),
    .B(net606));
 sg13g2_o21ai_1 _4471_ (.B1(_1351_),
    .Y(_0147_),
    .A1(_0917_),
    .A2(_1345_));
 sg13g2_nand2_1 _4472_ (.Y(_1352_),
    .A(net467),
    .B(net606));
 sg13g2_o21ai_1 _4473_ (.B1(_1352_),
    .Y(_0148_),
    .A1(_0935_),
    .A2(net608));
 sg13g2_nand2_1 _4474_ (.Y(_1353_),
    .A(net733),
    .B(net606));
 sg13g2_o21ai_1 _4475_ (.B1(_1353_),
    .Y(_0149_),
    .A1(_0953_),
    .A2(net608));
 sg13g2_nand2_1 _4476_ (.Y(_1354_),
    .A(net802),
    .B(net606));
 sg13g2_o21ai_1 _4477_ (.B1(_1354_),
    .Y(_0150_),
    .A1(_0964_),
    .A2(net608));
 sg13g2_nand2_1 _4478_ (.Y(_1355_),
    .A(net496),
    .B(net606));
 sg13g2_o21ai_1 _4479_ (.B1(_1355_),
    .Y(_0151_),
    .A1(_0978_),
    .A2(net608));
 sg13g2_nand2_1 _4480_ (.Y(_1356_),
    .A(net823),
    .B(net606));
 sg13g2_o21ai_1 _4481_ (.B1(_1356_),
    .Y(_0152_),
    .A1(_0984_),
    .A2(net608));
 sg13g2_nand2_1 _4482_ (.Y(_1357_),
    .A(net818),
    .B(net606));
 sg13g2_o21ai_1 _4483_ (.B1(_1357_),
    .Y(_0153_),
    .A1(_0986_),
    .A2(net608));
 sg13g2_and2_1 _4484_ (.A(net448),
    .B(net606),
    .X(_0154_));
 sg13g2_nand2b_1 _4485_ (.Y(_0155_),
    .B(net699),
    .A_N(net793));
 sg13g2_nor2b_2 _4486_ (.A(\project_audio.f_counter[2] ),
    .B_N(net624),
    .Y(_1358_));
 sg13g2_nand2_2 _4487_ (.Y(_1359_),
    .A(_0500_),
    .B(_1358_));
 sg13g2_a21oi_1 _4488_ (.A1(_0500_),
    .A2(_1358_),
    .Y(_1360_),
    .B1(net683));
 sg13g2_nand2_1 _4489_ (.Y(_1361_),
    .A(net470),
    .B(net604));
 sg13g2_o21ai_1 _4490_ (.B1(_1361_),
    .Y(_0156_),
    .A1(_0808_),
    .A2(_1359_));
 sg13g2_nand2_1 _4491_ (.Y(_1362_),
    .A(net501),
    .B(net604));
 sg13g2_o21ai_1 _4492_ (.B1(_1362_),
    .Y(_0157_),
    .A1(_0837_),
    .A2(_1359_));
 sg13g2_nand2_1 _4493_ (.Y(_1363_),
    .A(net725),
    .B(net604));
 sg13g2_o21ai_1 _4494_ (.B1(_1363_),
    .Y(_0158_),
    .A1(_0866_),
    .A2(_1359_));
 sg13g2_nand2_1 _4495_ (.Y(_1364_),
    .A(net831),
    .B(net603));
 sg13g2_o21ai_1 _4496_ (.B1(_1364_),
    .Y(_0159_),
    .A1(_0892_),
    .A2(net605));
 sg13g2_nand2_1 _4497_ (.Y(_1365_),
    .A(net799),
    .B(net604));
 sg13g2_o21ai_1 _4498_ (.B1(_1365_),
    .Y(_0160_),
    .A1(_0917_),
    .A2(net605));
 sg13g2_nand2_1 _4499_ (.Y(_1366_),
    .A(net491),
    .B(net603));
 sg13g2_o21ai_1 _4500_ (.B1(_1366_),
    .Y(_0161_),
    .A1(_0935_),
    .A2(net605));
 sg13g2_nand2_1 _4501_ (.Y(_1367_),
    .A(net844),
    .B(net603));
 sg13g2_o21ai_1 _4502_ (.B1(_1367_),
    .Y(_0162_),
    .A1(_0953_),
    .A2(net605));
 sg13g2_nand2_1 _4503_ (.Y(_1368_),
    .A(net765),
    .B(net603));
 sg13g2_o21ai_1 _4504_ (.B1(_1368_),
    .Y(_0163_),
    .A1(_0964_),
    .A2(net605));
 sg13g2_nand2_1 _4505_ (.Y(_1369_),
    .A(net769),
    .B(net603));
 sg13g2_o21ai_1 _4506_ (.B1(_1369_),
    .Y(_0164_),
    .A1(_0978_),
    .A2(net605));
 sg13g2_nand2_1 _4507_ (.Y(_1370_),
    .A(net843),
    .B(net603));
 sg13g2_o21ai_1 _4508_ (.B1(_1370_),
    .Y(_0165_),
    .A1(_0984_),
    .A2(net605));
 sg13g2_nand2_1 _4509_ (.Y(_1371_),
    .A(net724),
    .B(net603));
 sg13g2_o21ai_1 _4510_ (.B1(_1371_),
    .Y(_0166_),
    .A1(_0986_),
    .A2(net605));
 sg13g2_and2_1 _4511_ (.A(net454),
    .B(net603),
    .X(_0167_));
 sg13g2_nor2_2 _4512_ (.A(\project_audio.f_counter[2] ),
    .B(net624),
    .Y(_1372_));
 sg13g2_nand2_2 _4513_ (.Y(_1373_),
    .A(_0987_),
    .B(_1372_));
 sg13g2_a21oi_1 _4514_ (.A1(_0987_),
    .A2(_1372_),
    .Y(_1374_),
    .B1(net683));
 sg13g2_nand2_1 _4515_ (.Y(_1375_),
    .A(net479),
    .B(net600));
 sg13g2_o21ai_1 _4516_ (.B1(_1375_),
    .Y(_0168_),
    .A1(_0808_),
    .A2(net602));
 sg13g2_nand2_1 _4517_ (.Y(_1376_),
    .A(net728),
    .B(net600));
 sg13g2_o21ai_1 _4518_ (.B1(_1376_),
    .Y(_0169_),
    .A1(_0837_),
    .A2(net602));
 sg13g2_nand2_1 _4519_ (.Y(_1377_),
    .A(net534),
    .B(net600));
 sg13g2_o21ai_1 _4520_ (.B1(_1377_),
    .Y(_0170_),
    .A1(_0866_),
    .A2(net602));
 sg13g2_nand2_1 _4521_ (.Y(_1378_),
    .A(net741),
    .B(net601));
 sg13g2_o21ai_1 _4522_ (.B1(_1378_),
    .Y(_0171_),
    .A1(_0892_),
    .A2(_1373_));
 sg13g2_nand2_1 _4523_ (.Y(_1379_),
    .A(net817),
    .B(net600));
 sg13g2_o21ai_1 _4524_ (.B1(_1379_),
    .Y(_0172_),
    .A1(_0917_),
    .A2(_1373_));
 sg13g2_nand2_1 _4525_ (.Y(_1380_),
    .A(net463),
    .B(net600));
 sg13g2_o21ai_1 _4526_ (.B1(_1380_),
    .Y(_0173_),
    .A1(_0935_),
    .A2(_1373_));
 sg13g2_nand2_1 _4527_ (.Y(_1381_),
    .A(net757),
    .B(net600));
 sg13g2_o21ai_1 _4528_ (.B1(_1381_),
    .Y(_0174_),
    .A1(_0953_),
    .A2(net602));
 sg13g2_nand2_1 _4529_ (.Y(_1382_),
    .A(net529),
    .B(net601));
 sg13g2_o21ai_1 _4530_ (.B1(_1382_),
    .Y(_0175_),
    .A1(_0964_),
    .A2(net602));
 sg13g2_nand2_1 _4531_ (.Y(_1383_),
    .A(net784),
    .B(net601));
 sg13g2_o21ai_1 _4532_ (.B1(_1383_),
    .Y(_0176_),
    .A1(_0978_),
    .A2(net602));
 sg13g2_nand2_1 _4533_ (.Y(_1384_),
    .A(net836),
    .B(net601));
 sg13g2_o21ai_1 _4534_ (.B1(_1384_),
    .Y(_0177_),
    .A1(_0984_),
    .A2(net602));
 sg13g2_nand2_1 _4535_ (.Y(_1385_),
    .A(net832),
    .B(net600));
 sg13g2_o21ai_1 _4536_ (.B1(_1385_),
    .Y(_0178_),
    .A1(_0986_),
    .A2(net602));
 sg13g2_and2_1 _4537_ (.A(net785),
    .B(net600),
    .X(_0179_));
 sg13g2_nand2_2 _4538_ (.Y(_1386_),
    .A(_0987_),
    .B(_1358_));
 sg13g2_a21oi_1 _4539_ (.A1(_0987_),
    .A2(_1358_),
    .Y(_1387_),
    .B1(net683));
 sg13g2_nand2_1 _4540_ (.Y(_1388_),
    .A(net472),
    .B(net597));
 sg13g2_o21ai_1 _4541_ (.B1(_1388_),
    .Y(_0180_),
    .A1(_0808_),
    .A2(net599));
 sg13g2_nand2_1 _4542_ (.Y(_1389_),
    .A(net515),
    .B(net597));
 sg13g2_o21ai_1 _4543_ (.B1(_1389_),
    .Y(_0181_),
    .A1(_0837_),
    .A2(_1386_));
 sg13g2_nand2_1 _4544_ (.Y(_1390_),
    .A(net746),
    .B(net598));
 sg13g2_o21ai_1 _4545_ (.B1(_1390_),
    .Y(_0182_),
    .A1(_0866_),
    .A2(_1386_));
 sg13g2_nand2_1 _4546_ (.Y(_1391_),
    .A(net789),
    .B(net598));
 sg13g2_o21ai_1 _4547_ (.B1(_1391_),
    .Y(_0183_),
    .A1(_0892_),
    .A2(net599));
 sg13g2_nand2_1 _4548_ (.Y(_1392_),
    .A(net742),
    .B(net598));
 sg13g2_o21ai_1 _4549_ (.B1(_1392_),
    .Y(_0184_),
    .A1(_0917_),
    .A2(_1386_));
 sg13g2_nand2_1 _4550_ (.Y(_1393_),
    .A(net532),
    .B(net598));
 sg13g2_o21ai_1 _4551_ (.B1(_1393_),
    .Y(_0185_),
    .A1(_0935_),
    .A2(net599));
 sg13g2_nand2_1 _4552_ (.Y(_1394_),
    .A(net732),
    .B(net597));
 sg13g2_o21ai_1 _4553_ (.B1(_1394_),
    .Y(_0186_),
    .A1(_0953_),
    .A2(net599));
 sg13g2_nand2_1 _4554_ (.Y(_1395_),
    .A(net773),
    .B(net597));
 sg13g2_o21ai_1 _4555_ (.B1(_1395_),
    .Y(_0187_),
    .A1(_0964_),
    .A2(net599));
 sg13g2_nand2_1 _4556_ (.Y(_1396_),
    .A(net734),
    .B(net597));
 sg13g2_o21ai_1 _4557_ (.B1(_1396_),
    .Y(_0188_),
    .A1(_0978_),
    .A2(net599));
 sg13g2_nand2_1 _4558_ (.Y(_1397_),
    .A(net824),
    .B(net597));
 sg13g2_o21ai_1 _4559_ (.B1(_1397_),
    .Y(_0189_),
    .A1(_0984_),
    .A2(net599));
 sg13g2_nand2_1 _4560_ (.Y(_1398_),
    .A(net737),
    .B(net597));
 sg13g2_o21ai_1 _4561_ (.B1(_1398_),
    .Y(_0190_),
    .A1(_0986_),
    .A2(net599));
 sg13g2_and2_1 _4562_ (.A(net445),
    .B(net597),
    .X(_0191_));
 sg13g2_nand3_1 _4563_ (.B(net569),
    .C(net559),
    .A(net959),
    .Y(_1399_));
 sg13g2_o21ai_1 _4564_ (.B1(_1399_),
    .Y(_0192_),
    .A1(_2505_),
    .A2(net569));
 sg13g2_nand3_1 _4565_ (.B(net569),
    .C(net559),
    .A(net1062),
    .Y(_1400_));
 sg13g2_o21ai_1 _4566_ (.B1(_1400_),
    .Y(_0193_),
    .A1(_2504_),
    .A2(net569));
 sg13g2_nand3_1 _4567_ (.B(net569),
    .C(net559),
    .A(net887),
    .Y(_1401_));
 sg13g2_o21ai_1 _4568_ (.B1(_1401_),
    .Y(_0194_),
    .A1(_2503_),
    .A2(net568));
 sg13g2_nand3_1 _4569_ (.B(net568),
    .C(net557),
    .A(net1023),
    .Y(_1402_));
 sg13g2_o21ai_1 _4570_ (.B1(_1402_),
    .Y(_0195_),
    .A1(_2502_),
    .A2(net568));
 sg13g2_nand3_1 _4571_ (.B(net568),
    .C(net557),
    .A(net948),
    .Y(_1403_));
 sg13g2_o21ai_1 _4572_ (.B1(_1403_),
    .Y(_0196_),
    .A1(_2501_),
    .A2(net568));
 sg13g2_nand3_1 _4573_ (.B(net568),
    .C(net555),
    .A(net891),
    .Y(_1404_));
 sg13g2_o21ai_1 _4574_ (.B1(_1404_),
    .Y(_0197_),
    .A1(_2500_),
    .A2(net568));
 sg13g2_nand3_1 _4575_ (.B(net572),
    .C(net557),
    .A(net819),
    .Y(_1405_));
 sg13g2_o21ai_1 _4576_ (.B1(_1405_),
    .Y(_0198_),
    .A1(_2499_),
    .A2(net572));
 sg13g2_nand3_1 _4577_ (.B(net567),
    .C(net555),
    .A(net852),
    .Y(_1406_));
 sg13g2_o21ai_1 _4578_ (.B1(_1406_),
    .Y(_0199_),
    .A1(_2498_),
    .A2(net574));
 sg13g2_nand3_1 _4579_ (.B(net573),
    .C(net557),
    .A(net927),
    .Y(_1407_));
 sg13g2_o21ai_1 _4580_ (.B1(_1407_),
    .Y(_0200_),
    .A1(_2497_),
    .A2(net573));
 sg13g2_nand3_1 _4581_ (.B(net573),
    .C(net557),
    .A(net867),
    .Y(_1408_));
 sg13g2_o21ai_1 _4582_ (.B1(_1408_),
    .Y(_0201_),
    .A1(_2496_),
    .A2(net573));
 sg13g2_nand3_1 _4583_ (.B(net573),
    .C(net560),
    .A(net933),
    .Y(_1409_));
 sg13g2_o21ai_1 _4584_ (.B1(_1409_),
    .Y(_0202_),
    .A1(_2495_),
    .A2(net576));
 sg13g2_nand3_1 _4585_ (.B(net576),
    .C(net560),
    .A(net800),
    .Y(_1410_));
 sg13g2_o21ai_1 _4586_ (.B1(_1410_),
    .Y(_0203_),
    .A1(_2494_),
    .A2(net574));
 sg13g2_nand3_1 _4587_ (.B(net576),
    .C(net560),
    .A(\project_audio.iter.mult1_shift[29] ),
    .Y(_1411_));
 sg13g2_o21ai_1 _4588_ (.B1(_1411_),
    .Y(_0204_),
    .A1(_2493_),
    .A2(net574));
 sg13g2_nand3_1 _4589_ (.B(net575),
    .C(net560),
    .A(\project_audio.iter.mult1_shift[30] ),
    .Y(_1412_));
 sg13g2_o21ai_1 _4590_ (.B1(_1412_),
    .Y(_0205_),
    .A1(_2519_),
    .A2(net575));
 sg13g2_o21ai_1 _4591_ (.B1(net569),
    .Y(_1413_),
    .A1(\project_audio.iter.mult2_shift[0] ),
    .A2(net554));
 sg13g2_o21ai_1 _4592_ (.B1(net803),
    .Y(_1414_),
    .A1(_2553_),
    .A2(net547));
 sg13g2_nand2b_1 _4593_ (.Y(_1415_),
    .B(\project_audio.iter.mult1_shift[0] ),
    .A_N(net803));
 sg13g2_and3_1 _4594_ (.X(_1416_),
    .A(\project_audio.iter.mult2_shift[0] ),
    .B(net569),
    .C(net559));
 sg13g2_nand3_1 _4595_ (.B(net570),
    .C(net559),
    .A(\project_audio.iter.mult2_shift[0] ),
    .Y(_1417_));
 sg13g2_o21ai_1 _4596_ (.B1(net804),
    .Y(_0206_),
    .A1(_1415_),
    .A2(net541));
 sg13g2_nand2_1 _4597_ (.Y(_1418_),
    .A(net779),
    .B(net545));
 sg13g2_nand2_1 _4598_ (.Y(_1419_),
    .A(\project_audio.iter.mult1_shift[0] ),
    .B(\project_audio.iter.mult_accum[0] ));
 sg13g2_nand2_1 _4599_ (.Y(_1420_),
    .A(\project_audio.iter.mult1_shift[1] ),
    .B(\project_audio.iter.mult_accum[1] ));
 sg13g2_xnor2_1 _4600_ (.Y(_1421_),
    .A(\project_audio.iter.mult1_shift[1] ),
    .B(net779));
 sg13g2_xnor2_1 _4601_ (.Y(_1422_),
    .A(_1419_),
    .B(_1421_));
 sg13g2_o21ai_1 _4602_ (.B1(_1418_),
    .Y(_0207_),
    .A1(net540),
    .A2(_1422_));
 sg13g2_nand2_1 _4603_ (.Y(_1423_),
    .A(net808),
    .B(net545));
 sg13g2_o21ai_1 _4604_ (.B1(_1420_),
    .Y(_1424_),
    .A1(_1419_),
    .A2(_1421_));
 sg13g2_and2_1 _4605_ (.A(\project_audio.iter.mult1_shift[2] ),
    .B(net1244),
    .X(_1425_));
 sg13g2_xor2_1 _4606_ (.B(net808),
    .A(\project_audio.iter.mult1_shift[2] ),
    .X(_1426_));
 sg13g2_xnor2_1 _4607_ (.Y(_1427_),
    .A(_1424_),
    .B(_1426_));
 sg13g2_o21ai_1 _4608_ (.B1(_1423_),
    .Y(_0208_),
    .A1(net540),
    .A2(_1427_));
 sg13g2_nand2_1 _4609_ (.Y(_1428_),
    .A(net759),
    .B(net545));
 sg13g2_a21oi_1 _4610_ (.A1(_1424_),
    .A2(_1426_),
    .Y(_1429_),
    .B1(_1425_));
 sg13g2_nand2_1 _4611_ (.Y(_1430_),
    .A(\project_audio.iter.mult1_shift[3] ),
    .B(\project_audio.iter.mult_accum[3] ));
 sg13g2_xnor2_1 _4612_ (.Y(_1431_),
    .A(\project_audio.iter.mult1_shift[3] ),
    .B(net759));
 sg13g2_xnor2_1 _4613_ (.Y(_1432_),
    .A(_1429_),
    .B(_1431_));
 sg13g2_o21ai_1 _4614_ (.B1(_1428_),
    .Y(_0209_),
    .A1(net540),
    .A2(_1432_));
 sg13g2_nand2_1 _4615_ (.Y(_1433_),
    .A(net516),
    .B(net545));
 sg13g2_o21ai_1 _4616_ (.B1(_1430_),
    .Y(_1434_),
    .A1(_1429_),
    .A2(_1431_));
 sg13g2_and2_1 _4617_ (.A(\project_audio.iter.mult1_shift[4] ),
    .B(\project_audio.iter.mult_accum[4] ),
    .X(_1435_));
 sg13g2_xor2_1 _4618_ (.B(net516),
    .A(net1240),
    .X(_1436_));
 sg13g2_xnor2_1 _4619_ (.Y(_1437_),
    .A(_1434_),
    .B(_1436_));
 sg13g2_o21ai_1 _4620_ (.B1(_1433_),
    .Y(_0210_),
    .A1(net540),
    .A2(net1241));
 sg13g2_nand2_1 _4621_ (.Y(_1438_),
    .A(net839),
    .B(net545));
 sg13g2_a21oi_1 _4622_ (.A1(_1434_),
    .A2(_1436_),
    .Y(_1439_),
    .B1(_1435_));
 sg13g2_nor2_2 _4623_ (.A(\project_audio.iter.mult1_shift[5] ),
    .B(net839),
    .Y(_1440_));
 sg13g2_and2_1 _4624_ (.A(\project_audio.iter.mult1_shift[5] ),
    .B(\project_audio.iter.mult_accum[5] ),
    .X(_1441_));
 sg13g2_nor3_1 _4625_ (.A(_1439_),
    .B(_1440_),
    .C(_1441_),
    .Y(_1442_));
 sg13g2_o21ai_1 _4626_ (.B1(_1439_),
    .Y(_1443_),
    .A1(_1440_),
    .A2(_1441_));
 sg13g2_nand2_1 _4627_ (.Y(_1444_),
    .A(net544),
    .B(_1443_));
 sg13g2_o21ai_1 _4628_ (.B1(_1438_),
    .Y(_0211_),
    .A1(_1442_),
    .A2(_1444_));
 sg13g2_nand2_1 _4629_ (.Y(_1445_),
    .A(net730),
    .B(net545));
 sg13g2_nand2_1 _4630_ (.Y(_1446_),
    .A(\project_audio.iter.mult1_shift[6] ),
    .B(net730));
 sg13g2_xnor2_1 _4631_ (.Y(_1447_),
    .A(\project_audio.iter.mult1_shift[6] ),
    .B(net730));
 sg13g2_a221oi_1 _4632_ (.B2(_1436_),
    .C1(_1435_),
    .B1(_1434_),
    .A1(\project_audio.iter.mult1_shift[5] ),
    .Y(_1448_),
    .A2(\project_audio.iter.mult_accum[5] ));
 sg13g2_or3_1 _4633_ (.A(_1440_),
    .B(_1447_),
    .C(_1448_),
    .X(_1449_));
 sg13g2_o21ai_1 _4634_ (.B1(_1447_),
    .Y(_1450_),
    .A1(_1440_),
    .A2(_1448_));
 sg13g2_nand3_1 _4635_ (.B(_1449_),
    .C(_1450_),
    .A(net544),
    .Y(_1451_));
 sg13g2_nand2_1 _4636_ (.Y(_0212_),
    .A(_1445_),
    .B(_1451_));
 sg13g2_nand2_1 _4637_ (.Y(_1452_),
    .A(net738),
    .B(net545));
 sg13g2_and2_1 _4638_ (.A(\project_audio.iter.mult1_shift[7] ),
    .B(\project_audio.iter.mult_accum[7] ),
    .X(_1453_));
 sg13g2_xor2_1 _4639_ (.B(\project_audio.iter.mult_accum[7] ),
    .A(\project_audio.iter.mult1_shift[7] ),
    .X(_1454_));
 sg13g2_inv_1 _4640_ (.Y(_1455_),
    .A(_1454_));
 sg13g2_a21oi_1 _4641_ (.A1(_1446_),
    .A2(_1449_),
    .Y(_1456_),
    .B1(_1455_));
 sg13g2_nand3_1 _4642_ (.B(_1449_),
    .C(_1455_),
    .A(_1446_),
    .Y(_1457_));
 sg13g2_nand3b_1 _4643_ (.B(_1457_),
    .C(net544),
    .Y(_1458_),
    .A_N(_1456_));
 sg13g2_nand2_1 _4644_ (.Y(_0213_),
    .A(_1452_),
    .B(_1458_));
 sg13g2_nand2_1 _4645_ (.Y(_1459_),
    .A(net838),
    .B(net545));
 sg13g2_nor2_1 _4646_ (.A(_1453_),
    .B(_1456_),
    .Y(_1460_));
 sg13g2_xnor2_1 _4647_ (.Y(_1461_),
    .A(\project_audio.iter.mult1_shift[8] ),
    .B(\project_audio.iter.mult_accum[8] ));
 sg13g2_nor2_1 _4648_ (.A(_1460_),
    .B(_1461_),
    .Y(_1462_));
 sg13g2_a21o_1 _4649_ (.A2(_1461_),
    .A1(_1460_),
    .B1(net540),
    .X(_1463_));
 sg13g2_o21ai_1 _4650_ (.B1(_1459_),
    .Y(_0214_),
    .A1(_1462_),
    .A2(_1463_));
 sg13g2_or2_1 _4651_ (.X(_1464_),
    .B(\project_audio.iter.mult_accum[9] ),
    .A(\project_audio.iter.mult1_shift[9] ));
 sg13g2_xnor2_1 _4652_ (.Y(_1465_),
    .A(\project_audio.iter.mult1_shift[9] ),
    .B(\project_audio.iter.mult_accum[9] ));
 sg13g2_a21oi_1 _4653_ (.A1(\project_audio.iter.mult1_shift[8] ),
    .A2(\project_audio.iter.mult_accum[8] ),
    .Y(_1466_),
    .B1(_1462_));
 sg13g2_o21ai_1 _4654_ (.B1(net544),
    .Y(_1467_),
    .A1(_1465_),
    .A2(_1466_));
 sg13g2_a21oi_1 _4655_ (.A1(_1465_),
    .A2(_1466_),
    .Y(_1468_),
    .B1(_1467_));
 sg13g2_a21o_1 _4656_ (.A2(net546),
    .A1(net941),
    .B1(_1468_),
    .X(_0215_));
 sg13g2_nand2_1 _4657_ (.Y(_1469_),
    .A(net854),
    .B(net546));
 sg13g2_nor2_1 _4658_ (.A(_1461_),
    .B(_1465_),
    .Y(_1470_));
 sg13g2_o21ai_1 _4659_ (.B1(_1470_),
    .Y(_1471_),
    .A1(_1453_),
    .A2(_1456_));
 sg13g2_and3_1 _4660_ (.X(_1472_),
    .A(\project_audio.iter.mult1_shift[8] ),
    .B(\project_audio.iter.mult_accum[8] ),
    .C(_1464_));
 sg13g2_a21oi_1 _4661_ (.A1(\project_audio.iter.mult1_shift[9] ),
    .A2(\project_audio.iter.mult_accum[9] ),
    .Y(_1473_),
    .B1(_1472_));
 sg13g2_nand2_1 _4662_ (.Y(_1474_),
    .A(_1471_),
    .B(_1473_));
 sg13g2_nand2_1 _4663_ (.Y(_1475_),
    .A(\project_audio.iter.mult1_shift[10] ),
    .B(\project_audio.iter.mult_accum[10] ));
 sg13g2_xor2_1 _4664_ (.B(\project_audio.iter.mult_accum[10] ),
    .A(\project_audio.iter.mult1_shift[10] ),
    .X(_1476_));
 sg13g2_and2_1 _4665_ (.A(_1474_),
    .B(_1476_),
    .X(_1477_));
 sg13g2_o21ai_1 _4666_ (.B1(net544),
    .Y(_1478_),
    .A1(_1474_),
    .A2(_1476_));
 sg13g2_o21ai_1 _4667_ (.B1(_1469_),
    .Y(_0216_),
    .A1(_1477_),
    .A2(_1478_));
 sg13g2_nand2_1 _4668_ (.Y(_1479_),
    .A(\project_audio.iter.mult1_shift[11] ),
    .B(\project_audio.iter.mult_accum[11] ));
 sg13g2_nor2_1 _4669_ (.A(\project_audio.iter.mult1_shift[11] ),
    .B(\project_audio.iter.mult_accum[11] ),
    .Y(_1480_));
 sg13g2_xnor2_1 _4670_ (.Y(_1481_),
    .A(\project_audio.iter.mult1_shift[11] ),
    .B(net943));
 sg13g2_a21oi_1 _4671_ (.A1(\project_audio.iter.mult1_shift[10] ),
    .A2(\project_audio.iter.mult_accum[10] ),
    .Y(_1482_),
    .B1(_1477_));
 sg13g2_o21ai_1 _4672_ (.B1(net544),
    .Y(_1483_),
    .A1(_1481_),
    .A2(_1482_));
 sg13g2_a21oi_1 _4673_ (.A1(_1481_),
    .A2(_1482_),
    .Y(_1484_),
    .B1(_1483_));
 sg13g2_a21o_1 _4674_ (.A2(net546),
    .A1(net943),
    .B1(_1484_),
    .X(_0217_));
 sg13g2_nand3b_1 _4675_ (.B(_1476_),
    .C(_1479_),
    .Y(_1485_),
    .A_N(_1480_));
 sg13g2_a21oi_1 _4676_ (.A1(_1471_),
    .A2(_1473_),
    .Y(_1486_),
    .B1(_1485_));
 sg13g2_o21ai_1 _4677_ (.B1(_1479_),
    .Y(_1487_),
    .A1(_1475_),
    .A2(_1480_));
 sg13g2_nor2_1 _4678_ (.A(_1486_),
    .B(_1487_),
    .Y(_1488_));
 sg13g2_xnor2_1 _4679_ (.Y(_1489_),
    .A(\project_audio.iter.mult1_shift[12] ),
    .B(\project_audio.iter.mult_accum[12] ));
 sg13g2_nor2_1 _4680_ (.A(_1488_),
    .B(_1489_),
    .Y(_1490_));
 sg13g2_o21ai_1 _4681_ (.B1(net544),
    .Y(_1491_),
    .A1(_1488_),
    .A2(_1489_));
 sg13g2_a21oi_1 _4682_ (.A1(_1488_),
    .A2(_1489_),
    .Y(_1492_),
    .B1(_1491_));
 sg13g2_a21o_1 _4683_ (.A2(net546),
    .A1(net992),
    .B1(_1492_),
    .X(_0218_));
 sg13g2_nor2_1 _4684_ (.A(\project_audio.iter.mult1_shift[13] ),
    .B(\project_audio.iter.mult_accum[13] ),
    .Y(_1493_));
 sg13g2_xnor2_1 _4685_ (.Y(_1494_),
    .A(\project_audio.iter.mult1_shift[13] ),
    .B(\project_audio.iter.mult_accum[13] ));
 sg13g2_a21oi_1 _4686_ (.A1(net1242),
    .A2(\project_audio.iter.mult_accum[12] ),
    .Y(_1495_),
    .B1(_1490_));
 sg13g2_o21ai_1 _4687_ (.B1(net544),
    .Y(_1496_),
    .A1(_1494_),
    .A2(_1495_));
 sg13g2_a21oi_1 _4688_ (.A1(_1494_),
    .A2(_1495_),
    .Y(_1497_),
    .B1(_1496_));
 sg13g2_a21o_1 _4689_ (.A2(net546),
    .A1(net952),
    .B1(_1497_),
    .X(_0219_));
 sg13g2_nand2_1 _4690_ (.Y(_1498_),
    .A(net811),
    .B(net548));
 sg13g2_nor2_1 _4691_ (.A(\project_audio.iter.mult1_shift[14] ),
    .B(\project_audio.iter.mult_accum[14] ),
    .Y(_1499_));
 sg13g2_nand2_1 _4692_ (.Y(_1500_),
    .A(\project_audio.iter.mult1_shift[14] ),
    .B(\project_audio.iter.mult_accum[14] ));
 sg13g2_nor2b_1 _4693_ (.A(_1499_),
    .B_N(_1500_),
    .Y(_1501_));
 sg13g2_nor2_1 _4694_ (.A(_1489_),
    .B(_1494_),
    .Y(_1502_));
 sg13g2_o21ai_1 _4695_ (.B1(_1502_),
    .Y(_1503_),
    .A1(_1486_),
    .A2(_1487_));
 sg13g2_a22oi_1 _4696_ (.Y(_1504_),
    .B1(\project_audio.iter.mult_accum[13] ),
    .B2(\project_audio.iter.mult1_shift[13] ),
    .A2(\project_audio.iter.mult_accum[12] ),
    .A1(\project_audio.iter.mult1_shift[12] ));
 sg13g2_nor2_1 _4697_ (.A(_1493_),
    .B(_1504_),
    .Y(_1505_));
 sg13g2_o21ai_1 _4698_ (.B1(_1503_),
    .Y(_1506_),
    .A1(_1493_),
    .A2(_1504_));
 sg13g2_and2_1 _4699_ (.A(_1501_),
    .B(_1506_),
    .X(_1507_));
 sg13g2_o21ai_1 _4700_ (.B1(net542),
    .Y(_1508_),
    .A1(_1501_),
    .A2(_1506_));
 sg13g2_o21ai_1 _4701_ (.B1(_1498_),
    .Y(_0220_),
    .A1(_1507_),
    .A2(_1508_));
 sg13g2_nand2_1 _4702_ (.Y(_1509_),
    .A(net770),
    .B(net548));
 sg13g2_nor2_1 _4703_ (.A(\project_audio.iter.mult1_shift[15] ),
    .B(\project_audio.iter.mult_accum[15] ),
    .Y(_1510_));
 sg13g2_and2_1 _4704_ (.A(\project_audio.iter.mult1_shift[15] ),
    .B(\project_audio.iter.mult_accum[15] ),
    .X(_1511_));
 sg13g2_nand2_1 _4705_ (.Y(_1512_),
    .A(\project_audio.iter.mult1_shift[15] ),
    .B(\project_audio.iter.mult_accum[15] ));
 sg13g2_a21oi_1 _4706_ (.A1(\project_audio.iter.mult1_shift[14] ),
    .A2(\project_audio.iter.mult_accum[14] ),
    .Y(_1513_),
    .B1(_1507_));
 sg13g2_nor3_1 _4707_ (.A(_1510_),
    .B(_1511_),
    .C(_1513_),
    .Y(_1514_));
 sg13g2_o21ai_1 _4708_ (.B1(_1513_),
    .Y(_1515_),
    .A1(_1510_),
    .A2(_1511_));
 sg13g2_nand2_1 _4709_ (.Y(_1516_),
    .A(net542),
    .B(_1515_));
 sg13g2_o21ai_1 _4710_ (.B1(_1509_),
    .Y(_0221_),
    .A1(_1514_),
    .A2(_1516_));
 sg13g2_a21oi_1 _4711_ (.A1(_1500_),
    .A2(_1512_),
    .Y(_1517_),
    .B1(_1510_));
 sg13g2_nor2_1 _4712_ (.A(_1505_),
    .B(_1517_),
    .Y(_1518_));
 sg13g2_a221oi_1 _4713_ (.B2(_1503_),
    .C1(_1510_),
    .B1(_1518_),
    .A1(_1499_),
    .Y(_1519_),
    .A2(_1512_));
 sg13g2_xor2_1 _4714_ (.B(\project_audio.iter.mult1_shift[16] ),
    .A(\project_audio.iter.mult_accum[16] ),
    .X(_1520_));
 sg13g2_nand2_1 _4715_ (.Y(_1521_),
    .A(_1519_),
    .B(_1520_));
 sg13g2_o21ai_1 _4716_ (.B1(net542),
    .Y(_1522_),
    .A1(_1519_),
    .A2(_1520_));
 sg13g2_nor2b_1 _4717_ (.A(_1522_),
    .B_N(_1521_),
    .Y(_1523_));
 sg13g2_a21o_1 _4718_ (.A2(net549),
    .A1(net1082),
    .B1(_1523_),
    .X(_0222_));
 sg13g2_nor2_1 _4719_ (.A(\project_audio.iter.mult_accum[17] ),
    .B(\project_audio.iter.mult1_shift[17] ),
    .Y(_1524_));
 sg13g2_xor2_1 _4720_ (.B(\project_audio.iter.mult1_shift[17] ),
    .A(\project_audio.iter.mult_accum[17] ),
    .X(_1525_));
 sg13g2_o21ai_1 _4721_ (.B1(_1521_),
    .Y(_1526_),
    .A1(_2470_),
    .A2(_2516_));
 sg13g2_o21ai_1 _4722_ (.B1(net542),
    .Y(_1527_),
    .A1(_1525_),
    .A2(_1526_));
 sg13g2_a21oi_1 _4723_ (.A1(_1525_),
    .A2(_1526_),
    .Y(_1528_),
    .B1(_1527_));
 sg13g2_a21o_1 _4724_ (.A2(net547),
    .A1(net1194),
    .B1(_1528_),
    .X(_0223_));
 sg13g2_nand2_1 _4725_ (.Y(_1529_),
    .A(net1176),
    .B(net547));
 sg13g2_xor2_1 _4726_ (.B(\project_audio.iter.mult1_shift[18] ),
    .A(\project_audio.iter.mult_accum[18] ),
    .X(_1530_));
 sg13g2_a22oi_1 _4727_ (.Y(_1531_),
    .B1(\project_audio.iter.mult1_shift[16] ),
    .B2(\project_audio.iter.mult_accum[16] ),
    .A2(\project_audio.iter.mult1_shift[17] ),
    .A1(\project_audio.iter.mult_accum[17] ));
 sg13g2_a21oi_1 _4728_ (.A1(_1521_),
    .A2(_1531_),
    .Y(_1532_),
    .B1(_1524_));
 sg13g2_and2_1 _4729_ (.A(_1530_),
    .B(_1532_),
    .X(_1533_));
 sg13g2_o21ai_1 _4730_ (.B1(net542),
    .Y(_1534_),
    .A1(_1530_),
    .A2(_1532_));
 sg13g2_o21ai_1 _4731_ (.B1(_1529_),
    .Y(_0224_),
    .A1(_1533_),
    .A2(_1534_));
 sg13g2_nor2_1 _4732_ (.A(\project_audio.iter.mult_accum[19] ),
    .B(\project_audio.iter.mult1_shift[19] ),
    .Y(_1535_));
 sg13g2_xnor2_1 _4733_ (.Y(_1536_),
    .A(\project_audio.iter.mult_accum[19] ),
    .B(\project_audio.iter.mult1_shift[19] ));
 sg13g2_inv_1 _4734_ (.Y(_1537_),
    .A(_1536_));
 sg13g2_a21oi_1 _4735_ (.A1(\project_audio.iter.mult_accum[18] ),
    .A2(\project_audio.iter.mult1_shift[18] ),
    .Y(_1538_),
    .B1(_1533_));
 sg13g2_o21ai_1 _4736_ (.B1(net542),
    .Y(_1539_),
    .A1(_1536_),
    .A2(_1538_));
 sg13g2_a21oi_1 _4737_ (.A1(_1536_),
    .A2(_1538_),
    .Y(_1540_),
    .B1(_1539_));
 sg13g2_a21o_1 _4738_ (.A2(net547),
    .A1(net1185),
    .B1(_1540_),
    .X(_0225_));
 sg13g2_and4_1 _4739_ (.A(_1520_),
    .B(_1525_),
    .C(_1530_),
    .D(_1537_),
    .X(_1541_));
 sg13g2_a22oi_1 _4740_ (.Y(_1542_),
    .B1(\project_audio.iter.mult1_shift[18] ),
    .B2(\project_audio.iter.mult_accum[18] ),
    .A2(\project_audio.iter.mult1_shift[19] ),
    .A1(\project_audio.iter.mult_accum[19] ));
 sg13g2_nor2_1 _4741_ (.A(_1524_),
    .B(_1531_),
    .Y(_1543_));
 sg13g2_nand3_1 _4742_ (.B(_1537_),
    .C(_1543_),
    .A(_1530_),
    .Y(_1544_));
 sg13g2_o21ai_1 _4743_ (.B1(_1544_),
    .Y(_1545_),
    .A1(_1535_),
    .A2(_1542_));
 sg13g2_a21oi_1 _4744_ (.A1(_1519_),
    .A2(_1541_),
    .Y(_1546_),
    .B1(_1545_));
 sg13g2_nand2_1 _4745_ (.Y(_1547_),
    .A(\project_audio.iter.mult_accum[20] ),
    .B(\project_audio.iter.mult1_shift[20] ));
 sg13g2_xnor2_1 _4746_ (.Y(_1548_),
    .A(\project_audio.iter.mult_accum[20] ),
    .B(\project_audio.iter.mult1_shift[20] ));
 sg13g2_or2_1 _4747_ (.X(_1549_),
    .B(_1548_),
    .A(_1546_));
 sg13g2_a21oi_1 _4748_ (.A1(_1546_),
    .A2(_1548_),
    .Y(_1550_),
    .B1(net541));
 sg13g2_a22oi_1 _4749_ (.Y(_1551_),
    .B1(_1549_),
    .B2(_1550_),
    .A2(net547),
    .A1(net1205));
 sg13g2_inv_1 _4750_ (.Y(_0226_),
    .A(_1551_));
 sg13g2_nand2_1 _4751_ (.Y(_1552_),
    .A(net1177),
    .B(net547));
 sg13g2_nor2_1 _4752_ (.A(\project_audio.iter.mult_accum[21] ),
    .B(\project_audio.iter.mult1_shift[21] ),
    .Y(_1553_));
 sg13g2_xnor2_1 _4753_ (.Y(_1554_),
    .A(\project_audio.iter.mult_accum[21] ),
    .B(\project_audio.iter.mult1_shift[21] ));
 sg13g2_and2_1 _4754_ (.A(_1547_),
    .B(_1549_),
    .X(_1555_));
 sg13g2_a21oi_1 _4755_ (.A1(_1554_),
    .A2(_1555_),
    .Y(_1556_),
    .B1(net541));
 sg13g2_o21ai_1 _4756_ (.B1(_1556_),
    .Y(_1557_),
    .A1(_1554_),
    .A2(_1555_));
 sg13g2_nand2_1 _4757_ (.Y(_0227_),
    .A(_1552_),
    .B(_1557_));
 sg13g2_nand2_1 _4758_ (.Y(_1558_),
    .A(net1162),
    .B(net547));
 sg13g2_nand2_1 _4759_ (.Y(_1559_),
    .A(\project_audio.iter.mult_accum[22] ),
    .B(\project_audio.iter.mult1_shift[22] ));
 sg13g2_xnor2_1 _4760_ (.Y(_1560_),
    .A(\project_audio.iter.mult_accum[22] ),
    .B(\project_audio.iter.mult1_shift[22] ));
 sg13g2_a22oi_1 _4761_ (.Y(_1561_),
    .B1(\project_audio.iter.mult1_shift[20] ),
    .B2(\project_audio.iter.mult_accum[20] ),
    .A2(\project_audio.iter.mult1_shift[21] ),
    .A1(\project_audio.iter.mult_accum[21] ));
 sg13g2_a21o_1 _4762_ (.A2(_1561_),
    .A1(_1549_),
    .B1(_1553_),
    .X(_1562_));
 sg13g2_nor2_1 _4763_ (.A(_1560_),
    .B(_1562_),
    .Y(_1563_));
 sg13g2_a21o_1 _4764_ (.A2(_1562_),
    .A1(_1560_),
    .B1(net541),
    .X(_1564_));
 sg13g2_o21ai_1 _4765_ (.B1(_1558_),
    .Y(_0228_),
    .A1(_1563_),
    .A2(_1564_));
 sg13g2_nor2_1 _4766_ (.A(\project_audio.iter.mult_accum[23] ),
    .B(\project_audio.iter.mult1_shift[23] ),
    .Y(_1565_));
 sg13g2_nand2_1 _4767_ (.Y(_1566_),
    .A(\project_audio.iter.mult_accum[23] ),
    .B(\project_audio.iter.mult1_shift[23] ));
 sg13g2_nand2b_1 _4768_ (.Y(_1567_),
    .B(_1566_),
    .A_N(_1565_));
 sg13g2_a21oi_1 _4769_ (.A1(\project_audio.iter.mult_accum[22] ),
    .A2(\project_audio.iter.mult1_shift[22] ),
    .Y(_1568_),
    .B1(_1563_));
 sg13g2_o21ai_1 _4770_ (.B1(net542),
    .Y(_1569_),
    .A1(_1567_),
    .A2(_1568_));
 sg13g2_a21oi_1 _4771_ (.A1(_1567_),
    .A2(_1568_),
    .Y(_1570_),
    .B1(_1569_));
 sg13g2_a21o_1 _4772_ (.A2(net547),
    .A1(net1169),
    .B1(_1570_),
    .X(_0229_));
 sg13g2_nand2_1 _4773_ (.Y(_1571_),
    .A(net1006),
    .B(net549));
 sg13g2_or4_1 _4774_ (.A(_1548_),
    .B(_1554_),
    .C(_1560_),
    .D(_1567_),
    .X(_1572_));
 sg13g2_nor4_1 _4775_ (.A(_1553_),
    .B(_1560_),
    .C(_1561_),
    .D(_1567_),
    .Y(_1573_));
 sg13g2_o21ai_1 _4776_ (.B1(_1566_),
    .Y(_1574_),
    .A1(_1559_),
    .A2(_1565_));
 sg13g2_nor2_1 _4777_ (.A(_1573_),
    .B(_1574_),
    .Y(_1575_));
 sg13g2_o21ai_1 _4778_ (.B1(_1575_),
    .Y(_1576_),
    .A1(_1546_),
    .A2(_1572_));
 sg13g2_nand2_1 _4779_ (.Y(_1577_),
    .A(\project_audio.iter.mult_accum[24] ),
    .B(\project_audio.iter.mult1_shift[24] ));
 sg13g2_xor2_1 _4780_ (.B(\project_audio.iter.mult1_shift[24] ),
    .A(\project_audio.iter.mult_accum[24] ),
    .X(_1578_));
 sg13g2_inv_1 _4781_ (.Y(_1579_),
    .A(_1578_));
 sg13g2_nand2_1 _4782_ (.Y(_1580_),
    .A(_1576_),
    .B(_1578_));
 sg13g2_xnor2_1 _4783_ (.Y(_1581_),
    .A(_1576_),
    .B(_1578_));
 sg13g2_o21ai_1 _4784_ (.B1(_1571_),
    .Y(_0230_),
    .A1(net540),
    .A2(_1581_));
 sg13g2_nor2_1 _4785_ (.A(\project_audio.iter.mult_accum[25] ),
    .B(\project_audio.iter.mult1_shift[25] ),
    .Y(_1582_));
 sg13g2_xnor2_1 _4786_ (.Y(_1583_),
    .A(\project_audio.iter.mult_accum[25] ),
    .B(\project_audio.iter.mult1_shift[25] ));
 sg13g2_and2_1 _4787_ (.A(_1577_),
    .B(_1580_),
    .X(_1584_));
 sg13g2_o21ai_1 _4788_ (.B1(net542),
    .Y(_1585_),
    .A1(_1583_),
    .A2(_1584_));
 sg13g2_a21oi_1 _4789_ (.A1(_1583_),
    .A2(_1584_),
    .Y(_1586_),
    .B1(_1585_));
 sg13g2_a21o_1 _4790_ (.A2(net549),
    .A1(net1184),
    .B1(_1586_),
    .X(_0231_));
 sg13g2_nand2_1 _4791_ (.Y(_1587_),
    .A(net901),
    .B(net548));
 sg13g2_nor2_1 _4792_ (.A(_1579_),
    .B(_1583_),
    .Y(_1588_));
 sg13g2_nor2_1 _4793_ (.A(_1577_),
    .B(_1582_),
    .Y(_1589_));
 sg13g2_a221oi_1 _4794_ (.B2(_1588_),
    .C1(_1589_),
    .B1(_1576_),
    .A1(\project_audio.iter.mult_accum[25] ),
    .Y(_1590_),
    .A2(\project_audio.iter.mult1_shift[25] ));
 sg13g2_nand2_1 _4795_ (.Y(_1591_),
    .A(\project_audio.iter.mult_accum[26] ),
    .B(\project_audio.iter.mult1_shift[26] ));
 sg13g2_xnor2_1 _4796_ (.Y(_1592_),
    .A(\project_audio.iter.mult_accum[26] ),
    .B(net931));
 sg13g2_xnor2_1 _4797_ (.Y(_1593_),
    .A(_1590_),
    .B(net932));
 sg13g2_o21ai_1 _4798_ (.B1(_1587_),
    .Y(_0232_),
    .A1(net540),
    .A2(_1593_));
 sg13g2_nor2_1 _4799_ (.A(\project_audio.iter.mult_accum[27] ),
    .B(\project_audio.iter.mult1_shift[27] ),
    .Y(_1594_));
 sg13g2_xor2_1 _4800_ (.B(\project_audio.iter.mult1_shift[27] ),
    .A(\project_audio.iter.mult_accum[27] ),
    .X(_1595_));
 sg13g2_o21ai_1 _4801_ (.B1(_1591_),
    .Y(_1596_),
    .A1(_1590_),
    .A2(_1592_));
 sg13g2_o21ai_1 _4802_ (.B1(net543),
    .Y(_1597_),
    .A1(_1595_),
    .A2(_1596_));
 sg13g2_a21oi_1 _4803_ (.A1(_1595_),
    .A2(_1596_),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_a21o_1 _4804_ (.A2(net548),
    .A1(net1181),
    .B1(_1598_),
    .X(_0233_));
 sg13g2_and2_1 _4805_ (.A(\project_audio.iter.mult_accum[28] ),
    .B(\project_audio.iter.mult1_shift[28] ),
    .X(_1599_));
 sg13g2_xor2_1 _4806_ (.B(\project_audio.iter.mult1_shift[28] ),
    .A(\project_audio.iter.mult_accum[28] ),
    .X(_1600_));
 sg13g2_nand2b_1 _4807_ (.Y(_1601_),
    .B(_1595_),
    .A_N(_1592_));
 sg13g2_or2_1 _4808_ (.X(_1602_),
    .B(_1594_),
    .A(_1591_));
 sg13g2_inv_1 _4809_ (.Y(_1603_),
    .A(_1602_));
 sg13g2_a21oi_1 _4810_ (.A1(\project_audio.iter.mult_accum[27] ),
    .A2(\project_audio.iter.mult1_shift[27] ),
    .Y(_1604_),
    .B1(_1603_));
 sg13g2_o21ai_1 _4811_ (.B1(_1604_),
    .Y(_1605_),
    .A1(_1590_),
    .A2(_1601_));
 sg13g2_o21ai_1 _4812_ (.B1(net543),
    .Y(_1606_),
    .A1(_1600_),
    .A2(_1605_));
 sg13g2_a21oi_1 _4813_ (.A1(_1600_),
    .A2(_1605_),
    .Y(_1607_),
    .B1(_1606_));
 sg13g2_a21o_1 _4814_ (.A2(net548),
    .A1(net1146),
    .B1(_1607_),
    .X(_0234_));
 sg13g2_nand2_1 _4815_ (.Y(_1608_),
    .A(net1106),
    .B(net548));
 sg13g2_a21oi_1 _4816_ (.A1(_1600_),
    .A2(_1605_),
    .Y(_1609_),
    .B1(_1599_));
 sg13g2_nor2_1 _4817_ (.A(\project_audio.iter.mult_accum[29] ),
    .B(\project_audio.iter.mult1_shift[29] ),
    .Y(_1610_));
 sg13g2_xnor2_1 _4818_ (.Y(_1611_),
    .A(\project_audio.iter.mult_accum[29] ),
    .B(\project_audio.iter.mult1_shift[29] ));
 sg13g2_xnor2_1 _4819_ (.Y(_1612_),
    .A(_1609_),
    .B(_1611_));
 sg13g2_o21ai_1 _4820_ (.B1(_1608_),
    .Y(_0235_),
    .A1(net540),
    .A2(_1612_));
 sg13g2_nand2_1 _4821_ (.Y(_1613_),
    .A(net949),
    .B(net548));
 sg13g2_xnor2_1 _4822_ (.Y(_1614_),
    .A(\project_audio.iter.mult_accum[30] ),
    .B(\project_audio.iter.mult1_shift[30] ));
 sg13g2_a221oi_1 _4823_ (.B2(_1605_),
    .C1(_1599_),
    .B1(_1600_),
    .A1(\project_audio.iter.mult_accum[29] ),
    .Y(_1615_),
    .A2(\project_audio.iter.mult1_shift[29] ));
 sg13g2_nor3_1 _4824_ (.A(_1610_),
    .B(_1614_),
    .C(_1615_),
    .Y(_1616_));
 sg13g2_o21ai_1 _4825_ (.B1(_1614_),
    .Y(_1617_),
    .A1(_1610_),
    .A2(_1615_));
 sg13g2_nand2_1 _4826_ (.Y(_1618_),
    .A(net543),
    .B(_1617_));
 sg13g2_o21ai_1 _4827_ (.B1(_1613_),
    .Y(_0236_),
    .A1(_1616_),
    .A2(_1618_));
 sg13g2_nand2_1 _4828_ (.Y(_1619_),
    .A(net1030),
    .B(net548));
 sg13g2_a21oi_1 _4829_ (.A1(\project_audio.iter.mult_accum[30] ),
    .A2(\project_audio.iter.mult1_shift[30] ),
    .Y(_1620_),
    .B1(_1616_));
 sg13g2_xor2_1 _4830_ (.B(net760),
    .A(\project_audio.iter.mult_accum[31] ),
    .X(_1621_));
 sg13g2_inv_1 _4831_ (.Y(_1622_),
    .A(_1621_));
 sg13g2_and2_1 _4832_ (.A(_1620_),
    .B(_1622_),
    .X(_1623_));
 sg13g2_o21ai_1 _4833_ (.B1(net543),
    .Y(_1624_),
    .A1(_1620_),
    .A2(_1622_));
 sg13g2_o21ai_1 _4834_ (.B1(_1619_),
    .Y(_0237_),
    .A1(_1623_),
    .A2(_1624_));
 sg13g2_nor2b_1 _4835_ (.A(net535),
    .B_N(net633),
    .Y(_1625_));
 sg13g2_o21ai_1 _4836_ (.B1(net700),
    .Y(_1626_),
    .A1(net638),
    .A2(net908));
 sg13g2_nor2_1 _4837_ (.A(_1625_),
    .B(_1626_),
    .Y(_0238_));
 sg13g2_nand2_1 _4838_ (.Y(_1627_),
    .A(net652),
    .B(net528));
 sg13g2_nand2_1 _4839_ (.Y(_1628_),
    .A(net958),
    .B(net528));
 sg13g2_xor2_1 _4840_ (.B(_1627_),
    .A(net958),
    .X(_1629_));
 sg13g2_nor2_1 _4841_ (.A(net684),
    .B(_1629_),
    .Y(_0239_));
 sg13g2_nand2_1 _4842_ (.Y(_1630_),
    .A(\project_audio.genblk1[7].n_c_oh_my.phase[1] ),
    .B(\project_audio.freq[7][1] ));
 sg13g2_xnor2_1 _4843_ (.Y(_1631_),
    .A(net1014),
    .B(net777));
 sg13g2_xnor2_1 _4844_ (.Y(_1632_),
    .A(_1628_),
    .B(_1631_));
 sg13g2_o21ai_1 _4845_ (.B1(net701),
    .Y(_1633_),
    .A1(net652),
    .A2(net1014));
 sg13g2_a21oi_1 _4846_ (.A1(net652),
    .A2(_1632_),
    .Y(_0240_),
    .B1(_1633_));
 sg13g2_o21ai_1 _4847_ (.B1(_1630_),
    .Y(_1634_),
    .A1(_1628_),
    .A2(_1631_));
 sg13g2_and2_1 _4848_ (.A(\project_audio.genblk1[7].n_c_oh_my.phase[2] ),
    .B(\project_audio.freq[7][2] ),
    .X(_1635_));
 sg13g2_xor2_1 _4849_ (.B(net778),
    .A(net981),
    .X(_1636_));
 sg13g2_xnor2_1 _4850_ (.Y(_1637_),
    .A(_1634_),
    .B(_1636_));
 sg13g2_o21ai_1 _4851_ (.B1(net702),
    .Y(_1638_),
    .A1(net652),
    .A2(net981));
 sg13g2_a21oi_1 _4852_ (.A1(net652),
    .A2(_1637_),
    .Y(_0241_),
    .B1(_1638_));
 sg13g2_a21oi_1 _4853_ (.A1(_1634_),
    .A2(_1636_),
    .Y(_1639_),
    .B1(_1635_));
 sg13g2_nand2_1 _4854_ (.Y(_1640_),
    .A(\project_audio.genblk1[7].n_c_oh_my.phase[3] ),
    .B(\project_audio.freq[7][3] ));
 sg13g2_xnor2_1 _4855_ (.Y(_1641_),
    .A(net1040),
    .B(net806));
 sg13g2_xnor2_1 _4856_ (.Y(_1642_),
    .A(_1639_),
    .B(_1641_));
 sg13g2_o21ai_1 _4857_ (.B1(net702),
    .Y(_1643_),
    .A1(net657),
    .A2(net1040));
 sg13g2_a21oi_1 _4858_ (.A1(net657),
    .A2(_1642_),
    .Y(_0242_),
    .B1(_1643_));
 sg13g2_o21ai_1 _4859_ (.B1(_1640_),
    .Y(_1644_),
    .A1(_1639_),
    .A2(_1641_));
 sg13g2_and2_1 _4860_ (.A(\project_audio.genblk1[7].n_c_oh_my.phase[4] ),
    .B(\project_audio.freq[7][4] ),
    .X(_1645_));
 sg13g2_xor2_1 _4861_ (.B(net499),
    .A(net1068),
    .X(_1646_));
 sg13g2_xnor2_1 _4862_ (.Y(_1647_),
    .A(_1644_),
    .B(_1646_));
 sg13g2_o21ai_1 _4863_ (.B1(net702),
    .Y(_1648_),
    .A1(net653),
    .A2(net1068));
 sg13g2_a21oi_1 _4864_ (.A1(net653),
    .A2(_1647_),
    .Y(_0243_),
    .B1(_1648_));
 sg13g2_a21o_1 _4865_ (.A2(_1646_),
    .A1(_1644_),
    .B1(_1645_),
    .X(_1649_));
 sg13g2_or2_1 _4866_ (.X(_1650_),
    .B(\project_audio.freq[7][5] ),
    .A(\project_audio.genblk1[7].n_c_oh_my.phase[5] ));
 sg13g2_and2_1 _4867_ (.A(\project_audio.genblk1[7].n_c_oh_my.phase[5] ),
    .B(\project_audio.freq[7][5] ),
    .X(_1651_));
 sg13g2_xnor2_1 _4868_ (.Y(_1652_),
    .A(net1174),
    .B(net810));
 sg13g2_o21ai_1 _4869_ (.B1(net653),
    .Y(_1653_),
    .A1(_1649_),
    .A2(_1652_));
 sg13g2_a21oi_1 _4870_ (.A1(_1649_),
    .A2(_1652_),
    .Y(_1654_),
    .B1(_1653_));
 sg13g2_o21ai_1 _4871_ (.B1(net702),
    .Y(_1655_),
    .A1(net653),
    .A2(net1174));
 sg13g2_nor2_1 _4872_ (.A(_1654_),
    .B(_1655_),
    .Y(_0244_));
 sg13g2_xnor2_1 _4873_ (.Y(_1656_),
    .A(\project_audio.genblk1[7].n_c_oh_my.phase[6] ),
    .B(net829));
 sg13g2_a21oi_1 _4874_ (.A1(_1649_),
    .A2(_1650_),
    .Y(_1657_),
    .B1(_1651_));
 sg13g2_nor2_1 _4875_ (.A(_1656_),
    .B(_1657_),
    .Y(_1658_));
 sg13g2_xnor2_1 _4876_ (.Y(_1659_),
    .A(_1656_),
    .B(_1657_));
 sg13g2_o21ai_1 _4877_ (.B1(net702),
    .Y(_1660_),
    .A1(net653),
    .A2(net1115));
 sg13g2_a21oi_1 _4878_ (.A1(net653),
    .A2(_1659_),
    .Y(_0245_),
    .B1(_1660_));
 sg13g2_a21oi_1 _4879_ (.A1(\project_audio.genblk1[7].n_c_oh_my.phase[6] ),
    .A2(net829),
    .Y(_1661_),
    .B1(_1658_));
 sg13g2_nand2_1 _4880_ (.Y(_1662_),
    .A(net989),
    .B(net727));
 sg13g2_xnor2_1 _4881_ (.Y(_1663_),
    .A(net989),
    .B(net727));
 sg13g2_or2_1 _4882_ (.X(_1664_),
    .B(_1663_),
    .A(_1661_));
 sg13g2_xnor2_1 _4883_ (.Y(_1665_),
    .A(_1661_),
    .B(_1663_));
 sg13g2_o21ai_1 _4884_ (.B1(net702),
    .Y(_1666_),
    .A1(net654),
    .A2(net989));
 sg13g2_a21oi_1 _4885_ (.A1(net654),
    .A2(_1665_),
    .Y(_0246_),
    .B1(_1666_));
 sg13g2_xnor2_1 _4886_ (.Y(_1667_),
    .A(\project_audio.genblk1[7].n_c_oh_my.phase[8] ),
    .B(\project_audio.freq[7][8] ));
 sg13g2_a21oi_1 _4887_ (.A1(_1662_),
    .A2(_1664_),
    .Y(_1668_),
    .B1(_1667_));
 sg13g2_nand3_1 _4888_ (.B(_1664_),
    .C(_1667_),
    .A(_1662_),
    .Y(_1669_));
 sg13g2_nand2b_1 _4889_ (.Y(_1670_),
    .B(_1669_),
    .A_N(_1668_));
 sg13g2_o21ai_1 _4890_ (.B1(net702),
    .Y(_1671_),
    .A1(net654),
    .A2(net1086));
 sg13g2_a21oi_1 _4891_ (.A1(net654),
    .A2(_1670_),
    .Y(_0247_),
    .B1(_1671_));
 sg13g2_a21o_1 _4892_ (.A2(\project_audio.freq[7][8] ),
    .A1(\project_audio.genblk1[7].n_c_oh_my.phase[8] ),
    .B1(_1668_),
    .X(_1672_));
 sg13g2_nor2_1 _4893_ (.A(\project_audio.genblk1[7].n_c_oh_my.phase[9] ),
    .B(\project_audio.freq[7][9] ),
    .Y(_1673_));
 sg13g2_xor2_1 _4894_ (.B(net851),
    .A(net1114),
    .X(_1674_));
 sg13g2_xnor2_1 _4895_ (.Y(_1675_),
    .A(_1672_),
    .B(_1674_));
 sg13g2_o21ai_1 _4896_ (.B1(net701),
    .Y(_1676_),
    .A1(net653),
    .A2(net1114));
 sg13g2_a21oi_1 _4897_ (.A1(net652),
    .A2(_1675_),
    .Y(_0248_),
    .B1(_1676_));
 sg13g2_xnor2_1 _4898_ (.Y(_1677_),
    .A(net1017),
    .B(net717));
 sg13g2_a21oi_1 _4899_ (.A1(\project_audio.genblk1[7].n_c_oh_my.phase[9] ),
    .A2(\project_audio.freq[7][9] ),
    .Y(_1678_),
    .B1(_1672_));
 sg13g2_nor3_1 _4900_ (.A(_1673_),
    .B(_1677_),
    .C(_1678_),
    .Y(_1679_));
 sg13g2_o21ai_1 _4901_ (.B1(_1677_),
    .Y(_1680_),
    .A1(_1673_),
    .A2(_1678_));
 sg13g2_nand2b_1 _4902_ (.Y(_1681_),
    .B(_1680_),
    .A_N(_1679_));
 sg13g2_o21ai_1 _4903_ (.B1(net701),
    .Y(_1682_),
    .A1(net652),
    .A2(net1017));
 sg13g2_a21oi_1 _4904_ (.A1(net652),
    .A2(_1681_),
    .Y(_0249_),
    .B1(_1682_));
 sg13g2_a21oi_1 _4905_ (.A1(\project_audio.genblk1[7].n_c_oh_my.phase[10] ),
    .A2(net717),
    .Y(_1683_),
    .B1(_1679_));
 sg13g2_nor2_1 _4906_ (.A(\project_audio.genblk1[7].n_c_oh_my.phase[11] ),
    .B(\project_audio.freq[7][11] ),
    .Y(_1684_));
 sg13g2_nand2_1 _4907_ (.Y(_1685_),
    .A(net969),
    .B(net447));
 sg13g2_nand2b_1 _4908_ (.Y(_1686_),
    .B(_1685_),
    .A_N(_1684_));
 sg13g2_xnor2_1 _4909_ (.Y(_1687_),
    .A(_1683_),
    .B(_1686_));
 sg13g2_o21ai_1 _4910_ (.B1(net710),
    .Y(_1688_),
    .A1(net656),
    .A2(net969));
 sg13g2_a21oi_1 _4911_ (.A1(net656),
    .A2(_1687_),
    .Y(_0250_),
    .B1(_1688_));
 sg13g2_o21ai_1 _4912_ (.B1(_1685_),
    .Y(_1689_),
    .A1(_1683_),
    .A2(_1684_));
 sg13g2_a21oi_1 _4913_ (.A1(net632),
    .A2(_1689_),
    .Y(_1690_),
    .B1(net473));
 sg13g2_nand3_1 _4914_ (.B(net473),
    .C(_1689_),
    .A(net632),
    .Y(_1691_));
 sg13g2_inv_1 _4915_ (.Y(_1692_),
    .A(_1691_));
 sg13g2_nor3_1 _4916_ (.A(net680),
    .B(_1690_),
    .C(_1692_),
    .Y(_0251_));
 sg13g2_nand2_1 _4917_ (.Y(_1693_),
    .A(net524),
    .B(_1692_));
 sg13g2_nand2_1 _4918_ (.Y(_1694_),
    .A(net694),
    .B(_1693_));
 sg13g2_a21oi_1 _4919_ (.A1(_2492_),
    .A2(_1691_),
    .Y(_0252_),
    .B1(_1694_));
 sg13g2_o21ai_1 _4920_ (.B1(net694),
    .Y(_1695_),
    .A1(_2491_),
    .A2(_1693_));
 sg13g2_a21oi_1 _4921_ (.A1(_2491_),
    .A2(_1693_),
    .Y(_0253_),
    .B1(_1695_));
 sg13g2_and4_1 _4922_ (.A(\project_audio.genblk1[7].n_c_oh_my.phase[14] ),
    .B(net524),
    .C(net473),
    .D(net694),
    .X(_1696_));
 sg13g2_nand3_1 _4923_ (.B(_1689_),
    .C(_1696_),
    .A(_1625_),
    .Y(_1697_));
 sg13g2_o21ai_1 _4924_ (.B1(_1697_),
    .Y(_0254_),
    .A1(_2490_),
    .A2(_1695_));
 sg13g2_nor2b_1 _4925_ (.A(net530),
    .B_N(net640),
    .Y(_1698_));
 sg13g2_o21ai_1 _4926_ (.B1(net697),
    .Y(_1699_),
    .A1(net641),
    .A2(net957));
 sg13g2_nor2_1 _4927_ (.A(_1698_),
    .B(_1699_),
    .Y(_0255_));
 sg13g2_nand2_1 _4928_ (.Y(_1700_),
    .A(net662),
    .B(net749));
 sg13g2_nand2_1 _4929_ (.Y(_1701_),
    .A(net900),
    .B(net749));
 sg13g2_xor2_1 _4930_ (.B(_1700_),
    .A(net900),
    .X(_1702_));
 sg13g2_nor2_1 _4931_ (.A(net683),
    .B(_1702_),
    .Y(_0256_));
 sg13g2_nand2_1 _4932_ (.Y(_1703_),
    .A(\project_audio.genblk1[6].n_c_oh_my.phase[1] ),
    .B(\project_audio.freq[6][1] ));
 sg13g2_xnor2_1 _4933_ (.Y(_1704_),
    .A(net1087),
    .B(net807));
 sg13g2_xnor2_1 _4934_ (.Y(_1705_),
    .A(_1701_),
    .B(_1704_));
 sg13g2_o21ai_1 _4935_ (.B1(net712),
    .Y(_1706_),
    .A1(net664),
    .A2(net1087));
 sg13g2_a21oi_1 _4936_ (.A1(net662),
    .A2(_1705_),
    .Y(_0257_),
    .B1(_1706_));
 sg13g2_o21ai_1 _4937_ (.B1(_1703_),
    .Y(_1707_),
    .A1(_1701_),
    .A2(_1704_));
 sg13g2_and2_1 _4938_ (.A(\project_audio.genblk1[6].n_c_oh_my.phase[2] ),
    .B(\project_audio.freq[6][2] ),
    .X(_1708_));
 sg13g2_xor2_1 _4939_ (.B(net509),
    .A(\project_audio.genblk1[6].n_c_oh_my.phase[2] ),
    .X(_1709_));
 sg13g2_xnor2_1 _4940_ (.Y(_1710_),
    .A(_1707_),
    .B(_1709_));
 sg13g2_o21ai_1 _4941_ (.B1(net709),
    .Y(_1711_),
    .A1(net662),
    .A2(net1092));
 sg13g2_a21oi_1 _4942_ (.A1(net664),
    .A2(_1710_),
    .Y(_0258_),
    .B1(_1711_));
 sg13g2_a21oi_2 _4943_ (.B1(_1708_),
    .Y(_1712_),
    .A2(_1709_),
    .A1(_1707_));
 sg13g2_nand2_1 _4944_ (.Y(_1713_),
    .A(\project_audio.genblk1[6].n_c_oh_my.phase[3] ),
    .B(\project_audio.freq[6][3] ));
 sg13g2_xnor2_1 _4945_ (.Y(_1714_),
    .A(net1102),
    .B(net792));
 sg13g2_xnor2_1 _4946_ (.Y(_1715_),
    .A(_1712_),
    .B(_1714_));
 sg13g2_o21ai_1 _4947_ (.B1(net709),
    .Y(_1716_),
    .A1(net663),
    .A2(net1102));
 sg13g2_a21oi_1 _4948_ (.A1(net663),
    .A2(_1715_),
    .Y(_0259_),
    .B1(_1716_));
 sg13g2_o21ai_1 _4949_ (.B1(_1713_),
    .Y(_1717_),
    .A1(_1712_),
    .A2(_1714_));
 sg13g2_and2_1 _4950_ (.A(\project_audio.genblk1[6].n_c_oh_my.phase[4] ),
    .B(\project_audio.freq[6][4] ),
    .X(_1718_));
 sg13g2_xor2_1 _4951_ (.B(net533),
    .A(net1088),
    .X(_1719_));
 sg13g2_xnor2_1 _4952_ (.Y(_1720_),
    .A(_1717_),
    .B(_1719_));
 sg13g2_o21ai_1 _4953_ (.B1(net712),
    .Y(_1721_),
    .A1(net664),
    .A2(net1088));
 sg13g2_a21oi_1 _4954_ (.A1(net664),
    .A2(_1720_),
    .Y(_0260_),
    .B1(_1721_));
 sg13g2_a21o_1 _4955_ (.A2(_1719_),
    .A1(_1717_),
    .B1(_1718_),
    .X(_1722_));
 sg13g2_or2_1 _4956_ (.X(_1723_),
    .B(\project_audio.freq[6][5] ),
    .A(\project_audio.genblk1[6].n_c_oh_my.phase[5] ));
 sg13g2_nand2_1 _4957_ (.Y(_1724_),
    .A(net906),
    .B(net475));
 sg13g2_nand2_1 _4958_ (.Y(_1725_),
    .A(_1723_),
    .B(_1724_));
 sg13g2_xor2_1 _4959_ (.B(_1725_),
    .A(_1722_),
    .X(_1726_));
 sg13g2_o21ai_1 _4960_ (.B1(net712),
    .Y(_1727_),
    .A1(net665),
    .A2(net906));
 sg13g2_a21oi_1 _4961_ (.A1(net665),
    .A2(_1726_),
    .Y(_0261_),
    .B1(_1727_));
 sg13g2_xnor2_1 _4962_ (.Y(_1728_),
    .A(\project_audio.genblk1[6].n_c_oh_my.phase[6] ),
    .B(\project_audio.freq[6][6] ));
 sg13g2_nand2_1 _4963_ (.Y(_1729_),
    .A(_1722_),
    .B(_1723_));
 sg13g2_a21oi_1 _4964_ (.A1(_1724_),
    .A2(_1729_),
    .Y(_1730_),
    .B1(_1728_));
 sg13g2_nand3_1 _4965_ (.B(_1728_),
    .C(_1729_),
    .A(_1724_),
    .Y(_1731_));
 sg13g2_nand2b_1 _4966_ (.Y(_1732_),
    .B(_1731_),
    .A_N(_1730_));
 sg13g2_o21ai_1 _4967_ (.B1(net712),
    .Y(_1733_),
    .A1(net665),
    .A2(net1144));
 sg13g2_a21oi_1 _4968_ (.A1(net665),
    .A2(_1732_),
    .Y(_0262_),
    .B1(_1733_));
 sg13g2_a21oi_1 _4969_ (.A1(\project_audio.genblk1[6].n_c_oh_my.phase[6] ),
    .A2(net772),
    .Y(_1734_),
    .B1(_1730_));
 sg13g2_nand2_1 _4970_ (.Y(_1735_),
    .A(net1112),
    .B(net743));
 sg13g2_xnor2_1 _4971_ (.Y(_1736_),
    .A(net1112),
    .B(net743));
 sg13g2_or2_1 _4972_ (.X(_1737_),
    .B(_1736_),
    .A(_1734_));
 sg13g2_xnor2_1 _4973_ (.Y(_1738_),
    .A(_1734_),
    .B(_1736_));
 sg13g2_o21ai_1 _4974_ (.B1(net712),
    .Y(_1739_),
    .A1(net666),
    .A2(net1112));
 sg13g2_a21oi_1 _4975_ (.A1(net665),
    .A2(_1738_),
    .Y(_0263_),
    .B1(_1739_));
 sg13g2_xnor2_1 _4976_ (.Y(_1740_),
    .A(\project_audio.genblk1[6].n_c_oh_my.phase[8] ),
    .B(\project_audio.freq[6][8] ));
 sg13g2_a21oi_1 _4977_ (.A1(_1735_),
    .A2(_1737_),
    .Y(_1741_),
    .B1(_1740_));
 sg13g2_nand3_1 _4978_ (.B(_1737_),
    .C(_1740_),
    .A(_1735_),
    .Y(_1742_));
 sg13g2_nand2b_1 _4979_ (.Y(_1743_),
    .B(_1742_),
    .A_N(_1741_));
 sg13g2_o21ai_1 _4980_ (.B1(net712),
    .Y(_1744_),
    .A1(net665),
    .A2(net1149));
 sg13g2_a21oi_1 _4981_ (.A1(net667),
    .A2(_1743_),
    .Y(_0264_),
    .B1(_1744_));
 sg13g2_a21o_1 _4982_ (.A2(\project_audio.freq[6][8] ),
    .A1(\project_audio.genblk1[6].n_c_oh_my.phase[8] ),
    .B1(_1741_),
    .X(_1745_));
 sg13g2_nor2_1 _4983_ (.A(\project_audio.genblk1[6].n_c_oh_my.phase[9] ),
    .B(\project_audio.freq[6][9] ),
    .Y(_1746_));
 sg13g2_xor2_1 _4984_ (.B(net812),
    .A(net1126),
    .X(_1747_));
 sg13g2_xnor2_1 _4985_ (.Y(_1748_),
    .A(_1745_),
    .B(_1747_));
 sg13g2_o21ai_1 _4986_ (.B1(net713),
    .Y(_1749_),
    .A1(net665),
    .A2(net1126));
 sg13g2_a21oi_1 _4987_ (.A1(net665),
    .A2(_1748_),
    .Y(_0265_),
    .B1(_1749_));
 sg13g2_xnor2_1 _4988_ (.Y(_1750_),
    .A(net973),
    .B(net794));
 sg13g2_a21oi_1 _4989_ (.A1(\project_audio.genblk1[6].n_c_oh_my.phase[9] ),
    .A2(\project_audio.freq[6][9] ),
    .Y(_1751_),
    .B1(_1745_));
 sg13g2_nor3_1 _4990_ (.A(_1746_),
    .B(_1750_),
    .C(_1751_),
    .Y(_1752_));
 sg13g2_o21ai_1 _4991_ (.B1(_1750_),
    .Y(_1753_),
    .A1(_1746_),
    .A2(_1751_));
 sg13g2_nand2b_1 _4992_ (.Y(_1754_),
    .B(_1753_),
    .A_N(_1752_));
 sg13g2_o21ai_1 _4993_ (.B1(net712),
    .Y(_1755_),
    .A1(net666),
    .A2(net973));
 sg13g2_a21oi_1 _4994_ (.A1(net666),
    .A2(_1754_),
    .Y(_0266_),
    .B1(_1755_));
 sg13g2_a21oi_1 _4995_ (.A1(\project_audio.genblk1[6].n_c_oh_my.phase[10] ),
    .A2(net794),
    .Y(_1756_),
    .B1(_1752_));
 sg13g2_nor2_1 _4996_ (.A(\project_audio.genblk1[6].n_c_oh_my.phase[11] ),
    .B(\project_audio.freq[6][11] ),
    .Y(_1757_));
 sg13g2_nand2_1 _4997_ (.Y(_1758_),
    .A(net925),
    .B(net444));
 sg13g2_nand2b_1 _4998_ (.Y(_1759_),
    .B(_1758_),
    .A_N(_1757_));
 sg13g2_xnor2_1 _4999_ (.Y(_1760_),
    .A(_1756_),
    .B(_1759_));
 sg13g2_o21ai_1 _5000_ (.B1(net711),
    .Y(_1761_),
    .A1(net666),
    .A2(net925));
 sg13g2_a21oi_1 _5001_ (.A1(net666),
    .A2(_1760_),
    .Y(_0267_),
    .B1(_1761_));
 sg13g2_o21ai_1 _5002_ (.B1(_1758_),
    .Y(_1762_),
    .A1(_1756_),
    .A2(_1757_));
 sg13g2_a21oi_1 _5003_ (.A1(net640),
    .A2(_1762_),
    .Y(_1763_),
    .B1(net731));
 sg13g2_nand3_1 _5004_ (.B(net731),
    .C(_1762_),
    .A(net640),
    .Y(_1764_));
 sg13g2_inv_1 _5005_ (.Y(_1765_),
    .A(_1764_));
 sg13g2_nor3_1 _5006_ (.A(net681),
    .B(_1763_),
    .C(_1765_),
    .Y(_0268_));
 sg13g2_nand2_1 _5007_ (.Y(_1766_),
    .A(net503),
    .B(_1765_));
 sg13g2_nand2_1 _5008_ (.Y(_1767_),
    .A(net698),
    .B(_1766_));
 sg13g2_a21oi_1 _5009_ (.A1(_2489_),
    .A2(_1764_),
    .Y(_0269_),
    .B1(_1767_));
 sg13g2_o21ai_1 _5010_ (.B1(net698),
    .Y(_1768_),
    .A1(_2488_),
    .A2(_1766_));
 sg13g2_a21oi_1 _5011_ (.A1(_2488_),
    .A2(_1766_),
    .Y(_0270_),
    .B1(_1768_));
 sg13g2_and4_1 _5012_ (.A(\project_audio.genblk1[6].n_c_oh_my.phase[14] ),
    .B(net503),
    .C(\project_audio.genblk1[6].n_c_oh_my.phase[12] ),
    .D(net698),
    .X(_1769_));
 sg13g2_nand3_1 _5013_ (.B(_1762_),
    .C(_1769_),
    .A(_1698_),
    .Y(_1770_));
 sg13g2_o21ai_1 _5014_ (.B1(_1770_),
    .Y(_0271_),
    .A1(_2487_),
    .A2(_1768_));
 sg13g2_nor2b_1 _5015_ (.A(net494),
    .B_N(net632),
    .Y(_1771_));
 sg13g2_o21ai_1 _5016_ (.B1(net694),
    .Y(_1772_),
    .A1(net632),
    .A2(net837));
 sg13g2_nor2_1 _5017_ (.A(_1771_),
    .B(_1772_),
    .Y(_0272_));
 sg13g2_nand2_1 _5018_ (.Y(_1773_),
    .A(net648),
    .B(net474));
 sg13g2_nand2_1 _5019_ (.Y(_1774_),
    .A(net937),
    .B(net474));
 sg13g2_xor2_1 _5020_ (.B(_1773_),
    .A(net937),
    .X(_1775_));
 sg13g2_nor2_1 _5021_ (.A(net684),
    .B(_1775_),
    .Y(_0273_));
 sg13g2_nand2_1 _5022_ (.Y(_1776_),
    .A(\project_audio.genblk1[5].n_c_oh_my.phase[1] ),
    .B(\project_audio.freq[5][1] ));
 sg13g2_xnor2_1 _5023_ (.Y(_1777_),
    .A(net1097),
    .B(net718));
 sg13g2_xnor2_1 _5024_ (.Y(_1778_),
    .A(_1774_),
    .B(_1777_));
 sg13g2_o21ai_1 _5025_ (.B1(net703),
    .Y(_1779_),
    .A1(net648),
    .A2(net1097));
 sg13g2_a21oi_1 _5026_ (.A1(net648),
    .A2(_1778_),
    .Y(_0274_),
    .B1(_1779_));
 sg13g2_o21ai_1 _5027_ (.B1(_1776_),
    .Y(_1780_),
    .A1(_1774_),
    .A2(_1777_));
 sg13g2_and2_1 _5028_ (.A(\project_audio.genblk1[5].n_c_oh_my.phase[2] ),
    .B(\project_audio.freq[5][2] ),
    .X(_1781_));
 sg13g2_xor2_1 _5029_ (.B(net754),
    .A(net975),
    .X(_1782_));
 sg13g2_xnor2_1 _5030_ (.Y(_1783_),
    .A(_1780_),
    .B(_1782_));
 sg13g2_o21ai_1 _5031_ (.B1(net701),
    .Y(_1784_),
    .A1(net649),
    .A2(net975));
 sg13g2_a21oi_1 _5032_ (.A1(net649),
    .A2(_1783_),
    .Y(_0275_),
    .B1(_1784_));
 sg13g2_a21oi_1 _5033_ (.A1(_1780_),
    .A2(_1782_),
    .Y(_1785_),
    .B1(_1781_));
 sg13g2_nand2_1 _5034_ (.Y(_1786_),
    .A(\project_audio.genblk1[5].n_c_oh_my.phase[3] ),
    .B(\project_audio.freq[5][3] ));
 sg13g2_xnor2_1 _5035_ (.Y(_1787_),
    .A(net1019),
    .B(net729));
 sg13g2_xnor2_1 _5036_ (.Y(_1788_),
    .A(_1785_),
    .B(_1787_));
 sg13g2_o21ai_1 _5037_ (.B1(net701),
    .Y(_1789_),
    .A1(net649),
    .A2(net1019));
 sg13g2_a21oi_1 _5038_ (.A1(net649),
    .A2(_1788_),
    .Y(_0276_),
    .B1(_1789_));
 sg13g2_o21ai_1 _5039_ (.B1(_1786_),
    .Y(_1790_),
    .A1(_1785_),
    .A2(_1787_));
 sg13g2_and2_1 _5040_ (.A(\project_audio.genblk1[5].n_c_oh_my.phase[4] ),
    .B(\project_audio.freq[5][4] ),
    .X(_1791_));
 sg13g2_xor2_1 _5041_ (.B(net517),
    .A(net1027),
    .X(_1792_));
 sg13g2_xnor2_1 _5042_ (.Y(_1793_),
    .A(_1790_),
    .B(_1792_));
 sg13g2_o21ai_1 _5043_ (.B1(net701),
    .Y(_1794_),
    .A1(net649),
    .A2(net1027));
 sg13g2_a21oi_1 _5044_ (.A1(net649),
    .A2(_1793_),
    .Y(_0277_),
    .B1(_1794_));
 sg13g2_a21o_1 _5045_ (.A2(_1792_),
    .A1(_1790_),
    .B1(_1791_),
    .X(_1795_));
 sg13g2_or2_1 _5046_ (.X(_1796_),
    .B(\project_audio.freq[5][5] ),
    .A(\project_audio.genblk1[5].n_c_oh_my.phase[5] ));
 sg13g2_nand2_1 _5047_ (.Y(_1797_),
    .A(net880),
    .B(net469));
 sg13g2_nand2_1 _5048_ (.Y(_1798_),
    .A(_1796_),
    .B(_1797_));
 sg13g2_xor2_1 _5049_ (.B(_1798_),
    .A(_1795_),
    .X(_1799_));
 sg13g2_o21ai_1 _5050_ (.B1(net701),
    .Y(_1800_),
    .A1(net649),
    .A2(net880));
 sg13g2_a21oi_1 _5051_ (.A1(net648),
    .A2(_1799_),
    .Y(_0278_),
    .B1(_1800_));
 sg13g2_xnor2_1 _5052_ (.Y(_1801_),
    .A(\project_audio.genblk1[5].n_c_oh_my.phase[6] ),
    .B(\project_audio.freq[5][6] ));
 sg13g2_nand2_1 _5053_ (.Y(_1802_),
    .A(_1795_),
    .B(_1796_));
 sg13g2_a21oi_1 _5054_ (.A1(_1797_),
    .A2(_1802_),
    .Y(_1803_),
    .B1(_1801_));
 sg13g2_nand3_1 _5055_ (.B(_1801_),
    .C(_1802_),
    .A(_1797_),
    .Y(_1804_));
 sg13g2_nand2b_1 _5056_ (.Y(_1805_),
    .B(_1804_),
    .A_N(_1803_));
 sg13g2_o21ai_1 _5057_ (.B1(net703),
    .Y(_1806_),
    .A1(net648),
    .A2(net999));
 sg13g2_a21oi_1 _5058_ (.A1(net648),
    .A2(_1805_),
    .Y(_0279_),
    .B1(_1806_));
 sg13g2_a21oi_1 _5059_ (.A1(\project_audio.genblk1[5].n_c_oh_my.phase[6] ),
    .A2(\project_audio.freq[5][6] ),
    .Y(_1807_),
    .B1(_1803_));
 sg13g2_nand2_1 _5060_ (.Y(_1808_),
    .A(\project_audio.genblk1[5].n_c_oh_my.phase[7] ),
    .B(net744));
 sg13g2_xnor2_1 _5061_ (.Y(_1809_),
    .A(net1094),
    .B(net744));
 sg13g2_or2_1 _5062_ (.X(_1810_),
    .B(_1809_),
    .A(_1807_));
 sg13g2_xnor2_1 _5063_ (.Y(_1811_),
    .A(_1807_),
    .B(_1809_));
 sg13g2_o21ai_1 _5064_ (.B1(net703),
    .Y(_1812_),
    .A1(net648),
    .A2(net1094));
 sg13g2_a21oi_1 _5065_ (.A1(net648),
    .A2(_1811_),
    .Y(_0280_),
    .B1(_1812_));
 sg13g2_xnor2_1 _5066_ (.Y(_1813_),
    .A(\project_audio.genblk1[5].n_c_oh_my.phase[8] ),
    .B(\project_audio.freq[5][8] ));
 sg13g2_a21oi_1 _5067_ (.A1(_1808_),
    .A2(_1810_),
    .Y(_1814_),
    .B1(_1813_));
 sg13g2_nand3_1 _5068_ (.B(_1810_),
    .C(_1813_),
    .A(_1808_),
    .Y(_1815_));
 sg13g2_nand2b_1 _5069_ (.Y(_1816_),
    .B(_1815_),
    .A_N(_1814_));
 sg13g2_o21ai_1 _5070_ (.B1(net703),
    .Y(_1817_),
    .A1(net637),
    .A2(net955));
 sg13g2_a21oi_1 _5071_ (.A1(net637),
    .A2(_1816_),
    .Y(_0281_),
    .B1(_1817_));
 sg13g2_a21o_1 _5072_ (.A2(\project_audio.freq[5][8] ),
    .A1(net955),
    .B1(_1814_),
    .X(_1818_));
 sg13g2_nor2_1 _5073_ (.A(\project_audio.genblk1[5].n_c_oh_my.phase[9] ),
    .B(\project_audio.freq[5][9] ),
    .Y(_1819_));
 sg13g2_xor2_1 _5074_ (.B(net830),
    .A(net1157),
    .X(_1820_));
 sg13g2_xnor2_1 _5075_ (.Y(_1821_),
    .A(_1818_),
    .B(_1820_));
 sg13g2_o21ai_1 _5076_ (.B1(net703),
    .Y(_1822_),
    .A1(net637),
    .A2(net1157));
 sg13g2_a21oi_1 _5077_ (.A1(net637),
    .A2(_1821_),
    .Y(_0282_),
    .B1(_1822_));
 sg13g2_xnor2_1 _5078_ (.Y(_1823_),
    .A(net1038),
    .B(net798));
 sg13g2_a21oi_1 _5079_ (.A1(\project_audio.genblk1[5].n_c_oh_my.phase[9] ),
    .A2(\project_audio.freq[5][9] ),
    .Y(_1824_),
    .B1(_1818_));
 sg13g2_nor3_1 _5080_ (.A(_1819_),
    .B(_1823_),
    .C(_1824_),
    .Y(_1825_));
 sg13g2_o21ai_1 _5081_ (.B1(_1823_),
    .Y(_1826_),
    .A1(_1819_),
    .A2(_1824_));
 sg13g2_nand2b_1 _5082_ (.Y(_1827_),
    .B(_1826_),
    .A_N(_1825_));
 sg13g2_o21ai_1 _5083_ (.B1(net703),
    .Y(_1828_),
    .A1(net635),
    .A2(net1038));
 sg13g2_a21oi_1 _5084_ (.A1(net635),
    .A2(_1827_),
    .Y(_0283_),
    .B1(_1828_));
 sg13g2_a21oi_1 _5085_ (.A1(net1038),
    .A2(net798),
    .Y(_1829_),
    .B1(_1825_));
 sg13g2_nor2_1 _5086_ (.A(\project_audio.genblk1[5].n_c_oh_my.phase[11] ),
    .B(\project_audio.freq[5][11] ),
    .Y(_1830_));
 sg13g2_nand2_1 _5087_ (.Y(_1831_),
    .A(net1063),
    .B(\project_audio.freq[5][11] ));
 sg13g2_nand2b_1 _5088_ (.Y(_1832_),
    .B(_1831_),
    .A_N(_1830_));
 sg13g2_xnor2_1 _5089_ (.Y(_1833_),
    .A(_1829_),
    .B(_1832_));
 sg13g2_o21ai_1 _5090_ (.B1(net703),
    .Y(_1834_),
    .A1(net634),
    .A2(net1063));
 sg13g2_a21oi_1 _5091_ (.A1(net634),
    .A2(_1833_),
    .Y(_0284_),
    .B1(_1834_));
 sg13g2_o21ai_1 _5092_ (.B1(_1831_),
    .Y(_1835_),
    .A1(_1829_),
    .A2(_1830_));
 sg13g2_a21oi_1 _5093_ (.A1(net634),
    .A2(_1835_),
    .Y(_1836_),
    .B1(net508));
 sg13g2_nand3_1 _5094_ (.B(net508),
    .C(_1835_),
    .A(net634),
    .Y(_1837_));
 sg13g2_inv_1 _5095_ (.Y(_1838_),
    .A(_1837_));
 sg13g2_nor3_1 _5096_ (.A(net682),
    .B(_1836_),
    .C(_1838_),
    .Y(_0285_));
 sg13g2_nand2_1 _5097_ (.Y(_1839_),
    .A(net510),
    .B(_1838_));
 sg13g2_nand2_1 _5098_ (.Y(_1840_),
    .A(net688),
    .B(_1839_));
 sg13g2_a21oi_1 _5099_ (.A1(_2486_),
    .A2(_1837_),
    .Y(_0286_),
    .B1(_1840_));
 sg13g2_o21ai_1 _5100_ (.B1(net688),
    .Y(_1841_),
    .A1(_2485_),
    .A2(_1839_));
 sg13g2_a21oi_1 _5101_ (.A1(_2485_),
    .A2(_1839_),
    .Y(_0287_),
    .B1(_1841_));
 sg13g2_and4_1 _5102_ (.A(\project_audio.genblk1[5].n_c_oh_my.phase[14] ),
    .B(\project_audio.genblk1[5].n_c_oh_my.phase[13] ),
    .C(\project_audio.genblk1[5].n_c_oh_my.phase[12] ),
    .D(net688),
    .X(_1842_));
 sg13g2_nand3_1 _5103_ (.B(_1835_),
    .C(_1842_),
    .A(_1771_),
    .Y(_1843_));
 sg13g2_o21ai_1 _5104_ (.B1(_1843_),
    .Y(_0288_),
    .A1(_2484_),
    .A2(_1841_));
 sg13g2_nor2b_1 _5105_ (.A(net492),
    .B_N(net638),
    .Y(_1844_));
 sg13g2_o21ai_1 _5106_ (.B1(net694),
    .Y(_1845_),
    .A1(net638),
    .A2(net967));
 sg13g2_nor2_1 _5107_ (.A(_1844_),
    .B(_1845_),
    .Y(_0289_));
 sg13g2_nand2_1 _5108_ (.Y(_1846_),
    .A(net650),
    .B(net482));
 sg13g2_nand2_1 _5109_ (.Y(_1847_),
    .A(net892),
    .B(net482));
 sg13g2_xor2_1 _5110_ (.B(_1846_),
    .A(net892),
    .X(_1848_));
 sg13g2_nor2_1 _5111_ (.A(net684),
    .B(_1848_),
    .Y(_0290_));
 sg13g2_nand2_1 _5112_ (.Y(_1849_),
    .A(\project_audio.genblk1[4].n_c_oh_my.phase[1] ),
    .B(\project_audio.freq[4][1] ));
 sg13g2_xnor2_1 _5113_ (.Y(_1850_),
    .A(net1117),
    .B(net764));
 sg13g2_xnor2_1 _5114_ (.Y(_1851_),
    .A(_1847_),
    .B(_1850_));
 sg13g2_o21ai_1 _5115_ (.B1(net710),
    .Y(_1852_),
    .A1(net651),
    .A2(net1117));
 sg13g2_a21oi_1 _5116_ (.A1(net651),
    .A2(_1851_),
    .Y(_0291_),
    .B1(_1852_));
 sg13g2_o21ai_1 _5117_ (.B1(_1849_),
    .Y(_1853_),
    .A1(_1847_),
    .A2(_1850_));
 sg13g2_and2_1 _5118_ (.A(\project_audio.genblk1[4].n_c_oh_my.phase[2] ),
    .B(\project_audio.freq[4][2] ),
    .X(_1854_));
 sg13g2_xor2_1 _5119_ (.B(net518),
    .A(net987),
    .X(_1855_));
 sg13g2_xnor2_1 _5120_ (.Y(_1856_),
    .A(_1853_),
    .B(_1855_));
 sg13g2_o21ai_1 _5121_ (.B1(net710),
    .Y(_1857_),
    .A1(net650),
    .A2(net987));
 sg13g2_a21oi_1 _5122_ (.A1(net650),
    .A2(_1856_),
    .Y(_0292_),
    .B1(_1857_));
 sg13g2_a21oi_1 _5123_ (.A1(_1853_),
    .A2(_1855_),
    .Y(_1858_),
    .B1(_1854_));
 sg13g2_nand2_1 _5124_ (.Y(_1859_),
    .A(net1005),
    .B(\project_audio.freq[4][3] ));
 sg13g2_xnor2_1 _5125_ (.Y(_1860_),
    .A(net1005),
    .B(net796));
 sg13g2_xnor2_1 _5126_ (.Y(_1861_),
    .A(_1858_),
    .B(_1860_));
 sg13g2_o21ai_1 _5127_ (.B1(net705),
    .Y(_1862_),
    .A1(net650),
    .A2(net1005));
 sg13g2_a21oi_1 _5128_ (.A1(net650),
    .A2(_1861_),
    .Y(_0293_),
    .B1(_1862_));
 sg13g2_o21ai_1 _5129_ (.B1(_1859_),
    .Y(_1863_),
    .A1(_1858_),
    .A2(_1860_));
 sg13g2_and2_1 _5130_ (.A(\project_audio.genblk1[4].n_c_oh_my.phase[4] ),
    .B(\project_audio.freq[4][4] ),
    .X(_1864_));
 sg13g2_xor2_1 _5131_ (.B(net520),
    .A(net1034),
    .X(_1865_));
 sg13g2_xnor2_1 _5132_ (.Y(_1866_),
    .A(_1863_),
    .B(_1865_));
 sg13g2_o21ai_1 _5133_ (.B1(net705),
    .Y(_1867_),
    .A1(net650),
    .A2(net1034));
 sg13g2_a21oi_1 _5134_ (.A1(net650),
    .A2(_1866_),
    .Y(_0294_),
    .B1(_1867_));
 sg13g2_a21o_1 _5135_ (.A2(_1865_),
    .A1(_1863_),
    .B1(_1864_),
    .X(_1868_));
 sg13g2_or2_1 _5136_ (.X(_1869_),
    .B(\project_audio.freq[4][5] ),
    .A(\project_audio.genblk1[4].n_c_oh_my.phase[5] ));
 sg13g2_nand2_1 _5137_ (.Y(_1870_),
    .A(net903),
    .B(net467));
 sg13g2_nand2_1 _5138_ (.Y(_1871_),
    .A(_1869_),
    .B(_1870_));
 sg13g2_xor2_1 _5139_ (.B(_1871_),
    .A(_1868_),
    .X(_1872_));
 sg13g2_o21ai_1 _5140_ (.B1(net705),
    .Y(_1873_),
    .A1(net636),
    .A2(net903));
 sg13g2_a21oi_1 _5141_ (.A1(net636),
    .A2(_1872_),
    .Y(_0295_),
    .B1(_1873_));
 sg13g2_xnor2_1 _5142_ (.Y(_1874_),
    .A(\project_audio.genblk1[4].n_c_oh_my.phase[6] ),
    .B(\project_audio.freq[4][6] ));
 sg13g2_nand2_1 _5143_ (.Y(_1875_),
    .A(_1868_),
    .B(_1869_));
 sg13g2_a21oi_1 _5144_ (.A1(_1870_),
    .A2(_1875_),
    .Y(_1876_),
    .B1(_1874_));
 sg13g2_nand3_1 _5145_ (.B(_1874_),
    .C(_1875_),
    .A(_1870_),
    .Y(_1877_));
 sg13g2_nand2b_1 _5146_ (.Y(_1878_),
    .B(_1877_),
    .A_N(_1876_));
 sg13g2_o21ai_1 _5147_ (.B1(net704),
    .Y(_1879_),
    .A1(net636),
    .A2(net968));
 sg13g2_a21oi_1 _5148_ (.A1(net636),
    .A2(_1878_),
    .Y(_0296_),
    .B1(_1879_));
 sg13g2_a21oi_1 _5149_ (.A1(net968),
    .A2(net733),
    .Y(_1880_),
    .B1(_1876_));
 sg13g2_nand2_1 _5150_ (.Y(_1881_),
    .A(\project_audio.genblk1[4].n_c_oh_my.phase[7] ),
    .B(net802));
 sg13g2_xnor2_1 _5151_ (.Y(_1882_),
    .A(net1042),
    .B(net802));
 sg13g2_or2_1 _5152_ (.X(_1883_),
    .B(_1882_),
    .A(_1880_));
 sg13g2_xnor2_1 _5153_ (.Y(_1884_),
    .A(_1880_),
    .B(_1882_));
 sg13g2_o21ai_1 _5154_ (.B1(net704),
    .Y(_1885_),
    .A1(net635),
    .A2(net1042));
 sg13g2_a21oi_1 _5155_ (.A1(net635),
    .A2(_1884_),
    .Y(_0297_),
    .B1(_1885_));
 sg13g2_xnor2_1 _5156_ (.Y(_1886_),
    .A(\project_audio.genblk1[4].n_c_oh_my.phase[8] ),
    .B(\project_audio.freq[4][8] ));
 sg13g2_a21oi_1 _5157_ (.A1(_1881_),
    .A2(_1883_),
    .Y(_1887_),
    .B1(_1886_));
 sg13g2_nand3_1 _5158_ (.B(_1883_),
    .C(_1886_),
    .A(_1881_),
    .Y(_1888_));
 sg13g2_nand2b_1 _5159_ (.Y(_1889_),
    .B(_1888_),
    .A_N(_1887_));
 sg13g2_o21ai_1 _5160_ (.B1(net704),
    .Y(_1890_),
    .A1(net635),
    .A2(net995));
 sg13g2_a21oi_1 _5161_ (.A1(net635),
    .A2(_1889_),
    .Y(_0298_),
    .B1(_1890_));
 sg13g2_a21o_1 _5162_ (.A2(\project_audio.freq[4][8] ),
    .A1(\project_audio.genblk1[4].n_c_oh_my.phase[8] ),
    .B1(_1887_),
    .X(_1891_));
 sg13g2_nor2_1 _5163_ (.A(\project_audio.genblk1[4].n_c_oh_my.phase[9] ),
    .B(\project_audio.freq[4][9] ),
    .Y(_1892_));
 sg13g2_xor2_1 _5164_ (.B(net823),
    .A(net1160),
    .X(_1893_));
 sg13g2_xnor2_1 _5165_ (.Y(_1894_),
    .A(_1891_),
    .B(_1893_));
 sg13g2_o21ai_1 _5166_ (.B1(net695),
    .Y(_1895_),
    .A1(net633),
    .A2(net1160));
 sg13g2_a21oi_1 _5167_ (.A1(net633),
    .A2(_1894_),
    .Y(_0299_),
    .B1(_1895_));
 sg13g2_xnor2_1 _5168_ (.Y(_1896_),
    .A(net1084),
    .B(net818));
 sg13g2_a21oi_1 _5169_ (.A1(\project_audio.genblk1[4].n_c_oh_my.phase[9] ),
    .A2(\project_audio.freq[4][9] ),
    .Y(_1897_),
    .B1(_1891_));
 sg13g2_nor3_1 _5170_ (.A(_1892_),
    .B(_1896_),
    .C(_1897_),
    .Y(_1898_));
 sg13g2_o21ai_1 _5171_ (.B1(_1896_),
    .Y(_1899_),
    .A1(_1892_),
    .A2(_1897_));
 sg13g2_nand2b_1 _5172_ (.Y(_1900_),
    .B(_1899_),
    .A_N(_1898_));
 sg13g2_o21ai_1 _5173_ (.B1(net695),
    .Y(_1901_),
    .A1(net633),
    .A2(net1084));
 sg13g2_a21oi_1 _5174_ (.A1(net633),
    .A2(_1900_),
    .Y(_0300_),
    .B1(_1901_));
 sg13g2_a21oi_1 _5175_ (.A1(\project_audio.genblk1[4].n_c_oh_my.phase[10] ),
    .A2(net818),
    .Y(_1902_),
    .B1(_1898_));
 sg13g2_nor2_1 _5176_ (.A(\project_audio.genblk1[4].n_c_oh_my.phase[11] ),
    .B(\project_audio.freq[4][11] ),
    .Y(_1903_));
 sg13g2_nand2_1 _5177_ (.Y(_1904_),
    .A(net939),
    .B(net448));
 sg13g2_nand2b_1 _5178_ (.Y(_1905_),
    .B(_1904_),
    .A_N(_1903_));
 sg13g2_xnor2_1 _5179_ (.Y(_1906_),
    .A(_1902_),
    .B(_1905_));
 sg13g2_o21ai_1 _5180_ (.B1(net695),
    .Y(_1907_),
    .A1(net632),
    .A2(net939));
 sg13g2_a21oi_1 _5181_ (.A1(net632),
    .A2(_1906_),
    .Y(_0301_),
    .B1(_1907_));
 sg13g2_o21ai_1 _5182_ (.B1(_1904_),
    .Y(_1908_),
    .A1(_1902_),
    .A2(_1903_));
 sg13g2_a21oi_1 _5183_ (.A1(net632),
    .A2(_1908_),
    .Y(_1909_),
    .B1(net537));
 sg13g2_nand3_1 _5184_ (.B(net537),
    .C(_1908_),
    .A(net632),
    .Y(_1910_));
 sg13g2_inv_1 _5185_ (.Y(_1911_),
    .A(_1910_));
 sg13g2_nor3_1 _5186_ (.A(net680),
    .B(_1909_),
    .C(_1911_),
    .Y(_0302_));
 sg13g2_nand2_1 _5187_ (.Y(_1912_),
    .A(net487),
    .B(_1911_));
 sg13g2_nand2_1 _5188_ (.Y(_1913_),
    .A(net694),
    .B(_1912_));
 sg13g2_a21oi_1 _5189_ (.A1(_2483_),
    .A2(_1910_),
    .Y(_0303_),
    .B1(_1913_));
 sg13g2_o21ai_1 _5190_ (.B1(net694),
    .Y(_1914_),
    .A1(_2482_),
    .A2(_1912_));
 sg13g2_a21oi_1 _5191_ (.A1(_2482_),
    .A2(_1912_),
    .Y(_0304_),
    .B1(_1914_));
 sg13g2_and4_1 _5192_ (.A(\project_audio.genblk1[4].n_c_oh_my.phase[14] ),
    .B(net487),
    .C(\project_audio.genblk1[4].n_c_oh_my.phase[12] ),
    .D(net694),
    .X(_1915_));
 sg13g2_nand3_1 _5193_ (.B(_1908_),
    .C(_1915_),
    .A(_1844_),
    .Y(_1916_));
 sg13g2_o21ai_1 _5194_ (.B1(_1916_),
    .Y(_0305_),
    .A1(_2481_),
    .A2(_1914_));
 sg13g2_nor2b_1 _5195_ (.A(net525),
    .B_N(net639),
    .Y(_1917_));
 sg13g2_o21ai_1 _5196_ (.B1(net697),
    .Y(_1918_),
    .A1(net638),
    .A2(net1029));
 sg13g2_nor2_1 _5197_ (.A(_1917_),
    .B(_1918_),
    .Y(_0306_));
 sg13g2_nand2_1 _5198_ (.Y(_1919_),
    .A(net658),
    .B(net470));
 sg13g2_nand2_1 _5199_ (.Y(_1920_),
    .A(net909),
    .B(net470));
 sg13g2_xor2_1 _5200_ (.B(_1919_),
    .A(net909),
    .X(_1921_));
 sg13g2_nor2_1 _5201_ (.A(net684),
    .B(_1921_),
    .Y(_0307_));
 sg13g2_nand2_1 _5202_ (.Y(_1922_),
    .A(\project_audio.genblk1[3].n_c_oh_my.phase[1] ),
    .B(\project_audio.freq[3][1] ));
 sg13g2_xnor2_1 _5203_ (.Y(_1923_),
    .A(net977),
    .B(net501));
 sg13g2_xnor2_1 _5204_ (.Y(_1924_),
    .A(_1920_),
    .B(_1923_));
 sg13g2_o21ai_1 _5205_ (.B1(net705),
    .Y(_1925_),
    .A1(net658),
    .A2(net977));
 sg13g2_a21oi_1 _5206_ (.A1(net658),
    .A2(_1924_),
    .Y(_0308_),
    .B1(_1925_));
 sg13g2_o21ai_1 _5207_ (.B1(_1922_),
    .Y(_1926_),
    .A1(_1920_),
    .A2(_1923_));
 sg13g2_and2_1 _5208_ (.A(\project_audio.genblk1[3].n_c_oh_my.phase[2] ),
    .B(\project_audio.freq[3][2] ),
    .X(_1927_));
 sg13g2_xor2_1 _5209_ (.B(net725),
    .A(net1031),
    .X(_1928_));
 sg13g2_xnor2_1 _5210_ (.Y(_1929_),
    .A(_1926_),
    .B(_1928_));
 sg13g2_o21ai_1 _5211_ (.B1(net705),
    .Y(_1930_),
    .A1(net636),
    .A2(net1031));
 sg13g2_a21oi_1 _5212_ (.A1(net636),
    .A2(_1929_),
    .Y(_0309_),
    .B1(_1930_));
 sg13g2_a21oi_2 _5213_ (.B1(_1927_),
    .Y(_1931_),
    .A2(_1928_),
    .A1(_1926_));
 sg13g2_nand2_1 _5214_ (.Y(_1932_),
    .A(\project_audio.genblk1[3].n_c_oh_my.phase[3] ),
    .B(\project_audio.freq[3][3] ));
 sg13g2_xnor2_1 _5215_ (.Y(_1933_),
    .A(net1033),
    .B(net831));
 sg13g2_xnor2_1 _5216_ (.Y(_1934_),
    .A(_1931_),
    .B(_1933_));
 sg13g2_o21ai_1 _5217_ (.B1(net704),
    .Y(_1935_),
    .A1(net635),
    .A2(net1033));
 sg13g2_a21oi_1 _5218_ (.A1(net635),
    .A2(_1934_),
    .Y(_0310_),
    .B1(_1935_));
 sg13g2_o21ai_1 _5219_ (.B1(_1932_),
    .Y(_1936_),
    .A1(_1931_),
    .A2(_1933_));
 sg13g2_and2_1 _5220_ (.A(\project_audio.genblk1[3].n_c_oh_my.phase[4] ),
    .B(\project_audio.freq[3][4] ),
    .X(_1937_));
 sg13g2_xor2_1 _5221_ (.B(net799),
    .A(net1043),
    .X(_1938_));
 sg13g2_xnor2_1 _5222_ (.Y(_1939_),
    .A(_1936_),
    .B(_1938_));
 sg13g2_o21ai_1 _5223_ (.B1(net704),
    .Y(_1940_),
    .A1(net643),
    .A2(net1043));
 sg13g2_a21oi_1 _5224_ (.A1(net643),
    .A2(_1939_),
    .Y(_0311_),
    .B1(_1940_));
 sg13g2_a21o_1 _5225_ (.A2(_1938_),
    .A1(_1936_),
    .B1(_1937_),
    .X(_1941_));
 sg13g2_or2_1 _5226_ (.X(_1942_),
    .B(\project_audio.freq[3][5] ),
    .A(\project_audio.genblk1[3].n_c_oh_my.phase[5] ));
 sg13g2_nand2_1 _5227_ (.Y(_1943_),
    .A(net938),
    .B(net491));
 sg13g2_nand2_1 _5228_ (.Y(_1944_),
    .A(_1942_),
    .B(_1943_));
 sg13g2_xor2_1 _5229_ (.B(_1944_),
    .A(_1941_),
    .X(_1945_));
 sg13g2_o21ai_1 _5230_ (.B1(net704),
    .Y(_1946_),
    .A1(net643),
    .A2(net938));
 sg13g2_a21oi_1 _5231_ (.A1(net643),
    .A2(_1945_),
    .Y(_0312_),
    .B1(_1946_));
 sg13g2_xnor2_1 _5232_ (.Y(_1947_),
    .A(\project_audio.genblk1[3].n_c_oh_my.phase[6] ),
    .B(\project_audio.freq[3][6] ));
 sg13g2_nand2_1 _5233_ (.Y(_1948_),
    .A(_1941_),
    .B(_1942_));
 sg13g2_a21oi_1 _5234_ (.A1(_1943_),
    .A2(_1948_),
    .Y(_1949_),
    .B1(_1947_));
 sg13g2_nand3_1 _5235_ (.B(_1947_),
    .C(_1948_),
    .A(_1943_),
    .Y(_1950_));
 sg13g2_nand2b_1 _5236_ (.Y(_1951_),
    .B(_1950_),
    .A_N(_1949_));
 sg13g2_o21ai_1 _5237_ (.B1(net704),
    .Y(_1952_),
    .A1(net643),
    .A2(net1025));
 sg13g2_a21oi_1 _5238_ (.A1(net643),
    .A2(_1951_),
    .Y(_0313_),
    .B1(_1952_));
 sg13g2_a21oi_1 _5239_ (.A1(net1025),
    .A2(net844),
    .Y(_1953_),
    .B1(_1949_));
 sg13g2_nand2_1 _5240_ (.Y(_1954_),
    .A(\project_audio.genblk1[3].n_c_oh_my.phase[7] ),
    .B(net765));
 sg13g2_xnor2_1 _5241_ (.Y(_1955_),
    .A(net1065),
    .B(net765));
 sg13g2_or2_1 _5242_ (.X(_1956_),
    .B(_1955_),
    .A(_1953_));
 sg13g2_xnor2_1 _5243_ (.Y(_1957_),
    .A(_1953_),
    .B(_1955_));
 sg13g2_o21ai_1 _5244_ (.B1(net704),
    .Y(_1958_),
    .A1(net644),
    .A2(net1065));
 sg13g2_a21oi_1 _5245_ (.A1(net644),
    .A2(_1957_),
    .Y(_0314_),
    .B1(_1958_));
 sg13g2_xnor2_1 _5246_ (.Y(_1959_),
    .A(\project_audio.genblk1[3].n_c_oh_my.phase[8] ),
    .B(\project_audio.freq[3][8] ));
 sg13g2_a21oi_1 _5247_ (.A1(_1954_),
    .A2(_1956_),
    .Y(_1960_),
    .B1(_1959_));
 sg13g2_nand3_1 _5248_ (.B(_1956_),
    .C(_1959_),
    .A(_1954_),
    .Y(_1961_));
 sg13g2_nand2b_1 _5249_ (.Y(_1962_),
    .B(_1961_),
    .A_N(_1960_));
 sg13g2_o21ai_1 _5250_ (.B1(net695),
    .Y(_1963_),
    .A1(net639),
    .A2(net1015));
 sg13g2_a21oi_1 _5251_ (.A1(net639),
    .A2(_1962_),
    .Y(_0315_),
    .B1(_1963_));
 sg13g2_a21o_1 _5252_ (.A2(\project_audio.freq[3][8] ),
    .A1(\project_audio.genblk1[3].n_c_oh_my.phase[8] ),
    .B1(_1960_),
    .X(_1964_));
 sg13g2_nor2_1 _5253_ (.A(\project_audio.genblk1[3].n_c_oh_my.phase[9] ),
    .B(\project_audio.freq[3][9] ),
    .Y(_1965_));
 sg13g2_xor2_1 _5254_ (.B(net843),
    .A(net1165),
    .X(_1966_));
 sg13g2_xnor2_1 _5255_ (.Y(_1967_),
    .A(_1964_),
    .B(_1966_));
 sg13g2_o21ai_1 _5256_ (.B1(net700),
    .Y(_1968_),
    .A1(net642),
    .A2(net1165));
 sg13g2_a21oi_1 _5257_ (.A1(net639),
    .A2(_1967_),
    .Y(_0316_),
    .B1(_1968_));
 sg13g2_xnor2_1 _5258_ (.Y(_1969_),
    .A(\project_audio.genblk1[3].n_c_oh_my.phase[10] ),
    .B(\project_audio.freq[3][10] ));
 sg13g2_a21oi_1 _5259_ (.A1(\project_audio.genblk1[3].n_c_oh_my.phase[9] ),
    .A2(\project_audio.freq[3][9] ),
    .Y(_1970_),
    .B1(_1964_));
 sg13g2_nor3_1 _5260_ (.A(_1965_),
    .B(_1969_),
    .C(_1970_),
    .Y(_1971_));
 sg13g2_o21ai_1 _5261_ (.B1(_1969_),
    .Y(_1972_),
    .A1(_1965_),
    .A2(_1970_));
 sg13g2_nand2b_1 _5262_ (.Y(_1973_),
    .B(_1972_),
    .A_N(_1971_));
 sg13g2_o21ai_1 _5263_ (.B1(net695),
    .Y(_1974_),
    .A1(net639),
    .A2(net1008));
 sg13g2_a21oi_1 _5264_ (.A1(net639),
    .A2(_1973_),
    .Y(_0317_),
    .B1(_1974_));
 sg13g2_a21oi_1 _5265_ (.A1(\project_audio.genblk1[3].n_c_oh_my.phase[10] ),
    .A2(net724),
    .Y(_1975_),
    .B1(_1971_));
 sg13g2_nor2_1 _5266_ (.A(\project_audio.genblk1[3].n_c_oh_my.phase[11] ),
    .B(\project_audio.freq[3][11] ),
    .Y(_1976_));
 sg13g2_nand2_1 _5267_ (.Y(_1977_),
    .A(net946),
    .B(net454));
 sg13g2_nand2b_1 _5268_ (.Y(_1978_),
    .B(_1977_),
    .A_N(_1976_));
 sg13g2_xnor2_1 _5269_ (.Y(_1979_),
    .A(_1975_),
    .B(_1978_));
 sg13g2_o21ai_1 _5270_ (.B1(net700),
    .Y(_1980_),
    .A1(net638),
    .A2(net946));
 sg13g2_a21oi_1 _5271_ (.A1(net638),
    .A2(_1979_),
    .Y(_0318_),
    .B1(_1980_));
 sg13g2_o21ai_1 _5272_ (.B1(_1977_),
    .Y(_1981_),
    .A1(_1975_),
    .A2(_1976_));
 sg13g2_a21oi_1 _5273_ (.A1(net638),
    .A2(_1981_),
    .Y(_1982_),
    .B1(net513));
 sg13g2_nand3_1 _5274_ (.B(net513),
    .C(_1981_),
    .A(net638),
    .Y(_1983_));
 sg13g2_inv_1 _5275_ (.Y(_1984_),
    .A(_1983_));
 sg13g2_nor3_1 _5276_ (.A(net681),
    .B(_1982_),
    .C(_1984_),
    .Y(_0319_));
 sg13g2_nand2_1 _5277_ (.Y(_1985_),
    .A(net480),
    .B(_1984_));
 sg13g2_nand2_1 _5278_ (.Y(_1986_),
    .A(net695),
    .B(_1985_));
 sg13g2_a21oi_1 _5279_ (.A1(_2480_),
    .A2(_1983_),
    .Y(_0320_),
    .B1(_1986_));
 sg13g2_o21ai_1 _5280_ (.B1(net696),
    .Y(_1987_),
    .A1(_2479_),
    .A2(_1985_));
 sg13g2_a21oi_1 _5281_ (.A1(_2479_),
    .A2(_1985_),
    .Y(_0321_),
    .B1(_1987_));
 sg13g2_and4_1 _5282_ (.A(\project_audio.genblk1[3].n_c_oh_my.phase[14] ),
    .B(net480),
    .C(net513),
    .D(net695),
    .X(_1988_));
 sg13g2_nand3_1 _5283_ (.B(_1981_),
    .C(_1988_),
    .A(_1917_),
    .Y(_1989_));
 sg13g2_o21ai_1 _5284_ (.B1(_1989_),
    .Y(_0322_),
    .A1(_2478_),
    .A2(_1987_));
 sg13g2_nor2b_1 _5285_ (.A(net511),
    .B_N(net641),
    .Y(_1990_));
 sg13g2_o21ai_1 _5286_ (.B1(net696),
    .Y(_1991_),
    .A1(net641),
    .A2(net980));
 sg13g2_nor2_1 _5287_ (.A(_1990_),
    .B(_1991_),
    .Y(_0323_));
 sg13g2_nand2_1 _5288_ (.Y(_1992_),
    .A(net658),
    .B(net472));
 sg13g2_nand2_1 _5289_ (.Y(_1993_),
    .A(net883),
    .B(net472));
 sg13g2_xor2_1 _5290_ (.B(_1992_),
    .A(net883),
    .X(_1994_));
 sg13g2_nor2_1 _5291_ (.A(net683),
    .B(_1994_),
    .Y(_0324_));
 sg13g2_nand2_1 _5292_ (.Y(_1995_),
    .A(\project_audio.genblk1[2].n_c_oh_my.phase[1] ),
    .B(\project_audio.freq[2][1] ));
 sg13g2_xnor2_1 _5293_ (.Y(_1996_),
    .A(net1024),
    .B(net515));
 sg13g2_xnor2_1 _5294_ (.Y(_1997_),
    .A(_1993_),
    .B(_1996_));
 sg13g2_o21ai_1 _5295_ (.B1(net707),
    .Y(_1998_),
    .A1(net644),
    .A2(net1024));
 sg13g2_a21oi_1 _5296_ (.A1(net644),
    .A2(_1997_),
    .Y(_0325_),
    .B1(_1998_));
 sg13g2_o21ai_1 _5297_ (.B1(_1995_),
    .Y(_1999_),
    .A1(_1993_),
    .A2(_1996_));
 sg13g2_and2_1 _5298_ (.A(net1243),
    .B(\project_audio.freq[2][2] ),
    .X(_2000_));
 sg13g2_xor2_1 _5299_ (.B(net746),
    .A(net1100),
    .X(_2001_));
 sg13g2_xnor2_1 _5300_ (.Y(_2002_),
    .A(_1999_),
    .B(_2001_));
 sg13g2_o21ai_1 _5301_ (.B1(net706),
    .Y(_2003_),
    .A1(net644),
    .A2(net1100));
 sg13g2_a21oi_1 _5302_ (.A1(net644),
    .A2(_2002_),
    .Y(_0326_),
    .B1(_2003_));
 sg13g2_a21oi_1 _5303_ (.A1(_1999_),
    .A2(_2001_),
    .Y(_2004_),
    .B1(_2000_));
 sg13g2_nand2_1 _5304_ (.Y(_2005_),
    .A(\project_audio.genblk1[2].n_c_oh_my.phase[3] ),
    .B(\project_audio.freq[2][3] ));
 sg13g2_xnor2_1 _5305_ (.Y(_2006_),
    .A(net1079),
    .B(net789));
 sg13g2_xnor2_1 _5306_ (.Y(_2007_),
    .A(_2004_),
    .B(_2006_));
 sg13g2_o21ai_1 _5307_ (.B1(net706),
    .Y(_2008_),
    .A1(net643),
    .A2(net1079));
 sg13g2_a21oi_1 _5308_ (.A1(net643),
    .A2(_2007_),
    .Y(_0327_),
    .B1(_2008_));
 sg13g2_o21ai_1 _5309_ (.B1(_2005_),
    .Y(_2009_),
    .A1(_2004_),
    .A2(_2006_));
 sg13g2_and2_1 _5310_ (.A(\project_audio.genblk1[2].n_c_oh_my.phase[4] ),
    .B(\project_audio.freq[2][4] ),
    .X(_2010_));
 sg13g2_xor2_1 _5311_ (.B(net742),
    .A(net1003),
    .X(_2011_));
 sg13g2_xnor2_1 _5312_ (.Y(_2012_),
    .A(_2009_),
    .B(_2011_));
 sg13g2_o21ai_1 _5313_ (.B1(net706),
    .Y(_2013_),
    .A1(net646),
    .A2(net1003));
 sg13g2_a21oi_1 _5314_ (.A1(net646),
    .A2(_2012_),
    .Y(_0328_),
    .B1(_2013_));
 sg13g2_a21o_1 _5315_ (.A2(_2011_),
    .A1(_2009_),
    .B1(_2010_),
    .X(_2014_));
 sg13g2_or2_1 _5316_ (.X(_2015_),
    .B(\project_audio.freq[2][5] ),
    .A(\project_audio.genblk1[2].n_c_oh_my.phase[5] ));
 sg13g2_nand2_1 _5317_ (.Y(_2016_),
    .A(net1007),
    .B(net532));
 sg13g2_nand2_1 _5318_ (.Y(_2017_),
    .A(_2015_),
    .B(_2016_));
 sg13g2_xor2_1 _5319_ (.B(_2017_),
    .A(_2014_),
    .X(_2018_));
 sg13g2_o21ai_1 _5320_ (.B1(net706),
    .Y(_2019_),
    .A1(net646),
    .A2(net1007));
 sg13g2_a21oi_1 _5321_ (.A1(net646),
    .A2(_2018_),
    .Y(_0329_),
    .B1(_2019_));
 sg13g2_xnor2_1 _5322_ (.Y(_2020_),
    .A(\project_audio.genblk1[2].n_c_oh_my.phase[6] ),
    .B(\project_audio.freq[2][6] ));
 sg13g2_nand2_1 _5323_ (.Y(_2021_),
    .A(_2014_),
    .B(_2015_));
 sg13g2_a21oi_1 _5324_ (.A1(_2016_),
    .A2(_2021_),
    .Y(_2022_),
    .B1(_2020_));
 sg13g2_nand3_1 _5325_ (.B(_2020_),
    .C(_2021_),
    .A(_2016_),
    .Y(_2023_));
 sg13g2_nand2b_1 _5326_ (.Y(_2024_),
    .B(_2023_),
    .A_N(_2022_));
 sg13g2_o21ai_1 _5327_ (.B1(net706),
    .Y(_2025_),
    .A1(net646),
    .A2(net1110));
 sg13g2_a21oi_1 _5328_ (.A1(net646),
    .A2(_2024_),
    .Y(_0330_),
    .B1(_2025_));
 sg13g2_a21oi_1 _5329_ (.A1(net1110),
    .A2(net732),
    .Y(_2026_),
    .B1(_2022_));
 sg13g2_nand2_1 _5330_ (.Y(_2027_),
    .A(\project_audio.genblk1[2].n_c_oh_my.phase[7] ),
    .B(net773));
 sg13g2_xnor2_1 _5331_ (.Y(_2028_),
    .A(net1118),
    .B(net773));
 sg13g2_or2_1 _5332_ (.X(_2029_),
    .B(_2028_),
    .A(_2026_));
 sg13g2_xnor2_1 _5333_ (.Y(_2030_),
    .A(_2026_),
    .B(_2028_));
 sg13g2_o21ai_1 _5334_ (.B1(net706),
    .Y(_2031_),
    .A1(net645),
    .A2(net1118));
 sg13g2_a21oi_1 _5335_ (.A1(net645),
    .A2(_2030_),
    .Y(_0331_),
    .B1(_2031_));
 sg13g2_xnor2_1 _5336_ (.Y(_2032_),
    .A(\project_audio.genblk1[2].n_c_oh_my.phase[8] ),
    .B(\project_audio.freq[2][8] ));
 sg13g2_a21oi_1 _5337_ (.A1(_2027_),
    .A2(_2029_),
    .Y(_2033_),
    .B1(_2032_));
 sg13g2_nand3_1 _5338_ (.B(_2029_),
    .C(_2032_),
    .A(_2027_),
    .Y(_2034_));
 sg13g2_nand2b_1 _5339_ (.Y(_2035_),
    .B(_2034_),
    .A_N(_2033_));
 sg13g2_o21ai_1 _5340_ (.B1(net706),
    .Y(_2036_),
    .A1(net645),
    .A2(net997));
 sg13g2_a21oi_1 _5341_ (.A1(net645),
    .A2(_2035_),
    .Y(_0332_),
    .B1(_2036_));
 sg13g2_a21o_1 _5342_ (.A2(\project_audio.freq[2][8] ),
    .A1(\project_audio.genblk1[2].n_c_oh_my.phase[8] ),
    .B1(_2033_),
    .X(_2037_));
 sg13g2_nor2_1 _5343_ (.A(\project_audio.genblk1[2].n_c_oh_my.phase[9] ),
    .B(net824),
    .Y(_2038_));
 sg13g2_xor2_1 _5344_ (.B(net824),
    .A(net1153),
    .X(_2039_));
 sg13g2_xnor2_1 _5345_ (.Y(_2040_),
    .A(_2037_),
    .B(_2039_));
 sg13g2_o21ai_1 _5346_ (.B1(net697),
    .Y(_2041_),
    .A1(net640),
    .A2(net1153));
 sg13g2_a21oi_1 _5347_ (.A1(net640),
    .A2(_2040_),
    .Y(_0333_),
    .B1(_2041_));
 sg13g2_xnor2_1 _5348_ (.Y(_2042_),
    .A(net978),
    .B(net737));
 sg13g2_a21oi_1 _5349_ (.A1(\project_audio.genblk1[2].n_c_oh_my.phase[9] ),
    .A2(\project_audio.freq[2][9] ),
    .Y(_2043_),
    .B1(_2037_));
 sg13g2_nor3_1 _5350_ (.A(_2038_),
    .B(_2042_),
    .C(_2043_),
    .Y(_2044_));
 sg13g2_o21ai_1 _5351_ (.B1(_2042_),
    .Y(_2045_),
    .A1(_2038_),
    .A2(_2043_));
 sg13g2_nand2b_1 _5352_ (.Y(_2046_),
    .B(_2045_),
    .A_N(_2044_));
 sg13g2_o21ai_1 _5353_ (.B1(net698),
    .Y(_2047_),
    .A1(net641),
    .A2(net978));
 sg13g2_a21oi_1 _5354_ (.A1(net640),
    .A2(_2046_),
    .Y(_0334_),
    .B1(_2047_));
 sg13g2_a21oi_1 _5355_ (.A1(\project_audio.genblk1[2].n_c_oh_my.phase[10] ),
    .A2(net737),
    .Y(_2048_),
    .B1(_2044_));
 sg13g2_nor2_1 _5356_ (.A(\project_audio.genblk1[2].n_c_oh_my.phase[11] ),
    .B(net445),
    .Y(_2049_));
 sg13g2_nand2_1 _5357_ (.Y(_2050_),
    .A(net953),
    .B(net445));
 sg13g2_nand2b_1 _5358_ (.Y(_2051_),
    .B(_2050_),
    .A_N(_2049_));
 sg13g2_xnor2_1 _5359_ (.Y(_2052_),
    .A(_2048_),
    .B(_2051_));
 sg13g2_o21ai_1 _5360_ (.B1(net697),
    .Y(_2053_),
    .A1(net640),
    .A2(net953));
 sg13g2_a21oi_1 _5361_ (.A1(net640),
    .A2(_2052_),
    .Y(_0335_),
    .B1(_2053_));
 sg13g2_o21ai_1 _5362_ (.B1(_2050_),
    .Y(_2054_),
    .A1(_2048_),
    .A2(_2049_));
 sg13g2_a21oi_1 _5363_ (.A1(net641),
    .A2(_2054_),
    .Y(_2055_),
    .B1(net514));
 sg13g2_nand3_1 _5364_ (.B(net514),
    .C(_2054_),
    .A(net641),
    .Y(_2056_));
 sg13g2_inv_1 _5365_ (.Y(_2057_),
    .A(_2056_));
 sg13g2_nor3_1 _5366_ (.A(net680),
    .B(_2055_),
    .C(_2057_),
    .Y(_0336_));
 sg13g2_nand2_1 _5367_ (.Y(_2058_),
    .A(net476),
    .B(_2057_));
 sg13g2_nand2_1 _5368_ (.Y(_2059_),
    .A(net696),
    .B(_2058_));
 sg13g2_a21oi_1 _5369_ (.A1(_2477_),
    .A2(_2056_),
    .Y(_0337_),
    .B1(_2059_));
 sg13g2_o21ai_1 _5370_ (.B1(net696),
    .Y(_2060_),
    .A1(_2476_),
    .A2(_2058_));
 sg13g2_a21oi_1 _5371_ (.A1(_2476_),
    .A2(_2058_),
    .Y(_0338_),
    .B1(_2060_));
 sg13g2_and4_1 _5372_ (.A(\project_audio.genblk1[2].n_c_oh_my.phase[14] ),
    .B(net476),
    .C(\project_audio.genblk1[2].n_c_oh_my.phase[12] ),
    .D(net696),
    .X(_2061_));
 sg13g2_nand3_1 _5373_ (.B(_2054_),
    .C(_2061_),
    .A(_1990_),
    .Y(_2062_));
 sg13g2_o21ai_1 _5374_ (.B1(_2062_),
    .Y(_0339_),
    .A1(_2475_),
    .A2(_2060_));
 sg13g2_nor2b_1 _5375_ (.A(net740),
    .B_N(net639),
    .Y(_2063_));
 sg13g2_o21ai_1 _5376_ (.B1(net697),
    .Y(_2064_),
    .A1(net642),
    .A2(net991));
 sg13g2_nor2_1 _5377_ (.A(_2063_),
    .B(_2064_),
    .Y(_0340_));
 sg13g2_nand2_1 _5378_ (.Y(_2065_),
    .A(net661),
    .B(net468));
 sg13g2_nand2_1 _5379_ (.Y(_2066_),
    .A(net919),
    .B(net468));
 sg13g2_xor2_1 _5380_ (.B(_2065_),
    .A(net919),
    .X(_2067_));
 sg13g2_nor2_1 _5381_ (.A(net683),
    .B(_2067_),
    .Y(_0341_));
 sg13g2_nand2_1 _5382_ (.Y(_2068_),
    .A(\project_audio.genblk1[1].n_c_oh_my.phase[1] ),
    .B(\project_audio.freq[1][1] ));
 sg13g2_xnor2_1 _5383_ (.Y(_2069_),
    .A(\project_audio.genblk1[1].n_c_oh_my.phase[1] ),
    .B(net747));
 sg13g2_xnor2_1 _5384_ (.Y(_2070_),
    .A(_2066_),
    .B(_2069_));
 sg13g2_o21ai_1 _5385_ (.B1(net710),
    .Y(_2071_),
    .A1(net658),
    .A2(net1021));
 sg13g2_a21oi_1 _5386_ (.A1(net658),
    .A2(_2070_),
    .Y(_0342_),
    .B1(_2071_));
 sg13g2_o21ai_1 _5387_ (.B1(_2068_),
    .Y(_2072_),
    .A1(_2066_),
    .A2(_2069_));
 sg13g2_and2_1 _5388_ (.A(\project_audio.genblk1[1].n_c_oh_my.phase[2] ),
    .B(\project_audio.freq[1][2] ),
    .X(_2073_));
 sg13g2_xor2_1 _5389_ (.B(\project_audio.freq[1][2] ),
    .A(\project_audio.genblk1[1].n_c_oh_my.phase[2] ),
    .X(_2074_));
 sg13g2_xnor2_1 _5390_ (.Y(_2075_),
    .A(_2072_),
    .B(_2074_));
 sg13g2_o21ai_1 _5391_ (.B1(net710),
    .Y(_2076_),
    .A1(net658),
    .A2(net985));
 sg13g2_a21oi_1 _5392_ (.A1(net658),
    .A2(_2075_),
    .Y(_0343_),
    .B1(_2076_));
 sg13g2_a21oi_2 _5393_ (.B1(_2073_),
    .Y(_2077_),
    .A2(_2074_),
    .A1(_2072_));
 sg13g2_nand2_1 _5394_ (.Y(_2078_),
    .A(\project_audio.genblk1[1].n_c_oh_my.phase[3] ),
    .B(\project_audio.freq[1][3] ));
 sg13g2_xnor2_1 _5395_ (.Y(_2079_),
    .A(net951),
    .B(net768));
 sg13g2_xnor2_1 _5396_ (.Y(_2080_),
    .A(_2077_),
    .B(_2079_));
 sg13g2_o21ai_1 _5397_ (.B1(net711),
    .Y(_2081_),
    .A1(net661),
    .A2(net951));
 sg13g2_a21oi_1 _5398_ (.A1(net661),
    .A2(_2080_),
    .Y(_0344_),
    .B1(_2081_));
 sg13g2_o21ai_1 _5399_ (.B1(_2078_),
    .Y(_2082_),
    .A1(_2077_),
    .A2(_2079_));
 sg13g2_and2_1 _5400_ (.A(\project_audio.genblk1[1].n_c_oh_my.phase[4] ),
    .B(\project_audio.freq[1][4] ),
    .X(_2083_));
 sg13g2_xor2_1 _5401_ (.B(net500),
    .A(net1108),
    .X(_2084_));
 sg13g2_xnor2_1 _5402_ (.Y(_2085_),
    .A(_2082_),
    .B(_2084_));
 sg13g2_o21ai_1 _5403_ (.B1(net711),
    .Y(_2086_),
    .A1(net660),
    .A2(net1108));
 sg13g2_a21oi_1 _5404_ (.A1(net660),
    .A2(_2085_),
    .Y(_0345_),
    .B1(_2086_));
 sg13g2_a21o_1 _5405_ (.A2(_2084_),
    .A1(_2082_),
    .B1(_2083_),
    .X(_2087_));
 sg13g2_or2_1 _5406_ (.X(_2088_),
    .B(\project_audio.freq[1][5] ),
    .A(\project_audio.genblk1[1].n_c_oh_my.phase[5] ));
 sg13g2_nand2_1 _5407_ (.Y(_2089_),
    .A(net896),
    .B(net478));
 sg13g2_nand2_1 _5408_ (.Y(_2090_),
    .A(_2088_),
    .B(_2089_));
 sg13g2_xor2_1 _5409_ (.B(_2090_),
    .A(_2087_),
    .X(_2091_));
 sg13g2_o21ai_1 _5410_ (.B1(net711),
    .Y(_2092_),
    .A1(net666),
    .A2(net896));
 sg13g2_a21oi_1 _5411_ (.A1(net666),
    .A2(_2091_),
    .Y(_0346_),
    .B1(_2092_));
 sg13g2_xnor2_1 _5412_ (.Y(_2093_),
    .A(\project_audio.genblk1[1].n_c_oh_my.phase[6] ),
    .B(\project_audio.freq[1][6] ));
 sg13g2_nand2_1 _5413_ (.Y(_2094_),
    .A(_2087_),
    .B(_2088_));
 sg13g2_a21oi_1 _5414_ (.A1(_2089_),
    .A2(_2094_),
    .Y(_2095_),
    .B1(_2093_));
 sg13g2_nand3_1 _5415_ (.B(_2093_),
    .C(_2094_),
    .A(_2089_),
    .Y(_2096_));
 sg13g2_nand2b_1 _5416_ (.Y(_2097_),
    .B(_2096_),
    .A_N(_2095_));
 sg13g2_o21ai_1 _5417_ (.B1(net711),
    .Y(_2098_),
    .A1(net660),
    .A2(net1012));
 sg13g2_a21oi_1 _5418_ (.A1(net660),
    .A2(_2097_),
    .Y(_0347_),
    .B1(_2098_));
 sg13g2_a21oi_1 _5419_ (.A1(\project_audio.genblk1[1].n_c_oh_my.phase[6] ),
    .A2(net750),
    .Y(_2099_),
    .B1(_2095_));
 sg13g2_nand2_1 _5420_ (.Y(_2100_),
    .A(\project_audio.genblk1[1].n_c_oh_my.phase[7] ),
    .B(net722));
 sg13g2_xnor2_1 _5421_ (.Y(_2101_),
    .A(net1010),
    .B(net722));
 sg13g2_or2_1 _5422_ (.X(_2102_),
    .B(_2101_),
    .A(_2099_));
 sg13g2_xnor2_1 _5423_ (.Y(_2103_),
    .A(_2099_),
    .B(_2101_));
 sg13g2_o21ai_1 _5424_ (.B1(net713),
    .Y(_2104_),
    .A1(net660),
    .A2(net1010));
 sg13g2_a21oi_1 _5425_ (.A1(net660),
    .A2(_2103_),
    .Y(_0348_),
    .B1(_2104_));
 sg13g2_xnor2_1 _5426_ (.Y(_2105_),
    .A(\project_audio.genblk1[1].n_c_oh_my.phase[8] ),
    .B(\project_audio.freq[1][8] ));
 sg13g2_a21oi_1 _5427_ (.A1(_2100_),
    .A2(_2102_),
    .Y(_2106_),
    .B1(_2105_));
 sg13g2_nand3_1 _5428_ (.B(_2102_),
    .C(_2105_),
    .A(_2100_),
    .Y(_2107_));
 sg13g2_nand2b_1 _5429_ (.Y(_2108_),
    .B(_2107_),
    .A_N(_2106_));
 sg13g2_o21ai_1 _5430_ (.B1(net711),
    .Y(_2109_),
    .A1(net659),
    .A2(net983));
 sg13g2_a21oi_1 _5431_ (.A1(net659),
    .A2(_2108_),
    .Y(_0349_),
    .B1(_2109_));
 sg13g2_a21o_1 _5432_ (.A2(\project_audio.freq[1][8] ),
    .A1(\project_audio.genblk1[1].n_c_oh_my.phase[8] ),
    .B1(_2106_),
    .X(_2110_));
 sg13g2_nor2_1 _5433_ (.A(\project_audio.genblk1[1].n_c_oh_my.phase[9] ),
    .B(\project_audio.freq[1][9] ),
    .Y(_2111_));
 sg13g2_xor2_1 _5434_ (.B(net825),
    .A(net1178),
    .X(_2112_));
 sg13g2_xnor2_1 _5435_ (.Y(_2113_),
    .A(_2110_),
    .B(_2112_));
 sg13g2_o21ai_1 _5436_ (.B1(net707),
    .Y(_2114_),
    .A1(net659),
    .A2(net1178));
 sg13g2_a21oi_1 _5437_ (.A1(net659),
    .A2(_2113_),
    .Y(_0350_),
    .B1(_2114_));
 sg13g2_xnor2_1 _5438_ (.Y(_2115_),
    .A(\project_audio.genblk1[1].n_c_oh_my.phase[10] ),
    .B(net522));
 sg13g2_a21oi_1 _5439_ (.A1(\project_audio.genblk1[1].n_c_oh_my.phase[9] ),
    .A2(\project_audio.freq[1][9] ),
    .Y(_2116_),
    .B1(_2110_));
 sg13g2_nor3_1 _5440_ (.A(_2111_),
    .B(_2115_),
    .C(_2116_),
    .Y(_2117_));
 sg13g2_o21ai_1 _5441_ (.B1(_2115_),
    .Y(_2118_),
    .A1(_2111_),
    .A2(_2116_));
 sg13g2_nand2b_1 _5442_ (.Y(_2119_),
    .B(_2118_),
    .A_N(_2117_));
 sg13g2_o21ai_1 _5443_ (.B1(net707),
    .Y(_2120_),
    .A1(net659),
    .A2(net1073));
 sg13g2_a21oi_1 _5444_ (.A1(net659),
    .A2(_2119_),
    .Y(_0351_),
    .B1(_2120_));
 sg13g2_a21oi_1 _5445_ (.A1(\project_audio.genblk1[1].n_c_oh_my.phase[10] ),
    .A2(\project_audio.freq[1][10] ),
    .Y(_2121_),
    .B1(_2117_));
 sg13g2_nor2_1 _5446_ (.A(\project_audio.genblk1[1].n_c_oh_my.phase[11] ),
    .B(\project_audio.freq[1][11] ),
    .Y(_2122_));
 sg13g2_nand2_1 _5447_ (.Y(_2123_),
    .A(net965),
    .B(\project_audio.freq[1][11] ));
 sg13g2_nand2b_1 _5448_ (.Y(_2124_),
    .B(_2123_),
    .A_N(_2122_));
 sg13g2_xnor2_1 _5449_ (.Y(_2125_),
    .A(_2121_),
    .B(_2124_));
 sg13g2_o21ai_1 _5450_ (.B1(net707),
    .Y(_2126_),
    .A1(net659),
    .A2(net965));
 sg13g2_a21oi_1 _5451_ (.A1(net659),
    .A2(_2125_),
    .Y(_0352_),
    .B1(_2126_));
 sg13g2_o21ai_1 _5452_ (.B1(_2123_),
    .Y(_2127_),
    .A1(_2121_),
    .A2(_2122_));
 sg13g2_a21oi_1 _5453_ (.A1(net645),
    .A2(_2127_),
    .Y(_2128_),
    .B1(net723));
 sg13g2_nand3_1 _5454_ (.B(net723),
    .C(_2127_),
    .A(net645),
    .Y(_2129_));
 sg13g2_inv_1 _5455_ (.Y(_2130_),
    .A(_2129_));
 sg13g2_nor3_1 _5456_ (.A(net683),
    .B(_2128_),
    .C(_2130_),
    .Y(_0353_));
 sg13g2_nand2_1 _5457_ (.Y(_2131_),
    .A(net483),
    .B(_2130_));
 sg13g2_nand2_1 _5458_ (.Y(_2132_),
    .A(net697),
    .B(_2131_));
 sg13g2_a21oi_1 _5459_ (.A1(_2474_),
    .A2(_2129_),
    .Y(_0354_),
    .B1(_2132_));
 sg13g2_o21ai_1 _5460_ (.B1(net697),
    .Y(_2133_),
    .A1(_2473_),
    .A2(_2131_));
 sg13g2_a21oi_1 _5461_ (.A1(_2473_),
    .A2(_2131_),
    .Y(_0355_),
    .B1(_2133_));
 sg13g2_and4_1 _5462_ (.A(net538),
    .B(net483),
    .C(net723),
    .D(net697),
    .X(_2134_));
 sg13g2_nand3_1 _5463_ (.B(_2127_),
    .C(_2134_),
    .A(_2063_),
    .Y(_2135_));
 sg13g2_o21ai_1 _5464_ (.B1(_2135_),
    .Y(_0356_),
    .A1(_2472_),
    .A2(_2133_));
 sg13g2_o21ai_1 _5465_ (.B1(net706),
    .Y(_2136_),
    .A1(net645),
    .A2(net758));
 sg13g2_a21oi_1 _5466_ (.A1(_2471_),
    .A2(net645),
    .Y(_0357_),
    .B1(_2136_));
 sg13g2_nand2_1 _5467_ (.Y(_2137_),
    .A(net650),
    .B(net479));
 sg13g2_nand2_1 _5468_ (.Y(_2138_),
    .A(net907),
    .B(net479));
 sg13g2_xor2_1 _5469_ (.B(_2137_),
    .A(net907),
    .X(_2139_));
 sg13g2_nor2_1 _5470_ (.A(net685),
    .B(_2139_),
    .Y(_0358_));
 sg13g2_nand2_1 _5471_ (.Y(_2140_),
    .A(\project_audio.genblk1[0].n_c_oh_my.phase[1] ),
    .B(\project_audio.freq[0][1] ));
 sg13g2_xnor2_1 _5472_ (.Y(_2141_),
    .A(net1096),
    .B(net728));
 sg13g2_xnor2_1 _5473_ (.Y(_2142_),
    .A(_2138_),
    .B(_2141_));
 sg13g2_o21ai_1 _5474_ (.B1(net710),
    .Y(_2143_),
    .A1(net656),
    .A2(net1096));
 sg13g2_a21oi_1 _5475_ (.A1(net656),
    .A2(_2142_),
    .Y(_0359_),
    .B1(_2143_));
 sg13g2_o21ai_1 _5476_ (.B1(_2140_),
    .Y(_2144_),
    .A1(_2138_),
    .A2(_2141_));
 sg13g2_and2_1 _5477_ (.A(\project_audio.genblk1[0].n_c_oh_my.phase[2] ),
    .B(\project_audio.freq[0][2] ),
    .X(_2145_));
 sg13g2_xor2_1 _5478_ (.B(net534),
    .A(net1053),
    .X(_2146_));
 sg13g2_xnor2_1 _5479_ (.Y(_2147_),
    .A(_2144_),
    .B(_2146_));
 sg13g2_o21ai_1 _5480_ (.B1(net709),
    .Y(_2148_),
    .A1(net656),
    .A2(net1053));
 sg13g2_a21oi_1 _5481_ (.A1(net656),
    .A2(_2147_),
    .Y(_0360_),
    .B1(_2148_));
 sg13g2_a21oi_1 _5482_ (.A1(_2144_),
    .A2(_2146_),
    .Y(_2149_),
    .B1(_2145_));
 sg13g2_nand2_1 _5483_ (.Y(_2150_),
    .A(\project_audio.genblk1[0].n_c_oh_my.phase[3] ),
    .B(\project_audio.freq[0][3] ));
 sg13g2_xnor2_1 _5484_ (.Y(_2151_),
    .A(net961),
    .B(net741));
 sg13g2_xnor2_1 _5485_ (.Y(_2152_),
    .A(_2149_),
    .B(_2151_));
 sg13g2_o21ai_1 _5486_ (.B1(net709),
    .Y(_2153_),
    .A1(net654),
    .A2(net961));
 sg13g2_a21oi_1 _5487_ (.A1(net654),
    .A2(_2152_),
    .Y(_0361_),
    .B1(_2153_));
 sg13g2_o21ai_1 _5488_ (.B1(_2150_),
    .Y(_2154_),
    .A1(_2149_),
    .A2(_2151_));
 sg13g2_and2_1 _5489_ (.A(\project_audio.genblk1[0].n_c_oh_my.phase[4] ),
    .B(\project_audio.freq[0][4] ),
    .X(_2155_));
 sg13g2_xor2_1 _5490_ (.B(net817),
    .A(net1036),
    .X(_2156_));
 sg13g2_xnor2_1 _5491_ (.Y(_2157_),
    .A(_2154_),
    .B(_2156_));
 sg13g2_o21ai_1 _5492_ (.B1(net709),
    .Y(_2158_),
    .A1(net654),
    .A2(net1036));
 sg13g2_a21oi_1 _5493_ (.A1(net654),
    .A2(_2157_),
    .Y(_0362_),
    .B1(_2158_));
 sg13g2_a21o_1 _5494_ (.A2(_2156_),
    .A1(_2154_),
    .B1(_2155_),
    .X(_2159_));
 sg13g2_or2_1 _5495_ (.X(_2160_),
    .B(\project_audio.freq[0][5] ),
    .A(\project_audio.genblk1[0].n_c_oh_my.phase[5] ));
 sg13g2_nand2_1 _5496_ (.Y(_2161_),
    .A(net928),
    .B(net463));
 sg13g2_nand2_1 _5497_ (.Y(_2162_),
    .A(_2160_),
    .B(_2161_));
 sg13g2_xor2_1 _5498_ (.B(_2162_),
    .A(_2159_),
    .X(_2163_));
 sg13g2_o21ai_1 _5499_ (.B1(net709),
    .Y(_2164_),
    .A1(net655),
    .A2(net928));
 sg13g2_a21oi_1 _5500_ (.A1(net655),
    .A2(_2163_),
    .Y(_0363_),
    .B1(_2164_));
 sg13g2_xnor2_1 _5501_ (.Y(_2165_),
    .A(\project_audio.genblk1[0].n_c_oh_my.phase[6] ),
    .B(\project_audio.freq[0][6] ));
 sg13g2_nand2_1 _5502_ (.Y(_2166_),
    .A(_2159_),
    .B(_2160_));
 sg13g2_a21oi_1 _5503_ (.A1(_2161_),
    .A2(_2166_),
    .Y(_2167_),
    .B1(_2165_));
 sg13g2_nand3_1 _5504_ (.B(_2165_),
    .C(_2166_),
    .A(_2161_),
    .Y(_2168_));
 sg13g2_nand2b_1 _5505_ (.Y(_2169_),
    .B(_2168_),
    .A_N(_2167_));
 sg13g2_o21ai_1 _5506_ (.B1(net709),
    .Y(_2170_),
    .A1(net655),
    .A2(net1091));
 sg13g2_a21oi_1 _5507_ (.A1(net655),
    .A2(_2169_),
    .Y(_0364_),
    .B1(_2170_));
 sg13g2_a21oi_1 _5508_ (.A1(\project_audio.genblk1[0].n_c_oh_my.phase[6] ),
    .A2(\project_audio.freq[0][6] ),
    .Y(_2171_),
    .B1(_2167_));
 sg13g2_nand2_1 _5509_ (.Y(_2172_),
    .A(\project_audio.genblk1[0].n_c_oh_my.phase[7] ),
    .B(net529));
 sg13g2_xnor2_1 _5510_ (.Y(_2173_),
    .A(net1075),
    .B(net529));
 sg13g2_or2_1 _5511_ (.X(_2174_),
    .B(_2173_),
    .A(_2171_));
 sg13g2_xnor2_1 _5512_ (.Y(_2175_),
    .A(_2171_),
    .B(_2173_));
 sg13g2_o21ai_1 _5513_ (.B1(net714),
    .Y(_2176_),
    .A1(net663),
    .A2(net1075));
 sg13g2_a21oi_1 _5514_ (.A1(net663),
    .A2(_2175_),
    .Y(_0365_),
    .B1(_2176_));
 sg13g2_xnor2_1 _5515_ (.Y(_2177_),
    .A(\project_audio.genblk1[0].n_c_oh_my.phase[8] ),
    .B(\project_audio.freq[0][8] ));
 sg13g2_a21oi_1 _5516_ (.A1(_2172_),
    .A2(_2174_),
    .Y(_2178_),
    .B1(_2177_));
 sg13g2_nand3_1 _5517_ (.B(_2174_),
    .C(_2177_),
    .A(_2172_),
    .Y(_2179_));
 sg13g2_nand2b_1 _5518_ (.Y(_2180_),
    .B(_2179_),
    .A_N(_2178_));
 sg13g2_o21ai_1 _5519_ (.B1(net714),
    .Y(_2181_),
    .A1(net663),
    .A2(net993));
 sg13g2_a21oi_1 _5520_ (.A1(net663),
    .A2(_2180_),
    .Y(_0366_),
    .B1(_2181_));
 sg13g2_a21o_1 _5521_ (.A2(\project_audio.freq[0][8] ),
    .A1(\project_audio.genblk1[0].n_c_oh_my.phase[8] ),
    .B1(_2178_),
    .X(_2182_));
 sg13g2_nor2_1 _5522_ (.A(\project_audio.genblk1[0].n_c_oh_my.phase[9] ),
    .B(\project_audio.freq[0][9] ),
    .Y(_2183_));
 sg13g2_xor2_1 _5523_ (.B(net836),
    .A(net1180),
    .X(_2184_));
 sg13g2_xnor2_1 _5524_ (.Y(_2185_),
    .A(_2182_),
    .B(_2184_));
 sg13g2_o21ai_1 _5525_ (.B1(net714),
    .Y(_2186_),
    .A1(net663),
    .A2(net1180));
 sg13g2_a21oi_1 _5526_ (.A1(net663),
    .A2(_2185_),
    .Y(_0367_),
    .B1(_2186_));
 sg13g2_xnor2_1 _5527_ (.Y(_2187_),
    .A(\project_audio.genblk1[0].n_c_oh_my.phase[10] ),
    .B(net832));
 sg13g2_a21oi_1 _5528_ (.A1(\project_audio.genblk1[0].n_c_oh_my.phase[9] ),
    .A2(\project_audio.freq[0][9] ),
    .Y(_2188_),
    .B1(_2182_));
 sg13g2_nor3_1 _5529_ (.A(_2183_),
    .B(_2187_),
    .C(_2188_),
    .Y(_2189_));
 sg13g2_o21ai_1 _5530_ (.B1(_2187_),
    .Y(_2190_),
    .A1(_2183_),
    .A2(_2188_));
 sg13g2_nand2b_1 _5531_ (.Y(_2191_),
    .B(_2190_),
    .A_N(_2189_));
 sg13g2_o21ai_1 _5532_ (.B1(net709),
    .Y(_2192_),
    .A1(net662),
    .A2(net1127));
 sg13g2_a21oi_1 _5533_ (.A1(net662),
    .A2(_2191_),
    .Y(_0368_),
    .B1(_2192_));
 sg13g2_a21oi_2 _5534_ (.B1(_2189_),
    .Y(_2193_),
    .A2(net832),
    .A1(\project_audio.genblk1[0].n_c_oh_my.phase[10] ));
 sg13g2_nand2_1 _5535_ (.Y(_2194_),
    .A(\project_audio.genblk1[0].n_c_oh_my.phase[11] ),
    .B(\project_audio.freq[0][11] ));
 sg13g2_xnor2_1 _5536_ (.Y(_2195_),
    .A(net1124),
    .B(net785));
 sg13g2_xnor2_1 _5537_ (.Y(_2196_),
    .A(_2193_),
    .B(_2195_));
 sg13g2_o21ai_1 _5538_ (.B1(net710),
    .Y(_2197_),
    .A1(net662),
    .A2(net1124));
 sg13g2_a21oi_1 _5539_ (.A1(net662),
    .A2(_2196_),
    .Y(_0369_),
    .B1(_2197_));
 sg13g2_o21ai_1 _5540_ (.B1(net662),
    .Y(_2198_),
    .A1(\project_audio.genblk1[0].n_c_oh_my.phase[11] ),
    .A2(\project_audio.freq[0][11] ));
 sg13g2_a21oi_2 _5541_ (.B1(_2198_),
    .Y(_2199_),
    .A2(_2194_),
    .A1(_2193_));
 sg13g2_and2_1 _5542_ (.A(net889),
    .B(_2199_),
    .X(_2200_));
 sg13g2_o21ai_1 _5543_ (.B1(net711),
    .Y(_2201_),
    .A1(net889),
    .A2(_2199_));
 sg13g2_nor2_1 _5544_ (.A(_2200_),
    .B(net890),
    .Y(_0370_));
 sg13g2_o21ai_1 _5545_ (.B1(net711),
    .Y(_2202_),
    .A1(net489),
    .A2(_2200_));
 sg13g2_a21oi_1 _5546_ (.A1(net489),
    .A2(_2200_),
    .Y(_0371_),
    .B1(_2202_));
 sg13g2_a21oi_1 _5547_ (.A1(\project_audio.genblk1[0].n_c_oh_my.phase[13] ),
    .A2(_2200_),
    .Y(_2203_),
    .B1(net449));
 sg13g2_and3_1 _5548_ (.X(_2204_),
    .A(net449),
    .B(\project_audio.genblk1[0].n_c_oh_my.phase[13] ),
    .C(_2200_));
 sg13g2_nor3_1 _5549_ (.A(net684),
    .B(net450),
    .C(_2204_),
    .Y(_0372_));
 sg13g2_o21ai_1 _5550_ (.B1(net707),
    .Y(_2205_),
    .A1(net455),
    .A2(_2204_));
 sg13g2_a21oi_1 _5551_ (.A1(net455),
    .A2(_2204_),
    .Y(_0373_),
    .B1(_2205_));
 sg13g2_nand2b_1 _5552_ (.Y(_2206_),
    .B(net578),
    .A_N(_0025_));
 sg13g2_o21ai_1 _5553_ (.B1(_2206_),
    .Y(_2207_),
    .A1(\project_audio.iter.mult2_shift[0] ),
    .A2(net569));
 sg13g2_nand2_1 _5554_ (.Y(_2208_),
    .A(net1082),
    .B(net553));
 sg13g2_a21oi_1 _5555_ (.A1(net884),
    .A2(net558),
    .Y(_2209_),
    .B1(net564));
 sg13g2_a21oi_1 _5556_ (.A1(_2208_),
    .A2(_2209_),
    .Y(_0374_),
    .B1(_2207_));
 sg13g2_nand2b_1 _5557_ (.Y(_2210_),
    .B(net579),
    .A_N(_0026_));
 sg13g2_o21ai_1 _5558_ (.B1(_2210_),
    .Y(_2211_),
    .A1(net884),
    .A2(net570));
 sg13g2_nand2_1 _5559_ (.Y(_2212_),
    .A(\project_audio.iter.mult_accum[17] ),
    .B(net553));
 sg13g2_a21oi_1 _5560_ (.A1(net845),
    .A2(net558),
    .Y(_2213_),
    .B1(net564));
 sg13g2_a21oi_1 _5561_ (.A1(_2212_),
    .A2(_2213_),
    .Y(_0375_),
    .B1(net885));
 sg13g2_a22oi_1 _5562_ (.Y(_2214_),
    .B1(net579),
    .B2(_0027_),
    .A2(net583),
    .A1(net845));
 sg13g2_nor2b_1 _5563_ (.A(\project_audio.iter.mult2_shift[3] ),
    .B_N(net558),
    .Y(_2215_));
 sg13g2_o21ai_1 _5564_ (.B1(_2549_),
    .Y(_2216_),
    .A1(\project_audio.iter.mult_accum[18] ),
    .A2(net558));
 sg13g2_o21ai_1 _5565_ (.B1(net846),
    .Y(_0376_),
    .A1(_2215_),
    .A2(_2216_));
 sg13g2_nand2b_1 _5566_ (.Y(_2217_),
    .B(net578),
    .A_N(_0028_));
 sg13g2_o21ai_1 _5567_ (.B1(_2217_),
    .Y(_2218_),
    .A1(net934),
    .A2(net570));
 sg13g2_nand2_1 _5568_ (.Y(_2219_),
    .A(\project_audio.iter.mult_accum[19] ),
    .B(net553));
 sg13g2_a21oi_1 _5569_ (.A1(net855),
    .A2(net558),
    .Y(_2220_),
    .B1(net564));
 sg13g2_a21oi_1 _5570_ (.A1(_2219_),
    .A2(_2220_),
    .Y(_0377_),
    .B1(net935));
 sg13g2_nand2b_1 _5571_ (.Y(_2221_),
    .B(net578),
    .A_N(_0029_));
 sg13g2_o21ai_1 _5572_ (.B1(_2221_),
    .Y(_2222_),
    .A1(net855),
    .A2(net571));
 sg13g2_nand2_1 _5573_ (.Y(_2223_),
    .A(\project_audio.iter.mult_accum[20] ),
    .B(net553));
 sg13g2_a21oi_1 _5574_ (.A1(\project_audio.iter.mult2_shift[5] ),
    .A2(net558),
    .Y(_2224_),
    .B1(net564));
 sg13g2_a21oi_1 _5575_ (.A1(_2223_),
    .A2(_2224_),
    .Y(_0378_),
    .B1(net856));
 sg13g2_nand2b_1 _5576_ (.Y(_2225_),
    .B(net578),
    .A_N(_0030_));
 sg13g2_o21ai_1 _5577_ (.B1(_2225_),
    .Y(_2226_),
    .A1(net897),
    .A2(net571));
 sg13g2_nand2_1 _5578_ (.Y(_2227_),
    .A(\project_audio.iter.mult_accum[21] ),
    .B(net553));
 sg13g2_a21oi_1 _5579_ (.A1(net893),
    .A2(net558),
    .Y(_2228_),
    .B1(net564));
 sg13g2_a21oi_1 _5580_ (.A1(_2227_),
    .A2(_2228_),
    .Y(_0379_),
    .B1(net898));
 sg13g2_nand2b_1 _5581_ (.Y(_2229_),
    .B(net578),
    .A_N(_0031_));
 sg13g2_o21ai_1 _5582_ (.B1(_2229_),
    .Y(_2230_),
    .A1(net893),
    .A2(net571));
 sg13g2_nand2_1 _5583_ (.Y(_2231_),
    .A(\project_audio.iter.mult_accum[22] ),
    .B(net553));
 sg13g2_a21oi_1 _5584_ (.A1(\project_audio.iter.mult2_shift[7] ),
    .A2(net559),
    .Y(_2232_),
    .B1(net564));
 sg13g2_a21oi_1 _5585_ (.A1(_2231_),
    .A2(_2232_),
    .Y(_0380_),
    .B1(net894));
 sg13g2_nand2b_1 _5586_ (.Y(_2233_),
    .B(net578),
    .A_N(_0032_));
 sg13g2_o21ai_1 _5587_ (.B1(_2233_),
    .Y(_2234_),
    .A1(net914),
    .A2(net571));
 sg13g2_nand2_1 _5588_ (.Y(_2235_),
    .A(\project_audio.iter.mult_accum[23] ),
    .B(net553));
 sg13g2_a21oi_1 _5589_ (.A1(net833),
    .A2(net558),
    .Y(_2236_),
    .B1(net564));
 sg13g2_a21oi_1 _5590_ (.A1(_2235_),
    .A2(_2236_),
    .Y(_0381_),
    .B1(net915));
 sg13g2_a22oi_1 _5591_ (.Y(_2237_),
    .B1(net578),
    .B2(_0033_),
    .A2(net583),
    .A1(net833));
 sg13g2_nor2b_1 _5592_ (.A(\project_audio.iter.mult2_shift[9] ),
    .B_N(net561),
    .Y(_2238_));
 sg13g2_o21ai_1 _5593_ (.B1(_2549_),
    .Y(_2239_),
    .A1(\project_audio.iter.mult_accum[24] ),
    .A2(net559));
 sg13g2_o21ai_1 _5594_ (.B1(net834),
    .Y(_0382_),
    .A1(_2238_),
    .A2(_2239_));
 sg13g2_nand2b_1 _5595_ (.Y(_2240_),
    .B(net579),
    .A_N(_0034_));
 sg13g2_o21ai_1 _5596_ (.B1(_2240_),
    .Y(_2241_),
    .A1(\project_audio.iter.mult2_shift[9] ),
    .A2(net575));
 sg13g2_nand2_1 _5597_ (.Y(_2242_),
    .A(\project_audio.iter.mult_accum[25] ),
    .B(net554));
 sg13g2_a21oi_1 _5598_ (.A1(net878),
    .A2(net561),
    .Y(_2243_),
    .B1(net564));
 sg13g2_a21oi_1 _5599_ (.A1(_2242_),
    .A2(_2243_),
    .Y(_0383_),
    .B1(_2241_));
 sg13g2_nand2b_1 _5600_ (.Y(_2244_),
    .B(net579),
    .A_N(_0035_));
 sg13g2_o21ai_1 _5601_ (.B1(_2244_),
    .Y(_2245_),
    .A1(net878),
    .A2(net575));
 sg13g2_nand2_1 _5602_ (.Y(_2246_),
    .A(net901),
    .B(net554));
 sg13g2_a21oi_1 _5603_ (.A1(net872),
    .A2(net561),
    .Y(_2247_),
    .B1(net565));
 sg13g2_a21oi_1 _5604_ (.A1(_2246_),
    .A2(_2247_),
    .Y(_0384_),
    .B1(_2245_));
 sg13g2_nand2b_1 _5605_ (.Y(_2248_),
    .B(net580),
    .A_N(_0036_));
 sg13g2_o21ai_1 _5606_ (.B1(_2248_),
    .Y(_2249_),
    .A1(net872),
    .A2(net575));
 sg13g2_nand2_1 _5607_ (.Y(_2250_),
    .A(\project_audio.iter.mult_accum[27] ),
    .B(net554));
 sg13g2_a21oi_1 _5608_ (.A1(net869),
    .A2(net560),
    .Y(_2251_),
    .B1(net565));
 sg13g2_a21oi_1 _5609_ (.A1(_2250_),
    .A2(_2251_),
    .Y(_0385_),
    .B1(net873));
 sg13g2_nand2b_1 _5610_ (.Y(_2252_),
    .B(net579),
    .A_N(_0037_));
 sg13g2_o21ai_1 _5611_ (.B1(_2252_),
    .Y(_2253_),
    .A1(net869),
    .A2(net575));
 sg13g2_nand2_1 _5612_ (.Y(_2254_),
    .A(\project_audio.iter.mult_accum[28] ),
    .B(net554));
 sg13g2_a21oi_1 _5613_ (.A1(\project_audio.iter.mult2_shift[13] ),
    .A2(net560),
    .Y(_2255_),
    .B1(net565));
 sg13g2_a21oi_1 _5614_ (.A1(_2254_),
    .A2(_2255_),
    .Y(_0386_),
    .B1(net870));
 sg13g2_nand2b_1 _5615_ (.Y(_2256_),
    .B(net579),
    .A_N(_0038_));
 sg13g2_o21ai_1 _5616_ (.B1(_2256_),
    .Y(_2257_),
    .A1(net922),
    .A2(net575));
 sg13g2_nand2_1 _5617_ (.Y(_2258_),
    .A(\project_audio.iter.mult_accum[29] ),
    .B(net554));
 sg13g2_a21oi_1 _5618_ (.A1(\project_audio.iter.mult2_shift[14] ),
    .A2(net560),
    .Y(_2259_),
    .B1(net565));
 sg13g2_a21oi_1 _5619_ (.A1(_2258_),
    .A2(_2259_),
    .Y(_0387_),
    .B1(net923));
 sg13g2_nand2b_1 _5620_ (.Y(_2260_),
    .B(net579),
    .A_N(_0039_));
 sg13g2_o21ai_1 _5621_ (.B1(_2260_),
    .Y(_2261_),
    .A1(\project_audio.iter.mult2_shift[14] ),
    .A2(net575));
 sg13g2_nand2_1 _5622_ (.Y(_2262_),
    .A(\project_audio.iter.mult_accum[30] ),
    .B(net554));
 sg13g2_a21oi_1 _5623_ (.A1(net863),
    .A2(net560),
    .Y(_2263_),
    .B1(net565));
 sg13g2_a21oi_1 _5624_ (.A1(_2262_),
    .A2(_2263_),
    .Y(_0388_),
    .B1(_2261_));
 sg13g2_nand3_1 _5625_ (.B(_2537_),
    .C(net576),
    .A(\project_audio.iter.mult_accum[31] ),
    .Y(_2264_));
 sg13g2_a22oi_1 _5626_ (.Y(_2265_),
    .B1(net580),
    .B2(net505),
    .A2(net583),
    .A1(\project_audio.iter.mult2_shift[15] ));
 sg13g2_nand2_1 _5627_ (.Y(_0389_),
    .A(_2264_),
    .B(net506));
 sg13g2_nand2_1 _5628_ (.Y(_2266_),
    .A(\project_audio.genblk1[3].n_c_oh_my.snd ),
    .B(\project_audio.genblk1[4].n_c_oh_my.snd ));
 sg13g2_xor2_1 _5629_ (.B(\project_audio.genblk1[4].n_c_oh_my.snd ),
    .A(\project_audio.genblk1[3].n_c_oh_my.snd ),
    .X(_2267_));
 sg13g2_nand2_1 _5630_ (.Y(_2268_),
    .A(\project_audio.genblk1[1].n_c_oh_my.snd ),
    .B(_2267_));
 sg13g2_nand4_1 _5631_ (.B(\project_audio.iter.r[13] ),
    .C(\project_audio.iter.r[12] ),
    .A(\project_audio.iter.r[16] ),
    .Y(_2269_),
    .D(\project_audio.iter.r[11] ));
 sg13g2_nand2b_1 _5632_ (.Y(_2270_),
    .B(\project_audio.iter.r[15] ),
    .A_N(\project_audio.iter.r[14] ));
 sg13g2_nor3_2 _5633_ (.A(_0004_),
    .B(_2269_),
    .C(_2270_),
    .Y(_2271_));
 sg13g2_nand2_1 _5634_ (.Y(_2272_),
    .A(\project_audio.iter.r[11] ),
    .B(\project_audio.iter.r[10] ));
 sg13g2_nand2_1 _5635_ (.Y(_2273_),
    .A(\project_audio.iter.r[15] ),
    .B(\project_audio.iter.r[14] ));
 sg13g2_nand4_1 _5636_ (.B(\project_audio.iter.r[14] ),
    .C(\project_audio.iter.r[12] ),
    .A(\project_audio.iter.r[15] ),
    .Y(_2274_),
    .D(_2272_));
 sg13g2_nand2b_1 _5637_ (.Y(_2275_),
    .B(_2274_),
    .A_N(\project_audio.iter.r[13] ));
 sg13g2_and2_1 _5638_ (.A(\project_audio.iter.r[17] ),
    .B(\project_audio.iter.r[16] ),
    .X(_2276_));
 sg13g2_nand2_2 _5639_ (.Y(_2277_),
    .A(\project_audio.iter.r[17] ),
    .B(\project_audio.iter.r[16] ));
 sg13g2_or4_1 _5640_ (.A(\project_audio.iter.r[12] ),
    .B(\project_audio.iter.r[11] ),
    .C(\project_audio.iter.r[10] ),
    .D(_2270_),
    .X(_2278_));
 sg13g2_a21oi_1 _5641_ (.A1(\project_audio.iter.r[13] ),
    .A2(_2278_),
    .Y(_2279_),
    .B1(_2277_));
 sg13g2_a21oi_2 _5642_ (.B1(_2271_),
    .Y(_2280_),
    .A2(_2279_),
    .A1(_2275_));
 sg13g2_inv_1 _5643_ (.Y(_2281_),
    .A(_2280_));
 sg13g2_xor2_1 _5644_ (.B(_2267_),
    .A(\project_audio.genblk1[1].n_c_oh_my.snd ),
    .X(_2282_));
 sg13g2_nand3_1 _5645_ (.B(_2280_),
    .C(_2282_),
    .A(\project_audio.genblk1[6].n_c_oh_my.snd ),
    .Y(_2283_));
 sg13g2_nand2b_2 _5646_ (.Y(_2284_),
    .B(\project_audio.genblk1[5].n_c_oh_my.snd ),
    .A_N(_2271_));
 sg13g2_a21o_1 _5647_ (.A2(_2280_),
    .A1(\project_audio.genblk1[6].n_c_oh_my.snd ),
    .B1(_2282_),
    .X(_2285_));
 sg13g2_and2_1 _5648_ (.A(_2283_),
    .B(_2285_),
    .X(_2286_));
 sg13g2_nand2b_1 _5649_ (.Y(_2287_),
    .B(_2286_),
    .A_N(_2284_));
 sg13g2_a22oi_1 _5650_ (.Y(_2288_),
    .B1(_2283_),
    .B2(_2287_),
    .A2(_2268_),
    .A1(_2266_));
 sg13g2_nand4_1 _5651_ (.B(_2268_),
    .C(_2283_),
    .A(_2266_),
    .Y(_2289_),
    .D(_2287_));
 sg13g2_nand2b_1 _5652_ (.Y(_2290_),
    .B(_2289_),
    .A_N(_2288_));
 sg13g2_xnor2_1 _5653_ (.Y(_2291_),
    .A(_2284_),
    .B(_2286_));
 sg13g2_nand2_1 _5654_ (.Y(_2292_),
    .A(\project_audio.genblk1[0].n_c_oh_my.snd ),
    .B(_2291_));
 sg13g2_nand2_1 _5655_ (.Y(_2293_),
    .A(\project_audio.genblk1[7].n_c_oh_my.snd ),
    .B(_2280_));
 sg13g2_nor2_1 _5656_ (.A(\project_audio.genblk1[0].n_c_oh_my.snd ),
    .B(_2291_),
    .Y(_2294_));
 sg13g2_xor2_1 _5657_ (.B(_2291_),
    .A(\project_audio.genblk1[0].n_c_oh_my.snd ),
    .X(_2295_));
 sg13g2_o21ai_1 _5658_ (.B1(_2292_),
    .Y(_2296_),
    .A1(_2293_),
    .A2(_2294_));
 sg13g2_nand2b_1 _5659_ (.Y(_2297_),
    .B(_2296_),
    .A_N(_2290_));
 sg13g2_xnor2_1 _5660_ (.Y(_2298_),
    .A(_2293_),
    .B(_2295_));
 sg13g2_nand2_1 _5661_ (.Y(_2299_),
    .A(\project_audio.genblk1[2].n_c_oh_my.snd ),
    .B(_2298_));
 sg13g2_xor2_1 _5662_ (.B(_2296_),
    .A(_2290_),
    .X(_2300_));
 sg13g2_o21ai_1 _5663_ (.B1(_2297_),
    .Y(_2301_),
    .A1(_2299_),
    .A2(_2300_));
 sg13g2_inv_1 _5664_ (.Y(_2302_),
    .A(_2301_));
 sg13g2_a21oi_1 _5665_ (.A1(net875),
    .A2(_2302_),
    .Y(_2303_),
    .B1(net766));
 sg13g2_nor2_1 _5666_ (.A(\project_audio.mixer.counter[2] ),
    .B(_2302_),
    .Y(_2304_));
 sg13g2_o21ai_1 _5667_ (.B1(_2303_),
    .Y(_2305_),
    .A1(_2288_),
    .A2(_2304_));
 sg13g2_xnor2_1 _5668_ (.Y(_2306_),
    .A(_2299_),
    .B(_2300_));
 sg13g2_nor2_1 _5669_ (.A(\project_audio.mixer.counter[1] ),
    .B(_2306_),
    .Y(_2307_));
 sg13g2_xor2_1 _5670_ (.B(_2298_),
    .A(\project_audio.genblk1[2].n_c_oh_my.snd ),
    .X(_2308_));
 sg13g2_nor3_1 _5671_ (.A(\project_audio.mixer.counter[0] ),
    .B(_0041_),
    .C(_2308_),
    .Y(_2309_));
 sg13g2_a21o_1 _5672_ (.A2(_2308_),
    .A1(_0041_),
    .B1(_2309_),
    .X(_2310_));
 sg13g2_nand2_1 _5673_ (.Y(_2311_),
    .A(net1214),
    .B(_2306_));
 sg13g2_o21ai_1 _5674_ (.B1(_2311_),
    .Y(_2312_),
    .A1(_2307_),
    .A2(_2310_));
 sg13g2_and2_1 _5675_ (.A(_2305_),
    .B(_2312_),
    .X(_2313_));
 sg13g2_o21ai_1 _5676_ (.B1(net766),
    .Y(_2314_),
    .A1(net875),
    .A2(_2302_));
 sg13g2_a21oi_1 _5677_ (.A1(_2288_),
    .A2(_2314_),
    .Y(_2315_),
    .B1(_2303_));
 sg13g2_nor3_1 _5678_ (.A(net681),
    .B(net1215),
    .C(_2315_),
    .Y(_0390_));
 sg13g2_and2_1 _5679_ (.A(net696),
    .B(net443),
    .X(_0391_));
 sg13g2_o21ai_1 _5680_ (.B1(net696),
    .Y(_2316_),
    .A1(net865),
    .A2(\project_audio.mixer.counter[0] ));
 sg13g2_a21oi_1 _5681_ (.A1(net865),
    .A2(\project_audio.mixer.counter[0] ),
    .Y(_0392_),
    .B1(_2316_));
 sg13g2_a21oi_1 _5682_ (.A1(net865),
    .A2(\project_audio.mixer.counter[0] ),
    .Y(_2317_),
    .B1(net875));
 sg13g2_and3_1 _5683_ (.X(_2318_),
    .A(net875),
    .B(net865),
    .C(\project_audio.mixer.counter[0] ));
 sg13g2_nor3_1 _5684_ (.A(net681),
    .B(net876),
    .C(_2318_),
    .Y(_0393_));
 sg13g2_o21ai_1 _5685_ (.B1(net696),
    .Y(_2319_),
    .A1(net766),
    .A2(_2318_));
 sg13g2_a21oi_1 _5686_ (.A1(net766),
    .A2(_2318_),
    .Y(_0394_),
    .B1(_2319_));
 sg13g2_or4_1 _5687_ (.A(\project_audio.nco_increment_gen.counter[5] ),
    .B(\project_audio.nco_increment_gen.counter[4] ),
    .C(\project_audio.nco_increment_gen.counter[3] ),
    .D(net464),
    .X(_2320_));
 sg13g2_or3_1 _5688_ (.A(net459),
    .B(\project_audio.nco_increment_gen.counter[6] ),
    .C(_1335_),
    .X(_2321_));
 sg13g2_nor4_1 _5689_ (.A(\project_audio.nco_increment_gen.counter[0] ),
    .B(net497),
    .C(_2320_),
    .D(_2321_),
    .Y(_0395_));
 sg13g2_a21oi_1 _5690_ (.A1(_2452_),
    .A2(net552),
    .Y(_2322_),
    .B1(net562));
 sg13g2_o21ai_1 _5691_ (.B1(_2322_),
    .Y(_2323_),
    .A1(net1170),
    .A2(net552));
 sg13g2_o21ai_1 _5692_ (.B1(_2323_),
    .Y(_0396_),
    .A1(_2516_),
    .A2(net567));
 sg13g2_nand2_1 _5693_ (.Y(_2324_),
    .A(net959),
    .B(net583));
 sg13g2_o21ai_1 _5694_ (.B1(_2549_),
    .Y(_2325_),
    .A1(\project_audio.iter.r[17] ),
    .A2(net555));
 sg13g2_nor2_1 _5695_ (.A(\project_audio.iter.mult1_shift[16] ),
    .B(net553),
    .Y(_2326_));
 sg13g2_o21ai_1 _5696_ (.B1(_2324_),
    .Y(_0397_),
    .A1(_2325_),
    .A2(_2326_));
 sg13g2_nand4_1 _5697_ (.B(_2511_),
    .C(\project_audio.iter.counter[5] ),
    .A(\project_audio.iter.counter[1] ),
    .Y(_2327_),
    .D(_2521_));
 sg13g2_or2_1 _5698_ (.X(_2328_),
    .B(_2327_),
    .A(_2526_));
 sg13g2_o21ai_1 _5699_ (.B1(net686),
    .Y(_2329_),
    .A1(net1082),
    .A2(net586));
 sg13g2_a21oi_1 _5700_ (.A1(_2469_),
    .A2(net586),
    .Y(_0398_),
    .B1(_2329_));
 sg13g2_o21ai_1 _5701_ (.B1(net687),
    .Y(_2330_),
    .A1(net1194),
    .A2(net584));
 sg13g2_a21oi_1 _5702_ (.A1(_2468_),
    .A2(net584),
    .Y(_0399_),
    .B1(_2330_));
 sg13g2_o21ai_1 _5703_ (.B1(net686),
    .Y(_2331_),
    .A1(net1176),
    .A2(net585));
 sg13g2_a21oi_1 _5704_ (.A1(_2467_),
    .A2(net584),
    .Y(_0400_),
    .B1(_2331_));
 sg13g2_o21ai_1 _5705_ (.B1(net686),
    .Y(_2332_),
    .A1(\project_audio.iter.mult_accum[19] ),
    .A2(net584));
 sg13g2_a21oi_1 _5706_ (.A1(_2466_),
    .A2(net584),
    .Y(_0401_),
    .B1(_2332_));
 sg13g2_o21ai_1 _5707_ (.B1(net687),
    .Y(_2333_),
    .A1(net1205),
    .A2(net584));
 sg13g2_a21oi_1 _5708_ (.A1(_2465_),
    .A2(net584),
    .Y(_0402_),
    .B1(_2333_));
 sg13g2_o21ai_1 _5709_ (.B1(net687),
    .Y(_2334_),
    .A1(net1177),
    .A2(net584));
 sg13g2_a21oi_1 _5710_ (.A1(_2464_),
    .A2(net586),
    .Y(_0403_),
    .B1(_2334_));
 sg13g2_o21ai_1 _5711_ (.B1(net686),
    .Y(_2335_),
    .A1(net1162),
    .A2(net586));
 sg13g2_a21oi_1 _5712_ (.A1(_2463_),
    .A2(net586),
    .Y(_0404_),
    .B1(_2335_));
 sg13g2_o21ai_1 _5713_ (.B1(net686),
    .Y(_2336_),
    .A1(\project_audio.iter.mult_accum[23] ),
    .A2(net585));
 sg13g2_a21oi_1 _5714_ (.A1(_2462_),
    .A2(net585),
    .Y(_0405_),
    .B1(_2336_));
 sg13g2_o21ai_1 _5715_ (.B1(net686),
    .Y(_2337_),
    .A1(net1006),
    .A2(net585));
 sg13g2_a21oi_1 _5716_ (.A1(_2461_),
    .A2(net585),
    .Y(_0406_),
    .B1(_2337_));
 sg13g2_o21ai_1 _5717_ (.B1(net686),
    .Y(_2338_),
    .A1(net1184),
    .A2(net585));
 sg13g2_a21oi_1 _5718_ (.A1(_2460_),
    .A2(net585),
    .Y(_0407_),
    .B1(_2338_));
 sg13g2_o21ai_1 _5719_ (.B1(net687),
    .Y(_2339_),
    .A1(net901),
    .A2(net587));
 sg13g2_a21oi_1 _5720_ (.A1(_2459_),
    .A2(net587),
    .Y(_0408_),
    .B1(_2339_));
 sg13g2_o21ai_1 _5721_ (.B1(net686),
    .Y(_2340_),
    .A1(net1181),
    .A2(net587));
 sg13g2_a21oi_1 _5722_ (.A1(_2458_),
    .A2(net587),
    .Y(_0409_),
    .B1(_2340_));
 sg13g2_a21oi_1 _5723_ (.A1(net629),
    .A2(net588),
    .Y(_2341_),
    .B1(net682));
 sg13g2_o21ai_1 _5724_ (.B1(_2341_),
    .Y(_0410_),
    .A1(_2457_),
    .A2(net588));
 sg13g2_o21ai_1 _5725_ (.B1(net688),
    .Y(_2342_),
    .A1(net1106),
    .A2(net588));
 sg13g2_a21oi_1 _5726_ (.A1(_2455_),
    .A2(net588),
    .Y(_0411_),
    .B1(_2342_));
 sg13g2_o21ai_1 _5727_ (.B1(net689),
    .Y(_2343_),
    .A1(net949),
    .A2(net587));
 sg13g2_a21oi_1 _5728_ (.A1(_2454_),
    .A2(net587),
    .Y(_0412_),
    .B1(_2343_));
 sg13g2_o21ai_1 _5729_ (.B1(net688),
    .Y(_2344_),
    .A1(net1030),
    .A2(net587));
 sg13g2_a21oi_1 _5730_ (.A1(_2453_),
    .A2(net587),
    .Y(_0413_),
    .B1(_2344_));
 sg13g2_nor2_1 _5731_ (.A(net682),
    .B(net589),
    .Y(_0414_));
 sg13g2_nand4_1 _5732_ (.B(\project_audio.iter.counter[10] ),
    .C(\project_audio.iter.counter[13] ),
    .A(\project_audio.iter.counter[11] ),
    .Y(_2345_),
    .D(\project_audio.iter.counter[12] ));
 sg13g2_nand2_1 _5733_ (.Y(_2346_),
    .A(net690),
    .B(_2345_));
 sg13g2_and3_1 _5734_ (.X(_0415_),
    .A(net690),
    .B(net437),
    .C(_2345_));
 sg13g2_and2_1 _5735_ (.A(\project_audio.iter.counter[1] ),
    .B(net1211),
    .X(_2347_));
 sg13g2_nor3_1 _5736_ (.A(_2535_),
    .B(net617),
    .C(net1212),
    .Y(_0416_));
 sg13g2_and2_1 _5737_ (.A(net944),
    .B(_2347_),
    .X(_2348_));
 sg13g2_nor2_1 _5738_ (.A(net944),
    .B(_2347_),
    .Y(_2349_));
 sg13g2_nor3_1 _5739_ (.A(net617),
    .B(_2348_),
    .C(net945),
    .Y(_0417_));
 sg13g2_nor2_1 _5740_ (.A(net1090),
    .B(_2348_),
    .Y(_2350_));
 sg13g2_and2_1 _5741_ (.A(net1090),
    .B(_2348_),
    .X(_2351_));
 sg13g2_nor3_1 _5742_ (.A(net617),
    .B(_2350_),
    .C(_2351_),
    .Y(_0418_));
 sg13g2_nor2_1 _5743_ (.A(net1161),
    .B(_2351_),
    .Y(_2352_));
 sg13g2_and2_1 _5744_ (.A(net1161),
    .B(_2351_),
    .X(_2353_));
 sg13g2_nor3_1 _5745_ (.A(net617),
    .B(_2352_),
    .C(_2353_),
    .Y(_0419_));
 sg13g2_nor2_1 _5746_ (.A(net1098),
    .B(_2353_),
    .Y(_2354_));
 sg13g2_and2_1 _5747_ (.A(net1098),
    .B(_2353_),
    .X(_2355_));
 sg13g2_nor3_1 _5748_ (.A(net617),
    .B(net1099),
    .C(_2355_),
    .Y(_0420_));
 sg13g2_nor2_1 _5749_ (.A(net1046),
    .B(_2355_),
    .Y(_2356_));
 sg13g2_and2_1 _5750_ (.A(net1046),
    .B(_2355_),
    .X(_2357_));
 sg13g2_nor3_1 _5751_ (.A(net616),
    .B(net1047),
    .C(_2357_),
    .Y(_0421_));
 sg13g2_nor2_1 _5752_ (.A(net1050),
    .B(_2357_),
    .Y(_2358_));
 sg13g2_and2_1 _5753_ (.A(net1050),
    .B(_2357_),
    .X(_2359_));
 sg13g2_nor3_1 _5754_ (.A(net616),
    .B(_2358_),
    .C(_2359_),
    .Y(_0422_));
 sg13g2_nor2_1 _5755_ (.A(net971),
    .B(_2359_),
    .Y(_2360_));
 sg13g2_and2_1 _5756_ (.A(net971),
    .B(_2359_),
    .X(_2361_));
 sg13g2_nor3_1 _5757_ (.A(net616),
    .B(net972),
    .C(_2361_),
    .Y(_0423_));
 sg13g2_nor2_1 _5758_ (.A(net841),
    .B(_2361_),
    .Y(_2362_));
 sg13g2_and2_1 _5759_ (.A(net841),
    .B(_2361_),
    .X(_2363_));
 sg13g2_nor3_1 _5760_ (.A(net616),
    .B(net842),
    .C(_2363_),
    .Y(_0424_));
 sg13g2_nor2_1 _5761_ (.A(net1066),
    .B(_2363_),
    .Y(_2364_));
 sg13g2_and2_1 _5762_ (.A(net1066),
    .B(_2363_),
    .X(_2365_));
 sg13g2_nor3_1 _5763_ (.A(net616),
    .B(_2364_),
    .C(_2365_),
    .Y(_0425_));
 sg13g2_nor2_1 _5764_ (.A(net1048),
    .B(_2365_),
    .Y(_2366_));
 sg13g2_and2_1 _5765_ (.A(net1048),
    .B(_2365_),
    .X(_2367_));
 sg13g2_nor3_1 _5766_ (.A(net616),
    .B(net1049),
    .C(_2367_),
    .Y(_0426_));
 sg13g2_xnor2_1 _5767_ (.Y(_2368_),
    .A(net1061),
    .B(_2367_));
 sg13g2_nor2_1 _5768_ (.A(net616),
    .B(_2368_),
    .Y(_0427_));
 sg13g2_a21oi_1 _5769_ (.A1(\project_audio.iter.counter[12] ),
    .A2(_2367_),
    .Y(_2369_),
    .B1(net774));
 sg13g2_nor2_1 _5770_ (.A(net616),
    .B(net775),
    .Y(_0428_));
 sg13g2_nor2_1 _5771_ (.A(\project_audio.iter.next_ready ),
    .B(net682),
    .Y(_2370_));
 sg13g2_a22oi_1 _5772_ (.Y(_2371_),
    .B1(_2370_),
    .B2(\project_audio.r_counter ),
    .A2(_0498_),
    .A1(net441));
 sg13g2_inv_1 _5773_ (.Y(_0429_),
    .A(net442));
 sg13g2_and2_2 _5774_ (.A(\project_audio.iter.next_ready ),
    .B(\project_audio.r_counter ),
    .X(_2372_));
 sg13g2_nand2_2 _5775_ (.Y(_2373_),
    .A(\project_audio.iter.next_ready ),
    .B(\project_audio.r_counter ));
 sg13g2_nor2_1 _5776_ (.A(_2277_),
    .B(_2373_),
    .Y(_2374_));
 sg13g2_o21ai_1 _5777_ (.B1(net690),
    .Y(_2375_),
    .A1(net452),
    .A2(_2374_));
 sg13g2_a21oi_1 _5778_ (.A1(net452),
    .A2(_2374_),
    .Y(_0430_),
    .B1(_2375_));
 sg13g2_nor2_1 _5779_ (.A(_2272_),
    .B(_2277_),
    .Y(_2376_));
 sg13g2_nand3_1 _5780_ (.B(\project_audio.iter.r[5] ),
    .C(net1155),
    .A(net1059),
    .Y(_2377_));
 sg13g2_nand4_1 _5781_ (.B(\project_audio.iter.r[2] ),
    .C(\project_audio.iter.r[1] ),
    .A(\project_audio.iter.r[3] ),
    .Y(_2378_),
    .D(\project_audio.iter.r[0] ));
 sg13g2_nand4_1 _5782_ (.B(\project_audio.iter.r[6] ),
    .C(\project_audio.iter.r[5] ),
    .A(\project_audio.iter.r[7] ),
    .Y(_2379_),
    .D(\project_audio.iter.r[4] ));
 sg13g2_nand4_1 _5783_ (.B(\project_audio.iter.r[14] ),
    .C(\project_audio.iter.r[13] ),
    .A(\project_audio.iter.r[15] ),
    .Y(_2380_),
    .D(\project_audio.iter.r[12] ));
 sg13g2_nor3_1 _5784_ (.A(_2378_),
    .B(_2379_),
    .C(_2380_),
    .Y(_2381_));
 sg13g2_nand4_1 _5785_ (.B(\project_audio.iter.r[8] ),
    .C(_2376_),
    .A(\project_audio.iter.r[9] ),
    .Y(_2382_),
    .D(_2381_));
 sg13g2_and2_1 _5786_ (.A(_2372_),
    .B(_2382_),
    .X(_2383_));
 sg13g2_nor2_1 _5787_ (.A(_0002_),
    .B(_2277_),
    .Y(_2384_));
 sg13g2_xnor2_1 _5788_ (.Y(_2385_),
    .A(_0005_),
    .B(_2384_));
 sg13g2_a22oi_1 _5789_ (.Y(_2386_),
    .B1(_2383_),
    .B2(_2385_),
    .A2(_2373_),
    .A1(net881));
 sg13g2_nor2_1 _5790_ (.A(net682),
    .B(net882),
    .Y(_0431_));
 sg13g2_o21ai_1 _5791_ (.B1(net690),
    .Y(_2387_),
    .A1(_2373_),
    .A2(_2382_));
 sg13g2_inv_2 _5792_ (.Y(_2388_),
    .A(_2387_));
 sg13g2_o21ai_1 _5793_ (.B1(_2276_),
    .Y(_2389_),
    .A1(_0002_),
    .A2(_0005_));
 sg13g2_nand2_1 _5794_ (.Y(_2390_),
    .A(net720),
    .B(_2389_));
 sg13g2_nor2_1 _5795_ (.A(_2373_),
    .B(_2390_),
    .Y(_2391_));
 sg13g2_a21oi_1 _5796_ (.A1(_2372_),
    .A2(_2389_),
    .Y(_2392_),
    .B1(net720));
 sg13g2_nor3_1 _5797_ (.A(_2387_),
    .B(_2391_),
    .C(net721),
    .Y(_0432_));
 sg13g2_o21ai_1 _5798_ (.B1(_2388_),
    .Y(_2393_),
    .A1(net485),
    .A2(_2391_));
 sg13g2_a21oi_1 _5799_ (.A1(net485),
    .A2(_2391_),
    .Y(_0433_),
    .B1(_2393_));
 sg13g2_nor3_1 _5800_ (.A(net848),
    .B(_2373_),
    .C(_2390_),
    .Y(_2394_));
 sg13g2_nor2_1 _5801_ (.A(\project_audio.iter.r[4] ),
    .B(_2394_),
    .Y(_2395_));
 sg13g2_and2_1 _5802_ (.A(net1155),
    .B(_2394_),
    .X(_2396_));
 sg13g2_nor3_1 _5803_ (.A(_2387_),
    .B(net849),
    .C(_2396_),
    .Y(_0434_));
 sg13g2_and2_1 _5804_ (.A(net1166),
    .B(_2396_),
    .X(_2397_));
 sg13g2_o21ai_1 _5805_ (.B1(_2388_),
    .Y(_2398_),
    .A1(net1166),
    .A2(_2396_));
 sg13g2_nor2_1 _5806_ (.A(_2397_),
    .B(_2398_),
    .Y(_0435_));
 sg13g2_nor3_1 _5807_ (.A(net848),
    .B(_2377_),
    .C(_2390_),
    .Y(_2399_));
 sg13g2_and2_1 _5808_ (.A(_2372_),
    .B(_2399_),
    .X(_2400_));
 sg13g2_o21ai_1 _5809_ (.B1(_2388_),
    .Y(_2401_),
    .A1(net1059),
    .A2(_2397_));
 sg13g2_nor2_1 _5810_ (.A(_2400_),
    .B(_2401_),
    .Y(_0436_));
 sg13g2_and2_1 _5811_ (.A(\project_audio.iter.r[7] ),
    .B(_2399_),
    .X(_2402_));
 sg13g2_inv_1 _5812_ (.Y(_2403_),
    .A(_2402_));
 sg13g2_a22oi_1 _5813_ (.Y(_2404_),
    .B1(_2383_),
    .B2(_2403_),
    .A2(_2373_),
    .A1(net1137));
 sg13g2_o21ai_1 _5814_ (.B1(net690),
    .Y(_2405_),
    .A1(net1137),
    .A2(_2399_));
 sg13g2_nor2_1 _5815_ (.A(_2404_),
    .B(_2405_),
    .Y(_0437_));
 sg13g2_a21oi_1 _5816_ (.A1(\project_audio.iter.r[7] ),
    .A2(_2400_),
    .Y(_2406_),
    .B1(net904));
 sg13g2_and3_1 _5817_ (.X(_2407_),
    .A(net904),
    .B(_2372_),
    .C(_2402_));
 sg13g2_nor3_1 _5818_ (.A(_2387_),
    .B(net905),
    .C(_2407_),
    .Y(_0438_));
 sg13g2_o21ai_1 _5819_ (.B1(_2388_),
    .Y(_2408_),
    .A1(net1203),
    .A2(_2407_));
 sg13g2_and2_1 _5820_ (.A(net1203),
    .B(_2407_),
    .X(_2409_));
 sg13g2_nor2_1 _5821_ (.A(_2408_),
    .B(_2409_),
    .Y(_0439_));
 sg13g2_nand2_1 _5822_ (.Y(_2410_),
    .A(\project_audio.iter.r[10] ),
    .B(\project_audio.iter.r[9] ));
 sg13g2_o21ai_1 _5823_ (.B1(_2388_),
    .Y(_2411_),
    .A1(net1152),
    .A2(_2409_));
 sg13g2_a21oi_1 _5824_ (.A1(net1152),
    .A2(_2409_),
    .Y(_0440_),
    .B1(_2411_));
 sg13g2_a21oi_1 _5825_ (.A1(\project_audio.iter.r[10] ),
    .A2(_2409_),
    .Y(_2412_),
    .B1(net1000));
 sg13g2_nor2b_2 _5826_ (.A(_2272_),
    .B_N(_2409_),
    .Y(_2413_));
 sg13g2_nor3_1 _5827_ (.A(_2387_),
    .B(net1001),
    .C(_2413_),
    .Y(_0441_));
 sg13g2_xnor2_1 _5828_ (.Y(_2414_),
    .A(net1230),
    .B(_2413_));
 sg13g2_nand2_1 _5829_ (.Y(_0442_),
    .A(_2388_),
    .B(net1231));
 sg13g2_a21oi_1 _5830_ (.A1(\project_audio.iter.r[12] ),
    .A2(_2413_),
    .Y(_2415_),
    .B1(net1150));
 sg13g2_and3_1 _5831_ (.X(_2416_),
    .A(\project_audio.iter.r[13] ),
    .B(\project_audio.iter.r[12] ),
    .C(_2413_));
 sg13g2_nor3_1 _5832_ (.A(_2387_),
    .B(net1151),
    .C(_2416_),
    .Y(_0443_));
 sg13g2_o21ai_1 _5833_ (.B1(_2388_),
    .Y(_2417_),
    .A1(net1193),
    .A2(_2416_));
 sg13g2_a21oi_1 _5834_ (.A1(net1193),
    .A2(_2416_),
    .Y(_0444_),
    .B1(_2417_));
 sg13g2_a21oi_1 _5835_ (.A1(\project_audio.iter.r[14] ),
    .A2(_2416_),
    .Y(_2418_),
    .B1(net1139));
 sg13g2_nor2b_1 _5836_ (.A(_2273_),
    .B_N(_2416_),
    .Y(_2419_));
 sg13g2_nor3_1 _5837_ (.A(_2387_),
    .B(net1140),
    .C(_2419_),
    .Y(_0445_));
 sg13g2_a21oi_1 _5838_ (.A1(_2452_),
    .A2(_2419_),
    .Y(_2420_),
    .B1(_2387_));
 sg13g2_o21ai_1 _5839_ (.B1(_2420_),
    .Y(_0446_),
    .A1(_2452_),
    .A2(_2419_));
 sg13g2_nand2_1 _5840_ (.Y(_2421_),
    .A(net1132),
    .B(_2373_));
 sg13g2_nor3_1 _5841_ (.A(_2269_),
    .B(_2273_),
    .C(_2410_),
    .Y(_2422_));
 sg13g2_nand3_1 _5842_ (.B(_2402_),
    .C(_2422_),
    .A(net904),
    .Y(_2423_));
 sg13g2_xor2_1 _5843_ (.B(_2423_),
    .A(_0004_),
    .X(_2424_));
 sg13g2_nand2_1 _5844_ (.Y(_2425_),
    .A(_2383_),
    .B(_2424_));
 sg13g2_a21oi_1 _5845_ (.A1(net1133),
    .A2(_2425_),
    .Y(_0447_),
    .B1(net682));
 sg13g2_a22oi_1 _5846_ (.Y(_2426_),
    .B1(_2281_),
    .B2(net624),
    .A2(_2271_),
    .A1(\project_audio.f_counter[0] ));
 sg13g2_nand2b_1 _5847_ (.Y(_2427_),
    .B(\project_audio.f_counter[2] ),
    .A_N(_2426_));
 sg13g2_a21oi_1 _5848_ (.A1(_2512_),
    .A2(_2271_),
    .Y(_2428_),
    .B1(_0003_));
 sg13g2_o21ai_1 _5849_ (.B1(_2428_),
    .Y(_2429_),
    .A1(_2512_),
    .A2(_2271_));
 sg13g2_xor2_1 _5850_ (.B(_2280_),
    .A(net624),
    .X(_2430_));
 sg13g2_o21ai_1 _5851_ (.B1(_2427_),
    .Y(_2431_),
    .A1(_2429_),
    .A2(_2430_));
 sg13g2_nor3_1 _5852_ (.A(net1129),
    .B(_0499_),
    .C(_2431_),
    .Y(_2432_));
 sg13g2_a21o_1 _5853_ (.A2(_2370_),
    .A1(net1129),
    .B1(_2432_),
    .X(_0448_));
 sg13g2_nand2_1 _5854_ (.Y(_2433_),
    .A(net624),
    .B(\project_audio.f_counter[0] ));
 sg13g2_nand2b_1 _5855_ (.Y(_2434_),
    .B(_2433_),
    .A_N(_2431_));
 sg13g2_a22oi_1 _5856_ (.Y(_2435_),
    .B1(_0498_),
    .B2(net1129),
    .A2(net688),
    .A1(net624));
 sg13g2_a21oi_1 _5857_ (.A1(\project_audio.iter.next_ready ),
    .A2(_2434_),
    .Y(_0449_),
    .B1(net1130));
 sg13g2_nand2_1 _5858_ (.Y(_2436_),
    .A(\project_audio.f_counter[2] ),
    .B(_2370_));
 sg13g2_a21oi_1 _5859_ (.A1(net1070),
    .A2(_2433_),
    .Y(_2437_),
    .B1(_0499_));
 sg13g2_o21ai_1 _5860_ (.B1(_2437_),
    .Y(_2438_),
    .A1(net1070),
    .A2(_2433_));
 sg13g2_o21ai_1 _5861_ (.B1(_2436_),
    .Y(_0450_),
    .A1(_2431_),
    .A2(net1071));
 sg13g2_nand2_2 _5862_ (.Y(_2439_),
    .A(_0500_),
    .B(_1372_));
 sg13g2_a21oi_1 _5863_ (.A1(_0500_),
    .A2(_1372_),
    .Y(_2440_),
    .B1(net683));
 sg13g2_nand2_1 _5864_ (.Y(_2441_),
    .A(net468),
    .B(net594));
 sg13g2_o21ai_1 _5865_ (.B1(_2441_),
    .Y(_0451_),
    .A1(_0808_),
    .A2(net596));
 sg13g2_nand2_1 _5866_ (.Y(_2442_),
    .A(net747),
    .B(net594));
 sg13g2_o21ai_1 _5867_ (.B1(_2442_),
    .Y(_0452_),
    .A1(_0837_),
    .A2(net596));
 sg13g2_nand2_1 _5868_ (.Y(_2443_),
    .A(net787),
    .B(net594));
 sg13g2_o21ai_1 _5869_ (.B1(_2443_),
    .Y(_0453_),
    .A1(_0866_),
    .A2(net596));
 sg13g2_nand2_1 _5870_ (.Y(_2444_),
    .A(net768),
    .B(net594));
 sg13g2_o21ai_1 _5871_ (.B1(_2444_),
    .Y(_0454_),
    .A1(_0892_),
    .A2(net596));
 sg13g2_nand2_1 _5872_ (.Y(_2445_),
    .A(net500),
    .B(net595));
 sg13g2_o21ai_1 _5873_ (.B1(_2445_),
    .Y(_0455_),
    .A1(_0917_),
    .A2(net596));
 sg13g2_nand2_1 _5874_ (.Y(_2446_),
    .A(net478),
    .B(net595));
 sg13g2_o21ai_1 _5875_ (.B1(_2446_),
    .Y(_0456_),
    .A1(_0935_),
    .A2(net596));
 sg13g2_nand2_1 _5876_ (.Y(_2447_),
    .A(net750),
    .B(net595));
 sg13g2_o21ai_1 _5877_ (.B1(_2447_),
    .Y(_0457_),
    .A1(_0953_),
    .A2(net596));
 sg13g2_nand2_1 _5878_ (.Y(_2448_),
    .A(net722),
    .B(net594));
 sg13g2_o21ai_1 _5879_ (.B1(_2448_),
    .Y(_0458_),
    .A1(_0964_),
    .A2(net596));
 sg13g2_nand2_1 _5880_ (.Y(_2449_),
    .A(net762),
    .B(net595));
 sg13g2_o21ai_1 _5881_ (.B1(_2449_),
    .Y(_0459_),
    .A1(_0978_),
    .A2(_2439_));
 sg13g2_nand2_1 _5882_ (.Y(_2450_),
    .A(net825),
    .B(net594));
 sg13g2_o21ai_1 _5883_ (.B1(_2450_),
    .Y(_0460_),
    .A1(_0984_),
    .A2(_2439_));
 sg13g2_nand2_1 _5884_ (.Y(_2451_),
    .A(net522),
    .B(net594));
 sg13g2_o21ai_1 _5885_ (.B1(_2451_),
    .Y(_0461_),
    .A1(_0986_),
    .A2(_2439_));
 sg13g2_and2_1 _5886_ (.A(net446),
    .B(net594),
    .X(_0462_));
 sg13g2_and2_1 _5887_ (.A(_0109_),
    .B(_1278_),
    .X(_0108_));
 sg13g2_dfrbp_1 _5888_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net297),
    .D(net1121),
    .Q_N(_2943_),
    .Q(\project_audio.iter.mult1_shift[0] ));
 sg13g2_dfrbp_1 _5889_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net267),
    .D(_0046_),
    .Q_N(_2942_),
    .Q(\project_audio.iter.mult1_shift[1] ));
 sg13g2_dfrbp_1 _5890_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net266),
    .D(_0047_),
    .Q_N(_2941_),
    .Q(\project_audio.iter.mult1_shift[2] ));
 sg13g2_dfrbp_1 _5891_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net265),
    .D(net913),
    .Q_N(_2940_),
    .Q(\project_audio.iter.mult1_shift[3] ));
 sg13g2_dfrbp_1 _5892_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net264),
    .D(net1081),
    .Q_N(_2939_),
    .Q(\project_audio.iter.mult1_shift[4] ));
 sg13g2_dfrbp_1 _5893_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net263),
    .D(net1143),
    .Q_N(_2938_),
    .Q(\project_audio.iter.mult1_shift[5] ));
 sg13g2_dfrbp_1 _5894_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net262),
    .D(net1060),
    .Q_N(_2937_),
    .Q(\project_audio.iter.mult1_shift[6] ));
 sg13g2_dfrbp_1 _5895_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net261),
    .D(net1138),
    .Q_N(_2936_),
    .Q(\project_audio.iter.mult1_shift[7] ));
 sg13g2_dfrbp_1 _5896_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net260),
    .D(net1078),
    .Q_N(_2935_),
    .Q(\project_audio.iter.mult1_shift[8] ));
 sg13g2_dfrbp_1 _5897_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net259),
    .D(net1136),
    .Q_N(_2934_),
    .Q(\project_audio.iter.mult1_shift[9] ));
 sg13g2_dfrbp_1 _5898_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net258),
    .D(net1168),
    .Q_N(_2933_),
    .Q(\project_audio.iter.mult1_shift[10] ));
 sg13g2_dfrbp_1 _5899_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net257),
    .D(net1058),
    .Q_N(_2932_),
    .Q(\project_audio.iter.mult1_shift[11] ));
 sg13g2_dfrbp_1 _5900_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net256),
    .D(net1148),
    .Q_N(_2931_),
    .Q(\project_audio.iter.mult1_shift[12] ));
 sg13g2_dfrbp_1 _5901_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net255),
    .D(_0058_),
    .Q_N(_2930_),
    .Q(\project_audio.iter.mult1_shift[13] ));
 sg13g2_dfrbp_1 _5902_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net254),
    .D(net1191),
    .Q_N(_2929_),
    .Q(\project_audio.iter.mult1_shift[14] ));
 sg13g2_dfrbp_1 _5903_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net253),
    .D(net1171),
    .Q_N(_2928_),
    .Q(\project_audio.iter.mult1_shift[15] ));
 sg13g2_dfrbp_1 _5904_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net252),
    .D(_0061_),
    .Q_N(_2927_),
    .Q(\project_audio.freq[5][0] ));
 sg13g2_dfrbp_1 _5905_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net250),
    .D(net719),
    .Q_N(_2926_),
    .Q(\project_audio.freq[5][1] ));
 sg13g2_dfrbp_1 _5906_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net248),
    .D(net755),
    .Q_N(_2925_),
    .Q(\project_audio.freq[5][2] ));
 sg13g2_dfrbp_1 _5907_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net246),
    .D(_0064_),
    .Q_N(_2924_),
    .Q(\project_audio.freq[5][3] ));
 sg13g2_dfrbp_1 _5908_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net244),
    .D(_0065_),
    .Q_N(_2923_),
    .Q(\project_audio.freq[5][4] ));
 sg13g2_dfrbp_1 _5909_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net242),
    .D(_0066_),
    .Q_N(_2922_),
    .Q(\project_audio.freq[5][5] ));
 sg13g2_dfrbp_1 _5910_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net240),
    .D(_0067_),
    .Q_N(_2921_),
    .Q(\project_audio.freq[5][6] ));
 sg13g2_dfrbp_1 _5911_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net238),
    .D(net745),
    .Q_N(_2920_),
    .Q(\project_audio.freq[5][7] ));
 sg13g2_dfrbp_1 _5912_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net236),
    .D(_0069_),
    .Q_N(_2919_),
    .Q(\project_audio.freq[5][8] ));
 sg13g2_dfrbp_1 _5913_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net234),
    .D(_0070_),
    .Q_N(_2918_),
    .Q(\project_audio.freq[5][9] ));
 sg13g2_dfrbp_1 _5914_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net232),
    .D(_0071_),
    .Q_N(_2917_),
    .Q(\project_audio.freq[5][10] ));
 sg13g2_dfrbp_1 _5915_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net230),
    .D(_0072_),
    .Q_N(_2916_),
    .Q(\project_audio.freq[5][11] ));
 sg13g2_dfrbp_1 _5916_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net228),
    .D(_0073_),
    .Q_N(_2915_),
    .Q(\project_audio.freq[6][0] ));
 sg13g2_dfrbp_1 _5917_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net226),
    .D(_0074_),
    .Q_N(_2914_),
    .Q(\project_audio.freq[6][1] ));
 sg13g2_dfrbp_1 _5918_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net224),
    .D(_0075_),
    .Q_N(_2913_),
    .Q(\project_audio.freq[6][2] ));
 sg13g2_dfrbp_1 _5919_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net222),
    .D(_0076_),
    .Q_N(_2912_),
    .Q(\project_audio.freq[6][3] ));
 sg13g2_dfrbp_1 _5920_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net220),
    .D(_0077_),
    .Q_N(_2911_),
    .Q(\project_audio.freq[6][4] ));
 sg13g2_dfrbp_1 _5921_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net218),
    .D(_0078_),
    .Q_N(_2910_),
    .Q(\project_audio.freq[6][5] ));
 sg13g2_dfrbp_1 _5922_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net216),
    .D(_0079_),
    .Q_N(_2909_),
    .Q(\project_audio.freq[6][6] ));
 sg13g2_dfrbp_1 _5923_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net214),
    .D(_0080_),
    .Q_N(_2908_),
    .Q(\project_audio.freq[6][7] ));
 sg13g2_dfrbp_1 _5924_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net212),
    .D(_0081_),
    .Q_N(_2907_),
    .Q(\project_audio.freq[6][8] ));
 sg13g2_dfrbp_1 _5925_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net210),
    .D(_0082_),
    .Q_N(_2906_),
    .Q(\project_audio.freq[6][9] ));
 sg13g2_dfrbp_1 _5926_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net208),
    .D(_0083_),
    .Q_N(_2905_),
    .Q(\project_audio.freq[6][10] ));
 sg13g2_dfrbp_1 _5927_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net206),
    .D(_0084_),
    .Q_N(_2904_),
    .Q(\project_audio.freq[6][11] ));
 sg13g2_dfrbp_1 _5928_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net204),
    .D(_0085_),
    .Q_N(_2903_),
    .Q(\project_audio.freq[7][0] ));
 sg13g2_dfrbp_1 _5929_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net202),
    .D(_0086_),
    .Q_N(_2902_),
    .Q(\project_audio.freq[7][1] ));
 sg13g2_dfrbp_1 _5930_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net200),
    .D(_0087_),
    .Q_N(_2901_),
    .Q(\project_audio.freq[7][2] ));
 sg13g2_dfrbp_1 _5931_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net198),
    .D(_0088_),
    .Q_N(_2900_),
    .Q(\project_audio.freq[7][3] ));
 sg13g2_dfrbp_1 _5932_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net196),
    .D(_0089_),
    .Q_N(_2899_),
    .Q(\project_audio.freq[7][4] ));
 sg13g2_dfrbp_1 _5933_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net194),
    .D(_0090_),
    .Q_N(_2898_),
    .Q(\project_audio.freq[7][5] ));
 sg13g2_dfrbp_1 _5934_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net192),
    .D(_0091_),
    .Q_N(_2897_),
    .Q(\project_audio.freq[7][6] ));
 sg13g2_dfrbp_1 _5935_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net190),
    .D(_0092_),
    .Q_N(_2896_),
    .Q(\project_audio.freq[7][7] ));
 sg13g2_dfrbp_1 _5936_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net188),
    .D(_0093_),
    .Q_N(_2895_),
    .Q(\project_audio.freq[7][8] ));
 sg13g2_dfrbp_1 _5937_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net186),
    .D(_0094_),
    .Q_N(_2894_),
    .Q(\project_audio.freq[7][9] ));
 sg13g2_dfrbp_1 _5938_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net184),
    .D(_0095_),
    .Q_N(_2893_),
    .Q(\project_audio.freq[7][10] ));
 sg13g2_dfrbp_1 _5939_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net182),
    .D(_0096_),
    .Q_N(_2892_),
    .Q(\project_audio.freq[7][11] ));
 sg13g2_dfrbp_1 _5940_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net180),
    .D(_0097_),
    .Q_N(_0044_),
    .Q(\hpos[0] ));
 sg13g2_dfrbp_1 _5941_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net179),
    .D(net1210),
    .Q_N(_0007_),
    .Q(\hpos[1] ));
 sg13g2_dfrbp_1 _5942_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net178),
    .D(_0099_),
    .Q_N(_0008_),
    .Q(\hpos[2] ));
 sg13g2_dfrbp_1 _5943_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net177),
    .D(_0100_),
    .Q_N(_0009_),
    .Q(\hpos[3] ));
 sg13g2_dfrbp_1 _5944_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net176),
    .D(_0101_),
    .Q_N(_0010_),
    .Q(\hpos[4] ));
 sg13g2_dfrbp_1 _5945_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net175),
    .D(_0102_),
    .Q_N(_0011_),
    .Q(\hpos[5] ));
 sg13g2_dfrbp_1 _5946_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net174),
    .D(net822),
    .Q_N(_0012_),
    .Q(\hpos[6] ));
 sg13g2_dfrbp_1 _5947_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net173),
    .D(_0104_),
    .Q_N(_0013_),
    .Q(\hpos[7] ));
 sg13g2_dfrbp_1 _5948_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net172),
    .D(_0105_),
    .Q_N(_0023_),
    .Q(\hpos[8] ));
 sg13g2_dfrbp_1 _5949_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net171),
    .D(_0106_),
    .Q_N(_2891_),
    .Q(\hpos[9] ));
 sg13g2_dfrbp_1 _5950_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net170),
    .D(_0107_),
    .Q_N(_2890_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _5951_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net169),
    .D(_0108_),
    .Q_N(_2889_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _5952_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net168),
    .D(_0109_),
    .Q_N(_2888_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _5953_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net167),
    .D(_0110_),
    .Q_N(_2887_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _5954_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net166),
    .D(net440),
    .Q_N(_0043_),
    .Q(\frame_no[0] ));
 sg13g2_dfrbp_1 _5955_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net164),
    .D(_0112_),
    .Q_N(_2886_),
    .Q(\frame_no[1] ));
 sg13g2_dfrbp_1 _5956_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net162),
    .D(net1237),
    .Q_N(_0014_),
    .Q(\frame_no[2] ));
 sg13g2_dfrbp_1 _5957_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net160),
    .D(net1207),
    .Q_N(_0015_),
    .Q(\frame_no[3] ));
 sg13g2_dfrbp_1 _5958_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net158),
    .D(_0115_),
    .Q_N(_0017_),
    .Q(\frame_no[4] ));
 sg13g2_dfrbp_1 _5959_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net156),
    .D(net1233),
    .Q_N(_0016_),
    .Q(\frame_no[5] ));
 sg13g2_dfrbp_1 _5960_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net154),
    .D(_0117_),
    .Q_N(_0018_),
    .Q(\frame_no[6] ));
 sg13g2_dfrbp_1 _5961_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net152),
    .D(net1123),
    .Q_N(_0019_),
    .Q(\frame_no[7] ));
 sg13g2_dfrbp_1 _5962_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net150),
    .D(net458),
    .Q_N(_0020_),
    .Q(\frame_no[8] ));
 sg13g2_dfrbp_1 _5963_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net148),
    .D(_0120_),
    .Q_N(_2885_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _5964_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net147),
    .D(_0121_),
    .Q_N(_2884_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _5965_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net146),
    .D(net1197),
    .Q_N(_2883_),
    .Q(\sync_gen.vpos[0] ));
 sg13g2_dfrbp_1 _5966_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net144),
    .D(_0123_),
    .Q_N(_2882_),
    .Q(\sync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _5967_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net142),
    .D(_0124_),
    .Q_N(_2881_),
    .Q(\sync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _5968_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net140),
    .D(_0125_),
    .Q_N(_2880_),
    .Q(\sync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _5969_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net138),
    .D(_0126_),
    .Q_N(_2879_),
    .Q(\sync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _5970_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net136),
    .D(_0127_),
    .Q_N(_0022_),
    .Q(\sync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _5971_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net134),
    .D(_0128_),
    .Q_N(_2878_),
    .Q(\sync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _5972_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net132),
    .D(_0129_),
    .Q_N(_2877_),
    .Q(\sync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _5973_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net130),
    .D(_0130_),
    .Q_N(_2876_),
    .Q(\sync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _5974_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net128),
    .D(_0131_),
    .Q_N(_2875_),
    .Q(\sync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _5975_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net126),
    .D(net1164),
    .Q_N(_2874_),
    .Q(hsync));
 sg13g2_dfrbp_1 _5976_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net125),
    .D(net1227),
    .Q_N(_2873_),
    .Q(\sync_gen.vsync ));
 sg13g2_dfrbp_1 _5977_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net124),
    .D(net436),
    .Q_N(_0042_),
    .Q(\project_audio.nco_increment_gen.counter[0] ));
 sg13g2_dfrbp_1 _5978_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net123),
    .D(net964),
    .Q_N(_2872_),
    .Q(\project_audio.nco_increment_gen.counter[1] ));
 sg13g2_dfrbp_1 _5979_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net122),
    .D(net466),
    .Q_N(_2871_),
    .Q(\project_audio.nco_increment_gen.counter[2] ));
 sg13g2_dfrbp_1 _5980_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net121),
    .D(net753),
    .Q_N(_2870_),
    .Q(\project_audio.nco_increment_gen.counter[3] ));
 sg13g2_dfrbp_1 _5981_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net120),
    .D(net791),
    .Q_N(_2869_),
    .Q(\project_audio.nco_increment_gen.counter[4] ));
 sg13g2_dfrbp_1 _5982_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net119),
    .D(_0139_),
    .Q_N(_2868_),
    .Q(\project_audio.nco_increment_gen.counter[5] ));
 sg13g2_dfrbp_1 _5983_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net118),
    .D(net783),
    .Q_N(_2867_),
    .Q(\project_audio.nco_increment_gen.counter[6] ));
 sg13g2_dfrbp_1 _5984_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net117),
    .D(net461),
    .Q_N(_2866_),
    .Q(\project_audio.nco_increment_gen.counter[7] ));
 sg13g2_dfrbp_1 _5985_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net116),
    .D(net828),
    .Q_N(_0024_),
    .Q(\project_audio.nco_increment_gen.counter[8] ));
 sg13g2_dfrbp_1 _5986_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net115),
    .D(_0143_),
    .Q_N(_2865_),
    .Q(\project_audio.freq[4][0] ));
 sg13g2_dfrbp_1 _5987_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net113),
    .D(_0144_),
    .Q_N(_2864_),
    .Q(\project_audio.freq[4][1] ));
 sg13g2_dfrbp_1 _5988_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net111),
    .D(net519),
    .Q_N(_2863_),
    .Q(\project_audio.freq[4][2] ));
 sg13g2_dfrbp_1 _5989_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net109),
    .D(net797),
    .Q_N(_2862_),
    .Q(\project_audio.freq[4][3] ));
 sg13g2_dfrbp_1 _5990_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net107),
    .D(net521),
    .Q_N(_2861_),
    .Q(\project_audio.freq[4][4] ));
 sg13g2_dfrbp_1 _5991_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net105),
    .D(_0148_),
    .Q_N(_2860_),
    .Q(\project_audio.freq[4][5] ));
 sg13g2_dfrbp_1 _5992_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net103),
    .D(_0149_),
    .Q_N(_2859_),
    .Q(\project_audio.freq[4][6] ));
 sg13g2_dfrbp_1 _5993_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net101),
    .D(_0150_),
    .Q_N(_2858_),
    .Q(\project_audio.freq[4][7] ));
 sg13g2_dfrbp_1 _5994_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net99),
    .D(_0151_),
    .Q_N(_2857_),
    .Q(\project_audio.freq[4][8] ));
 sg13g2_dfrbp_1 _5995_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net97),
    .D(_0152_),
    .Q_N(_2856_),
    .Q(\project_audio.freq[4][9] ));
 sg13g2_dfrbp_1 _5996_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net95),
    .D(_0153_),
    .Q_N(_2855_),
    .Q(\project_audio.freq[4][10] ));
 sg13g2_dfrbp_1 _5997_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net93),
    .D(_0154_),
    .Q_N(_2854_),
    .Q(\project_audio.freq[4][11] ));
 sg13g2_dfrbp_1 _5998_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net91),
    .D(_0155_),
    .Q_N(_2853_),
    .Q(prev_vsync));
 sg13g2_dfrbp_1 _5999_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net90),
    .D(net471),
    .Q_N(_2852_),
    .Q(\project_audio.freq[3][0] ));
 sg13g2_dfrbp_1 _6000_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net88),
    .D(net502),
    .Q_N(_2851_),
    .Q(\project_audio.freq[3][1] ));
 sg13g2_dfrbp_1 _6001_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net86),
    .D(net726),
    .Q_N(_2850_),
    .Q(\project_audio.freq[3][2] ));
 sg13g2_dfrbp_1 _6002_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net84),
    .D(_0159_),
    .Q_N(_2849_),
    .Q(\project_audio.freq[3][3] ));
 sg13g2_dfrbp_1 _6003_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net82),
    .D(_0160_),
    .Q_N(_2848_),
    .Q(\project_audio.freq[3][4] ));
 sg13g2_dfrbp_1 _6004_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net80),
    .D(_0161_),
    .Q_N(_2847_),
    .Q(\project_audio.freq[3][5] ));
 sg13g2_dfrbp_1 _6005_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net78),
    .D(_0162_),
    .Q_N(_2846_),
    .Q(\project_audio.freq[3][6] ));
 sg13g2_dfrbp_1 _6006_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net76),
    .D(_0163_),
    .Q_N(_2845_),
    .Q(\project_audio.freq[3][7] ));
 sg13g2_dfrbp_1 _6007_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net74),
    .D(_0164_),
    .Q_N(_2844_),
    .Q(\project_audio.freq[3][8] ));
 sg13g2_dfrbp_1 _6008_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net72),
    .D(_0165_),
    .Q_N(_2843_),
    .Q(\project_audio.freq[3][9] ));
 sg13g2_dfrbp_1 _6009_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net70),
    .D(_0166_),
    .Q_N(_2842_),
    .Q(\project_audio.freq[3][10] ));
 sg13g2_dfrbp_1 _6010_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net68),
    .D(_0167_),
    .Q_N(_2841_),
    .Q(\project_audio.freq[3][11] ));
 sg13g2_dfrbp_1 _6011_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net66),
    .D(_0168_),
    .Q_N(_2840_),
    .Q(\project_audio.freq[0][0] ));
 sg13g2_dfrbp_1 _6012_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net64),
    .D(_0169_),
    .Q_N(_2839_),
    .Q(\project_audio.freq[0][1] ));
 sg13g2_dfrbp_1 _6013_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net62),
    .D(_0170_),
    .Q_N(_2838_),
    .Q(\project_audio.freq[0][2] ));
 sg13g2_dfrbp_1 _6014_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net60),
    .D(_0171_),
    .Q_N(_2837_),
    .Q(\project_audio.freq[0][3] ));
 sg13g2_dfrbp_1 _6015_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net58),
    .D(_0172_),
    .Q_N(_2836_),
    .Q(\project_audio.freq[0][4] ));
 sg13g2_dfrbp_1 _6016_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net56),
    .D(_0173_),
    .Q_N(_2835_),
    .Q(\project_audio.freq[0][5] ));
 sg13g2_dfrbp_1 _6017_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net54),
    .D(_0174_),
    .Q_N(_2834_),
    .Q(\project_audio.freq[0][6] ));
 sg13g2_dfrbp_1 _6018_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net52),
    .D(_0175_),
    .Q_N(_2833_),
    .Q(\project_audio.freq[0][7] ));
 sg13g2_dfrbp_1 _6019_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net50),
    .D(_0176_),
    .Q_N(_2832_),
    .Q(\project_audio.freq[0][8] ));
 sg13g2_dfrbp_1 _6020_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net48),
    .D(_0177_),
    .Q_N(_2831_),
    .Q(\project_audio.freq[0][9] ));
 sg13g2_dfrbp_1 _6021_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net46),
    .D(_0178_),
    .Q_N(_2830_),
    .Q(\project_audio.freq[0][10] ));
 sg13g2_dfrbp_1 _6022_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net44),
    .D(_0179_),
    .Q_N(_2829_),
    .Q(\project_audio.freq[0][11] ));
 sg13g2_dfrbp_1 _6023_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net42),
    .D(_0180_),
    .Q_N(_2828_),
    .Q(\project_audio.freq[2][0] ));
 sg13g2_dfrbp_1 _6024_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net40),
    .D(_0181_),
    .Q_N(_2827_),
    .Q(\project_audio.freq[2][1] ));
 sg13g2_dfrbp_1 _6025_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net38),
    .D(_0182_),
    .Q_N(_2826_),
    .Q(\project_audio.freq[2][2] ));
 sg13g2_dfrbp_1 _6026_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net36),
    .D(_0183_),
    .Q_N(_2825_),
    .Q(\project_audio.freq[2][3] ));
 sg13g2_dfrbp_1 _6027_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net34),
    .D(_0184_),
    .Q_N(_2824_),
    .Q(\project_audio.freq[2][4] ));
 sg13g2_dfrbp_1 _6028_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net32),
    .D(_0185_),
    .Q_N(_2823_),
    .Q(\project_audio.freq[2][5] ));
 sg13g2_dfrbp_1 _6029_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net30),
    .D(_0186_),
    .Q_N(_2822_),
    .Q(\project_audio.freq[2][6] ));
 sg13g2_dfrbp_1 _6030_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net28),
    .D(_0187_),
    .Q_N(_2821_),
    .Q(\project_audio.freq[2][7] ));
 sg13g2_dfrbp_1 _6031_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net26),
    .D(_0188_),
    .Q_N(_2820_),
    .Q(\project_audio.freq[2][8] ));
 sg13g2_dfrbp_1 _6032_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net24),
    .D(_0189_),
    .Q_N(_2819_),
    .Q(\project_audio.freq[2][9] ));
 sg13g2_dfrbp_1 _6033_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net22),
    .D(_0190_),
    .Q_N(_2818_),
    .Q(\project_audio.freq[2][10] ));
 sg13g2_dfrbp_1 _6034_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net20),
    .D(_0191_),
    .Q_N(_2817_),
    .Q(\project_audio.freq[2][11] ));
 sg13g2_dfrbp_1 _6035_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net18),
    .D(_0192_),
    .Q_N(_2816_),
    .Q(\project_audio.iter.mult1_shift[18] ));
 sg13g2_dfrbp_1 _6036_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net16),
    .D(_0193_),
    .Q_N(_2815_),
    .Q(\project_audio.iter.mult1_shift[19] ));
 sg13g2_dfrbp_1 _6037_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net432),
    .D(net888),
    .Q_N(_2814_),
    .Q(\project_audio.iter.mult1_shift[20] ));
 sg13g2_dfrbp_1 _6038_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net430),
    .D(_0195_),
    .Q_N(_2813_),
    .Q(\project_audio.iter.mult1_shift[21] ));
 sg13g2_dfrbp_1 _6039_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net428),
    .D(_0196_),
    .Q_N(_2812_),
    .Q(\project_audio.iter.mult1_shift[22] ));
 sg13g2_dfrbp_1 _6040_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net426),
    .D(_0197_),
    .Q_N(_2811_),
    .Q(\project_audio.iter.mult1_shift[23] ));
 sg13g2_dfrbp_1 _6041_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net424),
    .D(net820),
    .Q_N(_2810_),
    .Q(\project_audio.iter.mult1_shift[24] ));
 sg13g2_dfrbp_1 _6042_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net422),
    .D(net853),
    .Q_N(_2809_),
    .Q(\project_audio.iter.mult1_shift[25] ));
 sg13g2_dfrbp_1 _6043_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net420),
    .D(_0200_),
    .Q_N(_2808_),
    .Q(\project_audio.iter.mult1_shift[26] ));
 sg13g2_dfrbp_1 _6044_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net418),
    .D(net868),
    .Q_N(_2807_),
    .Q(\project_audio.iter.mult1_shift[27] ));
 sg13g2_dfrbp_1 _6045_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net416),
    .D(_0202_),
    .Q_N(_2806_),
    .Q(\project_audio.iter.mult1_shift[28] ));
 sg13g2_dfrbp_1 _6046_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net414),
    .D(net801),
    .Q_N(_2805_),
    .Q(\project_audio.iter.mult1_shift[29] ));
 sg13g2_dfrbp_1 _6047_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net412),
    .D(net1056),
    .Q_N(_2804_),
    .Q(\project_audio.iter.mult1_shift[30] ));
 sg13g2_dfrbp_1 _6048_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net410),
    .D(net761),
    .Q_N(_2803_),
    .Q(\project_audio.iter.mult1_shift[31] ));
 sg13g2_dfrbp_1 _6049_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net408),
    .D(net805),
    .Q_N(_2802_),
    .Q(\project_audio.iter.mult_accum[0] ));
 sg13g2_dfrbp_1 _6050_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net406),
    .D(net780),
    .Q_N(_2801_),
    .Q(\project_audio.iter.mult_accum[1] ));
 sg13g2_dfrbp_1 _6051_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net404),
    .D(net809),
    .Q_N(_2800_),
    .Q(\project_audio.iter.mult_accum[2] ));
 sg13g2_dfrbp_1 _6052_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net402),
    .D(_0209_),
    .Q_N(_2799_),
    .Q(\project_audio.iter.mult_accum[3] ));
 sg13g2_dfrbp_1 _6053_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net400),
    .D(_0210_),
    .Q_N(_2798_),
    .Q(\project_audio.iter.mult_accum[4] ));
 sg13g2_dfrbp_1 _6054_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net398),
    .D(net840),
    .Q_N(_2797_),
    .Q(\project_audio.iter.mult_accum[5] ));
 sg13g2_dfrbp_1 _6055_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net396),
    .D(_0212_),
    .Q_N(_2796_),
    .Q(\project_audio.iter.mult_accum[6] ));
 sg13g2_dfrbp_1 _6056_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net394),
    .D(net739),
    .Q_N(_2795_),
    .Q(\project_audio.iter.mult_accum[7] ));
 sg13g2_dfrbp_1 _6057_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net392),
    .D(_0214_),
    .Q_N(_2794_),
    .Q(\project_audio.iter.mult_accum[8] ));
 sg13g2_dfrbp_1 _6058_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net390),
    .D(net942),
    .Q_N(_2793_),
    .Q(\project_audio.iter.mult_accum[9] ));
 sg13g2_dfrbp_1 _6059_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net388),
    .D(_0216_),
    .Q_N(_2792_),
    .Q(\project_audio.iter.mult_accum[10] ));
 sg13g2_dfrbp_1 _6060_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net386),
    .D(_0217_),
    .Q_N(_2791_),
    .Q(\project_audio.iter.mult_accum[11] ));
 sg13g2_dfrbp_1 _6061_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net384),
    .D(_0218_),
    .Q_N(_2790_),
    .Q(\project_audio.iter.mult_accum[12] ));
 sg13g2_dfrbp_1 _6062_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net382),
    .D(_0219_),
    .Q_N(_2789_),
    .Q(\project_audio.iter.mult_accum[13] ));
 sg13g2_dfrbp_1 _6063_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net380),
    .D(_0220_),
    .Q_N(_2788_),
    .Q(\project_audio.iter.mult_accum[14] ));
 sg13g2_dfrbp_1 _6064_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net378),
    .D(net771),
    .Q_N(_2787_),
    .Q(\project_audio.iter.mult_accum[15] ));
 sg13g2_dfrbp_1 _6065_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net376),
    .D(_0222_),
    .Q_N(_2786_),
    .Q(\project_audio.iter.mult_accum[16] ));
 sg13g2_dfrbp_1 _6066_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net374),
    .D(_0223_),
    .Q_N(_2785_),
    .Q(\project_audio.iter.mult_accum[17] ));
 sg13g2_dfrbp_1 _6067_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net372),
    .D(_0224_),
    .Q_N(_2784_),
    .Q(\project_audio.iter.mult_accum[18] ));
 sg13g2_dfrbp_1 _6068_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net370),
    .D(_0225_),
    .Q_N(_2783_),
    .Q(\project_audio.iter.mult_accum[19] ));
 sg13g2_dfrbp_1 _6069_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net368),
    .D(_0226_),
    .Q_N(_2782_),
    .Q(\project_audio.iter.mult_accum[20] ));
 sg13g2_dfrbp_1 _6070_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net366),
    .D(_0227_),
    .Q_N(_2781_),
    .Q(\project_audio.iter.mult_accum[21] ));
 sg13g2_dfrbp_1 _6071_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net364),
    .D(_0228_),
    .Q_N(_2780_),
    .Q(\project_audio.iter.mult_accum[22] ));
 sg13g2_dfrbp_1 _6072_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net362),
    .D(_0229_),
    .Q_N(_2779_),
    .Q(\project_audio.iter.mult_accum[23] ));
 sg13g2_dfrbp_1 _6073_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net360),
    .D(_0230_),
    .Q_N(_2778_),
    .Q(\project_audio.iter.mult_accum[24] ));
 sg13g2_dfrbp_1 _6074_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net358),
    .D(_0231_),
    .Q_N(_2777_),
    .Q(\project_audio.iter.mult_accum[25] ));
 sg13g2_dfrbp_1 _6075_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net356),
    .D(_0232_),
    .Q_N(_2776_),
    .Q(\project_audio.iter.mult_accum[26] ));
 sg13g2_dfrbp_1 _6076_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net354),
    .D(_0233_),
    .Q_N(_2775_),
    .Q(\project_audio.iter.mult_accum[27] ));
 sg13g2_dfrbp_1 _6077_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net352),
    .D(_0234_),
    .Q_N(_2774_),
    .Q(\project_audio.iter.mult_accum[28] ));
 sg13g2_dfrbp_1 _6078_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net350),
    .D(net1107),
    .Q_N(_2773_),
    .Q(\project_audio.iter.mult_accum[29] ));
 sg13g2_dfrbp_1 _6079_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net348),
    .D(net950),
    .Q_N(_2772_),
    .Q(\project_audio.iter.mult_accum[30] ));
 sg13g2_dfrbp_1 _6080_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net346),
    .D(_0237_),
    .Q_N(_2771_),
    .Q(\project_audio.iter.mult_accum[31] ));
 sg13g2_dfrbp_1 _6081_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net344),
    .D(_0238_),
    .Q_N(_2770_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.snd ));
 sg13g2_dfrbp_1 _6082_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net342),
    .D(_0239_),
    .Q_N(_2769_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[0] ));
 sg13g2_dfrbp_1 _6083_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net340),
    .D(_0240_),
    .Q_N(_2768_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[1] ));
 sg13g2_dfrbp_1 _6084_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net338),
    .D(net982),
    .Q_N(_2767_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[2] ));
 sg13g2_dfrbp_1 _6085_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net336),
    .D(net1041),
    .Q_N(_2766_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[3] ));
 sg13g2_dfrbp_1 _6086_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net334),
    .D(net1069),
    .Q_N(_2765_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[4] ));
 sg13g2_dfrbp_1 _6087_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net332),
    .D(net1175),
    .Q_N(_2764_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[5] ));
 sg13g2_dfrbp_1 _6088_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net330),
    .D(net1116),
    .Q_N(_2763_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[6] ));
 sg13g2_dfrbp_1 _6089_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net328),
    .D(net990),
    .Q_N(_2762_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[7] ));
 sg13g2_dfrbp_1 _6090_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net326),
    .D(_0247_),
    .Q_N(_2761_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[8] ));
 sg13g2_dfrbp_1 _6091_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net324),
    .D(_0248_),
    .Q_N(_2760_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[9] ));
 sg13g2_dfrbp_1 _6092_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net322),
    .D(net1018),
    .Q_N(_2759_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[10] ));
 sg13g2_dfrbp_1 _6093_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net320),
    .D(net970),
    .Q_N(_2758_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[11] ));
 sg13g2_dfrbp_1 _6094_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net318),
    .D(_0251_),
    .Q_N(_2757_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[12] ));
 sg13g2_dfrbp_1 _6095_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net316),
    .D(_0252_),
    .Q_N(_2756_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[13] ));
 sg13g2_dfrbp_1 _6096_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net314),
    .D(_0253_),
    .Q_N(_2755_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[14] ));
 sg13g2_dfrbp_1 _6097_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net312),
    .D(net536),
    .Q_N(_2754_),
    .Q(\project_audio.genblk1[7].n_c_oh_my.phase[15] ));
 sg13g2_dfrbp_1 _6098_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net310),
    .D(_0255_),
    .Q_N(_2753_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.snd ));
 sg13g2_dfrbp_1 _6099_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net308),
    .D(_0256_),
    .Q_N(_2752_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[0] ));
 sg13g2_dfrbp_1 _6100_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net306),
    .D(_0257_),
    .Q_N(_2751_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[1] ));
 sg13g2_dfrbp_1 _6101_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net304),
    .D(net1093),
    .Q_N(_2750_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[2] ));
 sg13g2_dfrbp_1 _6102_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net302),
    .D(net1103),
    .Q_N(_2749_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[3] ));
 sg13g2_dfrbp_1 _6103_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net300),
    .D(net1089),
    .Q_N(_2748_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[4] ));
 sg13g2_dfrbp_1 _6104_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net298),
    .D(_0261_),
    .Q_N(_2747_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[5] ));
 sg13g2_dfrbp_1 _6105_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net296),
    .D(net1145),
    .Q_N(_2746_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[6] ));
 sg13g2_dfrbp_1 _6106_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net294),
    .D(net1113),
    .Q_N(_2745_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[7] ));
 sg13g2_dfrbp_1 _6107_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net292),
    .D(_0264_),
    .Q_N(_2744_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[8] ));
 sg13g2_dfrbp_1 _6108_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net290),
    .D(_0265_),
    .Q_N(_2743_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[9] ));
 sg13g2_dfrbp_1 _6109_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net288),
    .D(net974),
    .Q_N(_2742_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[10] ));
 sg13g2_dfrbp_1 _6110_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net286),
    .D(net926),
    .Q_N(_2741_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[11] ));
 sg13g2_dfrbp_1 _6111_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net284),
    .D(_0268_),
    .Q_N(_2740_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[12] ));
 sg13g2_dfrbp_1 _6112_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net282),
    .D(net504),
    .Q_N(_2739_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[13] ));
 sg13g2_dfrbp_1 _6113_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net280),
    .D(_0270_),
    .Q_N(_2738_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[14] ));
 sg13g2_dfrbp_1 _6114_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net278),
    .D(net531),
    .Q_N(_2737_),
    .Q(\project_audio.genblk1[6].n_c_oh_my.phase[15] ));
 sg13g2_dfrbp_1 _6115_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net276),
    .D(_0272_),
    .Q_N(_2736_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.snd ));
 sg13g2_dfrbp_1 _6116_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net274),
    .D(_0273_),
    .Q_N(_2735_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[0] ));
 sg13g2_dfrbp_1 _6117_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net272),
    .D(_0274_),
    .Q_N(_2734_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[1] ));
 sg13g2_dfrbp_1 _6118_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net270),
    .D(net976),
    .Q_N(_2733_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[2] ));
 sg13g2_dfrbp_1 _6119_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net268),
    .D(net1020),
    .Q_N(_2732_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[3] ));
 sg13g2_dfrbp_1 _6120_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net249),
    .D(net1028),
    .Q_N(_2731_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[4] ));
 sg13g2_dfrbp_1 _6121_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net245),
    .D(_0278_),
    .Q_N(_2730_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[5] ));
 sg13g2_dfrbp_1 _6122_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net241),
    .D(_0279_),
    .Q_N(_2729_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[6] ));
 sg13g2_dfrbp_1 _6123_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net237),
    .D(net1095),
    .Q_N(_2728_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[7] ));
 sg13g2_dfrbp_1 _6124_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net233),
    .D(net956),
    .Q_N(_2727_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[8] ));
 sg13g2_dfrbp_1 _6125_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net229),
    .D(_0282_),
    .Q_N(_2726_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[9] ));
 sg13g2_dfrbp_1 _6126_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net225),
    .D(net1039),
    .Q_N(_2725_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[10] ));
 sg13g2_dfrbp_1 _6127_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net221),
    .D(net1064),
    .Q_N(_2724_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[11] ));
 sg13g2_dfrbp_1 _6128_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net217),
    .D(_0285_),
    .Q_N(_2723_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[12] ));
 sg13g2_dfrbp_1 _6129_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net213),
    .D(_0286_),
    .Q_N(_2722_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[13] ));
 sg13g2_dfrbp_1 _6130_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net209),
    .D(_0287_),
    .Q_N(_2721_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[14] ));
 sg13g2_dfrbp_1 _6131_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net205),
    .D(net495),
    .Q_N(_2720_),
    .Q(\project_audio.genblk1[5].n_c_oh_my.phase[15] ));
 sg13g2_dfrbp_1 _6132_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net201),
    .D(_0289_),
    .Q_N(_2719_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.snd ));
 sg13g2_dfrbp_1 _6133_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net197),
    .D(_0290_),
    .Q_N(_2718_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[0] ));
 sg13g2_dfrbp_1 _6134_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net193),
    .D(_0291_),
    .Q_N(_2717_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[1] ));
 sg13g2_dfrbp_1 _6135_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net189),
    .D(net988),
    .Q_N(_2716_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[2] ));
 sg13g2_dfrbp_1 _6136_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net185),
    .D(_0293_),
    .Q_N(_2715_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[3] ));
 sg13g2_dfrbp_1 _6137_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net181),
    .D(net1035),
    .Q_N(_2714_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[4] ));
 sg13g2_dfrbp_1 _6138_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net163),
    .D(_0295_),
    .Q_N(_2713_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[5] ));
 sg13g2_dfrbp_1 _6139_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net159),
    .D(_0296_),
    .Q_N(_2712_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[6] ));
 sg13g2_dfrbp_1 _6140_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net155),
    .D(_0297_),
    .Q_N(_2711_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[7] ));
 sg13g2_dfrbp_1 _6141_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net151),
    .D(net996),
    .Q_N(_2710_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[8] ));
 sg13g2_dfrbp_1 _6142_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net145),
    .D(_0299_),
    .Q_N(_2709_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[9] ));
 sg13g2_dfrbp_1 _6143_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net141),
    .D(net1085),
    .Q_N(_2708_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[10] ));
 sg13g2_dfrbp_1 _6144_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net137),
    .D(net940),
    .Q_N(_2707_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[11] ));
 sg13g2_dfrbp_1 _6145_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net133),
    .D(_0302_),
    .Q_N(_2706_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[12] ));
 sg13g2_dfrbp_1 _6146_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net129),
    .D(net488),
    .Q_N(_2705_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[13] ));
 sg13g2_dfrbp_1 _6147_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net114),
    .D(_0304_),
    .Q_N(_2704_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[14] ));
 sg13g2_dfrbp_1 _6148_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net110),
    .D(net493),
    .Q_N(_2703_),
    .Q(\project_audio.genblk1[4].n_c_oh_my.phase[15] ));
 sg13g2_dfrbp_1 _6149_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net106),
    .D(_0306_),
    .Q_N(_2702_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.snd ));
 sg13g2_dfrbp_1 _6150_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net102),
    .D(_0307_),
    .Q_N(_2701_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[0] ));
 sg13g2_dfrbp_1 _6151_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net98),
    .D(_0308_),
    .Q_N(_2700_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[1] ));
 sg13g2_dfrbp_1 _6152_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net94),
    .D(net1032),
    .Q_N(_2699_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[2] ));
 sg13g2_dfrbp_1 _6153_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net89),
    .D(_0310_),
    .Q_N(_2698_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[3] ));
 sg13g2_dfrbp_1 _6154_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net85),
    .D(net1044),
    .Q_N(_2697_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[4] ));
 sg13g2_dfrbp_1 _6155_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net81),
    .D(_0312_),
    .Q_N(_2696_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[5] ));
 sg13g2_dfrbp_1 _6156_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net77),
    .D(net1026),
    .Q_N(_2695_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[6] ));
 sg13g2_dfrbp_1 _6157_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net73),
    .D(_0314_),
    .Q_N(_2694_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[7] ));
 sg13g2_dfrbp_1 _6158_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net69),
    .D(net1016),
    .Q_N(_2693_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[8] ));
 sg13g2_dfrbp_1 _6159_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net65),
    .D(_0316_),
    .Q_N(_2692_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[9] ));
 sg13g2_dfrbp_1 _6160_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net61),
    .D(net1009),
    .Q_N(_2691_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[10] ));
 sg13g2_dfrbp_1 _6161_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net57),
    .D(net947),
    .Q_N(_2690_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[11] ));
 sg13g2_dfrbp_1 _6162_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net53),
    .D(_0319_),
    .Q_N(_2689_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[12] ));
 sg13g2_dfrbp_1 _6163_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net49),
    .D(net481),
    .Q_N(_2688_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[13] ));
 sg13g2_dfrbp_1 _6164_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net45),
    .D(_0321_),
    .Q_N(_2687_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[14] ));
 sg13g2_dfrbp_1 _6165_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net41),
    .D(net526),
    .Q_N(_2686_),
    .Q(\project_audio.genblk1[3].n_c_oh_my.phase[15] ));
 sg13g2_dfrbp_1 _6166_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net37),
    .D(_0323_),
    .Q_N(_2685_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.snd ));
 sg13g2_dfrbp_1 _6167_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net33),
    .D(_0324_),
    .Q_N(_2684_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[0] ));
 sg13g2_dfrbp_1 _6168_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net29),
    .D(_0325_),
    .Q_N(_2683_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[1] ));
 sg13g2_dfrbp_1 _6169_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net25),
    .D(net1101),
    .Q_N(_2682_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[2] ));
 sg13g2_dfrbp_1 _6170_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net21),
    .D(_0327_),
    .Q_N(_2681_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[3] ));
 sg13g2_dfrbp_1 _6171_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net17),
    .D(net1004),
    .Q_N(_2680_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[4] ));
 sg13g2_dfrbp_1 _6172_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net431),
    .D(_0329_),
    .Q_N(_2679_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[5] ));
 sg13g2_dfrbp_1 _6173_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net427),
    .D(net1111),
    .Q_N(_2678_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[6] ));
 sg13g2_dfrbp_1 _6174_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net423),
    .D(_0331_),
    .Q_N(_2677_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[7] ));
 sg13g2_dfrbp_1 _6175_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net419),
    .D(net998),
    .Q_N(_2676_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[8] ));
 sg13g2_dfrbp_1 _6176_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net415),
    .D(net1154),
    .Q_N(_2675_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[9] ));
 sg13g2_dfrbp_1 _6177_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net411),
    .D(net979),
    .Q_N(_2674_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[10] ));
 sg13g2_dfrbp_1 _6178_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net407),
    .D(net954),
    .Q_N(_2673_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[11] ));
 sg13g2_dfrbp_1 _6179_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net403),
    .D(_0336_),
    .Q_N(_2672_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[12] ));
 sg13g2_dfrbp_1 _6180_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net399),
    .D(net477),
    .Q_N(_2671_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[13] ));
 sg13g2_dfrbp_1 _6181_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net395),
    .D(_0338_),
    .Q_N(_2670_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[14] ));
 sg13g2_dfrbp_1 _6182_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net391),
    .D(net512),
    .Q_N(_2669_),
    .Q(\project_audio.genblk1[2].n_c_oh_my.phase[15] ));
 sg13g2_dfrbp_1 _6183_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net387),
    .D(_0340_),
    .Q_N(_2668_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.snd ));
 sg13g2_dfrbp_1 _6184_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net383),
    .D(_0341_),
    .Q_N(_2667_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[0] ));
 sg13g2_dfrbp_1 _6185_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net379),
    .D(net1022),
    .Q_N(_2666_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[1] ));
 sg13g2_dfrbp_1 _6186_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net375),
    .D(net986),
    .Q_N(_2665_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[2] ));
 sg13g2_dfrbp_1 _6187_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net371),
    .D(_0344_),
    .Q_N(_2664_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[3] ));
 sg13g2_dfrbp_1 _6188_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net367),
    .D(net1109),
    .Q_N(_2663_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[4] ));
 sg13g2_dfrbp_1 _6189_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net363),
    .D(_0346_),
    .Q_N(_2662_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[5] ));
 sg13g2_dfrbp_1 _6190_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net359),
    .D(net1013),
    .Q_N(_2661_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[6] ));
 sg13g2_dfrbp_1 _6191_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net355),
    .D(net1011),
    .Q_N(_2660_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[7] ));
 sg13g2_dfrbp_1 _6192_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net351),
    .D(net984),
    .Q_N(_2659_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[8] ));
 sg13g2_dfrbp_1 _6193_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net347),
    .D(net1179),
    .Q_N(_2658_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[9] ));
 sg13g2_dfrbp_1 _6194_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net343),
    .D(net1074),
    .Q_N(_2657_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[10] ));
 sg13g2_dfrbp_1 _6195_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net339),
    .D(net966),
    .Q_N(_2656_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[11] ));
 sg13g2_dfrbp_1 _6196_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net335),
    .D(_0353_),
    .Q_N(_2655_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[12] ));
 sg13g2_dfrbp_1 _6197_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net331),
    .D(net484),
    .Q_N(_2654_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[13] ));
 sg13g2_dfrbp_1 _6198_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net327),
    .D(net539),
    .Q_N(_2653_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[14] ));
 sg13g2_dfrbp_1 _6199_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net323),
    .D(_0356_),
    .Q_N(_2652_),
    .Q(\project_audio.genblk1[1].n_c_oh_my.phase[15] ));
 sg13g2_dfrbp_1 _6200_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net319),
    .D(_0357_),
    .Q_N(_2651_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.snd ));
 sg13g2_dfrbp_1 _6201_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net315),
    .D(_0358_),
    .Q_N(_2650_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[0] ));
 sg13g2_dfrbp_1 _6202_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net311),
    .D(_0359_),
    .Q_N(_2649_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[1] ));
 sg13g2_dfrbp_1 _6203_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net307),
    .D(net1054),
    .Q_N(_2648_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[2] ));
 sg13g2_dfrbp_1 _6204_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net303),
    .D(net962),
    .Q_N(_2647_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[3] ));
 sg13g2_dfrbp_1 _6205_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net299),
    .D(net1037),
    .Q_N(_2646_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[4] ));
 sg13g2_dfrbp_1 _6206_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net295),
    .D(_0363_),
    .Q_N(_2645_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[5] ));
 sg13g2_dfrbp_1 _6207_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net291),
    .D(_0364_),
    .Q_N(_2644_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[6] ));
 sg13g2_dfrbp_1 _6208_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net287),
    .D(net1076),
    .Q_N(_2643_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[7] ));
 sg13g2_dfrbp_1 _6209_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net283),
    .D(net994),
    .Q_N(_2642_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[8] ));
 sg13g2_dfrbp_1 _6210_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net279),
    .D(_0367_),
    .Q_N(_2641_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[9] ));
 sg13g2_dfrbp_1 _6211_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net275),
    .D(net1128),
    .Q_N(_2640_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[10] ));
 sg13g2_dfrbp_1 _6212_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net271),
    .D(net1125),
    .Q_N(_2639_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[11] ));
 sg13g2_dfrbp_1 _6213_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net251),
    .D(_0370_),
    .Q_N(_2638_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[12] ));
 sg13g2_dfrbp_1 _6214_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net243),
    .D(net490),
    .Q_N(_2637_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[13] ));
 sg13g2_dfrbp_1 _6215_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net235),
    .D(net451),
    .Q_N(_2636_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[14] ));
 sg13g2_dfrbp_1 _6216_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net227),
    .D(net456),
    .Q_N(_2635_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.phase[15] ));
 sg13g2_dfrbp_1 _6217_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net219),
    .D(net1083),
    .Q_N(_2634_),
    .Q(\project_audio.iter.mult2_shift[0] ));
 sg13g2_dfrbp_1 _6218_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net215),
    .D(net886),
    .Q_N(_2633_),
    .Q(\project_audio.iter.mult2_shift[1] ));
 sg13g2_dfrbp_1 _6219_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net211),
    .D(net847),
    .Q_N(_2632_),
    .Q(\project_audio.iter.mult2_shift[2] ));
 sg13g2_dfrbp_1 _6220_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net207),
    .D(net936),
    .Q_N(_2631_),
    .Q(\project_audio.iter.mult2_shift[3] ));
 sg13g2_dfrbp_1 _6221_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net203),
    .D(net857),
    .Q_N(_2630_),
    .Q(\project_audio.iter.mult2_shift[4] ));
 sg13g2_dfrbp_1 _6222_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net199),
    .D(net899),
    .Q_N(_2629_),
    .Q(\project_audio.iter.mult2_shift[5] ));
 sg13g2_dfrbp_1 _6223_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net195),
    .D(net895),
    .Q_N(_2628_),
    .Q(\project_audio.iter.mult2_shift[6] ));
 sg13g2_dfrbp_1 _6224_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net191),
    .D(net916),
    .Q_N(_2627_),
    .Q(\project_audio.iter.mult2_shift[7] ));
 sg13g2_dfrbp_1 _6225_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net187),
    .D(net835),
    .Q_N(_2626_),
    .Q(\project_audio.iter.mult2_shift[8] ));
 sg13g2_dfrbp_1 _6226_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net183),
    .D(net879),
    .Q_N(_2625_),
    .Q(\project_audio.iter.mult2_shift[9] ));
 sg13g2_dfrbp_1 _6227_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net165),
    .D(net902),
    .Q_N(_2624_),
    .Q(\project_audio.iter.mult2_shift[10] ));
 sg13g2_dfrbp_1 _6228_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net161),
    .D(net874),
    .Q_N(_2623_),
    .Q(\project_audio.iter.mult2_shift[11] ));
 sg13g2_dfrbp_1 _6229_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net157),
    .D(net871),
    .Q_N(_2622_),
    .Q(\project_audio.iter.mult2_shift[12] ));
 sg13g2_dfrbp_1 _6230_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net153),
    .D(net924),
    .Q_N(_2621_),
    .Q(\project_audio.iter.mult2_shift[13] ));
 sg13g2_dfrbp_1 _6231_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net149),
    .D(net864),
    .Q_N(_2620_),
    .Q(\project_audio.iter.mult2_shift[14] ));
 sg13g2_dfrbp_1 _6232_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net143),
    .D(net507),
    .Q_N(_2619_),
    .Q(\project_audio.iter.mult2_shift[15] ));
 sg13g2_dfrbp_1 _6233_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net139),
    .D(_0390_),
    .Q_N(_2618_),
    .Q(\project_audio.mixer.audio_out ));
 sg13g2_dfrbp_1 _6234_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net135),
    .D(_0391_),
    .Q_N(_0041_),
    .Q(\project_audio.mixer.counter[0] ));
 sg13g2_dfrbp_1 _6235_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net131),
    .D(net866),
    .Q_N(_2617_),
    .Q(\project_audio.mixer.counter[1] ));
 sg13g2_dfrbp_1 _6236_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net127),
    .D(net877),
    .Q_N(_2616_),
    .Q(\project_audio.mixer.counter[2] ));
 sg13g2_dfrbp_1 _6237_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net112),
    .D(net767),
    .Q_N(_2615_),
    .Q(\project_audio.mixer.counter[3] ));
 sg13g2_dfrbp_1 _6238_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net108),
    .D(net498),
    .Q_N(_2614_),
    .Q(\project_audio.genblk1[0].n_c_oh_my.step ));
 sg13g2_dfrbp_1 _6239_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net104),
    .D(_0396_),
    .Q_N(_2613_),
    .Q(\project_audio.iter.mult1_shift[16] ));
 sg13g2_dfrbp_1 _6240_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net96),
    .D(net960),
    .Q_N(_2612_),
    .Q(\project_audio.iter.mult1_shift[17] ));
 sg13g2_dfrbp_1 _6241_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net87),
    .D(_0398_),
    .Q_N(_0025_),
    .Q(\project_audio.iter.x[0] ));
 sg13g2_dfrbp_1 _6242_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net79),
    .D(_0399_),
    .Q_N(_0026_),
    .Q(\project_audio.iter.x[1] ));
 sg13g2_dfrbp_1 _6243_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net71),
    .D(_0400_),
    .Q_N(_0027_),
    .Q(\project_audio.iter.x[2] ));
 sg13g2_dfrbp_1 _6244_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net63),
    .D(net859),
    .Q_N(_0028_),
    .Q(\project_audio.iter.x[3] ));
 sg13g2_dfrbp_1 _6245_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net55),
    .D(_0402_),
    .Q_N(_0029_),
    .Q(\project_audio.iter.x[4] ));
 sg13g2_dfrbp_1 _6246_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net47),
    .D(_0403_),
    .Q_N(_0030_),
    .Q(\project_audio.iter.x[5] ));
 sg13g2_dfrbp_1 _6247_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net39),
    .D(_0404_),
    .Q_N(_0031_),
    .Q(\project_audio.iter.x[6] ));
 sg13g2_dfrbp_1 _6248_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net31),
    .D(net1159),
    .Q_N(_0032_),
    .Q(\project_audio.iter.x[7] ));
 sg13g2_dfrbp_1 _6249_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net23),
    .D(_0406_),
    .Q_N(_0033_),
    .Q(\project_audio.iter.x[8] ));
 sg13g2_dfrbp_1 _6250_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net15),
    .D(_0407_),
    .Q_N(_0034_),
    .Q(\project_audio.iter.x[9] ));
 sg13g2_dfrbp_1 _6251_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net425),
    .D(_0408_),
    .Q_N(_0035_),
    .Q(\project_audio.iter.x[10] ));
 sg13g2_dfrbp_1 _6252_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net417),
    .D(_0409_),
    .Q_N(_0036_),
    .Q(\project_audio.iter.x[11] ));
 sg13g2_dfrbp_1 _6253_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net409),
    .D(_0410_),
    .Q_N(_0037_),
    .Q(\project_audio.iter.x[12] ));
 sg13g2_dfrbp_1 _6254_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net401),
    .D(_0411_),
    .Q_N(_0038_),
    .Q(\project_audio.iter.x[13] ));
 sg13g2_dfrbp_1 _6255_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net393),
    .D(_0412_),
    .Q_N(_0039_),
    .Q(\project_audio.iter.x[14] ));
 sg13g2_dfrbp_1 _6256_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net385),
    .D(_0413_),
    .Q_N(_0001_),
    .Q(\project_audio.iter.x[15] ));
 sg13g2_dfrbp_1 _6257_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net377),
    .D(_0414_),
    .Q_N(_2611_),
    .Q(\project_audio.iter.next_ready ));
 sg13g2_dfrbp_1 _6258_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net373),
    .D(net438),
    .Q_N(_0040_),
    .Q(\project_audio.iter.counter[0] ));
 sg13g2_dfrbp_1 _6259_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net369),
    .D(net1213),
    .Q_N(_2610_),
    .Q(\project_audio.iter.counter[1] ));
 sg13g2_dfrbp_1 _6260_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net365),
    .D(_0417_),
    .Q_N(_2609_),
    .Q(\project_audio.iter.counter[2] ));
 sg13g2_dfrbp_1 _6261_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net361),
    .D(_0418_),
    .Q_N(_2608_),
    .Q(\project_audio.iter.counter[3] ));
 sg13g2_dfrbp_1 _6262_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net357),
    .D(_0419_),
    .Q_N(_2607_),
    .Q(\project_audio.iter.counter[4] ));
 sg13g2_dfrbp_1 _6263_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net353),
    .D(_0420_),
    .Q_N(_2606_),
    .Q(\project_audio.iter.counter[5] ));
 sg13g2_dfrbp_1 _6264_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net349),
    .D(_0421_),
    .Q_N(_2605_),
    .Q(\project_audio.iter.counter[6] ));
 sg13g2_dfrbp_1 _6265_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net345),
    .D(_0422_),
    .Q_N(_2604_),
    .Q(\project_audio.iter.counter[7] ));
 sg13g2_dfrbp_1 _6266_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net341),
    .D(_0423_),
    .Q_N(_2603_),
    .Q(\project_audio.iter.counter[8] ));
 sg13g2_dfrbp_1 _6267_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net337),
    .D(_0424_),
    .Q_N(_2602_),
    .Q(\project_audio.iter.counter[9] ));
 sg13g2_dfrbp_1 _6268_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net333),
    .D(_0425_),
    .Q_N(_2601_),
    .Q(\project_audio.iter.counter[10] ));
 sg13g2_dfrbp_1 _6269_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net329),
    .D(_0426_),
    .Q_N(_2600_),
    .Q(\project_audio.iter.counter[11] ));
 sg13g2_dfrbp_1 _6270_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net325),
    .D(_0427_),
    .Q_N(_2599_),
    .Q(\project_audio.iter.counter[12] ));
 sg13g2_dfrbp_1 _6271_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net321),
    .D(_0428_),
    .Q_N(_2598_),
    .Q(\project_audio.iter.counter[13] ));
 sg13g2_dfrbp_1 _6272_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net317),
    .D(_0429_),
    .Q_N(_0000_),
    .Q(\project_audio.r_counter ));
 sg13g2_dfrbp_1 _6273_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net309),
    .D(net453),
    .Q_N(_0002_),
    .Q(\project_audio.iter.r[0] ));
 sg13g2_dfrbp_1 _6274_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net301),
    .D(_0431_),
    .Q_N(_0005_),
    .Q(\project_audio.iter.r[1] ));
 sg13g2_dfrbp_1 _6275_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net293),
    .D(_0432_),
    .Q_N(_2597_),
    .Q(\project_audio.iter.r[2] ));
 sg13g2_dfrbp_1 _6276_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net285),
    .D(net486),
    .Q_N(_0006_),
    .Q(\project_audio.iter.r[3] ));
 sg13g2_dfrbp_1 _6277_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net277),
    .D(net850),
    .Q_N(_2596_),
    .Q(\project_audio.iter.r[4] ));
 sg13g2_dfrbp_1 _6278_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net269),
    .D(_0435_),
    .Q_N(_2595_),
    .Q(\project_audio.iter.r[5] ));
 sg13g2_dfrbp_1 _6279_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net239),
    .D(_0436_),
    .Q_N(_2594_),
    .Q(\project_audio.iter.r[6] ));
 sg13g2_dfrbp_1 _6280_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net223),
    .D(net1156),
    .Q_N(_2593_),
    .Q(\project_audio.iter.r[7] ));
 sg13g2_dfrbp_1 _6281_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net92),
    .D(_0438_),
    .Q_N(_2592_),
    .Q(\project_audio.iter.r[8] ));
 sg13g2_dfrbp_1 _6282_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net75),
    .D(_0439_),
    .Q_N(_2591_),
    .Q(\project_audio.iter.r[9] ));
 sg13g2_dfrbp_1 _6283_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net59),
    .D(_0440_),
    .Q_N(_2590_),
    .Q(\project_audio.iter.r[10] ));
 sg13g2_dfrbp_1 _6284_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net43),
    .D(net1002),
    .Q_N(_2589_),
    .Q(\project_audio.iter.r[11] ));
 sg13g2_dfrbp_1 _6285_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net27),
    .D(_0442_),
    .Q_N(_2588_),
    .Q(\project_audio.iter.r[12] ));
 sg13g2_dfrbp_1 _6286_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net429),
    .D(_0443_),
    .Q_N(_2587_),
    .Q(\project_audio.iter.r[13] ));
 sg13g2_dfrbp_1 _6287_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net413),
    .D(_0444_),
    .Q_N(_2586_),
    .Q(\project_audio.iter.r[14] ));
 sg13g2_dfrbp_1 _6288_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net397),
    .D(net1141),
    .Q_N(_2585_),
    .Q(\project_audio.iter.r[15] ));
 sg13g2_dfrbp_1 _6289_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net381),
    .D(net1217),
    .Q_N(_2584_),
    .Q(\project_audio.iter.r[16] ));
 sg13g2_dfrbp_1 _6290_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net305),
    .D(net1134),
    .Q_N(_0004_),
    .Q(\project_audio.iter.r[17] ));
 sg13g2_dfrbp_1 _6291_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net289),
    .D(net1183),
    .Q_N(_0021_),
    .Q(\project_audio.f_counter[0] ));
 sg13g2_dfrbp_1 _6292_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net273),
    .D(net1131),
    .Q_N(_2583_),
    .Q(\project_audio.f_counter[1] ));
 sg13g2_dfrbp_1 _6293_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net231),
    .D(net1072),
    .Q_N(_0003_),
    .Q(\project_audio.f_counter[2] ));
 sg13g2_dfrbp_1 _6294_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net83),
    .D(_0451_),
    .Q_N(_2582_),
    .Q(\project_audio.freq[1][0] ));
 sg13g2_dfrbp_1 _6295_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net51),
    .D(_0452_),
    .Q_N(_2581_),
    .Q(\project_audio.freq[1][1] ));
 sg13g2_dfrbp_1 _6296_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net19),
    .D(_0453_),
    .Q_N(_2580_),
    .Q(\project_audio.freq[1][2] ));
 sg13g2_dfrbp_1 _6297_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net405),
    .D(_0454_),
    .Q_N(_2579_),
    .Q(\project_audio.freq[1][3] ));
 sg13g2_dfrbp_1 _6298_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net313),
    .D(_0455_),
    .Q_N(_2578_),
    .Q(\project_audio.freq[1][4] ));
 sg13g2_dfrbp_1 _6299_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net281),
    .D(_0456_),
    .Q_N(_2577_),
    .Q(\project_audio.freq[1][5] ));
 sg13g2_dfrbp_1 _6300_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net100),
    .D(_0457_),
    .Q_N(_2576_),
    .Q(\project_audio.freq[1][6] ));
 sg13g2_dfrbp_1 _6301_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net35),
    .D(_0458_),
    .Q_N(_2575_),
    .Q(\project_audio.freq[1][7] ));
 sg13g2_dfrbp_1 _6302_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net389),
    .D(net763),
    .Q_N(_2574_),
    .Q(\project_audio.freq[1][8] ));
 sg13g2_dfrbp_1 _6303_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net247),
    .D(net826),
    .Q_N(_2573_),
    .Q(\project_audio.freq[1][9] ));
 sg13g2_dfrbp_1 _6304_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net421),
    .D(net523),
    .Q_N(_2572_),
    .Q(\project_audio.freq[1][10] ));
 sg13g2_dfrbp_1 _6305_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net67),
    .D(_0462_),
    .Q_N(_2571_),
    .Q(\project_audio.freq[1][11] ));
 sg13g2_tiehi _6036__16 (.L_HI(net16));
 sg13g2_tiehi _6171__17 (.L_HI(net17));
 sg13g2_tiehi _6035__18 (.L_HI(net18));
 sg13g2_tiehi _6296__19 (.L_HI(net19));
 sg13g2_tiehi _6034__20 (.L_HI(net20));
 sg13g2_tiehi _6170__21 (.L_HI(net21));
 sg13g2_tiehi _6033__22 (.L_HI(net22));
 sg13g2_tiehi _6249__23 (.L_HI(net23));
 sg13g2_tiehi _6032__24 (.L_HI(net24));
 sg13g2_tiehi _6169__25 (.L_HI(net25));
 sg13g2_tiehi _6031__26 (.L_HI(net26));
 sg13g2_tiehi _6285__27 (.L_HI(net27));
 sg13g2_tiehi _6030__28 (.L_HI(net28));
 sg13g2_tiehi _6168__29 (.L_HI(net29));
 sg13g2_tiehi _6029__30 (.L_HI(net30));
 sg13g2_tiehi _6248__31 (.L_HI(net31));
 sg13g2_tiehi _6028__32 (.L_HI(net32));
 sg13g2_tiehi _6167__33 (.L_HI(net33));
 sg13g2_tiehi _6027__34 (.L_HI(net34));
 sg13g2_tiehi _6301__35 (.L_HI(net35));
 sg13g2_tiehi _6026__36 (.L_HI(net36));
 sg13g2_tiehi _6166__37 (.L_HI(net37));
 sg13g2_tiehi _6025__38 (.L_HI(net38));
 sg13g2_tiehi _6247__39 (.L_HI(net39));
 sg13g2_tiehi _6024__40 (.L_HI(net40));
 sg13g2_tiehi _6165__41 (.L_HI(net41));
 sg13g2_tiehi _6023__42 (.L_HI(net42));
 sg13g2_tiehi _6284__43 (.L_HI(net43));
 sg13g2_tiehi _6022__44 (.L_HI(net44));
 sg13g2_tiehi _6164__45 (.L_HI(net45));
 sg13g2_tiehi _6021__46 (.L_HI(net46));
 sg13g2_tiehi _6246__47 (.L_HI(net47));
 sg13g2_tiehi _6020__48 (.L_HI(net48));
 sg13g2_tiehi _6163__49 (.L_HI(net49));
 sg13g2_tiehi _6019__50 (.L_HI(net50));
 sg13g2_tiehi _6295__51 (.L_HI(net51));
 sg13g2_tiehi _6018__52 (.L_HI(net52));
 sg13g2_tiehi _6162__53 (.L_HI(net53));
 sg13g2_tiehi _6017__54 (.L_HI(net54));
 sg13g2_tiehi _6245__55 (.L_HI(net55));
 sg13g2_tiehi _6016__56 (.L_HI(net56));
 sg13g2_tiehi _6161__57 (.L_HI(net57));
 sg13g2_tiehi _6015__58 (.L_HI(net58));
 sg13g2_tiehi _6283__59 (.L_HI(net59));
 sg13g2_tiehi _6014__60 (.L_HI(net60));
 sg13g2_tiehi _6160__61 (.L_HI(net61));
 sg13g2_tiehi _6013__62 (.L_HI(net62));
 sg13g2_tiehi _6244__63 (.L_HI(net63));
 sg13g2_tiehi _6012__64 (.L_HI(net64));
 sg13g2_tiehi _6159__65 (.L_HI(net65));
 sg13g2_tiehi _6011__66 (.L_HI(net66));
 sg13g2_tiehi _6305__67 (.L_HI(net67));
 sg13g2_tiehi _6010__68 (.L_HI(net68));
 sg13g2_tiehi _6158__69 (.L_HI(net69));
 sg13g2_tiehi _6009__70 (.L_HI(net70));
 sg13g2_tiehi _6243__71 (.L_HI(net71));
 sg13g2_tiehi _6008__72 (.L_HI(net72));
 sg13g2_tiehi _6157__73 (.L_HI(net73));
 sg13g2_tiehi _6007__74 (.L_HI(net74));
 sg13g2_tiehi _6282__75 (.L_HI(net75));
 sg13g2_tiehi _6006__76 (.L_HI(net76));
 sg13g2_tiehi _6156__77 (.L_HI(net77));
 sg13g2_tiehi _6005__78 (.L_HI(net78));
 sg13g2_tiehi _6242__79 (.L_HI(net79));
 sg13g2_tiehi _6004__80 (.L_HI(net80));
 sg13g2_tiehi _6155__81 (.L_HI(net81));
 sg13g2_tiehi _6003__82 (.L_HI(net82));
 sg13g2_tiehi _6294__83 (.L_HI(net83));
 sg13g2_tiehi _6002__84 (.L_HI(net84));
 sg13g2_tiehi _6154__85 (.L_HI(net85));
 sg13g2_tiehi _6001__86 (.L_HI(net86));
 sg13g2_tiehi _6241__87 (.L_HI(net87));
 sg13g2_tiehi _6000__88 (.L_HI(net88));
 sg13g2_tiehi _6153__89 (.L_HI(net89));
 sg13g2_tiehi _5999__90 (.L_HI(net90));
 sg13g2_tiehi _5998__91 (.L_HI(net91));
 sg13g2_tiehi _6281__92 (.L_HI(net92));
 sg13g2_tiehi _5997__93 (.L_HI(net93));
 sg13g2_tiehi _6152__94 (.L_HI(net94));
 sg13g2_tiehi _5996__95 (.L_HI(net95));
 sg13g2_tiehi _6240__96 (.L_HI(net96));
 sg13g2_tiehi _5995__97 (.L_HI(net97));
 sg13g2_tiehi _6151__98 (.L_HI(net98));
 sg13g2_tiehi _5994__99 (.L_HI(net99));
 sg13g2_tiehi _6300__100 (.L_HI(net100));
 sg13g2_tiehi _5993__101 (.L_HI(net101));
 sg13g2_tiehi _6150__102 (.L_HI(net102));
 sg13g2_tiehi _5992__103 (.L_HI(net103));
 sg13g2_tiehi _6239__104 (.L_HI(net104));
 sg13g2_tiehi _5991__105 (.L_HI(net105));
 sg13g2_tiehi _6149__106 (.L_HI(net106));
 sg13g2_tiehi _5990__107 (.L_HI(net107));
 sg13g2_tiehi _6238__108 (.L_HI(net108));
 sg13g2_tiehi _5989__109 (.L_HI(net109));
 sg13g2_tiehi _6148__110 (.L_HI(net110));
 sg13g2_tiehi _5988__111 (.L_HI(net111));
 sg13g2_tiehi _6237__112 (.L_HI(net112));
 sg13g2_tiehi _5987__113 (.L_HI(net113));
 sg13g2_tiehi _6147__114 (.L_HI(net114));
 sg13g2_tiehi _5986__115 (.L_HI(net115));
 sg13g2_tiehi _5985__116 (.L_HI(net116));
 sg13g2_tiehi _5984__117 (.L_HI(net117));
 sg13g2_tiehi _5983__118 (.L_HI(net118));
 sg13g2_tiehi _5982__119 (.L_HI(net119));
 sg13g2_tiehi _5981__120 (.L_HI(net120));
 sg13g2_tiehi _5980__121 (.L_HI(net121));
 sg13g2_tiehi _5979__122 (.L_HI(net122));
 sg13g2_tiehi _5978__123 (.L_HI(net123));
 sg13g2_tiehi _5977__124 (.L_HI(net124));
 sg13g2_tiehi _5976__125 (.L_HI(net125));
 sg13g2_tiehi _5975__126 (.L_HI(net126));
 sg13g2_tiehi _6236__127 (.L_HI(net127));
 sg13g2_tiehi _5974__128 (.L_HI(net128));
 sg13g2_tiehi _6146__129 (.L_HI(net129));
 sg13g2_tiehi _5973__130 (.L_HI(net130));
 sg13g2_tiehi _6235__131 (.L_HI(net131));
 sg13g2_tiehi _5972__132 (.L_HI(net132));
 sg13g2_tiehi _6145__133 (.L_HI(net133));
 sg13g2_tiehi _5971__134 (.L_HI(net134));
 sg13g2_tiehi _6234__135 (.L_HI(net135));
 sg13g2_tiehi _5970__136 (.L_HI(net136));
 sg13g2_tiehi _6144__137 (.L_HI(net137));
 sg13g2_tiehi _5969__138 (.L_HI(net138));
 sg13g2_tiehi _6233__139 (.L_HI(net139));
 sg13g2_tiehi _5968__140 (.L_HI(net140));
 sg13g2_tiehi _6143__141 (.L_HI(net141));
 sg13g2_tiehi _5967__142 (.L_HI(net142));
 sg13g2_tiehi _6232__143 (.L_HI(net143));
 sg13g2_tiehi _5966__144 (.L_HI(net144));
 sg13g2_tiehi _6142__145 (.L_HI(net145));
 sg13g2_tiehi _5965__146 (.L_HI(net146));
 sg13g2_tiehi _5964__147 (.L_HI(net147));
 sg13g2_tiehi _5963__148 (.L_HI(net148));
 sg13g2_tiehi _6231__149 (.L_HI(net149));
 sg13g2_tiehi _5962__150 (.L_HI(net150));
 sg13g2_tiehi _6141__151 (.L_HI(net151));
 sg13g2_tiehi _5961__152 (.L_HI(net152));
 sg13g2_tiehi _6230__153 (.L_HI(net153));
 sg13g2_tiehi _5960__154 (.L_HI(net154));
 sg13g2_tiehi _6140__155 (.L_HI(net155));
 sg13g2_tiehi _5959__156 (.L_HI(net156));
 sg13g2_tiehi _6229__157 (.L_HI(net157));
 sg13g2_tiehi _5958__158 (.L_HI(net158));
 sg13g2_tiehi _6139__159 (.L_HI(net159));
 sg13g2_tiehi _5957__160 (.L_HI(net160));
 sg13g2_tiehi _6228__161 (.L_HI(net161));
 sg13g2_tiehi _5956__162 (.L_HI(net162));
 sg13g2_tiehi _6138__163 (.L_HI(net163));
 sg13g2_tiehi _5955__164 (.L_HI(net164));
 sg13g2_tiehi _6227__165 (.L_HI(net165));
 sg13g2_tiehi _5954__166 (.L_HI(net166));
 sg13g2_tiehi _5953__167 (.L_HI(net167));
 sg13g2_tiehi _5952__168 (.L_HI(net168));
 sg13g2_tiehi _5951__169 (.L_HI(net169));
 sg13g2_tiehi _5950__170 (.L_HI(net170));
 sg13g2_tiehi _5949__171 (.L_HI(net171));
 sg13g2_tiehi _5948__172 (.L_HI(net172));
 sg13g2_tiehi _5947__173 (.L_HI(net173));
 sg13g2_tiehi _5946__174 (.L_HI(net174));
 sg13g2_tiehi _5945__175 (.L_HI(net175));
 sg13g2_tiehi _5944__176 (.L_HI(net176));
 sg13g2_tiehi _5943__177 (.L_HI(net177));
 sg13g2_tiehi _5942__178 (.L_HI(net178));
 sg13g2_tiehi _5941__179 (.L_HI(net179));
 sg13g2_tiehi _5940__180 (.L_HI(net180));
 sg13g2_tiehi _6137__181 (.L_HI(net181));
 sg13g2_tiehi _5939__182 (.L_HI(net182));
 sg13g2_tiehi _6226__183 (.L_HI(net183));
 sg13g2_tiehi _5938__184 (.L_HI(net184));
 sg13g2_tiehi _6136__185 (.L_HI(net185));
 sg13g2_tiehi _5937__186 (.L_HI(net186));
 sg13g2_tiehi _6225__187 (.L_HI(net187));
 sg13g2_tiehi _5936__188 (.L_HI(net188));
 sg13g2_tiehi _6135__189 (.L_HI(net189));
 sg13g2_tiehi _5935__190 (.L_HI(net190));
 sg13g2_tiehi _6224__191 (.L_HI(net191));
 sg13g2_tiehi _5934__192 (.L_HI(net192));
 sg13g2_tiehi _6134__193 (.L_HI(net193));
 sg13g2_tiehi _5933__194 (.L_HI(net194));
 sg13g2_tiehi _6223__195 (.L_HI(net195));
 sg13g2_tiehi _5932__196 (.L_HI(net196));
 sg13g2_tiehi _6133__197 (.L_HI(net197));
 sg13g2_tiehi _5931__198 (.L_HI(net198));
 sg13g2_tiehi _6222__199 (.L_HI(net199));
 sg13g2_tiehi _5930__200 (.L_HI(net200));
 sg13g2_tiehi _6132__201 (.L_HI(net201));
 sg13g2_tiehi _5929__202 (.L_HI(net202));
 sg13g2_tiehi _6221__203 (.L_HI(net203));
 sg13g2_tiehi _5928__204 (.L_HI(net204));
 sg13g2_tiehi _6131__205 (.L_HI(net205));
 sg13g2_tiehi _5927__206 (.L_HI(net206));
 sg13g2_tiehi _6220__207 (.L_HI(net207));
 sg13g2_tiehi _5926__208 (.L_HI(net208));
 sg13g2_tiehi _6130__209 (.L_HI(net209));
 sg13g2_tiehi _5925__210 (.L_HI(net210));
 sg13g2_tiehi _6219__211 (.L_HI(net211));
 sg13g2_tiehi _5924__212 (.L_HI(net212));
 sg13g2_tiehi _6129__213 (.L_HI(net213));
 sg13g2_tiehi _5923__214 (.L_HI(net214));
 sg13g2_tiehi _6218__215 (.L_HI(net215));
 sg13g2_tiehi _5922__216 (.L_HI(net216));
 sg13g2_tiehi _6128__217 (.L_HI(net217));
 sg13g2_tiehi _5921__218 (.L_HI(net218));
 sg13g2_tiehi _6217__219 (.L_HI(net219));
 sg13g2_tiehi _5920__220 (.L_HI(net220));
 sg13g2_tiehi _6127__221 (.L_HI(net221));
 sg13g2_tiehi _5919__222 (.L_HI(net222));
 sg13g2_tiehi _6280__223 (.L_HI(net223));
 sg13g2_tiehi _5918__224 (.L_HI(net224));
 sg13g2_tiehi _6126__225 (.L_HI(net225));
 sg13g2_tiehi _5917__226 (.L_HI(net226));
 sg13g2_tiehi _6216__227 (.L_HI(net227));
 sg13g2_tiehi _5916__228 (.L_HI(net228));
 sg13g2_tiehi _6125__229 (.L_HI(net229));
 sg13g2_tiehi _5915__230 (.L_HI(net230));
 sg13g2_tiehi _6293__231 (.L_HI(net231));
 sg13g2_tiehi _5914__232 (.L_HI(net232));
 sg13g2_tiehi _6124__233 (.L_HI(net233));
 sg13g2_tiehi _5913__234 (.L_HI(net234));
 sg13g2_tiehi _6215__235 (.L_HI(net235));
 sg13g2_tiehi _5912__236 (.L_HI(net236));
 sg13g2_tiehi _6123__237 (.L_HI(net237));
 sg13g2_tiehi _5911__238 (.L_HI(net238));
 sg13g2_tiehi _6279__239 (.L_HI(net239));
 sg13g2_tiehi _5910__240 (.L_HI(net240));
 sg13g2_tiehi _6122__241 (.L_HI(net241));
 sg13g2_tiehi _5909__242 (.L_HI(net242));
 sg13g2_tiehi _6214__243 (.L_HI(net243));
 sg13g2_tiehi _5908__244 (.L_HI(net244));
 sg13g2_tiehi _6121__245 (.L_HI(net245));
 sg13g2_tiehi _5907__246 (.L_HI(net246));
 sg13g2_tiehi _6303__247 (.L_HI(net247));
 sg13g2_tiehi _5906__248 (.L_HI(net248));
 sg13g2_tiehi _6120__249 (.L_HI(net249));
 sg13g2_tiehi _5905__250 (.L_HI(net250));
 sg13g2_tiehi _6213__251 (.L_HI(net251));
 sg13g2_tiehi _5904__252 (.L_HI(net252));
 sg13g2_tiehi _5903__253 (.L_HI(net253));
 sg13g2_tiehi _5902__254 (.L_HI(net254));
 sg13g2_tiehi _5901__255 (.L_HI(net255));
 sg13g2_tiehi _5900__256 (.L_HI(net256));
 sg13g2_tiehi _5899__257 (.L_HI(net257));
 sg13g2_tiehi _5898__258 (.L_HI(net258));
 sg13g2_tiehi _5897__259 (.L_HI(net259));
 sg13g2_tiehi _5896__260 (.L_HI(net260));
 sg13g2_tiehi _5895__261 (.L_HI(net261));
 sg13g2_tiehi _5894__262 (.L_HI(net262));
 sg13g2_tiehi _5893__263 (.L_HI(net263));
 sg13g2_tiehi _5892__264 (.L_HI(net264));
 sg13g2_tiehi _5891__265 (.L_HI(net265));
 sg13g2_tiehi _5890__266 (.L_HI(net266));
 sg13g2_tiehi _5889__267 (.L_HI(net267));
 sg13g2_tiehi _6119__268 (.L_HI(net268));
 sg13g2_tiehi _6278__269 (.L_HI(net269));
 sg13g2_tiehi _6118__270 (.L_HI(net270));
 sg13g2_tiehi _6212__271 (.L_HI(net271));
 sg13g2_tiehi _6117__272 (.L_HI(net272));
 sg13g2_tiehi _6292__273 (.L_HI(net273));
 sg13g2_tiehi _6116__274 (.L_HI(net274));
 sg13g2_tiehi _6211__275 (.L_HI(net275));
 sg13g2_tiehi _6115__276 (.L_HI(net276));
 sg13g2_tiehi _6277__277 (.L_HI(net277));
 sg13g2_tiehi _6114__278 (.L_HI(net278));
 sg13g2_tiehi _6210__279 (.L_HI(net279));
 sg13g2_tiehi _6113__280 (.L_HI(net280));
 sg13g2_tiehi _6299__281 (.L_HI(net281));
 sg13g2_tiehi _6112__282 (.L_HI(net282));
 sg13g2_tiehi _6209__283 (.L_HI(net283));
 sg13g2_tiehi _6111__284 (.L_HI(net284));
 sg13g2_tiehi _6276__285 (.L_HI(net285));
 sg13g2_tiehi _6110__286 (.L_HI(net286));
 sg13g2_tiehi _6208__287 (.L_HI(net287));
 sg13g2_tiehi _6109__288 (.L_HI(net288));
 sg13g2_tiehi _6291__289 (.L_HI(net289));
 sg13g2_tiehi _6108__290 (.L_HI(net290));
 sg13g2_tiehi _6207__291 (.L_HI(net291));
 sg13g2_tiehi _6107__292 (.L_HI(net292));
 sg13g2_tiehi _6275__293 (.L_HI(net293));
 sg13g2_tiehi _6106__294 (.L_HI(net294));
 sg13g2_tiehi _6206__295 (.L_HI(net295));
 sg13g2_tiehi _6105__296 (.L_HI(net296));
 sg13g2_tiehi _5888__297 (.L_HI(net297));
 sg13g2_tiehi _6104__298 (.L_HI(net298));
 sg13g2_tiehi _6205__299 (.L_HI(net299));
 sg13g2_tiehi _6103__300 (.L_HI(net300));
 sg13g2_tiehi _6274__301 (.L_HI(net301));
 sg13g2_tiehi _6102__302 (.L_HI(net302));
 sg13g2_tiehi _6204__303 (.L_HI(net303));
 sg13g2_tiehi _6101__304 (.L_HI(net304));
 sg13g2_tiehi _6290__305 (.L_HI(net305));
 sg13g2_tiehi _6100__306 (.L_HI(net306));
 sg13g2_tiehi _6203__307 (.L_HI(net307));
 sg13g2_tiehi _6099__308 (.L_HI(net308));
 sg13g2_tiehi _6273__309 (.L_HI(net309));
 sg13g2_tiehi _6098__310 (.L_HI(net310));
 sg13g2_tiehi _6202__311 (.L_HI(net311));
 sg13g2_tiehi _6097__312 (.L_HI(net312));
 sg13g2_tiehi _6298__313 (.L_HI(net313));
 sg13g2_tiehi _6096__314 (.L_HI(net314));
 sg13g2_tiehi _6201__315 (.L_HI(net315));
 sg13g2_tiehi _6095__316 (.L_HI(net316));
 sg13g2_tiehi _6272__317 (.L_HI(net317));
 sg13g2_tiehi _6094__318 (.L_HI(net318));
 sg13g2_tiehi _6200__319 (.L_HI(net319));
 sg13g2_tiehi _6093__320 (.L_HI(net320));
 sg13g2_tiehi _6271__321 (.L_HI(net321));
 sg13g2_tiehi _6092__322 (.L_HI(net322));
 sg13g2_tiehi _6199__323 (.L_HI(net323));
 sg13g2_tiehi _6091__324 (.L_HI(net324));
 sg13g2_tiehi _6270__325 (.L_HI(net325));
 sg13g2_tiehi _6090__326 (.L_HI(net326));
 sg13g2_tiehi _6198__327 (.L_HI(net327));
 sg13g2_tiehi _6089__328 (.L_HI(net328));
 sg13g2_tiehi _6269__329 (.L_HI(net329));
 sg13g2_tiehi _6088__330 (.L_HI(net330));
 sg13g2_tiehi _6197__331 (.L_HI(net331));
 sg13g2_tiehi _6087__332 (.L_HI(net332));
 sg13g2_tiehi _6268__333 (.L_HI(net333));
 sg13g2_tiehi _6086__334 (.L_HI(net334));
 sg13g2_tiehi _6196__335 (.L_HI(net335));
 sg13g2_tiehi _6085__336 (.L_HI(net336));
 sg13g2_tiehi _6267__337 (.L_HI(net337));
 sg13g2_tiehi _6084__338 (.L_HI(net338));
 sg13g2_tiehi _6195__339 (.L_HI(net339));
 sg13g2_tiehi _6083__340 (.L_HI(net340));
 sg13g2_tiehi _6266__341 (.L_HI(net341));
 sg13g2_tiehi _6082__342 (.L_HI(net342));
 sg13g2_tiehi _6194__343 (.L_HI(net343));
 sg13g2_tiehi _6081__344 (.L_HI(net344));
 sg13g2_tiehi _6265__345 (.L_HI(net345));
 sg13g2_tiehi _6080__346 (.L_HI(net346));
 sg13g2_tiehi _6193__347 (.L_HI(net347));
 sg13g2_tiehi _6079__348 (.L_HI(net348));
 sg13g2_tiehi _6264__349 (.L_HI(net349));
 sg13g2_tiehi _6078__350 (.L_HI(net350));
 sg13g2_tiehi _6192__351 (.L_HI(net351));
 sg13g2_tiehi _6077__352 (.L_HI(net352));
 sg13g2_tiehi _6263__353 (.L_HI(net353));
 sg13g2_tiehi _6076__354 (.L_HI(net354));
 sg13g2_tiehi _6191__355 (.L_HI(net355));
 sg13g2_tiehi _6075__356 (.L_HI(net356));
 sg13g2_tiehi _6262__357 (.L_HI(net357));
 sg13g2_tiehi _6074__358 (.L_HI(net358));
 sg13g2_tiehi _6190__359 (.L_HI(net359));
 sg13g2_tiehi _6073__360 (.L_HI(net360));
 sg13g2_tiehi _6261__361 (.L_HI(net361));
 sg13g2_tiehi _6072__362 (.L_HI(net362));
 sg13g2_tiehi _6189__363 (.L_HI(net363));
 sg13g2_tiehi _6071__364 (.L_HI(net364));
 sg13g2_tiehi _6260__365 (.L_HI(net365));
 sg13g2_tiehi _6070__366 (.L_HI(net366));
 sg13g2_tiehi _6188__367 (.L_HI(net367));
 sg13g2_tiehi _6069__368 (.L_HI(net368));
 sg13g2_tiehi _6259__369 (.L_HI(net369));
 sg13g2_tiehi _6068__370 (.L_HI(net370));
 sg13g2_tiehi _6187__371 (.L_HI(net371));
 sg13g2_tiehi _6067__372 (.L_HI(net372));
 sg13g2_tiehi _6258__373 (.L_HI(net373));
 sg13g2_tiehi _6066__374 (.L_HI(net374));
 sg13g2_tiehi _6186__375 (.L_HI(net375));
 sg13g2_tiehi _6065__376 (.L_HI(net376));
 sg13g2_tiehi _6257__377 (.L_HI(net377));
 sg13g2_tiehi _6064__378 (.L_HI(net378));
 sg13g2_tiehi _6185__379 (.L_HI(net379));
 sg13g2_tiehi _6063__380 (.L_HI(net380));
 sg13g2_tiehi _6289__381 (.L_HI(net381));
 sg13g2_tiehi _6062__382 (.L_HI(net382));
 sg13g2_tiehi _6184__383 (.L_HI(net383));
 sg13g2_tiehi _6061__384 (.L_HI(net384));
 sg13g2_tiehi _6256__385 (.L_HI(net385));
 sg13g2_tiehi _6060__386 (.L_HI(net386));
 sg13g2_tiehi _6183__387 (.L_HI(net387));
 sg13g2_tiehi _6059__388 (.L_HI(net388));
 sg13g2_tiehi _6302__389 (.L_HI(net389));
 sg13g2_tiehi _6058__390 (.L_HI(net390));
 sg13g2_tiehi _6182__391 (.L_HI(net391));
 sg13g2_tiehi _6057__392 (.L_HI(net392));
 sg13g2_tiehi _6255__393 (.L_HI(net393));
 sg13g2_tiehi _6056__394 (.L_HI(net394));
 sg13g2_tiehi _6181__395 (.L_HI(net395));
 sg13g2_tiehi _6055__396 (.L_HI(net396));
 sg13g2_tiehi _6288__397 (.L_HI(net397));
 sg13g2_tiehi _6054__398 (.L_HI(net398));
 sg13g2_tiehi _6180__399 (.L_HI(net399));
 sg13g2_tiehi _6053__400 (.L_HI(net400));
 sg13g2_tiehi _6254__401 (.L_HI(net401));
 sg13g2_tiehi _6052__402 (.L_HI(net402));
 sg13g2_tiehi _6179__403 (.L_HI(net403));
 sg13g2_tiehi _6051__404 (.L_HI(net404));
 sg13g2_tiehi _6297__405 (.L_HI(net405));
 sg13g2_tiehi _6050__406 (.L_HI(net406));
 sg13g2_tiehi _6178__407 (.L_HI(net407));
 sg13g2_tiehi _6049__408 (.L_HI(net408));
 sg13g2_tiehi _6253__409 (.L_HI(net409));
 sg13g2_tiehi _6048__410 (.L_HI(net410));
 sg13g2_tiehi _6177__411 (.L_HI(net411));
 sg13g2_tiehi _6047__412 (.L_HI(net412));
 sg13g2_tiehi _6287__413 (.L_HI(net413));
 sg13g2_tiehi _6046__414 (.L_HI(net414));
 sg13g2_tiehi _6176__415 (.L_HI(net415));
 sg13g2_tiehi _6045__416 (.L_HI(net416));
 sg13g2_tiehi _6252__417 (.L_HI(net417));
 sg13g2_tiehi _6044__418 (.L_HI(net418));
 sg13g2_tiehi _6175__419 (.L_HI(net419));
 sg13g2_tiehi _6043__420 (.L_HI(net420));
 sg13g2_tiehi _6304__421 (.L_HI(net421));
 sg13g2_tiehi _6042__422 (.L_HI(net422));
 sg13g2_tiehi _6174__423 (.L_HI(net423));
 sg13g2_tiehi _6041__424 (.L_HI(net424));
 sg13g2_tiehi _6251__425 (.L_HI(net425));
 sg13g2_tiehi _6040__426 (.L_HI(net426));
 sg13g2_tiehi _6173__427 (.L_HI(net427));
 sg13g2_tiehi _6039__428 (.L_HI(net428));
 sg13g2_tiehi _6286__429 (.L_HI(net429));
 sg13g2_tiehi _6038__430 (.L_HI(net430));
 sg13g2_tiehi _6172__431 (.L_HI(net431));
 sg13g2_tiehi _6037__432 (.L_HI(net432));
 sg13g2_tiehi tt_um_zec_square1_433 (.L_HI(net433));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_zec_square1_2 (.L_LO(net2));
 sg13g2_tielo tt_um_zec_square1_3 (.L_LO(net3));
 sg13g2_tielo tt_um_zec_square1_4 (.L_LO(net4));
 sg13g2_tielo tt_um_zec_square1_5 (.L_LO(net5));
 sg13g2_tielo tt_um_zec_square1_6 (.L_LO(net6));
 sg13g2_tielo tt_um_zec_square1_7 (.L_LO(net7));
 sg13g2_tielo tt_um_zec_square1_8 (.L_LO(net8));
 sg13g2_tielo tt_um_zec_square1_9 (.L_LO(net9));
 sg13g2_tielo tt_um_zec_square1_10 (.L_LO(net10));
 sg13g2_tielo tt_um_zec_square1_11 (.L_LO(net11));
 sg13g2_tielo tt_um_zec_square1_12 (.L_LO(net12));
 sg13g2_tielo tt_um_zec_square1_13 (.L_LO(net13));
 sg13g2_tielo tt_um_zec_square1_14 (.L_LO(net14));
 sg13g2_tiehi _6250__15 (.L_HI(net15));
 sg13g2_buf_2 _6739_ (.A(\project_audio.mixer.audio_out ),
    .X(uio_out[7]));
 sg13g2_buf_1 _6740_ (.A(\sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _6741_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(_1417_));
 sg13g2_buf_1 fanout541 (.A(_1417_),
    .X(net541));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(_1416_));
 sg13g2_buf_2 fanout543 (.A(_1416_),
    .X(net543));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(_1416_));
 sg13g2_buf_2 fanout545 (.A(_1413_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_1413_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(net549),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_1413_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net551),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_2552_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(_2552_));
 sg13g2_buf_2 fanout555 (.A(net557),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(net557),
    .X(net556));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(_2551_));
 sg13g2_buf_2 fanout558 (.A(net559),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(net561),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_2551_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(net566),
    .X(net562));
 sg13g2_buf_1 fanout563 (.A(net566),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(net566),
    .X(net564));
 sg13g2_buf_1 fanout565 (.A(net566),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_2550_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net572),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_1 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_1 fanout572 (.A(_2538_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net576),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_2538_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net580),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_2544_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_1 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(_2539_));
 sg13g2_buf_2 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(net589),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net589),
    .X(net587));
 sg13g2_buf_1 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(_2328_));
 sg13g2_buf_2 fanout590 (.A(_1002_),
    .X(net590));
 sg13g2_buf_1 fanout591 (.A(_1002_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_0989_),
    .X(net592));
 sg13g2_buf_1 fanout593 (.A(_0989_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_2440_),
    .X(net594));
 sg13g2_buf_1 fanout595 (.A(_2440_),
    .X(net595));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(_2439_));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(_1387_));
 sg13g2_buf_1 fanout598 (.A(_1387_),
    .X(net598));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(_1386_));
 sg13g2_buf_2 fanout600 (.A(_1374_),
    .X(net600));
 sg13g2_buf_1 fanout601 (.A(_1374_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_1373_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_1360_),
    .X(net603));
 sg13g2_buf_1 fanout604 (.A(_1360_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_1359_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_1346_),
    .X(net606));
 sg13g2_buf_1 fanout607 (.A(_1346_),
    .X(net607));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(_1345_));
 sg13g2_buf_2 fanout609 (.A(_1001_),
    .X(net609));
 sg13g2_buf_1 fanout610 (.A(_1001_),
    .X(net610));
 sg13g2_buf_4 fanout611 (.X(net611),
    .A(_0988_));
 sg13g2_buf_1 fanout612 (.A(_0988_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_0503_),
    .X(net614));
 sg13g2_buf_4 fanout615 (.X(net615),
    .A(_0502_));
 sg13g2_buf_2 fanout616 (.A(_2346_),
    .X(net616));
 sg13g2_buf_1 fanout617 (.A(_2346_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_1072_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_1067_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_1061_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_1 fanout623 (.A(_1052_),
    .X(net623));
 sg13g2_buf_4 fanout624 (.X(net624),
    .A(\project_audio.f_counter[1] ));
 sg13g2_buf_2 fanout625 (.A(net626),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(net1192),
    .X(net626));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(net1199));
 sg13g2_buf_4 fanout628 (.X(net628),
    .A(net629));
 sg13g2_buf_2 fanout629 (.A(net1172),
    .X(net629));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(\project_audio.iter.x[7] ));
 sg13g2_buf_2 fanout631 (.A(\project_audio.iter.x[3] ),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(net634),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net668),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(net637),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net637),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(net668),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(net642),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(net647),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(net647),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(net647),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(net647),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(net668),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(net651),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(net651),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(net668),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(net657),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(net656),
    .X(net654));
 sg13g2_buf_1 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(net657),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(net668),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(net661),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(net661),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(net667),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(net664),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(net664),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net667),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(net666),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(\project_audio.genblk1[0].n_c_oh_my.step ));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(net1239));
 sg13g2_buf_2 fanout670 (.A(net1232),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(net674),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(net1206),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(net676),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(\frame_no[2] ),
    .X(net676));
 sg13g2_buf_4 fanout677 (.X(net677),
    .A(net1221));
 sg13g2_buf_1 fanout678 (.A(\frame_no[1] ),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(\frame_no[0] ),
    .X(net679));
 sg13g2_buf_4 fanout680 (.X(net680),
    .A(net685));
 sg13g2_buf_2 fanout681 (.A(net685),
    .X(net681));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(net685));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(net684));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(net685));
 sg13g2_buf_2 fanout685 (.A(_2513_),
    .X(net685));
 sg13g2_buf_4 fanout686 (.X(net686),
    .A(net689));
 sg13g2_buf_2 fanout687 (.A(net689),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(net689),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(net716));
 sg13g2_buf_4 fanout691 (.X(net691),
    .A(net693));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_4 fanout693 (.X(net693),
    .A(net716));
 sg13g2_buf_2 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(net700));
 sg13g2_buf_2 fanout696 (.A(net699),
    .X(net696));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(net699));
 sg13g2_buf_1 fanout698 (.A(net699),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(net716),
    .X(net700));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(net703));
 sg13g2_buf_2 fanout702 (.A(net715),
    .X(net702));
 sg13g2_buf_4 fanout703 (.X(net703),
    .A(net715));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(net708));
 sg13g2_buf_2 fanout705 (.A(net708),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(net708),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(net715),
    .X(net708));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(net710));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(net714));
 sg13g2_buf_2 fanout711 (.A(net713),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(net715),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(rst_n),
    .X(net716));
 sg13g2_tielo tt_um_zec_square1_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_4_11_0_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_4_13_0_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_56_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_57_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_55_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_11_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_16_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_19_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_40_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_35_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_47_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_48_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_36_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_24_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_42_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_49_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_25_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_29_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_31_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0044_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0042_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0134_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0040_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0415_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0043_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0111_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0000_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold9 (.A(_2371_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0041_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold11 (.A(\project_audio.freq[6][11] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold12 (.A(\project_audio.freq[2][11] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold13 (.A(\project_audio.freq[1][11] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold14 (.A(\project_audio.freq[7][11] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold15 (.A(\project_audio.freq[4][11] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold16 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[14] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold17 (.A(_2203_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0372_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold19 (.A(\project_audio.iter.r[0] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0430_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold21 (.A(\project_audio.freq[3][11] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold22 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[15] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0373_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold24 (.A(\frame_no[8] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0119_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold26 (.A(\project_audio.nco_increment_gen.counter[7] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold27 (.A(_1343_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0141_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold29 (.A(\project_audio.freq[5][11] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold30 (.A(\project_audio.freq[0][5] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold31 (.A(\project_audio.nco_increment_gen.counter[2] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold32 (.A(_1338_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0136_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold34 (.A(\project_audio.freq[4][5] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold35 (.A(\project_audio.freq[1][0] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold36 (.A(\project_audio.freq[5][5] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold37 (.A(\project_audio.freq[3][0] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0156_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold39 (.A(\project_audio.freq[2][0] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold40 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[12] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold41 (.A(\project_audio.freq[5][0] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold42 (.A(\project_audio.freq[6][5] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold43 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[13] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0337_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold45 (.A(\project_audio.freq[1][5] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold46 (.A(\project_audio.freq[0][0] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold47 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[13] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0320_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold49 (.A(\project_audio.freq[4][0] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold50 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[13] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0354_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold52 (.A(\project_audio.iter.r[3] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0433_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold54 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[13] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0303_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold56 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[13] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0371_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold58 (.A(\project_audio.freq[3][5] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold59 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[15] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0305_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold61 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[15] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0288_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold63 (.A(\project_audio.freq[4][8] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold64 (.A(\project_audio.nco_increment_gen.counter[1] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0395_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold66 (.A(\project_audio.freq[7][4] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold67 (.A(\project_audio.freq[1][4] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold68 (.A(\project_audio.freq[3][1] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0157_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold70 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[13] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0269_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0001_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold73 (.A(_2265_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0389_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold75 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[12] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold76 (.A(\project_audio.freq[6][2] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold77 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[13] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold78 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[15] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0339_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold80 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[12] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold81 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[12] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold82 (.A(\project_audio.freq[2][1] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold83 (.A(\project_audio.iter.mult_accum[4] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold84 (.A(\project_audio.freq[5][4] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold85 (.A(\project_audio.freq[4][2] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0145_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold87 (.A(\project_audio.freq[4][4] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0147_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold89 (.A(\project_audio.freq[1][10] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0461_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold91 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[13] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold92 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[15] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0322_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold94 (.A(\project_audio.freq[5][6] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold95 (.A(\project_audio.freq[7][0] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold96 (.A(\project_audio.freq[0][7] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold97 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[15] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0271_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold99 (.A(\project_audio.freq[2][5] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold100 (.A(\project_audio.freq[6][4] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold101 (.A(\project_audio.freq[0][2] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold102 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[15] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0254_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold104 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[12] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold105 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[14] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0355_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold107 (.A(\project_audio.freq[7][10] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold108 (.A(\project_audio.freq[5][1] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0062_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold110 (.A(\project_audio.iter.r[2] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold111 (.A(_2392_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold112 (.A(\project_audio.freq[1][7] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold113 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[12] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold114 (.A(\project_audio.freq[3][10] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold115 (.A(\project_audio.freq[3][2] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0158_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold117 (.A(\project_audio.freq[7][7] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold118 (.A(\project_audio.freq[0][1] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold119 (.A(\project_audio.freq[5][3] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold120 (.A(\project_audio.iter.mult_accum[6] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold121 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[12] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold122 (.A(\project_audio.freq[2][6] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold123 (.A(\project_audio.freq[4][6] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold124 (.A(\project_audio.freq[2][8] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold125 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[14] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold126 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[14] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold127 (.A(\project_audio.freq[2][10] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold128 (.A(\project_audio.iter.mult_accum[7] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0213_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold130 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[15] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold131 (.A(\project_audio.freq[0][3] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold132 (.A(\project_audio.freq[2][4] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold133 (.A(\project_audio.freq[6][7] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold134 (.A(\project_audio.freq[5][7] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0068_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold136 (.A(\project_audio.freq[2][2] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold137 (.A(\project_audio.freq[1][1] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold138 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[14] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold139 (.A(\project_audio.freq[6][0] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold140 (.A(\project_audio.freq[1][6] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold141 (.A(\project_audio.nco_increment_gen.counter[3] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold142 (.A(_1339_),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0137_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold144 (.A(\project_audio.freq[5][2] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0063_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold146 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[14] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold147 (.A(\project_audio.freq[0][6] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold148 (.A(\project_audio.genblk1[0].n_c_oh_my.snd ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold149 (.A(\project_audio.iter.mult_accum[3] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold150 (.A(\project_audio.iter.mult1_shift[31] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0205_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold152 (.A(\project_audio.freq[1][8] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0459_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold154 (.A(\project_audio.freq[4][1] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold155 (.A(\project_audio.freq[3][7] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold156 (.A(\project_audio.mixer.counter[3] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0394_),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold158 (.A(\project_audio.freq[1][3] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold159 (.A(\project_audio.freq[3][8] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold160 (.A(\project_audio.iter.mult_accum[15] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0221_),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold162 (.A(\project_audio.freq[6][6] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold163 (.A(\project_audio.freq[2][7] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold164 (.A(\project_audio.iter.counter[13] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold165 (.A(_2369_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold166 (.A(\project_audio.freq[6][8] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold167 (.A(\project_audio.freq[7][1] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold168 (.A(\project_audio.freq[7][2] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold169 (.A(\project_audio.iter.mult_accum[1] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0207_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold171 (.A(\project_audio.freq[7][8] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold172 (.A(\project_audio.nco_increment_gen.counter[6] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0140_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold174 (.A(\project_audio.freq[0][8] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold175 (.A(\project_audio.freq[0][11] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold176 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[14] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold177 (.A(\project_audio.freq[1][2] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold178 (.A(\project_audio.freq[5][8] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold179 (.A(\project_audio.freq[2][3] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold180 (.A(\project_audio.nco_increment_gen.counter[4] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0138_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold182 (.A(\project_audio.freq[6][3] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold183 (.A(\sync_gen.vsync ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold184 (.A(\project_audio.freq[6][10] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold185 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[14] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold186 (.A(\project_audio.freq[4][3] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0146_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold188 (.A(\project_audio.freq[5][10] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold189 (.A(\project_audio.freq[3][4] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold190 (.A(\project_audio.iter.mult1_shift[28] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0203_),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold192 (.A(\project_audio.freq[4][7] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold193 (.A(\project_audio.iter.mult_accum[0] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold194 (.A(_1414_),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0206_),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold196 (.A(\project_audio.freq[7][3] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold197 (.A(\project_audio.freq[6][1] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold198 (.A(\project_audio.iter.mult_accum[2] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0208_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold200 (.A(\project_audio.freq[7][5] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold201 (.A(\project_audio.iter.mult_accum[14] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold202 (.A(\project_audio.freq[6][9] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold203 (.A(\hpos[3] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold204 (.A(_1026_),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold205 (.A(\sync_gen.vpos[9] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold206 (.A(_1322_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold207 (.A(\project_audio.freq[0][4] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold208 (.A(\project_audio.freq[4][10] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold209 (.A(\project_audio.iter.mult1_shift[23] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0198_),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold211 (.A(\hpos[6] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0103_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold213 (.A(\project_audio.freq[4][9] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold214 (.A(\project_audio.freq[2][9] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold215 (.A(\project_audio.freq[1][9] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0460_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold217 (.A(\project_audio.nco_increment_gen.counter[8] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0142_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold219 (.A(\project_audio.freq[7][6] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold220 (.A(\project_audio.freq[5][9] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold221 (.A(\project_audio.freq[3][3] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold222 (.A(\project_audio.freq[0][10] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold223 (.A(\project_audio.iter.mult2_shift[8] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold224 (.A(_2237_),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0382_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold226 (.A(\project_audio.freq[0][9] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold227 (.A(\project_audio.genblk1[5].n_c_oh_my.snd ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold228 (.A(\project_audio.iter.mult_accum[8] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold229 (.A(\project_audio.iter.mult_accum[5] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0211_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold231 (.A(\project_audio.iter.counter[9] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold232 (.A(_2362_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold233 (.A(\project_audio.freq[3][9] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold234 (.A(\project_audio.freq[3][6] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold235 (.A(\project_audio.iter.mult2_shift[2] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold236 (.A(_2214_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0376_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0006_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold239 (.A(_2395_),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0434_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold241 (.A(\project_audio.freq[7][9] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold242 (.A(\project_audio.iter.mult1_shift[24] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0199_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold244 (.A(\project_audio.iter.mult_accum[10] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold245 (.A(\project_audio.iter.mult2_shift[4] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold246 (.A(_2222_),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0378_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold248 (.A(\project_audio.iter.x[3] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0401_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0010_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold251 (.A(_1029_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold252 (.A(\project_audio.nco_increment_gen.counter[5] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold253 (.A(\project_audio.iter.mult2_shift[15] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0388_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold255 (.A(\project_audio.mixer.counter[1] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0392_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold257 (.A(\project_audio.iter.mult1_shift[26] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0201_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold259 (.A(\project_audio.iter.mult2_shift[12] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold260 (.A(_2253_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0386_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold262 (.A(\project_audio.iter.mult2_shift[11] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold263 (.A(_2249_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0385_),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold265 (.A(\project_audio.mixer.counter[2] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold266 (.A(_2317_),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0393_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold268 (.A(\project_audio.iter.mult2_shift[10] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0383_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold270 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[5] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold271 (.A(\project_audio.iter.r[1] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold272 (.A(_2386_),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold273 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[0] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold274 (.A(\project_audio.iter.mult2_shift[1] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold275 (.A(_2211_),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0375_),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold277 (.A(\project_audio.iter.mult1_shift[19] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0194_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold279 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[12] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold280 (.A(_2201_),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold281 (.A(\project_audio.iter.mult1_shift[22] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold282 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[0] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold283 (.A(\project_audio.iter.mult2_shift[6] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold284 (.A(_2230_),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0380_),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold286 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[5] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold287 (.A(\project_audio.iter.mult2_shift[5] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold288 (.A(_2226_),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0379_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold290 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[0] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold291 (.A(\project_audio.iter.mult_accum[26] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0384_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold293 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[5] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold294 (.A(\project_audio.iter.r[8] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold295 (.A(_2406_),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold296 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[5] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold297 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[0] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold298 (.A(\project_audio.genblk1[7].n_c_oh_my.snd ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold299 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[0] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold300 (.A(\hpos[2] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold301 (.A(_1024_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold302 (.A(\project_audio.iter.mult1_shift[2] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0048_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold304 (.A(\project_audio.iter.mult2_shift[7] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold305 (.A(_2234_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0381_),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold307 (.A(\sync_gen.vpos[4] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold308 (.A(_1310_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold309 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[0] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold310 (.A(\hpos[4] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold311 (.A(_1027_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold312 (.A(\project_audio.iter.mult2_shift[13] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold313 (.A(_2257_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0387_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold315 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[11] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0267_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold317 (.A(\project_audio.iter.mult1_shift[25] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold318 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[5] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold319 (.A(\hpos[9] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold320 (.A(_1038_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold321 (.A(\project_audio.iter.mult1_shift[26] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold322 (.A(_1592_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold323 (.A(\project_audio.iter.mult1_shift[27] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold324 (.A(\project_audio.iter.mult2_shift[3] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold325 (.A(_2218_),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0377_),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold327 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[0] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold328 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[5] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold329 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[11] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0301_),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold331 (.A(\project_audio.iter.mult_accum[9] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0215_),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold333 (.A(\project_audio.iter.mult_accum[11] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold334 (.A(\project_audio.iter.counter[2] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold335 (.A(_2349_),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold336 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[11] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0318_),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold338 (.A(\project_audio.iter.mult1_shift[21] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold339 (.A(\project_audio.iter.mult_accum[30] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0236_),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold341 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[3] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold342 (.A(\project_audio.iter.mult_accum[13] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold343 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[11] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0335_),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold345 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[8] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0281_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold347 (.A(\project_audio.genblk1[6].n_c_oh_my.snd ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold348 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[0] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold349 (.A(\project_audio.iter.mult1_shift[17] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0397_),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold351 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[3] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0361_),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold353 (.A(\project_audio.nco_increment_gen.counter[0] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0135_),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold355 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[11] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0352_),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold357 (.A(\project_audio.genblk1[4].n_c_oh_my.snd ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold358 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[6] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold359 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[11] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0250_),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold361 (.A(\project_audio.iter.counter[8] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold362 (.A(_2360_),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold363 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[10] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0266_),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold365 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[2] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0275_),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold367 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[1] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold368 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[10] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0334_),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold370 (.A(\project_audio.genblk1[2].n_c_oh_my.snd ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold371 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[2] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0241_),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold373 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[8] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0349_),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold375 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[2] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0343_),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold377 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[2] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0292_),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold379 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[7] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0246_),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold381 (.A(\project_audio.genblk1[1].n_c_oh_my.snd ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold382 (.A(\project_audio.iter.mult_accum[12] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold383 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[8] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0366_),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold385 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[8] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0298_),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold387 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[8] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0332_),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold389 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[6] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold390 (.A(\project_audio.iter.r[11] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold391 (.A(_2412_),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0441_),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold393 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[4] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0328_),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold395 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[3] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold396 (.A(\project_audio.iter.mult_accum[24] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold397 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[5] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold398 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[10] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0317_),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold400 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[7] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0348_),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold402 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[6] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0347_),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold404 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[1] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold405 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[8] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0315_),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold407 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[10] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0249_),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold409 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[3] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0276_),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold411 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[1] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0342_),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold413 (.A(\project_audio.iter.mult1_shift[20] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold414 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[1] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold415 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[6] ),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0313_),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold417 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[4] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0277_),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold419 (.A(\project_audio.genblk1[3].n_c_oh_my.snd ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold420 (.A(\project_audio.iter.mult_accum[31] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold421 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[2] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold422 (.A(_0309_),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold423 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[3] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold424 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[4] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0294_),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold426 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[4] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0362_),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold428 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[10] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0283_),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold430 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[3] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold431 (.A(_0242_),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold432 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[7] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold433 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[4] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0311_),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold435 (.A(\project_audio.iter.mult1_shift[1] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold436 (.A(\project_audio.iter.counter[6] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold437 (.A(_2356_),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold438 (.A(\project_audio.iter.counter[11] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold439 (.A(_2366_),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold440 (.A(\project_audio.iter.counter[7] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold441 (.A(\hpos[7] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold442 (.A(_1034_),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold443 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[2] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0360_),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold445 (.A(\project_audio.iter.mult1_shift[30] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0204_),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold447 (.A(\project_audio.iter.mult1_shift[11] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0056_),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold449 (.A(\project_audio.iter.r[6] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0051_),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold451 (.A(\project_audio.iter.counter[12] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold452 (.A(\project_audio.iter.mult1_shift[18] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold453 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[11] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0284_),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold455 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[7] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold456 (.A(\project_audio.iter.counter[10] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold457 (.A(\hpos[8] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold458 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[4] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold459 (.A(_0243_),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0003_),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold461 (.A(_2438_),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold462 (.A(_0450_),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold463 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[10] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0351_),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold465 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[7] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0365_),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold467 (.A(\project_audio.iter.mult1_shift[7] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0053_),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold469 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[3] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold470 (.A(\project_audio.iter.mult1_shift[4] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0049_),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold472 (.A(\project_audio.iter.mult_accum[16] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0374_),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold474 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[10] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0300_),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold476 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[8] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold477 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[1] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold478 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[4] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0260_),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold480 (.A(\project_audio.iter.counter[3] ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold481 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[6] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold482 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[2] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0258_),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold484 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[7] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold485 (.A(_0280_),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold486 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[1] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold487 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[1] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold488 (.A(\project_audio.iter.counter[5] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold489 (.A(_2354_),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold490 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[2] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold491 (.A(_0326_),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold492 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[3] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0259_),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold494 (.A(\sync_gen.vpos[2] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold495 (.A(_1307_),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold496 (.A(\project_audio.iter.mult_accum[29] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0235_),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold498 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[4] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0345_),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold500 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[6] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0330_),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold502 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[7] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0263_),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold504 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[9] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold505 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[6] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold506 (.A(_0245_),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold507 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[1] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold508 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[7] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold509 (.A(\project_audio.iter.mult1_shift[0] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold510 (.A(_2545_),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0045_),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold512 (.A(_0018_),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold513 (.A(_0118_),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold514 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[11] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold515 (.A(_0369_),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold516 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[9] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold517 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[10] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold518 (.A(_0368_),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold519 (.A(\project_audio.f_counter[0] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold520 (.A(_2435_),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold521 (.A(_0449_),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold522 (.A(\project_audio.iter.r[17] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold523 (.A(_2421_),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold524 (.A(_0447_),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold525 (.A(\project_audio.iter.mult1_shift[8] ),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0054_),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold527 (.A(\project_audio.iter.r[7] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0052_),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold529 (.A(\project_audio.iter.r[15] ),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold530 (.A(_2418_),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0445_),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold532 (.A(\project_audio.iter.mult1_shift[5] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0050_),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold534 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[6] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold535 (.A(_0262_),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold536 (.A(\project_audio.iter.mult_accum[28] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold537 (.A(\project_audio.iter.mult1_shift[12] ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold538 (.A(_0057_),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold539 (.A(\project_audio.genblk1[6].n_c_oh_my.phase[8] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold540 (.A(\project_audio.iter.r[13] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold541 (.A(_2415_),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold542 (.A(\project_audio.iter.r[10] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold543 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[9] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0333_),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold545 (.A(\project_audio.iter.r[4] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0437_),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold547 (.A(\project_audio.genblk1[5].n_c_oh_my.phase[9] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold548 (.A(\project_audio.iter.x[7] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold549 (.A(_0405_),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold550 (.A(\project_audio.genblk1[4].n_c_oh_my.phase[9] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold551 (.A(\project_audio.iter.counter[4] ),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold552 (.A(\project_audio.iter.mult_accum[22] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold553 (.A(\hpos[4] ),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold554 (.A(_0132_),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold555 (.A(\project_audio.genblk1[3].n_c_oh_my.phase[9] ),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold556 (.A(\project_audio.iter.r[5] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold557 (.A(\project_audio.iter.mult1_shift[10] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold558 (.A(_0055_),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold559 (.A(\project_audio.iter.mult_accum[23] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold560 (.A(\project_audio.iter.mult1_shift[15] ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0060_),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold562 (.A(\project_audio.iter.x[12] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold563 (.A(\project_audio.iter.mult1_shift[13] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold564 (.A(\project_audio.genblk1[7].n_c_oh_my.phase[5] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold565 (.A(_0244_),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold566 (.A(\project_audio.iter.mult_accum[18] ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold567 (.A(\project_audio.iter.mult_accum[21] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold568 (.A(\project_audio.genblk1[1].n_c_oh_my.phase[9] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold569 (.A(_0350_),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold570 (.A(\project_audio.genblk1[0].n_c_oh_my.phase[9] ),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold571 (.A(\project_audio.iter.mult_accum[27] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold572 (.A(\project_audio.iter.next_ready ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0448_),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold574 (.A(\project_audio.iter.mult_accum[25] ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold575 (.A(\project_audio.iter.mult_accum[19] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold576 (.A(\project_audio.iter.x[8] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold577 (.A(\sync_gen.vpos[5] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold578 (.A(_1315_),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold579 (.A(\project_audio.iter.mult1_shift[16] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold580 (.A(\project_audio.iter.mult1_shift[14] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold581 (.A(_0059_),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold582 (.A(\project_audio.iter.x[14] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold583 (.A(\project_audio.iter.r[14] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold584 (.A(\project_audio.iter.mult_accum[17] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold585 (.A(\sync_gen.vpos[0] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold586 (.A(_1303_),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold587 (.A(_0122_),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold588 (.A(\project_audio.iter.x[15] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold589 (.A(\project_audio.iter.x[13] ),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold590 (.A(\project_audio.iter.x[10] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold591 (.A(\sync_gen.vpos[7] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold592 (.A(_1319_),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold593 (.A(\project_audio.iter.r[9] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold594 (.A(\project_audio.iter.x[11] ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold595 (.A(\project_audio.iter.mult_accum[20] ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold596 (.A(\frame_no[3] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold597 (.A(_0114_),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold598 (.A(\hpos[1] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold599 (.A(_1023_),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold600 (.A(_0098_),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold601 (.A(\project_audio.iter.counter[0] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold602 (.A(_2347_),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold603 (.A(_0416_),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold604 (.A(\project_audio.mixer.counter[1] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold605 (.A(_2313_),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold606 (.A(\project_audio.iter.r[16] ),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold607 (.A(_0446_),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold608 (.A(\project_audio.iter.x[9] ),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold609 (.A(\project_audio.iter.x[0] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold610 (.A(\sync_gen.vpos[3] ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold611 (.A(\frame_no[1] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold612 (.A(_1282_),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold613 (.A(\project_audio.iter.x[1] ),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold614 (.A(\project_audio.iter.x[2] ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold615 (.A(\sync_gen.vpos[6] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold616 (.A(_1040_),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold617 (.A(_0133_),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold618 (.A(\sync_gen.vpos[8] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold619 (.A(\project_audio.iter.x[6] ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold620 (.A(\project_audio.iter.r[12] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold621 (.A(_2414_),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold622 (.A(\frame_no[5] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold623 (.A(_0116_),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold624 (.A(\project_audio.iter.x[4] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold625 (.A(\sync_gen.vpos[1] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold626 (.A(prev_vsync),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold627 (.A(_0113_),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold628 (.A(\project_audio.iter.x[5] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold629 (.A(\frame_no[6] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold630 (.A(\project_audio.iter.mult1_shift[4] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold631 (.A(_1437_),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold632 (.A(\project_audio.iter.mult1_shift[12] ),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold633 (.A(\project_audio.genblk1[2].n_c_oh_my.phase[2] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold634 (.A(\project_audio.iter.mult_accum[2] ),
    .X(net1244));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_fill_1 FILLER_13_52 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_fill_1 FILLER_13_77 ();
 sg13g2_fill_2 FILLER_13_82 ();
 sg13g2_decap_8 FILLER_13_88 ();
 sg13g2_decap_4 FILLER_13_95 ();
 sg13g2_fill_2 FILLER_13_99 ();
 sg13g2_fill_1 FILLER_13_109 ();
 sg13g2_decap_4 FILLER_13_119 ();
 sg13g2_fill_1 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_132 ();
 sg13g2_decap_8 FILLER_13_139 ();
 sg13g2_decap_8 FILLER_13_146 ();
 sg13g2_decap_8 FILLER_13_153 ();
 sg13g2_decap_8 FILLER_13_160 ();
 sg13g2_decap_8 FILLER_13_167 ();
 sg13g2_decap_8 FILLER_13_174 ();
 sg13g2_decap_8 FILLER_13_181 ();
 sg13g2_decap_8 FILLER_13_188 ();
 sg13g2_decap_4 FILLER_13_195 ();
 sg13g2_fill_1 FILLER_13_199 ();
 sg13g2_decap_8 FILLER_13_204 ();
 sg13g2_decap_8 FILLER_13_211 ();
 sg13g2_decap_8 FILLER_13_218 ();
 sg13g2_decap_8 FILLER_13_225 ();
 sg13g2_decap_8 FILLER_13_232 ();
 sg13g2_decap_8 FILLER_13_239 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_250 ();
 sg13g2_decap_8 FILLER_13_254 ();
 sg13g2_decap_8 FILLER_13_261 ();
 sg13g2_decap_8 FILLER_13_268 ();
 sg13g2_decap_8 FILLER_13_275 ();
 sg13g2_decap_8 FILLER_13_282 ();
 sg13g2_decap_8 FILLER_13_289 ();
 sg13g2_decap_8 FILLER_13_296 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_decap_8 FILLER_13_310 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_352 ();
 sg13g2_fill_1 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_4 FILLER_13_385 ();
 sg13g2_fill_2 FILLER_13_389 ();
 sg13g2_fill_2 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_13_412 ();
 sg13g2_decap_8 FILLER_13_419 ();
 sg13g2_decap_8 FILLER_13_426 ();
 sg13g2_decap_8 FILLER_13_433 ();
 sg13g2_decap_8 FILLER_13_440 ();
 sg13g2_decap_8 FILLER_13_447 ();
 sg13g2_decap_8 FILLER_13_454 ();
 sg13g2_decap_8 FILLER_13_461 ();
 sg13g2_decap_8 FILLER_13_468 ();
 sg13g2_decap_8 FILLER_13_475 ();
 sg13g2_decap_8 FILLER_13_482 ();
 sg13g2_decap_8 FILLER_13_489 ();
 sg13g2_decap_8 FILLER_13_496 ();
 sg13g2_decap_8 FILLER_13_503 ();
 sg13g2_decap_8 FILLER_13_510 ();
 sg13g2_decap_8 FILLER_13_517 ();
 sg13g2_decap_8 FILLER_13_524 ();
 sg13g2_decap_8 FILLER_13_531 ();
 sg13g2_decap_8 FILLER_13_538 ();
 sg13g2_decap_8 FILLER_13_545 ();
 sg13g2_decap_8 FILLER_13_552 ();
 sg13g2_decap_8 FILLER_13_559 ();
 sg13g2_decap_8 FILLER_13_566 ();
 sg13g2_decap_8 FILLER_13_573 ();
 sg13g2_decap_8 FILLER_13_580 ();
 sg13g2_decap_8 FILLER_13_587 ();
 sg13g2_decap_8 FILLER_13_594 ();
 sg13g2_decap_8 FILLER_13_601 ();
 sg13g2_decap_8 FILLER_13_608 ();
 sg13g2_decap_8 FILLER_13_615 ();
 sg13g2_decap_8 FILLER_13_622 ();
 sg13g2_decap_8 FILLER_13_629 ();
 sg13g2_decap_8 FILLER_13_636 ();
 sg13g2_decap_8 FILLER_13_643 ();
 sg13g2_decap_8 FILLER_13_650 ();
 sg13g2_decap_8 FILLER_13_657 ();
 sg13g2_decap_8 FILLER_13_664 ();
 sg13g2_decap_8 FILLER_13_671 ();
 sg13g2_decap_8 FILLER_13_678 ();
 sg13g2_decap_8 FILLER_13_685 ();
 sg13g2_decap_8 FILLER_13_692 ();
 sg13g2_decap_8 FILLER_13_699 ();
 sg13g2_decap_8 FILLER_13_706 ();
 sg13g2_decap_8 FILLER_13_713 ();
 sg13g2_decap_8 FILLER_13_720 ();
 sg13g2_decap_8 FILLER_13_727 ();
 sg13g2_decap_8 FILLER_13_734 ();
 sg13g2_decap_8 FILLER_13_741 ();
 sg13g2_decap_8 FILLER_13_748 ();
 sg13g2_decap_8 FILLER_13_755 ();
 sg13g2_decap_8 FILLER_13_762 ();
 sg13g2_decap_8 FILLER_13_769 ();
 sg13g2_decap_8 FILLER_13_776 ();
 sg13g2_decap_8 FILLER_13_783 ();
 sg13g2_decap_8 FILLER_13_790 ();
 sg13g2_decap_8 FILLER_13_797 ();
 sg13g2_decap_8 FILLER_13_804 ();
 sg13g2_decap_8 FILLER_13_811 ();
 sg13g2_decap_8 FILLER_13_818 ();
 sg13g2_decap_8 FILLER_13_825 ();
 sg13g2_decap_8 FILLER_13_832 ();
 sg13g2_decap_8 FILLER_13_839 ();
 sg13g2_decap_8 FILLER_13_846 ();
 sg13g2_decap_8 FILLER_13_853 ();
 sg13g2_fill_2 FILLER_13_860 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_4 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_29 ();
 sg13g2_fill_1 FILLER_14_31 ();
 sg13g2_fill_2 FILLER_14_115 ();
 sg13g2_fill_1 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_fill_2 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_174 ();
 sg13g2_fill_2 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_181 ();
 sg13g2_decap_4 FILLER_14_216 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_232 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_fill_1 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_302 ();
 sg13g2_decap_8 FILLER_14_309 ();
 sg13g2_decap_8 FILLER_14_316 ();
 sg13g2_decap_8 FILLER_14_323 ();
 sg13g2_decap_8 FILLER_14_330 ();
 sg13g2_decap_8 FILLER_14_337 ();
 sg13g2_decap_8 FILLER_14_344 ();
 sg13g2_fill_2 FILLER_14_351 ();
 sg13g2_fill_2 FILLER_14_359 ();
 sg13g2_fill_2 FILLER_14_365 ();
 sg13g2_fill_1 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_4 FILLER_14_380 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_411 ();
 sg13g2_decap_4 FILLER_14_418 ();
 sg13g2_decap_8 FILLER_14_433 ();
 sg13g2_decap_8 FILLER_14_444 ();
 sg13g2_decap_8 FILLER_14_451 ();
 sg13g2_decap_8 FILLER_14_458 ();
 sg13g2_decap_8 FILLER_14_465 ();
 sg13g2_decap_8 FILLER_14_472 ();
 sg13g2_decap_8 FILLER_14_479 ();
 sg13g2_decap_8 FILLER_14_486 ();
 sg13g2_decap_8 FILLER_14_493 ();
 sg13g2_decap_8 FILLER_14_500 ();
 sg13g2_decap_8 FILLER_14_507 ();
 sg13g2_decap_8 FILLER_14_514 ();
 sg13g2_decap_8 FILLER_14_521 ();
 sg13g2_decap_8 FILLER_14_528 ();
 sg13g2_decap_8 FILLER_14_535 ();
 sg13g2_decap_8 FILLER_14_542 ();
 sg13g2_decap_8 FILLER_14_549 ();
 sg13g2_decap_8 FILLER_14_556 ();
 sg13g2_decap_8 FILLER_14_563 ();
 sg13g2_decap_8 FILLER_14_570 ();
 sg13g2_decap_8 FILLER_14_577 ();
 sg13g2_decap_8 FILLER_14_584 ();
 sg13g2_decap_8 FILLER_14_591 ();
 sg13g2_decap_8 FILLER_14_598 ();
 sg13g2_decap_8 FILLER_14_605 ();
 sg13g2_decap_8 FILLER_14_612 ();
 sg13g2_decap_8 FILLER_14_619 ();
 sg13g2_decap_8 FILLER_14_626 ();
 sg13g2_decap_8 FILLER_14_633 ();
 sg13g2_decap_8 FILLER_14_640 ();
 sg13g2_decap_8 FILLER_14_647 ();
 sg13g2_decap_8 FILLER_14_654 ();
 sg13g2_decap_8 FILLER_14_661 ();
 sg13g2_decap_8 FILLER_14_668 ();
 sg13g2_decap_8 FILLER_14_675 ();
 sg13g2_decap_8 FILLER_14_682 ();
 sg13g2_decap_8 FILLER_14_689 ();
 sg13g2_decap_8 FILLER_14_696 ();
 sg13g2_decap_8 FILLER_14_703 ();
 sg13g2_decap_8 FILLER_14_710 ();
 sg13g2_decap_8 FILLER_14_717 ();
 sg13g2_decap_8 FILLER_14_724 ();
 sg13g2_decap_8 FILLER_14_731 ();
 sg13g2_decap_8 FILLER_14_738 ();
 sg13g2_decap_8 FILLER_14_745 ();
 sg13g2_decap_8 FILLER_14_752 ();
 sg13g2_decap_8 FILLER_14_759 ();
 sg13g2_decap_8 FILLER_14_766 ();
 sg13g2_decap_8 FILLER_14_773 ();
 sg13g2_decap_8 FILLER_14_780 ();
 sg13g2_decap_8 FILLER_14_787 ();
 sg13g2_decap_8 FILLER_14_794 ();
 sg13g2_decap_8 FILLER_14_801 ();
 sg13g2_decap_8 FILLER_14_808 ();
 sg13g2_decap_8 FILLER_14_815 ();
 sg13g2_decap_8 FILLER_14_822 ();
 sg13g2_decap_8 FILLER_14_829 ();
 sg13g2_decap_8 FILLER_14_836 ();
 sg13g2_decap_8 FILLER_14_843 ();
 sg13g2_decap_8 FILLER_14_850 ();
 sg13g2_decap_4 FILLER_14_857 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_40 ();
 sg13g2_fill_2 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_fill_2 FILLER_15_162 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_fill_2 FILLER_15_238 ();
 sg13g2_fill_2 FILLER_15_259 ();
 sg13g2_fill_1 FILLER_15_279 ();
 sg13g2_fill_1 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_331 ();
 sg13g2_decap_8 FILLER_15_338 ();
 sg13g2_decap_4 FILLER_15_345 ();
 sg13g2_fill_1 FILLER_15_349 ();
 sg13g2_fill_2 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_fill_1 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_435 ();
 sg13g2_decap_8 FILLER_15_464 ();
 sg13g2_decap_4 FILLER_15_471 ();
 sg13g2_fill_1 FILLER_15_475 ();
 sg13g2_decap_8 FILLER_15_486 ();
 sg13g2_decap_8 FILLER_15_493 ();
 sg13g2_decap_8 FILLER_15_500 ();
 sg13g2_decap_8 FILLER_15_507 ();
 sg13g2_decap_8 FILLER_15_514 ();
 sg13g2_decap_8 FILLER_15_521 ();
 sg13g2_decap_8 FILLER_15_528 ();
 sg13g2_decap_8 FILLER_15_535 ();
 sg13g2_decap_8 FILLER_15_542 ();
 sg13g2_decap_8 FILLER_15_549 ();
 sg13g2_decap_8 FILLER_15_556 ();
 sg13g2_decap_8 FILLER_15_563 ();
 sg13g2_decap_8 FILLER_15_570 ();
 sg13g2_decap_8 FILLER_15_577 ();
 sg13g2_decap_8 FILLER_15_584 ();
 sg13g2_decap_8 FILLER_15_591 ();
 sg13g2_decap_8 FILLER_15_598 ();
 sg13g2_decap_8 FILLER_15_605 ();
 sg13g2_decap_8 FILLER_15_612 ();
 sg13g2_decap_8 FILLER_15_619 ();
 sg13g2_decap_8 FILLER_15_626 ();
 sg13g2_decap_8 FILLER_15_633 ();
 sg13g2_decap_8 FILLER_15_640 ();
 sg13g2_decap_8 FILLER_15_647 ();
 sg13g2_decap_8 FILLER_15_654 ();
 sg13g2_decap_8 FILLER_15_661 ();
 sg13g2_decap_8 FILLER_15_668 ();
 sg13g2_decap_8 FILLER_15_675 ();
 sg13g2_decap_8 FILLER_15_682 ();
 sg13g2_decap_8 FILLER_15_689 ();
 sg13g2_decap_8 FILLER_15_696 ();
 sg13g2_decap_8 FILLER_15_703 ();
 sg13g2_decap_8 FILLER_15_710 ();
 sg13g2_decap_8 FILLER_15_717 ();
 sg13g2_decap_8 FILLER_15_724 ();
 sg13g2_decap_8 FILLER_15_731 ();
 sg13g2_decap_8 FILLER_15_738 ();
 sg13g2_decap_8 FILLER_15_745 ();
 sg13g2_decap_8 FILLER_15_752 ();
 sg13g2_decap_8 FILLER_15_759 ();
 sg13g2_decap_8 FILLER_15_766 ();
 sg13g2_decap_8 FILLER_15_773 ();
 sg13g2_decap_8 FILLER_15_780 ();
 sg13g2_decap_8 FILLER_15_787 ();
 sg13g2_decap_8 FILLER_15_794 ();
 sg13g2_decap_8 FILLER_15_801 ();
 sg13g2_decap_8 FILLER_15_808 ();
 sg13g2_decap_8 FILLER_15_815 ();
 sg13g2_decap_8 FILLER_15_822 ();
 sg13g2_decap_8 FILLER_15_829 ();
 sg13g2_decap_8 FILLER_15_836 ();
 sg13g2_decap_8 FILLER_15_843 ();
 sg13g2_decap_8 FILLER_15_850 ();
 sg13g2_decap_4 FILLER_15_857 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_4 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_53 ();
 sg13g2_fill_1 FILLER_16_55 ();
 sg13g2_fill_2 FILLER_16_83 ();
 sg13g2_fill_1 FILLER_16_85 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_171 ();
 sg13g2_fill_1 FILLER_16_173 ();
 sg13g2_fill_2 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_fill_1 FILLER_16_234 ();
 sg13g2_fill_2 FILLER_16_249 ();
 sg13g2_fill_2 FILLER_16_278 ();
 sg13g2_fill_1 FILLER_16_292 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_fill_2 FILLER_16_349 ();
 sg13g2_decap_4 FILLER_16_359 ();
 sg13g2_fill_1 FILLER_16_373 ();
 sg13g2_fill_2 FILLER_16_383 ();
 sg13g2_fill_2 FILLER_16_395 ();
 sg13g2_fill_2 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_403 ();
 sg13g2_fill_1 FILLER_16_414 ();
 sg13g2_decap_8 FILLER_16_423 ();
 sg13g2_decap_8 FILLER_16_430 ();
 sg13g2_decap_4 FILLER_16_437 ();
 sg13g2_fill_1 FILLER_16_441 ();
 sg13g2_fill_2 FILLER_16_450 ();
 sg13g2_fill_2 FILLER_16_456 ();
 sg13g2_fill_1 FILLER_16_458 ();
 sg13g2_fill_1 FILLER_16_471 ();
 sg13g2_decap_8 FILLER_16_491 ();
 sg13g2_decap_8 FILLER_16_498 ();
 sg13g2_decap_8 FILLER_16_505 ();
 sg13g2_decap_8 FILLER_16_512 ();
 sg13g2_decap_8 FILLER_16_519 ();
 sg13g2_decap_8 FILLER_16_526 ();
 sg13g2_decap_8 FILLER_16_533 ();
 sg13g2_decap_8 FILLER_16_540 ();
 sg13g2_decap_8 FILLER_16_547 ();
 sg13g2_decap_8 FILLER_16_554 ();
 sg13g2_decap_8 FILLER_16_561 ();
 sg13g2_decap_8 FILLER_16_568 ();
 sg13g2_decap_8 FILLER_16_575 ();
 sg13g2_decap_8 FILLER_16_582 ();
 sg13g2_decap_8 FILLER_16_589 ();
 sg13g2_decap_8 FILLER_16_596 ();
 sg13g2_decap_8 FILLER_16_603 ();
 sg13g2_decap_8 FILLER_16_610 ();
 sg13g2_decap_8 FILLER_16_617 ();
 sg13g2_decap_8 FILLER_16_624 ();
 sg13g2_decap_8 FILLER_16_631 ();
 sg13g2_decap_8 FILLER_16_638 ();
 sg13g2_decap_8 FILLER_16_645 ();
 sg13g2_decap_8 FILLER_16_652 ();
 sg13g2_decap_8 FILLER_16_659 ();
 sg13g2_decap_8 FILLER_16_666 ();
 sg13g2_decap_8 FILLER_16_673 ();
 sg13g2_decap_8 FILLER_16_680 ();
 sg13g2_decap_8 FILLER_16_687 ();
 sg13g2_decap_8 FILLER_16_694 ();
 sg13g2_decap_8 FILLER_16_701 ();
 sg13g2_decap_8 FILLER_16_708 ();
 sg13g2_decap_8 FILLER_16_715 ();
 sg13g2_decap_8 FILLER_16_722 ();
 sg13g2_decap_8 FILLER_16_729 ();
 sg13g2_decap_8 FILLER_16_736 ();
 sg13g2_decap_8 FILLER_16_743 ();
 sg13g2_decap_8 FILLER_16_750 ();
 sg13g2_decap_8 FILLER_16_757 ();
 sg13g2_decap_8 FILLER_16_764 ();
 sg13g2_decap_8 FILLER_16_771 ();
 sg13g2_decap_8 FILLER_16_778 ();
 sg13g2_decap_8 FILLER_16_785 ();
 sg13g2_decap_8 FILLER_16_792 ();
 sg13g2_decap_8 FILLER_16_799 ();
 sg13g2_decap_8 FILLER_16_806 ();
 sg13g2_decap_8 FILLER_16_813 ();
 sg13g2_decap_8 FILLER_16_820 ();
 sg13g2_decap_8 FILLER_16_827 ();
 sg13g2_decap_8 FILLER_16_834 ();
 sg13g2_decap_8 FILLER_16_841 ();
 sg13g2_decap_8 FILLER_16_848 ();
 sg13g2_decap_8 FILLER_16_855 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_11 ();
 sg13g2_fill_2 FILLER_17_38 ();
 sg13g2_fill_1 FILLER_17_114 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_fill_2 FILLER_17_196 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_1 FILLER_17_209 ();
 sg13g2_fill_2 FILLER_17_216 ();
 sg13g2_fill_2 FILLER_17_223 ();
 sg13g2_fill_1 FILLER_17_225 ();
 sg13g2_fill_1 FILLER_17_252 ();
 sg13g2_fill_2 FILLER_17_257 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_decap_4 FILLER_17_341 ();
 sg13g2_fill_2 FILLER_17_359 ();
 sg13g2_fill_2 FILLER_17_380 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_fill_1 FILLER_17_409 ();
 sg13g2_fill_1 FILLER_17_414 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_1 FILLER_17_427 ();
 sg13g2_fill_2 FILLER_17_436 ();
 sg13g2_fill_1 FILLER_17_451 ();
 sg13g2_decap_8 FILLER_17_457 ();
 sg13g2_fill_2 FILLER_17_464 ();
 sg13g2_fill_2 FILLER_17_480 ();
 sg13g2_decap_8 FILLER_17_491 ();
 sg13g2_decap_8 FILLER_17_498 ();
 sg13g2_decap_8 FILLER_17_505 ();
 sg13g2_decap_8 FILLER_17_512 ();
 sg13g2_decap_8 FILLER_17_519 ();
 sg13g2_decap_8 FILLER_17_526 ();
 sg13g2_decap_8 FILLER_17_533 ();
 sg13g2_decap_8 FILLER_17_540 ();
 sg13g2_decap_8 FILLER_17_547 ();
 sg13g2_decap_8 FILLER_17_554 ();
 sg13g2_decap_8 FILLER_17_561 ();
 sg13g2_decap_8 FILLER_17_568 ();
 sg13g2_decap_8 FILLER_17_575 ();
 sg13g2_decap_8 FILLER_17_582 ();
 sg13g2_decap_8 FILLER_17_589 ();
 sg13g2_decap_8 FILLER_17_596 ();
 sg13g2_decap_8 FILLER_17_603 ();
 sg13g2_decap_8 FILLER_17_610 ();
 sg13g2_decap_8 FILLER_17_617 ();
 sg13g2_decap_8 FILLER_17_624 ();
 sg13g2_decap_8 FILLER_17_631 ();
 sg13g2_decap_8 FILLER_17_638 ();
 sg13g2_decap_8 FILLER_17_645 ();
 sg13g2_decap_8 FILLER_17_652 ();
 sg13g2_decap_8 FILLER_17_659 ();
 sg13g2_decap_8 FILLER_17_666 ();
 sg13g2_decap_8 FILLER_17_673 ();
 sg13g2_decap_8 FILLER_17_680 ();
 sg13g2_decap_8 FILLER_17_687 ();
 sg13g2_decap_8 FILLER_17_694 ();
 sg13g2_decap_8 FILLER_17_701 ();
 sg13g2_decap_8 FILLER_17_708 ();
 sg13g2_decap_8 FILLER_17_715 ();
 sg13g2_decap_8 FILLER_17_722 ();
 sg13g2_decap_8 FILLER_17_729 ();
 sg13g2_decap_8 FILLER_17_736 ();
 sg13g2_decap_8 FILLER_17_743 ();
 sg13g2_decap_8 FILLER_17_750 ();
 sg13g2_decap_8 FILLER_17_757 ();
 sg13g2_decap_8 FILLER_17_764 ();
 sg13g2_decap_8 FILLER_17_771 ();
 sg13g2_decap_8 FILLER_17_778 ();
 sg13g2_decap_8 FILLER_17_785 ();
 sg13g2_decap_8 FILLER_17_792 ();
 sg13g2_decap_8 FILLER_17_799 ();
 sg13g2_decap_8 FILLER_17_806 ();
 sg13g2_decap_8 FILLER_17_813 ();
 sg13g2_decap_8 FILLER_17_820 ();
 sg13g2_decap_8 FILLER_17_827 ();
 sg13g2_decap_8 FILLER_17_834 ();
 sg13g2_decap_8 FILLER_17_841 ();
 sg13g2_decap_8 FILLER_17_848 ();
 sg13g2_decap_8 FILLER_17_855 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_27 ();
 sg13g2_fill_1 FILLER_18_29 ();
 sg13g2_fill_1 FILLER_18_55 ();
 sg13g2_fill_2 FILLER_18_102 ();
 sg13g2_fill_1 FILLER_18_104 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_fill_1 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_153 ();
 sg13g2_decap_4 FILLER_18_160 ();
 sg13g2_fill_2 FILLER_18_164 ();
 sg13g2_decap_8 FILLER_18_170 ();
 sg13g2_fill_2 FILLER_18_177 ();
 sg13g2_fill_1 FILLER_18_179 ();
 sg13g2_fill_2 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_229 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_241 ();
 sg13g2_decap_8 FILLER_18_268 ();
 sg13g2_fill_2 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_291 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_decap_4 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_fill_2 FILLER_18_400 ();
 sg13g2_fill_1 FILLER_18_417 ();
 sg13g2_fill_2 FILLER_18_426 ();
 sg13g2_fill_1 FILLER_18_428 ();
 sg13g2_fill_1 FILLER_18_453 ();
 sg13g2_fill_1 FILLER_18_462 ();
 sg13g2_fill_2 FILLER_18_467 ();
 sg13g2_fill_2 FILLER_18_473 ();
 sg13g2_fill_1 FILLER_18_475 ();
 sg13g2_decap_8 FILLER_18_498 ();
 sg13g2_decap_8 FILLER_18_505 ();
 sg13g2_decap_8 FILLER_18_512 ();
 sg13g2_decap_8 FILLER_18_519 ();
 sg13g2_decap_8 FILLER_18_526 ();
 sg13g2_decap_8 FILLER_18_533 ();
 sg13g2_decap_8 FILLER_18_540 ();
 sg13g2_decap_8 FILLER_18_547 ();
 sg13g2_decap_8 FILLER_18_554 ();
 sg13g2_decap_8 FILLER_18_561 ();
 sg13g2_decap_8 FILLER_18_568 ();
 sg13g2_decap_8 FILLER_18_575 ();
 sg13g2_decap_8 FILLER_18_582 ();
 sg13g2_decap_8 FILLER_18_589 ();
 sg13g2_decap_8 FILLER_18_596 ();
 sg13g2_decap_8 FILLER_18_603 ();
 sg13g2_decap_8 FILLER_18_610 ();
 sg13g2_decap_8 FILLER_18_617 ();
 sg13g2_decap_8 FILLER_18_624 ();
 sg13g2_decap_8 FILLER_18_631 ();
 sg13g2_decap_8 FILLER_18_638 ();
 sg13g2_decap_8 FILLER_18_645 ();
 sg13g2_decap_8 FILLER_18_652 ();
 sg13g2_decap_8 FILLER_18_659 ();
 sg13g2_decap_8 FILLER_18_666 ();
 sg13g2_decap_8 FILLER_18_673 ();
 sg13g2_decap_8 FILLER_18_680 ();
 sg13g2_decap_8 FILLER_18_687 ();
 sg13g2_decap_8 FILLER_18_694 ();
 sg13g2_decap_8 FILLER_18_701 ();
 sg13g2_decap_8 FILLER_18_708 ();
 sg13g2_decap_8 FILLER_18_715 ();
 sg13g2_decap_8 FILLER_18_722 ();
 sg13g2_decap_8 FILLER_18_729 ();
 sg13g2_decap_8 FILLER_18_736 ();
 sg13g2_decap_8 FILLER_18_743 ();
 sg13g2_decap_8 FILLER_18_750 ();
 sg13g2_decap_8 FILLER_18_757 ();
 sg13g2_decap_8 FILLER_18_764 ();
 sg13g2_decap_8 FILLER_18_771 ();
 sg13g2_decap_8 FILLER_18_778 ();
 sg13g2_decap_8 FILLER_18_785 ();
 sg13g2_decap_8 FILLER_18_792 ();
 sg13g2_decap_8 FILLER_18_799 ();
 sg13g2_decap_8 FILLER_18_806 ();
 sg13g2_decap_8 FILLER_18_813 ();
 sg13g2_decap_8 FILLER_18_820 ();
 sg13g2_decap_8 FILLER_18_827 ();
 sg13g2_decap_8 FILLER_18_834 ();
 sg13g2_decap_8 FILLER_18_841 ();
 sg13g2_decap_8 FILLER_18_848 ();
 sg13g2_decap_8 FILLER_18_855 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_42 ();
 sg13g2_fill_1 FILLER_19_44 ();
 sg13g2_fill_2 FILLER_19_80 ();
 sg13g2_fill_1 FILLER_19_91 ();
 sg13g2_fill_2 FILLER_19_136 ();
 sg13g2_fill_1 FILLER_19_138 ();
 sg13g2_decap_4 FILLER_19_150 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_198 ();
 sg13g2_decap_4 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_213 ();
 sg13g2_decap_8 FILLER_19_219 ();
 sg13g2_decap_8 FILLER_19_226 ();
 sg13g2_decap_4 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_274 ();
 sg13g2_fill_1 FILLER_19_276 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_341 ();
 sg13g2_fill_1 FILLER_19_343 ();
 sg13g2_decap_4 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_379 ();
 sg13g2_decap_4 FILLER_19_393 ();
 sg13g2_fill_2 FILLER_19_400 ();
 sg13g2_fill_1 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_431 ();
 sg13g2_fill_1 FILLER_19_433 ();
 sg13g2_fill_2 FILLER_19_452 ();
 sg13g2_fill_2 FILLER_19_473 ();
 sg13g2_decap_4 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_fill_2 FILLER_20_68 ();
 sg13g2_fill_1 FILLER_20_70 ();
 sg13g2_fill_2 FILLER_20_83 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_fill_1 FILLER_20_326 ();
 sg13g2_fill_1 FILLER_20_332 ();
 sg13g2_fill_2 FILLER_20_372 ();
 sg13g2_fill_1 FILLER_20_374 ();
 sg13g2_decap_4 FILLER_20_383 ();
 sg13g2_fill_2 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_4 FILLER_20_427 ();
 sg13g2_decap_4 FILLER_20_436 ();
 sg13g2_fill_2 FILLER_20_440 ();
 sg13g2_fill_2 FILLER_20_455 ();
 sg13g2_fill_1 FILLER_20_461 ();
 sg13g2_decap_8 FILLER_20_480 ();
 sg13g2_decap_8 FILLER_20_496 ();
 sg13g2_decap_8 FILLER_20_503 ();
 sg13g2_decap_8 FILLER_20_510 ();
 sg13g2_decap_8 FILLER_20_517 ();
 sg13g2_decap_8 FILLER_20_524 ();
 sg13g2_decap_8 FILLER_20_531 ();
 sg13g2_decap_8 FILLER_20_538 ();
 sg13g2_decap_8 FILLER_20_545 ();
 sg13g2_decap_8 FILLER_20_552 ();
 sg13g2_decap_8 FILLER_20_559 ();
 sg13g2_decap_8 FILLER_20_566 ();
 sg13g2_decap_8 FILLER_20_573 ();
 sg13g2_decap_8 FILLER_20_580 ();
 sg13g2_decap_8 FILLER_20_587 ();
 sg13g2_decap_8 FILLER_20_594 ();
 sg13g2_decap_8 FILLER_20_601 ();
 sg13g2_decap_8 FILLER_20_608 ();
 sg13g2_decap_8 FILLER_20_615 ();
 sg13g2_decap_8 FILLER_20_622 ();
 sg13g2_decap_8 FILLER_20_629 ();
 sg13g2_decap_8 FILLER_20_636 ();
 sg13g2_decap_8 FILLER_20_643 ();
 sg13g2_decap_8 FILLER_20_650 ();
 sg13g2_decap_8 FILLER_20_657 ();
 sg13g2_decap_8 FILLER_20_664 ();
 sg13g2_decap_8 FILLER_20_671 ();
 sg13g2_decap_8 FILLER_20_678 ();
 sg13g2_decap_8 FILLER_20_685 ();
 sg13g2_decap_8 FILLER_20_692 ();
 sg13g2_decap_8 FILLER_20_699 ();
 sg13g2_decap_8 FILLER_20_706 ();
 sg13g2_decap_8 FILLER_20_713 ();
 sg13g2_decap_8 FILLER_20_720 ();
 sg13g2_decap_8 FILLER_20_727 ();
 sg13g2_decap_8 FILLER_20_734 ();
 sg13g2_decap_8 FILLER_20_741 ();
 sg13g2_decap_8 FILLER_20_748 ();
 sg13g2_decap_8 FILLER_20_755 ();
 sg13g2_decap_8 FILLER_20_762 ();
 sg13g2_decap_8 FILLER_20_769 ();
 sg13g2_decap_8 FILLER_20_776 ();
 sg13g2_decap_8 FILLER_20_783 ();
 sg13g2_decap_8 FILLER_20_790 ();
 sg13g2_decap_8 FILLER_20_797 ();
 sg13g2_decap_8 FILLER_20_804 ();
 sg13g2_decap_8 FILLER_20_811 ();
 sg13g2_decap_8 FILLER_20_818 ();
 sg13g2_decap_8 FILLER_20_825 ();
 sg13g2_decap_8 FILLER_20_832 ();
 sg13g2_decap_8 FILLER_20_839 ();
 sg13g2_decap_8 FILLER_20_846 ();
 sg13g2_decap_8 FILLER_20_853 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_decap_4 FILLER_21_127 ();
 sg13g2_fill_1 FILLER_21_131 ();
 sg13g2_fill_1 FILLER_21_147 ();
 sg13g2_fill_1 FILLER_21_160 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_fill_2 FILLER_21_194 ();
 sg13g2_fill_1 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_fill_2 FILLER_21_230 ();
 sg13g2_fill_2 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_297 ();
 sg13g2_fill_2 FILLER_21_313 ();
 sg13g2_fill_1 FILLER_21_315 ();
 sg13g2_fill_2 FILLER_21_335 ();
 sg13g2_fill_2 FILLER_21_347 ();
 sg13g2_fill_2 FILLER_21_353 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_fill_2 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_414 ();
 sg13g2_fill_1 FILLER_21_446 ();
 sg13g2_decap_8 FILLER_21_466 ();
 sg13g2_fill_2 FILLER_21_473 ();
 sg13g2_fill_1 FILLER_21_475 ();
 sg13g2_decap_8 FILLER_21_503 ();
 sg13g2_decap_8 FILLER_21_510 ();
 sg13g2_decap_8 FILLER_21_517 ();
 sg13g2_decap_8 FILLER_21_524 ();
 sg13g2_decap_8 FILLER_21_531 ();
 sg13g2_decap_8 FILLER_21_538 ();
 sg13g2_decap_8 FILLER_21_545 ();
 sg13g2_decap_8 FILLER_21_552 ();
 sg13g2_decap_8 FILLER_21_559 ();
 sg13g2_decap_8 FILLER_21_566 ();
 sg13g2_decap_8 FILLER_21_573 ();
 sg13g2_decap_8 FILLER_21_580 ();
 sg13g2_decap_8 FILLER_21_587 ();
 sg13g2_decap_8 FILLER_21_594 ();
 sg13g2_decap_8 FILLER_21_601 ();
 sg13g2_decap_8 FILLER_21_608 ();
 sg13g2_decap_8 FILLER_21_615 ();
 sg13g2_decap_8 FILLER_21_622 ();
 sg13g2_decap_8 FILLER_21_629 ();
 sg13g2_decap_8 FILLER_21_636 ();
 sg13g2_decap_8 FILLER_21_643 ();
 sg13g2_decap_8 FILLER_21_650 ();
 sg13g2_decap_8 FILLER_21_657 ();
 sg13g2_decap_8 FILLER_21_664 ();
 sg13g2_decap_8 FILLER_21_671 ();
 sg13g2_decap_8 FILLER_21_678 ();
 sg13g2_decap_8 FILLER_21_685 ();
 sg13g2_decap_8 FILLER_21_692 ();
 sg13g2_decap_8 FILLER_21_699 ();
 sg13g2_decap_8 FILLER_21_706 ();
 sg13g2_decap_8 FILLER_21_713 ();
 sg13g2_decap_8 FILLER_21_720 ();
 sg13g2_decap_8 FILLER_21_727 ();
 sg13g2_decap_8 FILLER_21_734 ();
 sg13g2_decap_8 FILLER_21_741 ();
 sg13g2_decap_8 FILLER_21_748 ();
 sg13g2_decap_8 FILLER_21_755 ();
 sg13g2_decap_8 FILLER_21_762 ();
 sg13g2_decap_8 FILLER_21_769 ();
 sg13g2_decap_8 FILLER_21_776 ();
 sg13g2_decap_8 FILLER_21_783 ();
 sg13g2_decap_8 FILLER_21_790 ();
 sg13g2_decap_8 FILLER_21_797 ();
 sg13g2_decap_8 FILLER_21_804 ();
 sg13g2_decap_8 FILLER_21_811 ();
 sg13g2_decap_8 FILLER_21_818 ();
 sg13g2_decap_8 FILLER_21_825 ();
 sg13g2_decap_8 FILLER_21_832 ();
 sg13g2_decap_8 FILLER_21_839 ();
 sg13g2_decap_8 FILLER_21_846 ();
 sg13g2_decap_8 FILLER_21_853 ();
 sg13g2_fill_2 FILLER_21_860 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_fill_2 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_36 ();
 sg13g2_fill_2 FILLER_22_46 ();
 sg13g2_fill_2 FILLER_22_74 ();
 sg13g2_fill_1 FILLER_22_76 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_fill_1 FILLER_22_111 ();
 sg13g2_fill_2 FILLER_22_125 ();
 sg13g2_decap_8 FILLER_22_131 ();
 sg13g2_fill_1 FILLER_22_138 ();
 sg13g2_fill_2 FILLER_22_160 ();
 sg13g2_fill_1 FILLER_22_162 ();
 sg13g2_fill_2 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_281 ();
 sg13g2_fill_2 FILLER_22_311 ();
 sg13g2_fill_2 FILLER_22_327 ();
 sg13g2_fill_1 FILLER_22_373 ();
 sg13g2_fill_2 FILLER_22_382 ();
 sg13g2_fill_2 FILLER_22_388 ();
 sg13g2_fill_2 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_fill_2 FILLER_22_424 ();
 sg13g2_fill_1 FILLER_22_426 ();
 sg13g2_fill_1 FILLER_22_448 ();
 sg13g2_decap_4 FILLER_22_458 ();
 sg13g2_fill_1 FILLER_22_462 ();
 sg13g2_fill_2 FILLER_22_471 ();
 sg13g2_fill_2 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_512 ();
 sg13g2_decap_8 FILLER_22_519 ();
 sg13g2_decap_8 FILLER_22_526 ();
 sg13g2_decap_8 FILLER_22_533 ();
 sg13g2_decap_8 FILLER_22_540 ();
 sg13g2_decap_8 FILLER_22_547 ();
 sg13g2_decap_8 FILLER_22_554 ();
 sg13g2_decap_8 FILLER_22_561 ();
 sg13g2_decap_8 FILLER_22_568 ();
 sg13g2_decap_8 FILLER_22_575 ();
 sg13g2_decap_8 FILLER_22_582 ();
 sg13g2_decap_8 FILLER_22_589 ();
 sg13g2_decap_8 FILLER_22_596 ();
 sg13g2_decap_8 FILLER_22_603 ();
 sg13g2_decap_8 FILLER_22_610 ();
 sg13g2_decap_8 FILLER_22_617 ();
 sg13g2_decap_8 FILLER_22_624 ();
 sg13g2_decap_8 FILLER_22_631 ();
 sg13g2_decap_8 FILLER_22_638 ();
 sg13g2_decap_8 FILLER_22_645 ();
 sg13g2_decap_8 FILLER_22_652 ();
 sg13g2_decap_8 FILLER_22_659 ();
 sg13g2_decap_8 FILLER_22_666 ();
 sg13g2_decap_8 FILLER_22_673 ();
 sg13g2_decap_8 FILLER_22_680 ();
 sg13g2_decap_8 FILLER_22_687 ();
 sg13g2_decap_8 FILLER_22_694 ();
 sg13g2_decap_8 FILLER_22_701 ();
 sg13g2_decap_8 FILLER_22_708 ();
 sg13g2_decap_8 FILLER_22_715 ();
 sg13g2_decap_8 FILLER_22_722 ();
 sg13g2_decap_8 FILLER_22_729 ();
 sg13g2_decap_8 FILLER_22_736 ();
 sg13g2_decap_8 FILLER_22_743 ();
 sg13g2_decap_8 FILLER_22_750 ();
 sg13g2_decap_8 FILLER_22_757 ();
 sg13g2_decap_8 FILLER_22_764 ();
 sg13g2_decap_8 FILLER_22_771 ();
 sg13g2_decap_8 FILLER_22_778 ();
 sg13g2_decap_8 FILLER_22_785 ();
 sg13g2_decap_8 FILLER_22_792 ();
 sg13g2_decap_8 FILLER_22_799 ();
 sg13g2_decap_8 FILLER_22_806 ();
 sg13g2_decap_8 FILLER_22_813 ();
 sg13g2_decap_8 FILLER_22_820 ();
 sg13g2_decap_8 FILLER_22_827 ();
 sg13g2_decap_8 FILLER_22_834 ();
 sg13g2_decap_8 FILLER_22_841 ();
 sg13g2_decap_8 FILLER_22_848 ();
 sg13g2_decap_8 FILLER_22_855 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_11 ();
 sg13g2_fill_2 FILLER_23_60 ();
 sg13g2_fill_1 FILLER_23_71 ();
 sg13g2_fill_2 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_195 ();
 sg13g2_decap_4 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_325 ();
 sg13g2_fill_2 FILLER_23_331 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_387 ();
 sg13g2_decap_4 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_416 ();
 sg13g2_fill_1 FILLER_23_423 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_fill_2 FILLER_23_452 ();
 sg13g2_decap_8 FILLER_23_472 ();
 sg13g2_decap_8 FILLER_23_479 ();
 sg13g2_decap_4 FILLER_23_486 ();
 sg13g2_decap_8 FILLER_23_509 ();
 sg13g2_decap_8 FILLER_23_516 ();
 sg13g2_decap_8 FILLER_23_523 ();
 sg13g2_decap_8 FILLER_23_530 ();
 sg13g2_decap_8 FILLER_23_537 ();
 sg13g2_decap_8 FILLER_23_544 ();
 sg13g2_decap_8 FILLER_23_551 ();
 sg13g2_decap_8 FILLER_23_558 ();
 sg13g2_decap_8 FILLER_23_565 ();
 sg13g2_decap_8 FILLER_23_572 ();
 sg13g2_decap_8 FILLER_23_579 ();
 sg13g2_decap_8 FILLER_23_586 ();
 sg13g2_decap_8 FILLER_23_593 ();
 sg13g2_decap_8 FILLER_23_600 ();
 sg13g2_decap_8 FILLER_23_607 ();
 sg13g2_decap_8 FILLER_23_614 ();
 sg13g2_decap_8 FILLER_23_621 ();
 sg13g2_decap_8 FILLER_23_628 ();
 sg13g2_decap_8 FILLER_23_635 ();
 sg13g2_decap_8 FILLER_23_642 ();
 sg13g2_decap_8 FILLER_23_649 ();
 sg13g2_decap_8 FILLER_23_656 ();
 sg13g2_decap_8 FILLER_23_663 ();
 sg13g2_decap_8 FILLER_23_670 ();
 sg13g2_decap_8 FILLER_23_677 ();
 sg13g2_decap_8 FILLER_23_684 ();
 sg13g2_decap_8 FILLER_23_691 ();
 sg13g2_decap_8 FILLER_23_698 ();
 sg13g2_decap_8 FILLER_23_705 ();
 sg13g2_decap_8 FILLER_23_712 ();
 sg13g2_decap_8 FILLER_23_719 ();
 sg13g2_decap_8 FILLER_23_726 ();
 sg13g2_decap_8 FILLER_23_733 ();
 sg13g2_decap_8 FILLER_23_740 ();
 sg13g2_decap_8 FILLER_23_747 ();
 sg13g2_decap_8 FILLER_23_754 ();
 sg13g2_decap_8 FILLER_23_761 ();
 sg13g2_decap_8 FILLER_23_768 ();
 sg13g2_decap_8 FILLER_23_775 ();
 sg13g2_decap_8 FILLER_23_782 ();
 sg13g2_decap_8 FILLER_23_789 ();
 sg13g2_decap_8 FILLER_23_796 ();
 sg13g2_decap_8 FILLER_23_803 ();
 sg13g2_decap_8 FILLER_23_810 ();
 sg13g2_decap_8 FILLER_23_817 ();
 sg13g2_decap_8 FILLER_23_824 ();
 sg13g2_decap_8 FILLER_23_831 ();
 sg13g2_decap_8 FILLER_23_838 ();
 sg13g2_decap_8 FILLER_23_845 ();
 sg13g2_decap_8 FILLER_23_852 ();
 sg13g2_fill_2 FILLER_23_859 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_55 ();
 sg13g2_decap_4 FILLER_24_95 ();
 sg13g2_fill_2 FILLER_24_107 ();
 sg13g2_fill_2 FILLER_24_149 ();
 sg13g2_fill_1 FILLER_24_151 ();
 sg13g2_fill_2 FILLER_24_179 ();
 sg13g2_fill_1 FILLER_24_233 ();
 sg13g2_fill_2 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_326 ();
 sg13g2_fill_2 FILLER_24_337 ();
 sg13g2_fill_1 FILLER_24_365 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_fill_1 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_411 ();
 sg13g2_decap_4 FILLER_24_418 ();
 sg13g2_fill_1 FILLER_24_422 ();
 sg13g2_decap_8 FILLER_24_439 ();
 sg13g2_decap_8 FILLER_24_446 ();
 sg13g2_decap_8 FILLER_24_453 ();
 sg13g2_decap_8 FILLER_24_516 ();
 sg13g2_decap_8 FILLER_24_523 ();
 sg13g2_decap_8 FILLER_24_530 ();
 sg13g2_decap_8 FILLER_24_537 ();
 sg13g2_decap_8 FILLER_24_544 ();
 sg13g2_decap_8 FILLER_24_551 ();
 sg13g2_decap_8 FILLER_24_558 ();
 sg13g2_decap_8 FILLER_24_565 ();
 sg13g2_decap_8 FILLER_24_572 ();
 sg13g2_decap_8 FILLER_24_579 ();
 sg13g2_decap_8 FILLER_24_586 ();
 sg13g2_decap_8 FILLER_24_593 ();
 sg13g2_decap_8 FILLER_24_600 ();
 sg13g2_decap_8 FILLER_24_607 ();
 sg13g2_decap_8 FILLER_24_614 ();
 sg13g2_decap_8 FILLER_24_621 ();
 sg13g2_decap_8 FILLER_24_628 ();
 sg13g2_decap_8 FILLER_24_635 ();
 sg13g2_decap_8 FILLER_24_642 ();
 sg13g2_decap_8 FILLER_24_649 ();
 sg13g2_decap_8 FILLER_24_656 ();
 sg13g2_decap_8 FILLER_24_663 ();
 sg13g2_decap_8 FILLER_24_670 ();
 sg13g2_decap_8 FILLER_24_677 ();
 sg13g2_decap_8 FILLER_24_684 ();
 sg13g2_decap_8 FILLER_24_691 ();
 sg13g2_decap_8 FILLER_24_698 ();
 sg13g2_decap_8 FILLER_24_705 ();
 sg13g2_decap_8 FILLER_24_712 ();
 sg13g2_decap_8 FILLER_24_719 ();
 sg13g2_decap_8 FILLER_24_726 ();
 sg13g2_decap_8 FILLER_24_733 ();
 sg13g2_decap_8 FILLER_24_740 ();
 sg13g2_decap_8 FILLER_24_747 ();
 sg13g2_decap_8 FILLER_24_754 ();
 sg13g2_decap_8 FILLER_24_761 ();
 sg13g2_decap_8 FILLER_24_768 ();
 sg13g2_decap_8 FILLER_24_775 ();
 sg13g2_decap_8 FILLER_24_782 ();
 sg13g2_decap_8 FILLER_24_789 ();
 sg13g2_decap_8 FILLER_24_796 ();
 sg13g2_decap_8 FILLER_24_803 ();
 sg13g2_decap_8 FILLER_24_810 ();
 sg13g2_decap_8 FILLER_24_817 ();
 sg13g2_decap_8 FILLER_24_824 ();
 sg13g2_decap_8 FILLER_24_831 ();
 sg13g2_decap_8 FILLER_24_838 ();
 sg13g2_decap_8 FILLER_24_845 ();
 sg13g2_decap_8 FILLER_24_852 ();
 sg13g2_fill_2 FILLER_24_859 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_30 ();
 sg13g2_decap_4 FILLER_25_71 ();
 sg13g2_fill_1 FILLER_25_75 ();
 sg13g2_decap_4 FILLER_25_84 ();
 sg13g2_fill_2 FILLER_25_88 ();
 sg13g2_fill_1 FILLER_25_116 ();
 sg13g2_fill_2 FILLER_25_140 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_fill_2 FILLER_25_149 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_fill_1 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_217 ();
 sg13g2_fill_2 FILLER_25_291 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_fill_1 FILLER_25_319 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_327 ();
 sg13g2_fill_1 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_fill_2 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_fill_2 FILLER_25_416 ();
 sg13g2_fill_1 FILLER_25_418 ();
 sg13g2_decap_8 FILLER_25_442 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_4 FILLER_25_476 ();
 sg13g2_fill_2 FILLER_25_492 ();
 sg13g2_fill_1 FILLER_25_494 ();
 sg13g2_decap_8 FILLER_25_505 ();
 sg13g2_decap_8 FILLER_25_512 ();
 sg13g2_decap_8 FILLER_25_519 ();
 sg13g2_decap_8 FILLER_25_526 ();
 sg13g2_decap_8 FILLER_25_533 ();
 sg13g2_decap_8 FILLER_25_540 ();
 sg13g2_decap_8 FILLER_25_547 ();
 sg13g2_decap_8 FILLER_25_554 ();
 sg13g2_decap_8 FILLER_25_561 ();
 sg13g2_decap_8 FILLER_25_568 ();
 sg13g2_decap_8 FILLER_25_575 ();
 sg13g2_decap_8 FILLER_25_582 ();
 sg13g2_decap_8 FILLER_25_589 ();
 sg13g2_decap_8 FILLER_25_596 ();
 sg13g2_decap_8 FILLER_25_603 ();
 sg13g2_decap_8 FILLER_25_610 ();
 sg13g2_decap_8 FILLER_25_617 ();
 sg13g2_decap_8 FILLER_25_624 ();
 sg13g2_decap_8 FILLER_25_631 ();
 sg13g2_decap_8 FILLER_25_638 ();
 sg13g2_decap_8 FILLER_25_645 ();
 sg13g2_decap_8 FILLER_25_652 ();
 sg13g2_decap_8 FILLER_25_659 ();
 sg13g2_decap_8 FILLER_25_666 ();
 sg13g2_decap_8 FILLER_25_673 ();
 sg13g2_decap_8 FILLER_25_680 ();
 sg13g2_decap_8 FILLER_25_687 ();
 sg13g2_decap_8 FILLER_25_694 ();
 sg13g2_decap_8 FILLER_25_701 ();
 sg13g2_decap_8 FILLER_25_708 ();
 sg13g2_decap_8 FILLER_25_715 ();
 sg13g2_decap_8 FILLER_25_722 ();
 sg13g2_decap_8 FILLER_25_729 ();
 sg13g2_decap_8 FILLER_25_736 ();
 sg13g2_decap_8 FILLER_25_743 ();
 sg13g2_decap_8 FILLER_25_750 ();
 sg13g2_decap_8 FILLER_25_757 ();
 sg13g2_decap_8 FILLER_25_764 ();
 sg13g2_decap_8 FILLER_25_771 ();
 sg13g2_decap_8 FILLER_25_778 ();
 sg13g2_decap_8 FILLER_25_785 ();
 sg13g2_decap_8 FILLER_25_792 ();
 sg13g2_decap_8 FILLER_25_799 ();
 sg13g2_decap_8 FILLER_25_806 ();
 sg13g2_decap_8 FILLER_25_813 ();
 sg13g2_decap_8 FILLER_25_820 ();
 sg13g2_decap_8 FILLER_25_827 ();
 sg13g2_decap_8 FILLER_25_834 ();
 sg13g2_decap_8 FILLER_25_841 ();
 sg13g2_decap_8 FILLER_25_848 ();
 sg13g2_decap_8 FILLER_25_855 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_fill_2 FILLER_26_37 ();
 sg13g2_fill_1 FILLER_26_39 ();
 sg13g2_fill_2 FILLER_26_53 ();
 sg13g2_fill_1 FILLER_26_55 ();
 sg13g2_fill_1 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_fill_1 FILLER_26_111 ();
 sg13g2_fill_1 FILLER_26_143 ();
 sg13g2_fill_2 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_225 ();
 sg13g2_fill_2 FILLER_26_381 ();
 sg13g2_fill_1 FILLER_26_383 ();
 sg13g2_decap_4 FILLER_26_392 ();
 sg13g2_fill_1 FILLER_26_396 ();
 sg13g2_fill_2 FILLER_26_402 ();
 sg13g2_fill_1 FILLER_26_404 ();
 sg13g2_decap_4 FILLER_26_409 ();
 sg13g2_decap_8 FILLER_26_421 ();
 sg13g2_fill_1 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_26_453 ();
 sg13g2_decap_4 FILLER_26_460 ();
 sg13g2_fill_2 FILLER_26_464 ();
 sg13g2_fill_2 FILLER_26_471 ();
 sg13g2_fill_1 FILLER_26_473 ();
 sg13g2_decap_4 FILLER_26_491 ();
 sg13g2_fill_1 FILLER_26_495 ();
 sg13g2_decap_8 FILLER_26_519 ();
 sg13g2_decap_8 FILLER_26_526 ();
 sg13g2_decap_8 FILLER_26_533 ();
 sg13g2_decap_8 FILLER_26_540 ();
 sg13g2_decap_8 FILLER_26_547 ();
 sg13g2_decap_8 FILLER_26_554 ();
 sg13g2_decap_8 FILLER_26_561 ();
 sg13g2_decap_8 FILLER_26_568 ();
 sg13g2_decap_8 FILLER_26_575 ();
 sg13g2_decap_8 FILLER_26_582 ();
 sg13g2_decap_8 FILLER_26_589 ();
 sg13g2_decap_8 FILLER_26_596 ();
 sg13g2_decap_8 FILLER_26_603 ();
 sg13g2_decap_8 FILLER_26_610 ();
 sg13g2_decap_8 FILLER_26_617 ();
 sg13g2_decap_8 FILLER_26_624 ();
 sg13g2_decap_8 FILLER_26_631 ();
 sg13g2_decap_8 FILLER_26_638 ();
 sg13g2_decap_8 FILLER_26_645 ();
 sg13g2_decap_8 FILLER_26_652 ();
 sg13g2_decap_8 FILLER_26_659 ();
 sg13g2_decap_8 FILLER_26_666 ();
 sg13g2_decap_8 FILLER_26_673 ();
 sg13g2_decap_8 FILLER_26_680 ();
 sg13g2_decap_8 FILLER_26_687 ();
 sg13g2_decap_8 FILLER_26_694 ();
 sg13g2_decap_8 FILLER_26_701 ();
 sg13g2_decap_8 FILLER_26_708 ();
 sg13g2_decap_8 FILLER_26_715 ();
 sg13g2_decap_8 FILLER_26_722 ();
 sg13g2_decap_8 FILLER_26_729 ();
 sg13g2_decap_8 FILLER_26_736 ();
 sg13g2_decap_8 FILLER_26_743 ();
 sg13g2_decap_8 FILLER_26_750 ();
 sg13g2_decap_8 FILLER_26_757 ();
 sg13g2_decap_8 FILLER_26_764 ();
 sg13g2_decap_8 FILLER_26_771 ();
 sg13g2_decap_8 FILLER_26_778 ();
 sg13g2_decap_8 FILLER_26_785 ();
 sg13g2_decap_8 FILLER_26_792 ();
 sg13g2_decap_8 FILLER_26_799 ();
 sg13g2_decap_8 FILLER_26_806 ();
 sg13g2_decap_8 FILLER_26_813 ();
 sg13g2_decap_8 FILLER_26_820 ();
 sg13g2_decap_8 FILLER_26_827 ();
 sg13g2_decap_8 FILLER_26_834 ();
 sg13g2_decap_8 FILLER_26_841 ();
 sg13g2_decap_8 FILLER_26_848 ();
 sg13g2_decap_8 FILLER_26_855 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_2 FILLER_27_29 ();
 sg13g2_fill_1 FILLER_27_31 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_decap_4 FILLER_27_68 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_121 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_fill_2 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_fill_2 FILLER_27_218 ();
 sg13g2_fill_1 FILLER_27_220 ();
 sg13g2_fill_2 FILLER_27_229 ();
 sg13g2_fill_1 FILLER_27_231 ();
 sg13g2_fill_2 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_304 ();
 sg13g2_decap_4 FILLER_27_366 ();
 sg13g2_fill_2 FILLER_27_370 ();
 sg13g2_fill_1 FILLER_27_376 ();
 sg13g2_fill_1 FILLER_27_396 ();
 sg13g2_decap_8 FILLER_27_418 ();
 sg13g2_decap_8 FILLER_27_425 ();
 sg13g2_fill_1 FILLER_27_432 ();
 sg13g2_fill_2 FILLER_27_441 ();
 sg13g2_fill_2 FILLER_27_448 ();
 sg13g2_fill_1 FILLER_27_450 ();
 sg13g2_decap_4 FILLER_27_461 ();
 sg13g2_fill_1 FILLER_27_465 ();
 sg13g2_fill_2 FILLER_27_474 ();
 sg13g2_fill_2 FILLER_27_492 ();
 sg13g2_fill_1 FILLER_27_494 ();
 sg13g2_fill_2 FILLER_27_502 ();
 sg13g2_fill_1 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_522 ();
 sg13g2_decap_8 FILLER_27_529 ();
 sg13g2_decap_8 FILLER_27_536 ();
 sg13g2_decap_8 FILLER_27_543 ();
 sg13g2_decap_8 FILLER_27_550 ();
 sg13g2_decap_8 FILLER_27_557 ();
 sg13g2_decap_8 FILLER_27_564 ();
 sg13g2_decap_8 FILLER_27_571 ();
 sg13g2_decap_8 FILLER_27_578 ();
 sg13g2_decap_8 FILLER_27_585 ();
 sg13g2_decap_8 FILLER_27_592 ();
 sg13g2_decap_8 FILLER_27_599 ();
 sg13g2_decap_8 FILLER_27_606 ();
 sg13g2_decap_8 FILLER_27_613 ();
 sg13g2_decap_8 FILLER_27_620 ();
 sg13g2_decap_8 FILLER_27_627 ();
 sg13g2_decap_8 FILLER_27_634 ();
 sg13g2_decap_8 FILLER_27_641 ();
 sg13g2_decap_8 FILLER_27_648 ();
 sg13g2_decap_8 FILLER_27_655 ();
 sg13g2_decap_8 FILLER_27_662 ();
 sg13g2_decap_8 FILLER_27_669 ();
 sg13g2_decap_8 FILLER_27_676 ();
 sg13g2_decap_8 FILLER_27_683 ();
 sg13g2_decap_8 FILLER_27_690 ();
 sg13g2_decap_8 FILLER_27_697 ();
 sg13g2_decap_8 FILLER_27_704 ();
 sg13g2_decap_8 FILLER_27_711 ();
 sg13g2_decap_8 FILLER_27_718 ();
 sg13g2_decap_8 FILLER_27_725 ();
 sg13g2_decap_8 FILLER_27_732 ();
 sg13g2_decap_8 FILLER_27_739 ();
 sg13g2_decap_8 FILLER_27_746 ();
 sg13g2_decap_8 FILLER_27_753 ();
 sg13g2_decap_8 FILLER_27_760 ();
 sg13g2_decap_8 FILLER_27_767 ();
 sg13g2_decap_8 FILLER_27_774 ();
 sg13g2_decap_8 FILLER_27_781 ();
 sg13g2_decap_8 FILLER_27_788 ();
 sg13g2_decap_8 FILLER_27_795 ();
 sg13g2_decap_8 FILLER_27_802 ();
 sg13g2_decap_8 FILLER_27_809 ();
 sg13g2_decap_8 FILLER_27_816 ();
 sg13g2_decap_8 FILLER_27_823 ();
 sg13g2_decap_8 FILLER_27_830 ();
 sg13g2_decap_8 FILLER_27_837 ();
 sg13g2_decap_8 FILLER_27_844 ();
 sg13g2_decap_8 FILLER_27_851 ();
 sg13g2_decap_4 FILLER_27_858 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_64 ();
 sg13g2_fill_1 FILLER_28_82 ();
 sg13g2_fill_1 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_164 ();
 sg13g2_fill_1 FILLER_28_170 ();
 sg13g2_decap_8 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_183 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_decap_4 FILLER_28_190 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_296 ();
 sg13g2_fill_2 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_fill_2 FILLER_28_382 ();
 sg13g2_fill_1 FILLER_28_402 ();
 sg13g2_decap_4 FILLER_28_411 ();
 sg13g2_fill_2 FILLER_28_415 ();
 sg13g2_decap_4 FILLER_28_438 ();
 sg13g2_fill_1 FILLER_28_442 ();
 sg13g2_fill_2 FILLER_28_491 ();
 sg13g2_fill_2 FILLER_28_497 ();
 sg13g2_fill_1 FILLER_28_499 ();
 sg13g2_decap_8 FILLER_28_518 ();
 sg13g2_decap_8 FILLER_28_525 ();
 sg13g2_decap_8 FILLER_28_532 ();
 sg13g2_decap_8 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_546 ();
 sg13g2_decap_8 FILLER_28_553 ();
 sg13g2_decap_8 FILLER_28_560 ();
 sg13g2_decap_8 FILLER_28_567 ();
 sg13g2_decap_8 FILLER_28_574 ();
 sg13g2_decap_8 FILLER_28_581 ();
 sg13g2_decap_8 FILLER_28_588 ();
 sg13g2_decap_8 FILLER_28_595 ();
 sg13g2_decap_8 FILLER_28_602 ();
 sg13g2_decap_8 FILLER_28_609 ();
 sg13g2_decap_8 FILLER_28_616 ();
 sg13g2_decap_8 FILLER_28_623 ();
 sg13g2_decap_8 FILLER_28_630 ();
 sg13g2_decap_8 FILLER_28_637 ();
 sg13g2_decap_8 FILLER_28_644 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_decap_8 FILLER_28_665 ();
 sg13g2_decap_8 FILLER_28_672 ();
 sg13g2_decap_8 FILLER_28_679 ();
 sg13g2_decap_8 FILLER_28_686 ();
 sg13g2_decap_8 FILLER_28_693 ();
 sg13g2_decap_8 FILLER_28_700 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_11 ();
 sg13g2_fill_2 FILLER_29_26 ();
 sg13g2_fill_1 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_47 ();
 sg13g2_fill_2 FILLER_29_51 ();
 sg13g2_fill_2 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_fill_1 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_333 ();
 sg13g2_fill_2 FILLER_29_339 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_fill_2 FILLER_29_377 ();
 sg13g2_fill_1 FILLER_29_379 ();
 sg13g2_fill_1 FILLER_29_400 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_fill_2 FILLER_29_441 ();
 sg13g2_fill_1 FILLER_29_466 ();
 sg13g2_decap_4 FILLER_29_479 ();
 sg13g2_fill_1 FILLER_29_483 ();
 sg13g2_fill_2 FILLER_29_501 ();
 sg13g2_decap_8 FILLER_29_520 ();
 sg13g2_decap_8 FILLER_29_527 ();
 sg13g2_decap_8 FILLER_29_534 ();
 sg13g2_decap_8 FILLER_29_541 ();
 sg13g2_decap_8 FILLER_29_548 ();
 sg13g2_decap_8 FILLER_29_555 ();
 sg13g2_decap_8 FILLER_29_562 ();
 sg13g2_decap_8 FILLER_29_569 ();
 sg13g2_decap_8 FILLER_29_576 ();
 sg13g2_decap_8 FILLER_29_583 ();
 sg13g2_decap_8 FILLER_29_590 ();
 sg13g2_decap_8 FILLER_29_597 ();
 sg13g2_decap_8 FILLER_29_604 ();
 sg13g2_decap_8 FILLER_29_611 ();
 sg13g2_decap_8 FILLER_29_618 ();
 sg13g2_decap_8 FILLER_29_625 ();
 sg13g2_decap_8 FILLER_29_632 ();
 sg13g2_decap_8 FILLER_29_639 ();
 sg13g2_decap_8 FILLER_29_646 ();
 sg13g2_decap_8 FILLER_29_653 ();
 sg13g2_decap_8 FILLER_29_660 ();
 sg13g2_decap_8 FILLER_29_667 ();
 sg13g2_decap_8 FILLER_29_674 ();
 sg13g2_decap_8 FILLER_29_681 ();
 sg13g2_decap_8 FILLER_29_688 ();
 sg13g2_decap_8 FILLER_29_695 ();
 sg13g2_decap_8 FILLER_29_702 ();
 sg13g2_decap_8 FILLER_29_709 ();
 sg13g2_decap_8 FILLER_29_716 ();
 sg13g2_decap_8 FILLER_29_723 ();
 sg13g2_decap_8 FILLER_29_730 ();
 sg13g2_decap_8 FILLER_29_737 ();
 sg13g2_decap_8 FILLER_29_744 ();
 sg13g2_decap_8 FILLER_29_751 ();
 sg13g2_decap_8 FILLER_29_758 ();
 sg13g2_decap_8 FILLER_29_765 ();
 sg13g2_decap_8 FILLER_29_772 ();
 sg13g2_decap_8 FILLER_29_779 ();
 sg13g2_decap_8 FILLER_29_786 ();
 sg13g2_decap_8 FILLER_29_793 ();
 sg13g2_decap_8 FILLER_29_800 ();
 sg13g2_decap_8 FILLER_29_807 ();
 sg13g2_decap_8 FILLER_29_814 ();
 sg13g2_decap_8 FILLER_29_821 ();
 sg13g2_decap_8 FILLER_29_828 ();
 sg13g2_decap_8 FILLER_29_835 ();
 sg13g2_decap_8 FILLER_29_842 ();
 sg13g2_decap_8 FILLER_29_849 ();
 sg13g2_decap_4 FILLER_29_856 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_2 FILLER_30_29 ();
 sg13g2_fill_1 FILLER_30_31 ();
 sg13g2_fill_1 FILLER_30_47 ();
 sg13g2_fill_1 FILLER_30_52 ();
 sg13g2_fill_1 FILLER_30_70 ();
 sg13g2_decap_4 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_fill_2 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_311 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_decap_4 FILLER_30_346 ();
 sg13g2_fill_2 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_356 ();
 sg13g2_decap_4 FILLER_30_363 ();
 sg13g2_fill_1 FILLER_30_367 ();
 sg13g2_fill_2 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_435 ();
 sg13g2_fill_2 FILLER_30_451 ();
 sg13g2_fill_1 FILLER_30_453 ();
 sg13g2_fill_1 FILLER_30_459 ();
 sg13g2_decap_8 FILLER_30_473 ();
 sg13g2_decap_8 FILLER_30_480 ();
 sg13g2_fill_2 FILLER_30_487 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_decap_4 FILLER_30_504 ();
 sg13g2_fill_1 FILLER_30_508 ();
 sg13g2_decap_8 FILLER_30_517 ();
 sg13g2_decap_8 FILLER_30_524 ();
 sg13g2_decap_8 FILLER_30_531 ();
 sg13g2_decap_8 FILLER_30_538 ();
 sg13g2_decap_8 FILLER_30_545 ();
 sg13g2_decap_8 FILLER_30_552 ();
 sg13g2_decap_8 FILLER_30_559 ();
 sg13g2_decap_8 FILLER_30_566 ();
 sg13g2_decap_8 FILLER_30_573 ();
 sg13g2_decap_8 FILLER_30_580 ();
 sg13g2_decap_8 FILLER_30_587 ();
 sg13g2_decap_8 FILLER_30_594 ();
 sg13g2_decap_8 FILLER_30_601 ();
 sg13g2_decap_8 FILLER_30_608 ();
 sg13g2_decap_8 FILLER_30_615 ();
 sg13g2_decap_8 FILLER_30_622 ();
 sg13g2_decap_8 FILLER_30_629 ();
 sg13g2_decap_8 FILLER_30_636 ();
 sg13g2_decap_8 FILLER_30_643 ();
 sg13g2_decap_8 FILLER_30_650 ();
 sg13g2_decap_8 FILLER_30_657 ();
 sg13g2_decap_8 FILLER_30_664 ();
 sg13g2_decap_8 FILLER_30_671 ();
 sg13g2_decap_8 FILLER_30_678 ();
 sg13g2_decap_8 FILLER_30_685 ();
 sg13g2_decap_8 FILLER_30_692 ();
 sg13g2_decap_8 FILLER_30_699 ();
 sg13g2_decap_8 FILLER_30_706 ();
 sg13g2_decap_8 FILLER_30_713 ();
 sg13g2_decap_8 FILLER_30_720 ();
 sg13g2_decap_8 FILLER_30_727 ();
 sg13g2_decap_8 FILLER_30_734 ();
 sg13g2_decap_8 FILLER_30_741 ();
 sg13g2_decap_8 FILLER_30_748 ();
 sg13g2_decap_8 FILLER_30_755 ();
 sg13g2_decap_8 FILLER_30_762 ();
 sg13g2_decap_8 FILLER_30_769 ();
 sg13g2_decap_8 FILLER_30_776 ();
 sg13g2_decap_8 FILLER_30_783 ();
 sg13g2_decap_8 FILLER_30_790 ();
 sg13g2_decap_8 FILLER_30_797 ();
 sg13g2_decap_8 FILLER_30_804 ();
 sg13g2_decap_8 FILLER_30_811 ();
 sg13g2_decap_8 FILLER_30_818 ();
 sg13g2_decap_8 FILLER_30_825 ();
 sg13g2_decap_8 FILLER_30_832 ();
 sg13g2_decap_8 FILLER_30_839 ();
 sg13g2_decap_8 FILLER_30_846 ();
 sg13g2_decap_8 FILLER_30_853 ();
 sg13g2_fill_2 FILLER_30_860 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_9 ();
 sg13g2_decap_4 FILLER_31_27 ();
 sg13g2_fill_1 FILLER_31_31 ();
 sg13g2_decap_4 FILLER_31_62 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_163 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_180 ();
 sg13g2_fill_2 FILLER_31_197 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_fill_1 FILLER_31_215 ();
 sg13g2_fill_1 FILLER_31_242 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_decap_4 FILLER_31_326 ();
 sg13g2_fill_1 FILLER_31_330 ();
 sg13g2_fill_2 FILLER_31_382 ();
 sg13g2_fill_1 FILLER_31_402 ();
 sg13g2_fill_1 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_4 FILLER_31_427 ();
 sg13g2_fill_1 FILLER_31_431 ();
 sg13g2_decap_4 FILLER_31_457 ();
 sg13g2_fill_2 FILLER_31_461 ();
 sg13g2_decap_4 FILLER_31_468 ();
 sg13g2_decap_4 FILLER_31_480 ();
 sg13g2_fill_2 FILLER_31_484 ();
 sg13g2_decap_8 FILLER_31_503 ();
 sg13g2_decap_8 FILLER_31_510 ();
 sg13g2_decap_8 FILLER_31_517 ();
 sg13g2_decap_8 FILLER_31_524 ();
 sg13g2_decap_8 FILLER_31_531 ();
 sg13g2_decap_8 FILLER_31_538 ();
 sg13g2_decap_8 FILLER_31_545 ();
 sg13g2_decap_8 FILLER_31_552 ();
 sg13g2_decap_8 FILLER_31_559 ();
 sg13g2_decap_8 FILLER_31_566 ();
 sg13g2_decap_8 FILLER_31_573 ();
 sg13g2_decap_8 FILLER_31_580 ();
 sg13g2_decap_8 FILLER_31_587 ();
 sg13g2_decap_8 FILLER_31_594 ();
 sg13g2_decap_8 FILLER_31_601 ();
 sg13g2_decap_8 FILLER_31_608 ();
 sg13g2_decap_8 FILLER_31_615 ();
 sg13g2_decap_8 FILLER_31_622 ();
 sg13g2_decap_8 FILLER_31_629 ();
 sg13g2_decap_8 FILLER_31_636 ();
 sg13g2_decap_8 FILLER_31_643 ();
 sg13g2_decap_8 FILLER_31_650 ();
 sg13g2_decap_8 FILLER_31_657 ();
 sg13g2_decap_8 FILLER_31_664 ();
 sg13g2_decap_8 FILLER_31_671 ();
 sg13g2_decap_8 FILLER_31_678 ();
 sg13g2_decap_8 FILLER_31_685 ();
 sg13g2_decap_8 FILLER_31_692 ();
 sg13g2_decap_8 FILLER_31_699 ();
 sg13g2_decap_8 FILLER_31_706 ();
 sg13g2_decap_8 FILLER_31_713 ();
 sg13g2_decap_8 FILLER_31_720 ();
 sg13g2_decap_8 FILLER_31_727 ();
 sg13g2_decap_8 FILLER_31_734 ();
 sg13g2_decap_8 FILLER_31_741 ();
 sg13g2_decap_8 FILLER_31_748 ();
 sg13g2_decap_8 FILLER_31_755 ();
 sg13g2_decap_8 FILLER_31_762 ();
 sg13g2_decap_8 FILLER_31_769 ();
 sg13g2_decap_8 FILLER_31_776 ();
 sg13g2_decap_8 FILLER_31_783 ();
 sg13g2_decap_8 FILLER_31_790 ();
 sg13g2_decap_8 FILLER_31_797 ();
 sg13g2_decap_8 FILLER_31_804 ();
 sg13g2_decap_8 FILLER_31_811 ();
 sg13g2_decap_8 FILLER_31_818 ();
 sg13g2_decap_8 FILLER_31_825 ();
 sg13g2_decap_8 FILLER_31_832 ();
 sg13g2_decap_8 FILLER_31_839 ();
 sg13g2_decap_8 FILLER_31_846 ();
 sg13g2_decap_8 FILLER_31_853 ();
 sg13g2_fill_2 FILLER_31_860 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_59 ();
 sg13g2_decap_8 FILLER_32_66 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_fill_2 FILLER_32_136 ();
 sg13g2_decap_8 FILLER_32_162 ();
 sg13g2_fill_2 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_fill_1 FILLER_32_225 ();
 sg13g2_fill_2 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_fill_2 FILLER_32_326 ();
 sg13g2_fill_1 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_360 ();
 sg13g2_decap_4 FILLER_32_378 ();
 sg13g2_fill_2 FILLER_32_390 ();
 sg13g2_fill_1 FILLER_32_392 ();
 sg13g2_fill_2 FILLER_32_411 ();
 sg13g2_decap_4 FILLER_32_429 ();
 sg13g2_fill_2 FILLER_32_433 ();
 sg13g2_fill_2 FILLER_32_449 ();
 sg13g2_fill_1 FILLER_32_451 ();
 sg13g2_fill_1 FILLER_32_462 ();
 sg13g2_decap_4 FILLER_32_479 ();
 sg13g2_fill_1 FILLER_32_483 ();
 sg13g2_decap_8 FILLER_32_505 ();
 sg13g2_decap_8 FILLER_32_512 ();
 sg13g2_decap_8 FILLER_32_519 ();
 sg13g2_decap_8 FILLER_32_526 ();
 sg13g2_decap_8 FILLER_32_533 ();
 sg13g2_decap_8 FILLER_32_540 ();
 sg13g2_decap_8 FILLER_32_547 ();
 sg13g2_decap_8 FILLER_32_554 ();
 sg13g2_decap_8 FILLER_32_561 ();
 sg13g2_decap_4 FILLER_32_568 ();
 sg13g2_decap_8 FILLER_32_577 ();
 sg13g2_decap_8 FILLER_32_584 ();
 sg13g2_decap_8 FILLER_32_591 ();
 sg13g2_decap_8 FILLER_32_598 ();
 sg13g2_decap_8 FILLER_32_605 ();
 sg13g2_decap_8 FILLER_32_612 ();
 sg13g2_decap_8 FILLER_32_619 ();
 sg13g2_decap_8 FILLER_32_626 ();
 sg13g2_decap_8 FILLER_32_633 ();
 sg13g2_decap_8 FILLER_32_640 ();
 sg13g2_decap_8 FILLER_32_647 ();
 sg13g2_decap_8 FILLER_32_654 ();
 sg13g2_decap_8 FILLER_32_661 ();
 sg13g2_decap_8 FILLER_32_668 ();
 sg13g2_decap_8 FILLER_32_675 ();
 sg13g2_decap_8 FILLER_32_682 ();
 sg13g2_decap_8 FILLER_32_689 ();
 sg13g2_decap_8 FILLER_32_696 ();
 sg13g2_decap_8 FILLER_32_703 ();
 sg13g2_decap_8 FILLER_32_710 ();
 sg13g2_decap_8 FILLER_32_717 ();
 sg13g2_decap_8 FILLER_32_724 ();
 sg13g2_decap_8 FILLER_32_731 ();
 sg13g2_decap_8 FILLER_32_738 ();
 sg13g2_decap_8 FILLER_32_745 ();
 sg13g2_decap_8 FILLER_32_752 ();
 sg13g2_decap_8 FILLER_32_759 ();
 sg13g2_decap_8 FILLER_32_766 ();
 sg13g2_decap_8 FILLER_32_773 ();
 sg13g2_decap_8 FILLER_32_780 ();
 sg13g2_decap_8 FILLER_32_787 ();
 sg13g2_decap_8 FILLER_32_794 ();
 sg13g2_decap_8 FILLER_32_801 ();
 sg13g2_decap_8 FILLER_32_808 ();
 sg13g2_decap_8 FILLER_32_815 ();
 sg13g2_decap_8 FILLER_32_822 ();
 sg13g2_decap_8 FILLER_32_829 ();
 sg13g2_decap_8 FILLER_32_836 ();
 sg13g2_decap_8 FILLER_32_843 ();
 sg13g2_decap_8 FILLER_32_850 ();
 sg13g2_decap_4 FILLER_32_857 ();
 sg13g2_fill_1 FILLER_32_861 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_20 ();
 sg13g2_fill_1 FILLER_33_27 ();
 sg13g2_fill_1 FILLER_33_51 ();
 sg13g2_fill_2 FILLER_33_57 ();
 sg13g2_fill_2 FILLER_33_82 ();
 sg13g2_fill_1 FILLER_33_102 ();
 sg13g2_fill_2 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_224 ();
 sg13g2_fill_2 FILLER_33_260 ();
 sg13g2_fill_1 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_277 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_decap_8 FILLER_33_334 ();
 sg13g2_decap_4 FILLER_33_341 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_356 ();
 sg13g2_decap_4 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_367 ();
 sg13g2_fill_2 FILLER_33_394 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_4 FILLER_33_414 ();
 sg13g2_fill_2 FILLER_33_418 ();
 sg13g2_fill_2 FILLER_33_425 ();
 sg13g2_decap_8 FILLER_33_436 ();
 sg13g2_fill_2 FILLER_33_443 ();
 sg13g2_decap_4 FILLER_33_450 ();
 sg13g2_fill_2 FILLER_33_462 ();
 sg13g2_fill_1 FILLER_33_464 ();
 sg13g2_fill_2 FILLER_33_477 ();
 sg13g2_fill_1 FILLER_33_479 ();
 sg13g2_decap_8 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_fill_2 FILLER_33_536 ();
 sg13g2_fill_1 FILLER_33_538 ();
 sg13g2_fill_1 FILLER_33_591 ();
 sg13g2_decap_8 FILLER_33_606 ();
 sg13g2_decap_8 FILLER_33_613 ();
 sg13g2_decap_8 FILLER_33_620 ();
 sg13g2_decap_8 FILLER_33_627 ();
 sg13g2_decap_8 FILLER_33_634 ();
 sg13g2_decap_8 FILLER_33_641 ();
 sg13g2_decap_8 FILLER_33_648 ();
 sg13g2_decap_8 FILLER_33_655 ();
 sg13g2_decap_8 FILLER_33_662 ();
 sg13g2_decap_8 FILLER_33_669 ();
 sg13g2_decap_8 FILLER_33_676 ();
 sg13g2_decap_8 FILLER_33_683 ();
 sg13g2_decap_8 FILLER_33_690 ();
 sg13g2_decap_8 FILLER_33_697 ();
 sg13g2_decap_8 FILLER_33_704 ();
 sg13g2_decap_8 FILLER_33_711 ();
 sg13g2_decap_8 FILLER_33_718 ();
 sg13g2_decap_8 FILLER_33_725 ();
 sg13g2_decap_8 FILLER_33_732 ();
 sg13g2_decap_8 FILLER_33_739 ();
 sg13g2_decap_8 FILLER_33_746 ();
 sg13g2_decap_8 FILLER_33_753 ();
 sg13g2_decap_8 FILLER_33_760 ();
 sg13g2_decap_8 FILLER_33_767 ();
 sg13g2_decap_8 FILLER_33_774 ();
 sg13g2_decap_8 FILLER_33_781 ();
 sg13g2_decap_8 FILLER_33_788 ();
 sg13g2_decap_8 FILLER_33_795 ();
 sg13g2_decap_8 FILLER_33_802 ();
 sg13g2_decap_8 FILLER_33_809 ();
 sg13g2_decap_8 FILLER_33_816 ();
 sg13g2_decap_8 FILLER_33_823 ();
 sg13g2_decap_8 FILLER_33_830 ();
 sg13g2_decap_8 FILLER_33_837 ();
 sg13g2_decap_8 FILLER_33_844 ();
 sg13g2_decap_8 FILLER_33_851 ();
 sg13g2_decap_4 FILLER_33_858 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_4 ();
 sg13g2_fill_2 FILLER_34_62 ();
 sg13g2_fill_1 FILLER_34_64 ();
 sg13g2_fill_2 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_fill_2 FILLER_34_134 ();
 sg13g2_fill_2 FILLER_34_152 ();
 sg13g2_fill_1 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_285 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_357 ();
 sg13g2_fill_2 FILLER_34_371 ();
 sg13g2_decap_4 FILLER_34_390 ();
 sg13g2_decap_4 FILLER_34_412 ();
 sg13g2_fill_2 FILLER_34_416 ();
 sg13g2_decap_4 FILLER_34_443 ();
 sg13g2_fill_2 FILLER_34_460 ();
 sg13g2_decap_8 FILLER_34_470 ();
 sg13g2_fill_2 FILLER_34_484 ();
 sg13g2_decap_4 FILLER_34_516 ();
 sg13g2_fill_1 FILLER_34_520 ();
 sg13g2_fill_2 FILLER_34_565 ();
 sg13g2_fill_2 FILLER_34_594 ();
 sg13g2_fill_1 FILLER_34_596 ();
 sg13g2_decap_8 FILLER_34_623 ();
 sg13g2_decap_8 FILLER_34_630 ();
 sg13g2_decap_8 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_644 ();
 sg13g2_decap_8 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_662 ();
 sg13g2_decap_8 FILLER_34_669 ();
 sg13g2_decap_8 FILLER_34_676 ();
 sg13g2_decap_8 FILLER_34_683 ();
 sg13g2_decap_8 FILLER_34_690 ();
 sg13g2_decap_8 FILLER_34_697 ();
 sg13g2_decap_8 FILLER_34_708 ();
 sg13g2_decap_8 FILLER_34_715 ();
 sg13g2_decap_8 FILLER_34_722 ();
 sg13g2_decap_8 FILLER_34_729 ();
 sg13g2_decap_8 FILLER_34_736 ();
 sg13g2_decap_8 FILLER_34_743 ();
 sg13g2_decap_8 FILLER_34_750 ();
 sg13g2_decap_8 FILLER_34_757 ();
 sg13g2_decap_8 FILLER_34_764 ();
 sg13g2_decap_8 FILLER_34_771 ();
 sg13g2_decap_8 FILLER_34_778 ();
 sg13g2_decap_8 FILLER_34_785 ();
 sg13g2_decap_8 FILLER_34_792 ();
 sg13g2_decap_8 FILLER_34_799 ();
 sg13g2_decap_8 FILLER_34_806 ();
 sg13g2_decap_8 FILLER_34_813 ();
 sg13g2_decap_8 FILLER_34_820 ();
 sg13g2_decap_8 FILLER_34_827 ();
 sg13g2_decap_8 FILLER_34_834 ();
 sg13g2_decap_8 FILLER_34_841 ();
 sg13g2_decap_8 FILLER_34_848 ();
 sg13g2_decap_8 FILLER_34_855 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_11 ();
 sg13g2_fill_2 FILLER_35_26 ();
 sg13g2_fill_1 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_57 ();
 sg13g2_fill_2 FILLER_35_74 ();
 sg13g2_fill_1 FILLER_35_76 ();
 sg13g2_fill_2 FILLER_35_86 ();
 sg13g2_fill_1 FILLER_35_88 ();
 sg13g2_fill_1 FILLER_35_124 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_fill_1 FILLER_35_153 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_221 ();
 sg13g2_fill_1 FILLER_35_231 ();
 sg13g2_fill_2 FILLER_35_242 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_2 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_332 ();
 sg13g2_fill_2 FILLER_35_339 ();
 sg13g2_fill_1 FILLER_35_341 ();
 sg13g2_fill_2 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_360 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_decap_4 FILLER_35_397 ();
 sg13g2_fill_2 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_414 ();
 sg13g2_decap_8 FILLER_35_421 ();
 sg13g2_fill_1 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_35_447 ();
 sg13g2_fill_2 FILLER_35_454 ();
 sg13g2_decap_8 FILLER_35_472 ();
 sg13g2_fill_2 FILLER_35_479 ();
 sg13g2_fill_1 FILLER_35_481 ();
 sg13g2_decap_4 FILLER_35_492 ();
 sg13g2_fill_2 FILLER_35_496 ();
 sg13g2_fill_2 FILLER_35_501 ();
 sg13g2_fill_1 FILLER_35_503 ();
 sg13g2_decap_4 FILLER_35_529 ();
 sg13g2_decap_4 FILLER_35_537 ();
 sg13g2_decap_4 FILLER_35_560 ();
 sg13g2_fill_2 FILLER_35_616 ();
 sg13g2_fill_1 FILLER_35_618 ();
 sg13g2_fill_1 FILLER_35_645 ();
 sg13g2_fill_2 FILLER_35_651 ();
 sg13g2_decap_4 FILLER_35_684 ();
 sg13g2_decap_8 FILLER_35_718 ();
 sg13g2_decap_8 FILLER_35_725 ();
 sg13g2_decap_8 FILLER_35_732 ();
 sg13g2_decap_8 FILLER_35_739 ();
 sg13g2_decap_8 FILLER_35_746 ();
 sg13g2_decap_8 FILLER_35_753 ();
 sg13g2_decap_8 FILLER_35_760 ();
 sg13g2_decap_8 FILLER_35_767 ();
 sg13g2_decap_8 FILLER_35_774 ();
 sg13g2_decap_8 FILLER_35_781 ();
 sg13g2_decap_8 FILLER_35_788 ();
 sg13g2_decap_8 FILLER_35_795 ();
 sg13g2_decap_8 FILLER_35_802 ();
 sg13g2_decap_8 FILLER_35_809 ();
 sg13g2_decap_8 FILLER_35_816 ();
 sg13g2_decap_8 FILLER_35_823 ();
 sg13g2_decap_8 FILLER_35_830 ();
 sg13g2_decap_8 FILLER_35_837 ();
 sg13g2_decap_8 FILLER_35_844 ();
 sg13g2_decap_8 FILLER_35_851 ();
 sg13g2_decap_4 FILLER_35_858 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_4 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_18 ();
 sg13g2_fill_2 FILLER_36_54 ();
 sg13g2_fill_1 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_fill_1 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_145 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_234 ();
 sg13g2_fill_2 FILLER_36_250 ();
 sg13g2_fill_2 FILLER_36_297 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_fill_2 FILLER_36_380 ();
 sg13g2_fill_2 FILLER_36_391 ();
 sg13g2_fill_1 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_424 ();
 sg13g2_fill_1 FILLER_36_431 ();
 sg13g2_decap_8 FILLER_36_445 ();
 sg13g2_decap_4 FILLER_36_452 ();
 sg13g2_fill_2 FILLER_36_456 ();
 sg13g2_decap_4 FILLER_36_468 ();
 sg13g2_fill_2 FILLER_36_472 ();
 sg13g2_fill_2 FILLER_36_478 ();
 sg13g2_decap_8 FILLER_36_488 ();
 sg13g2_decap_8 FILLER_36_495 ();
 sg13g2_fill_1 FILLER_36_502 ();
 sg13g2_fill_1 FILLER_36_520 ();
 sg13g2_fill_2 FILLER_36_547 ();
 sg13g2_fill_2 FILLER_36_583 ();
 sg13g2_fill_1 FILLER_36_601 ();
 sg13g2_decap_8 FILLER_36_614 ();
 sg13g2_decap_8 FILLER_36_621 ();
 sg13g2_fill_1 FILLER_36_640 ();
 sg13g2_fill_1 FILLER_36_646 ();
 sg13g2_fill_2 FILLER_36_656 ();
 sg13g2_fill_1 FILLER_36_658 ();
 sg13g2_fill_2 FILLER_36_676 ();
 sg13g2_decap_4 FILLER_36_687 ();
 sg13g2_fill_2 FILLER_36_704 ();
 sg13g2_fill_1 FILLER_36_706 ();
 sg13g2_decap_4 FILLER_36_732 ();
 sg13g2_fill_1 FILLER_36_736 ();
 sg13g2_fill_1 FILLER_36_750 ();
 sg13g2_fill_2 FILLER_36_756 ();
 sg13g2_fill_1 FILLER_36_758 ();
 sg13g2_decap_8 FILLER_36_768 ();
 sg13g2_decap_8 FILLER_36_775 ();
 sg13g2_decap_8 FILLER_36_782 ();
 sg13g2_decap_8 FILLER_36_789 ();
 sg13g2_decap_8 FILLER_36_796 ();
 sg13g2_decap_8 FILLER_36_803 ();
 sg13g2_decap_8 FILLER_36_810 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_decap_8 FILLER_36_824 ();
 sg13g2_decap_8 FILLER_36_831 ();
 sg13g2_decap_8 FILLER_36_838 ();
 sg13g2_decap_8 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_852 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_1 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_33 ();
 sg13g2_decap_4 FILLER_37_40 ();
 sg13g2_fill_2 FILLER_37_74 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_fill_2 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_144 ();
 sg13g2_decap_4 FILLER_37_180 ();
 sg13g2_fill_1 FILLER_37_184 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_201 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_210 ();
 sg13g2_decap_4 FILLER_37_224 ();
 sg13g2_fill_2 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_1 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_fill_2 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_388 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_fill_1 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_414 ();
 sg13g2_fill_2 FILLER_37_429 ();
 sg13g2_fill_1 FILLER_37_431 ();
 sg13g2_fill_2 FILLER_37_461 ();
 sg13g2_fill_1 FILLER_37_463 ();
 sg13g2_fill_1 FILLER_37_472 ();
 sg13g2_decap_8 FILLER_37_486 ();
 sg13g2_fill_1 FILLER_37_493 ();
 sg13g2_fill_2 FILLER_37_510 ();
 sg13g2_fill_2 FILLER_37_516 ();
 sg13g2_fill_2 FILLER_37_540 ();
 sg13g2_fill_1 FILLER_37_542 ();
 sg13g2_fill_1 FILLER_37_552 ();
 sg13g2_fill_1 FILLER_37_563 ();
 sg13g2_fill_2 FILLER_37_604 ();
 sg13g2_fill_1 FILLER_37_661 ();
 sg13g2_fill_1 FILLER_37_685 ();
 sg13g2_fill_2 FILLER_37_717 ();
 sg13g2_decap_8 FILLER_37_773 ();
 sg13g2_decap_8 FILLER_37_780 ();
 sg13g2_decap_8 FILLER_37_787 ();
 sg13g2_decap_8 FILLER_37_794 ();
 sg13g2_decap_8 FILLER_37_801 ();
 sg13g2_decap_8 FILLER_37_808 ();
 sg13g2_decap_8 FILLER_37_815 ();
 sg13g2_decap_8 FILLER_37_822 ();
 sg13g2_decap_8 FILLER_37_829 ();
 sg13g2_decap_8 FILLER_37_836 ();
 sg13g2_decap_8 FILLER_37_843 ();
 sg13g2_decap_8 FILLER_37_850 ();
 sg13g2_decap_4 FILLER_37_857 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_37 ();
 sg13g2_fill_2 FILLER_38_105 ();
 sg13g2_fill_1 FILLER_38_107 ();
 sg13g2_fill_2 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_125 ();
 sg13g2_fill_1 FILLER_38_132 ();
 sg13g2_fill_2 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_144 ();
 sg13g2_fill_1 FILLER_38_160 ();
 sg13g2_fill_1 FILLER_38_170 ();
 sg13g2_decap_4 FILLER_38_184 ();
 sg13g2_fill_1 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_214 ();
 sg13g2_decap_4 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_225 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_280 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_decap_4 FILLER_38_351 ();
 sg13g2_fill_1 FILLER_38_371 ();
 sg13g2_fill_1 FILLER_38_380 ();
 sg13g2_decap_4 FILLER_38_402 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_429 ();
 sg13g2_decap_4 FILLER_38_436 ();
 sg13g2_fill_1 FILLER_38_444 ();
 sg13g2_decap_4 FILLER_38_462 ();
 sg13g2_fill_1 FILLER_38_466 ();
 sg13g2_decap_8 FILLER_38_483 ();
 sg13g2_decap_8 FILLER_38_490 ();
 sg13g2_fill_2 FILLER_38_528 ();
 sg13g2_fill_1 FILLER_38_530 ();
 sg13g2_fill_2 FILLER_38_561 ();
 sg13g2_fill_1 FILLER_38_571 ();
 sg13g2_fill_1 FILLER_38_577 ();
 sg13g2_fill_2 FILLER_38_586 ();
 sg13g2_fill_1 FILLER_38_588 ();
 sg13g2_fill_1 FILLER_38_598 ();
 sg13g2_decap_4 FILLER_38_625 ();
 sg13g2_fill_1 FILLER_38_652 ();
 sg13g2_decap_4 FILLER_38_674 ();
 sg13g2_fill_2 FILLER_38_678 ();
 sg13g2_decap_4 FILLER_38_685 ();
 sg13g2_fill_1 FILLER_38_689 ();
 sg13g2_fill_2 FILLER_38_734 ();
 sg13g2_decap_4 FILLER_38_746 ();
 sg13g2_fill_2 FILLER_38_759 ();
 sg13g2_fill_1 FILLER_38_761 ();
 sg13g2_decap_8 FILLER_38_775 ();
 sg13g2_decap_8 FILLER_38_782 ();
 sg13g2_decap_8 FILLER_38_789 ();
 sg13g2_decap_8 FILLER_38_796 ();
 sg13g2_decap_8 FILLER_38_803 ();
 sg13g2_decap_8 FILLER_38_810 ();
 sg13g2_decap_8 FILLER_38_817 ();
 sg13g2_decap_8 FILLER_38_824 ();
 sg13g2_decap_8 FILLER_38_831 ();
 sg13g2_decap_8 FILLER_38_838 ();
 sg13g2_decap_8 FILLER_38_845 ();
 sg13g2_decap_8 FILLER_38_852 ();
 sg13g2_fill_2 FILLER_38_859 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_4 FILLER_39_35 ();
 sg13g2_fill_1 FILLER_39_39 ();
 sg13g2_fill_2 FILLER_39_66 ();
 sg13g2_fill_1 FILLER_39_68 ();
 sg13g2_fill_2 FILLER_39_83 ();
 sg13g2_fill_2 FILLER_39_107 ();
 sg13g2_fill_1 FILLER_39_109 ();
 sg13g2_fill_2 FILLER_39_124 ();
 sg13g2_decap_4 FILLER_39_189 ();
 sg13g2_fill_2 FILLER_39_219 ();
 sg13g2_fill_1 FILLER_39_221 ();
 sg13g2_fill_2 FILLER_39_232 ();
 sg13g2_fill_2 FILLER_39_257 ();
 sg13g2_fill_2 FILLER_39_319 ();
 sg13g2_fill_1 FILLER_39_321 ();
 sg13g2_fill_2 FILLER_39_327 ();
 sg13g2_decap_8 FILLER_39_339 ();
 sg13g2_decap_4 FILLER_39_346 ();
 sg13g2_fill_1 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_355 ();
 sg13g2_fill_1 FILLER_39_362 ();
 sg13g2_fill_2 FILLER_39_370 ();
 sg13g2_fill_1 FILLER_39_372 ();
 sg13g2_fill_2 FILLER_39_389 ();
 sg13g2_fill_2 FILLER_39_396 ();
 sg13g2_fill_1 FILLER_39_398 ();
 sg13g2_decap_8 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_432 ();
 sg13g2_fill_1 FILLER_39_437 ();
 sg13g2_fill_2 FILLER_39_455 ();
 sg13g2_fill_2 FILLER_39_512 ();
 sg13g2_fill_1 FILLER_39_514 ();
 sg13g2_fill_2 FILLER_39_536 ();
 sg13g2_fill_1 FILLER_39_538 ();
 sg13g2_fill_2 FILLER_39_599 ();
 sg13g2_fill_2 FILLER_39_614 ();
 sg13g2_fill_2 FILLER_39_677 ();
 sg13g2_decap_4 FILLER_39_718 ();
 sg13g2_fill_2 FILLER_39_749 ();
 sg13g2_fill_1 FILLER_39_751 ();
 sg13g2_decap_8 FILLER_39_778 ();
 sg13g2_decap_8 FILLER_39_785 ();
 sg13g2_decap_8 FILLER_39_792 ();
 sg13g2_decap_8 FILLER_39_799 ();
 sg13g2_decap_8 FILLER_39_806 ();
 sg13g2_decap_8 FILLER_39_813 ();
 sg13g2_decap_8 FILLER_39_820 ();
 sg13g2_decap_8 FILLER_39_827 ();
 sg13g2_decap_8 FILLER_39_834 ();
 sg13g2_decap_8 FILLER_39_841 ();
 sg13g2_decap_8 FILLER_39_848 ();
 sg13g2_decap_8 FILLER_39_855 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_fill_1 FILLER_40_75 ();
 sg13g2_fill_2 FILLER_40_85 ();
 sg13g2_fill_1 FILLER_40_87 ();
 sg13g2_fill_2 FILLER_40_102 ();
 sg13g2_fill_2 FILLER_40_139 ();
 sg13g2_fill_1 FILLER_40_141 ();
 sg13g2_fill_1 FILLER_40_180 ();
 sg13g2_decap_4 FILLER_40_188 ();
 sg13g2_fill_1 FILLER_40_192 ();
 sg13g2_fill_1 FILLER_40_211 ();
 sg13g2_fill_2 FILLER_40_229 ();
 sg13g2_fill_1 FILLER_40_243 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_fill_2 FILLER_40_314 ();
 sg13g2_fill_1 FILLER_40_316 ();
 sg13g2_fill_1 FILLER_40_326 ();
 sg13g2_decap_4 FILLER_40_336 ();
 sg13g2_fill_2 FILLER_40_379 ();
 sg13g2_decap_8 FILLER_40_393 ();
 sg13g2_fill_2 FILLER_40_400 ();
 sg13g2_fill_1 FILLER_40_402 ();
 sg13g2_decap_8 FILLER_40_417 ();
 sg13g2_fill_1 FILLER_40_424 ();
 sg13g2_decap_8 FILLER_40_438 ();
 sg13g2_decap_8 FILLER_40_445 ();
 sg13g2_decap_8 FILLER_40_452 ();
 sg13g2_fill_2 FILLER_40_464 ();
 sg13g2_fill_1 FILLER_40_466 ();
 sg13g2_fill_1 FILLER_40_480 ();
 sg13g2_fill_2 FILLER_40_508 ();
 sg13g2_fill_2 FILLER_40_540 ();
 sg13g2_fill_1 FILLER_40_556 ();
 sg13g2_fill_1 FILLER_40_565 ();
 sg13g2_decap_8 FILLER_40_571 ();
 sg13g2_decap_8 FILLER_40_578 ();
 sg13g2_fill_1 FILLER_40_585 ();
 sg13g2_fill_1 FILLER_40_595 ();
 sg13g2_fill_1 FILLER_40_601 ();
 sg13g2_decap_8 FILLER_40_611 ();
 sg13g2_decap_8 FILLER_40_618 ();
 sg13g2_decap_4 FILLER_40_625 ();
 sg13g2_fill_2 FILLER_40_634 ();
 sg13g2_decap_4 FILLER_40_640 ();
 sg13g2_fill_2 FILLER_40_644 ();
 sg13g2_decap_4 FILLER_40_655 ();
 sg13g2_fill_1 FILLER_40_659 ();
 sg13g2_decap_4 FILLER_40_664 ();
 sg13g2_fill_1 FILLER_40_668 ();
 sg13g2_decap_4 FILLER_40_733 ();
 sg13g2_fill_1 FILLER_40_742 ();
 sg13g2_fill_1 FILLER_40_753 ();
 sg13g2_decap_8 FILLER_40_767 ();
 sg13g2_decap_8 FILLER_40_774 ();
 sg13g2_decap_8 FILLER_40_781 ();
 sg13g2_decap_8 FILLER_40_788 ();
 sg13g2_decap_8 FILLER_40_795 ();
 sg13g2_decap_8 FILLER_40_802 ();
 sg13g2_decap_8 FILLER_40_809 ();
 sg13g2_decap_8 FILLER_40_816 ();
 sg13g2_decap_8 FILLER_40_823 ();
 sg13g2_decap_8 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_40_837 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_4 FILLER_40_858 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_fill_2 FILLER_41_56 ();
 sg13g2_fill_2 FILLER_41_88 ();
 sg13g2_fill_2 FILLER_41_105 ();
 sg13g2_fill_2 FILLER_41_126 ();
 sg13g2_fill_1 FILLER_41_128 ();
 sg13g2_fill_2 FILLER_41_186 ();
 sg13g2_fill_2 FILLER_41_332 ();
 sg13g2_fill_2 FILLER_41_360 ();
 sg13g2_fill_1 FILLER_41_362 ();
 sg13g2_decap_4 FILLER_41_375 ();
 sg13g2_decap_4 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_429 ();
 sg13g2_fill_2 FILLER_41_436 ();
 sg13g2_fill_2 FILLER_41_442 ();
 sg13g2_decap_4 FILLER_41_448 ();
 sg13g2_fill_2 FILLER_41_452 ();
 sg13g2_fill_2 FILLER_41_480 ();
 sg13g2_fill_2 FILLER_41_508 ();
 sg13g2_fill_1 FILLER_41_591 ();
 sg13g2_fill_1 FILLER_41_639 ();
 sg13g2_fill_2 FILLER_41_645 ();
 sg13g2_fill_1 FILLER_41_647 ();
 sg13g2_fill_1 FILLER_41_684 ();
 sg13g2_decap_4 FILLER_41_711 ();
 sg13g2_fill_2 FILLER_41_715 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_fill_2 FILLER_41_728 ();
 sg13g2_fill_1 FILLER_41_730 ();
 sg13g2_fill_2 FILLER_41_758 ();
 sg13g2_decap_8 FILLER_41_773 ();
 sg13g2_decap_8 FILLER_41_780 ();
 sg13g2_decap_8 FILLER_41_787 ();
 sg13g2_decap_8 FILLER_41_794 ();
 sg13g2_decap_8 FILLER_41_801 ();
 sg13g2_decap_8 FILLER_41_808 ();
 sg13g2_decap_8 FILLER_41_815 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_decap_8 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_850 ();
 sg13g2_decap_4 FILLER_41_857 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_fill_2 FILLER_42_63 ();
 sg13g2_fill_2 FILLER_42_77 ();
 sg13g2_fill_1 FILLER_42_79 ();
 sg13g2_decap_4 FILLER_42_143 ();
 sg13g2_fill_2 FILLER_42_190 ();
 sg13g2_fill_1 FILLER_42_192 ();
 sg13g2_fill_2 FILLER_42_197 ();
 sg13g2_fill_2 FILLER_42_203 ();
 sg13g2_fill_2 FILLER_42_248 ();
 sg13g2_fill_1 FILLER_42_250 ();
 sg13g2_fill_1 FILLER_42_256 ();
 sg13g2_decap_4 FILLER_42_278 ();
 sg13g2_fill_2 FILLER_42_282 ();
 sg13g2_decap_4 FILLER_42_287 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_fill_1 FILLER_42_323 ();
 sg13g2_fill_1 FILLER_42_331 ();
 sg13g2_fill_2 FILLER_42_341 ();
 sg13g2_fill_1 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_352 ();
 sg13g2_decap_8 FILLER_42_359 ();
 sg13g2_decap_4 FILLER_42_366 ();
 sg13g2_decap_8 FILLER_42_403 ();
 sg13g2_fill_1 FILLER_42_414 ();
 sg13g2_fill_2 FILLER_42_419 ();
 sg13g2_fill_2 FILLER_42_426 ();
 sg13g2_decap_4 FILLER_42_459 ();
 sg13g2_fill_2 FILLER_42_463 ();
 sg13g2_fill_2 FILLER_42_469 ();
 sg13g2_fill_1 FILLER_42_471 ();
 sg13g2_fill_2 FILLER_42_490 ();
 sg13g2_fill_1 FILLER_42_492 ();
 sg13g2_fill_1 FILLER_42_497 ();
 sg13g2_fill_2 FILLER_42_502 ();
 sg13g2_decap_4 FILLER_42_513 ();
 sg13g2_fill_1 FILLER_42_517 ();
 sg13g2_fill_2 FILLER_42_544 ();
 sg13g2_decap_8 FILLER_42_577 ();
 sg13g2_fill_1 FILLER_42_584 ();
 sg13g2_fill_1 FILLER_42_593 ();
 sg13g2_decap_8 FILLER_42_604 ();
 sg13g2_fill_2 FILLER_42_615 ();
 sg13g2_fill_1 FILLER_42_617 ();
 sg13g2_fill_1 FILLER_42_658 ();
 sg13g2_fill_2 FILLER_42_664 ();
 sg13g2_fill_1 FILLER_42_691 ();
 sg13g2_fill_2 FILLER_42_696 ();
 sg13g2_fill_2 FILLER_42_733 ();
 sg13g2_decap_8 FILLER_42_775 ();
 sg13g2_decap_8 FILLER_42_782 ();
 sg13g2_decap_8 FILLER_42_789 ();
 sg13g2_decap_8 FILLER_42_796 ();
 sg13g2_decap_8 FILLER_42_803 ();
 sg13g2_decap_8 FILLER_42_810 ();
 sg13g2_decap_8 FILLER_42_817 ();
 sg13g2_decap_8 FILLER_42_824 ();
 sg13g2_decap_8 FILLER_42_831 ();
 sg13g2_decap_8 FILLER_42_838 ();
 sg13g2_decap_8 FILLER_42_845 ();
 sg13g2_decap_8 FILLER_42_852 ();
 sg13g2_fill_2 FILLER_42_859 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_fill_2 FILLER_43_63 ();
 sg13g2_fill_1 FILLER_43_65 ();
 sg13g2_fill_1 FILLER_43_113 ();
 sg13g2_fill_1 FILLER_43_122 ();
 sg13g2_fill_1 FILLER_43_131 ();
 sg13g2_fill_2 FILLER_43_163 ();
 sg13g2_fill_2 FILLER_43_174 ();
 sg13g2_fill_1 FILLER_43_176 ();
 sg13g2_fill_1 FILLER_43_208 ();
 sg13g2_fill_2 FILLER_43_213 ();
 sg13g2_fill_1 FILLER_43_215 ();
 sg13g2_fill_1 FILLER_43_220 ();
 sg13g2_decap_4 FILLER_43_225 ();
 sg13g2_fill_1 FILLER_43_229 ();
 sg13g2_fill_2 FILLER_43_247 ();
 sg13g2_fill_1 FILLER_43_310 ();
 sg13g2_decap_4 FILLER_43_401 ();
 sg13g2_fill_2 FILLER_43_435 ();
 sg13g2_fill_2 FILLER_43_463 ();
 sg13g2_fill_1 FILLER_43_465 ();
 sg13g2_fill_1 FILLER_43_484 ();
 sg13g2_decap_8 FILLER_43_495 ();
 sg13g2_fill_2 FILLER_43_543 ();
 sg13g2_fill_1 FILLER_43_545 ();
 sg13g2_decap_4 FILLER_43_607 ();
 sg13g2_fill_2 FILLER_43_637 ();
 sg13g2_fill_2 FILLER_43_662 ();
 sg13g2_fill_1 FILLER_43_664 ();
 sg13g2_decap_4 FILLER_43_678 ();
 sg13g2_fill_1 FILLER_43_687 ();
 sg13g2_fill_2 FILLER_43_700 ();
 sg13g2_decap_4 FILLER_43_711 ();
 sg13g2_fill_2 FILLER_43_733 ();
 sg13g2_fill_1 FILLER_43_739 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_4 FILLER_44_81 ();
 sg13g2_fill_1 FILLER_44_85 ();
 sg13g2_fill_2 FILLER_44_125 ();
 sg13g2_fill_1 FILLER_44_127 ();
 sg13g2_fill_1 FILLER_44_140 ();
 sg13g2_fill_1 FILLER_44_196 ();
 sg13g2_fill_2 FILLER_44_236 ();
 sg13g2_fill_2 FILLER_44_292 ();
 sg13g2_fill_1 FILLER_44_334 ();
 sg13g2_fill_2 FILLER_44_358 ();
 sg13g2_fill_1 FILLER_44_360 ();
 sg13g2_decap_8 FILLER_44_369 ();
 sg13g2_decap_8 FILLER_44_376 ();
 sg13g2_fill_2 FILLER_44_383 ();
 sg13g2_decap_4 FILLER_44_411 ();
 sg13g2_fill_2 FILLER_44_415 ();
 sg13g2_fill_1 FILLER_44_430 ();
 sg13g2_fill_2 FILLER_44_440 ();
 sg13g2_fill_1 FILLER_44_442 ();
 sg13g2_fill_1 FILLER_44_499 ();
 sg13g2_fill_1 FILLER_44_518 ();
 sg13g2_fill_1 FILLER_44_524 ();
 sg13g2_fill_2 FILLER_44_551 ();
 sg13g2_fill_1 FILLER_44_553 ();
 sg13g2_fill_1 FILLER_44_563 ();
 sg13g2_fill_2 FILLER_44_569 ();
 sg13g2_fill_2 FILLER_44_592 ();
 sg13g2_decap_8 FILLER_44_608 ();
 sg13g2_decap_4 FILLER_44_615 ();
 sg13g2_fill_1 FILLER_44_619 ();
 sg13g2_fill_2 FILLER_44_633 ();
 sg13g2_fill_1 FILLER_44_635 ();
 sg13g2_fill_1 FILLER_44_655 ();
 sg13g2_fill_2 FILLER_44_682 ();
 sg13g2_fill_1 FILLER_44_684 ();
 sg13g2_fill_1 FILLER_44_735 ();
 sg13g2_fill_2 FILLER_44_744 ();
 sg13g2_fill_1 FILLER_44_746 ();
 sg13g2_decap_8 FILLER_44_773 ();
 sg13g2_decap_8 FILLER_44_780 ();
 sg13g2_decap_8 FILLER_44_787 ();
 sg13g2_decap_8 FILLER_44_794 ();
 sg13g2_decap_8 FILLER_44_801 ();
 sg13g2_decap_8 FILLER_44_808 ();
 sg13g2_decap_8 FILLER_44_815 ();
 sg13g2_decap_8 FILLER_44_822 ();
 sg13g2_decap_8 FILLER_44_829 ();
 sg13g2_decap_8 FILLER_44_836 ();
 sg13g2_decap_8 FILLER_44_843 ();
 sg13g2_decap_8 FILLER_44_850 ();
 sg13g2_decap_4 FILLER_44_857 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_fill_2 FILLER_45_77 ();
 sg13g2_decap_4 FILLER_45_83 ();
 sg13g2_fill_2 FILLER_45_96 ();
 sg13g2_fill_1 FILLER_45_103 ();
 sg13g2_decap_8 FILLER_45_207 ();
 sg13g2_decap_8 FILLER_45_214 ();
 sg13g2_decap_8 FILLER_45_221 ();
 sg13g2_decap_8 FILLER_45_228 ();
 sg13g2_decap_4 FILLER_45_235 ();
 sg13g2_fill_2 FILLER_45_239 ();
 sg13g2_decap_4 FILLER_45_245 ();
 sg13g2_fill_1 FILLER_45_253 ();
 sg13g2_fill_1 FILLER_45_309 ();
 sg13g2_fill_2 FILLER_45_391 ();
 sg13g2_fill_1 FILLER_45_393 ();
 sg13g2_fill_2 FILLER_45_403 ();
 sg13g2_fill_1 FILLER_45_405 ();
 sg13g2_fill_2 FILLER_45_435 ();
 sg13g2_fill_1 FILLER_45_469 ();
 sg13g2_fill_1 FILLER_45_498 ();
 sg13g2_fill_2 FILLER_45_513 ();
 sg13g2_fill_1 FILLER_45_515 ();
 sg13g2_decap_8 FILLER_45_623 ();
 sg13g2_fill_1 FILLER_45_630 ();
 sg13g2_fill_2 FILLER_45_636 ();
 sg13g2_fill_1 FILLER_45_638 ();
 sg13g2_fill_1 FILLER_45_652 ();
 sg13g2_fill_2 FILLER_45_670 ();
 sg13g2_fill_1 FILLER_45_672 ();
 sg13g2_decap_4 FILLER_45_682 ();
 sg13g2_decap_4 FILLER_45_691 ();
 sg13g2_fill_1 FILLER_45_695 ();
 sg13g2_fill_2 FILLER_45_700 ();
 sg13g2_fill_2 FILLER_45_728 ();
 sg13g2_fill_2 FILLER_45_745 ();
 sg13g2_fill_1 FILLER_45_747 ();
 sg13g2_fill_1 FILLER_45_757 ();
 sg13g2_decap_8 FILLER_45_771 ();
 sg13g2_decap_8 FILLER_45_778 ();
 sg13g2_decap_8 FILLER_45_785 ();
 sg13g2_decap_8 FILLER_45_792 ();
 sg13g2_decap_8 FILLER_45_799 ();
 sg13g2_decap_8 FILLER_45_806 ();
 sg13g2_decap_8 FILLER_45_813 ();
 sg13g2_decap_8 FILLER_45_820 ();
 sg13g2_decap_8 FILLER_45_827 ();
 sg13g2_decap_8 FILLER_45_834 ();
 sg13g2_decap_8 FILLER_45_841 ();
 sg13g2_decap_8 FILLER_45_848 ();
 sg13g2_decap_8 FILLER_45_855 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_fill_2 FILLER_46_91 ();
 sg13g2_decap_4 FILLER_46_102 ();
 sg13g2_fill_2 FILLER_46_115 ();
 sg13g2_fill_2 FILLER_46_147 ();
 sg13g2_fill_1 FILLER_46_149 ();
 sg13g2_fill_2 FILLER_46_159 ();
 sg13g2_decap_8 FILLER_46_201 ();
 sg13g2_decap_8 FILLER_46_208 ();
 sg13g2_decap_8 FILLER_46_215 ();
 sg13g2_decap_8 FILLER_46_222 ();
 sg13g2_fill_1 FILLER_46_229 ();
 sg13g2_fill_1 FILLER_46_300 ();
 sg13g2_fill_1 FILLER_46_312 ();
 sg13g2_fill_1 FILLER_46_332 ();
 sg13g2_fill_1 FILLER_46_347 ();
 sg13g2_decap_8 FILLER_46_367 ();
 sg13g2_decap_8 FILLER_46_444 ();
 sg13g2_decap_8 FILLER_46_451 ();
 sg13g2_fill_1 FILLER_46_458 ();
 sg13g2_fill_2 FILLER_46_498 ();
 sg13g2_decap_8 FILLER_46_531 ();
 sg13g2_fill_1 FILLER_46_538 ();
 sg13g2_fill_1 FILLER_46_547 ();
 sg13g2_fill_2 FILLER_46_557 ();
 sg13g2_fill_1 FILLER_46_559 ();
 sg13g2_fill_2 FILLER_46_577 ();
 sg13g2_fill_1 FILLER_46_579 ();
 sg13g2_decap_4 FILLER_46_589 ();
 sg13g2_fill_1 FILLER_46_616 ();
 sg13g2_fill_2 FILLER_46_652 ();
 sg13g2_fill_1 FILLER_46_654 ();
 sg13g2_decap_8 FILLER_46_696 ();
 sg13g2_decap_8 FILLER_46_703 ();
 sg13g2_fill_1 FILLER_46_723 ();
 sg13g2_fill_2 FILLER_46_729 ();
 sg13g2_fill_1 FILLER_46_741 ();
 sg13g2_decap_8 FILLER_46_765 ();
 sg13g2_decap_8 FILLER_46_772 ();
 sg13g2_decap_8 FILLER_46_779 ();
 sg13g2_decap_8 FILLER_46_786 ();
 sg13g2_decap_8 FILLER_46_793 ();
 sg13g2_decap_8 FILLER_46_800 ();
 sg13g2_decap_8 FILLER_46_807 ();
 sg13g2_decap_8 FILLER_46_814 ();
 sg13g2_decap_8 FILLER_46_821 ();
 sg13g2_decap_8 FILLER_46_828 ();
 sg13g2_decap_8 FILLER_46_835 ();
 sg13g2_decap_8 FILLER_46_842 ();
 sg13g2_decap_8 FILLER_46_849 ();
 sg13g2_decap_4 FILLER_46_856 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_fill_1 FILLER_47_119 ();
 sg13g2_fill_1 FILLER_47_172 ();
 sg13g2_decap_8 FILLER_47_190 ();
 sg13g2_decap_8 FILLER_47_197 ();
 sg13g2_decap_8 FILLER_47_204 ();
 sg13g2_decap_8 FILLER_47_211 ();
 sg13g2_decap_8 FILLER_47_218 ();
 sg13g2_decap_8 FILLER_47_225 ();
 sg13g2_decap_8 FILLER_47_232 ();
 sg13g2_decap_8 FILLER_47_239 ();
 sg13g2_fill_1 FILLER_47_246 ();
 sg13g2_fill_1 FILLER_47_273 ();
 sg13g2_fill_2 FILLER_47_283 ();
 sg13g2_fill_1 FILLER_47_285 ();
 sg13g2_decap_4 FILLER_47_291 ();
 sg13g2_fill_1 FILLER_47_295 ();
 sg13g2_fill_2 FILLER_47_345 ();
 sg13g2_fill_1 FILLER_47_347 ();
 sg13g2_fill_1 FILLER_47_365 ();
 sg13g2_fill_1 FILLER_47_384 ();
 sg13g2_fill_2 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_425 ();
 sg13g2_fill_1 FILLER_47_435 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_fill_2 FILLER_47_469 ();
 sg13g2_fill_1 FILLER_47_471 ();
 sg13g2_fill_2 FILLER_47_500 ();
 sg13g2_fill_1 FILLER_47_502 ();
 sg13g2_fill_2 FILLER_47_534 ();
 sg13g2_fill_1 FILLER_47_536 ();
 sg13g2_fill_2 FILLER_47_547 ();
 sg13g2_fill_1 FILLER_47_596 ();
 sg13g2_decap_4 FILLER_47_623 ();
 sg13g2_fill_1 FILLER_47_627 ();
 sg13g2_fill_2 FILLER_47_632 ();
 sg13g2_fill_1 FILLER_47_638 ();
 sg13g2_fill_2 FILLER_47_648 ();
 sg13g2_fill_1 FILLER_47_739 ();
 sg13g2_decap_8 FILLER_47_766 ();
 sg13g2_decap_8 FILLER_47_773 ();
 sg13g2_decap_8 FILLER_47_780 ();
 sg13g2_decap_8 FILLER_47_787 ();
 sg13g2_decap_8 FILLER_47_794 ();
 sg13g2_decap_8 FILLER_47_801 ();
 sg13g2_decap_8 FILLER_47_808 ();
 sg13g2_decap_8 FILLER_47_815 ();
 sg13g2_decap_8 FILLER_47_822 ();
 sg13g2_decap_8 FILLER_47_829 ();
 sg13g2_decap_8 FILLER_47_836 ();
 sg13g2_decap_8 FILLER_47_843 ();
 sg13g2_decap_8 FILLER_47_850 ();
 sg13g2_decap_4 FILLER_47_857 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_4 FILLER_48_126 ();
 sg13g2_fill_2 FILLER_48_130 ();
 sg13g2_fill_2 FILLER_48_136 ();
 sg13g2_fill_2 FILLER_48_147 ();
 sg13g2_fill_2 FILLER_48_154 ();
 sg13g2_fill_1 FILLER_48_156 ();
 sg13g2_fill_1 FILLER_48_161 ();
 sg13g2_fill_1 FILLER_48_176 ();
 sg13g2_fill_1 FILLER_48_194 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_4 FILLER_48_245 ();
 sg13g2_fill_2 FILLER_48_249 ();
 sg13g2_fill_1 FILLER_48_268 ();
 sg13g2_decap_4 FILLER_48_314 ();
 sg13g2_fill_1 FILLER_48_326 ();
 sg13g2_fill_1 FILLER_48_452 ();
 sg13g2_fill_2 FILLER_48_479 ();
 sg13g2_decap_4 FILLER_48_506 ();
 sg13g2_decap_4 FILLER_48_514 ();
 sg13g2_fill_1 FILLER_48_518 ();
 sg13g2_fill_2 FILLER_48_532 ();
 sg13g2_fill_1 FILLER_48_581 ();
 sg13g2_fill_1 FILLER_48_587 ();
 sg13g2_fill_2 FILLER_48_593 ();
 sg13g2_fill_1 FILLER_48_595 ();
 sg13g2_fill_2 FILLER_48_610 ();
 sg13g2_decap_8 FILLER_48_656 ();
 sg13g2_fill_2 FILLER_48_663 ();
 sg13g2_fill_1 FILLER_48_665 ();
 sg13g2_decap_4 FILLER_48_697 ();
 sg13g2_fill_2 FILLER_48_748 ();
 sg13g2_fill_1 FILLER_48_750 ();
 sg13g2_decap_8 FILLER_48_765 ();
 sg13g2_decap_8 FILLER_48_772 ();
 sg13g2_decap_8 FILLER_48_779 ();
 sg13g2_decap_8 FILLER_48_786 ();
 sg13g2_decap_8 FILLER_48_793 ();
 sg13g2_decap_8 FILLER_48_800 ();
 sg13g2_decap_8 FILLER_48_807 ();
 sg13g2_decap_8 FILLER_48_814 ();
 sg13g2_decap_8 FILLER_48_821 ();
 sg13g2_decap_8 FILLER_48_828 ();
 sg13g2_decap_8 FILLER_48_835 ();
 sg13g2_decap_8 FILLER_48_842 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_decap_4 FILLER_48_856 ();
 sg13g2_fill_2 FILLER_48_860 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_4 FILLER_49_140 ();
 sg13g2_fill_2 FILLER_49_167 ();
 sg13g2_fill_1 FILLER_49_169 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_fill_1 FILLER_49_258 ();
 sg13g2_decap_4 FILLER_49_288 ();
 sg13g2_fill_1 FILLER_49_292 ();
 sg13g2_fill_2 FILLER_49_315 ();
 sg13g2_fill_2 FILLER_49_326 ();
 sg13g2_fill_1 FILLER_49_328 ();
 sg13g2_fill_2 FILLER_49_343 ();
 sg13g2_fill_1 FILLER_49_345 ();
 sg13g2_fill_1 FILLER_49_360 ();
 sg13g2_decap_8 FILLER_49_380 ();
 sg13g2_decap_4 FILLER_49_387 ();
 sg13g2_decap_4 FILLER_49_409 ();
 sg13g2_fill_1 FILLER_49_433 ();
 sg13g2_decap_8 FILLER_49_453 ();
 sg13g2_fill_2 FILLER_49_460 ();
 sg13g2_fill_1 FILLER_49_462 ();
 sg13g2_fill_1 FILLER_49_486 ();
 sg13g2_fill_2 FILLER_49_497 ();
 sg13g2_fill_1 FILLER_49_499 ();
 sg13g2_fill_1 FILLER_49_512 ();
 sg13g2_decap_4 FILLER_49_522 ();
 sg13g2_fill_2 FILLER_49_526 ();
 sg13g2_fill_2 FILLER_49_591 ();
 sg13g2_fill_2 FILLER_49_598 ();
 sg13g2_fill_1 FILLER_49_600 ();
 sg13g2_fill_2 FILLER_49_635 ();
 sg13g2_fill_1 FILLER_49_637 ();
 sg13g2_fill_1 FILLER_49_643 ();
 sg13g2_fill_1 FILLER_49_695 ();
 sg13g2_fill_1 FILLER_49_704 ();
 sg13g2_decap_4 FILLER_49_724 ();
 sg13g2_fill_1 FILLER_49_728 ();
 sg13g2_fill_1 FILLER_49_734 ();
 sg13g2_fill_1 FILLER_49_740 ();
 sg13g2_fill_1 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_783 ();
 sg13g2_decap_8 FILLER_49_790 ();
 sg13g2_decap_8 FILLER_49_797 ();
 sg13g2_decap_8 FILLER_49_804 ();
 sg13g2_decap_8 FILLER_49_811 ();
 sg13g2_decap_8 FILLER_49_818 ();
 sg13g2_decap_8 FILLER_49_825 ();
 sg13g2_decap_8 FILLER_49_832 ();
 sg13g2_decap_8 FILLER_49_839 ();
 sg13g2_decap_8 FILLER_49_846 ();
 sg13g2_decap_8 FILLER_49_853 ();
 sg13g2_fill_2 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_4 FILLER_50_140 ();
 sg13g2_fill_1 FILLER_50_144 ();
 sg13g2_fill_1 FILLER_50_184 ();
 sg13g2_decap_4 FILLER_50_229 ();
 sg13g2_decap_4 FILLER_50_237 ();
 sg13g2_fill_1 FILLER_50_241 ();
 sg13g2_fill_1 FILLER_50_296 ();
 sg13g2_fill_2 FILLER_50_349 ();
 sg13g2_fill_1 FILLER_50_351 ();
 sg13g2_fill_2 FILLER_50_431 ();
 sg13g2_decap_8 FILLER_50_459 ();
 sg13g2_fill_2 FILLER_50_466 ();
 sg13g2_fill_1 FILLER_50_468 ();
 sg13g2_fill_1 FILLER_50_474 ();
 sg13g2_decap_8 FILLER_50_479 ();
 sg13g2_decap_4 FILLER_50_486 ();
 sg13g2_fill_1 FILLER_50_490 ();
 sg13g2_fill_1 FILLER_50_500 ();
 sg13g2_decap_8 FILLER_50_532 ();
 sg13g2_decap_8 FILLER_50_605 ();
 sg13g2_fill_1 FILLER_50_616 ();
 sg13g2_fill_2 FILLER_50_639 ();
 sg13g2_fill_1 FILLER_50_646 ();
 sg13g2_fill_1 FILLER_50_666 ();
 sg13g2_fill_2 FILLER_50_685 ();
 sg13g2_fill_1 FILLER_50_743 ();
 sg13g2_fill_2 FILLER_50_765 ();
 sg13g2_decap_8 FILLER_50_780 ();
 sg13g2_decap_8 FILLER_50_787 ();
 sg13g2_decap_8 FILLER_50_794 ();
 sg13g2_decap_8 FILLER_50_801 ();
 sg13g2_decap_8 FILLER_50_808 ();
 sg13g2_decap_8 FILLER_50_815 ();
 sg13g2_decap_8 FILLER_50_822 ();
 sg13g2_decap_8 FILLER_50_829 ();
 sg13g2_decap_8 FILLER_50_836 ();
 sg13g2_decap_8 FILLER_50_843 ();
 sg13g2_decap_8 FILLER_50_850 ();
 sg13g2_decap_4 FILLER_50_857 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_fill_2 FILLER_51_140 ();
 sg13g2_fill_2 FILLER_51_159 ();
 sg13g2_fill_2 FILLER_51_179 ();
 sg13g2_fill_1 FILLER_51_181 ();
 sg13g2_decap_8 FILLER_51_234 ();
 sg13g2_fill_2 FILLER_51_253 ();
 sg13g2_fill_2 FILLER_51_264 ();
 sg13g2_fill_1 FILLER_51_266 ();
 sg13g2_fill_2 FILLER_51_300 ();
 sg13g2_fill_2 FILLER_51_358 ();
 sg13g2_fill_1 FILLER_51_360 ();
 sg13g2_fill_2 FILLER_51_366 ();
 sg13g2_fill_1 FILLER_51_368 ();
 sg13g2_fill_1 FILLER_51_378 ();
 sg13g2_decap_4 FILLER_51_387 ();
 sg13g2_fill_2 FILLER_51_431 ();
 sg13g2_fill_1 FILLER_51_433 ();
 sg13g2_fill_2 FILLER_51_496 ();
 sg13g2_fill_1 FILLER_51_498 ();
 sg13g2_fill_2 FILLER_51_518 ();
 sg13g2_fill_1 FILLER_51_536 ();
 sg13g2_fill_2 FILLER_51_541 ();
 sg13g2_fill_1 FILLER_51_543 ();
 sg13g2_fill_1 FILLER_51_558 ();
 sg13g2_fill_1 FILLER_51_585 ();
 sg13g2_decap_8 FILLER_51_594 ();
 sg13g2_fill_1 FILLER_51_601 ();
 sg13g2_fill_2 FILLER_51_628 ();
 sg13g2_fill_1 FILLER_51_630 ();
 sg13g2_fill_2 FILLER_51_697 ();
 sg13g2_fill_1 FILLER_51_699 ();
 sg13g2_fill_2 FILLER_51_726 ();
 sg13g2_fill_1 FILLER_51_728 ();
 sg13g2_fill_2 FILLER_51_738 ();
 sg13g2_fill_1 FILLER_51_745 ();
 sg13g2_decap_8 FILLER_51_774 ();
 sg13g2_decap_8 FILLER_51_781 ();
 sg13g2_decap_8 FILLER_51_788 ();
 sg13g2_decap_8 FILLER_51_795 ();
 sg13g2_decap_8 FILLER_51_802 ();
 sg13g2_decap_8 FILLER_51_809 ();
 sg13g2_decap_8 FILLER_51_816 ();
 sg13g2_decap_8 FILLER_51_823 ();
 sg13g2_decap_8 FILLER_51_830 ();
 sg13g2_decap_8 FILLER_51_837 ();
 sg13g2_decap_8 FILLER_51_844 ();
 sg13g2_decap_8 FILLER_51_851 ();
 sg13g2_decap_4 FILLER_51_858 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_fill_2 FILLER_52_133 ();
 sg13g2_fill_1 FILLER_52_177 ();
 sg13g2_fill_1 FILLER_52_195 ();
 sg13g2_fill_1 FILLER_52_231 ();
 sg13g2_fill_2 FILLER_52_272 ();
 sg13g2_fill_2 FILLER_52_317 ();
 sg13g2_fill_2 FILLER_52_350 ();
 sg13g2_fill_2 FILLER_52_392 ();
 sg13g2_fill_2 FILLER_52_420 ();
 sg13g2_fill_2 FILLER_52_435 ();
 sg13g2_decap_8 FILLER_52_463 ();
 sg13g2_fill_2 FILLER_52_470 ();
 sg13g2_decap_4 FILLER_52_476 ();
 sg13g2_fill_2 FILLER_52_485 ();
 sg13g2_fill_1 FILLER_52_487 ();
 sg13g2_fill_1 FILLER_52_531 ();
 sg13g2_fill_2 FILLER_52_546 ();
 sg13g2_fill_1 FILLER_52_570 ();
 sg13g2_decap_8 FILLER_52_605 ();
 sg13g2_fill_2 FILLER_52_639 ();
 sg13g2_fill_1 FILLER_52_641 ();
 sg13g2_decap_8 FILLER_52_659 ();
 sg13g2_fill_2 FILLER_52_756 ();
 sg13g2_fill_1 FILLER_52_758 ();
 sg13g2_decap_8 FILLER_52_785 ();
 sg13g2_decap_8 FILLER_52_792 ();
 sg13g2_decap_8 FILLER_52_799 ();
 sg13g2_decap_8 FILLER_52_806 ();
 sg13g2_decap_8 FILLER_52_813 ();
 sg13g2_decap_8 FILLER_52_820 ();
 sg13g2_decap_8 FILLER_52_827 ();
 sg13g2_decap_8 FILLER_52_834 ();
 sg13g2_decap_8 FILLER_52_841 ();
 sg13g2_decap_8 FILLER_52_848 ();
 sg13g2_decap_8 FILLER_52_855 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_4 FILLER_53_126 ();
 sg13g2_fill_1 FILLER_53_130 ();
 sg13g2_fill_2 FILLER_53_157 ();
 sg13g2_fill_1 FILLER_53_159 ();
 sg13g2_fill_1 FILLER_53_170 ();
 sg13g2_fill_1 FILLER_53_207 ();
 sg13g2_fill_2 FILLER_53_226 ();
 sg13g2_fill_2 FILLER_53_252 ();
 sg13g2_fill_1 FILLER_53_283 ();
 sg13g2_fill_1 FILLER_53_289 ();
 sg13g2_fill_2 FILLER_53_299 ();
 sg13g2_decap_4 FILLER_53_325 ();
 sg13g2_fill_1 FILLER_53_329 ();
 sg13g2_fill_2 FILLER_53_347 ();
 sg13g2_fill_1 FILLER_53_349 ();
 sg13g2_fill_2 FILLER_53_358 ();
 sg13g2_fill_1 FILLER_53_360 ();
 sg13g2_fill_2 FILLER_53_366 ();
 sg13g2_fill_1 FILLER_53_373 ();
 sg13g2_decap_8 FILLER_53_388 ();
 sg13g2_decap_8 FILLER_53_395 ();
 sg13g2_fill_1 FILLER_53_402 ();
 sg13g2_decap_8 FILLER_53_425 ();
 sg13g2_decap_4 FILLER_53_462 ();
 sg13g2_fill_2 FILLER_53_466 ();
 sg13g2_fill_2 FILLER_53_498 ();
 sg13g2_fill_1 FILLER_53_500 ();
 sg13g2_decap_4 FILLER_53_510 ();
 sg13g2_fill_2 FILLER_53_529 ();
 sg13g2_fill_1 FILLER_53_531 ();
 sg13g2_fill_1 FILLER_53_563 ();
 sg13g2_decap_8 FILLER_53_587 ();
 sg13g2_decap_4 FILLER_53_594 ();
 sg13g2_fill_2 FILLER_53_598 ();
 sg13g2_fill_1 FILLER_53_606 ();
 sg13g2_decap_4 FILLER_53_638 ();
 sg13g2_fill_2 FILLER_53_677 ();
 sg13g2_fill_1 FILLER_53_679 ();
 sg13g2_decap_4 FILLER_53_689 ();
 sg13g2_decap_4 FILLER_53_697 ();
 sg13g2_fill_2 FILLER_53_714 ();
 sg13g2_fill_1 FILLER_53_737 ();
 sg13g2_fill_2 FILLER_53_765 ();
 sg13g2_fill_1 FILLER_53_767 ();
 sg13g2_decap_8 FILLER_53_777 ();
 sg13g2_decap_8 FILLER_53_784 ();
 sg13g2_decap_8 FILLER_53_791 ();
 sg13g2_decap_8 FILLER_53_798 ();
 sg13g2_decap_8 FILLER_53_805 ();
 sg13g2_decap_8 FILLER_53_812 ();
 sg13g2_decap_8 FILLER_53_819 ();
 sg13g2_decap_8 FILLER_53_826 ();
 sg13g2_decap_8 FILLER_53_833 ();
 sg13g2_decap_8 FILLER_53_840 ();
 sg13g2_decap_8 FILLER_53_847 ();
 sg13g2_decap_8 FILLER_53_854 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_fill_2 FILLER_54_133 ();
 sg13g2_fill_1 FILLER_54_135 ();
 sg13g2_fill_2 FILLER_54_214 ();
 sg13g2_fill_2 FILLER_54_290 ();
 sg13g2_decap_4 FILLER_54_305 ();
 sg13g2_decap_4 FILLER_54_339 ();
 sg13g2_fill_1 FILLER_54_343 ();
 sg13g2_fill_2 FILLER_54_363 ();
 sg13g2_fill_1 FILLER_54_365 ();
 sg13g2_fill_1 FILLER_54_448 ();
 sg13g2_fill_1 FILLER_54_469 ();
 sg13g2_fill_2 FILLER_54_533 ();
 sg13g2_fill_2 FILLER_54_548 ();
 sg13g2_fill_2 FILLER_54_559 ();
 sg13g2_fill_1 FILLER_54_561 ();
 sg13g2_decap_8 FILLER_54_608 ();
 sg13g2_fill_1 FILLER_54_615 ();
 sg13g2_fill_2 FILLER_54_639 ();
 sg13g2_decap_8 FILLER_54_645 ();
 sg13g2_fill_1 FILLER_54_652 ();
 sg13g2_decap_4 FILLER_54_657 ();
 sg13g2_fill_2 FILLER_54_661 ();
 sg13g2_fill_1 FILLER_54_708 ();
 sg13g2_fill_2 FILLER_54_748 ();
 sg13g2_fill_1 FILLER_54_750 ();
 sg13g2_decap_8 FILLER_54_777 ();
 sg13g2_decap_8 FILLER_54_784 ();
 sg13g2_decap_8 FILLER_54_791 ();
 sg13g2_decap_8 FILLER_54_798 ();
 sg13g2_decap_8 FILLER_54_805 ();
 sg13g2_decap_8 FILLER_54_812 ();
 sg13g2_decap_8 FILLER_54_819 ();
 sg13g2_decap_8 FILLER_54_826 ();
 sg13g2_decap_8 FILLER_54_833 ();
 sg13g2_decap_8 FILLER_54_840 ();
 sg13g2_decap_8 FILLER_54_847 ();
 sg13g2_decap_8 FILLER_54_854 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_4 FILLER_55_147 ();
 sg13g2_decap_4 FILLER_55_186 ();
 sg13g2_fill_2 FILLER_55_199 ();
 sg13g2_decap_8 FILLER_55_209 ();
 sg13g2_decap_8 FILLER_55_216 ();
 sg13g2_decap_4 FILLER_55_223 ();
 sg13g2_decap_4 FILLER_55_315 ();
 sg13g2_fill_2 FILLER_55_319 ();
 sg13g2_fill_1 FILLER_55_330 ();
 sg13g2_decap_4 FILLER_55_340 ();
 sg13g2_fill_2 FILLER_55_370 ();
 sg13g2_fill_1 FILLER_55_372 ();
 sg13g2_fill_2 FILLER_55_382 ();
 sg13g2_fill_1 FILLER_55_384 ();
 sg13g2_fill_2 FILLER_55_399 ();
 sg13g2_fill_2 FILLER_55_410 ();
 sg13g2_fill_1 FILLER_55_412 ();
 sg13g2_fill_1 FILLER_55_431 ();
 sg13g2_fill_2 FILLER_55_441 ();
 sg13g2_fill_2 FILLER_55_461 ();
 sg13g2_fill_2 FILLER_55_477 ();
 sg13g2_fill_2 FILLER_55_489 ();
 sg13g2_fill_1 FILLER_55_491 ();
 sg13g2_fill_2 FILLER_55_497 ();
 sg13g2_fill_1 FILLER_55_524 ();
 sg13g2_fill_1 FILLER_55_534 ();
 sg13g2_decap_8 FILLER_55_616 ();
 sg13g2_fill_2 FILLER_55_623 ();
 sg13g2_decap_8 FILLER_55_641 ();
 sg13g2_decap_4 FILLER_55_648 ();
 sg13g2_fill_1 FILLER_55_652 ();
 sg13g2_decap_8 FILLER_55_657 ();
 sg13g2_fill_1 FILLER_55_664 ();
 sg13g2_fill_1 FILLER_55_673 ();
 sg13g2_fill_2 FILLER_55_679 ();
 sg13g2_fill_1 FILLER_55_686 ();
 sg13g2_fill_2 FILLER_55_696 ();
 sg13g2_fill_1 FILLER_55_698 ();
 sg13g2_fill_1 FILLER_55_734 ();
 sg13g2_fill_1 FILLER_55_744 ();
 sg13g2_fill_2 FILLER_55_750 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_decap_8 FILLER_55_777 ();
 sg13g2_decap_8 FILLER_55_784 ();
 sg13g2_decap_8 FILLER_55_791 ();
 sg13g2_decap_8 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_805 ();
 sg13g2_decap_8 FILLER_55_812 ();
 sg13g2_decap_8 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_826 ();
 sg13g2_decap_8 FILLER_55_833 ();
 sg13g2_decap_8 FILLER_55_840 ();
 sg13g2_decap_8 FILLER_55_847 ();
 sg13g2_decap_8 FILLER_55_854 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_4 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_180 ();
 sg13g2_decap_8 FILLER_56_187 ();
 sg13g2_decap_8 FILLER_56_194 ();
 sg13g2_decap_8 FILLER_56_201 ();
 sg13g2_fill_2 FILLER_56_208 ();
 sg13g2_fill_1 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_222 ();
 sg13g2_decap_8 FILLER_56_229 ();
 sg13g2_fill_2 FILLER_56_263 ();
 sg13g2_decap_4 FILLER_56_290 ();
 sg13g2_fill_2 FILLER_56_294 ();
 sg13g2_fill_1 FILLER_56_309 ();
 sg13g2_fill_2 FILLER_56_350 ();
 sg13g2_fill_1 FILLER_56_352 ();
 sg13g2_fill_2 FILLER_56_438 ();
 sg13g2_fill_2 FILLER_56_466 ();
 sg13g2_fill_1 FILLER_56_511 ();
 sg13g2_fill_2 FILLER_56_524 ();
 sg13g2_fill_2 FILLER_56_556 ();
 sg13g2_fill_2 FILLER_56_582 ();
 sg13g2_fill_2 FILLER_56_598 ();
 sg13g2_fill_2 FILLER_56_639 ();
 sg13g2_fill_1 FILLER_56_641 ();
 sg13g2_fill_2 FILLER_56_690 ();
 sg13g2_decap_8 FILLER_56_773 ();
 sg13g2_decap_8 FILLER_56_780 ();
 sg13g2_decap_8 FILLER_56_787 ();
 sg13g2_decap_8 FILLER_56_794 ();
 sg13g2_decap_8 FILLER_56_801 ();
 sg13g2_decap_8 FILLER_56_808 ();
 sg13g2_decap_8 FILLER_56_815 ();
 sg13g2_decap_8 FILLER_56_822 ();
 sg13g2_decap_8 FILLER_56_829 ();
 sg13g2_decap_8 FILLER_56_836 ();
 sg13g2_decap_8 FILLER_56_843 ();
 sg13g2_decap_8 FILLER_56_850 ();
 sg13g2_decap_4 FILLER_56_857 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_decap_8 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_189 ();
 sg13g2_decap_8 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_231 ();
 sg13g2_decap_4 FILLER_57_238 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_fill_2 FILLER_57_272 ();
 sg13g2_fill_1 FILLER_57_284 ();
 sg13g2_fill_2 FILLER_57_337 ();
 sg13g2_fill_2 FILLER_57_375 ();
 sg13g2_fill_2 FILLER_57_381 ();
 sg13g2_fill_1 FILLER_57_383 ();
 sg13g2_fill_2 FILLER_57_388 ();
 sg13g2_decap_8 FILLER_57_404 ();
 sg13g2_fill_2 FILLER_57_411 ();
 sg13g2_fill_1 FILLER_57_434 ();
 sg13g2_fill_2 FILLER_57_440 ();
 sg13g2_fill_1 FILLER_57_442 ();
 sg13g2_fill_2 FILLER_57_460 ();
 sg13g2_fill_1 FILLER_57_462 ();
 sg13g2_fill_1 FILLER_57_489 ();
 sg13g2_fill_1 FILLER_57_546 ();
 sg13g2_fill_2 FILLER_57_639 ();
 sg13g2_fill_1 FILLER_57_641 ();
 sg13g2_decap_4 FILLER_57_659 ();
 sg13g2_fill_1 FILLER_57_677 ();
 sg13g2_fill_2 FILLER_57_691 ();
 sg13g2_fill_2 FILLER_57_698 ();
 sg13g2_fill_2 FILLER_57_705 ();
 sg13g2_fill_1 FILLER_57_707 ();
 sg13g2_fill_1 FILLER_57_744 ();
 sg13g2_fill_2 FILLER_57_759 ();
 sg13g2_fill_1 FILLER_57_761 ();
 sg13g2_decap_8 FILLER_57_779 ();
 sg13g2_decap_8 FILLER_57_786 ();
 sg13g2_decap_8 FILLER_57_793 ();
 sg13g2_decap_8 FILLER_57_800 ();
 sg13g2_decap_8 FILLER_57_807 ();
 sg13g2_decap_8 FILLER_57_814 ();
 sg13g2_decap_8 FILLER_57_821 ();
 sg13g2_decap_8 FILLER_57_828 ();
 sg13g2_decap_8 FILLER_57_835 ();
 sg13g2_decap_8 FILLER_57_842 ();
 sg13g2_decap_8 FILLER_57_849 ();
 sg13g2_decap_4 FILLER_57_856 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_210 ();
 sg13g2_decap_8 FILLER_58_217 ();
 sg13g2_decap_8 FILLER_58_224 ();
 sg13g2_fill_2 FILLER_58_279 ();
 sg13g2_fill_1 FILLER_58_300 ();
 sg13g2_fill_1 FILLER_58_306 ();
 sg13g2_fill_1 FILLER_58_311 ();
 sg13g2_fill_2 FILLER_58_385 ();
 sg13g2_decap_8 FILLER_58_407 ();
 sg13g2_fill_2 FILLER_58_427 ();
 sg13g2_fill_1 FILLER_58_523 ();
 sg13g2_fill_1 FILLER_58_549 ();
 sg13g2_decap_8 FILLER_58_555 ();
 sg13g2_fill_2 FILLER_58_562 ();
 sg13g2_decap_8 FILLER_58_605 ();
 sg13g2_decap_4 FILLER_58_677 ();
 sg13g2_fill_2 FILLER_58_693 ();
 sg13g2_fill_2 FILLER_58_704 ();
 sg13g2_fill_2 FILLER_58_711 ();
 sg13g2_fill_2 FILLER_58_727 ();
 sg13g2_fill_2 FILLER_58_751 ();
 sg13g2_fill_1 FILLER_58_753 ();
 sg13g2_fill_2 FILLER_58_759 ();
 sg13g2_fill_1 FILLER_58_761 ();
 sg13g2_decap_8 FILLER_58_780 ();
 sg13g2_decap_8 FILLER_58_787 ();
 sg13g2_decap_8 FILLER_58_794 ();
 sg13g2_decap_8 FILLER_58_801 ();
 sg13g2_decap_8 FILLER_58_808 ();
 sg13g2_decap_8 FILLER_58_815 ();
 sg13g2_decap_8 FILLER_58_822 ();
 sg13g2_decap_8 FILLER_58_829 ();
 sg13g2_decap_8 FILLER_58_836 ();
 sg13g2_decap_8 FILLER_58_843 ();
 sg13g2_decap_8 FILLER_58_850 ();
 sg13g2_decap_4 FILLER_58_857 ();
 sg13g2_fill_1 FILLER_58_861 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_fill_1 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_97 ();
 sg13g2_decap_8 FILLER_59_104 ();
 sg13g2_fill_2 FILLER_59_111 ();
 sg13g2_fill_2 FILLER_59_173 ();
 sg13g2_decap_8 FILLER_59_179 ();
 sg13g2_decap_4 FILLER_59_186 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_decap_8 FILLER_59_210 ();
 sg13g2_decap_8 FILLER_59_217 ();
 sg13g2_decap_8 FILLER_59_224 ();
 sg13g2_decap_8 FILLER_59_231 ();
 sg13g2_fill_2 FILLER_59_268 ();
 sg13g2_fill_2 FILLER_59_278 ();
 sg13g2_fill_1 FILLER_59_306 ();
 sg13g2_fill_2 FILLER_59_333 ();
 sg13g2_fill_2 FILLER_59_352 ();
 sg13g2_fill_2 FILLER_59_373 ();
 sg13g2_fill_2 FILLER_59_394 ();
 sg13g2_fill_1 FILLER_59_396 ();
 sg13g2_fill_2 FILLER_59_428 ();
 sg13g2_fill_2 FILLER_59_435 ();
 sg13g2_fill_2 FILLER_59_442 ();
 sg13g2_decap_4 FILLER_59_449 ();
 sg13g2_decap_4 FILLER_59_457 ();
 sg13g2_fill_1 FILLER_59_461 ();
 sg13g2_fill_2 FILLER_59_480 ();
 sg13g2_fill_2 FILLER_59_504 ();
 sg13g2_fill_1 FILLER_59_506 ();
 sg13g2_fill_2 FILLER_59_533 ();
 sg13g2_fill_1 FILLER_59_535 ();
 sg13g2_fill_2 FILLER_59_566 ();
 sg13g2_decap_4 FILLER_59_572 ();
 sg13g2_fill_1 FILLER_59_576 ();
 sg13g2_fill_1 FILLER_59_598 ();
 sg13g2_fill_1 FILLER_59_653 ();
 sg13g2_fill_1 FILLER_59_671 ();
 sg13g2_fill_1 FILLER_59_694 ();
 sg13g2_fill_2 FILLER_59_747 ();
 sg13g2_fill_1 FILLER_59_749 ();
 sg13g2_decap_8 FILLER_59_776 ();
 sg13g2_decap_8 FILLER_59_783 ();
 sg13g2_decap_8 FILLER_59_790 ();
 sg13g2_decap_8 FILLER_59_797 ();
 sg13g2_decap_8 FILLER_59_804 ();
 sg13g2_decap_8 FILLER_59_811 ();
 sg13g2_decap_8 FILLER_59_818 ();
 sg13g2_decap_8 FILLER_59_825 ();
 sg13g2_decap_8 FILLER_59_832 ();
 sg13g2_decap_8 FILLER_59_839 ();
 sg13g2_decap_8 FILLER_59_846 ();
 sg13g2_decap_8 FILLER_59_853 ();
 sg13g2_fill_2 FILLER_59_860 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_4 FILLER_60_77 ();
 sg13g2_fill_2 FILLER_60_137 ();
 sg13g2_decap_8 FILLER_60_210 ();
 sg13g2_decap_8 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_238 ();
 sg13g2_decap_4 FILLER_60_245 ();
 sg13g2_fill_1 FILLER_60_249 ();
 sg13g2_fill_2 FILLER_60_295 ();
 sg13g2_fill_2 FILLER_60_311 ();
 sg13g2_fill_1 FILLER_60_313 ();
 sg13g2_fill_2 FILLER_60_336 ();
 sg13g2_fill_2 FILLER_60_342 ();
 sg13g2_fill_1 FILLER_60_344 ();
 sg13g2_decap_4 FILLER_60_407 ();
 sg13g2_fill_2 FILLER_60_411 ();
 sg13g2_decap_8 FILLER_60_417 ();
 sg13g2_fill_2 FILLER_60_424 ();
 sg13g2_fill_1 FILLER_60_426 ();
 sg13g2_fill_2 FILLER_60_431 ();
 sg13g2_fill_2 FILLER_60_442 ();
 sg13g2_fill_1 FILLER_60_453 ();
 sg13g2_fill_1 FILLER_60_507 ();
 sg13g2_decap_4 FILLER_60_542 ();
 sg13g2_fill_1 FILLER_60_546 ();
 sg13g2_fill_2 FILLER_60_551 ();
 sg13g2_fill_2 FILLER_60_571 ();
 sg13g2_fill_2 FILLER_60_594 ();
 sg13g2_decap_8 FILLER_60_601 ();
 sg13g2_fill_2 FILLER_60_608 ();
 sg13g2_decap_4 FILLER_60_614 ();
 sg13g2_decap_4 FILLER_60_670 ();
 sg13g2_fill_2 FILLER_60_694 ();
 sg13g2_fill_2 FILLER_60_710 ();
 sg13g2_fill_1 FILLER_60_721 ();
 sg13g2_fill_2 FILLER_60_735 ();
 sg13g2_fill_1 FILLER_60_750 ();
 sg13g2_decap_8 FILLER_60_769 ();
 sg13g2_decap_8 FILLER_60_776 ();
 sg13g2_decap_8 FILLER_60_783 ();
 sg13g2_decap_8 FILLER_60_790 ();
 sg13g2_decap_8 FILLER_60_797 ();
 sg13g2_decap_8 FILLER_60_804 ();
 sg13g2_decap_8 FILLER_60_811 ();
 sg13g2_decap_8 FILLER_60_818 ();
 sg13g2_decap_8 FILLER_60_825 ();
 sg13g2_decap_8 FILLER_60_832 ();
 sg13g2_decap_8 FILLER_60_839 ();
 sg13g2_decap_8 FILLER_60_846 ();
 sg13g2_decap_8 FILLER_60_853 ();
 sg13g2_fill_2 FILLER_60_860 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_4 FILLER_61_56 ();
 sg13g2_fill_1 FILLER_61_60 ();
 sg13g2_fill_1 FILLER_61_87 ();
 sg13g2_fill_2 FILLER_61_105 ();
 sg13g2_fill_1 FILLER_61_107 ();
 sg13g2_fill_2 FILLER_61_117 ();
 sg13g2_fill_1 FILLER_61_119 ();
 sg13g2_fill_2 FILLER_61_156 ();
 sg13g2_fill_2 FILLER_61_164 ();
 sg13g2_fill_1 FILLER_61_193 ();
 sg13g2_decap_8 FILLER_61_220 ();
 sg13g2_decap_8 FILLER_61_227 ();
 sg13g2_decap_4 FILLER_61_234 ();
 sg13g2_fill_2 FILLER_61_238 ();
 sg13g2_fill_1 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_fill_2 FILLER_61_350 ();
 sg13g2_fill_2 FILLER_61_357 ();
 sg13g2_fill_2 FILLER_61_394 ();
 sg13g2_decap_8 FILLER_61_409 ();
 sg13g2_fill_1 FILLER_61_416 ();
 sg13g2_fill_1 FILLER_61_464 ();
 sg13g2_decap_4 FILLER_61_469 ();
 sg13g2_fill_1 FILLER_61_517 ();
 sg13g2_fill_2 FILLER_61_612 ();
 sg13g2_fill_1 FILLER_61_614 ();
 sg13g2_decap_4 FILLER_61_619 ();
 sg13g2_fill_1 FILLER_61_623 ();
 sg13g2_fill_1 FILLER_61_628 ();
 sg13g2_decap_4 FILLER_61_633 ();
 sg13g2_fill_1 FILLER_61_637 ();
 sg13g2_fill_2 FILLER_61_659 ();
 sg13g2_fill_2 FILLER_61_698 ();
 sg13g2_fill_1 FILLER_61_700 ();
 sg13g2_fill_1 FILLER_61_732 ();
 sg13g2_fill_2 FILLER_61_746 ();
 sg13g2_decap_8 FILLER_61_774 ();
 sg13g2_decap_8 FILLER_61_781 ();
 sg13g2_decap_8 FILLER_61_788 ();
 sg13g2_decap_8 FILLER_61_795 ();
 sg13g2_decap_8 FILLER_61_802 ();
 sg13g2_decap_8 FILLER_61_809 ();
 sg13g2_decap_8 FILLER_61_816 ();
 sg13g2_decap_8 FILLER_61_823 ();
 sg13g2_decap_8 FILLER_61_830 ();
 sg13g2_decap_8 FILLER_61_837 ();
 sg13g2_decap_8 FILLER_61_844 ();
 sg13g2_decap_8 FILLER_61_851 ();
 sg13g2_decap_4 FILLER_61_858 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_4 FILLER_62_56 ();
 sg13g2_fill_2 FILLER_62_60 ();
 sg13g2_fill_2 FILLER_62_87 ();
 sg13g2_fill_2 FILLER_62_97 ();
 sg13g2_fill_1 FILLER_62_99 ();
 sg13g2_fill_1 FILLER_62_109 ();
 sg13g2_fill_1 FILLER_62_133 ();
 sg13g2_fill_1 FILLER_62_160 ();
 sg13g2_fill_1 FILLER_62_169 ();
 sg13g2_fill_2 FILLER_62_218 ();
 sg13g2_fill_1 FILLER_62_220 ();
 sg13g2_fill_1 FILLER_62_239 ();
 sg13g2_fill_1 FILLER_62_331 ();
 sg13g2_decap_8 FILLER_62_340 ();
 sg13g2_fill_2 FILLER_62_408 ();
 sg13g2_fill_2 FILLER_62_436 ();
 sg13g2_fill_1 FILLER_62_438 ();
 sg13g2_fill_2 FILLER_62_462 ();
 sg13g2_fill_2 FILLER_62_471 ();
 sg13g2_fill_1 FILLER_62_473 ();
 sg13g2_fill_2 FILLER_62_479 ();
 sg13g2_fill_1 FILLER_62_517 ();
 sg13g2_fill_2 FILLER_62_522 ();
 sg13g2_fill_2 FILLER_62_534 ();
 sg13g2_fill_1 FILLER_62_536 ();
 sg13g2_fill_1 FILLER_62_551 ();
 sg13g2_fill_2 FILLER_62_561 ();
 sg13g2_fill_2 FILLER_62_577 ();
 sg13g2_fill_2 FILLER_62_588 ();
 sg13g2_fill_2 FILLER_62_643 ();
 sg13g2_fill_1 FILLER_62_645 ();
 sg13g2_fill_2 FILLER_62_651 ();
 sg13g2_decap_8 FILLER_62_772 ();
 sg13g2_decap_8 FILLER_62_779 ();
 sg13g2_decap_8 FILLER_62_786 ();
 sg13g2_decap_8 FILLER_62_793 ();
 sg13g2_decap_8 FILLER_62_800 ();
 sg13g2_decap_8 FILLER_62_807 ();
 sg13g2_decap_8 FILLER_62_814 ();
 sg13g2_decap_8 FILLER_62_821 ();
 sg13g2_decap_8 FILLER_62_828 ();
 sg13g2_decap_8 FILLER_62_835 ();
 sg13g2_decap_8 FILLER_62_842 ();
 sg13g2_decap_8 FILLER_62_849 ();
 sg13g2_decap_4 FILLER_62_856 ();
 sg13g2_fill_2 FILLER_62_860 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_fill_2 FILLER_63_42 ();
 sg13g2_fill_1 FILLER_63_44 ();
 sg13g2_decap_4 FILLER_63_49 ();
 sg13g2_fill_1 FILLER_63_53 ();
 sg13g2_fill_1 FILLER_63_149 ();
 sg13g2_fill_2 FILLER_63_155 ();
 sg13g2_fill_1 FILLER_63_168 ();
 sg13g2_fill_2 FILLER_63_195 ();
 sg13g2_fill_1 FILLER_63_197 ();
 sg13g2_fill_1 FILLER_63_224 ();
 sg13g2_fill_1 FILLER_63_251 ();
 sg13g2_fill_2 FILLER_63_293 ();
 sg13g2_fill_1 FILLER_63_295 ();
 sg13g2_fill_1 FILLER_63_306 ();
 sg13g2_decap_4 FILLER_63_335 ();
 sg13g2_decap_4 FILLER_63_343 ();
 sg13g2_fill_1 FILLER_63_347 ();
 sg13g2_fill_1 FILLER_63_362 ();
 sg13g2_fill_1 FILLER_63_377 ();
 sg13g2_decap_8 FILLER_63_397 ();
 sg13g2_fill_1 FILLER_63_404 ();
 sg13g2_fill_1 FILLER_63_410 ();
 sg13g2_decap_8 FILLER_63_429 ();
 sg13g2_fill_2 FILLER_63_462 ();
 sg13g2_fill_2 FILLER_63_485 ();
 sg13g2_decap_4 FILLER_63_513 ();
 sg13g2_fill_2 FILLER_63_517 ();
 sg13g2_fill_2 FILLER_63_545 ();
 sg13g2_fill_2 FILLER_63_573 ();
 sg13g2_fill_1 FILLER_63_575 ();
 sg13g2_fill_2 FILLER_63_636 ();
 sg13g2_fill_1 FILLER_63_638 ();
 sg13g2_decap_4 FILLER_63_696 ();
 sg13g2_fill_2 FILLER_63_700 ();
 sg13g2_fill_2 FILLER_63_733 ();
 sg13g2_fill_1 FILLER_63_742 ();
 sg13g2_decap_4 FILLER_63_751 ();
 sg13g2_decap_8 FILLER_63_781 ();
 sg13g2_decap_8 FILLER_63_788 ();
 sg13g2_decap_8 FILLER_63_795 ();
 sg13g2_decap_8 FILLER_63_802 ();
 sg13g2_decap_8 FILLER_63_809 ();
 sg13g2_decap_8 FILLER_63_816 ();
 sg13g2_decap_8 FILLER_63_823 ();
 sg13g2_decap_8 FILLER_63_830 ();
 sg13g2_decap_8 FILLER_63_837 ();
 sg13g2_decap_8 FILLER_63_844 ();
 sg13g2_decap_8 FILLER_63_851 ();
 sg13g2_decap_4 FILLER_63_858 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_14 ();
 sg13g2_fill_2 FILLER_64_18 ();
 sg13g2_decap_8 FILLER_64_24 ();
 sg13g2_fill_2 FILLER_64_31 ();
 sg13g2_fill_2 FILLER_64_91 ();
 sg13g2_fill_1 FILLER_64_107 ();
 sg13g2_fill_1 FILLER_64_176 ();
 sg13g2_fill_2 FILLER_64_195 ();
 sg13g2_fill_1 FILLER_64_197 ();
 sg13g2_fill_2 FILLER_64_206 ();
 sg13g2_fill_1 FILLER_64_208 ();
 sg13g2_decap_8 FILLER_64_213 ();
 sg13g2_fill_1 FILLER_64_220 ();
 sg13g2_fill_2 FILLER_64_246 ();
 sg13g2_fill_1 FILLER_64_248 ();
 sg13g2_fill_2 FILLER_64_395 ();
 sg13g2_decap_8 FILLER_64_428 ();
 sg13g2_decap_4 FILLER_64_435 ();
 sg13g2_fill_2 FILLER_64_448 ();
 sg13g2_fill_1 FILLER_64_459 ();
 sg13g2_fill_1 FILLER_64_524 ();
 sg13g2_fill_1 FILLER_64_548 ();
 sg13g2_fill_1 FILLER_64_598 ();
 sg13g2_fill_2 FILLER_64_636 ();
 sg13g2_fill_1 FILLER_64_638 ();
 sg13g2_decap_8 FILLER_64_658 ();
 sg13g2_decap_8 FILLER_64_665 ();
 sg13g2_fill_2 FILLER_64_672 ();
 sg13g2_fill_2 FILLER_64_705 ();
 sg13g2_fill_1 FILLER_64_715 ();
 sg13g2_fill_2 FILLER_64_720 ();
 sg13g2_fill_1 FILLER_64_722 ();
 sg13g2_fill_2 FILLER_64_736 ();
 sg13g2_fill_1 FILLER_64_743 ();
 sg13g2_decap_8 FILLER_64_776 ();
 sg13g2_decap_8 FILLER_64_783 ();
 sg13g2_decap_8 FILLER_64_790 ();
 sg13g2_decap_8 FILLER_64_797 ();
 sg13g2_decap_8 FILLER_64_804 ();
 sg13g2_decap_8 FILLER_64_811 ();
 sg13g2_decap_8 FILLER_64_818 ();
 sg13g2_decap_8 FILLER_64_825 ();
 sg13g2_decap_8 FILLER_64_832 ();
 sg13g2_decap_8 FILLER_64_839 ();
 sg13g2_decap_8 FILLER_64_846 ();
 sg13g2_decap_8 FILLER_64_853 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_40 ();
 sg13g2_fill_2 FILLER_65_72 ();
 sg13g2_fill_1 FILLER_65_74 ();
 sg13g2_fill_1 FILLER_65_88 ();
 sg13g2_fill_1 FILLER_65_106 ();
 sg13g2_fill_2 FILLER_65_116 ();
 sg13g2_fill_1 FILLER_65_118 ();
 sg13g2_decap_4 FILLER_65_212 ();
 sg13g2_fill_1 FILLER_65_216 ();
 sg13g2_fill_2 FILLER_65_230 ();
 sg13g2_decap_8 FILLER_65_236 ();
 sg13g2_fill_2 FILLER_65_243 ();
 sg13g2_fill_1 FILLER_65_245 ();
 sg13g2_fill_2 FILLER_65_278 ();
 sg13g2_fill_2 FILLER_65_322 ();
 sg13g2_decap_8 FILLER_65_333 ();
 sg13g2_decap_8 FILLER_65_340 ();
 sg13g2_decap_4 FILLER_65_347 ();
 sg13g2_fill_1 FILLER_65_351 ();
 sg13g2_fill_1 FILLER_65_362 ();
 sg13g2_fill_2 FILLER_65_398 ();
 sg13g2_fill_1 FILLER_65_411 ();
 sg13g2_fill_1 FILLER_65_416 ();
 sg13g2_fill_1 FILLER_65_458 ();
 sg13g2_fill_2 FILLER_65_472 ();
 sg13g2_fill_1 FILLER_65_474 ();
 sg13g2_fill_2 FILLER_65_501 ();
 sg13g2_fill_1 FILLER_65_503 ();
 sg13g2_fill_1 FILLER_65_508 ();
 sg13g2_fill_2 FILLER_65_544 ();
 sg13g2_fill_1 FILLER_65_590 ();
 sg13g2_fill_2 FILLER_65_596 ();
 sg13g2_fill_1 FILLER_65_615 ();
 sg13g2_fill_2 FILLER_65_625 ();
 sg13g2_fill_1 FILLER_65_627 ();
 sg13g2_fill_1 FILLER_65_641 ();
 sg13g2_decap_8 FILLER_65_668 ();
 sg13g2_fill_2 FILLER_65_675 ();
 sg13g2_fill_2 FILLER_65_694 ();
 sg13g2_fill_2 FILLER_65_705 ();
 sg13g2_fill_2 FILLER_65_733 ();
 sg13g2_decap_4 FILLER_65_753 ();
 sg13g2_decap_8 FILLER_65_774 ();
 sg13g2_decap_8 FILLER_65_781 ();
 sg13g2_decap_8 FILLER_65_788 ();
 sg13g2_decap_8 FILLER_65_795 ();
 sg13g2_decap_8 FILLER_65_802 ();
 sg13g2_decap_8 FILLER_65_809 ();
 sg13g2_decap_8 FILLER_65_816 ();
 sg13g2_decap_8 FILLER_65_823 ();
 sg13g2_decap_8 FILLER_65_830 ();
 sg13g2_decap_8 FILLER_65_837 ();
 sg13g2_decap_8 FILLER_65_844 ();
 sg13g2_decap_8 FILLER_65_851 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_fill_2 FILLER_66_21 ();
 sg13g2_fill_1 FILLER_66_23 ();
 sg13g2_fill_2 FILLER_66_131 ();
 sg13g2_fill_2 FILLER_66_153 ();
 sg13g2_fill_2 FILLER_66_187 ();
 sg13g2_decap_4 FILLER_66_198 ();
 sg13g2_fill_2 FILLER_66_202 ();
 sg13g2_fill_1 FILLER_66_212 ();
 sg13g2_fill_2 FILLER_66_247 ();
 sg13g2_fill_2 FILLER_66_284 ();
 sg13g2_fill_1 FILLER_66_286 ();
 sg13g2_fill_2 FILLER_66_356 ();
 sg13g2_fill_1 FILLER_66_358 ();
 sg13g2_fill_1 FILLER_66_394 ();
 sg13g2_fill_2 FILLER_66_404 ();
 sg13g2_fill_1 FILLER_66_406 ();
 sg13g2_decap_4 FILLER_66_412 ();
 sg13g2_fill_1 FILLER_66_420 ();
 sg13g2_fill_1 FILLER_66_430 ();
 sg13g2_decap_8 FILLER_66_440 ();
 sg13g2_fill_2 FILLER_66_447 ();
 sg13g2_fill_1 FILLER_66_449 ();
 sg13g2_fill_2 FILLER_66_477 ();
 sg13g2_fill_1 FILLER_66_479 ();
 sg13g2_fill_1 FILLER_66_503 ();
 sg13g2_fill_2 FILLER_66_555 ();
 sg13g2_fill_2 FILLER_66_621 ();
 sg13g2_fill_1 FILLER_66_623 ();
 sg13g2_fill_1 FILLER_66_662 ();
 sg13g2_fill_2 FILLER_66_681 ();
 sg13g2_fill_2 FILLER_66_692 ();
 sg13g2_fill_1 FILLER_66_694 ();
 sg13g2_fill_2 FILLER_66_700 ();
 sg13g2_fill_1 FILLER_66_707 ();
 sg13g2_fill_2 FILLER_66_715 ();
 sg13g2_fill_1 FILLER_66_735 ();
 sg13g2_fill_2 FILLER_66_745 ();
 sg13g2_fill_1 FILLER_66_752 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_decap_8 FILLER_66_786 ();
 sg13g2_decap_8 FILLER_66_793 ();
 sg13g2_decap_8 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_807 ();
 sg13g2_decap_8 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_4 FILLER_66_856 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_69 ();
 sg13g2_fill_2 FILLER_67_107 ();
 sg13g2_fill_1 FILLER_67_109 ();
 sg13g2_fill_2 FILLER_67_118 ();
 sg13g2_fill_1 FILLER_67_120 ();
 sg13g2_fill_2 FILLER_67_147 ();
 sg13g2_fill_1 FILLER_67_149 ();
 sg13g2_fill_2 FILLER_67_167 ();
 sg13g2_fill_1 FILLER_67_169 ();
 sg13g2_fill_2 FILLER_67_194 ();
 sg13g2_fill_2 FILLER_67_212 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_fill_2 FILLER_67_252 ();
 sg13g2_fill_1 FILLER_67_280 ();
 sg13g2_fill_1 FILLER_67_286 ();
 sg13g2_fill_2 FILLER_67_296 ();
 sg13g2_decap_8 FILLER_67_302 ();
 sg13g2_decap_4 FILLER_67_309 ();
 sg13g2_fill_1 FILLER_67_326 ();
 sg13g2_fill_1 FILLER_67_336 ();
 sg13g2_fill_2 FILLER_67_350 ();
 sg13g2_fill_1 FILLER_67_430 ();
 sg13g2_fill_1 FILLER_67_457 ();
 sg13g2_fill_2 FILLER_67_485 ();
 sg13g2_fill_1 FILLER_67_487 ();
 sg13g2_fill_2 FILLER_67_540 ();
 sg13g2_fill_1 FILLER_67_556 ();
 sg13g2_fill_1 FILLER_67_565 ();
 sg13g2_fill_2 FILLER_67_583 ();
 sg13g2_fill_1 FILLER_67_585 ();
 sg13g2_fill_2 FILLER_67_611 ();
 sg13g2_fill_2 FILLER_67_649 ();
 sg13g2_fill_1 FILLER_67_730 ();
 sg13g2_decap_8 FILLER_67_765 ();
 sg13g2_decap_8 FILLER_67_772 ();
 sg13g2_decap_8 FILLER_67_779 ();
 sg13g2_decap_8 FILLER_67_786 ();
 sg13g2_decap_8 FILLER_67_793 ();
 sg13g2_decap_8 FILLER_67_800 ();
 sg13g2_decap_8 FILLER_67_807 ();
 sg13g2_decap_8 FILLER_67_814 ();
 sg13g2_decap_8 FILLER_67_821 ();
 sg13g2_decap_8 FILLER_67_828 ();
 sg13g2_decap_8 FILLER_67_835 ();
 sg13g2_decap_8 FILLER_67_842 ();
 sg13g2_decap_8 FILLER_67_849 ();
 sg13g2_decap_4 FILLER_67_856 ();
 sg13g2_fill_2 FILLER_67_860 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_fill_2 FILLER_68_21 ();
 sg13g2_fill_1 FILLER_68_23 ();
 sg13g2_fill_1 FILLER_68_90 ();
 sg13g2_decap_8 FILLER_68_109 ();
 sg13g2_fill_2 FILLER_68_116 ();
 sg13g2_fill_1 FILLER_68_118 ();
 sg13g2_fill_2 FILLER_68_149 ();
 sg13g2_decap_4 FILLER_68_159 ();
 sg13g2_fill_1 FILLER_68_163 ();
 sg13g2_decap_8 FILLER_68_169 ();
 sg13g2_decap_4 FILLER_68_176 ();
 sg13g2_fill_2 FILLER_68_180 ();
 sg13g2_fill_2 FILLER_68_208 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_fill_1 FILLER_68_219 ();
 sg13g2_fill_1 FILLER_68_255 ();
 sg13g2_decap_8 FILLER_68_296 ();
 sg13g2_decap_8 FILLER_68_303 ();
 sg13g2_decap_4 FILLER_68_310 ();
 sg13g2_fill_2 FILLER_68_339 ();
 sg13g2_fill_1 FILLER_68_346 ();
 sg13g2_fill_2 FILLER_68_357 ();
 sg13g2_fill_2 FILLER_68_373 ();
 sg13g2_fill_1 FILLER_68_375 ();
 sg13g2_fill_2 FILLER_68_385 ();
 sg13g2_fill_1 FILLER_68_387 ();
 sg13g2_decap_4 FILLER_68_409 ();
 sg13g2_fill_2 FILLER_68_464 ();
 sg13g2_fill_1 FILLER_68_466 ();
 sg13g2_fill_2 FILLER_68_477 ();
 sg13g2_decap_8 FILLER_68_510 ();
 sg13g2_decap_4 FILLER_68_517 ();
 sg13g2_fill_2 FILLER_68_521 ();
 sg13g2_fill_2 FILLER_68_546 ();
 sg13g2_fill_1 FILLER_68_548 ();
 sg13g2_fill_2 FILLER_68_575 ();
 sg13g2_fill_2 FILLER_68_627 ();
 sg13g2_fill_1 FILLER_68_629 ();
 sg13g2_fill_1 FILLER_68_635 ();
 sg13g2_decap_4 FILLER_68_662 ();
 sg13g2_decap_4 FILLER_68_671 ();
 sg13g2_fill_1 FILLER_68_675 ();
 sg13g2_decap_8 FILLER_68_684 ();
 sg13g2_fill_1 FILLER_68_691 ();
 sg13g2_fill_2 FILLER_68_713 ();
 sg13g2_fill_1 FILLER_68_715 ();
 sg13g2_fill_2 FILLER_68_730 ();
 sg13g2_fill_1 FILLER_68_732 ();
 sg13g2_decap_8 FILLER_68_768 ();
 sg13g2_decap_8 FILLER_68_775 ();
 sg13g2_decap_8 FILLER_68_782 ();
 sg13g2_decap_8 FILLER_68_789 ();
 sg13g2_decap_8 FILLER_68_796 ();
 sg13g2_decap_8 FILLER_68_803 ();
 sg13g2_decap_8 FILLER_68_810 ();
 sg13g2_decap_8 FILLER_68_817 ();
 sg13g2_decap_8 FILLER_68_824 ();
 sg13g2_decap_8 FILLER_68_831 ();
 sg13g2_decap_8 FILLER_68_838 ();
 sg13g2_decap_8 FILLER_68_845 ();
 sg13g2_decap_8 FILLER_68_852 ();
 sg13g2_fill_2 FILLER_68_859 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_11 ();
 sg13g2_fill_1 FILLER_69_51 ();
 sg13g2_fill_2 FILLER_69_83 ();
 sg13g2_fill_1 FILLER_69_85 ();
 sg13g2_decap_4 FILLER_69_94 ();
 sg13g2_fill_2 FILLER_69_106 ();
 sg13g2_fill_1 FILLER_69_108 ();
 sg13g2_fill_1 FILLER_69_113 ();
 sg13g2_fill_2 FILLER_69_139 ();
 sg13g2_fill_2 FILLER_69_159 ();
 sg13g2_decap_8 FILLER_69_179 ();
 sg13g2_fill_1 FILLER_69_186 ();
 sg13g2_decap_8 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_205 ();
 sg13g2_fill_2 FILLER_69_210 ();
 sg13g2_fill_1 FILLER_69_221 ();
 sg13g2_fill_1 FILLER_69_239 ();
 sg13g2_fill_2 FILLER_69_266 ();
 sg13g2_fill_2 FILLER_69_311 ();
 sg13g2_fill_1 FILLER_69_313 ();
 sg13g2_fill_2 FILLER_69_357 ();
 sg13g2_fill_1 FILLER_69_404 ();
 sg13g2_fill_2 FILLER_69_474 ();
 sg13g2_fill_1 FILLER_69_528 ();
 sg13g2_fill_2 FILLER_69_546 ();
 sg13g2_fill_1 FILLER_69_548 ();
 sg13g2_decap_4 FILLER_69_587 ();
 sg13g2_fill_2 FILLER_69_600 ();
 sg13g2_fill_1 FILLER_69_622 ();
 sg13g2_decap_8 FILLER_69_637 ();
 sg13g2_fill_2 FILLER_69_644 ();
 sg13g2_fill_1 FILLER_69_646 ();
 sg13g2_fill_1 FILLER_69_651 ();
 sg13g2_fill_2 FILLER_69_657 ();
 sg13g2_fill_2 FILLER_69_664 ();
 sg13g2_decap_4 FILLER_69_709 ();
 sg13g2_fill_2 FILLER_69_754 ();
 sg13g2_fill_1 FILLER_69_756 ();
 sg13g2_decap_8 FILLER_69_766 ();
 sg13g2_decap_8 FILLER_69_773 ();
 sg13g2_decap_8 FILLER_69_780 ();
 sg13g2_decap_8 FILLER_69_787 ();
 sg13g2_decap_8 FILLER_69_794 ();
 sg13g2_decap_8 FILLER_69_801 ();
 sg13g2_decap_8 FILLER_69_808 ();
 sg13g2_decap_8 FILLER_69_815 ();
 sg13g2_decap_8 FILLER_69_822 ();
 sg13g2_decap_8 FILLER_69_829 ();
 sg13g2_decap_8 FILLER_69_836 ();
 sg13g2_decap_8 FILLER_69_843 ();
 sg13g2_decap_8 FILLER_69_850 ();
 sg13g2_decap_4 FILLER_69_857 ();
 sg13g2_fill_1 FILLER_69_861 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_fill_2 FILLER_70_14 ();
 sg13g2_fill_1 FILLER_70_16 ();
 sg13g2_fill_2 FILLER_70_81 ();
 sg13g2_decap_8 FILLER_70_129 ();
 sg13g2_fill_2 FILLER_70_136 ();
 sg13g2_fill_2 FILLER_70_143 ();
 sg13g2_fill_1 FILLER_70_145 ();
 sg13g2_fill_2 FILLER_70_182 ();
 sg13g2_fill_1 FILLER_70_184 ();
 sg13g2_fill_2 FILLER_70_210 ();
 sg13g2_fill_2 FILLER_70_224 ();
 sg13g2_fill_1 FILLER_70_226 ();
 sg13g2_fill_1 FILLER_70_232 ();
 sg13g2_fill_2 FILLER_70_274 ();
 sg13g2_decap_4 FILLER_70_330 ();
 sg13g2_fill_2 FILLER_70_334 ();
 sg13g2_fill_1 FILLER_70_368 ();
 sg13g2_fill_2 FILLER_70_396 ();
 sg13g2_fill_1 FILLER_70_398 ();
 sg13g2_fill_2 FILLER_70_425 ();
 sg13g2_decap_8 FILLER_70_446 ();
 sg13g2_decap_8 FILLER_70_488 ();
 sg13g2_decap_4 FILLER_70_495 ();
 sg13g2_decap_4 FILLER_70_502 ();
 sg13g2_fill_1 FILLER_70_506 ();
 sg13g2_fill_1 FILLER_70_516 ();
 sg13g2_fill_2 FILLER_70_561 ();
 sg13g2_decap_4 FILLER_70_615 ();
 sg13g2_decap_4 FILLER_70_688 ();
 sg13g2_fill_2 FILLER_70_692 ();
 sg13g2_fill_1 FILLER_70_704 ();
 sg13g2_fill_1 FILLER_70_710 ();
 sg13g2_fill_1 FILLER_70_720 ();
 sg13g2_decap_8 FILLER_70_730 ();
 sg13g2_fill_2 FILLER_70_737 ();
 sg13g2_decap_8 FILLER_70_744 ();
 sg13g2_fill_2 FILLER_70_751 ();
 sg13g2_decap_8 FILLER_70_757 ();
 sg13g2_decap_8 FILLER_70_764 ();
 sg13g2_decap_8 FILLER_70_771 ();
 sg13g2_decap_8 FILLER_70_778 ();
 sg13g2_decap_8 FILLER_70_785 ();
 sg13g2_decap_8 FILLER_70_792 ();
 sg13g2_decap_8 FILLER_70_799 ();
 sg13g2_decap_8 FILLER_70_806 ();
 sg13g2_decap_8 FILLER_70_813 ();
 sg13g2_decap_8 FILLER_70_820 ();
 sg13g2_decap_8 FILLER_70_827 ();
 sg13g2_decap_8 FILLER_70_834 ();
 sg13g2_decap_8 FILLER_70_841 ();
 sg13g2_decap_8 FILLER_70_848 ();
 sg13g2_decap_8 FILLER_70_855 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_fill_2 FILLER_71_21 ();
 sg13g2_decap_4 FILLER_71_86 ();
 sg13g2_fill_2 FILLER_71_90 ();
 sg13g2_fill_2 FILLER_71_100 ();
 sg13g2_fill_1 FILLER_71_102 ();
 sg13g2_fill_1 FILLER_71_111 ();
 sg13g2_fill_2 FILLER_71_121 ();
 sg13g2_fill_2 FILLER_71_127 ();
 sg13g2_fill_1 FILLER_71_129 ();
 sg13g2_fill_2 FILLER_71_135 ();
 sg13g2_fill_1 FILLER_71_137 ();
 sg13g2_fill_1 FILLER_71_146 ();
 sg13g2_decap_4 FILLER_71_152 ();
 sg13g2_fill_1 FILLER_71_156 ();
 sg13g2_decap_4 FILLER_71_161 ();
 sg13g2_decap_4 FILLER_71_184 ();
 sg13g2_fill_2 FILLER_71_188 ();
 sg13g2_fill_1 FILLER_71_214 ();
 sg13g2_fill_2 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_242 ();
 sg13g2_fill_1 FILLER_71_249 ();
 sg13g2_decap_4 FILLER_71_291 ();
 sg13g2_fill_1 FILLER_71_295 ();
 sg13g2_fill_2 FILLER_71_304 ();
 sg13g2_decap_4 FILLER_71_311 ();
 sg13g2_fill_2 FILLER_71_319 ();
 sg13g2_fill_2 FILLER_71_343 ();
 sg13g2_fill_1 FILLER_71_345 ();
 sg13g2_fill_2 FILLER_71_382 ();
 sg13g2_decap_8 FILLER_71_410 ();
 sg13g2_decap_8 FILLER_71_417 ();
 sg13g2_fill_1 FILLER_71_424 ();
 sg13g2_decap_8 FILLER_71_430 ();
 sg13g2_decap_8 FILLER_71_437 ();
 sg13g2_decap_8 FILLER_71_444 ();
 sg13g2_decap_8 FILLER_71_451 ();
 sg13g2_decap_4 FILLER_71_458 ();
 sg13g2_fill_2 FILLER_71_462 ();
 sg13g2_decap_8 FILLER_71_468 ();
 sg13g2_decap_8 FILLER_71_475 ();
 sg13g2_fill_2 FILLER_71_482 ();
 sg13g2_fill_2 FILLER_71_510 ();
 sg13g2_fill_1 FILLER_71_562 ();
 sg13g2_fill_2 FILLER_71_605 ();
 sg13g2_fill_1 FILLER_71_607 ();
 sg13g2_fill_2 FILLER_71_631 ();
 sg13g2_fill_1 FILLER_71_633 ();
 sg13g2_decap_4 FILLER_71_660 ();
 sg13g2_fill_2 FILLER_71_686 ();
 sg13g2_decap_8 FILLER_71_730 ();
 sg13g2_decap_8 FILLER_71_737 ();
 sg13g2_decap_8 FILLER_71_744 ();
 sg13g2_decap_8 FILLER_71_751 ();
 sg13g2_decap_8 FILLER_71_758 ();
 sg13g2_decap_8 FILLER_71_765 ();
 sg13g2_decap_8 FILLER_71_772 ();
 sg13g2_decap_8 FILLER_71_779 ();
 sg13g2_decap_8 FILLER_71_786 ();
 sg13g2_decap_8 FILLER_71_793 ();
 sg13g2_decap_8 FILLER_71_800 ();
 sg13g2_decap_8 FILLER_71_807 ();
 sg13g2_decap_8 FILLER_71_814 ();
 sg13g2_decap_8 FILLER_71_821 ();
 sg13g2_decap_8 FILLER_71_828 ();
 sg13g2_decap_8 FILLER_71_835 ();
 sg13g2_decap_8 FILLER_71_842 ();
 sg13g2_decap_8 FILLER_71_849 ();
 sg13g2_decap_4 FILLER_71_856 ();
 sg13g2_fill_2 FILLER_71_860 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_1 FILLER_72_14 ();
 sg13g2_fill_2 FILLER_72_79 ();
 sg13g2_decap_4 FILLER_72_93 ();
 sg13g2_fill_1 FILLER_72_118 ();
 sg13g2_fill_2 FILLER_72_156 ();
 sg13g2_fill_1 FILLER_72_167 ();
 sg13g2_fill_1 FILLER_72_182 ();
 sg13g2_fill_1 FILLER_72_222 ();
 sg13g2_fill_2 FILLER_72_229 ();
 sg13g2_fill_1 FILLER_72_231 ();
 sg13g2_decap_8 FILLER_72_246 ();
 sg13g2_decap_8 FILLER_72_253 ();
 sg13g2_decap_4 FILLER_72_260 ();
 sg13g2_fill_1 FILLER_72_264 ();
 sg13g2_decap_4 FILLER_72_281 ();
 sg13g2_fill_2 FILLER_72_311 ();
 sg13g2_fill_2 FILLER_72_331 ();
 sg13g2_fill_1 FILLER_72_372 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_fill_2 FILLER_72_392 ();
 sg13g2_fill_1 FILLER_72_394 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_decap_8 FILLER_72_406 ();
 sg13g2_decap_8 FILLER_72_413 ();
 sg13g2_decap_8 FILLER_72_420 ();
 sg13g2_decap_8 FILLER_72_427 ();
 sg13g2_decap_8 FILLER_72_434 ();
 sg13g2_decap_8 FILLER_72_441 ();
 sg13g2_decap_8 FILLER_72_448 ();
 sg13g2_decap_8 FILLER_72_455 ();
 sg13g2_decap_8 FILLER_72_462 ();
 sg13g2_decap_8 FILLER_72_469 ();
 sg13g2_decap_8 FILLER_72_476 ();
 sg13g2_decap_8 FILLER_72_483 ();
 sg13g2_fill_2 FILLER_72_490 ();
 sg13g2_fill_2 FILLER_72_505 ();
 sg13g2_decap_4 FILLER_72_516 ();
 sg13g2_decap_4 FILLER_72_533 ();
 sg13g2_fill_2 FILLER_72_537 ();
 sg13g2_decap_8 FILLER_72_692 ();
 sg13g2_decap_8 FILLER_72_734 ();
 sg13g2_decap_8 FILLER_72_741 ();
 sg13g2_decap_8 FILLER_72_748 ();
 sg13g2_decap_8 FILLER_72_755 ();
 sg13g2_decap_8 FILLER_72_762 ();
 sg13g2_decap_8 FILLER_72_769 ();
 sg13g2_decap_8 FILLER_72_776 ();
 sg13g2_decap_8 FILLER_72_783 ();
 sg13g2_decap_8 FILLER_72_790 ();
 sg13g2_decap_8 FILLER_72_797 ();
 sg13g2_decap_8 FILLER_72_804 ();
 sg13g2_decap_8 FILLER_72_811 ();
 sg13g2_decap_8 FILLER_72_818 ();
 sg13g2_decap_8 FILLER_72_825 ();
 sg13g2_decap_8 FILLER_72_832 ();
 sg13g2_decap_8 FILLER_72_839 ();
 sg13g2_decap_8 FILLER_72_846 ();
 sg13g2_decap_8 FILLER_72_853 ();
 sg13g2_fill_2 FILLER_72_860 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_4 FILLER_73_28 ();
 sg13g2_fill_1 FILLER_73_32 ();
 sg13g2_fill_1 FILLER_73_69 ();
 sg13g2_decap_8 FILLER_73_96 ();
 sg13g2_fill_2 FILLER_73_103 ();
 sg13g2_decap_8 FILLER_73_115 ();
 sg13g2_decap_8 FILLER_73_122 ();
 sg13g2_fill_2 FILLER_73_129 ();
 sg13g2_decap_4 FILLER_73_153 ();
 sg13g2_decap_4 FILLER_73_162 ();
 sg13g2_fill_1 FILLER_73_166 ();
 sg13g2_fill_1 FILLER_73_171 ();
 sg13g2_decap_8 FILLER_73_181 ();
 sg13g2_fill_2 FILLER_73_188 ();
 sg13g2_fill_1 FILLER_73_197 ();
 sg13g2_decap_8 FILLER_73_208 ();
 sg13g2_fill_1 FILLER_73_215 ();
 sg13g2_fill_1 FILLER_73_221 ();
 sg13g2_fill_1 FILLER_73_230 ();
 sg13g2_decap_4 FILLER_73_236 ();
 sg13g2_fill_2 FILLER_73_240 ();
 sg13g2_decap_4 FILLER_73_245 ();
 sg13g2_fill_2 FILLER_73_306 ();
 sg13g2_fill_1 FILLER_73_308 ();
 sg13g2_fill_2 FILLER_73_329 ();
 sg13g2_fill_1 FILLER_73_336 ();
 sg13g2_decap_8 FILLER_73_367 ();
 sg13g2_decap_8 FILLER_73_374 ();
 sg13g2_decap_8 FILLER_73_381 ();
 sg13g2_decap_8 FILLER_73_388 ();
 sg13g2_decap_8 FILLER_73_395 ();
 sg13g2_decap_8 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_73_409 ();
 sg13g2_decap_8 FILLER_73_416 ();
 sg13g2_decap_8 FILLER_73_423 ();
 sg13g2_decap_8 FILLER_73_430 ();
 sg13g2_decap_8 FILLER_73_437 ();
 sg13g2_decap_8 FILLER_73_444 ();
 sg13g2_decap_8 FILLER_73_451 ();
 sg13g2_decap_8 FILLER_73_458 ();
 sg13g2_decap_8 FILLER_73_465 ();
 sg13g2_decap_8 FILLER_73_472 ();
 sg13g2_decap_8 FILLER_73_479 ();
 sg13g2_decap_8 FILLER_73_486 ();
 sg13g2_decap_8 FILLER_73_493 ();
 sg13g2_decap_4 FILLER_73_500 ();
 sg13g2_decap_8 FILLER_73_509 ();
 sg13g2_decap_8 FILLER_73_516 ();
 sg13g2_decap_8 FILLER_73_523 ();
 sg13g2_decap_8 FILLER_73_530 ();
 sg13g2_decap_8 FILLER_73_537 ();
 sg13g2_fill_2 FILLER_73_562 ();
 sg13g2_fill_1 FILLER_73_564 ();
 sg13g2_fill_2 FILLER_73_572 ();
 sg13g2_fill_1 FILLER_73_574 ();
 sg13g2_fill_2 FILLER_73_589 ();
 sg13g2_decap_8 FILLER_73_600 ();
 sg13g2_fill_2 FILLER_73_607 ();
 sg13g2_fill_1 FILLER_73_613 ();
 sg13g2_decap_8 FILLER_73_619 ();
 sg13g2_decap_8 FILLER_73_626 ();
 sg13g2_fill_1 FILLER_73_633 ();
 sg13g2_decap_8 FILLER_73_638 ();
 sg13g2_decap_4 FILLER_73_645 ();
 sg13g2_fill_2 FILLER_73_659 ();
 sg13g2_decap_8 FILLER_73_670 ();
 sg13g2_decap_8 FILLER_73_681 ();
 sg13g2_decap_8 FILLER_73_688 ();
 sg13g2_decap_8 FILLER_73_695 ();
 sg13g2_decap_8 FILLER_73_702 ();
 sg13g2_fill_1 FILLER_73_709 ();
 sg13g2_decap_8 FILLER_73_714 ();
 sg13g2_decap_8 FILLER_73_721 ();
 sg13g2_decap_8 FILLER_73_728 ();
 sg13g2_decap_8 FILLER_73_735 ();
 sg13g2_decap_8 FILLER_73_742 ();
 sg13g2_decap_8 FILLER_73_749 ();
 sg13g2_decap_8 FILLER_73_756 ();
 sg13g2_decap_8 FILLER_73_763 ();
 sg13g2_decap_8 FILLER_73_770 ();
 sg13g2_decap_8 FILLER_73_777 ();
 sg13g2_decap_8 FILLER_73_784 ();
 sg13g2_decap_8 FILLER_73_791 ();
 sg13g2_decap_8 FILLER_73_798 ();
 sg13g2_decap_8 FILLER_73_805 ();
 sg13g2_decap_8 FILLER_73_812 ();
 sg13g2_decap_8 FILLER_73_819 ();
 sg13g2_decap_8 FILLER_73_826 ();
 sg13g2_decap_8 FILLER_73_833 ();
 sg13g2_decap_8 FILLER_73_840 ();
 sg13g2_decap_8 FILLER_73_847 ();
 sg13g2_decap_8 FILLER_73_854 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_4 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_74 ();
 sg13g2_fill_2 FILLER_74_108 ();
 sg13g2_fill_1 FILLER_74_110 ();
 sg13g2_decap_4 FILLER_74_115 ();
 sg13g2_fill_2 FILLER_74_119 ();
 sg13g2_fill_1 FILLER_74_134 ();
 sg13g2_fill_2 FILLER_74_157 ();
 sg13g2_fill_2 FILLER_74_174 ();
 sg13g2_fill_1 FILLER_74_176 ();
 sg13g2_fill_2 FILLER_74_182 ();
 sg13g2_fill_2 FILLER_74_193 ();
 sg13g2_decap_4 FILLER_74_209 ();
 sg13g2_fill_1 FILLER_74_234 ();
 sg13g2_decap_4 FILLER_74_257 ();
 sg13g2_decap_4 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_269 ();
 sg13g2_fill_1 FILLER_74_278 ();
 sg13g2_fill_1 FILLER_74_284 ();
 sg13g2_fill_1 FILLER_74_351 ();
 sg13g2_decap_8 FILLER_74_356 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_decap_8 FILLER_74_370 ();
 sg13g2_decap_8 FILLER_74_377 ();
 sg13g2_decap_8 FILLER_74_384 ();
 sg13g2_decap_8 FILLER_74_391 ();
 sg13g2_decap_8 FILLER_74_398 ();
 sg13g2_decap_8 FILLER_74_405 ();
 sg13g2_decap_8 FILLER_74_412 ();
 sg13g2_decap_8 FILLER_74_419 ();
 sg13g2_decap_8 FILLER_74_426 ();
 sg13g2_decap_8 FILLER_74_433 ();
 sg13g2_decap_8 FILLER_74_440 ();
 sg13g2_decap_8 FILLER_74_447 ();
 sg13g2_decap_8 FILLER_74_454 ();
 sg13g2_decap_8 FILLER_74_461 ();
 sg13g2_decap_8 FILLER_74_468 ();
 sg13g2_decap_8 FILLER_74_475 ();
 sg13g2_decap_8 FILLER_74_482 ();
 sg13g2_decap_8 FILLER_74_489 ();
 sg13g2_decap_8 FILLER_74_496 ();
 sg13g2_decap_8 FILLER_74_503 ();
 sg13g2_decap_8 FILLER_74_510 ();
 sg13g2_decap_8 FILLER_74_517 ();
 sg13g2_decap_8 FILLER_74_524 ();
 sg13g2_decap_8 FILLER_74_531 ();
 sg13g2_decap_8 FILLER_74_538 ();
 sg13g2_decap_8 FILLER_74_545 ();
 sg13g2_decap_8 FILLER_74_552 ();
 sg13g2_fill_2 FILLER_74_559 ();
 sg13g2_decap_8 FILLER_74_566 ();
 sg13g2_fill_1 FILLER_74_573 ();
 sg13g2_decap_4 FILLER_74_578 ();
 sg13g2_decap_8 FILLER_74_591 ();
 sg13g2_decap_8 FILLER_74_598 ();
 sg13g2_decap_8 FILLER_74_605 ();
 sg13g2_decap_8 FILLER_74_612 ();
 sg13g2_decap_8 FILLER_74_619 ();
 sg13g2_decap_8 FILLER_74_626 ();
 sg13g2_decap_8 FILLER_74_633 ();
 sg13g2_decap_8 FILLER_74_640 ();
 sg13g2_decap_8 FILLER_74_647 ();
 sg13g2_decap_8 FILLER_74_658 ();
 sg13g2_decap_8 FILLER_74_665 ();
 sg13g2_decap_8 FILLER_74_672 ();
 sg13g2_decap_8 FILLER_74_679 ();
 sg13g2_decap_8 FILLER_74_686 ();
 sg13g2_decap_8 FILLER_74_693 ();
 sg13g2_decap_8 FILLER_74_700 ();
 sg13g2_decap_8 FILLER_74_707 ();
 sg13g2_decap_8 FILLER_74_714 ();
 sg13g2_decap_8 FILLER_74_721 ();
 sg13g2_decap_8 FILLER_74_728 ();
 sg13g2_decap_8 FILLER_74_735 ();
 sg13g2_decap_8 FILLER_74_742 ();
 sg13g2_decap_8 FILLER_74_749 ();
 sg13g2_decap_8 FILLER_74_756 ();
 sg13g2_decap_8 FILLER_74_763 ();
 sg13g2_decap_8 FILLER_74_770 ();
 sg13g2_decap_8 FILLER_74_777 ();
 sg13g2_decap_8 FILLER_74_784 ();
 sg13g2_decap_8 FILLER_74_791 ();
 sg13g2_decap_8 FILLER_74_798 ();
 sg13g2_decap_8 FILLER_74_805 ();
 sg13g2_decap_8 FILLER_74_812 ();
 sg13g2_decap_8 FILLER_74_819 ();
 sg13g2_decap_8 FILLER_74_826 ();
 sg13g2_decap_8 FILLER_74_833 ();
 sg13g2_decap_8 FILLER_74_840 ();
 sg13g2_decap_8 FILLER_74_847 ();
 sg13g2_decap_8 FILLER_74_854 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_fill_1 FILLER_75_42 ();
 sg13g2_fill_1 FILLER_75_62 ();
 sg13g2_fill_2 FILLER_75_77 ();
 sg13g2_fill_1 FILLER_75_79 ();
 sg13g2_decap_8 FILLER_75_100 ();
 sg13g2_fill_1 FILLER_75_107 ();
 sg13g2_fill_1 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_125 ();
 sg13g2_fill_2 FILLER_75_132 ();
 sg13g2_fill_1 FILLER_75_139 ();
 sg13g2_fill_2 FILLER_75_145 ();
 sg13g2_fill_1 FILLER_75_159 ();
 sg13g2_decap_8 FILLER_75_164 ();
 sg13g2_fill_1 FILLER_75_171 ();
 sg13g2_fill_1 FILLER_75_207 ();
 sg13g2_fill_2 FILLER_75_212 ();
 sg13g2_fill_2 FILLER_75_220 ();
 sg13g2_decap_8 FILLER_75_236 ();
 sg13g2_fill_1 FILLER_75_246 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_4 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_293 ();
 sg13g2_fill_1 FILLER_75_300 ();
 sg13g2_decap_8 FILLER_75_305 ();
 sg13g2_fill_2 FILLER_75_312 ();
 sg13g2_fill_1 FILLER_75_314 ();
 sg13g2_decap_8 FILLER_75_332 ();
 sg13g2_decap_8 FILLER_75_339 ();
 sg13g2_decap_8 FILLER_75_346 ();
 sg13g2_decap_8 FILLER_75_353 ();
 sg13g2_decap_8 FILLER_75_360 ();
 sg13g2_decap_8 FILLER_75_367 ();
 sg13g2_decap_8 FILLER_75_374 ();
 sg13g2_decap_8 FILLER_75_381 ();
 sg13g2_decap_8 FILLER_75_388 ();
 sg13g2_decap_8 FILLER_75_395 ();
 sg13g2_decap_8 FILLER_75_402 ();
 sg13g2_decap_8 FILLER_75_409 ();
 sg13g2_decap_8 FILLER_75_416 ();
 sg13g2_decap_8 FILLER_75_423 ();
 sg13g2_decap_8 FILLER_75_430 ();
 sg13g2_decap_8 FILLER_75_437 ();
 sg13g2_decap_8 FILLER_75_444 ();
 sg13g2_decap_8 FILLER_75_451 ();
 sg13g2_decap_8 FILLER_75_458 ();
 sg13g2_decap_8 FILLER_75_465 ();
 sg13g2_decap_8 FILLER_75_472 ();
 sg13g2_decap_8 FILLER_75_479 ();
 sg13g2_decap_8 FILLER_75_486 ();
 sg13g2_decap_8 FILLER_75_493 ();
 sg13g2_decap_8 FILLER_75_500 ();
 sg13g2_decap_8 FILLER_75_507 ();
 sg13g2_decap_8 FILLER_75_514 ();
 sg13g2_decap_8 FILLER_75_521 ();
 sg13g2_decap_8 FILLER_75_528 ();
 sg13g2_decap_8 FILLER_75_535 ();
 sg13g2_decap_8 FILLER_75_542 ();
 sg13g2_decap_8 FILLER_75_549 ();
 sg13g2_decap_8 FILLER_75_556 ();
 sg13g2_decap_8 FILLER_75_563 ();
 sg13g2_decap_8 FILLER_75_570 ();
 sg13g2_decap_8 FILLER_75_577 ();
 sg13g2_decap_8 FILLER_75_584 ();
 sg13g2_decap_8 FILLER_75_591 ();
 sg13g2_decap_8 FILLER_75_598 ();
 sg13g2_decap_8 FILLER_75_605 ();
 sg13g2_decap_8 FILLER_75_612 ();
 sg13g2_decap_8 FILLER_75_619 ();
 sg13g2_decap_8 FILLER_75_626 ();
 sg13g2_decap_8 FILLER_75_633 ();
 sg13g2_decap_8 FILLER_75_640 ();
 sg13g2_decap_8 FILLER_75_647 ();
 sg13g2_decap_8 FILLER_75_654 ();
 sg13g2_decap_8 FILLER_75_661 ();
 sg13g2_decap_8 FILLER_75_668 ();
 sg13g2_decap_8 FILLER_75_675 ();
 sg13g2_decap_8 FILLER_75_682 ();
 sg13g2_decap_8 FILLER_75_689 ();
 sg13g2_decap_8 FILLER_75_696 ();
 sg13g2_decap_8 FILLER_75_703 ();
 sg13g2_decap_8 FILLER_75_710 ();
 sg13g2_decap_8 FILLER_75_717 ();
 sg13g2_decap_8 FILLER_75_724 ();
 sg13g2_decap_8 FILLER_75_731 ();
 sg13g2_decap_8 FILLER_75_738 ();
 sg13g2_decap_8 FILLER_75_745 ();
 sg13g2_decap_8 FILLER_75_752 ();
 sg13g2_decap_8 FILLER_75_759 ();
 sg13g2_decap_8 FILLER_75_766 ();
 sg13g2_decap_8 FILLER_75_773 ();
 sg13g2_decap_8 FILLER_75_780 ();
 sg13g2_decap_8 FILLER_75_787 ();
 sg13g2_decap_8 FILLER_75_794 ();
 sg13g2_decap_8 FILLER_75_801 ();
 sg13g2_decap_8 FILLER_75_808 ();
 sg13g2_decap_8 FILLER_75_815 ();
 sg13g2_decap_8 FILLER_75_822 ();
 sg13g2_decap_8 FILLER_75_829 ();
 sg13g2_decap_8 FILLER_75_836 ();
 sg13g2_decap_8 FILLER_75_843 ();
 sg13g2_decap_8 FILLER_75_850 ();
 sg13g2_decap_4 FILLER_75_857 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_fill_1 FILLER_76_105 ();
 sg13g2_fill_1 FILLER_76_117 ();
 sg13g2_fill_2 FILLER_76_133 ();
 sg13g2_fill_1 FILLER_76_135 ();
 sg13g2_decap_8 FILLER_76_155 ();
 sg13g2_fill_2 FILLER_76_184 ();
 sg13g2_fill_1 FILLER_76_186 ();
 sg13g2_decap_8 FILLER_76_213 ();
 sg13g2_fill_1 FILLER_76_220 ();
 sg13g2_fill_2 FILLER_76_226 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_fill_1 FILLER_76_245 ();
 sg13g2_fill_1 FILLER_76_272 ();
 sg13g2_fill_1 FILLER_76_277 ();
 sg13g2_fill_2 FILLER_76_283 ();
 sg13g2_decap_8 FILLER_76_311 ();
 sg13g2_decap_8 FILLER_76_318 ();
 sg13g2_decap_8 FILLER_76_325 ();
 sg13g2_decap_8 FILLER_76_332 ();
 sg13g2_decap_8 FILLER_76_339 ();
 sg13g2_decap_8 FILLER_76_346 ();
 sg13g2_decap_8 FILLER_76_353 ();
 sg13g2_decap_8 FILLER_76_360 ();
 sg13g2_decap_8 FILLER_76_367 ();
 sg13g2_decap_8 FILLER_76_374 ();
 sg13g2_decap_8 FILLER_76_381 ();
 sg13g2_decap_8 FILLER_76_388 ();
 sg13g2_decap_8 FILLER_76_395 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_76_409 ();
 sg13g2_decap_8 FILLER_76_416 ();
 sg13g2_decap_8 FILLER_76_423 ();
 sg13g2_decap_8 FILLER_76_430 ();
 sg13g2_decap_8 FILLER_76_437 ();
 sg13g2_decap_8 FILLER_76_444 ();
 sg13g2_decap_8 FILLER_76_451 ();
 sg13g2_decap_8 FILLER_76_458 ();
 sg13g2_decap_8 FILLER_76_465 ();
 sg13g2_decap_8 FILLER_76_472 ();
 sg13g2_decap_8 FILLER_76_479 ();
 sg13g2_decap_8 FILLER_76_486 ();
 sg13g2_decap_8 FILLER_76_493 ();
 sg13g2_decap_8 FILLER_76_500 ();
 sg13g2_decap_8 FILLER_76_507 ();
 sg13g2_decap_8 FILLER_76_514 ();
 sg13g2_decap_8 FILLER_76_521 ();
 sg13g2_decap_8 FILLER_76_528 ();
 sg13g2_decap_8 FILLER_76_535 ();
 sg13g2_decap_8 FILLER_76_542 ();
 sg13g2_decap_8 FILLER_76_549 ();
 sg13g2_decap_8 FILLER_76_556 ();
 sg13g2_decap_8 FILLER_76_563 ();
 sg13g2_decap_8 FILLER_76_570 ();
 sg13g2_decap_8 FILLER_76_577 ();
 sg13g2_decap_8 FILLER_76_584 ();
 sg13g2_decap_8 FILLER_76_591 ();
 sg13g2_decap_8 FILLER_76_598 ();
 sg13g2_decap_8 FILLER_76_605 ();
 sg13g2_decap_8 FILLER_76_612 ();
 sg13g2_decap_8 FILLER_76_619 ();
 sg13g2_decap_8 FILLER_76_626 ();
 sg13g2_decap_8 FILLER_76_633 ();
 sg13g2_decap_8 FILLER_76_640 ();
 sg13g2_decap_8 FILLER_76_647 ();
 sg13g2_decap_8 FILLER_76_654 ();
 sg13g2_decap_8 FILLER_76_661 ();
 sg13g2_decap_8 FILLER_76_668 ();
 sg13g2_decap_8 FILLER_76_675 ();
 sg13g2_decap_8 FILLER_76_682 ();
 sg13g2_decap_8 FILLER_76_689 ();
 sg13g2_decap_8 FILLER_76_696 ();
 sg13g2_decap_8 FILLER_76_703 ();
 sg13g2_decap_8 FILLER_76_710 ();
 sg13g2_decap_8 FILLER_76_717 ();
 sg13g2_decap_8 FILLER_76_724 ();
 sg13g2_decap_8 FILLER_76_731 ();
 sg13g2_decap_8 FILLER_76_738 ();
 sg13g2_decap_8 FILLER_76_745 ();
 sg13g2_decap_8 FILLER_76_752 ();
 sg13g2_decap_8 FILLER_76_759 ();
 sg13g2_decap_8 FILLER_76_766 ();
 sg13g2_decap_8 FILLER_76_773 ();
 sg13g2_decap_8 FILLER_76_780 ();
 sg13g2_decap_8 FILLER_76_787 ();
 sg13g2_decap_8 FILLER_76_794 ();
 sg13g2_decap_8 FILLER_76_801 ();
 sg13g2_decap_8 FILLER_76_808 ();
 sg13g2_decap_8 FILLER_76_815 ();
 sg13g2_decap_8 FILLER_76_822 ();
 sg13g2_decap_8 FILLER_76_829 ();
 sg13g2_decap_8 FILLER_76_836 ();
 sg13g2_decap_8 FILLER_76_843 ();
 sg13g2_decap_8 FILLER_76_850 ();
 sg13g2_decap_4 FILLER_76_857 ();
 sg13g2_fill_1 FILLER_76_861 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_fill_1 FILLER_77_42 ();
 sg13g2_fill_1 FILLER_77_83 ();
 sg13g2_decap_4 FILLER_77_127 ();
 sg13g2_fill_2 FILLER_77_177 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_fill_2 FILLER_77_196 ();
 sg13g2_fill_2 FILLER_77_204 ();
 sg13g2_fill_1 FILLER_77_206 ();
 sg13g2_decap_4 FILLER_77_212 ();
 sg13g2_fill_2 FILLER_77_216 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_4 FILLER_77_252 ();
 sg13g2_fill_1 FILLER_77_256 ();
 sg13g2_decap_8 FILLER_77_261 ();
 sg13g2_decap_8 FILLER_77_268 ();
 sg13g2_decap_8 FILLER_77_275 ();
 sg13g2_decap_8 FILLER_77_282 ();
 sg13g2_decap_8 FILLER_77_289 ();
 sg13g2_decap_8 FILLER_77_300 ();
 sg13g2_decap_8 FILLER_77_307 ();
 sg13g2_decap_8 FILLER_77_314 ();
 sg13g2_decap_8 FILLER_77_321 ();
 sg13g2_decap_8 FILLER_77_328 ();
 sg13g2_decap_8 FILLER_77_335 ();
 sg13g2_decap_8 FILLER_77_342 ();
 sg13g2_decap_8 FILLER_77_349 ();
 sg13g2_decap_8 FILLER_77_356 ();
 sg13g2_decap_8 FILLER_77_363 ();
 sg13g2_decap_8 FILLER_77_370 ();
 sg13g2_decap_8 FILLER_77_377 ();
 sg13g2_decap_8 FILLER_77_384 ();
 sg13g2_decap_8 FILLER_77_391 ();
 sg13g2_decap_8 FILLER_77_398 ();
 sg13g2_decap_8 FILLER_77_405 ();
 sg13g2_decap_8 FILLER_77_412 ();
 sg13g2_decap_8 FILLER_77_419 ();
 sg13g2_decap_8 FILLER_77_426 ();
 sg13g2_decap_8 FILLER_77_433 ();
 sg13g2_decap_8 FILLER_77_440 ();
 sg13g2_decap_8 FILLER_77_447 ();
 sg13g2_decap_8 FILLER_77_454 ();
 sg13g2_decap_8 FILLER_77_461 ();
 sg13g2_decap_8 FILLER_77_468 ();
 sg13g2_decap_8 FILLER_77_475 ();
 sg13g2_decap_8 FILLER_77_482 ();
 sg13g2_decap_8 FILLER_77_489 ();
 sg13g2_decap_8 FILLER_77_496 ();
 sg13g2_decap_8 FILLER_77_503 ();
 sg13g2_decap_8 FILLER_77_510 ();
 sg13g2_decap_8 FILLER_77_517 ();
 sg13g2_decap_8 FILLER_77_524 ();
 sg13g2_decap_8 FILLER_77_531 ();
 sg13g2_decap_8 FILLER_77_538 ();
 sg13g2_decap_8 FILLER_77_545 ();
 sg13g2_decap_8 FILLER_77_552 ();
 sg13g2_decap_8 FILLER_77_559 ();
 sg13g2_decap_8 FILLER_77_566 ();
 sg13g2_decap_8 FILLER_77_573 ();
 sg13g2_decap_8 FILLER_77_580 ();
 sg13g2_decap_8 FILLER_77_587 ();
 sg13g2_decap_8 FILLER_77_594 ();
 sg13g2_decap_8 FILLER_77_601 ();
 sg13g2_decap_8 FILLER_77_608 ();
 sg13g2_decap_8 FILLER_77_615 ();
 sg13g2_decap_8 FILLER_77_622 ();
 sg13g2_decap_8 FILLER_77_629 ();
 sg13g2_decap_8 FILLER_77_636 ();
 sg13g2_decap_8 FILLER_77_643 ();
 sg13g2_decap_8 FILLER_77_650 ();
 sg13g2_decap_8 FILLER_77_657 ();
 sg13g2_decap_8 FILLER_77_664 ();
 sg13g2_decap_8 FILLER_77_671 ();
 sg13g2_decap_8 FILLER_77_678 ();
 sg13g2_decap_8 FILLER_77_685 ();
 sg13g2_decap_8 FILLER_77_692 ();
 sg13g2_decap_8 FILLER_77_699 ();
 sg13g2_decap_8 FILLER_77_706 ();
 sg13g2_decap_8 FILLER_77_713 ();
 sg13g2_decap_8 FILLER_77_720 ();
 sg13g2_decap_8 FILLER_77_727 ();
 sg13g2_decap_8 FILLER_77_734 ();
 sg13g2_decap_8 FILLER_77_741 ();
 sg13g2_decap_8 FILLER_77_748 ();
 sg13g2_decap_8 FILLER_77_755 ();
 sg13g2_decap_8 FILLER_77_762 ();
 sg13g2_decap_8 FILLER_77_769 ();
 sg13g2_decap_8 FILLER_77_776 ();
 sg13g2_decap_8 FILLER_77_783 ();
 sg13g2_decap_8 FILLER_77_790 ();
 sg13g2_decap_8 FILLER_77_797 ();
 sg13g2_decap_8 FILLER_77_804 ();
 sg13g2_decap_8 FILLER_77_811 ();
 sg13g2_decap_8 FILLER_77_818 ();
 sg13g2_decap_8 FILLER_77_825 ();
 sg13g2_decap_8 FILLER_77_832 ();
 sg13g2_decap_8 FILLER_77_839 ();
 sg13g2_decap_8 FILLER_77_846 ();
 sg13g2_decap_8 FILLER_77_853 ();
 sg13g2_fill_2 FILLER_77_860 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_fill_1 FILLER_78_56 ();
 sg13g2_fill_2 FILLER_78_75 ();
 sg13g2_fill_2 FILLER_78_90 ();
 sg13g2_fill_1 FILLER_78_92 ();
 sg13g2_decap_8 FILLER_78_108 ();
 sg13g2_decap_8 FILLER_78_115 ();
 sg13g2_decap_8 FILLER_78_122 ();
 sg13g2_fill_2 FILLER_78_129 ();
 sg13g2_fill_1 FILLER_78_131 ();
 sg13g2_fill_1 FILLER_78_137 ();
 sg13g2_fill_2 FILLER_78_159 ();
 sg13g2_fill_2 FILLER_78_187 ();
 sg13g2_fill_1 FILLER_78_189 ();
 sg13g2_decap_4 FILLER_78_195 ();
 sg13g2_fill_1 FILLER_78_199 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_441 ();
 sg13g2_decap_8 FILLER_78_448 ();
 sg13g2_decap_8 FILLER_78_455 ();
 sg13g2_decap_8 FILLER_78_462 ();
 sg13g2_decap_8 FILLER_78_469 ();
 sg13g2_decap_8 FILLER_78_476 ();
 sg13g2_decap_8 FILLER_78_483 ();
 sg13g2_decap_8 FILLER_78_490 ();
 sg13g2_decap_8 FILLER_78_497 ();
 sg13g2_decap_8 FILLER_78_504 ();
 sg13g2_decap_8 FILLER_78_511 ();
 sg13g2_decap_8 FILLER_78_518 ();
 sg13g2_decap_8 FILLER_78_525 ();
 sg13g2_decap_8 FILLER_78_532 ();
 sg13g2_decap_8 FILLER_78_539 ();
 sg13g2_decap_8 FILLER_78_546 ();
 sg13g2_decap_8 FILLER_78_553 ();
 sg13g2_decap_8 FILLER_78_560 ();
 sg13g2_decap_8 FILLER_78_567 ();
 sg13g2_decap_8 FILLER_78_574 ();
 sg13g2_decap_8 FILLER_78_581 ();
 sg13g2_decap_8 FILLER_78_588 ();
 sg13g2_decap_8 FILLER_78_595 ();
 sg13g2_decap_8 FILLER_78_602 ();
 sg13g2_decap_8 FILLER_78_609 ();
 sg13g2_decap_8 FILLER_78_616 ();
 sg13g2_decap_8 FILLER_78_623 ();
 sg13g2_decap_8 FILLER_78_630 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_decap_8 FILLER_78_644 ();
 sg13g2_decap_8 FILLER_78_651 ();
 sg13g2_decap_8 FILLER_78_658 ();
 sg13g2_decap_8 FILLER_78_665 ();
 sg13g2_decap_8 FILLER_78_672 ();
 sg13g2_decap_8 FILLER_78_679 ();
 sg13g2_decap_8 FILLER_78_686 ();
 sg13g2_decap_8 FILLER_78_693 ();
 sg13g2_decap_8 FILLER_78_700 ();
 sg13g2_decap_8 FILLER_78_707 ();
 sg13g2_decap_8 FILLER_78_714 ();
 sg13g2_decap_8 FILLER_78_721 ();
 sg13g2_decap_8 FILLER_78_728 ();
 sg13g2_decap_8 FILLER_78_735 ();
 sg13g2_decap_8 FILLER_78_742 ();
 sg13g2_decap_8 FILLER_78_749 ();
 sg13g2_decap_8 FILLER_78_756 ();
 sg13g2_decap_8 FILLER_78_763 ();
 sg13g2_decap_8 FILLER_78_770 ();
 sg13g2_decap_8 FILLER_78_777 ();
 sg13g2_decap_8 FILLER_78_784 ();
 sg13g2_decap_8 FILLER_78_791 ();
 sg13g2_decap_8 FILLER_78_798 ();
 sg13g2_decap_8 FILLER_78_805 ();
 sg13g2_decap_8 FILLER_78_812 ();
 sg13g2_decap_8 FILLER_78_819 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_decap_8 FILLER_78_833 ();
 sg13g2_decap_8 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_decap_8 FILLER_78_854 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_4 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_79 ();
 sg13g2_decap_8 FILLER_79_86 ();
 sg13g2_fill_1 FILLER_79_93 ();
 sg13g2_decap_8 FILLER_79_104 ();
 sg13g2_decap_8 FILLER_79_111 ();
 sg13g2_fill_1 FILLER_79_118 ();
 sg13g2_decap_8 FILLER_79_135 ();
 sg13g2_decap_4 FILLER_79_142 ();
 sg13g2_fill_1 FILLER_79_146 ();
 sg13g2_decap_4 FILLER_79_163 ();
 sg13g2_fill_1 FILLER_79_167 ();
 sg13g2_fill_1 FILLER_79_192 ();
 sg13g2_fill_2 FILLER_79_197 ();
 sg13g2_fill_1 FILLER_79_199 ();
 sg13g2_decap_8 FILLER_79_207 ();
 sg13g2_decap_8 FILLER_79_214 ();
 sg13g2_decap_8 FILLER_79_221 ();
 sg13g2_decap_8 FILLER_79_228 ();
 sg13g2_decap_8 FILLER_79_235 ();
 sg13g2_decap_8 FILLER_79_242 ();
 sg13g2_decap_8 FILLER_79_249 ();
 sg13g2_decap_8 FILLER_79_256 ();
 sg13g2_decap_8 FILLER_79_263 ();
 sg13g2_decap_8 FILLER_79_270 ();
 sg13g2_decap_8 FILLER_79_277 ();
 sg13g2_decap_8 FILLER_79_284 ();
 sg13g2_decap_8 FILLER_79_291 ();
 sg13g2_decap_8 FILLER_79_298 ();
 sg13g2_decap_8 FILLER_79_305 ();
 sg13g2_decap_8 FILLER_79_312 ();
 sg13g2_decap_8 FILLER_79_319 ();
 sg13g2_decap_8 FILLER_79_326 ();
 sg13g2_decap_8 FILLER_79_333 ();
 sg13g2_decap_8 FILLER_79_340 ();
 sg13g2_decap_8 FILLER_79_347 ();
 sg13g2_decap_8 FILLER_79_354 ();
 sg13g2_decap_8 FILLER_79_361 ();
 sg13g2_decap_8 FILLER_79_368 ();
 sg13g2_decap_8 FILLER_79_375 ();
 sg13g2_decap_8 FILLER_79_382 ();
 sg13g2_decap_8 FILLER_79_389 ();
 sg13g2_decap_8 FILLER_79_396 ();
 sg13g2_decap_8 FILLER_79_403 ();
 sg13g2_decap_8 FILLER_79_410 ();
 sg13g2_decap_8 FILLER_79_417 ();
 sg13g2_decap_8 FILLER_79_424 ();
 sg13g2_decap_8 FILLER_79_431 ();
 sg13g2_decap_8 FILLER_79_438 ();
 sg13g2_decap_8 FILLER_79_445 ();
 sg13g2_decap_8 FILLER_79_452 ();
 sg13g2_decap_8 FILLER_79_459 ();
 sg13g2_decap_8 FILLER_79_466 ();
 sg13g2_decap_8 FILLER_79_473 ();
 sg13g2_decap_8 FILLER_79_480 ();
 sg13g2_decap_8 FILLER_79_487 ();
 sg13g2_decap_8 FILLER_79_494 ();
 sg13g2_decap_8 FILLER_79_501 ();
 sg13g2_decap_8 FILLER_79_508 ();
 sg13g2_decap_8 FILLER_79_515 ();
 sg13g2_decap_8 FILLER_79_522 ();
 sg13g2_decap_8 FILLER_79_529 ();
 sg13g2_decap_8 FILLER_79_536 ();
 sg13g2_decap_8 FILLER_79_543 ();
 sg13g2_decap_8 FILLER_79_550 ();
 sg13g2_decap_8 FILLER_79_557 ();
 sg13g2_decap_8 FILLER_79_564 ();
 sg13g2_decap_8 FILLER_79_571 ();
 sg13g2_decap_8 FILLER_79_578 ();
 sg13g2_decap_8 FILLER_79_585 ();
 sg13g2_decap_8 FILLER_79_592 ();
 sg13g2_decap_8 FILLER_79_599 ();
 sg13g2_decap_8 FILLER_79_606 ();
 sg13g2_decap_8 FILLER_79_613 ();
 sg13g2_decap_8 FILLER_79_620 ();
 sg13g2_decap_8 FILLER_79_627 ();
 sg13g2_decap_8 FILLER_79_634 ();
 sg13g2_decap_8 FILLER_79_641 ();
 sg13g2_decap_8 FILLER_79_648 ();
 sg13g2_decap_8 FILLER_79_655 ();
 sg13g2_decap_8 FILLER_79_662 ();
 sg13g2_decap_8 FILLER_79_669 ();
 sg13g2_decap_8 FILLER_79_676 ();
 sg13g2_decap_8 FILLER_79_683 ();
 sg13g2_decap_8 FILLER_79_690 ();
 sg13g2_decap_8 FILLER_79_697 ();
 sg13g2_decap_8 FILLER_79_704 ();
 sg13g2_decap_8 FILLER_79_711 ();
 sg13g2_decap_8 FILLER_79_718 ();
 sg13g2_decap_8 FILLER_79_725 ();
 sg13g2_decap_8 FILLER_79_732 ();
 sg13g2_decap_8 FILLER_79_739 ();
 sg13g2_decap_8 FILLER_79_746 ();
 sg13g2_decap_8 FILLER_79_753 ();
 sg13g2_decap_8 FILLER_79_760 ();
 sg13g2_decap_8 FILLER_79_767 ();
 sg13g2_decap_8 FILLER_79_774 ();
 sg13g2_decap_8 FILLER_79_781 ();
 sg13g2_decap_8 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_795 ();
 sg13g2_decap_8 FILLER_79_802 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_851 ();
 sg13g2_decap_4 FILLER_79_858 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_fill_2 FILLER_80_157 ();
 sg13g2_fill_1 FILLER_80_159 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_fill_2 FILLER_80_176 ();
 sg13g2_decap_8 FILLER_80_186 ();
 sg13g2_decap_8 FILLER_80_193 ();
 sg13g2_decap_8 FILLER_80_200 ();
 sg13g2_decap_8 FILLER_80_207 ();
 sg13g2_decap_8 FILLER_80_214 ();
 sg13g2_decap_8 FILLER_80_221 ();
 sg13g2_decap_8 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_235 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_decap_8 FILLER_80_249 ();
 sg13g2_decap_8 FILLER_80_256 ();
 sg13g2_decap_8 FILLER_80_263 ();
 sg13g2_decap_8 FILLER_80_270 ();
 sg13g2_decap_8 FILLER_80_277 ();
 sg13g2_decap_8 FILLER_80_284 ();
 sg13g2_decap_8 FILLER_80_291 ();
 sg13g2_decap_8 FILLER_80_298 ();
 sg13g2_decap_8 FILLER_80_305 ();
 sg13g2_decap_8 FILLER_80_312 ();
 sg13g2_decap_8 FILLER_80_319 ();
 sg13g2_decap_8 FILLER_80_326 ();
 sg13g2_decap_8 FILLER_80_333 ();
 sg13g2_decap_8 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_347 ();
 sg13g2_decap_8 FILLER_80_354 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_decap_8 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_382 ();
 sg13g2_decap_8 FILLER_80_389 ();
 sg13g2_decap_8 FILLER_80_396 ();
 sg13g2_decap_8 FILLER_80_403 ();
 sg13g2_decap_8 FILLER_80_410 ();
 sg13g2_decap_8 FILLER_80_417 ();
 sg13g2_decap_8 FILLER_80_424 ();
 sg13g2_decap_8 FILLER_80_431 ();
 sg13g2_decap_8 FILLER_80_438 ();
 sg13g2_decap_8 FILLER_80_445 ();
 sg13g2_decap_8 FILLER_80_452 ();
 sg13g2_decap_8 FILLER_80_459 ();
 sg13g2_decap_8 FILLER_80_466 ();
 sg13g2_decap_8 FILLER_80_473 ();
 sg13g2_decap_8 FILLER_80_480 ();
 sg13g2_decap_8 FILLER_80_487 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_8 FILLER_80_508 ();
 sg13g2_decap_8 FILLER_80_515 ();
 sg13g2_decap_8 FILLER_80_522 ();
 sg13g2_decap_8 FILLER_80_529 ();
 sg13g2_decap_8 FILLER_80_536 ();
 sg13g2_decap_8 FILLER_80_543 ();
 sg13g2_decap_8 FILLER_80_550 ();
 sg13g2_decap_8 FILLER_80_557 ();
 sg13g2_decap_8 FILLER_80_564 ();
 sg13g2_decap_8 FILLER_80_571 ();
 sg13g2_decap_8 FILLER_80_578 ();
 sg13g2_decap_8 FILLER_80_585 ();
 sg13g2_decap_8 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_599 ();
 sg13g2_decap_8 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_613 ();
 sg13g2_decap_8 FILLER_80_620 ();
 sg13g2_decap_8 FILLER_80_627 ();
 sg13g2_decap_8 FILLER_80_634 ();
 sg13g2_decap_8 FILLER_80_641 ();
 sg13g2_decap_8 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_655 ();
 sg13g2_decap_8 FILLER_80_662 ();
 sg13g2_decap_8 FILLER_80_669 ();
 sg13g2_decap_8 FILLER_80_676 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_decap_8 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_697 ();
 sg13g2_decap_8 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_711 ();
 sg13g2_decap_8 FILLER_80_718 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_decap_8 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_739 ();
 sg13g2_decap_8 FILLER_80_746 ();
 sg13g2_decap_8 FILLER_80_753 ();
 sg13g2_decap_8 FILLER_80_760 ();
 sg13g2_decap_8 FILLER_80_767 ();
 sg13g2_decap_8 FILLER_80_774 ();
 sg13g2_decap_8 FILLER_80_781 ();
 sg13g2_decap_8 FILLER_80_788 ();
 sg13g2_decap_8 FILLER_80_795 ();
 sg13g2_decap_8 FILLER_80_802 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_decap_8 FILLER_80_830 ();
 sg13g2_decap_8 FILLER_80_837 ();
 sg13g2_decap_8 FILLER_80_844 ();
 sg13g2_decap_8 FILLER_80_851 ();
 sg13g2_decap_4 FILLER_80_858 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net433;
 assign uio_out[0] = net8;
 assign uio_out[1] = net9;
 assign uio_out[2] = net10;
 assign uio_out[3] = net11;
 assign uio_out[4] = net12;
 assign uio_out[5] = net13;
 assign uio_out[6] = net14;
endmodule

module tt_um_a1k0n_vgadonut (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire clknet_leaf_0_clk;
 wire hsync;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire \vgadonut.bayer_j[0] ;
 wire \vgadonut.bayer_j[1] ;
 wire \vgadonut.donut.cA[0] ;
 wire \vgadonut.donut.cA[10] ;
 wire \vgadonut.donut.cA[11] ;
 wire \vgadonut.donut.cA[12] ;
 wire \vgadonut.donut.cA[13] ;
 wire \vgadonut.donut.cA[14] ;
 wire \vgadonut.donut.cA[15] ;
 wire \vgadonut.donut.cA[1] ;
 wire \vgadonut.donut.cA[2] ;
 wire \vgadonut.donut.cA[3] ;
 wire \vgadonut.donut.cA[4] ;
 wire \vgadonut.donut.cA[5] ;
 wire \vgadonut.donut.cA[6] ;
 wire \vgadonut.donut.cA[7] ;
 wire \vgadonut.donut.cA[8] ;
 wire \vgadonut.donut.cA[9] ;
 wire \vgadonut.donut.cAcB[0] ;
 wire \vgadonut.donut.cAcB[10] ;
 wire \vgadonut.donut.cAcB[11] ;
 wire \vgadonut.donut.cAcB[12] ;
 wire \vgadonut.donut.cAcB[13] ;
 wire \vgadonut.donut.cAcB[14] ;
 wire \vgadonut.donut.cAcB[15] ;
 wire \vgadonut.donut.cAcB[1] ;
 wire \vgadonut.donut.cAcB[2] ;
 wire \vgadonut.donut.cAcB[3] ;
 wire \vgadonut.donut.cAcB[4] ;
 wire \vgadonut.donut.cAcB[5] ;
 wire \vgadonut.donut.cAcB[6] ;
 wire \vgadonut.donut.cAcB[7] ;
 wire \vgadonut.donut.cAcB[8] ;
 wire \vgadonut.donut.cAcB[9] ;
 wire \vgadonut.donut.cAsB[0] ;
 wire \vgadonut.donut.cAsB[10] ;
 wire \vgadonut.donut.cAsB[11] ;
 wire \vgadonut.donut.cAsB[12] ;
 wire \vgadonut.donut.cAsB[13] ;
 wire \vgadonut.donut.cAsB[14] ;
 wire \vgadonut.donut.cAsB[15] ;
 wire \vgadonut.donut.cAsB[1] ;
 wire \vgadonut.donut.cAsB[2] ;
 wire \vgadonut.donut.cAsB[3] ;
 wire \vgadonut.donut.cAsB[4] ;
 wire \vgadonut.donut.cAsB[5] ;
 wire \vgadonut.donut.cAsB[6] ;
 wire \vgadonut.donut.cAsB[7] ;
 wire \vgadonut.donut.cAsB[8] ;
 wire \vgadonut.donut.cAsB[9] ;
 wire \vgadonut.donut.cB[0] ;
 wire \vgadonut.donut.cB[10] ;
 wire \vgadonut.donut.cB[11] ;
 wire \vgadonut.donut.cB[12] ;
 wire \vgadonut.donut.cB[13] ;
 wire \vgadonut.donut.cB[14] ;
 wire \vgadonut.donut.cB[15] ;
 wire \vgadonut.donut.cB[1] ;
 wire \vgadonut.donut.cB[2] ;
 wire \vgadonut.donut.cB[3] ;
 wire \vgadonut.donut.cB[4] ;
 wire \vgadonut.donut.cB[5] ;
 wire \vgadonut.donut.cB[6] ;
 wire \vgadonut.donut.cB[7] ;
 wire \vgadonut.donut.cB[8] ;
 wire \vgadonut.donut.cB[9] ;
 wire \vgadonut.donut.donut_luma[0] ;
 wire \vgadonut.donut.donut_luma[1] ;
 wire \vgadonut.donut.donut_luma[2] ;
 wire \vgadonut.donut.donut_luma[3] ;
 wire \vgadonut.donut.donut_luma[4] ;
 wire \vgadonut.donut.donut_luma[5] ;
 wire \vgadonut.donut.donut_visible ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[0] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[10] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[11] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[12] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[13] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[1] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[2] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[3] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[4] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[5] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[6] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[7] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[8] ;
 wire \vgadonut.donut.donuthit.cordicxy.x2in[9] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[0] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[10] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[11] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[12] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[13] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[14] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[15] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[1] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[2] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[3] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[4] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[5] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[6] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[7] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[8] ;
 wire \vgadonut.donut.donuthit.cordicxy.xin[9] ;
 wire \vgadonut.donut.donuthit.cordicxy.xinvert ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[0] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[10] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[11] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[12] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[13] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[14] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[1] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[2] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[3] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[4] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[5] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[6] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[7] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[8] ;
 wire \vgadonut.donut.donuthit.cordicxy.yin[9] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[10] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[11] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[12] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[13] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[8] ;
 wire \vgadonut.donut.donuthit.cordicxz.x2out[9] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[0] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[10] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[11] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[12] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[13] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[14] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[15] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[1] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[2] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[3] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[4] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[5] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[6] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[7] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[8] ;
 wire \vgadonut.donut.donuthit.cordicxz.xin[9] ;
 wire \vgadonut.donut.donuthit.hit ;
 wire \vgadonut.donut.donuthit.light[10] ;
 wire \vgadonut.donut.donuthit.light[11] ;
 wire \vgadonut.donut.donuthit.light[12] ;
 wire \vgadonut.donut.donuthit.light[13] ;
 wire \vgadonut.donut.donuthit.light[8] ;
 wire \vgadonut.donut.donuthit.light[9] ;
 wire \vgadonut.donut.donuthit.rx[10] ;
 wire \vgadonut.donut.donuthit.rx[11] ;
 wire \vgadonut.donut.donuthit.rx[12] ;
 wire \vgadonut.donut.donuthit.rx[13] ;
 wire \vgadonut.donut.donuthit.rx[14] ;
 wire \vgadonut.donut.donuthit.rx[15] ;
 wire \vgadonut.donut.donuthit.rx[5] ;
 wire \vgadonut.donut.donuthit.rx[6] ;
 wire \vgadonut.donut.donuthit.rx[7] ;
 wire \vgadonut.donut.donuthit.rx[8] ;
 wire \vgadonut.donut.donuthit.rx[9] ;
 wire \vgadonut.donut.donuthit.rxin[0] ;
 wire \vgadonut.donut.donuthit.rxin[10] ;
 wire \vgadonut.donut.donuthit.rxin[11] ;
 wire \vgadonut.donut.donuthit.rxin[12] ;
 wire \vgadonut.donut.donuthit.rxin[13] ;
 wire \vgadonut.donut.donuthit.rxin[14] ;
 wire \vgadonut.donut.donuthit.rxin[15] ;
 wire \vgadonut.donut.donuthit.rxin[1] ;
 wire \vgadonut.donut.donuthit.rxin[2] ;
 wire \vgadonut.donut.donuthit.rxin[3] ;
 wire \vgadonut.donut.donuthit.rxin[4] ;
 wire \vgadonut.donut.donuthit.rxin[5] ;
 wire \vgadonut.donut.donuthit.rxin[6] ;
 wire \vgadonut.donut.donuthit.rxin[7] ;
 wire \vgadonut.donut.donuthit.rxin[8] ;
 wire \vgadonut.donut.donuthit.rxin[9] ;
 wire \vgadonut.donut.donuthit.ry[10] ;
 wire \vgadonut.donut.donuthit.ry[11] ;
 wire \vgadonut.donut.donuthit.ry[12] ;
 wire \vgadonut.donut.donuthit.ry[13] ;
 wire \vgadonut.donut.donuthit.ry[14] ;
 wire \vgadonut.donut.donuthit.ry[15] ;
 wire \vgadonut.donut.donuthit.ry[5] ;
 wire \vgadonut.donut.donuthit.ry[6] ;
 wire \vgadonut.donut.donuthit.ry[7] ;
 wire \vgadonut.donut.donuthit.ry[8] ;
 wire \vgadonut.donut.donuthit.ry[9] ;
 wire \vgadonut.donut.donuthit.ryin[0] ;
 wire \vgadonut.donut.donuthit.ryin[10] ;
 wire \vgadonut.donut.donuthit.ryin[11] ;
 wire \vgadonut.donut.donuthit.ryin[12] ;
 wire \vgadonut.donut.donuthit.ryin[13] ;
 wire \vgadonut.donut.donuthit.ryin[14] ;
 wire \vgadonut.donut.donuthit.ryin[15] ;
 wire \vgadonut.donut.donuthit.ryin[1] ;
 wire \vgadonut.donut.donuthit.ryin[2] ;
 wire \vgadonut.donut.donuthit.ryin[3] ;
 wire \vgadonut.donut.donuthit.ryin[4] ;
 wire \vgadonut.donut.donuthit.ryin[5] ;
 wire \vgadonut.donut.donuthit.ryin[6] ;
 wire \vgadonut.donut.donuthit.ryin[7] ;
 wire \vgadonut.donut.donuthit.ryin[8] ;
 wire \vgadonut.donut.donuthit.ryin[9] ;
 wire \vgadonut.donut.donuthit.rz[10] ;
 wire \vgadonut.donut.donuthit.rz[11] ;
 wire \vgadonut.donut.donuthit.rz[12] ;
 wire \vgadonut.donut.donuthit.rz[13] ;
 wire \vgadonut.donut.donuthit.rz[14] ;
 wire \vgadonut.donut.donuthit.rz[15] ;
 wire \vgadonut.donut.donuthit.rz[5] ;
 wire \vgadonut.donut.donuthit.rz[6] ;
 wire \vgadonut.donut.donuthit.rz[7] ;
 wire \vgadonut.donut.donuthit.rz[8] ;
 wire \vgadonut.donut.donuthit.rz[9] ;
 wire \vgadonut.donut.donuthit.rzin[0] ;
 wire \vgadonut.donut.donuthit.rzin[10] ;
 wire \vgadonut.donut.donuthit.rzin[11] ;
 wire \vgadonut.donut.donuthit.rzin[12] ;
 wire \vgadonut.donut.donuthit.rzin[13] ;
 wire \vgadonut.donut.donuthit.rzin[14] ;
 wire \vgadonut.donut.donuthit.rzin[15] ;
 wire \vgadonut.donut.donuthit.rzin[1] ;
 wire \vgadonut.donut.donuthit.rzin[2] ;
 wire \vgadonut.donut.donuthit.rzin[3] ;
 wire \vgadonut.donut.donuthit.rzin[4] ;
 wire \vgadonut.donut.donuthit.rzin[5] ;
 wire \vgadonut.donut.donuthit.rzin[6] ;
 wire \vgadonut.donut.donuthit.rzin[7] ;
 wire \vgadonut.donut.donuthit.rzin[8] ;
 wire \vgadonut.donut.donuthit.rzin[9] ;
 wire \vgadonut.donut.donuthit.t[0] ;
 wire \vgadonut.donut.donuthit.t[10] ;
 wire \vgadonut.donut.donuthit.t[11] ;
 wire \vgadonut.donut.donuthit.t[12] ;
 wire \vgadonut.donut.donuthit.t[13] ;
 wire \vgadonut.donut.donuthit.t[14] ;
 wire \vgadonut.donut.donuthit.t[15] ;
 wire \vgadonut.donut.donuthit.t[1] ;
 wire \vgadonut.donut.donuthit.t[2] ;
 wire \vgadonut.donut.donuthit.t[3] ;
 wire \vgadonut.donut.donuthit.t[4] ;
 wire \vgadonut.donut.donuthit.t[5] ;
 wire \vgadonut.donut.donuthit.t[6] ;
 wire \vgadonut.donut.donuthit.t[7] ;
 wire \vgadonut.donut.donuthit.t[8] ;
 wire \vgadonut.donut.donuthit.t[9] ;
 wire \vgadonut.donut.frame ;
 wire \vgadonut.donut.h_count[0] ;
 wire \vgadonut.donut.h_count[10] ;
 wire \vgadonut.donut.h_count[1] ;
 wire \vgadonut.donut.h_count[2] ;
 wire \vgadonut.donut.h_count[3] ;
 wire \vgadonut.donut.h_count[4] ;
 wire \vgadonut.donut.h_count[5] ;
 wire \vgadonut.donut.h_count[6] ;
 wire \vgadonut.donut.h_count[7] ;
 wire \vgadonut.donut.h_count[8] ;
 wire \vgadonut.donut.h_count[9] ;
 wire \vgadonut.donut.rx6[0] ;
 wire \vgadonut.donut.rx6[1] ;
 wire \vgadonut.donut.rx6[2] ;
 wire \vgadonut.donut.rx6[3] ;
 wire \vgadonut.donut.rx6[4] ;
 wire \vgadonut.donut.rx6[5] ;
 wire \vgadonut.donut.ry6[0] ;
 wire \vgadonut.donut.ry6[1] ;
 wire \vgadonut.donut.ry6[2] ;
 wire \vgadonut.donut.ry6[3] ;
 wire \vgadonut.donut.ry6[4] ;
 wire \vgadonut.donut.ry6[5] ;
 wire \vgadonut.donut.rz6[0] ;
 wire \vgadonut.donut.rz6[1] ;
 wire \vgadonut.donut.rz6[2] ;
 wire \vgadonut.donut.rz6[3] ;
 wire \vgadonut.donut.rz6[4] ;
 wire \vgadonut.donut.rz6[5] ;
 wire \vgadonut.donut.sA[0] ;
 wire \vgadonut.donut.sA[10] ;
 wire \vgadonut.donut.sA[11] ;
 wire \vgadonut.donut.sA[12] ;
 wire \vgadonut.donut.sA[13] ;
 wire \vgadonut.donut.sA[14] ;
 wire \vgadonut.donut.sA[15] ;
 wire \vgadonut.donut.sA[1] ;
 wire \vgadonut.donut.sA[2] ;
 wire \vgadonut.donut.sA[3] ;
 wire \vgadonut.donut.sA[4] ;
 wire \vgadonut.donut.sA[5] ;
 wire \vgadonut.donut.sA[6] ;
 wire \vgadonut.donut.sA[7] ;
 wire \vgadonut.donut.sA[8] ;
 wire \vgadonut.donut.sA[9] ;
 wire \vgadonut.donut.sAcB[0] ;
 wire \vgadonut.donut.sAcB[10] ;
 wire \vgadonut.donut.sAcB[11] ;
 wire \vgadonut.donut.sAcB[12] ;
 wire \vgadonut.donut.sAcB[13] ;
 wire \vgadonut.donut.sAcB[14] ;
 wire \vgadonut.donut.sAcB[15] ;
 wire \vgadonut.donut.sAcB[1] ;
 wire \vgadonut.donut.sAcB[2] ;
 wire \vgadonut.donut.sAcB[3] ;
 wire \vgadonut.donut.sAcB[4] ;
 wire \vgadonut.donut.sAcB[5] ;
 wire \vgadonut.donut.sAcB[6] ;
 wire \vgadonut.donut.sAcB[7] ;
 wire \vgadonut.donut.sAcB[8] ;
 wire \vgadonut.donut.sAcB[9] ;
 wire \vgadonut.donut.sAsB[0] ;
 wire \vgadonut.donut.sAsB[10] ;
 wire \vgadonut.donut.sAsB[11] ;
 wire \vgadonut.donut.sAsB[12] ;
 wire \vgadonut.donut.sAsB[13] ;
 wire \vgadonut.donut.sAsB[14] ;
 wire \vgadonut.donut.sAsB[15] ;
 wire \vgadonut.donut.sAsB[1] ;
 wire \vgadonut.donut.sAsB[2] ;
 wire \vgadonut.donut.sAsB[3] ;
 wire \vgadonut.donut.sAsB[4] ;
 wire \vgadonut.donut.sAsB[5] ;
 wire \vgadonut.donut.sAsB[6] ;
 wire \vgadonut.donut.sAsB[7] ;
 wire \vgadonut.donut.sAsB[8] ;
 wire \vgadonut.donut.sAsB[9] ;
 wire \vgadonut.donut.sB[0] ;
 wire \vgadonut.donut.sB[1] ;
 wire \vgadonut.donut.v_count[2] ;
 wire \vgadonut.donut.v_count[3] ;
 wire \vgadonut.donut.v_count[4] ;
 wire \vgadonut.donut.v_count[5] ;
 wire \vgadonut.donut.v_count[6] ;
 wire \vgadonut.donut.v_count[7] ;
 wire \vgadonut.donut.v_count[8] ;
 wire \vgadonut.donut.v_count[9] ;
 wire \vgadonut.donut.ycA[0] ;
 wire \vgadonut.donut.ycA[10] ;
 wire \vgadonut.donut.ycA[11] ;
 wire \vgadonut.donut.ycA[12] ;
 wire \vgadonut.donut.ycA[13] ;
 wire \vgadonut.donut.ycA[14] ;
 wire \vgadonut.donut.ycA[15] ;
 wire \vgadonut.donut.ycA[16] ;
 wire \vgadonut.donut.ycA[17] ;
 wire \vgadonut.donut.ycA[18] ;
 wire \vgadonut.donut.ycA[19] ;
 wire \vgadonut.donut.ycA[1] ;
 wire \vgadonut.donut.ycA[20] ;
 wire \vgadonut.donut.ycA[21] ;
 wire \vgadonut.donut.ycA[2] ;
 wire \vgadonut.donut.ycA[3] ;
 wire \vgadonut.donut.ycA[4] ;
 wire \vgadonut.donut.ycA[5] ;
 wire \vgadonut.donut.ycA[6] ;
 wire \vgadonut.donut.ycA[7] ;
 wire \vgadonut.donut.ycA[8] ;
 wire \vgadonut.donut.ycA[9] ;
 wire \vgadonut.donut.ysA[0] ;
 wire \vgadonut.donut.ysA[10] ;
 wire \vgadonut.donut.ysA[11] ;
 wire \vgadonut.donut.ysA[12] ;
 wire \vgadonut.donut.ysA[13] ;
 wire \vgadonut.donut.ysA[14] ;
 wire \vgadonut.donut.ysA[15] ;
 wire \vgadonut.donut.ysA[16] ;
 wire \vgadonut.donut.ysA[17] ;
 wire \vgadonut.donut.ysA[18] ;
 wire \vgadonut.donut.ysA[19] ;
 wire \vgadonut.donut.ysA[1] ;
 wire \vgadonut.donut.ysA[20] ;
 wire \vgadonut.donut.ysA[21] ;
 wire \vgadonut.donut.ysA[2] ;
 wire \vgadonut.donut.ysA[3] ;
 wire \vgadonut.donut.ysA[4] ;
 wire \vgadonut.donut.ysA[5] ;
 wire \vgadonut.donut.ysA[6] ;
 wire \vgadonut.donut.ysA[7] ;
 wire \vgadonut.donut.ysA[8] ;
 wire \vgadonut.donut.ysA[9] ;
 wire \vgadonut.frame[1] ;
 wire \vgadonut.frame[2] ;
 wire \vgadonut.frame[3] ;
 wire \vgadonut.frame[4] ;
 wire \vgadonut.frame[5] ;
 wire \vgadonut.frame[6] ;
 wire \vgadonut.frame[7] ;
 wire \vgadonut.vsync ;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;

 sg13g2_inv_1 _07444_ (.Y(_06847_),
    .A(net1914));
 sg13g2_inv_1 _07445_ (.Y(_06848_),
    .A(\vgadonut.donut.v_count[5] ));
 sg13g2_inv_1 _07446_ (.Y(_06849_),
    .A(net2235));
 sg13g2_inv_1 _07447_ (.Y(_06850_),
    .A(net2177));
 sg13g2_inv_1 _07448_ (.Y(_06851_),
    .A(\vgadonut.donut.ysA[4] ));
 sg13g2_inv_1 _07449_ (.Y(_06852_),
    .A(net2106));
 sg13g2_inv_1 _07450_ (.Y(_06853_),
    .A(net1908));
 sg13g2_inv_1 _07451_ (.Y(_06854_),
    .A(net2210));
 sg13g2_inv_1 _07452_ (.Y(_06855_),
    .A(net2107));
 sg13g2_inv_1 _07453_ (.Y(_06856_),
    .A(net1907));
 sg13g2_inv_1 _07454_ (.Y(_06857_),
    .A(net2086));
 sg13g2_inv_1 _07455_ (.Y(_06858_),
    .A(net2066));
 sg13g2_inv_1 _07456_ (.Y(_06859_),
    .A(\vgadonut.donut.cAsB[7] ));
 sg13g2_inv_1 _07457_ (.Y(_06860_),
    .A(\vgadonut.donut.cAcB[2] ));
 sg13g2_inv_1 _07458_ (.Y(_06861_),
    .A(net2174));
 sg13g2_inv_1 _07459_ (.Y(_06862_),
    .A(net2085));
 sg13g2_inv_1 _07460_ (.Y(_06863_),
    .A(net2188));
 sg13g2_inv_1 _07461_ (.Y(_06864_),
    .A(net2118));
 sg13g2_inv_1 _07462_ (.Y(_06865_),
    .A(net1902));
 sg13g2_inv_1 _07463_ (.Y(_06866_),
    .A(net2178));
 sg13g2_inv_1 _07464_ (.Y(_06867_),
    .A(net2264));
 sg13g2_inv_1 _07465_ (.Y(_06868_),
    .A(net2310));
 sg13g2_inv_1 _07466_ (.Y(_06869_),
    .A(net1950));
 sg13g2_inv_1 _07467_ (.Y(_06870_),
    .A(\vgadonut.donut.ysA[13] ));
 sg13g2_inv_1 _07468_ (.Y(_06871_),
    .A(net2152));
 sg13g2_inv_1 _07469_ (.Y(_06872_),
    .A(net2245));
 sg13g2_inv_1 _07470_ (.Y(_06873_),
    .A(net1947));
 sg13g2_inv_1 _07471_ (.Y(_06874_),
    .A(net2165));
 sg13g2_inv_1 _07472_ (.Y(_06875_),
    .A(net1895));
 sg13g2_inv_2 _07473_ (.Y(_06876_),
    .A(net2179));
 sg13g2_inv_1 _07474_ (.Y(_06877_),
    .A(net1943));
 sg13g2_inv_2 _07475_ (.Y(_06878_),
    .A(net2173));
 sg13g2_inv_1 _07476_ (.Y(_06879_),
    .A(net2140));
 sg13g2_inv_1 _07477_ (.Y(_06880_),
    .A(net2170));
 sg13g2_inv_2 _07478_ (.Y(_06881_),
    .A(net2151));
 sg13g2_inv_1 _07479_ (.Y(_06882_),
    .A(net2319));
 sg13g2_inv_1 _07480_ (.Y(_06883_),
    .A(net2091));
 sg13g2_inv_1 _07481_ (.Y(_06884_),
    .A(net2064));
 sg13g2_inv_1 _07482_ (.Y(_06885_),
    .A(net2031));
 sg13g2_inv_1 _07483_ (.Y(_06886_),
    .A(\vgadonut.donut.sAsB[3] ));
 sg13g2_inv_1 _07484_ (.Y(_06887_),
    .A(net2001));
 sg13g2_inv_2 _07485_ (.Y(_06888_),
    .A(net2263));
 sg13g2_inv_1 _07486_ (.Y(_06889_),
    .A(net2238));
 sg13g2_inv_1 _07487_ (.Y(_06890_),
    .A(net2109));
 sg13g2_inv_1 _07488_ (.Y(_06891_),
    .A(net2080));
 sg13g2_inv_1 _07489_ (.Y(_06892_),
    .A(\vgadonut.donut.ycA[7] ));
 sg13g2_inv_1 _07490_ (.Y(_06893_),
    .A(\vgadonut.donut.sAsB[7] ));
 sg13g2_inv_1 _07491_ (.Y(_06894_),
    .A(net2065));
 sg13g2_inv_1 _07492_ (.Y(_06895_),
    .A(\vgadonut.donut.ycA[8] ));
 sg13g2_inv_2 _07493_ (.Y(_06896_),
    .A(\vgadonut.donut.sAsB[8] ));
 sg13g2_inv_1 _07494_ (.Y(_06897_),
    .A(net2040));
 sg13g2_inv_2 _07495_ (.Y(_06898_),
    .A(\vgadonut.donut.sAcB[3] ));
 sg13g2_inv_1 _07496_ (.Y(_06899_),
    .A(net2247));
 sg13g2_inv_2 _07497_ (.Y(_06900_),
    .A(\vgadonut.donut.sAsB[9] ));
 sg13g2_inv_1 _07498_ (.Y(_06901_),
    .A(net2048));
 sg13g2_inv_1 _07499_ (.Y(_06902_),
    .A(\vgadonut.donut.ycA[10] ));
 sg13g2_inv_4 _07500_ (.A(\vgadonut.donut.sAsB[10] ),
    .Y(_06903_));
 sg13g2_inv_1 _07501_ (.Y(_06904_),
    .A(net2079));
 sg13g2_inv_1 _07502_ (.Y(_06905_),
    .A(net2277));
 sg13g2_inv_2 _07503_ (.Y(_06906_),
    .A(net2338));
 sg13g2_inv_1 _07504_ (.Y(_06907_),
    .A(net2041));
 sg13g2_inv_1 _07505_ (.Y(_06908_),
    .A(\vgadonut.donut.sAsB[13] ));
 sg13g2_inv_1 _07506_ (.Y(_06909_),
    .A(_00110_));
 sg13g2_inv_2 _07507_ (.Y(_06910_),
    .A(net1929));
 sg13g2_inv_1 _07508_ (.Y(_06911_),
    .A(net2133));
 sg13g2_inv_1 _07509_ (.Y(_06912_),
    .A(net2327));
 sg13g2_inv_1 _07510_ (.Y(_06913_),
    .A(net1928));
 sg13g2_inv_1 _07511_ (.Y(_06914_),
    .A(net2150));
 sg13g2_inv_4 _07512_ (.A(net1886),
    .Y(_00546_));
 sg13g2_inv_1 _07513_ (.Y(_00547_),
    .A(net2187));
 sg13g2_inv_1 _07514_ (.Y(_00548_),
    .A(net1926));
 sg13g2_inv_1 _07515_ (.Y(_00549_),
    .A(net2274));
 sg13g2_inv_1 _07516_ (.Y(_00550_),
    .A(net2234));
 sg13g2_inv_2 _07517_ (.Y(_00551_),
    .A(net2020));
 sg13g2_inv_1 _07518_ (.Y(_00552_),
    .A(net2209));
 sg13g2_inv_2 _07519_ (.Y(_00553_),
    .A(net1919));
 sg13g2_inv_1 _07520_ (.Y(_00554_),
    .A(net2096));
 sg13g2_inv_1 _07521_ (.Y(_00555_),
    .A(net2227));
 sg13g2_inv_1 _07522_ (.Y(_00556_),
    .A(net2345));
 sg13g2_inv_1 _07523_ (.Y(_00557_),
    .A(net1916));
 sg13g2_inv_1 _07524_ (.Y(_00558_),
    .A(net2032));
 sg13g2_inv_2 _07525_ (.Y(_00559_),
    .A(net2215));
 sg13g2_inv_1 _07526_ (.Y(_00560_),
    .A(net2011));
 sg13g2_inv_1 _07527_ (.Y(_00561_),
    .A(net1863));
 sg13g2_inv_1 _07528_ (.Y(_00562_),
    .A(net2098));
 sg13g2_inv_1 _07529_ (.Y(_00563_),
    .A(\vgadonut.donut.cB[5] ));
 sg13g2_inv_1 _07530_ (.Y(_00564_),
    .A(net2043));
 sg13g2_inv_1 _07531_ (.Y(_00565_),
    .A(net2084));
 sg13g2_inv_1 _07532_ (.Y(_00566_),
    .A(\vgadonut.donut.cB[7] ));
 sg13g2_inv_1 _07533_ (.Y(_00567_),
    .A(net2095));
 sg13g2_inv_1 _07534_ (.Y(_00568_),
    .A(\vgadonut.donut.cB[8] ));
 sg13g2_inv_1 _07535_ (.Y(_00569_),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[1] ));
 sg13g2_inv_1 _07536_ (.Y(_00570_),
    .A(net2099));
 sg13g2_inv_1 _07537_ (.Y(_00571_),
    .A(net2058));
 sg13g2_inv_1 _07538_ (.Y(_00572_),
    .A(\vgadonut.donut.cB[10] ));
 sg13g2_inv_2 _07539_ (.Y(_00573_),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[3] ));
 sg13g2_inv_1 _07540_ (.Y(_00574_),
    .A(net2332));
 sg13g2_inv_2 _07541_ (.Y(_00575_),
    .A(net2104));
 sg13g2_inv_1 _07542_ (.Y(_00576_),
    .A(\vgadonut.donut.cB[12] ));
 sg13g2_inv_2 _07543_ (.Y(_00577_),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[5] ));
 sg13g2_inv_1 _07544_ (.Y(_00578_),
    .A(net2299));
 sg13g2_inv_1 _07545_ (.Y(_00579_),
    .A(net1882));
 sg13g2_inv_1 _07546_ (.Y(_00580_),
    .A(net2244));
 sg13g2_inv_1 _07547_ (.Y(_00581_),
    .A(net2271));
 sg13g2_inv_2 _07548_ (.Y(_00582_),
    .A(net1859));
 sg13g2_inv_2 _07549_ (.Y(_00583_),
    .A(net2243));
 sg13g2_inv_2 _07550_ (.Y(_00584_),
    .A(net2206));
 sg13g2_inv_1 _07551_ (.Y(_00585_),
    .A(net1877));
 sg13g2_inv_1 _07552_ (.Y(_00586_),
    .A(net2214));
 sg13g2_inv_2 _07553_ (.Y(_00587_),
    .A(net1875));
 sg13g2_inv_1 _07554_ (.Y(_00588_),
    .A(net2308));
 sg13g2_inv_1 _07555_ (.Y(_00589_),
    .A(net1873));
 sg13g2_inv_1 _07556_ (.Y(_00590_),
    .A(net2192));
 sg13g2_inv_1 _07557_ (.Y(_00591_),
    .A(net2273));
 sg13g2_inv_1 _07558_ (.Y(_00592_),
    .A(net1870));
 sg13g2_inv_1 _07559_ (.Y(_00593_),
    .A(net2297));
 sg13g2_inv_2 _07560_ (.Y(_00594_),
    .A(net1846));
 sg13g2_inv_1 _07561_ (.Y(_00595_),
    .A(net1842));
 sg13g2_inv_1 _07562_ (.Y(_00596_),
    .A(net1840));
 sg13g2_inv_2 _07563_ (.Y(_00597_),
    .A(net1833));
 sg13g2_inv_1 _07564_ (.Y(_00598_),
    .A(net1831));
 sg13g2_inv_1 _07565_ (.Y(_00599_),
    .A(net1829));
 sg13g2_inv_2 _07566_ (.Y(_00600_),
    .A(\vgadonut.donut.cA[6] ));
 sg13g2_inv_2 _07567_ (.Y(_00601_),
    .A(\vgadonut.donut.cA[5] ));
 sg13g2_inv_1 _07568_ (.Y(_00602_),
    .A(\vgadonut.donut.cA[4] ));
 sg13g2_inv_1 _07569_ (.Y(_00603_),
    .A(\vgadonut.donut.cA[3] ));
 sg13g2_inv_2 _07570_ (.Y(_00604_),
    .A(\vgadonut.donut.cA[7] ));
 sg13g2_inv_2 _07571_ (.Y(_00605_),
    .A(\vgadonut.donut.cA[9] ));
 sg13g2_inv_2 _07572_ (.Y(_00606_),
    .A(net1821));
 sg13g2_inv_1 _07573_ (.Y(_00607_),
    .A(net1813));
 sg13g2_inv_1 _07574_ (.Y(_00608_),
    .A(_00126_));
 sg13g2_inv_1 _07575_ (.Y(_00609_),
    .A(_00128_));
 sg13g2_inv_1 _07576_ (.Y(_00610_),
    .A(_00129_));
 sg13g2_inv_1 _07577_ (.Y(_00611_),
    .A(_00131_));
 sg13g2_inv_1 _07578_ (.Y(_00612_),
    .A(_00132_));
 sg13g2_inv_1 _07579_ (.Y(_00613_),
    .A(_00133_));
 sg13g2_inv_1 _07580_ (.Y(_00614_),
    .A(_00134_));
 sg13g2_inv_1 _07581_ (.Y(_00615_),
    .A(_00135_));
 sg13g2_inv_1 _07582_ (.Y(_00616_),
    .A(_00136_));
 sg13g2_inv_1 _07583_ (.Y(_00617_),
    .A(_00138_));
 sg13g2_inv_1 _07584_ (.Y(_00618_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[13] ));
 sg13g2_inv_1 _07585_ (.Y(_00619_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[12] ));
 sg13g2_inv_1 _07586_ (.Y(_00620_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[12] ));
 sg13g2_inv_1 _07587_ (.Y(_00621_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[9] ));
 sg13g2_inv_1 _07588_ (.Y(_00622_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[7] ));
 sg13g2_inv_2 _07589_ (.Y(_00623_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[6] ));
 sg13g2_inv_1 _07590_ (.Y(_00624_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[2] ));
 sg13g2_inv_1 _07591_ (.Y(_00625_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[0] ));
 sg13g2_inv_1 _07592_ (.Y(_00626_),
    .A(_00143_));
 sg13g2_inv_2 _07593_ (.Y(_00627_),
    .A(_00144_));
 sg13g2_inv_1 _07594_ (.Y(_00628_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[9] ));
 sg13g2_inv_1 _07595_ (.Y(_00629_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[7] ));
 sg13g2_inv_1 _07596_ (.Y(_00630_),
    .A(_00148_));
 sg13g2_inv_1 _07597_ (.Y(_00631_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[4] ));
 sg13g2_inv_1 _07598_ (.Y(_00632_),
    .A(_00150_));
 sg13g2_inv_1 _07599_ (.Y(_00633_),
    .A(_00152_));
 sg13g2_inv_1 _07600_ (.Y(_00634_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[1] ));
 sg13g2_inv_1 _07601_ (.Y(_00635_),
    .A(_00153_));
 sg13g2_inv_2 _07602_ (.Y(_00636_),
    .A(_00157_));
 sg13g2_inv_1 _07603_ (.Y(_00637_),
    .A(_00165_));
 sg13g2_inv_1 _07604_ (.Y(_00638_),
    .A(net2307));
 sg13g2_inv_1 _07605_ (.Y(_00639_),
    .A(net2325));
 sg13g2_inv_1 _07606_ (.Y(_00640_),
    .A(net2252));
 sg13g2_inv_1 _07607_ (.Y(_00641_),
    .A(\vgadonut.donut.donuthit.t[3] ));
 sg13g2_inv_1 _07608_ (.Y(_00642_),
    .A(\vgadonut.donut.donuthit.t[9] ));
 sg13g2_inv_1 _07609_ (.Y(_00643_),
    .A(\vgadonut.donut.donuthit.t[12] ));
 sg13g2_inv_1 _07610_ (.Y(_00644_),
    .A(net2358));
 sg13g2_inv_2 _07611_ (.Y(_00645_),
    .A(net1857));
 sg13g2_inv_1 _07612_ (.Y(_00646_),
    .A(\vgadonut.frame[6] ));
 sg13g2_inv_1 _07613_ (.Y(_00647_),
    .A(net2082));
 sg13g2_nand2_1 _07614_ (.Y(_00648_),
    .A(\vgadonut.donut.h_count[3] ),
    .B(net1800));
 sg13g2_and2_1 _07615_ (.A(net1801),
    .B(\vgadonut.donut.h_count[3] ),
    .X(_00649_));
 sg13g2_nand4_1 _07616_ (.B(net1800),
    .C(\vgadonut.donut.h_count[7] ),
    .A(\vgadonut.donut.h_count[5] ),
    .Y(_00650_),
    .D(_00649_));
 sg13g2_nand2_1 _07617_ (.Y(_00651_),
    .A(net2076),
    .B(net2159));
 sg13g2_nor2_1 _07618_ (.A(\vgadonut.donut.h_count[9] ),
    .B(\vgadonut.donut.h_count[8] ),
    .Y(_00652_));
 sg13g2_nand3_1 _07619_ (.B(_00651_),
    .C(_00652_),
    .A(_00650_),
    .Y(_00653_));
 sg13g2_nand2_1 _07620_ (.Y(_00654_),
    .A(\vgadonut.donut.h_count[10] ),
    .B(_00653_));
 sg13g2_xnor2_1 _07621_ (.Y(_00655_),
    .A(\vgadonut.donut.frame ),
    .B(net1915));
 sg13g2_xnor2_1 _07622_ (.Y(_00656_),
    .A(_00178_),
    .B(_00655_));
 sg13g2_xor2_1 _07623_ (.B(net1802),
    .A(net1799),
    .X(_00657_));
 sg13g2_xnor2_1 _07624_ (.Y(_00658_),
    .A(net1799),
    .B(\vgadonut.donut.h_count[1] ));
 sg13g2_xnor2_1 _07625_ (.Y(_00659_),
    .A(\vgadonut.bayer_j[1] ),
    .B(_00657_));
 sg13g2_xor2_1 _07626_ (.B(net1915),
    .A(\vgadonut.donut.h_count[2] ),
    .X(_00660_));
 sg13g2_nor2_1 _07627_ (.A(\vgadonut.donut.h_count[0] ),
    .B(_00660_),
    .Y(_00661_));
 sg13g2_and4_1 _07628_ (.A(_00654_),
    .B(_00656_),
    .C(_00659_),
    .D(_00661_),
    .X(_00662_));
 sg13g2_nand4_1 _07629_ (.B(_00656_),
    .C(_00659_),
    .A(_00654_),
    .Y(_00663_),
    .D(_00661_));
 sg13g2_nand2_1 _07630_ (.Y(_00664_),
    .A(net1984),
    .B(net1689));
 sg13g2_nand2b_1 _07631_ (.Y(_00665_),
    .B(net1671),
    .A_N(\vgadonut.donut.donut_luma[4] ));
 sg13g2_o21ai_1 _07632_ (.B1(_00665_),
    .Y(_00666_),
    .A1(\vgadonut.donut.donuthit.light[12] ),
    .A2(net1671));
 sg13g2_inv_1 _07633_ (.Y(_00292_),
    .A(_00666_));
 sg13g2_nand2b_1 _07634_ (.Y(_00667_),
    .B(net1671),
    .A_N(\vgadonut.donut.donut_luma[2] ));
 sg13g2_o21ai_1 _07635_ (.B1(_00667_),
    .Y(_00668_),
    .A1(\vgadonut.donut.donuthit.light[10] ),
    .A2(net1672));
 sg13g2_inv_1 _07636_ (.Y(_00290_),
    .A(_00668_));
 sg13g2_mux2_1 _07637_ (.A0(net2007),
    .A1(\vgadonut.donut.donut_luma[0] ),
    .S(net1672),
    .X(_00288_));
 sg13g2_and2_2 _07638_ (.A(net1635),
    .B(net1647),
    .X(_00669_));
 sg13g2_nand2_2 _07639_ (.Y(_00670_),
    .A(net1635),
    .B(net1647));
 sg13g2_nor2_2 _07640_ (.A(net1635),
    .B(net1647),
    .Y(_00671_));
 sg13g2_or2_1 _07641_ (.X(_00672_),
    .B(_00671_),
    .A(_00669_));
 sg13g2_nand2b_1 _07642_ (.Y(_00673_),
    .B(net1672),
    .A_N(\vgadonut.donut.donut_luma[3] ));
 sg13g2_o21ai_1 _07643_ (.B1(_00673_),
    .Y(_00674_),
    .A1(net2154),
    .A2(net1672));
 sg13g2_inv_1 _07644_ (.Y(_00291_),
    .A(net2155));
 sg13g2_nand2_1 _07645_ (.Y(_00675_),
    .A(net1615),
    .B(net1645));
 sg13g2_nand2b_1 _07646_ (.Y(_00676_),
    .B(net1671),
    .A_N(\vgadonut.donut.donut_luma[1] ));
 sg13g2_o21ai_1 _07647_ (.B1(_00676_),
    .Y(_00677_),
    .A1(\vgadonut.donut.donuthit.light[9] ),
    .A2(net1671));
 sg13g2_inv_2 _07648_ (.Y(_00289_),
    .A(_00677_));
 sg13g2_nor2_1 _07649_ (.A(net1633),
    .B(_00677_),
    .Y(_00678_));
 sg13g2_o21ai_1 _07650_ (.B1(_00675_),
    .Y(_00679_),
    .A1(_00671_),
    .A2(_00678_));
 sg13g2_nand2b_1 _07651_ (.Y(_00680_),
    .B(net1671),
    .A_N(\vgadonut.donut.donut_luma[5] ));
 sg13g2_o21ai_1 _07652_ (.B1(_00680_),
    .Y(_00681_),
    .A1(net2335),
    .A2(net1671));
 sg13g2_inv_1 _07653_ (.Y(_00293_),
    .A(_00681_));
 sg13g2_nor2_2 _07654_ (.A(net1636),
    .B(_00289_),
    .Y(_00682_));
 sg13g2_nand2_1 _07655_ (.Y(_00683_),
    .A(_00668_),
    .B(_00677_));
 sg13g2_nor2_1 _07656_ (.A(net1647),
    .B(_00289_),
    .Y(_00684_));
 sg13g2_nand2_1 _07657_ (.Y(_00685_),
    .A(_00668_),
    .B(_00684_));
 sg13g2_nor2_1 _07658_ (.A(net1634),
    .B(_00685_),
    .Y(_00686_));
 sg13g2_nor2_1 _07659_ (.A(net1637),
    .B(net1642),
    .Y(_00687_));
 sg13g2_nand2_2 _07660_ (.Y(_00688_),
    .A(net1646),
    .B(net1630));
 sg13g2_o21ai_1 _07661_ (.B1(net1629),
    .Y(_00689_),
    .A1(net1646),
    .A2(_00686_));
 sg13g2_a21oi_1 _07662_ (.A1(net1646),
    .A2(_00679_),
    .Y(_00690_),
    .B1(_00689_));
 sg13g2_nor2_2 _07663_ (.A(net1646),
    .B(net1629),
    .Y(_00691_));
 sg13g2_nor2_2 _07664_ (.A(_00668_),
    .B(_00677_),
    .Y(_00692_));
 sg13g2_nand2_2 _07665_ (.Y(_00693_),
    .A(net1635),
    .B(_00289_));
 sg13g2_nand2_2 _07666_ (.Y(_00694_),
    .A(_00669_),
    .B(_00289_));
 sg13g2_nor2_2 _07667_ (.A(_00671_),
    .B(_00682_),
    .Y(_00695_));
 sg13g2_and2_1 _07668_ (.A(_00694_),
    .B(_00695_),
    .X(_00696_));
 sg13g2_nor2_1 _07669_ (.A(net1639),
    .B(net1635),
    .Y(_00697_));
 sg13g2_nor2_1 _07670_ (.A(net1643),
    .B(_00693_),
    .Y(_00698_));
 sg13g2_nand2_1 _07671_ (.Y(_00699_),
    .A(net1633),
    .B(_00692_));
 sg13g2_nand2_1 _07672_ (.Y(_00700_),
    .A(_00691_),
    .B(_00698_));
 sg13g2_nand2_1 _07673_ (.Y(_00701_),
    .A(_00696_),
    .B(_00699_));
 sg13g2_a221oi_1 _07674_ (.B2(_00691_),
    .C1(_00690_),
    .B1(_00701_),
    .A1(net2336),
    .Y(_00000_),
    .A2(_00697_));
 sg13g2_nand2_1 _07675_ (.Y(_00702_),
    .A(net1637),
    .B(_00699_));
 sg13g2_a21oi_1 _07676_ (.A1(net1643),
    .A2(_00694_),
    .Y(_00703_),
    .B1(_00702_));
 sg13g2_nor2_2 _07677_ (.A(net1637),
    .B(net1644),
    .Y(_00704_));
 sg13g2_nor3_1 _07678_ (.A(net1629),
    .B(_00703_),
    .C(_00704_),
    .Y(_00705_));
 sg13g2_nand2_1 _07679_ (.Y(_00706_),
    .A(net1645),
    .B(_00695_));
 sg13g2_nand2_1 _07680_ (.Y(_00707_),
    .A(net1643),
    .B(_00693_));
 sg13g2_nor2_1 _07681_ (.A(_00692_),
    .B(_00706_),
    .Y(_00708_));
 sg13g2_nor2_2 _07682_ (.A(net1636),
    .B(_00677_),
    .Y(_00709_));
 sg13g2_nor3_1 _07683_ (.A(_00669_),
    .B(net1643),
    .C(_00709_),
    .Y(_00710_));
 sg13g2_nor3_1 _07684_ (.A(_00688_),
    .B(_00708_),
    .C(_00710_),
    .Y(_00711_));
 sg13g2_nor2_1 _07685_ (.A(net1646),
    .B(net1642),
    .Y(_00712_));
 sg13g2_nand2b_2 _07686_ (.Y(_00713_),
    .B(_00289_),
    .A_N(net1647));
 sg13g2_and4_1 _07687_ (.A(net1615),
    .B(net1643),
    .C(_00712_),
    .D(_00713_),
    .X(_00714_));
 sg13g2_nor3_1 _07688_ (.A(_00705_),
    .B(_00711_),
    .C(_00714_),
    .Y(_00001_));
 sg13g2_nand3_1 _07689_ (.B(_00712_),
    .C(_00713_),
    .A(_00668_),
    .Y(_00715_));
 sg13g2_a22oi_1 _07690_ (.Y(_00716_),
    .B1(_00707_),
    .B2(net1629),
    .A2(_00699_),
    .A1(_00691_));
 sg13g2_nand2_2 _07691_ (.Y(_00717_),
    .A(net1647),
    .B(_00677_));
 sg13g2_nand2_1 _07692_ (.Y(_00718_),
    .A(_00713_),
    .B(_00717_));
 sg13g2_nor2_1 _07693_ (.A(_00668_),
    .B(_00718_),
    .Y(_00719_));
 sg13g2_nor2_1 _07694_ (.A(_00709_),
    .B(_00719_),
    .Y(_00720_));
 sg13g2_nor2_1 _07695_ (.A(net1643),
    .B(_00720_),
    .Y(_00721_));
 sg13g2_a22oi_1 _07696_ (.Y(_00002_),
    .B1(_00721_),
    .B2(_00687_),
    .A2(_00716_),
    .A1(_00715_));
 sg13g2_nor3_1 _07697_ (.A(net1646),
    .B(net1632),
    .C(_00719_),
    .Y(_00722_));
 sg13g2_a21oi_1 _07698_ (.A1(_00694_),
    .A2(_00704_),
    .Y(_00723_),
    .B1(_00722_));
 sg13g2_o21ai_1 _07699_ (.B1(net1629),
    .Y(_00724_),
    .A1(_00682_),
    .A2(_00723_));
 sg13g2_nand2_1 _07700_ (.Y(_00003_),
    .A(_00700_),
    .B(_00724_));
 sg13g2_nor3_1 _07701_ (.A(net1615),
    .B(net1644),
    .C(_00709_),
    .Y(_00725_));
 sg13g2_a21o_1 _07702_ (.A2(net1644),
    .A1(net1615),
    .B1(_00725_),
    .X(_00726_));
 sg13g2_nor2_1 _07703_ (.A(net1638),
    .B(net1632),
    .Y(_00727_));
 sg13g2_nand2_1 _07704_ (.Y(_00728_),
    .A(_00717_),
    .B(_00727_));
 sg13g2_a21oi_1 _07705_ (.A1(_00668_),
    .A2(_00713_),
    .Y(_00729_),
    .B1(_00728_));
 sg13g2_nor2_1 _07706_ (.A(net1615),
    .B(_00684_),
    .Y(_00730_));
 sg13g2_a221oi_1 _07707_ (.B2(_00704_),
    .C1(_00729_),
    .B1(_00730_),
    .A1(net1638),
    .Y(_00731_),
    .A2(_00726_));
 sg13g2_o21ai_1 _07708_ (.B1(_00712_),
    .Y(_00732_),
    .A1(net1632),
    .A2(_00683_));
 sg13g2_inv_1 _07709_ (.Y(_00225_),
    .A(_00732_));
 sg13g2_nor2_2 _07710_ (.A(net1644),
    .B(_00682_),
    .Y(_00733_));
 sg13g2_nand2_1 _07711_ (.Y(_00734_),
    .A(net1632),
    .B(_00683_));
 sg13g2_a22oi_1 _07712_ (.Y(_00735_),
    .B1(_00733_),
    .B2(_00670_),
    .A2(_00730_),
    .A1(net1643));
 sg13g2_a21oi_1 _07713_ (.A1(_00687_),
    .A2(_00735_),
    .Y(_00736_),
    .B1(_00225_));
 sg13g2_o21ai_1 _07714_ (.B1(_00736_),
    .Y(_00004_),
    .A1(net1629),
    .A2(_00731_));
 sg13g2_nor3_1 _07715_ (.A(_00672_),
    .B(net1632),
    .C(_00720_),
    .Y(_00737_));
 sg13g2_o21ai_1 _07716_ (.B1(_00720_),
    .Y(_00738_),
    .A1(_00672_),
    .A2(net1632));
 sg13g2_nand2_1 _07717_ (.Y(_00739_),
    .A(net1638),
    .B(_00738_));
 sg13g2_nor2_1 _07718_ (.A(_00669_),
    .B(_00707_),
    .Y(_00740_));
 sg13g2_nand3_1 _07719_ (.B(net1643),
    .C(_00693_),
    .A(_00670_),
    .Y(_00741_));
 sg13g2_nor2_1 _07720_ (.A(net1638),
    .B(_00741_),
    .Y(_00742_));
 sg13g2_o21ai_1 _07721_ (.B1(_00289_),
    .Y(_00743_),
    .A1(_00668_),
    .A2(net1647));
 sg13g2_a22oi_1 _07722_ (.Y(_00744_),
    .B1(_00743_),
    .B2(_00704_),
    .A2(_00742_),
    .A1(_00695_));
 sg13g2_o21ai_1 _07723_ (.B1(_00744_),
    .Y(_00745_),
    .A1(_00737_),
    .A2(_00739_));
 sg13g2_nand2_1 _07724_ (.Y(_00746_),
    .A(_00670_),
    .B(_00289_));
 sg13g2_nand2_1 _07725_ (.Y(_00747_),
    .A(net1644),
    .B(_00746_));
 sg13g2_o21ai_1 _07726_ (.B1(_00747_),
    .Y(_00748_),
    .A1(_00671_),
    .A2(_00719_));
 sg13g2_nor2_1 _07727_ (.A(net1632),
    .B(_00717_),
    .Y(_00749_));
 sg13g2_nor2_1 _07728_ (.A(_00688_),
    .B(_00749_),
    .Y(_00750_));
 sg13g2_a22oi_1 _07729_ (.Y(_00751_),
    .B1(_00748_),
    .B2(_00750_),
    .A2(_00745_),
    .A1(net1642));
 sg13g2_nand2_1 _07730_ (.Y(_00005_),
    .A(_00732_),
    .B(_00751_));
 sg13g2_a21oi_1 _07731_ (.A1(_00694_),
    .A2(_00733_),
    .Y(_00752_),
    .B1(net1637));
 sg13g2_a21oi_1 _07732_ (.A1(_00741_),
    .A2(_00752_),
    .Y(_00753_),
    .B1(net1630));
 sg13g2_a221oi_1 _07733_ (.B2(_00675_),
    .C1(_00689_),
    .B1(_00746_),
    .A1(net1644),
    .Y(_00754_),
    .A2(_00709_));
 sg13g2_o21ai_1 _07734_ (.B1(net1632),
    .Y(_00755_),
    .A1(_00669_),
    .A2(_00692_));
 sg13g2_nand2_1 _07735_ (.Y(_00756_),
    .A(net1637),
    .B(_00755_));
 sg13g2_inv_1 _07736_ (.Y(_00757_),
    .A(_00756_));
 sg13g2_nand3_1 _07737_ (.B(_00706_),
    .C(_00755_),
    .A(_00691_),
    .Y(_00758_));
 sg13g2_o21ai_1 _07738_ (.B1(_00758_),
    .Y(_00006_),
    .A1(_00753_),
    .A2(_00754_));
 sg13g2_o21ai_1 _07739_ (.B1(net1637),
    .Y(_00759_),
    .A1(net1634),
    .A2(_00695_));
 sg13g2_nand2b_1 _07740_ (.Y(_00760_),
    .B(_00755_),
    .A_N(_00759_));
 sg13g2_o21ai_1 _07741_ (.B1(_00760_),
    .Y(_00761_),
    .A1(net1637),
    .A2(_00733_));
 sg13g2_a21oi_1 _07742_ (.A1(_00693_),
    .A2(_00733_),
    .Y(_00762_),
    .B1(_00688_));
 sg13g2_a22oi_1 _07743_ (.Y(_00007_),
    .B1(_00762_),
    .B2(_00741_),
    .A2(_00761_),
    .A1(net1642));
 sg13g2_o21ai_1 _07744_ (.B1(net1629),
    .Y(_00763_),
    .A1(_00698_),
    .A2(_00740_));
 sg13g2_nand2_1 _07745_ (.Y(_00008_),
    .A(_00759_),
    .B(_00763_));
 sg13g2_a21oi_1 _07746_ (.A1(_00670_),
    .A2(_00713_),
    .Y(_00764_),
    .B1(net1633));
 sg13g2_nor2_1 _07747_ (.A(net1642),
    .B(_00764_),
    .Y(_00765_));
 sg13g2_o21ai_1 _07748_ (.B1(_00765_),
    .Y(_00766_),
    .A1(net1615),
    .A2(_00734_));
 sg13g2_xor2_1 _07749_ (.B(_00733_),
    .A(net1647),
    .X(_00767_));
 sg13g2_a21oi_1 _07750_ (.A1(_00681_),
    .A2(_00767_),
    .Y(_00768_),
    .B1(net1639));
 sg13g2_o21ai_1 _07751_ (.B1(net1644),
    .Y(_00769_),
    .A1(net1615),
    .A2(_00709_));
 sg13g2_nor2b_1 _07752_ (.A(_00725_),
    .B_N(_00691_),
    .Y(_00770_));
 sg13g2_a22oi_1 _07753_ (.Y(_00009_),
    .B1(_00769_),
    .B2(_00770_),
    .A2(_00768_),
    .A1(_00766_));
 sg13g2_a21oi_1 _07754_ (.A1(_00713_),
    .A2(_00717_),
    .Y(_00771_),
    .B1(_00682_));
 sg13g2_a21oi_1 _07755_ (.A1(_00769_),
    .A2(_00771_),
    .Y(_00772_),
    .B1(_00666_));
 sg13g2_o21ai_1 _07756_ (.B1(_00772_),
    .Y(_00773_),
    .A1(_00769_),
    .A2(_00771_));
 sg13g2_a221oi_1 _07757_ (.B2(_00771_),
    .C1(net1631),
    .B1(_00704_),
    .A1(_00666_),
    .Y(_00774_),
    .A2(_00678_));
 sg13g2_a21oi_1 _07758_ (.A1(net1636),
    .A2(net1644),
    .Y(_00775_),
    .B1(_00677_));
 sg13g2_nor3_1 _07759_ (.A(net1615),
    .B(_00688_),
    .C(_00775_),
    .Y(_00776_));
 sg13g2_a21oi_1 _07760_ (.A1(_00773_),
    .A2(_00774_),
    .Y(_00010_),
    .B1(_00776_));
 sg13g2_a21o_1 _07761_ (.A2(_00718_),
    .A1(net1633),
    .B1(net1635),
    .X(_00777_));
 sg13g2_a21o_1 _07762_ (.A2(_00777_),
    .A1(_00693_),
    .B1(_00686_),
    .X(_00778_));
 sg13g2_nor3_1 _07763_ (.A(_00669_),
    .B(_00692_),
    .C(_00734_),
    .Y(_00779_));
 sg13g2_o21ai_1 _07764_ (.B1(net1637),
    .Y(_00780_),
    .A1(_00708_),
    .A2(_00779_));
 sg13g2_a221oi_1 _07765_ (.B2(net1635),
    .C1(net1629),
    .B1(_00727_),
    .A1(_00696_),
    .Y(_00781_),
    .A2(_00704_));
 sg13g2_a22oi_1 _07766_ (.Y(_00011_),
    .B1(_00780_),
    .B2(_00781_),
    .A2(_00778_),
    .A1(_00687_));
 sg13g2_a221oi_1 _07767_ (.B2(_00757_),
    .C1(net1630),
    .B1(_00707_),
    .A1(_00694_),
    .Y(_00782_),
    .A2(_00704_));
 sg13g2_nor2_1 _07768_ (.A(net1635),
    .B(_00688_),
    .Y(_00783_));
 sg13g2_nand2_1 _07769_ (.Y(_00784_),
    .A(net1634),
    .B(_00684_));
 sg13g2_a21oi_1 _07770_ (.A1(_00783_),
    .A2(_00784_),
    .Y(_00012_),
    .B1(_00782_));
 sg13g2_nand3_1 _07771_ (.B(net1630),
    .C(_00685_),
    .A(net1634),
    .Y(_00785_));
 sg13g2_nand2b_1 _07772_ (.Y(_00786_),
    .B(_00704_),
    .A_N(_00694_));
 sg13g2_nand3_1 _07773_ (.B(_00785_),
    .C(_00786_),
    .A(_00756_),
    .Y(_00013_));
 sg13g2_xnor2_1 _07774_ (.Y(_00787_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[15] ),
    .B(net1808));
 sg13g2_xor2_1 _07775_ (.B(net1808),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[15] ),
    .X(_00788_));
 sg13g2_nor2_1 _07776_ (.A(_00619_),
    .B(_00620_),
    .Y(_00789_));
 sg13g2_nand2_1 _07777_ (.Y(_00790_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[12] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[12] ));
 sg13g2_xor2_1 _07778_ (.B(\vgadonut.donut.donuthit.cordicxy.xin[12] ),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[12] ),
    .X(_00791_));
 sg13g2_nor2_1 _07779_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[11] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[11] ),
    .Y(_00792_));
 sg13g2_xor2_1 _07780_ (.B(\vgadonut.donut.donuthit.cordicxy.xin[11] ),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[11] ),
    .X(_00793_));
 sg13g2_xnor2_1 _07781_ (.Y(_00794_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[11] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[11] ));
 sg13g2_nand2_1 _07782_ (.Y(_00795_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[10] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[10] ));
 sg13g2_xnor2_1 _07783_ (.Y(_00796_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[10] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[10] ));
 sg13g2_nor2_1 _07784_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[7] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[7] ),
    .Y(_00797_));
 sg13g2_nand2_1 _07785_ (.Y(_00798_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[7] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[7] ));
 sg13g2_xnor2_1 _07786_ (.Y(_00799_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[7] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[7] ));
 sg13g2_xnor2_1 _07787_ (.Y(_00800_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[6] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[6] ));
 sg13g2_nor2b_1 _07788_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[3] ),
    .B_N(\vgadonut.donut.donuthit.cordicxy.yin[3] ),
    .Y(_00801_));
 sg13g2_or2_1 _07789_ (.X(_00802_),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[3] ),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[3] ));
 sg13g2_and2_1 _07790_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[3] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[3] ),
    .X(_00803_));
 sg13g2_xnor2_1 _07791_ (.Y(_00804_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[3] ),
    .B(\vgadonut.donut.donuthit.cordicxy.yin[3] ));
 sg13g2_nor2b_1 _07792_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[2] ),
    .B_N(\vgadonut.donut.donuthit.cordicxy.yin[2] ),
    .Y(_00805_));
 sg13g2_and2_1 _07793_ (.A(net298),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[2] ),
    .X(_00806_));
 sg13g2_xor2_1 _07794_ (.B(\vgadonut.donut.donuthit.cordicxy.xin[2] ),
    .A(net297),
    .X(_00807_));
 sg13g2_xnor2_1 _07795_ (.Y(_00808_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[2] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[2] ));
 sg13g2_nor2b_1 _07796_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[1] ),
    .B_N(\vgadonut.donut.donuthit.cordicxy.yin[1] ),
    .Y(_00809_));
 sg13g2_xnor2_1 _07797_ (.Y(_00810_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[1] ),
    .B(\vgadonut.donut.donuthit.cordicxy.yin[1] ));
 sg13g2_nand2b_1 _07798_ (.Y(_00811_),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[0] ),
    .A_N(\vgadonut.donut.donuthit.cordicxy.yin[0] ));
 sg13g2_a21oi_2 _07799_ (.B1(_00809_),
    .Y(_00812_),
    .A2(_00811_),
    .A1(_00810_));
 sg13g2_nor2_1 _07800_ (.A(_00807_),
    .B(_00812_),
    .Y(_00813_));
 sg13g2_nor2_1 _07801_ (.A(_00805_),
    .B(_00813_),
    .Y(_00814_));
 sg13g2_nand2_1 _07802_ (.Y(_00815_),
    .A(_00804_),
    .B(_00808_));
 sg13g2_a21oi_1 _07803_ (.A1(net276),
    .A2(_00805_),
    .Y(_00816_),
    .B1(_00801_));
 sg13g2_o21ai_1 _07804_ (.B1(_00816_),
    .Y(_00817_),
    .A1(_00815_),
    .A2(_00812_));
 sg13g2_nand2b_1 _07805_ (.Y(_00818_),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[5] ),
    .A_N(\vgadonut.donut.donuthit.cordicxy.yin[5] ));
 sg13g2_nor2b_1 _07806_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[5] ),
    .B_N(net295),
    .Y(_00819_));
 sg13g2_xnor2_1 _07807_ (.Y(_00820_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[5] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[5] ));
 sg13g2_xor2_1 _07808_ (.B(\vgadonut.donut.donuthit.cordicxy.xin[5] ),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[5] ),
    .X(_00821_));
 sg13g2_nand2_1 _07809_ (.Y(_00822_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[4] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[4] ));
 sg13g2_xor2_1 _07810_ (.B(\vgadonut.donut.donuthit.cordicxy.xin[4] ),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[4] ),
    .X(_00823_));
 sg13g2_xnor2_1 _07811_ (.Y(_00824_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[4] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[4] ));
 sg13g2_nor2_1 _07812_ (.A(_00821_),
    .B(_00823_),
    .Y(_00825_));
 sg13g2_and3_1 _07813_ (.X(_00826_),
    .A(_00799_),
    .B(_00800_),
    .C(_00825_));
 sg13g2_nand2_1 _07814_ (.Y(_00827_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[7] ),
    .B(_00622_));
 sg13g2_nor2b_1 _07815_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[4] ),
    .B_N(\vgadonut.donut.donuthit.cordicxy.yin[4] ),
    .Y(_00828_));
 sg13g2_a221oi_1 _07816_ (.B2(_00828_),
    .C1(_00819_),
    .B1(_00818_),
    .A1(\vgadonut.donut.donuthit.cordicxy.yin[6] ),
    .Y(_00829_),
    .A2(_00623_));
 sg13g2_o21ai_1 _07817_ (.B1(_00799_),
    .Y(_00830_),
    .A1(\vgadonut.donut.donuthit.cordicxy.yin[6] ),
    .A2(_00623_));
 sg13g2_o21ai_1 _07818_ (.B1(_00827_),
    .Y(_00831_),
    .A1(_00829_),
    .A2(_00830_));
 sg13g2_a21o_2 _07819_ (.A2(_00817_),
    .A1(_00826_),
    .B1(_00831_),
    .X(_00832_));
 sg13g2_nor2b_1 _07820_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[9] ),
    .B_N(\vgadonut.donut.donuthit.cordicxy.xin[9] ),
    .Y(_00833_));
 sg13g2_nand2b_1 _07821_ (.Y(_00834_),
    .B(\vgadonut.donut.donuthit.cordicxy.yin[9] ),
    .A_N(\vgadonut.donut.donuthit.cordicxy.xin[9] ));
 sg13g2_nor2b_2 _07822_ (.A(_00833_),
    .B_N(_00834_),
    .Y(_00835_));
 sg13g2_nand2_1 _07823_ (.Y(_00836_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[8] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[8] ));
 sg13g2_xnor2_1 _07824_ (.Y(_00837_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[8] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[8] ));
 sg13g2_inv_1 _07825_ (.Y(_00838_),
    .A(_00837_));
 sg13g2_and2_1 _07826_ (.A(_00835_),
    .B(_00837_),
    .X(_00839_));
 sg13g2_and3_1 _07827_ (.X(_00840_),
    .A(_00794_),
    .B(_00796_),
    .C(_00839_));
 sg13g2_nand2b_1 _07828_ (.Y(_00841_),
    .B(\vgadonut.donut.donuthit.cordicxy.yin[11] ),
    .A_N(\vgadonut.donut.donuthit.cordicxy.xin[11] ));
 sg13g2_nor2b_1 _07829_ (.A(\vgadonut.donut.donuthit.cordicxy.xin[10] ),
    .B_N(\vgadonut.donut.donuthit.cordicxy.yin[10] ),
    .Y(_00842_));
 sg13g2_nand2b_1 _07830_ (.Y(_00843_),
    .B(\vgadonut.donut.donuthit.cordicxy.yin[8] ),
    .A_N(\vgadonut.donut.donuthit.cordicxy.xin[8] ));
 sg13g2_o21ai_1 _07831_ (.B1(_00834_),
    .Y(_00844_),
    .A1(_00833_),
    .A2(_00843_));
 sg13g2_a21oi_1 _07832_ (.A1(_00796_),
    .A2(_00844_),
    .Y(_00845_),
    .B1(_00842_));
 sg13g2_o21ai_1 _07833_ (.B1(_00841_),
    .Y(_00846_),
    .A1(_00793_),
    .A2(_00845_));
 sg13g2_a21o_1 _07834_ (.A2(_00840_),
    .A1(_00832_),
    .B1(_00846_),
    .X(_00847_));
 sg13g2_nor2b_1 _07835_ (.A(_00791_),
    .B_N(_00847_),
    .Y(_00848_));
 sg13g2_nor2_1 _07836_ (.A(\vgadonut.donut.donuthit.cordicxy.yin[13] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[13] ),
    .Y(_00849_));
 sg13g2_nand2_1 _07837_ (.Y(_00850_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[13] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[13] ));
 sg13g2_nor2b_2 _07838_ (.A(_00849_),
    .B_N(_00850_),
    .Y(_00851_));
 sg13g2_a21oi_1 _07839_ (.A1(\vgadonut.donut.donuthit.cordicxy.yin[12] ),
    .A2(_00620_),
    .Y(_00852_),
    .B1(_00848_));
 sg13g2_nor2_1 _07840_ (.A(_00791_),
    .B(_00851_),
    .Y(_00853_));
 sg13g2_nor3_1 _07841_ (.A(_00619_),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[12] ),
    .C(_00851_),
    .Y(_00854_));
 sg13g2_a221oi_1 _07842_ (.B2(_00847_),
    .C1(_00854_),
    .B1(_00853_),
    .A1(_00851_),
    .Y(_00855_),
    .A2(_00852_));
 sg13g2_nor2_1 _07843_ (.A(_00794_),
    .B(_00796_),
    .Y(_00856_));
 sg13g2_nor2_1 _07844_ (.A(_00792_),
    .B(_00795_),
    .Y(_00857_));
 sg13g2_nand2_1 _07845_ (.Y(_00858_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[9] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[9] ));
 sg13g2_nor2_1 _07846_ (.A(_00799_),
    .B(_00800_),
    .Y(_00859_));
 sg13g2_nand2_1 _07847_ (.Y(_00860_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[6] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[6] ));
 sg13g2_a21oi_2 _07848_ (.B1(_00797_),
    .Y(_00861_),
    .A2(_00860_),
    .A1(_00798_));
 sg13g2_and2_1 _07849_ (.A(net295),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[5] ),
    .X(_00862_));
 sg13g2_nand2_1 _07850_ (.Y(_00863_),
    .A(net293),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[1] ));
 sg13g2_nand2_1 _07851_ (.Y(_00864_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[0] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[0] ));
 sg13g2_o21ai_1 _07852_ (.B1(_00863_),
    .Y(_00865_),
    .A1(_00864_),
    .A2(_00810_));
 sg13g2_a21oi_1 _07853_ (.A1(_00807_),
    .A2(_00865_),
    .Y(_00866_),
    .B1(_00806_));
 sg13g2_nor2_1 _07854_ (.A(_00804_),
    .B(_00808_),
    .Y(_00867_));
 sg13g2_a221oi_1 _07855_ (.B2(_00865_),
    .C1(_00803_),
    .B1(_00867_),
    .A1(_00802_),
    .Y(_00868_),
    .A2(_00806_));
 sg13g2_nor2_1 _07856_ (.A(_00820_),
    .B(_00822_),
    .Y(_00869_));
 sg13g2_o21ai_1 _07857_ (.B1(_00859_),
    .Y(_00870_),
    .A1(_00862_),
    .A2(_00869_));
 sg13g2_nand3_1 _07858_ (.B(_00823_),
    .C(_00859_),
    .A(_00821_),
    .Y(_00871_));
 sg13g2_o21ai_1 _07859_ (.B1(_00870_),
    .Y(_00872_),
    .A1(_00871_),
    .A2(_00868_));
 sg13g2_nor2_1 _07860_ (.A(_00861_),
    .B(_00872_),
    .Y(_00873_));
 sg13g2_o21ai_1 _07861_ (.B1(_00838_),
    .Y(_00874_),
    .A1(_00861_),
    .A2(net280));
 sg13g2_nor4_1 _07862_ (.A(_00794_),
    .B(_00796_),
    .C(_00835_),
    .D(_00837_),
    .Y(_00875_));
 sg13g2_o21ai_1 _07863_ (.B1(_00875_),
    .Y(_00876_),
    .A1(_00872_),
    .A2(_00861_));
 sg13g2_o21ai_1 _07864_ (.B1(_00858_),
    .Y(_00877_),
    .A1(_00835_),
    .A2(_00836_));
 sg13g2_a221oi_1 _07865_ (.B2(_00877_),
    .C1(_00857_),
    .B1(_00856_),
    .A1(\vgadonut.donut.donuthit.cordicxy.yin[11] ),
    .Y(_00878_),
    .A2(\vgadonut.donut.donuthit.cordicxy.xin[11] ));
 sg13g2_nand2_1 _07866_ (.Y(_00879_),
    .A(net290),
    .B(_00878_));
 sg13g2_a21oi_1 _07867_ (.A1(_00791_),
    .A2(_00879_),
    .Y(_00880_),
    .B1(_00789_));
 sg13g2_xnor2_1 _07868_ (.Y(_00881_),
    .A(_00851_),
    .B(_00880_));
 sg13g2_mux2_1 _07869_ (.A0(_00855_),
    .A1(_00881_),
    .S(net1793),
    .X(_00882_));
 sg13g2_xnor2_1 _07870_ (.Y(_00883_),
    .A(net1806),
    .B(_00882_));
 sg13g2_nand2_1 _07871_ (.Y(_00884_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[14] ),
    .B(\vgadonut.donut.donuthit.cordicxy.xin[14] ));
 sg13g2_nand2b_1 _07872_ (.Y(_00885_),
    .B(\vgadonut.donut.donuthit.cordicxy.yin[14] ),
    .A_N(\vgadonut.donut.donuthit.cordicxy.xin[14] ));
 sg13g2_xor2_1 _07873_ (.B(\vgadonut.donut.donuthit.cordicxy.xin[14] ),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[14] ),
    .X(_00886_));
 sg13g2_nand2_1 _07874_ (.Y(_00887_),
    .A(_00791_),
    .B(_00851_));
 sg13g2_a21oi_2 _07875_ (.B1(_00887_),
    .Y(_00888_),
    .A2(_00878_),
    .A1(_00876_));
 sg13g2_o21ai_1 _07876_ (.B1(_00850_),
    .Y(_00889_),
    .A1(_00790_),
    .A2(_00849_));
 sg13g2_nor2_1 _07877_ (.A(_00888_),
    .B(_00889_),
    .Y(_00890_));
 sg13g2_o21ai_1 _07878_ (.B1(_00886_),
    .Y(_00891_),
    .A1(_00889_),
    .A2(_00888_));
 sg13g2_a221oi_1 _07879_ (.B2(_00853_),
    .C1(_00854_),
    .B1(_00847_),
    .A1(\vgadonut.donut.donuthit.cordicxy.yin[13] ),
    .Y(_00892_),
    .A2(_00618_));
 sg13g2_o21ai_1 _07880_ (.B1(_00885_),
    .Y(_00893_),
    .A1(_00892_),
    .A2(_00886_));
 sg13g2_and2_1 _07881_ (.A(net1792),
    .B(_00893_),
    .X(_00894_));
 sg13g2_nand2_2 _07882_ (.Y(_00895_),
    .A(_00893_),
    .B(net1792));
 sg13g2_a21oi_2 _07883_ (.B1(net1792),
    .Y(_00896_),
    .A2(_00891_),
    .A1(_00884_));
 sg13g2_a21o_1 _07884_ (.A2(_00884_),
    .A1(_00891_),
    .B1(net1792),
    .X(_00897_));
 sg13g2_nand2_1 _07885_ (.Y(_00898_),
    .A(_00895_),
    .B(_00897_));
 sg13g2_xnor2_1 _07886_ (.Y(_00899_),
    .A(_00886_),
    .B(_00890_));
 sg13g2_xnor2_1 _07887_ (.Y(_00900_),
    .A(_00886_),
    .B(_00892_));
 sg13g2_nor2_1 _07888_ (.A(net1782),
    .B(_00900_),
    .Y(_00901_));
 sg13g2_a21oi_2 _07889_ (.B1(_00901_),
    .Y(_00902_),
    .A2(_00899_),
    .A1(net1782));
 sg13g2_xnor2_1 _07890_ (.Y(_00903_),
    .A(net1625),
    .B(_00902_));
 sg13g2_nor2_1 _07891_ (.A(_00883_),
    .B(_00903_),
    .Y(_00904_));
 sg13g2_nor2_1 _07892_ (.A(net1793),
    .B(_00900_),
    .Y(_00905_));
 sg13g2_a21oi_1 _07893_ (.A1(net1793),
    .A2(_00899_),
    .Y(_00906_),
    .B1(_00905_));
 sg13g2_xnor2_1 _07894_ (.Y(_00907_),
    .A(net1806),
    .B(_00906_));
 sg13g2_xnor2_1 _07895_ (.Y(_00908_),
    .A(_00883_),
    .B(_00903_));
 sg13g2_xor2_1 _07896_ (.B(_00847_),
    .A(_00791_),
    .X(_00909_));
 sg13g2_nor2_1 _07897_ (.A(net1793),
    .B(_00909_),
    .Y(_00910_));
 sg13g2_xor2_1 _07898_ (.B(_00879_),
    .A(_00791_),
    .X(_00911_));
 sg13g2_a21oi_1 _07899_ (.A1(net1793),
    .A2(_00911_),
    .Y(_00912_),
    .B1(_00910_));
 sg13g2_xnor2_1 _07900_ (.Y(_00913_),
    .A(net1806),
    .B(_00912_));
 sg13g2_mux2_2 _07901_ (.A0(_00855_),
    .A1(_00881_),
    .S(net1783),
    .X(_00914_));
 sg13g2_inv_1 _07902_ (.Y(_00915_),
    .A(_00914_));
 sg13g2_xnor2_1 _07903_ (.Y(_00916_),
    .A(net1624),
    .B(_00914_));
 sg13g2_nand2_1 _07904_ (.Y(_00917_),
    .A(_00913_),
    .B(_00916_));
 sg13g2_xnor2_1 _07905_ (.Y(_00918_),
    .A(_00913_),
    .B(_00916_));
 sg13g2_a21oi_1 _07906_ (.A1(_00884_),
    .A2(_00891_),
    .Y(_00919_),
    .B1(net1782));
 sg13g2_a21o_2 _07907_ (.A2(_00893_),
    .A1(net1782),
    .B1(_00919_),
    .X(_00920_));
 sg13g2_xnor2_1 _07908_ (.Y(_00921_),
    .A(net1806),
    .B(net1627));
 sg13g2_xor2_1 _07909_ (.B(net1618),
    .A(_00920_),
    .X(_00922_));
 sg13g2_nor2_1 _07910_ (.A(_00902_),
    .B(_00922_),
    .Y(_00923_));
 sg13g2_xor2_1 _07911_ (.B(_00922_),
    .A(_00902_),
    .X(_00924_));
 sg13g2_a21oi_1 _07912_ (.A1(_00817_),
    .A2(_00824_),
    .Y(_00925_),
    .B1(_00828_));
 sg13g2_xnor2_1 _07913_ (.Y(_00926_),
    .A(_00820_),
    .B(_00925_));
 sg13g2_o21ai_1 _07914_ (.B1(_00822_),
    .Y(_00927_),
    .A1(_00824_),
    .A2(net278));
 sg13g2_xnor2_1 _07915_ (.Y(_00928_),
    .A(_00821_),
    .B(_00927_));
 sg13g2_nor2_1 _07916_ (.A(net1784),
    .B(_00928_),
    .Y(_00929_));
 sg13g2_a21oi_1 _07917_ (.A1(net1784),
    .A2(_00926_),
    .Y(_00930_),
    .B1(_00929_));
 sg13g2_xnor2_1 _07918_ (.Y(_00931_),
    .A(net1807),
    .B(_00930_));
 sg13g2_xor2_1 _07919_ (.B(_00931_),
    .A(net1623),
    .X(_00932_));
 sg13g2_xnor2_1 _07920_ (.Y(_00933_),
    .A(_00823_),
    .B(_00868_));
 sg13g2_nand2_1 _07921_ (.Y(_00934_),
    .A(net1784),
    .B(_00933_));
 sg13g2_xnor2_1 _07922_ (.Y(_00935_),
    .A(net286),
    .B(_00824_));
 sg13g2_o21ai_1 _07923_ (.B1(_00934_),
    .Y(_00936_),
    .A1(net1784),
    .A2(_00935_));
 sg13g2_nand2_1 _07924_ (.Y(_00937_),
    .A(_00932_),
    .B(_00936_));
 sg13g2_xor2_1 _07925_ (.B(_00936_),
    .A(_00932_),
    .X(_00938_));
 sg13g2_nand2_1 _07926_ (.Y(_00939_),
    .A(net1791),
    .B(_00933_));
 sg13g2_o21ai_1 _07927_ (.B1(_00939_),
    .Y(_00940_),
    .A1(net1792),
    .A2(_00935_));
 sg13g2_xor2_1 _07928_ (.B(_00940_),
    .A(net1807),
    .X(_00941_));
 sg13g2_xor2_1 _07929_ (.B(_00941_),
    .A(net1623),
    .X(_00942_));
 sg13g2_xor2_1 _07930_ (.B(_00866_),
    .A(net277),
    .X(_00943_));
 sg13g2_xor2_1 _07931_ (.B(_00814_),
    .A(net277),
    .X(_00944_));
 sg13g2_nor2_1 _07932_ (.A(net1785),
    .B(_00944_),
    .Y(_00945_));
 sg13g2_a21oi_2 _07933_ (.B1(_00945_),
    .Y(_00946_),
    .A2(_00943_),
    .A1(net1785));
 sg13g2_nor2b_2 _07934_ (.A(_00946_),
    .B_N(_00942_),
    .Y(_00947_));
 sg13g2_nand2b_1 _07935_ (.Y(_00948_),
    .B(_00946_),
    .A_N(_00942_));
 sg13g2_nor2_1 _07936_ (.A(net1785),
    .B(_00943_),
    .Y(_00949_));
 sg13g2_a21oi_1 _07937_ (.A1(net1785),
    .A2(_00944_),
    .Y(_00950_),
    .B1(_00949_));
 sg13g2_xnor2_1 _07938_ (.Y(_00951_),
    .A(net1807),
    .B(_00950_));
 sg13g2_inv_1 _07939_ (.Y(_00952_),
    .A(_00951_));
 sg13g2_nand3_1 _07940_ (.B(net283),
    .C(_00952_),
    .A(_00895_),
    .Y(_00953_));
 sg13g2_o21ai_1 _07941_ (.B1(_00951_),
    .Y(_00954_),
    .A1(_00894_),
    .A2(_00896_));
 sg13g2_xnor2_1 _07942_ (.Y(_00955_),
    .A(_00807_),
    .B(net285));
 sg13g2_nor2_1 _07943_ (.A(net1795),
    .B(_00955_),
    .Y(_00956_));
 sg13g2_xnor2_1 _07944_ (.Y(_00957_),
    .A(_00808_),
    .B(_00812_));
 sg13g2_a21oi_2 _07945_ (.B1(_00956_),
    .Y(_00958_),
    .A2(_00957_),
    .A1(net1795));
 sg13g2_inv_1 _07946_ (.Y(_00959_),
    .A(_00958_));
 sg13g2_a21oi_1 _07947_ (.A1(_00953_),
    .A2(_00954_),
    .Y(_00960_),
    .B1(_00958_));
 sg13g2_nand3_1 _07948_ (.B(_00954_),
    .C(_00959_),
    .A(_00953_),
    .Y(_00961_));
 sg13g2_a21o_1 _07949_ (.A2(_00954_),
    .A1(_00953_),
    .B1(_00959_),
    .X(_00962_));
 sg13g2_nand2_1 _07950_ (.Y(_00963_),
    .A(_00961_),
    .B(_00962_));
 sg13g2_xnor2_1 _07951_ (.Y(_00964_),
    .A(net275),
    .B(_00864_));
 sg13g2_xor2_1 _07952_ (.B(_00811_),
    .A(net274),
    .X(_00965_));
 sg13g2_nand2_1 _07953_ (.Y(_00966_),
    .A(net1795),
    .B(_00965_));
 sg13g2_o21ai_1 _07954_ (.B1(_00966_),
    .Y(_00967_),
    .A1(net1795),
    .A2(_00964_));
 sg13g2_nor2_1 _07955_ (.A(net1785),
    .B(_00955_),
    .Y(_00968_));
 sg13g2_a21oi_1 _07956_ (.A1(net1785),
    .A2(_00957_),
    .Y(_00969_),
    .B1(_00968_));
 sg13g2_xnor2_1 _07957_ (.Y(_00970_),
    .A(net1808),
    .B(_00969_));
 sg13g2_inv_1 _07958_ (.Y(_00971_),
    .A(_00970_));
 sg13g2_a21oi_1 _07959_ (.A1(_00895_),
    .A2(net283),
    .Y(_00972_),
    .B1(_00970_));
 sg13g2_nor3_1 _07960_ (.A(_00894_),
    .B(_00896_),
    .C(_00971_),
    .Y(_00973_));
 sg13g2_o21ai_1 _07961_ (.B1(_00967_),
    .Y(_00974_),
    .A1(_00972_),
    .A2(_00973_));
 sg13g2_nor3_1 _07962_ (.A(_00967_),
    .B(_00972_),
    .C(_00973_),
    .Y(_00975_));
 sg13g2_nand2_1 _07963_ (.Y(_00976_),
    .A(net1785),
    .B(_00965_));
 sg13g2_o21ai_1 _07964_ (.B1(_00976_),
    .Y(_00977_),
    .A1(net1785),
    .A2(_00964_));
 sg13g2_xor2_1 _07965_ (.B(_00977_),
    .A(net1808),
    .X(_00978_));
 sg13g2_o21ai_1 _07966_ (.B1(_00978_),
    .Y(_00979_),
    .A1(_00894_),
    .A2(_00896_));
 sg13g2_xor2_1 _07967_ (.B(\vgadonut.donut.donuthit.cordicxy.xin[0] ),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[0] ),
    .X(_00980_));
 sg13g2_nand3b_1 _07968_ (.B(net284),
    .C(_00895_),
    .Y(_00981_),
    .A_N(_00978_));
 sg13g2_nand3_1 _07969_ (.B(_00980_),
    .C(_00981_),
    .A(_00979_),
    .Y(_00982_));
 sg13g2_a21oi_1 _07970_ (.A1(_00974_),
    .A2(_00982_),
    .Y(_00983_),
    .B1(_00975_));
 sg13g2_a221oi_1 _07971_ (.B2(_00982_),
    .C1(_00975_),
    .B1(_00974_),
    .A1(_00961_),
    .Y(_00984_),
    .A2(_00962_));
 sg13g2_nor2_1 _07972_ (.A(_00960_),
    .B(_00984_),
    .Y(_00985_));
 sg13g2_or3_1 _07973_ (.A(_00947_),
    .B(_00960_),
    .C(_00984_),
    .X(_00986_));
 sg13g2_nand3_1 _07974_ (.B(_00948_),
    .C(_00986_),
    .A(_00938_),
    .Y(_00987_));
 sg13g2_a221oi_1 _07975_ (.B2(_00818_),
    .C1(_00819_),
    .B1(_00828_),
    .A1(_00817_),
    .Y(_00988_),
    .A2(_00825_));
 sg13g2_nor2b_1 _07976_ (.A(_00988_),
    .B_N(_00800_),
    .Y(_00989_));
 sg13g2_xnor2_1 _07977_ (.Y(_00990_),
    .A(_00800_),
    .B(_00988_));
 sg13g2_a21oi_1 _07978_ (.A1(_00821_),
    .A2(_00927_),
    .Y(_00991_),
    .B1(_00862_));
 sg13g2_xnor2_1 _07979_ (.Y(_00992_),
    .A(_00800_),
    .B(_00991_));
 sg13g2_nor2_1 _07980_ (.A(net1791),
    .B(_00990_),
    .Y(_00993_));
 sg13g2_a21oi_1 _07981_ (.A1(net1791),
    .A2(_00992_),
    .Y(_00994_),
    .B1(_00993_));
 sg13g2_xor2_1 _07982_ (.B(_00994_),
    .A(net1807),
    .X(_00995_));
 sg13g2_xor2_1 _07983_ (.B(_00995_),
    .A(net1623),
    .X(_00996_));
 sg13g2_inv_1 _07984_ (.Y(_00997_),
    .A(_00996_));
 sg13g2_nor2_1 _07985_ (.A(net1791),
    .B(_00928_),
    .Y(_00998_));
 sg13g2_a21oi_2 _07986_ (.B1(_00998_),
    .Y(_00999_),
    .A2(_00926_),
    .A1(net1792));
 sg13g2_nand2b_1 _07987_ (.Y(_01000_),
    .B(_00996_),
    .A_N(_00999_));
 sg13g2_and2_1 _07988_ (.A(_00937_),
    .B(_01000_),
    .X(_01001_));
 sg13g2_nor2b_1 _07989_ (.A(_00996_),
    .B_N(_00999_),
    .Y(_01002_));
 sg13g2_a21o_1 _07990_ (.A2(_01001_),
    .A1(_00987_),
    .B1(_01002_),
    .X(_01003_));
 sg13g2_a21oi_1 _07991_ (.A1(\vgadonut.donut.donuthit.cordicxy.yin[6] ),
    .A2(_00623_),
    .Y(_01004_),
    .B1(_00989_));
 sg13g2_xnor2_1 _07992_ (.Y(_01005_),
    .A(_00799_),
    .B(_01004_));
 sg13g2_o21ai_1 _07993_ (.B1(_00860_),
    .Y(_01006_),
    .A1(_00800_),
    .A2(_00991_));
 sg13g2_xor2_1 _07994_ (.B(_01006_),
    .A(_00799_),
    .X(_01007_));
 sg13g2_nor2_1 _07995_ (.A(net1784),
    .B(_01007_),
    .Y(_01008_));
 sg13g2_a21oi_1 _07996_ (.A1(net1784),
    .A2(_01005_),
    .Y(_01009_),
    .B1(_01008_));
 sg13g2_xnor2_1 _07997_ (.Y(_01010_),
    .A(_01009_),
    .B(net1807));
 sg13g2_xor2_1 _07998_ (.B(net1623),
    .A(_01010_),
    .X(_01011_));
 sg13g2_nor2_1 _07999_ (.A(net1791),
    .B(_00992_),
    .Y(_01012_));
 sg13g2_a21oi_2 _08000_ (.B1(_01012_),
    .Y(_01013_),
    .A2(_00990_),
    .A1(net1791));
 sg13g2_inv_1 _08001_ (.Y(_01014_),
    .A(_01013_));
 sg13g2_nor2_1 _08002_ (.A(_01011_),
    .B(_01014_),
    .Y(_01015_));
 sg13g2_nand2_1 _08003_ (.Y(_01016_),
    .A(_01011_),
    .B(_01014_));
 sg13g2_xnor2_1 _08004_ (.Y(_01017_),
    .A(_01011_),
    .B(_01013_));
 sg13g2_nand2_1 _08005_ (.Y(_01018_),
    .A(_00832_),
    .B(_00837_));
 sg13g2_xnor2_1 _08006_ (.Y(_01019_),
    .A(_00832_),
    .B(_00837_));
 sg13g2_nor2_1 _08007_ (.A(net1794),
    .B(_01019_),
    .Y(_01020_));
 sg13g2_xnor2_1 _08008_ (.Y(_01021_),
    .A(_00838_),
    .B(_00873_));
 sg13g2_a21oi_1 _08009_ (.A1(net1794),
    .A2(_01021_),
    .Y(_01022_),
    .B1(_01020_));
 sg13g2_xnor2_1 _08010_ (.Y(_01023_),
    .A(net1806),
    .B(_01022_));
 sg13g2_xor2_1 _08011_ (.B(_01023_),
    .A(net1623),
    .X(_01024_));
 sg13g2_nand2_1 _08012_ (.Y(_01025_),
    .A(net1791),
    .B(_01005_));
 sg13g2_o21ai_1 _08013_ (.B1(_01025_),
    .Y(_01026_),
    .A1(net1791),
    .A2(net287));
 sg13g2_nand2_1 _08014_ (.Y(_01027_),
    .A(_01024_),
    .B(_01026_));
 sg13g2_nor2_1 _08015_ (.A(_01024_),
    .B(_01026_),
    .Y(_01028_));
 sg13g2_xor2_1 _08016_ (.B(_01026_),
    .A(_01024_),
    .X(_01029_));
 sg13g2_nand2_1 _08017_ (.Y(_01030_),
    .A(_01017_),
    .B(_01029_));
 sg13g2_a221oi_1 _08018_ (.B2(_01001_),
    .C1(_01030_),
    .B1(_00987_),
    .A1(_00997_),
    .Y(_01031_),
    .A2(_00999_));
 sg13g2_a21oi_1 _08019_ (.A1(_01016_),
    .A2(_01027_),
    .Y(_01032_),
    .B1(_01028_));
 sg13g2_nor2_2 _08020_ (.A(net279),
    .B(_01032_),
    .Y(_01033_));
 sg13g2_a21o_1 _08021_ (.A2(_00839_),
    .A1(_00832_),
    .B1(_00844_),
    .X(_01034_));
 sg13g2_a21oi_1 _08022_ (.A1(_00796_),
    .A2(_01034_),
    .Y(_01035_),
    .B1(_00842_));
 sg13g2_xnor2_1 _08023_ (.Y(_01036_),
    .A(_00793_),
    .B(_01035_));
 sg13g2_nor2_1 _08024_ (.A(net1793),
    .B(_01036_),
    .Y(_01037_));
 sg13g2_a21oi_2 _08025_ (.B1(_00835_),
    .Y(_01038_),
    .A2(_00874_),
    .A1(_00836_));
 sg13g2_a21oi_2 _08026_ (.B1(_01038_),
    .Y(_01039_),
    .A2(\vgadonut.donut.donuthit.cordicxy.xin[9] ),
    .A1(\vgadonut.donut.donuthit.cordicxy.yin[9] ));
 sg13g2_o21ai_1 _08027_ (.B1(_00795_),
    .Y(_01040_),
    .A1(_00796_),
    .A2(_01039_));
 sg13g2_xnor2_1 _08028_ (.Y(_01041_),
    .A(_00794_),
    .B(_01040_));
 sg13g2_a21oi_2 _08029_ (.B1(_01037_),
    .Y(_01042_),
    .A2(_01041_),
    .A1(net1793));
 sg13g2_xnor2_1 _08030_ (.Y(_01043_),
    .A(net1806),
    .B(_01042_));
 sg13g2_xnor2_1 _08031_ (.Y(_01044_),
    .A(net1618),
    .B(_01042_));
 sg13g2_xor2_1 _08032_ (.B(_01039_),
    .A(_00796_),
    .X(_01045_));
 sg13g2_nand2_1 _08033_ (.Y(_01046_),
    .A(net1783),
    .B(_01045_));
 sg13g2_xnor2_1 _08034_ (.Y(_01047_),
    .A(_00796_),
    .B(_01034_));
 sg13g2_o21ai_1 _08035_ (.B1(_01046_),
    .Y(_01048_),
    .A1(net1783),
    .A2(_01047_));
 sg13g2_nand2b_1 _08036_ (.Y(_01049_),
    .B(_01048_),
    .A_N(_01044_));
 sg13g2_xor2_1 _08037_ (.B(_01048_),
    .A(_01044_),
    .X(_01050_));
 sg13g2_xor2_1 _08038_ (.B(_00913_),
    .A(net1625),
    .X(_01051_));
 sg13g2_inv_1 _08039_ (.Y(_01052_),
    .A(_01051_));
 sg13g2_nor2_1 _08040_ (.A(net1783),
    .B(_01036_),
    .Y(_01053_));
 sg13g2_a21oi_2 _08041_ (.B1(_01053_),
    .Y(_01054_),
    .A2(_01041_),
    .A1(net1783));
 sg13g2_nor2_1 _08042_ (.A(_01052_),
    .B(_01054_),
    .Y(_01055_));
 sg13g2_xor2_1 _08043_ (.B(_01054_),
    .A(_01051_),
    .X(_01056_));
 sg13g2_nand2_1 _08044_ (.Y(_01057_),
    .A(_00843_),
    .B(_01018_));
 sg13g2_xnor2_1 _08045_ (.Y(_01058_),
    .A(_00835_),
    .B(_01057_));
 sg13g2_nor2_1 _08046_ (.A(net1794),
    .B(_01058_),
    .Y(_01059_));
 sg13g2_nand3_1 _08047_ (.B(_00836_),
    .C(_00874_),
    .A(_00835_),
    .Y(_01060_));
 sg13g2_nor2b_2 _08048_ (.A(_01038_),
    .B_N(_01060_),
    .Y(_01061_));
 sg13g2_a21oi_1 _08049_ (.A1(net1793),
    .A2(_01061_),
    .Y(_01062_),
    .B1(_01059_));
 sg13g2_xnor2_1 _08050_ (.Y(_01063_),
    .A(net1806),
    .B(_01062_));
 sg13g2_xor2_1 _08051_ (.B(_01063_),
    .A(net1624),
    .X(_01064_));
 sg13g2_nor2_1 _08052_ (.A(net1783),
    .B(_01019_),
    .Y(_01065_));
 sg13g2_a21oi_2 _08053_ (.B1(_01065_),
    .Y(_01066_),
    .A2(_01021_),
    .A1(net1783));
 sg13g2_inv_1 _08054_ (.Y(_01067_),
    .A(_01066_));
 sg13g2_nand2_1 _08055_ (.Y(_01068_),
    .A(_01064_),
    .B(_01067_));
 sg13g2_xnor2_1 _08056_ (.Y(_01069_),
    .A(_01064_),
    .B(_01066_));
 sg13g2_inv_1 _08057_ (.Y(_01070_),
    .A(_01069_));
 sg13g2_nor2_1 _08058_ (.A(net1794),
    .B(_01047_),
    .Y(_01071_));
 sg13g2_a21oi_1 _08059_ (.A1(net1794),
    .A2(_01045_),
    .Y(_01072_),
    .B1(_01071_));
 sg13g2_xnor2_1 _08060_ (.Y(_01073_),
    .A(net1806),
    .B(_01072_));
 sg13g2_inv_1 _08061_ (.Y(_01074_),
    .A(_01073_));
 sg13g2_xor2_1 _08062_ (.B(_01073_),
    .A(net1625),
    .X(_01075_));
 sg13g2_nor2_1 _08063_ (.A(net1782),
    .B(_01058_),
    .Y(_01076_));
 sg13g2_a21oi_2 _08064_ (.B1(_01076_),
    .Y(_01077_),
    .A2(_01061_),
    .A1(net1784));
 sg13g2_a21o_1 _08065_ (.A2(_01061_),
    .A1(net1782),
    .B1(_01076_),
    .X(_01078_));
 sg13g2_nor2_1 _08066_ (.A(_01075_),
    .B(_01078_),
    .Y(_01079_));
 sg13g2_xnor2_1 _08067_ (.Y(_01080_),
    .A(_01075_),
    .B(_01077_));
 sg13g2_nand2_1 _08068_ (.Y(_01081_),
    .A(_01069_),
    .B(_01080_));
 sg13g2_nor3_1 _08069_ (.A(_01050_),
    .B(_01056_),
    .C(_01081_),
    .Y(_01082_));
 sg13g2_o21ai_1 _08070_ (.B1(_01082_),
    .Y(_01083_),
    .A1(_01031_),
    .A2(_01032_));
 sg13g2_a22oi_1 _08071_ (.Y(_01084_),
    .B1(_01075_),
    .B2(_01078_),
    .A2(_01067_),
    .A1(_01064_));
 sg13g2_or2_1 _08072_ (.X(_01085_),
    .B(_01084_),
    .A(_01079_));
 sg13g2_nor3_1 _08073_ (.A(_01050_),
    .B(_01056_),
    .C(_01085_),
    .Y(_01086_));
 sg13g2_a21oi_1 _08074_ (.A1(_01052_),
    .A2(_01054_),
    .Y(_01087_),
    .B1(_01049_));
 sg13g2_nor3_1 _08075_ (.A(_01055_),
    .B(_01086_),
    .C(_01087_),
    .Y(_01088_));
 sg13g2_nand2_1 _08076_ (.Y(_01089_),
    .A(_01083_),
    .B(_01088_));
 sg13g2_xnor2_1 _08077_ (.Y(_01090_),
    .A(_00883_),
    .B(net1624));
 sg13g2_nand2_1 _08078_ (.Y(_01091_),
    .A(net1782),
    .B(_00911_));
 sg13g2_o21ai_1 _08079_ (.B1(_01091_),
    .Y(_01092_),
    .A1(net1782),
    .A2(_00909_));
 sg13g2_nand2_1 _08080_ (.Y(_01093_),
    .A(_01090_),
    .B(_01092_));
 sg13g2_inv_1 _08081_ (.Y(_01094_),
    .A(_01093_));
 sg13g2_xor2_1 _08082_ (.B(_01092_),
    .A(_01090_),
    .X(_01095_));
 sg13g2_xnor2_1 _08083_ (.Y(_01096_),
    .A(net1624),
    .B(_00907_));
 sg13g2_nand2_1 _08084_ (.Y(_01097_),
    .A(_00915_),
    .B(_01096_));
 sg13g2_xnor2_1 _08085_ (.Y(_01098_),
    .A(_00914_),
    .B(_01096_));
 sg13g2_nand2_1 _08086_ (.Y(_01099_),
    .A(_01095_),
    .B(_01098_));
 sg13g2_a21oi_1 _08087_ (.A1(_01083_),
    .A2(_01088_),
    .Y(_01100_),
    .B1(_01099_));
 sg13g2_o21ai_1 _08088_ (.B1(_01093_),
    .Y(_01101_),
    .A1(_00915_),
    .A2(_01096_));
 sg13g2_a21o_1 _08089_ (.A2(_01101_),
    .A1(_01097_),
    .B1(_01100_),
    .X(_01102_));
 sg13g2_xnor2_1 _08090_ (.Y(_01103_),
    .A(_00924_),
    .B(_01102_));
 sg13g2_a21oi_1 _08091_ (.A1(_00924_),
    .A2(_01102_),
    .Y(_01104_),
    .B1(_00923_));
 sg13g2_xor2_1 _08092_ (.B(_00920_),
    .A(_00142_),
    .X(_01105_));
 sg13g2_xnor2_1 _08093_ (.Y(_01106_),
    .A(_01104_),
    .B(_01105_));
 sg13g2_xor2_1 _08094_ (.B(net1610),
    .A(_01103_),
    .X(_01107_));
 sg13g2_o21ai_1 _08095_ (.B1(_00917_),
    .Y(_01108_),
    .A1(_00918_),
    .A2(_01107_));
 sg13g2_nand2b_1 _08096_ (.Y(_01109_),
    .B(_01108_),
    .A_N(_00908_));
 sg13g2_xor2_1 _08097_ (.B(_01092_),
    .A(net1624),
    .X(_01110_));
 sg13g2_inv_1 _08098_ (.Y(_01111_),
    .A(_01110_));
 sg13g2_xnor2_1 _08099_ (.Y(_01112_),
    .A(_01043_),
    .B(_01110_));
 sg13g2_a21oi_1 _08100_ (.A1(_01089_),
    .A2(_01095_),
    .Y(_01113_),
    .B1(_01094_));
 sg13g2_xnor2_1 _08101_ (.Y(_01114_),
    .A(_01098_),
    .B(_01113_));
 sg13g2_xnor2_1 _08102_ (.Y(_01115_),
    .A(net1611),
    .B(_01114_));
 sg13g2_nor2b_1 _08103_ (.A(_01115_),
    .B_N(_01112_),
    .Y(_01116_));
 sg13g2_a21oi_1 _08104_ (.A1(_01043_),
    .A2(_01111_),
    .Y(_01117_),
    .B1(_01116_));
 sg13g2_xnor2_1 _08105_ (.Y(_01118_),
    .A(_00918_),
    .B(_01107_));
 sg13g2_nor2_1 _08106_ (.A(_01117_),
    .B(_01118_),
    .Y(_01119_));
 sg13g2_xnor2_1 _08107_ (.Y(_01120_),
    .A(_01117_),
    .B(_01118_));
 sg13g2_xnor2_1 _08108_ (.Y(_01121_),
    .A(net1624),
    .B(_01054_));
 sg13g2_nor2_1 _08109_ (.A(_01074_),
    .B(_01121_),
    .Y(_01122_));
 sg13g2_xnor2_1 _08110_ (.Y(_01123_),
    .A(_01074_),
    .B(_01121_));
 sg13g2_xor2_1 _08111_ (.B(_01095_),
    .A(_01089_),
    .X(_01124_));
 sg13g2_xnor2_1 _08112_ (.Y(_01125_),
    .A(net1611),
    .B(_01124_));
 sg13g2_nor2_1 _08113_ (.A(_01123_),
    .B(_01125_),
    .Y(_01126_));
 sg13g2_nor2_2 _08114_ (.A(_01122_),
    .B(_01126_),
    .Y(_01127_));
 sg13g2_xnor2_1 _08115_ (.Y(_01128_),
    .A(_01112_),
    .B(_01115_));
 sg13g2_inv_1 _08116_ (.Y(_01129_),
    .A(_01128_));
 sg13g2_nor2_1 _08117_ (.A(_01127_),
    .B(_01129_),
    .Y(_01130_));
 sg13g2_xnor2_1 _08118_ (.Y(_01131_),
    .A(_01123_),
    .B(_01125_));
 sg13g2_xor2_1 _08119_ (.B(_01048_),
    .A(net1625),
    .X(_01132_));
 sg13g2_nand2b_1 _08120_ (.Y(_01133_),
    .B(_01063_),
    .A_N(_01132_));
 sg13g2_xor2_1 _08121_ (.B(_01132_),
    .A(_01063_),
    .X(_01134_));
 sg13g2_o21ai_1 _08122_ (.B1(_01085_),
    .Y(_01135_),
    .A1(_01033_),
    .A2(_01081_));
 sg13g2_inv_1 _08123_ (.Y(_01136_),
    .A(_01135_));
 sg13g2_o21ai_1 _08124_ (.B1(_01049_),
    .Y(_01137_),
    .A1(_01050_),
    .A2(_01136_));
 sg13g2_xnor2_1 _08125_ (.Y(_01138_),
    .A(_01056_),
    .B(_01137_));
 sg13g2_xnor2_1 _08126_ (.Y(_01139_),
    .A(net1611),
    .B(_01138_));
 sg13g2_o21ai_1 _08127_ (.B1(_01133_),
    .Y(_01140_),
    .A1(_01134_),
    .A2(_01139_));
 sg13g2_nand2b_1 _08128_ (.Y(_01141_),
    .B(_01140_),
    .A_N(_01131_));
 sg13g2_xor2_1 _08129_ (.B(_01140_),
    .A(_01131_),
    .X(_01142_));
 sg13g2_xor2_1 _08130_ (.B(_01026_),
    .A(net1626),
    .X(_01143_));
 sg13g2_nand2b_1 _08131_ (.Y(_01144_),
    .B(_00995_),
    .A_N(_01143_));
 sg13g2_xor2_1 _08132_ (.B(_01143_),
    .A(_00995_),
    .X(_01145_));
 sg13g2_xnor2_1 _08133_ (.Y(_01146_),
    .A(_01033_),
    .B(_01069_));
 sg13g2_xnor2_1 _08134_ (.Y(_01147_),
    .A(net1610),
    .B(_01146_));
 sg13g2_xnor2_1 _08135_ (.Y(_01148_),
    .A(_01145_),
    .B(_01147_));
 sg13g2_xnor2_1 _08136_ (.Y(_01149_),
    .A(net1623),
    .B(_01013_));
 sg13g2_nand2b_1 _08137_ (.Y(_01150_),
    .B(_00931_),
    .A_N(_01149_));
 sg13g2_xor2_1 _08138_ (.B(_01149_),
    .A(_00931_),
    .X(_01151_));
 sg13g2_o21ai_1 _08139_ (.B1(_01016_),
    .Y(_01152_),
    .A1(_01003_),
    .A2(_01015_));
 sg13g2_xor2_1 _08140_ (.B(_01152_),
    .A(_01029_),
    .X(_01153_));
 sg13g2_xnor2_1 _08141_ (.Y(_01154_),
    .A(net1610),
    .B(_01153_));
 sg13g2_o21ai_1 _08142_ (.B1(_01150_),
    .Y(_01155_),
    .A1(_01151_),
    .A2(_01154_));
 sg13g2_nor2b_1 _08143_ (.A(_01148_),
    .B_N(_01155_),
    .Y(_01156_));
 sg13g2_inv_1 _08144_ (.Y(_01157_),
    .A(_01156_));
 sg13g2_xor2_1 _08145_ (.B(_01155_),
    .A(_01148_),
    .X(_01158_));
 sg13g2_o21ai_1 _08146_ (.B1(_01144_),
    .Y(_01159_),
    .A1(_01145_),
    .A2(_01147_));
 sg13g2_xnor2_1 _08147_ (.Y(_01160_),
    .A(net1624),
    .B(_01066_));
 sg13g2_nand2b_1 _08148_ (.Y(_01161_),
    .B(net289),
    .A_N(_01160_));
 sg13g2_xor2_1 _08149_ (.B(_01160_),
    .A(net288),
    .X(_01162_));
 sg13g2_o21ai_1 _08150_ (.B1(_01068_),
    .Y(_01163_),
    .A1(_01033_),
    .A2(_01070_));
 sg13g2_xor2_1 _08151_ (.B(_01163_),
    .A(_01080_),
    .X(_01164_));
 sg13g2_xnor2_1 _08152_ (.Y(_01165_),
    .A(net1610),
    .B(_01164_));
 sg13g2_xor2_1 _08153_ (.B(_01165_),
    .A(_01162_),
    .X(_01166_));
 sg13g2_nor2_1 _08154_ (.A(_01159_),
    .B(_01166_),
    .Y(_01167_));
 sg13g2_xnor2_1 _08155_ (.Y(_01168_),
    .A(_01159_),
    .B(_01166_));
 sg13g2_nor2_1 _08156_ (.A(_01158_),
    .B(_01168_),
    .Y(_01169_));
 sg13g2_or2_1 _08157_ (.X(_01170_),
    .B(_01168_),
    .A(_01158_));
 sg13g2_xnor2_1 _08158_ (.Y(_01171_),
    .A(net1626),
    .B(_00999_));
 sg13g2_inv_1 _08159_ (.Y(_01172_),
    .A(_01171_));
 sg13g2_nand2_1 _08160_ (.Y(_01173_),
    .A(_00941_),
    .B(_01172_));
 sg13g2_xnor2_1 _08161_ (.Y(_01174_),
    .A(_00941_),
    .B(_01171_));
 sg13g2_inv_1 _08162_ (.Y(_01175_),
    .A(_01174_));
 sg13g2_xnor2_1 _08163_ (.Y(_01176_),
    .A(_01003_),
    .B(_01017_));
 sg13g2_xnor2_1 _08164_ (.Y(_01177_),
    .A(net1610),
    .B(_01176_));
 sg13g2_o21ai_1 _08165_ (.B1(_01173_),
    .Y(_01178_),
    .A1(_01175_),
    .A2(_01177_));
 sg13g2_xor2_1 _08166_ (.B(_01154_),
    .A(_01151_),
    .X(_01179_));
 sg13g2_or2_1 _08167_ (.X(_01180_),
    .B(_01179_),
    .A(_01178_));
 sg13g2_and2_1 _08168_ (.A(_01178_),
    .B(_01179_),
    .X(_01181_));
 sg13g2_xnor2_1 _08169_ (.Y(_01182_),
    .A(_01174_),
    .B(_01177_));
 sg13g2_xor2_1 _08170_ (.B(_00936_),
    .A(net1623),
    .X(_01183_));
 sg13g2_nor2_1 _08171_ (.A(_00951_),
    .B(_01183_),
    .Y(_01184_));
 sg13g2_xnor2_1 _08172_ (.Y(_01185_),
    .A(_00952_),
    .B(_01183_));
 sg13g2_nand2_1 _08173_ (.Y(_01186_),
    .A(_00937_),
    .B(_00987_));
 sg13g2_xnor2_1 _08174_ (.Y(_01187_),
    .A(_00996_),
    .B(_00999_));
 sg13g2_xnor2_1 _08175_ (.Y(_01188_),
    .A(_01186_),
    .B(_01187_));
 sg13g2_xnor2_1 _08176_ (.Y(_01189_),
    .A(net1610),
    .B(_01188_));
 sg13g2_a21oi_1 _08177_ (.A1(_01185_),
    .A2(_01189_),
    .Y(_01190_),
    .B1(_01184_));
 sg13g2_nor2b_1 _08178_ (.A(_01190_),
    .B_N(_01182_),
    .Y(_01191_));
 sg13g2_a21o_1 _08179_ (.A2(_01191_),
    .A1(_01180_),
    .B1(_01181_),
    .X(_01192_));
 sg13g2_inv_1 _08180_ (.Y(_01193_),
    .A(_01192_));
 sg13g2_xnor2_1 _08181_ (.Y(_01194_),
    .A(net1623),
    .B(_00946_));
 sg13g2_xnor2_1 _08182_ (.Y(_01195_),
    .A(_00970_),
    .B(_01194_));
 sg13g2_a21o_1 _08183_ (.A2(_00986_),
    .A1(_00948_),
    .B1(_00938_),
    .X(_01196_));
 sg13g2_and2_1 _08184_ (.A(_00987_),
    .B(_01196_),
    .X(_01197_));
 sg13g2_xnor2_1 _08185_ (.Y(_01198_),
    .A(net1610),
    .B(_01197_));
 sg13g2_nand2b_1 _08186_ (.Y(_01199_),
    .B(_01195_),
    .A_N(_01198_));
 sg13g2_xnor2_1 _08187_ (.Y(_01200_),
    .A(_01195_),
    .B(_01198_));
 sg13g2_xnor2_1 _08188_ (.Y(_01201_),
    .A(net1627),
    .B(_00958_));
 sg13g2_inv_1 _08189_ (.Y(_01202_),
    .A(_01201_));
 sg13g2_nand2_1 _08190_ (.Y(_01203_),
    .A(_00978_),
    .B(_01202_));
 sg13g2_nor2_1 _08191_ (.A(_00978_),
    .B(_01202_),
    .Y(_01204_));
 sg13g2_xnor2_1 _08192_ (.Y(_01205_),
    .A(_00978_),
    .B(_01201_));
 sg13g2_nand2b_1 _08193_ (.Y(_01206_),
    .B(_00948_),
    .A_N(_00947_));
 sg13g2_xnor2_1 _08194_ (.Y(_01207_),
    .A(_00985_),
    .B(_01206_));
 sg13g2_xor2_1 _08195_ (.B(_01207_),
    .A(net1612),
    .X(_01208_));
 sg13g2_o21ai_1 _08196_ (.B1(_01203_),
    .Y(_01209_),
    .A1(_01204_),
    .A2(_01208_));
 sg13g2_and2_1 _08197_ (.A(_01200_),
    .B(_01209_),
    .X(_01210_));
 sg13g2_xor2_1 _08198_ (.B(_01209_),
    .A(_01200_),
    .X(_01211_));
 sg13g2_xnor2_1 _08199_ (.Y(_01212_),
    .A(_01205_),
    .B(_01208_));
 sg13g2_xnor2_1 _08200_ (.Y(_01213_),
    .A(net1808),
    .B(_00980_));
 sg13g2_xor2_1 _08201_ (.B(_00967_),
    .A(net1627),
    .X(_01214_));
 sg13g2_nand2_1 _08202_ (.Y(_01215_),
    .A(_01213_),
    .B(_01214_));
 sg13g2_xor2_1 _08203_ (.B(_00983_),
    .A(_00963_),
    .X(_01216_));
 sg13g2_xnor2_1 _08204_ (.Y(_01217_),
    .A(net1612),
    .B(_01216_));
 sg13g2_o21ai_1 _08205_ (.B1(_01217_),
    .Y(_01218_),
    .A1(_01213_),
    .A2(_01214_));
 sg13g2_and3_2 _08206_ (.X(_01219_),
    .A(_01212_),
    .B(_01215_),
    .C(_01218_));
 sg13g2_o21ai_1 _08207_ (.B1(_01199_),
    .Y(_01220_),
    .A1(_00971_),
    .A2(_01194_));
 sg13g2_xor2_1 _08208_ (.B(_01189_),
    .A(_01185_),
    .X(_01221_));
 sg13g2_a221oi_1 _08209_ (.B2(_01221_),
    .C1(_01210_),
    .B1(_01220_),
    .A1(_01219_),
    .Y(_01222_),
    .A2(_01211_));
 sg13g2_nor2_2 _08210_ (.A(_01220_),
    .B(_01221_),
    .Y(_01223_));
 sg13g2_xor2_1 _08211_ (.B(_01179_),
    .A(_01178_),
    .X(_01224_));
 sg13g2_xnor2_1 _08212_ (.Y(_01225_),
    .A(_01182_),
    .B(_01190_));
 sg13g2_inv_1 _08213_ (.Y(_01226_),
    .A(_01225_));
 sg13g2_nand2_1 _08214_ (.Y(_01227_),
    .A(_01224_),
    .B(_01225_));
 sg13g2_or3_1 _08215_ (.A(_01227_),
    .B(_01223_),
    .C(_01222_),
    .X(_01228_));
 sg13g2_nor2b_1 _08216_ (.A(_01167_),
    .B_N(_01156_),
    .Y(_01229_));
 sg13g2_a221oi_1 _08217_ (.B2(_01192_),
    .C1(_01229_),
    .B1(_01169_),
    .A1(_01159_),
    .Y(_01230_),
    .A2(_01166_));
 sg13g2_or4_2 _08218_ (.A(_01170_),
    .B(net272),
    .C(_01223_),
    .D(_01227_),
    .X(_01231_));
 sg13g2_xnor2_1 _08219_ (.Y(_01232_),
    .A(net1624),
    .B(_01077_));
 sg13g2_nand2b_1 _08220_ (.Y(_01233_),
    .B(_01023_),
    .A_N(_01232_));
 sg13g2_xor2_1 _08221_ (.B(_01232_),
    .A(_01023_),
    .X(_01234_));
 sg13g2_xnor2_1 _08222_ (.Y(_01235_),
    .A(_01050_),
    .B(_01135_));
 sg13g2_xnor2_1 _08223_ (.Y(_01236_),
    .A(net1610),
    .B(_01235_));
 sg13g2_o21ai_1 _08224_ (.B1(_01233_),
    .Y(_01237_),
    .A1(_01234_),
    .A2(_01236_));
 sg13g2_xor2_1 _08225_ (.B(_01139_),
    .A(_01134_),
    .X(_01238_));
 sg13g2_nand2_1 _08226_ (.Y(_01239_),
    .A(_01237_),
    .B(_01238_));
 sg13g2_xor2_1 _08227_ (.B(_01238_),
    .A(_01237_),
    .X(_01240_));
 sg13g2_inv_1 _08228_ (.Y(_01241_),
    .A(_01240_));
 sg13g2_xnor2_1 _08229_ (.Y(_01242_),
    .A(_01234_),
    .B(_01236_));
 sg13g2_o21ai_1 _08230_ (.B1(_01161_),
    .Y(_01243_),
    .A1(_01162_),
    .A2(_01165_));
 sg13g2_nor2b_1 _08231_ (.A(_01242_),
    .B_N(_01243_),
    .Y(_01244_));
 sg13g2_xor2_1 _08232_ (.B(_01243_),
    .A(_01242_),
    .X(_01245_));
 sg13g2_or2_1 _08233_ (.X(_01246_),
    .B(_01245_),
    .A(_01241_));
 sg13g2_a21o_1 _08234_ (.A2(_01231_),
    .A1(_01230_),
    .B1(_01246_),
    .X(_01247_));
 sg13g2_o21ai_1 _08235_ (.B1(_01244_),
    .Y(_01248_),
    .A1(_01237_),
    .A2(_01238_));
 sg13g2_and2_1 _08236_ (.A(_01239_),
    .B(_01248_),
    .X(_01249_));
 sg13g2_a21o_2 _08237_ (.A2(_01249_),
    .A1(_01247_),
    .B1(_01142_),
    .X(_01250_));
 sg13g2_nand2_1 _08238_ (.Y(_01251_),
    .A(_01141_),
    .B(_01250_));
 sg13g2_nor2b_1 _08239_ (.A(_01130_),
    .B_N(_01141_),
    .Y(_01252_));
 sg13g2_a22oi_1 _08240_ (.Y(_01253_),
    .B1(_01250_),
    .B2(_01252_),
    .A2(_01129_),
    .A1(_01127_));
 sg13g2_a221oi_1 _08241_ (.B2(_01252_),
    .C1(_01120_),
    .B1(_01250_),
    .A1(_01127_),
    .Y(_01254_),
    .A2(_01129_));
 sg13g2_xor2_1 _08242_ (.B(_01108_),
    .A(_00908_),
    .X(_01255_));
 sg13g2_inv_1 _08243_ (.Y(_01256_),
    .A(_01255_));
 sg13g2_o21ai_1 _08244_ (.B1(_01256_),
    .Y(_01257_),
    .A1(_01119_),
    .A2(_01254_));
 sg13g2_xnor2_1 _08245_ (.Y(_01258_),
    .A(_00904_),
    .B(_00907_));
 sg13g2_a21oi_1 _08246_ (.A1(_01109_),
    .A2(_01257_),
    .Y(_01259_),
    .B1(_01258_));
 sg13g2_a21oi_1 _08247_ (.A1(_00904_),
    .A2(_00907_),
    .Y(_01260_),
    .B1(_01259_));
 sg13g2_xor2_1 _08248_ (.B(_00920_),
    .A(net1807),
    .X(_01261_));
 sg13g2_xnor2_1 _08249_ (.Y(_01262_),
    .A(_01260_),
    .B(_01261_));
 sg13g2_nand3_1 _08250_ (.B(_01257_),
    .C(_01258_),
    .A(_01109_),
    .Y(_01263_));
 sg13g2_nand2b_2 _08251_ (.Y(_01264_),
    .B(_01263_),
    .A_N(_01259_));
 sg13g2_inv_1 _08252_ (.Y(_01265_),
    .A(_01264_));
 sg13g2_xnor2_1 _08253_ (.Y(_01266_),
    .A(_01120_),
    .B(_01253_));
 sg13g2_nor2_1 _08254_ (.A(_01265_),
    .B(_01266_),
    .Y(_01267_));
 sg13g2_or3_1 _08255_ (.A(_01119_),
    .B(_01254_),
    .C(_01256_),
    .X(_01268_));
 sg13g2_and2_2 _08256_ (.A(_01257_),
    .B(_01268_),
    .X(_01269_));
 sg13g2_nor2b_1 _08257_ (.A(_01262_),
    .B_N(_01269_),
    .Y(_01270_));
 sg13g2_xnor2_1 _08258_ (.Y(_01271_),
    .A(_01262_),
    .B(_01269_));
 sg13g2_nand2b_1 _08259_ (.Y(_01272_),
    .B(_01271_),
    .A_N(_01267_));
 sg13g2_nor2b_1 _08260_ (.A(_01271_),
    .B_N(_01267_),
    .Y(_01273_));
 sg13g2_xnor2_1 _08261_ (.Y(_01274_),
    .A(_01267_),
    .B(_01271_));
 sg13g2_xnor2_1 _08262_ (.Y(_01275_),
    .A(_01127_),
    .B(_01128_));
 sg13g2_xnor2_1 _08263_ (.Y(_01276_),
    .A(_01251_),
    .B(_01275_));
 sg13g2_nor2b_1 _08264_ (.A(_01269_),
    .B_N(_01276_),
    .Y(_01277_));
 sg13g2_xnor2_1 _08265_ (.Y(_01278_),
    .A(_01264_),
    .B(_01266_));
 sg13g2_nand2_1 _08266_ (.Y(_01279_),
    .A(_01277_),
    .B(_01278_));
 sg13g2_nand3_1 _08267_ (.B(_01247_),
    .C(_01249_),
    .A(_01142_),
    .Y(_01280_));
 sg13g2_and2_1 _08268_ (.A(_01250_),
    .B(_01280_),
    .X(_01281_));
 sg13g2_nor2_1 _08269_ (.A(_01266_),
    .B(_01281_),
    .Y(_01282_));
 sg13g2_xnor2_1 _08270_ (.Y(_01283_),
    .A(_01269_),
    .B(_01276_));
 sg13g2_nor2_1 _08271_ (.A(_01282_),
    .B(_01283_),
    .Y(_01284_));
 sg13g2_or2_1 _08272_ (.X(_01285_),
    .B(_01283_),
    .A(_01282_));
 sg13g2_xnor2_1 _08273_ (.Y(_01286_),
    .A(_01282_),
    .B(_01283_));
 sg13g2_a21oi_2 _08274_ (.B1(_01245_),
    .Y(_01287_),
    .A2(_01231_),
    .A1(_01230_));
 sg13g2_o21ai_1 _08275_ (.B1(_01240_),
    .Y(_01288_),
    .A1(_01244_),
    .A2(_01287_));
 sg13g2_or3_1 _08276_ (.A(_01240_),
    .B(_01244_),
    .C(_01287_),
    .X(_01289_));
 sg13g2_and2_2 _08277_ (.A(_01288_),
    .B(_01289_),
    .X(_01290_));
 sg13g2_nand2b_2 _08278_ (.Y(_01291_),
    .B(_01290_),
    .A_N(_01276_));
 sg13g2_xor2_1 _08279_ (.B(_01281_),
    .A(_01266_),
    .X(_01292_));
 sg13g2_a21o_1 _08280_ (.A2(_01228_),
    .A1(_01193_),
    .B1(_01158_),
    .X(_01293_));
 sg13g2_a21o_1 _08281_ (.A2(_01157_),
    .A1(_01293_),
    .B1(_01168_),
    .X(_01294_));
 sg13g2_nand3_1 _08282_ (.B(_01168_),
    .C(_01293_),
    .A(_01157_),
    .Y(_01295_));
 sg13g2_nand2_1 _08283_ (.Y(_01296_),
    .A(_01294_),
    .B(_01295_));
 sg13g2_nand4_1 _08284_ (.B(_01289_),
    .C(_01294_),
    .A(_01288_),
    .Y(_01297_),
    .D(_01295_));
 sg13g2_nand3_1 _08285_ (.B(_01231_),
    .C(_01245_),
    .A(_01230_),
    .Y(_01298_));
 sg13g2_nor2b_2 _08286_ (.A(_01287_),
    .B_N(_01298_),
    .Y(_01299_));
 sg13g2_and3_1 _08287_ (.X(_01300_),
    .A(_01250_),
    .B(_01280_),
    .C(_01299_));
 sg13g2_nand2_1 _08288_ (.Y(_01301_),
    .A(_01281_),
    .B(_01299_));
 sg13g2_a21oi_1 _08289_ (.A1(_01250_),
    .A2(_01280_),
    .Y(_01302_),
    .B1(_01299_));
 sg13g2_o21ai_1 _08290_ (.B1(_01297_),
    .Y(_01303_),
    .A1(_01300_),
    .A2(_01302_));
 sg13g2_nor3_1 _08291_ (.A(_01297_),
    .B(_01300_),
    .C(_01302_),
    .Y(_01304_));
 sg13g2_or3_1 _08292_ (.A(_01297_),
    .B(_01300_),
    .C(_01302_),
    .X(_01305_));
 sg13g2_nand3_1 _08293_ (.B(_01193_),
    .C(_01228_),
    .A(_01158_),
    .Y(_01306_));
 sg13g2_nand2_2 _08294_ (.Y(_01307_),
    .A(_01293_),
    .B(_01306_));
 sg13g2_and3_1 _08295_ (.X(_01308_),
    .A(_01293_),
    .B(_01299_),
    .C(_01306_));
 sg13g2_xnor2_1 _08296_ (.Y(_01309_),
    .A(_01290_),
    .B(_01296_));
 sg13g2_nand2_1 _08297_ (.Y(_01310_),
    .A(_01308_),
    .B(_01309_));
 sg13g2_nand3_1 _08298_ (.B(_01308_),
    .C(_01309_),
    .A(_01303_),
    .Y(_01311_));
 sg13g2_nor3_2 _08299_ (.A(_01226_),
    .B(_01223_),
    .C(_01222_),
    .Y(_01312_));
 sg13g2_or3_1 _08300_ (.A(_01222_),
    .B(_01223_),
    .C(_01226_),
    .X(_01313_));
 sg13g2_o21ai_1 _08301_ (.B1(_01224_),
    .Y(_01314_),
    .A1(_01312_),
    .A2(_01191_));
 sg13g2_or3_2 _08302_ (.A(_01191_),
    .B(_01224_),
    .C(_01312_),
    .X(_01315_));
 sg13g2_and2_1 _08303_ (.A(_01314_),
    .B(_01315_),
    .X(_01316_));
 sg13g2_nand3_1 _08304_ (.B(_01295_),
    .C(_01316_),
    .A(_01294_),
    .Y(_01317_));
 sg13g2_xor2_1 _08305_ (.B(_01299_),
    .A(_01307_),
    .X(_01318_));
 sg13g2_nor2_1 _08306_ (.A(_01317_),
    .B(_01318_),
    .Y(_01319_));
 sg13g2_nand2_1 _08307_ (.Y(_01320_),
    .A(_01317_),
    .B(_01318_));
 sg13g2_o21ai_1 _08308_ (.B1(_01226_),
    .Y(_01321_),
    .A1(_01222_),
    .A2(_01223_));
 sg13g2_and2_1 _08309_ (.A(_01313_),
    .B(_01321_),
    .X(_01322_));
 sg13g2_nor2b_1 _08310_ (.A(_01307_),
    .B_N(_01322_),
    .Y(_01323_));
 sg13g2_a21o_1 _08311_ (.A2(_01295_),
    .A1(_01294_),
    .B1(_01316_),
    .X(_01324_));
 sg13g2_and3_1 _08312_ (.X(_01325_),
    .A(net1444),
    .B(_01323_),
    .C(_01324_));
 sg13g2_nand3_1 _08313_ (.B(_01323_),
    .C(_01324_),
    .A(net273),
    .Y(_01326_));
 sg13g2_xor2_1 _08314_ (.B(_01221_),
    .A(_01220_),
    .X(_01327_));
 sg13g2_a21oi_1 _08315_ (.A1(_01211_),
    .A2(_01219_),
    .Y(_01328_),
    .B1(_01210_));
 sg13g2_xnor2_1 _08316_ (.Y(_01329_),
    .A(_01327_),
    .B(_01328_));
 sg13g2_and3_1 _08317_ (.X(_01330_),
    .A(_01314_),
    .B(_01315_),
    .C(_01329_));
 sg13g2_nand3_1 _08318_ (.B(_01315_),
    .C(_01329_),
    .A(_01314_),
    .Y(_01331_));
 sg13g2_a21oi_1 _08319_ (.A1(_01314_),
    .A2(_01315_),
    .Y(_01332_),
    .B1(_01329_));
 sg13g2_a21o_1 _08320_ (.A2(_01315_),
    .A1(_01314_),
    .B1(_01329_),
    .X(_01333_));
 sg13g2_xnor2_1 _08321_ (.Y(_01334_),
    .A(_01211_),
    .B(_01219_));
 sg13g2_inv_1 _08322_ (.Y(_01335_),
    .A(_01334_));
 sg13g2_and3_1 _08323_ (.X(_01336_),
    .A(_01313_),
    .B(_01321_),
    .C(_01335_));
 sg13g2_a21oi_1 _08324_ (.A1(_01313_),
    .A2(_01321_),
    .Y(_01337_),
    .B1(_01335_));
 sg13g2_a21o_1 _08325_ (.A2(_01321_),
    .A1(_01313_),
    .B1(_01335_),
    .X(_01338_));
 sg13g2_a21oi_1 _08326_ (.A1(_01215_),
    .A2(_01218_),
    .Y(_01339_),
    .B1(_01212_));
 sg13g2_nor2_2 _08327_ (.A(_01219_),
    .B(_01339_),
    .Y(_01340_));
 sg13g2_and2_1 _08328_ (.A(_01329_),
    .B(_01340_),
    .X(_01341_));
 sg13g2_nand2_1 _08329_ (.Y(_01342_),
    .A(_01329_),
    .B(_01340_));
 sg13g2_nand3b_1 _08330_ (.B(_01338_),
    .C(_01341_),
    .Y(_01343_),
    .A_N(_01336_));
 sg13g2_a21oi_1 _08331_ (.A1(_01338_),
    .A2(_01341_),
    .Y(_01344_),
    .B1(_01336_));
 sg13g2_nor3_2 _08332_ (.A(_01330_),
    .B(_01332_),
    .C(_01344_),
    .Y(_01345_));
 sg13g2_o21ai_1 _08333_ (.B1(_01331_),
    .Y(_01346_),
    .A1(_01332_),
    .A2(_01344_));
 sg13g2_xnor2_1 _08334_ (.Y(_01347_),
    .A(_01307_),
    .B(_01322_));
 sg13g2_and2_1 _08335_ (.A(_01346_),
    .B(_01347_),
    .X(_01348_));
 sg13g2_nand2_1 _08336_ (.Y(_01349_),
    .A(_01346_),
    .B(_01347_));
 sg13g2_a21oi_1 _08337_ (.A1(_01317_),
    .A2(_01324_),
    .Y(_01350_),
    .B1(_01323_));
 sg13g2_a21o_1 _08338_ (.A2(_01324_),
    .A1(net273),
    .B1(_01323_),
    .X(_01351_));
 sg13g2_nor3_2 _08339_ (.A(_01325_),
    .B(_01349_),
    .C(_01350_),
    .Y(_01352_));
 sg13g2_o21ai_1 _08340_ (.B1(_01326_),
    .Y(_01353_),
    .A1(_01349_),
    .A2(_01350_));
 sg13g2_xor2_1 _08341_ (.B(_01318_),
    .A(_01317_),
    .X(_01354_));
 sg13g2_nand4_1 _08342_ (.B(_01348_),
    .C(_01351_),
    .A(_01354_),
    .Y(_01355_),
    .D(_01326_));
 sg13g2_a21oi_1 _08343_ (.A1(_01320_),
    .A2(_01325_),
    .Y(_01356_),
    .B1(_01319_));
 sg13g2_and2_1 _08344_ (.A(_01355_),
    .B(_01356_),
    .X(_01357_));
 sg13g2_nand4_1 _08345_ (.B(_01311_),
    .C(_01305_),
    .A(_01355_),
    .Y(_01358_),
    .D(_01356_));
 sg13g2_or3_1 _08346_ (.A(_01304_),
    .B(_01308_),
    .C(_01309_),
    .X(_01359_));
 sg13g2_and2_1 _08347_ (.A(_01303_),
    .B(_01359_),
    .X(_01360_));
 sg13g2_xor2_1 _08348_ (.B(_01290_),
    .A(_01276_),
    .X(_01361_));
 sg13g2_nor2_1 _08349_ (.A(_01301_),
    .B(_01361_),
    .Y(_01362_));
 sg13g2_xnor2_1 _08350_ (.Y(_01363_),
    .A(_01300_),
    .B(_01361_));
 sg13g2_nand3_1 _08351_ (.B(_01358_),
    .C(_01363_),
    .A(_01360_),
    .Y(_01364_));
 sg13g2_nor2_1 _08352_ (.A(_01291_),
    .B(_01292_),
    .Y(_01365_));
 sg13g2_nor2_1 _08353_ (.A(_01362_),
    .B(_01365_),
    .Y(_01366_));
 sg13g2_xnor2_1 _08354_ (.Y(_01367_),
    .A(_01291_),
    .B(_01292_));
 sg13g2_a22oi_1 _08355_ (.Y(_01368_),
    .B1(_01364_),
    .B2(_01366_),
    .A2(_01292_),
    .A1(_01291_));
 sg13g2_a221oi_1 _08356_ (.B2(_01364_),
    .C1(_01286_),
    .B1(_01366_),
    .A1(_01291_),
    .Y(_01369_),
    .A2(_01292_));
 sg13g2_o21ai_1 _08357_ (.B1(_01285_),
    .Y(_01370_),
    .A1(_01277_),
    .A2(_01278_));
 sg13g2_o21ai_1 _08358_ (.B1(_01279_),
    .Y(_01371_),
    .A1(_01370_),
    .A2(_01369_));
 sg13g2_o21ai_1 _08359_ (.B1(_01272_),
    .Y(_01372_),
    .A1(_01371_),
    .A2(_01273_));
 sg13g2_nand2b_1 _08360_ (.Y(_01373_),
    .B(_01264_),
    .A_N(_01262_));
 sg13g2_nand2_1 _08361_ (.Y(_01374_),
    .A(_01262_),
    .B(_01265_));
 sg13g2_xnor2_1 _08362_ (.Y(_01375_),
    .A(_01265_),
    .B(_01270_));
 sg13g2_or3_1 _08363_ (.A(_01269_),
    .B(_01373_),
    .C(_01372_),
    .X(_01376_));
 sg13g2_nor2b_2 _08364_ (.A(_01262_),
    .B_N(_01376_),
    .Y(_01377_));
 sg13g2_xnor2_1 _08365_ (.Y(_01378_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[15] ),
    .B(_01377_));
 sg13g2_xor2_1 _08366_ (.B(net1596),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[15] ),
    .X(_01379_));
 sg13g2_xor2_1 _08367_ (.B(_01368_),
    .A(_01286_),
    .X(_01380_));
 sg13g2_nor2_1 _08368_ (.A(_00627_),
    .B(_01380_),
    .Y(_01381_));
 sg13g2_nand2_1 _08369_ (.Y(_01382_),
    .A(_00627_),
    .B(_01380_));
 sg13g2_xnor2_1 _08370_ (.Y(_01383_),
    .A(_00627_),
    .B(_01380_));
 sg13g2_nand2b_1 _08371_ (.Y(_01384_),
    .B(_01364_),
    .A_N(_01362_));
 sg13g2_xor2_1 _08372_ (.B(_01384_),
    .A(_01367_),
    .X(_01385_));
 sg13g2_nor2b_1 _08373_ (.A(_00145_),
    .B_N(_01385_),
    .Y(_01386_));
 sg13g2_nand2b_1 _08374_ (.Y(_01387_),
    .B(_00145_),
    .A_N(_01385_));
 sg13g2_a21o_1 _08375_ (.A2(_01360_),
    .A1(_01358_),
    .B1(_01363_),
    .X(_01388_));
 sg13g2_and2_2 _08376_ (.A(_01364_),
    .B(_01388_),
    .X(_01389_));
 sg13g2_nand2_1 _08377_ (.Y(_01390_),
    .A(_00146_),
    .B(_01389_));
 sg13g2_xnor2_1 _08378_ (.Y(_01391_),
    .A(_00146_),
    .B(_01389_));
 sg13g2_inv_1 _08379_ (.Y(_01392_),
    .A(_01391_));
 sg13g2_nand2_2 _08380_ (.Y(_01393_),
    .A(_01303_),
    .B(_01305_));
 sg13g2_xnor2_1 _08381_ (.Y(_01394_),
    .A(_01308_),
    .B(_01309_));
 sg13g2_o21ai_1 _08382_ (.B1(_01310_),
    .Y(_01395_),
    .A1(_01357_),
    .A2(_01394_));
 sg13g2_xnor2_1 _08383_ (.Y(_01396_),
    .A(_01393_),
    .B(_01395_));
 sg13g2_xor2_1 _08384_ (.B(_01395_),
    .A(_01393_),
    .X(_01397_));
 sg13g2_nand2_1 _08385_ (.Y(_01398_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[7] ),
    .B(_01397_));
 sg13g2_xnor2_1 _08386_ (.Y(_01399_),
    .A(_01357_),
    .B(_01394_));
 sg13g2_nor2_1 _08387_ (.A(_00630_),
    .B(_01399_),
    .Y(_01400_));
 sg13g2_xnor2_1 _08388_ (.Y(_01401_),
    .A(_01353_),
    .B(_01354_));
 sg13g2_or2_1 _08389_ (.X(_01402_),
    .B(_01401_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[5] ));
 sg13g2_or2_1 _08390_ (.X(_01403_),
    .B(_01401_),
    .A(_00149_));
 sg13g2_xor2_1 _08391_ (.B(_01401_),
    .A(_00149_),
    .X(_01404_));
 sg13g2_a21oi_2 _08392_ (.B1(_01348_),
    .Y(_01405_),
    .A2(_01351_),
    .A1(_01326_));
 sg13g2_nor3_1 _08393_ (.A(_00632_),
    .B(_01352_),
    .C(_01405_),
    .Y(_01406_));
 sg13g2_xnor2_1 _08394_ (.Y(_01407_),
    .A(_01346_),
    .B(_01347_));
 sg13g2_or2_1 _08395_ (.X(_01408_),
    .B(_01407_),
    .A(_00151_));
 sg13g2_xor2_1 _08396_ (.B(_01407_),
    .A(_00151_),
    .X(_01409_));
 sg13g2_a221oi_1 _08397_ (.B2(_01341_),
    .C1(_01336_),
    .B1(_01338_),
    .A1(_01331_),
    .Y(_01410_),
    .A2(_01333_));
 sg13g2_nor3_1 _08398_ (.A(_00633_),
    .B(_01345_),
    .C(_01410_),
    .Y(_01411_));
 sg13g2_o21ai_1 _08399_ (.B1(_01342_),
    .Y(_01412_),
    .A1(_01336_),
    .A2(_01337_));
 sg13g2_and3_1 _08400_ (.X(_01413_),
    .A(_00634_),
    .B(_01343_),
    .C(_01412_));
 sg13g2_nand3_1 _08401_ (.B(_01343_),
    .C(_01412_),
    .A(_00634_),
    .Y(_01414_));
 sg13g2_a21oi_1 _08402_ (.A1(_01343_),
    .A2(_01412_),
    .Y(_01415_),
    .B1(_00634_));
 sg13g2_nor2_1 _08403_ (.A(_01413_),
    .B(_01415_),
    .Y(_01416_));
 sg13g2_xor2_1 _08404_ (.B(_01340_),
    .A(_01329_),
    .X(_01417_));
 sg13g2_nor2_1 _08405_ (.A(_00154_),
    .B(_01417_),
    .Y(_01418_));
 sg13g2_o21ai_1 _08406_ (.B1(_01414_),
    .Y(_01419_),
    .A1(_01415_),
    .A2(_01418_));
 sg13g2_nor3_1 _08407_ (.A(_00152_),
    .B(_01345_),
    .C(_01410_),
    .Y(_01420_));
 sg13g2_o21ai_1 _08408_ (.B1(_00633_),
    .Y(_01421_),
    .A1(_01345_),
    .A2(_01410_));
 sg13g2_nand2b_1 _08409_ (.Y(_01422_),
    .B(_01421_),
    .A_N(_01411_));
 sg13g2_a21oi_1 _08410_ (.A1(_01419_),
    .A2(_01421_),
    .Y(_01423_),
    .B1(_01411_));
 sg13g2_or2_1 _08411_ (.X(_01424_),
    .B(_01407_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[3] ));
 sg13g2_o21ai_1 _08412_ (.B1(_01424_),
    .Y(_01425_),
    .A1(_01409_),
    .A2(_01423_));
 sg13g2_o21ai_1 _08413_ (.B1(_00632_),
    .Y(_01426_),
    .A1(_01352_),
    .A2(_01405_));
 sg13g2_nand2b_1 _08414_ (.Y(_01427_),
    .B(_01426_),
    .A_N(_01406_));
 sg13g2_a21oi_1 _08415_ (.A1(_01425_),
    .A2(_01426_),
    .Y(_01428_),
    .B1(_01406_));
 sg13g2_o21ai_1 _08416_ (.B1(_01402_),
    .Y(_01429_),
    .A1(_01404_),
    .A2(_01428_));
 sg13g2_nor2_1 _08417_ (.A(_00148_),
    .B(_01399_),
    .Y(_01430_));
 sg13g2_inv_1 _08418_ (.Y(_01431_),
    .A(_01430_));
 sg13g2_xnor2_1 _08419_ (.Y(_01432_),
    .A(_00148_),
    .B(_01399_));
 sg13g2_a21oi_1 _08420_ (.A1(_01429_),
    .A2(_01432_),
    .Y(_01433_),
    .B1(_01400_));
 sg13g2_a221oi_1 _08421_ (.B2(_01432_),
    .C1(_01400_),
    .B1(_01429_),
    .A1(_00629_),
    .Y(_01434_),
    .A2(_01396_));
 sg13g2_inv_1 _08422_ (.Y(_01435_),
    .A(_01434_));
 sg13g2_and3_1 _08423_ (.X(_01436_),
    .A(_01392_),
    .B(_01398_),
    .C(_01435_));
 sg13g2_nand3_1 _08424_ (.B(_01398_),
    .C(_01435_),
    .A(_01392_),
    .Y(_01437_));
 sg13g2_a21oi_1 _08425_ (.A1(_01387_),
    .A2(_01390_),
    .Y(_01438_),
    .B1(_01386_));
 sg13g2_nor2b_2 _08426_ (.A(_01386_),
    .B_N(_01387_),
    .Y(_01439_));
 sg13g2_a21o_1 _08427_ (.A2(_01439_),
    .A1(_01436_),
    .B1(_01438_),
    .X(_01440_));
 sg13g2_xnor2_1 _08428_ (.Y(_01441_),
    .A(_01383_),
    .B(_01440_));
 sg13g2_nand2b_1 _08429_ (.Y(_01442_),
    .B(_01389_),
    .A_N(_00146_));
 sg13g2_nor2_1 _08430_ (.A(_00147_),
    .B(_01397_),
    .Y(_01443_));
 sg13g2_nand2_1 _08431_ (.Y(_01444_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[0] ),
    .B(_01417_));
 sg13g2_inv_1 _08432_ (.Y(_01445_),
    .A(_01444_));
 sg13g2_o21ai_1 _08433_ (.B1(_01445_),
    .Y(_01446_),
    .A1(_01413_),
    .A2(_01415_));
 sg13g2_nand3_1 _08434_ (.B(_01343_),
    .C(_01412_),
    .A(_00635_),
    .Y(_01447_));
 sg13g2_o21ai_1 _08435_ (.B1(\vgadonut.donut.donuthit.cordicxz.xin[2] ),
    .Y(_01448_),
    .A1(_01345_),
    .A2(_01410_));
 sg13g2_or3_1 _08436_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[2] ),
    .B(_01345_),
    .C(_01410_),
    .X(_01449_));
 sg13g2_a22oi_1 _08437_ (.Y(_01450_),
    .B1(_01448_),
    .B2(_01449_),
    .A2(_01447_),
    .A1(_01446_));
 sg13g2_nor2_1 _08438_ (.A(_01420_),
    .B(_01450_),
    .Y(_01451_));
 sg13g2_o21ai_1 _08439_ (.B1(_01409_),
    .Y(_01452_),
    .A1(_01420_),
    .A2(_01450_));
 sg13g2_nand2_1 _08440_ (.Y(_01453_),
    .A(_01408_),
    .B(_01452_));
 sg13g2_o21ai_1 _08441_ (.B1(\vgadonut.donut.donuthit.cordicxz.xin[4] ),
    .Y(_01454_),
    .A1(_01352_),
    .A2(_01405_));
 sg13g2_or3_1 _08442_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[4] ),
    .B(_01352_),
    .C(_01405_),
    .X(_01455_));
 sg13g2_and2_1 _08443_ (.A(_01454_),
    .B(_01455_),
    .X(_01456_));
 sg13g2_a22oi_1 _08444_ (.Y(_01457_),
    .B1(_01454_),
    .B2(_01455_),
    .A2(_01452_),
    .A1(_01408_));
 sg13g2_nor3_1 _08445_ (.A(_00150_),
    .B(_01352_),
    .C(_01405_),
    .Y(_01458_));
 sg13g2_nor2_1 _08446_ (.A(_01457_),
    .B(_01458_),
    .Y(_01459_));
 sg13g2_o21ai_1 _08447_ (.B1(_01404_),
    .Y(_01460_),
    .A1(_01457_),
    .A2(_01458_));
 sg13g2_xor2_1 _08448_ (.B(_01399_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[6] ),
    .X(_01461_));
 sg13g2_a21o_1 _08449_ (.A2(_01460_),
    .A1(_01403_),
    .B1(_01461_),
    .X(_01462_));
 sg13g2_nand2_1 _08450_ (.Y(_01463_),
    .A(_01431_),
    .B(_01462_));
 sg13g2_xnor2_1 _08451_ (.Y(_01464_),
    .A(_00147_),
    .B(_01397_));
 sg13g2_a21oi_1 _08452_ (.A1(_01431_),
    .A2(_01462_),
    .Y(_01465_),
    .B1(_01464_));
 sg13g2_nor2_1 _08453_ (.A(_01443_),
    .B(_01465_),
    .Y(_01466_));
 sg13g2_o21ai_1 _08454_ (.B1(_01391_),
    .Y(_01467_),
    .A1(_01443_),
    .A2(_01465_));
 sg13g2_a21o_1 _08455_ (.A2(_01467_),
    .A1(_01442_),
    .B1(_01439_),
    .X(_01468_));
 sg13g2_o21ai_1 _08456_ (.B1(_01468_),
    .Y(_01469_),
    .A1(_00628_),
    .A2(_01385_));
 sg13g2_xor2_1 _08457_ (.B(_01380_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[10] ),
    .X(_01470_));
 sg13g2_inv_1 _08458_ (.Y(_01471_),
    .A(_01470_));
 sg13g2_xnor2_1 _08459_ (.Y(_01472_),
    .A(_01469_),
    .B(_01470_));
 sg13g2_mux2_1 _08460_ (.A0(_01441_),
    .A1(_01472_),
    .S(net1578),
    .X(_01473_));
 sg13g2_xor2_1 _08461_ (.B(_01473_),
    .A(net1596),
    .X(_01474_));
 sg13g2_nand3_1 _08462_ (.B(_01373_),
    .C(_01375_),
    .A(_01372_),
    .Y(_01475_));
 sg13g2_and3_2 _08463_ (.X(_01476_),
    .A(_01374_),
    .B(_01376_),
    .C(_01475_));
 sg13g2_nor2_1 _08464_ (.A(_00158_),
    .B(_01476_),
    .Y(_01477_));
 sg13g2_xor2_1 _08465_ (.B(_01372_),
    .A(_01375_),
    .X(_01478_));
 sg13g2_nand2b_1 _08466_ (.Y(_01479_),
    .B(net299),
    .A_N(\vgadonut.donut.donuthit.cordicxz.xin[13] ));
 sg13g2_xnor2_1 _08467_ (.Y(_01480_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[13] ),
    .B(net299));
 sg13g2_xor2_1 _08468_ (.B(_01278_),
    .A(_01277_),
    .X(_01481_));
 sg13g2_or3_2 _08469_ (.A(_01284_),
    .B(_01369_),
    .C(_01481_),
    .X(_01482_));
 sg13g2_o21ai_1 _08470_ (.B1(_01481_),
    .Y(_01483_),
    .A1(_01284_),
    .A2(_01369_));
 sg13g2_nand2_1 _08471_ (.Y(_01484_),
    .A(_01482_),
    .B(_01483_));
 sg13g2_a21o_1 _08472_ (.A2(_01483_),
    .A1(_01482_),
    .B1(_00626_),
    .X(_01485_));
 sg13g2_nor2_1 _08473_ (.A(_00143_),
    .B(_01484_),
    .Y(_01486_));
 sg13g2_nand3_1 _08474_ (.B(_01482_),
    .C(_01483_),
    .A(_00626_),
    .Y(_01487_));
 sg13g2_nand2b_1 _08475_ (.Y(_01488_),
    .B(_00627_),
    .A_N(_01380_));
 sg13g2_inv_1 _08476_ (.Y(_01489_),
    .A(_01488_));
 sg13g2_a21oi_1 _08477_ (.A1(_01469_),
    .A2(_01471_),
    .Y(_01490_),
    .B1(_01489_));
 sg13g2_and2_1 _08478_ (.A(_01485_),
    .B(_01487_),
    .X(_01491_));
 sg13g2_nand2_1 _08479_ (.Y(_01492_),
    .A(_01485_),
    .B(_01487_));
 sg13g2_nor2_1 _08480_ (.A(_01470_),
    .B(_01492_),
    .Y(_01493_));
 sg13g2_a221oi_1 _08481_ (.B2(_01469_),
    .C1(_01486_),
    .B1(_01493_),
    .A1(_01485_),
    .Y(_01494_),
    .A2(_01489_));
 sg13g2_xnor2_1 _08482_ (.Y(_01495_),
    .A(_01274_),
    .B(_01371_));
 sg13g2_nand2_1 _08483_ (.Y(_01496_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[12] ),
    .B(_01495_));
 sg13g2_xnor2_1 _08484_ (.Y(_01497_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[12] ),
    .B(_01495_));
 sg13g2_or2_1 _08485_ (.X(_01498_),
    .B(_01497_),
    .A(_01480_));
 sg13g2_nand2_1 _08486_ (.Y(_01499_),
    .A(_00636_),
    .B(net299));
 sg13g2_nor2_1 _08487_ (.A(_01480_),
    .B(_01496_),
    .Y(_01500_));
 sg13g2_a21oi_1 _08488_ (.A1(_00636_),
    .A2(net299),
    .Y(_01501_),
    .B1(_01500_));
 sg13g2_o21ai_1 _08489_ (.B1(_01501_),
    .Y(_01502_),
    .A1(_01494_),
    .A2(_01498_));
 sg13g2_xnor2_1 _08490_ (.Y(_01503_),
    .A(_00158_),
    .B(_01476_));
 sg13g2_inv_1 _08491_ (.Y(_01504_),
    .A(_01503_));
 sg13g2_a21oi_2 _08492_ (.B1(_01477_),
    .Y(_01505_),
    .A2(_01504_),
    .A1(_01502_));
 sg13g2_a21o_2 _08493_ (.A2(_01504_),
    .A1(_01502_),
    .B1(_01477_),
    .X(_01506_));
 sg13g2_or2_1 _08494_ (.X(_01507_),
    .B(_01476_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[14] ));
 sg13g2_nor2_1 _08495_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[11] ),
    .B(_01484_),
    .Y(_01508_));
 sg13g2_a21o_1 _08496_ (.A2(_01440_),
    .A1(_01382_),
    .B1(_01381_),
    .X(_01509_));
 sg13g2_a21oi_1 _08497_ (.A1(_01485_),
    .A2(_01487_),
    .Y(_01510_),
    .B1(_01383_));
 sg13g2_nand3_1 _08498_ (.B(_01439_),
    .C(_01510_),
    .A(_01436_),
    .Y(_01511_));
 sg13g2_a221oi_1 _08499_ (.B2(_01438_),
    .C1(_01508_),
    .B1(_01510_),
    .A1(_01381_),
    .Y(_01512_),
    .A2(_01492_));
 sg13g2_and2_1 _08500_ (.A(_01511_),
    .B(_01512_),
    .X(_01513_));
 sg13g2_nand2b_1 _08501_ (.Y(_01514_),
    .B(_00157_),
    .A_N(net299));
 sg13g2_xnor2_1 _08502_ (.Y(_01515_),
    .A(net299),
    .B(_00157_));
 sg13g2_nand2_1 _08503_ (.Y(_01516_),
    .A(_00155_),
    .B(_01495_));
 sg13g2_xnor2_1 _08504_ (.Y(_01517_),
    .A(_00155_),
    .B(_01495_));
 sg13g2_a221oi_1 _08505_ (.B2(_01499_),
    .C1(_01517_),
    .B1(_01514_),
    .A1(_01511_),
    .Y(_01518_),
    .A2(_01512_));
 sg13g2_o21ai_1 _08506_ (.B1(_01479_),
    .Y(_01519_),
    .A1(_01515_),
    .A2(_01516_));
 sg13g2_xor2_1 _08507_ (.B(_01476_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[14] ),
    .X(_01520_));
 sg13g2_o21ai_1 _08508_ (.B1(_01520_),
    .Y(_01521_),
    .A1(_01519_),
    .A2(_01518_));
 sg13g2_xor2_1 _08509_ (.B(net1596),
    .A(_00156_),
    .X(_01522_));
 sg13g2_and3_1 _08510_ (.X(_01523_),
    .A(_01507_),
    .B(_01521_),
    .C(_01522_));
 sg13g2_nand3_1 _08511_ (.B(_01521_),
    .C(_01522_),
    .A(_01507_),
    .Y(_01524_));
 sg13g2_a21oi_1 _08512_ (.A1(_01507_),
    .A2(_01521_),
    .Y(_01525_),
    .B1(_01522_));
 sg13g2_a21o_1 _08513_ (.A2(_01507_),
    .A1(_01521_),
    .B1(_01522_),
    .X(_01526_));
 sg13g2_nor3_2 _08514_ (.A(net1590),
    .B(_01523_),
    .C(_01525_),
    .Y(_01527_));
 sg13g2_a21oi_2 _08515_ (.B1(net1589),
    .Y(_01528_),
    .A2(_01526_),
    .A1(_01524_));
 sg13g2_a21oi_2 _08516_ (.B1(_01527_),
    .Y(_01529_),
    .A2(_01505_),
    .A1(net1587));
 sg13g2_a21oi_2 _08517_ (.B1(_01528_),
    .Y(_01530_),
    .A2(_01506_),
    .A1(net1587));
 sg13g2_xnor2_1 _08518_ (.Y(_01531_),
    .A(_01491_),
    .B(_01509_));
 sg13g2_and2_1 _08519_ (.A(net1580),
    .B(_01531_),
    .X(_01532_));
 sg13g2_xnor2_1 _08520_ (.Y(_01533_),
    .A(_01490_),
    .B(_01491_));
 sg13g2_a21oi_1 _08521_ (.A1(net1589),
    .A2(_01533_),
    .Y(_01534_),
    .B1(_01532_));
 sg13g2_xnor2_1 _08522_ (.Y(_01535_),
    .A(net1550),
    .B(_01534_));
 sg13g2_inv_1 _08523_ (.Y(_01536_),
    .A(_01535_));
 sg13g2_nor2_1 _08524_ (.A(_01474_),
    .B(_01536_),
    .Y(_01537_));
 sg13g2_nand2_1 _08525_ (.Y(_01538_),
    .A(_01474_),
    .B(_01536_));
 sg13g2_nand2b_1 _08526_ (.Y(_01539_),
    .B(_01538_),
    .A_N(_01537_));
 sg13g2_nand3_1 _08527_ (.B(_01442_),
    .C(_01467_),
    .A(_01439_),
    .Y(_01540_));
 sg13g2_nand2_1 _08528_ (.Y(_01541_),
    .A(_01468_),
    .B(_01540_));
 sg13g2_and2_1 _08529_ (.A(_01390_),
    .B(_01437_),
    .X(_01542_));
 sg13g2_xor2_1 _08530_ (.B(_01542_),
    .A(_01439_),
    .X(_01543_));
 sg13g2_mux2_1 _08531_ (.A0(_01541_),
    .A1(_01543_),
    .S(net1589),
    .X(_01544_));
 sg13g2_xnor2_1 _08532_ (.Y(_01545_),
    .A(net1596),
    .B(_01544_));
 sg13g2_and2_1 _08533_ (.A(net1578),
    .B(_01441_),
    .X(_01546_));
 sg13g2_a21oi_1 _08534_ (.A1(net1589),
    .A2(_01472_),
    .Y(_01547_),
    .B1(_01546_));
 sg13g2_xnor2_1 _08535_ (.Y(_01548_),
    .A(net1550),
    .B(_01547_));
 sg13g2_xnor2_1 _08536_ (.Y(_01549_),
    .A(_01416_),
    .B(_01418_));
 sg13g2_xnor2_1 _08537_ (.Y(_01550_),
    .A(_01416_),
    .B(_01445_));
 sg13g2_mux2_1 _08538_ (.A0(_01549_),
    .A1(_01550_),
    .S(net1577),
    .X(_01551_));
 sg13g2_xnor2_1 _08539_ (.Y(_01552_),
    .A(net1594),
    .B(_01551_));
 sg13g2_inv_1 _08540_ (.Y(_01553_),
    .A(_01552_));
 sg13g2_xnor2_1 _08541_ (.Y(_01554_),
    .A(_01419_),
    .B(_01422_));
 sg13g2_nand2_1 _08542_ (.Y(_01555_),
    .A(net1577),
    .B(_01554_));
 sg13g2_nand4_1 _08543_ (.B(_01447_),
    .C(_01448_),
    .A(_01446_),
    .Y(_01556_),
    .D(_01449_));
 sg13g2_nor2b_1 _08544_ (.A(_01450_),
    .B_N(_01556_),
    .Y(_01557_));
 sg13g2_nand2_1 _08545_ (.Y(_01558_),
    .A(net1588),
    .B(_01557_));
 sg13g2_or2_1 _08546_ (.X(_01559_),
    .B(_01554_),
    .A(net1588));
 sg13g2_nand2b_1 _08547_ (.Y(_01560_),
    .B(net1588),
    .A_N(_01557_));
 sg13g2_a221oi_1 _08548_ (.B2(_01558_),
    .C1(_01528_),
    .B1(_01555_),
    .A1(net1585),
    .Y(_01561_),
    .A2(_01506_));
 sg13g2_a221oi_1 _08549_ (.B2(_01560_),
    .C1(_01527_),
    .B1(_01559_),
    .A1(net1585),
    .Y(_01562_),
    .A2(_01505_));
 sg13g2_nor3_1 _08550_ (.A(_01553_),
    .B(_01561_),
    .C(_01562_),
    .Y(_01563_));
 sg13g2_nand2_1 _08551_ (.Y(_01564_),
    .A(net1588),
    .B(_01550_));
 sg13g2_nand2_1 _08552_ (.Y(_01565_),
    .A(net1577),
    .B(_01549_));
 sg13g2_or2_1 _08553_ (.X(_01566_),
    .B(_01549_),
    .A(net1588));
 sg13g2_nand2b_1 _08554_ (.Y(_01567_),
    .B(net1588),
    .A_N(_01550_));
 sg13g2_a221oi_1 _08555_ (.B2(_01567_),
    .C1(_01527_),
    .B1(_01566_),
    .A1(net1585),
    .Y(_01568_),
    .A2(_01505_));
 sg13g2_xnor2_1 _08556_ (.Y(_01569_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[0] ),
    .B(_01417_));
 sg13g2_xnor2_1 _08557_ (.Y(_01570_),
    .A(net1594),
    .B(_01569_));
 sg13g2_a221oi_1 _08558_ (.B2(_01565_),
    .C1(_01528_),
    .B1(_01564_),
    .A1(net1585),
    .Y(_01571_),
    .A2(_01506_));
 sg13g2_nor3_2 _08559_ (.A(_01568_),
    .B(_01570_),
    .C(_01571_),
    .Y(_01572_));
 sg13g2_o21ai_1 _08560_ (.B1(_01553_),
    .Y(_01573_),
    .A1(_01561_),
    .A2(_01562_));
 sg13g2_nor2b_1 _08561_ (.A(_01563_),
    .B_N(_01573_),
    .Y(_01574_));
 sg13g2_a21oi_2 _08562_ (.B1(_01563_),
    .Y(_01575_),
    .A2(_01573_),
    .A1(_01572_));
 sg13g2_xnor2_1 _08563_ (.Y(_01576_),
    .A(_01409_),
    .B(_01423_));
 sg13g2_xor2_1 _08564_ (.B(_01451_),
    .A(_01409_),
    .X(_01577_));
 sg13g2_mux2_1 _08565_ (.A0(_01576_),
    .A1(_01577_),
    .S(net1577),
    .X(_01578_));
 sg13g2_xnor2_1 _08566_ (.Y(_01579_),
    .A(net1594),
    .B(_01578_));
 sg13g2_xnor2_1 _08567_ (.Y(_01580_),
    .A(_01425_),
    .B(_01427_));
 sg13g2_nand2_1 _08568_ (.Y(_01581_),
    .A(net1576),
    .B(_01580_));
 sg13g2_xnor2_1 _08569_ (.Y(_01582_),
    .A(_01453_),
    .B(_01456_));
 sg13g2_nand2_1 _08570_ (.Y(_01583_),
    .A(net1586),
    .B(_01582_));
 sg13g2_or2_1 _08571_ (.X(_01584_),
    .B(_01580_),
    .A(net1586));
 sg13g2_nand2b_1 _08572_ (.Y(_01585_),
    .B(net1586),
    .A_N(_01582_));
 sg13g2_a221oi_1 _08573_ (.B2(_01585_),
    .C1(_01527_),
    .B1(_01584_),
    .A1(net1586),
    .Y(_01586_),
    .A2(_01505_));
 sg13g2_a221oi_1 _08574_ (.B2(_01583_),
    .C1(_01528_),
    .B1(_01581_),
    .A1(net1585),
    .Y(_01587_),
    .A2(_01506_));
 sg13g2_nor3_1 _08575_ (.A(_01579_),
    .B(_01586_),
    .C(_01587_),
    .Y(_01588_));
 sg13g2_or3_1 _08576_ (.A(_01579_),
    .B(_01586_),
    .C(_01587_),
    .X(_01589_));
 sg13g2_o21ai_1 _08577_ (.B1(_01579_),
    .Y(_01590_),
    .A1(_01586_),
    .A2(_01587_));
 sg13g2_nand2_1 _08578_ (.Y(_01591_),
    .A(_01589_),
    .B(_01590_));
 sg13g2_mux2_1 _08579_ (.A0(_01554_),
    .A1(_01557_),
    .S(net1577),
    .X(_01592_));
 sg13g2_xor2_1 _08580_ (.B(_01592_),
    .A(net1594),
    .X(_01593_));
 sg13g2_or2_1 _08581_ (.X(_01594_),
    .B(_01577_),
    .A(net1577));
 sg13g2_nand2b_1 _08582_ (.Y(_01595_),
    .B(net1576),
    .A_N(_01576_));
 sg13g2_nand2_1 _08583_ (.Y(_01596_),
    .A(net1576),
    .B(_01576_));
 sg13g2_nand2_1 _08584_ (.Y(_01597_),
    .A(net1585),
    .B(_01577_));
 sg13g2_a221oi_1 _08585_ (.B2(_01597_),
    .C1(_01527_),
    .B1(_01596_),
    .A1(net1585),
    .Y(_01598_),
    .A2(_01505_));
 sg13g2_a221oi_1 _08586_ (.B2(_01594_),
    .C1(_01528_),
    .B1(_01595_),
    .A1(net1585),
    .Y(_01599_),
    .A2(_01506_));
 sg13g2_nor3_1 _08587_ (.A(_01593_),
    .B(_01598_),
    .C(_01599_),
    .Y(_01600_));
 sg13g2_or3_1 _08588_ (.A(_01599_),
    .B(_01598_),
    .C(_01593_),
    .X(_01601_));
 sg13g2_o21ai_1 _08589_ (.B1(_01593_),
    .Y(_01602_),
    .A1(_01598_),
    .A2(_01599_));
 sg13g2_nand2_1 _08590_ (.Y(_01603_),
    .A(_01601_),
    .B(_01602_));
 sg13g2_nand4_1 _08591_ (.B(_01590_),
    .C(_01601_),
    .A(_01589_),
    .Y(_01604_),
    .D(_01602_));
 sg13g2_a21oi_1 _08592_ (.A1(_01590_),
    .A2(_01600_),
    .Y(_01605_),
    .B1(_01588_));
 sg13g2_o21ai_1 _08593_ (.B1(_01605_),
    .Y(_01606_),
    .A1(_01604_),
    .A2(_01575_));
 sg13g2_xnor2_1 _08594_ (.Y(_01607_),
    .A(_01404_),
    .B(_01428_));
 sg13g2_xor2_1 _08595_ (.B(_01459_),
    .A(_01404_),
    .X(_01608_));
 sg13g2_mux2_1 _08596_ (.A0(_01607_),
    .A1(_01608_),
    .S(net1576),
    .X(_01609_));
 sg13g2_xor2_1 _08597_ (.B(_01609_),
    .A(net1594),
    .X(_01610_));
 sg13g2_xor2_1 _08598_ (.B(_01432_),
    .A(_01429_),
    .X(_01611_));
 sg13g2_nand3_1 _08599_ (.B(_01460_),
    .C(_01461_),
    .A(_01403_),
    .Y(_01612_));
 sg13g2_and2_1 _08600_ (.A(_01462_),
    .B(_01612_),
    .X(_01613_));
 sg13g2_and2_1 _08601_ (.A(net1588),
    .B(_01613_),
    .X(_01614_));
 sg13g2_a21oi_1 _08602_ (.A1(net1576),
    .A2(_01611_),
    .Y(_01615_),
    .B1(_01614_));
 sg13g2_xnor2_1 _08603_ (.Y(_01616_),
    .A(net1550),
    .B(_01615_));
 sg13g2_nor2_1 _08604_ (.A(_01610_),
    .B(_01616_),
    .Y(_01617_));
 sg13g2_xnor2_1 _08605_ (.Y(_01618_),
    .A(_01616_),
    .B(_01610_));
 sg13g2_xor2_1 _08606_ (.B(_01464_),
    .A(_01463_),
    .X(_01619_));
 sg13g2_xnor2_1 _08607_ (.Y(_01620_),
    .A(_00629_),
    .B(_01396_));
 sg13g2_xnor2_1 _08608_ (.Y(_01621_),
    .A(_01433_),
    .B(_01620_));
 sg13g2_mux2_1 _08609_ (.A0(_01619_),
    .A1(_01621_),
    .S(net1590),
    .X(_01622_));
 sg13g2_xnor2_1 _08610_ (.Y(_01623_),
    .A(net1596),
    .B(_01622_));
 sg13g2_inv_1 _08611_ (.Y(_01624_),
    .A(_01623_));
 sg13g2_xnor2_1 _08612_ (.Y(_01625_),
    .A(_01391_),
    .B(_01466_));
 sg13g2_a21o_1 _08613_ (.A2(_01435_),
    .A1(_01398_),
    .B1(_01392_),
    .X(_01626_));
 sg13g2_nand2_1 _08614_ (.Y(_01627_),
    .A(_01437_),
    .B(_01626_));
 sg13g2_nor2_1 _08615_ (.A(net1590),
    .B(_01627_),
    .Y(_01628_));
 sg13g2_a21oi_1 _08616_ (.A1(net1590),
    .A2(_01625_),
    .Y(_01629_),
    .B1(_01628_));
 sg13g2_xnor2_1 _08617_ (.Y(_01630_),
    .A(_01530_),
    .B(_01629_));
 sg13g2_nor2_1 _08618_ (.A(_01624_),
    .B(_01630_),
    .Y(_01631_));
 sg13g2_and2_1 _08619_ (.A(_01624_),
    .B(_01630_),
    .X(_01632_));
 sg13g2_xnor2_1 _08620_ (.Y(_01633_),
    .A(_01624_),
    .B(_01630_));
 sg13g2_mux2_1 _08621_ (.A0(_01580_),
    .A1(_01582_),
    .S(net1576),
    .X(_01634_));
 sg13g2_xor2_1 _08622_ (.B(_01634_),
    .A(net1594),
    .X(_01635_));
 sg13g2_inv_1 _08623_ (.Y(_01636_),
    .A(_01635_));
 sg13g2_mux2_1 _08624_ (.A0(_01607_),
    .A1(_01608_),
    .S(net1586),
    .X(_01637_));
 sg13g2_xnor2_1 _08625_ (.Y(_01638_),
    .A(_01529_),
    .B(_01637_));
 sg13g2_xnor2_1 _08626_ (.Y(_01639_),
    .A(net1550),
    .B(_01637_));
 sg13g2_nor2_1 _08627_ (.A(_01635_),
    .B(_01638_),
    .Y(_01640_));
 sg13g2_xnor2_1 _08628_ (.Y(_01641_),
    .A(_01635_),
    .B(_01638_));
 sg13g2_inv_1 _08629_ (.Y(_01642_),
    .A(_01641_));
 sg13g2_mux2_1 _08630_ (.A0(_01611_),
    .A1(_01613_),
    .S(net1576),
    .X(_01643_));
 sg13g2_xor2_1 _08631_ (.B(_01643_),
    .A(net1594),
    .X(_01644_));
 sg13g2_inv_1 _08632_ (.Y(_01645_),
    .A(_01644_));
 sg13g2_mux2_1 _08633_ (.A0(_01619_),
    .A1(_01621_),
    .S(net1576),
    .X(_01646_));
 sg13g2_xnor2_1 _08634_ (.Y(_01647_),
    .A(net1550),
    .B(_01646_));
 sg13g2_nor2_1 _08635_ (.A(_01645_),
    .B(_01647_),
    .Y(_01648_));
 sg13g2_nand2_1 _08636_ (.Y(_01649_),
    .A(_01645_),
    .B(_01647_));
 sg13g2_xnor2_1 _08637_ (.Y(_01650_),
    .A(_01645_),
    .B(_01647_));
 sg13g2_nor2_1 _08638_ (.A(_01618_),
    .B(_01641_),
    .Y(_01651_));
 sg13g2_nor4_1 _08639_ (.A(_01618_),
    .B(_01633_),
    .C(_01641_),
    .D(_01650_),
    .Y(_01652_));
 sg13g2_a22oi_1 _08640_ (.Y(_01653_),
    .B1(_01636_),
    .B2(_01639_),
    .A2(_01616_),
    .A1(_01610_));
 sg13g2_nor2_1 _08641_ (.A(_01617_),
    .B(_01653_),
    .Y(_01654_));
 sg13g2_o21ai_1 _08642_ (.B1(_01649_),
    .Y(_01655_),
    .A1(_01617_),
    .A2(_01653_));
 sg13g2_nor2_1 _08643_ (.A(_01631_),
    .B(_01648_),
    .Y(_01656_));
 sg13g2_a221oi_1 _08644_ (.B2(_01656_),
    .C1(_01632_),
    .B1(_01655_),
    .A1(_01652_),
    .Y(_01657_),
    .A2(_01606_));
 sg13g2_nor2_1 _08645_ (.A(net1578),
    .B(_01627_),
    .Y(_01658_));
 sg13g2_a21oi_1 _08646_ (.A1(net1579),
    .A2(_01625_),
    .Y(_01659_),
    .B1(_01658_));
 sg13g2_xnor2_1 _08647_ (.Y(_01660_),
    .A(net1595),
    .B(_01659_));
 sg13g2_mux2_1 _08648_ (.A0(_01541_),
    .A1(_01543_),
    .S(net1578),
    .X(_01661_));
 sg13g2_xnor2_1 _08649_ (.Y(_01662_),
    .A(net1550),
    .B(_01661_));
 sg13g2_nor2b_1 _08650_ (.A(_01660_),
    .B_N(_01662_),
    .Y(_01663_));
 sg13g2_inv_1 _08651_ (.Y(_01664_),
    .A(_01663_));
 sg13g2_xor2_1 _08652_ (.B(_01662_),
    .A(_01660_),
    .X(_01665_));
 sg13g2_nor2b_1 _08653_ (.A(_01545_),
    .B_N(_01548_),
    .Y(_01666_));
 sg13g2_xnor2_1 _08654_ (.Y(_01667_),
    .A(_01545_),
    .B(_01548_));
 sg13g2_nand2b_1 _08655_ (.Y(_01668_),
    .B(_01667_),
    .A_N(_01665_));
 sg13g2_a21oi_1 _08656_ (.A1(_01663_),
    .A2(_01667_),
    .Y(_01669_),
    .B1(_01666_));
 sg13g2_o21ai_1 _08657_ (.B1(_01669_),
    .Y(_01670_),
    .A1(_01668_),
    .A2(_01657_));
 sg13g2_xnor2_1 _08658_ (.Y(_01671_),
    .A(_01539_),
    .B(_01670_));
 sg13g2_o21ai_1 _08659_ (.B1(_01496_),
    .Y(_01672_),
    .A1(_01494_),
    .A2(_01497_));
 sg13g2_xor2_1 _08660_ (.B(_01672_),
    .A(_01480_),
    .X(_01673_));
 sg13g2_o21ai_1 _08661_ (.B1(_01516_),
    .Y(_01674_),
    .A1(_01513_),
    .A2(_01517_));
 sg13g2_xor2_1 _08662_ (.B(_01674_),
    .A(_01515_),
    .X(_01675_));
 sg13g2_mux2_1 _08663_ (.A0(_01673_),
    .A1(_01675_),
    .S(net1579),
    .X(_01676_));
 sg13g2_xnor2_1 _08664_ (.Y(_01677_),
    .A(_01529_),
    .B(_01676_));
 sg13g2_xor2_1 _08665_ (.B(_01497_),
    .A(_01494_),
    .X(_01678_));
 sg13g2_xor2_1 _08666_ (.B(_01517_),
    .A(_01513_),
    .X(_01679_));
 sg13g2_and2_1 _08667_ (.A(net1589),
    .B(_01679_),
    .X(_01680_));
 sg13g2_a21oi_1 _08668_ (.A1(net1578),
    .A2(_01678_),
    .Y(_01681_),
    .B1(_01680_));
 sg13g2_xnor2_1 _08669_ (.Y(_01682_),
    .A(net1596),
    .B(_01681_));
 sg13g2_nor2_1 _08670_ (.A(_01677_),
    .B(_01682_),
    .Y(_01683_));
 sg13g2_xor2_1 _08671_ (.B(_01682_),
    .A(_01677_),
    .X(_01684_));
 sg13g2_mux2_1 _08672_ (.A0(_01531_),
    .A1(_01533_),
    .S(net1580),
    .X(_01685_));
 sg13g2_xnor2_1 _08673_ (.Y(_01686_),
    .A(net1595),
    .B(_01685_));
 sg13g2_and2_1 _08674_ (.A(net1578),
    .B(_01679_),
    .X(_01687_));
 sg13g2_a21oi_1 _08675_ (.A1(net1589),
    .A2(_01678_),
    .Y(_01688_),
    .B1(_01687_));
 sg13g2_xnor2_1 _08676_ (.Y(_01689_),
    .A(net1550),
    .B(_01688_));
 sg13g2_nand2_1 _08677_ (.Y(_01690_),
    .A(_01686_),
    .B(_01689_));
 sg13g2_nor2_1 _08678_ (.A(_01686_),
    .B(_01689_),
    .Y(_01691_));
 sg13g2_a21oi_2 _08679_ (.B1(_01537_),
    .Y(_01692_),
    .A2(_01538_),
    .A1(_01670_));
 sg13g2_o21ai_1 _08680_ (.B1(_01690_),
    .Y(_01693_),
    .A1(_01692_),
    .A2(_01691_));
 sg13g2_xor2_1 _08681_ (.B(_01684_),
    .A(_01693_),
    .X(_01694_));
 sg13g2_nor2_2 _08682_ (.A(_01671_),
    .B(_01694_),
    .Y(_01695_));
 sg13g2_a21oi_1 _08683_ (.A1(_01684_),
    .A2(_01693_),
    .Y(_01696_),
    .B1(_01683_));
 sg13g2_mux2_1 _08684_ (.A0(_01673_),
    .A1(_01675_),
    .S(net1589),
    .X(_01697_));
 sg13g2_xnor2_1 _08685_ (.Y(_01698_),
    .A(net1595),
    .B(_01697_));
 sg13g2_or3_1 _08686_ (.A(_01518_),
    .B(_01519_),
    .C(_01520_),
    .X(_01699_));
 sg13g2_nand2_1 _08687_ (.Y(_01700_),
    .A(_01521_),
    .B(_01699_));
 sg13g2_xnor2_1 _08688_ (.Y(_01701_),
    .A(_01502_),
    .B(_01504_));
 sg13g2_mux2_1 _08689_ (.A0(_01700_),
    .A1(_01701_),
    .S(net1589),
    .X(_01702_));
 sg13g2_xnor2_1 _08690_ (.Y(_01703_),
    .A(net1550),
    .B(_01702_));
 sg13g2_nand2b_1 _08691_ (.Y(_01704_),
    .B(_01703_),
    .A_N(_01698_));
 sg13g2_xnor2_1 _08692_ (.Y(_01705_),
    .A(_01698_),
    .B(_01703_));
 sg13g2_nand2b_1 _08693_ (.Y(_01706_),
    .B(_01705_),
    .A_N(_01696_));
 sg13g2_xnor2_1 _08694_ (.Y(_01707_),
    .A(_01696_),
    .B(_01705_));
 sg13g2_xor2_1 _08695_ (.B(_01689_),
    .A(_01686_),
    .X(_01708_));
 sg13g2_xnor2_1 _08696_ (.Y(_01709_),
    .A(_01692_),
    .B(_01708_));
 sg13g2_nor2_1 _08697_ (.A(_01707_),
    .B(_01709_),
    .Y(_01710_));
 sg13g2_xor2_1 _08698_ (.B(_01709_),
    .A(_01707_),
    .X(_01711_));
 sg13g2_nor2_1 _08699_ (.A(_01695_),
    .B(_01711_),
    .Y(_01712_));
 sg13g2_xor2_1 _08700_ (.B(_01711_),
    .A(_01695_),
    .X(_01713_));
 sg13g2_xnor2_1 _08701_ (.Y(_01714_),
    .A(_01695_),
    .B(_01711_));
 sg13g2_a21oi_1 _08702_ (.A1(_01606_),
    .A2(_01651_),
    .Y(_01715_),
    .B1(_01654_));
 sg13g2_o21ai_1 _08703_ (.B1(_01649_),
    .Y(_01716_),
    .A1(_01650_),
    .A2(_01715_));
 sg13g2_xnor2_1 _08704_ (.Y(_01717_),
    .A(_01633_),
    .B(_01716_));
 sg13g2_a21oi_1 _08705_ (.A1(_01606_),
    .A2(_01642_),
    .Y(_01718_),
    .B1(_01640_));
 sg13g2_xnor2_1 _08706_ (.Y(_01719_),
    .A(_01618_),
    .B(_01718_));
 sg13g2_xor2_1 _08707_ (.B(_01718_),
    .A(_01618_),
    .X(_01720_));
 sg13g2_nand2_1 _08708_ (.Y(_01721_),
    .A(_01717_),
    .B(_01720_));
 sg13g2_xor2_1 _08709_ (.B(_01665_),
    .A(_01657_),
    .X(_01722_));
 sg13g2_xor2_1 _08710_ (.B(_01715_),
    .A(_01650_),
    .X(_01723_));
 sg13g2_inv_1 _08711_ (.Y(_01724_),
    .A(_01723_));
 sg13g2_nand2_1 _08712_ (.Y(_01725_),
    .A(_01722_),
    .B(_01723_));
 sg13g2_xnor2_1 _08713_ (.Y(_01726_),
    .A(_01722_),
    .B(_01723_));
 sg13g2_nor2_1 _08714_ (.A(_01721_),
    .B(_01726_),
    .Y(_01727_));
 sg13g2_nand2_1 _08715_ (.Y(_01728_),
    .A(_01721_),
    .B(_01726_));
 sg13g2_nor2b_1 _08716_ (.A(_01727_),
    .B_N(_01728_),
    .Y(_01729_));
 sg13g2_o21ai_1 _08717_ (.B1(_01601_),
    .Y(_01730_),
    .A1(_01575_),
    .A2(_01603_));
 sg13g2_xor2_1 _08718_ (.B(_01730_),
    .A(_01591_),
    .X(_01731_));
 sg13g2_nor2_1 _08719_ (.A(_01719_),
    .B(_01731_),
    .Y(_01732_));
 sg13g2_xnor2_1 _08720_ (.Y(_01733_),
    .A(_01606_),
    .B(_01642_));
 sg13g2_nor2_2 _08721_ (.A(_01724_),
    .B(_01733_),
    .Y(_01734_));
 sg13g2_xnor2_1 _08722_ (.Y(_01735_),
    .A(_01723_),
    .B(_01733_));
 sg13g2_and2_1 _08723_ (.A(_01732_),
    .B(_01735_),
    .X(_01736_));
 sg13g2_inv_1 _08724_ (.Y(_01737_),
    .A(_01736_));
 sg13g2_xor2_1 _08725_ (.B(_01603_),
    .A(_01575_),
    .X(_01738_));
 sg13g2_inv_1 _08726_ (.Y(_01739_),
    .A(_01738_));
 sg13g2_nor2_1 _08727_ (.A(_01733_),
    .B(_01739_),
    .Y(_01740_));
 sg13g2_xnor2_1 _08728_ (.Y(_01741_),
    .A(_01719_),
    .B(_01731_));
 sg13g2_nor3_1 _08729_ (.A(_01733_),
    .B(_01739_),
    .C(_01741_),
    .Y(_01742_));
 sg13g2_and2_1 _08730_ (.A(_01733_),
    .B(_01739_),
    .X(_01743_));
 sg13g2_nor2_1 _08731_ (.A(_01740_),
    .B(_01743_),
    .Y(_01744_));
 sg13g2_xnor2_1 _08732_ (.Y(_01745_),
    .A(_01572_),
    .B(_01574_));
 sg13g2_nor2_1 _08733_ (.A(_01731_),
    .B(_01745_),
    .Y(_01746_));
 sg13g2_inv_1 _08734_ (.Y(_01747_),
    .A(_01746_));
 sg13g2_nand2_1 _08735_ (.Y(_01748_),
    .A(_01744_),
    .B(_01746_));
 sg13g2_xnor2_1 _08736_ (.Y(_01749_),
    .A(_01740_),
    .B(_01741_));
 sg13g2_nor4_1 _08737_ (.A(_01740_),
    .B(_01741_),
    .C(_01743_),
    .D(_01747_),
    .Y(_01750_));
 sg13g2_or2_1 _08738_ (.X(_01751_),
    .B(_01750_),
    .A(_01742_));
 sg13g2_xor2_1 _08739_ (.B(_01735_),
    .A(_01732_),
    .X(_01752_));
 sg13g2_o21ai_1 _08740_ (.B1(_01752_),
    .Y(_01753_),
    .A1(_01742_),
    .A2(_01750_));
 sg13g2_and2_1 _08741_ (.A(_01737_),
    .B(_01753_),
    .X(_01754_));
 sg13g2_xnor2_1 _08742_ (.Y(_01755_),
    .A(_01717_),
    .B(_01719_));
 sg13g2_and2_1 _08743_ (.A(_01734_),
    .B(_01755_),
    .X(_01756_));
 sg13g2_xor2_1 _08744_ (.B(_01755_),
    .A(_01734_),
    .X(_01757_));
 sg13g2_xnor2_1 _08745_ (.Y(_01758_),
    .A(_01734_),
    .B(_01755_));
 sg13g2_a21oi_1 _08746_ (.A1(_01737_),
    .A2(_01753_),
    .Y(_01759_),
    .B1(_01758_));
 sg13g2_or2_1 _08747_ (.X(_01760_),
    .B(_01756_),
    .A(_01727_));
 sg13g2_a21o_1 _08748_ (.A2(_01756_),
    .A1(_01728_),
    .B1(_01727_),
    .X(_01761_));
 sg13g2_o21ai_1 _08749_ (.B1(_01664_),
    .Y(_01762_),
    .A1(_01657_),
    .A2(_01665_));
 sg13g2_xor2_1 _08750_ (.B(_01762_),
    .A(_01667_),
    .X(_01763_));
 sg13g2_nand2_1 _08751_ (.Y(_01764_),
    .A(_01717_),
    .B(_01763_));
 sg13g2_nand2_1 _08752_ (.Y(_01765_),
    .A(_01671_),
    .B(_01722_));
 sg13g2_xnor2_1 _08753_ (.Y(_01766_),
    .A(_01671_),
    .B(_01722_));
 sg13g2_nand2_1 _08754_ (.Y(_01767_),
    .A(_01764_),
    .B(_01766_));
 sg13g2_xnor2_1 _08755_ (.Y(_01768_),
    .A(_01717_),
    .B(_01763_));
 sg13g2_nor2_1 _08756_ (.A(_01725_),
    .B(_01768_),
    .Y(_01769_));
 sg13g2_nor2_1 _08757_ (.A(_01764_),
    .B(_01766_),
    .Y(_01770_));
 sg13g2_a21o_1 _08758_ (.A2(_01769_),
    .A1(_01767_),
    .B1(_01770_),
    .X(_01771_));
 sg13g2_a221oi_1 _08759_ (.B2(_01728_),
    .C1(_01771_),
    .B1(_01760_),
    .A1(_01729_),
    .Y(_01772_),
    .A2(_01759_));
 sg13g2_xor2_1 _08760_ (.B(_01768_),
    .A(_01725_),
    .X(_01773_));
 sg13g2_xor2_1 _08761_ (.B(_01766_),
    .A(_01764_),
    .X(_01774_));
 sg13g2_a21oi_2 _08762_ (.B1(_01771_),
    .Y(_01775_),
    .A2(_01774_),
    .A1(_01773_));
 sg13g2_or2_2 _08763_ (.X(_01776_),
    .B(_01763_),
    .A(_01709_));
 sg13g2_xnor2_1 _08764_ (.Y(_01777_),
    .A(_01709_),
    .B(_01763_));
 sg13g2_nor2b_2 _08765_ (.A(_01765_),
    .B_N(_01777_),
    .Y(_01778_));
 sg13g2_inv_1 _08766_ (.Y(_01779_),
    .A(_01778_));
 sg13g2_xor2_1 _08767_ (.B(_01777_),
    .A(_01765_),
    .X(_01780_));
 sg13g2_xnor2_1 _08768_ (.Y(_01781_),
    .A(_01694_),
    .B(_01671_));
 sg13g2_nand2_1 _08769_ (.Y(_01782_),
    .A(_01776_),
    .B(_01781_));
 sg13g2_xor2_1 _08770_ (.B(_01781_),
    .A(_01776_),
    .X(_01783_));
 sg13g2_xnor2_1 _08771_ (.Y(_01784_),
    .A(_01781_),
    .B(_01776_));
 sg13g2_nor4_2 _08772_ (.A(_01772_),
    .B(_01775_),
    .C(_01780_),
    .Y(_01785_),
    .D(_01784_));
 sg13g2_or4_1 _08773_ (.A(_01772_),
    .B(_01775_),
    .C(_01780_),
    .D(_01784_),
    .X(_01786_));
 sg13g2_o21ai_1 _08774_ (.B1(_01778_),
    .Y(_01787_),
    .A1(_01776_),
    .A2(_01781_));
 sg13g2_and2_1 _08775_ (.A(_01782_),
    .B(_01787_),
    .X(_01788_));
 sg13g2_nand2_1 _08776_ (.Y(_01789_),
    .A(_01782_),
    .B(_01787_));
 sg13g2_a21oi_2 _08777_ (.B1(_01714_),
    .Y(_01790_),
    .A2(_01788_),
    .A1(_01786_));
 sg13g2_o21ai_1 _08778_ (.B1(_01713_),
    .Y(_01791_),
    .A1(_01785_),
    .A2(_01789_));
 sg13g2_nor3_2 _08779_ (.A(_01713_),
    .B(_01785_),
    .C(_01789_),
    .Y(_01792_));
 sg13g2_nand3_1 _08780_ (.B(_01786_),
    .C(_01788_),
    .A(_01714_),
    .Y(_01793_));
 sg13g2_o21ai_1 _08781_ (.B1(_01714_),
    .Y(_01794_),
    .A1(_01785_),
    .A2(_01789_));
 sg13g2_nand3_1 _08782_ (.B(_01786_),
    .C(_01788_),
    .A(_01713_),
    .Y(_01795_));
 sg13g2_nand2_1 _08783_ (.Y(_01796_),
    .A(net1544),
    .B(net1541));
 sg13g2_xnor2_1 _08784_ (.Y(_01797_),
    .A(\vgadonut.donut.donuthit.rx[14] ),
    .B(net1536));
 sg13g2_xor2_1 _08785_ (.B(net1536),
    .A(\vgadonut.donut.donuthit.rx[14] ),
    .X(_01798_));
 sg13g2_xnor2_1 _08786_ (.Y(_01799_),
    .A(_01748_),
    .B(_01749_));
 sg13g2_o21ai_1 _08787_ (.B1(_01799_),
    .Y(_01800_),
    .A1(net1545),
    .A2(net1542));
 sg13g2_or3_1 _08788_ (.A(net1545),
    .B(net1542),
    .C(_01799_),
    .X(_01801_));
 sg13g2_and2_1 _08789_ (.A(_01800_),
    .B(_01801_),
    .X(_01802_));
 sg13g2_nand2_1 _08790_ (.Y(_01803_),
    .A(_01800_),
    .B(_01801_));
 sg13g2_xnor2_1 _08791_ (.Y(_01804_),
    .A(_01751_),
    .B(_01752_));
 sg13g2_nand3b_1 _08792_ (.B(net1540),
    .C(net1543),
    .Y(_01805_),
    .A_N(_01804_));
 sg13g2_o21ai_1 _08793_ (.B1(_01804_),
    .Y(_01806_),
    .A1(net1545),
    .A2(net1542));
 sg13g2_and2_2 _08794_ (.A(_01805_),
    .B(_01806_),
    .X(_01807_));
 sg13g2_nor3_1 _08795_ (.A(_01772_),
    .B(_01775_),
    .C(_01780_),
    .Y(_01808_));
 sg13g2_or3_1 _08796_ (.A(_01772_),
    .B(_01775_),
    .C(_01780_),
    .X(_01809_));
 sg13g2_nand3_1 _08797_ (.B(_01784_),
    .C(_01809_),
    .A(_01779_),
    .Y(_01810_));
 sg13g2_o21ai_1 _08798_ (.B1(_01783_),
    .Y(_01811_),
    .A1(_01778_),
    .A2(_01808_));
 sg13g2_o21ai_1 _08799_ (.B1(_01784_),
    .Y(_01812_),
    .A1(_01778_),
    .A2(_01808_));
 sg13g2_nand3_1 _08800_ (.B(_01783_),
    .C(_01809_),
    .A(_01779_),
    .Y(_01813_));
 sg13g2_nand2_1 _08801_ (.Y(_01814_),
    .A(_01810_),
    .B(_01811_));
 sg13g2_a22oi_1 _08802_ (.Y(_01815_),
    .B1(_01810_),
    .B2(_01811_),
    .A2(_01795_),
    .A1(_01794_));
 sg13g2_nand4_1 _08803_ (.B(net1544),
    .C(_01812_),
    .A(net1541),
    .Y(_01816_),
    .D(_01813_));
 sg13g2_a22oi_1 _08804_ (.Y(_01817_),
    .B1(_01812_),
    .B2(_01813_),
    .A2(net1541),
    .A1(net1544));
 sg13g2_nand4_1 _08805_ (.B(_01795_),
    .C(_01810_),
    .A(_01794_),
    .Y(_01818_),
    .D(_01811_));
 sg13g2_nor2_1 _08806_ (.A(_01815_),
    .B(_01817_),
    .Y(_01819_));
 sg13g2_nand2_1 _08807_ (.Y(_01820_),
    .A(_01816_),
    .B(_01818_));
 sg13g2_o21ai_1 _08808_ (.B1(_01780_),
    .Y(_01821_),
    .A1(_01772_),
    .A2(_01775_));
 sg13g2_and2_2 _08809_ (.A(_01809_),
    .B(_01821_),
    .X(_01822_));
 sg13g2_o21ai_1 _08810_ (.B1(_01822_),
    .Y(_01823_),
    .A1(net1545),
    .A2(net1542));
 sg13g2_or3_1 _08811_ (.A(net1545),
    .B(net1542),
    .C(_01822_),
    .X(_01824_));
 sg13g2_nand2_1 _08812_ (.Y(_01825_),
    .A(_01823_),
    .B(_01824_));
 sg13g2_and4_1 _08813_ (.A(_01816_),
    .B(_01824_),
    .C(_01823_),
    .D(_01818_),
    .X(_01826_));
 sg13g2_a21o_1 _08814_ (.A2(_01759_),
    .A1(_01729_),
    .B1(_01761_),
    .X(_01827_));
 sg13g2_xor2_1 _08815_ (.B(_01827_),
    .A(_01773_),
    .X(_01828_));
 sg13g2_inv_1 _08816_ (.Y(_01829_),
    .A(_01828_));
 sg13g2_a21oi_1 _08817_ (.A1(net1543),
    .A2(net1540),
    .Y(_01830_),
    .B1(_01828_));
 sg13g2_nor3_1 _08818_ (.A(_01790_),
    .B(_01792_),
    .C(_01829_),
    .Y(_01831_));
 sg13g2_nor3_1 _08819_ (.A(_01790_),
    .B(net1542),
    .C(_01828_),
    .Y(_01832_));
 sg13g2_a21oi_1 _08820_ (.A1(net1543),
    .A2(net1540),
    .Y(_01833_),
    .B1(_01829_));
 sg13g2_a21oi_2 _08821_ (.B1(_01769_),
    .Y(_01834_),
    .A2(_01827_),
    .A1(_01773_));
 sg13g2_xor2_1 _08822_ (.B(_01834_),
    .A(_01774_),
    .X(_01835_));
 sg13g2_xnor2_1 _08823_ (.Y(_01836_),
    .A(_01774_),
    .B(_01834_));
 sg13g2_a21oi_1 _08824_ (.A1(net1543),
    .A2(net1540),
    .Y(_01837_),
    .B1(_01835_));
 sg13g2_nor3_2 _08825_ (.A(_01790_),
    .B(net1542),
    .C(_01836_),
    .Y(_01838_));
 sg13g2_or2_1 _08826_ (.X(_01839_),
    .B(_01838_),
    .A(_01837_));
 sg13g2_nor4_1 _08827_ (.A(_01832_),
    .B(_01833_),
    .C(_01837_),
    .D(_01838_),
    .Y(_01840_));
 sg13g2_nor2_1 _08828_ (.A(_01756_),
    .B(_01759_),
    .Y(_01841_));
 sg13g2_xnor2_1 _08829_ (.Y(_01842_),
    .A(_01729_),
    .B(_01841_));
 sg13g2_nand3_1 _08830_ (.B(net1540),
    .C(_01842_),
    .A(net1543),
    .Y(_01843_));
 sg13g2_a21o_1 _08831_ (.A2(net1540),
    .A1(net1543),
    .B1(_01842_),
    .X(_01844_));
 sg13g2_and2_2 _08832_ (.A(_01843_),
    .B(_01844_),
    .X(_01845_));
 sg13g2_xnor2_1 _08833_ (.Y(_01846_),
    .A(_01754_),
    .B(_01757_));
 sg13g2_or3_1 _08834_ (.A(net1545),
    .B(_01792_),
    .C(_01846_),
    .X(_01847_));
 sg13g2_o21ai_1 _08835_ (.B1(_01846_),
    .Y(_01848_),
    .A1(net1545),
    .A2(net1542));
 sg13g2_nand3_1 _08836_ (.B(net1540),
    .C(_01846_),
    .A(net1543),
    .Y(_01849_));
 sg13g2_a21o_1 _08837_ (.A2(net1540),
    .A1(net1543),
    .B1(_01846_),
    .X(_01850_));
 sg13g2_a22oi_1 _08838_ (.Y(_01851_),
    .B1(_01849_),
    .B2(_01850_),
    .A2(_01844_),
    .A1(_01843_));
 sg13g2_nand3b_1 _08839_ (.B(net1511),
    .C(net1521),
    .Y(_01852_),
    .A_N(_01851_));
 sg13g2_nand3_1 _08840_ (.B(net1512),
    .C(_01851_),
    .A(net1521),
    .Y(_01853_));
 sg13g2_nor3_2 _08841_ (.A(_01802_),
    .B(_01807_),
    .C(net1508),
    .Y(_01854_));
 sg13g2_and4_2 _08842_ (.A(_01807_),
    .B(net1521),
    .C(net1511),
    .D(_01851_),
    .X(_01855_));
 sg13g2_nand4_1 _08843_ (.B(_01807_),
    .C(net1511),
    .A(net1521),
    .Y(_01856_),
    .D(_01851_));
 sg13g2_xnor2_1 _08844_ (.Y(_01857_),
    .A(\vgadonut.donut.donuthit.rx[13] ),
    .B(net1535));
 sg13g2_xor2_1 _08845_ (.B(net1535),
    .A(\vgadonut.donut.donuthit.rx[13] ),
    .X(_01858_));
 sg13g2_and2_1 _08846_ (.A(net1521),
    .B(net1514),
    .X(_01859_));
 sg13g2_xnor2_1 _08847_ (.Y(_01860_),
    .A(\vgadonut.donut.donuthit.rx[9] ),
    .B(net1536));
 sg13g2_nand3_1 _08848_ (.B(net1514),
    .C(_01860_),
    .A(net1520),
    .Y(_01861_));
 sg13g2_and2_1 _08849_ (.A(net1531),
    .B(net1525),
    .X(_01862_));
 sg13g2_nand2_2 _08850_ (.Y(_01863_),
    .A(net1531),
    .B(net1525));
 sg13g2_xnor2_1 _08851_ (.Y(_01864_),
    .A(\vgadonut.donut.donuthit.rx[8] ),
    .B(net1536));
 sg13g2_nand3_1 _08852_ (.B(net1525),
    .C(_01864_),
    .A(net1531),
    .Y(_01865_));
 sg13g2_xnor2_1 _08853_ (.Y(_01866_),
    .A(\vgadonut.donut.donuthit.rx[7] ),
    .B(net1535));
 sg13g2_nand2_1 _08854_ (.Y(_01867_),
    .A(net1529),
    .B(_01866_));
 sg13g2_nor4_2 _08855_ (.A(_01830_),
    .B(_01831_),
    .C(_01837_),
    .Y(_01868_),
    .D(_01838_));
 sg13g2_and2_1 _08856_ (.A(net1521),
    .B(net1509),
    .X(_01869_));
 sg13g2_xnor2_1 _08857_ (.Y(_01870_),
    .A(\vgadonut.donut.donuthit.rx[10] ),
    .B(net1537));
 sg13g2_nand3_1 _08858_ (.B(_01868_),
    .C(_01870_),
    .A(net1520),
    .Y(_01871_));
 sg13g2_nand4_1 _08859_ (.B(_01865_),
    .C(_01867_),
    .A(_01861_),
    .Y(_01872_),
    .D(_01871_));
 sg13g2_and3_1 _08860_ (.X(_01873_),
    .A(net1522),
    .B(net1512),
    .C(_01845_));
 sg13g2_xnor2_1 _08861_ (.Y(_01874_),
    .A(\vgadonut.donut.donuthit.rx[11] ),
    .B(net1537));
 sg13g2_nand4_1 _08862_ (.B(net1512),
    .C(_01845_),
    .A(net1519),
    .Y(_01875_),
    .D(_01874_));
 sg13g2_a22oi_1 _08863_ (.Y(_01876_),
    .B1(_01847_),
    .B2(_01848_),
    .A2(_01844_),
    .A1(_01843_));
 sg13g2_and3_1 _08864_ (.X(_01877_),
    .A(net1521),
    .B(net1512),
    .C(_01876_));
 sg13g2_nand3_1 _08865_ (.B(net1511),
    .C(_01876_),
    .A(net1518),
    .Y(_01878_));
 sg13g2_xnor2_1 _08866_ (.Y(_01879_),
    .A(\vgadonut.donut.donuthit.rx[12] ),
    .B(net1535));
 sg13g2_xor2_1 _08867_ (.B(net1535),
    .A(\vgadonut.donut.donuthit.rx[12] ),
    .X(_01880_));
 sg13g2_nor2_1 _08868_ (.A(_01878_),
    .B(_01880_),
    .Y(_01881_));
 sg13g2_a22oi_1 _08869_ (.Y(_01882_),
    .B1(_01805_),
    .B2(_01806_),
    .A2(_01801_),
    .A1(_01800_));
 sg13g2_and4_1 _08870_ (.A(net1521),
    .B(net1511),
    .C(_01851_),
    .D(_01882_),
    .X(_01883_));
 sg13g2_nand4_1 _08871_ (.B(net1511),
    .C(_01851_),
    .A(net1522),
    .Y(_01884_),
    .D(_01882_));
 sg13g2_nor2_1 _08872_ (.A(_01798_),
    .B(net1496),
    .Y(_01885_));
 sg13g2_o21ai_1 _08873_ (.B1(_01875_),
    .Y(_01886_),
    .A1(_01856_),
    .A2(_01858_));
 sg13g2_nor4_2 _08874_ (.A(_01872_),
    .B(_01881_),
    .C(_01885_),
    .Y(_01887_),
    .D(_01886_));
 sg13g2_nand2_1 _08875_ (.Y(_01888_),
    .A(\vgadonut.donut.donuthit.rx[15] ),
    .B(net1535));
 sg13g2_or2_1 _08876_ (.X(_01889_),
    .B(net1535),
    .A(\vgadonut.donut.donuthit.rx[15] ));
 sg13g2_and2_2 _08877_ (.A(_01888_),
    .B(_01889_),
    .X(_01890_));
 sg13g2_nand2_2 _08878_ (.Y(_01891_),
    .A(_01888_),
    .B(_01889_));
 sg13g2_xor2_1 _08879_ (.B(_01745_),
    .A(_01731_),
    .X(_01892_));
 sg13g2_mux2_1 _08880_ (.A0(_01805_),
    .A1(_01806_),
    .S(_01892_),
    .X(_01893_));
 sg13g2_xnor2_1 _08881_ (.Y(_01894_),
    .A(_01744_),
    .B(_01746_));
 sg13g2_xnor2_1 _08882_ (.Y(_01895_),
    .A(net1539),
    .B(_01894_));
 sg13g2_nand3b_1 _08883_ (.B(_01895_),
    .C(_01802_),
    .Y(_01896_),
    .A_N(_01893_));
 sg13g2_nor2_2 _08884_ (.A(net1508),
    .B(net1495),
    .Y(_01897_));
 sg13g2_or2_2 _08885_ (.X(_01898_),
    .B(_01895_),
    .A(_01803_));
 sg13g2_nor3_2 _08886_ (.A(_01807_),
    .B(net1507),
    .C(_01898_),
    .Y(_01899_));
 sg13g2_or3_2 _08887_ (.A(_01803_),
    .B(_01807_),
    .C(_01895_),
    .X(_01900_));
 sg13g2_a21o_1 _08888_ (.A2(_01900_),
    .A1(net1495),
    .B1(net1507),
    .X(_01901_));
 sg13g2_a21oi_2 _08889_ (.B1(net1507),
    .Y(_01902_),
    .A2(_01900_),
    .A1(net1495));
 sg13g2_a221oi_1 _08890_ (.B2(_01900_),
    .C1(net1507),
    .B1(net1495),
    .A1(_01888_),
    .Y(_01903_),
    .A2(_01889_));
 sg13g2_nand2_2 _08891_ (.Y(_01904_),
    .A(_01891_),
    .B(_01902_));
 sg13g2_nand3_1 _08892_ (.B(net1514),
    .C(_01866_),
    .A(net1520),
    .Y(_01905_));
 sg13g2_nand3_1 _08893_ (.B(_01864_),
    .C(_01868_),
    .A(net1519),
    .Y(_01906_));
 sg13g2_nand2_1 _08894_ (.Y(_01907_),
    .A(\vgadonut.donut.donuthit.rx[5] ),
    .B(_01818_));
 sg13g2_o21ai_1 _08895_ (.B1(_01907_),
    .Y(_01908_),
    .A1(\vgadonut.donut.donuthit.rx[5] ),
    .A2(_01815_));
 sg13g2_xnor2_1 _08896_ (.Y(_01909_),
    .A(\vgadonut.donut.donuthit.rx[6] ),
    .B(net1535));
 sg13g2_nand3_1 _08897_ (.B(net1525),
    .C(_01909_),
    .A(net1531),
    .Y(_01910_));
 sg13g2_nand4_1 _08898_ (.B(_01906_),
    .C(_01908_),
    .A(_01905_),
    .Y(_01911_),
    .D(_01910_));
 sg13g2_nor3_1 _08899_ (.A(_01798_),
    .B(net1507),
    .C(net1495),
    .Y(_01912_));
 sg13g2_and2_1 _08900_ (.A(_01855_),
    .B(_01874_),
    .X(_01913_));
 sg13g2_nor4_1 _08901_ (.A(_01807_),
    .B(net1507),
    .C(_01858_),
    .D(_01898_),
    .Y(_01914_));
 sg13g2_a221oi_1 _08902_ (.B2(_01870_),
    .C1(_01913_),
    .B1(net1497),
    .A1(_01860_),
    .Y(_01915_),
    .A2(net1498));
 sg13g2_nor2_1 _08903_ (.A(_01880_),
    .B(net1496),
    .Y(_01916_));
 sg13g2_nor4_2 _08904_ (.A(_01911_),
    .B(_01912_),
    .C(_01914_),
    .Y(_01917_),
    .D(_01916_));
 sg13g2_a22oi_1 _08905_ (.Y(_01918_),
    .B1(_01915_),
    .B2(_01917_),
    .A2(_01904_),
    .A1(_01887_));
 sg13g2_nand4_1 _08906_ (.B(_01904_),
    .C(_01915_),
    .A(_01887_),
    .Y(_01919_),
    .D(_01917_));
 sg13g2_nor2b_1 _08907_ (.A(_01918_),
    .B_N(_01919_),
    .Y(_01920_));
 sg13g2_and2_1 _08908_ (.A(net2275),
    .B(_01920_),
    .X(_01921_));
 sg13g2_o21ai_1 _08909_ (.B1(net1677),
    .Y(_01922_),
    .A1(net2275),
    .A2(_01920_));
 sg13g2_xor2_1 _08910_ (.B(\vgadonut.donut.donuthit.cordicxy.x2in[4] ),
    .A(net1884),
    .X(_01923_));
 sg13g2_o21ai_1 _08911_ (.B1(\vgadonut.donut.sB[1] ),
    .Y(_01924_),
    .A1(\vgadonut.donut.donuthit.cordicxy.x2in[0] ),
    .A2(\vgadonut.donut.donuthit.cordicxy.x2in[2] ));
 sg13g2_nand2_1 _08912_ (.Y(_01925_),
    .A(_00573_),
    .B(_01924_));
 sg13g2_o21ai_1 _08913_ (.B1(\vgadonut.donut.donuthit.cordicxy.x2in[3] ),
    .Y(_01926_),
    .A1(\vgadonut.donut.sB[1] ),
    .A2(\vgadonut.donut.donuthit.cordicxy.x2in[2] ));
 sg13g2_nor2_1 _08914_ (.A(\vgadonut.donut.sB[0] ),
    .B(net1884),
    .Y(_01927_));
 sg13g2_a21oi_1 _08915_ (.A1(_00569_),
    .A2(_01926_),
    .Y(_01928_),
    .B1(_01927_));
 sg13g2_a22oi_1 _08916_ (.Y(_01929_),
    .B1(_01928_),
    .B2(\vgadonut.donut.donuthit.cordicxy.x2in[0] ),
    .A2(_01925_),
    .A1(\vgadonut.donut.donuthit.cordicxy.x2in[1] ));
 sg13g2_nor2b_1 _08917_ (.A(_01929_),
    .B_N(_01923_),
    .Y(_01930_));
 sg13g2_xnor2_1 _08918_ (.Y(_01931_),
    .A(_01923_),
    .B(_01929_));
 sg13g2_or2_1 _08919_ (.X(_01932_),
    .B(_01931_),
    .A(\vgadonut.donut.donuthit.rxin[5] ));
 sg13g2_nand2_1 _08920_ (.Y(_01933_),
    .A(\vgadonut.donut.donuthit.rxin[5] ),
    .B(_01931_));
 sg13g2_nand3_1 _08921_ (.B(_01932_),
    .C(_01933_),
    .A(net1690),
    .Y(_01934_));
 sg13g2_o21ai_1 _08922_ (.B1(_01934_),
    .Y(_00046_),
    .A1(_01921_),
    .A2(_01922_));
 sg13g2_a21oi_1 _08923_ (.A1(\vgadonut.donut.donuthit.cordicxy.xin[0] ),
    .A2(_01919_),
    .Y(_01935_),
    .B1(_01918_));
 sg13g2_nand3_1 _08924_ (.B(_01868_),
    .C(_01874_),
    .A(net1519),
    .Y(_01936_));
 sg13g2_nand2_1 _08925_ (.Y(_01937_),
    .A(net1526),
    .B(_01864_));
 sg13g2_nand3_1 _08926_ (.B(net1525),
    .C(_01860_),
    .A(net1531),
    .Y(_01938_));
 sg13g2_nand3_1 _08927_ (.B(net1514),
    .C(_01870_),
    .A(net1519),
    .Y(_01939_));
 sg13g2_nand4_1 _08928_ (.B(_01937_),
    .C(_01938_),
    .A(_01936_),
    .Y(_01940_),
    .D(_01939_));
 sg13g2_nand4_1 _08929_ (.B(net1512),
    .C(_01845_),
    .A(net1519),
    .Y(_01941_),
    .D(_01879_));
 sg13g2_nand4_1 _08930_ (.B(net1510),
    .C(_01857_),
    .A(net1519),
    .Y(_01942_),
    .D(_01876_));
 sg13g2_o21ai_1 _08931_ (.B1(_01941_),
    .Y(_01943_),
    .A1(net1496),
    .A2(_01890_));
 sg13g2_o21ai_1 _08932_ (.B1(_01942_),
    .Y(_01944_),
    .A1(_01798_),
    .A2(_01856_));
 sg13g2_nor4_2 _08933_ (.A(_01903_),
    .B(_01940_),
    .C(_01943_),
    .Y(_01945_),
    .D(_01944_));
 sg13g2_nand2_1 _08934_ (.Y(_01946_),
    .A(_01860_),
    .B(net1500));
 sg13g2_nand2_1 _08935_ (.Y(_01947_),
    .A(net1526),
    .B(_01909_));
 sg13g2_a22oi_1 _08936_ (.Y(_01948_),
    .B1(_01866_),
    .B2(net1503),
    .A2(_01864_),
    .A1(net1505));
 sg13g2_nand4_1 _08937_ (.B(net1510),
    .C(_01845_),
    .A(net1519),
    .Y(_01949_),
    .D(_01870_));
 sg13g2_a22oi_1 _08938_ (.Y(_01950_),
    .B1(_01879_),
    .B2(_01855_),
    .A2(net1497),
    .A1(_01874_));
 sg13g2_and4_1 _08939_ (.A(_01946_),
    .B(_01947_),
    .C(_01948_),
    .D(_01950_),
    .X(_01951_));
 sg13g2_o21ai_1 _08940_ (.B1(_01949_),
    .Y(_01952_),
    .A1(_01858_),
    .A2(net1496));
 sg13g2_a221oi_1 _08941_ (.B2(_01797_),
    .C1(_01952_),
    .B1(_01899_),
    .A1(_01891_),
    .Y(_01953_),
    .A2(_01897_));
 sg13g2_a21oi_1 _08942_ (.A1(_01951_),
    .A2(_01953_),
    .Y(_01954_),
    .B1(_01945_));
 sg13g2_a21o_1 _08943_ (.A2(_01953_),
    .A1(_01951_),
    .B1(_01945_),
    .X(_01955_));
 sg13g2_nand3_1 _08944_ (.B(_01951_),
    .C(_01953_),
    .A(_01945_),
    .Y(_01956_));
 sg13g2_and3_1 _08945_ (.X(_01957_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[1] ),
    .B(_01955_),
    .C(_01956_));
 sg13g2_a21oi_1 _08946_ (.A1(_01955_),
    .A2(_01956_),
    .Y(_01958_),
    .B1(\vgadonut.donut.donuthit.cordicxy.xin[1] ));
 sg13g2_nor3_2 _08947_ (.A(_01935_),
    .B(_01957_),
    .C(_01958_),
    .Y(_01959_));
 sg13g2_o21ai_1 _08948_ (.B1(_01935_),
    .Y(_01960_),
    .A1(_01957_),
    .A2(_01958_));
 sg13g2_nand2_1 _08949_ (.Y(_01961_),
    .A(net1676),
    .B(_01960_));
 sg13g2_nor2_1 _08950_ (.A(_01959_),
    .B(_01961_),
    .Y(_01962_));
 sg13g2_a21o_1 _08951_ (.A2(\vgadonut.donut.donuthit.cordicxy.x2in[4] ),
    .A1(net1884),
    .B1(_01930_),
    .X(_01963_));
 sg13g2_nor2_1 _08952_ (.A(_00573_),
    .B(_00577_),
    .Y(_01964_));
 sg13g2_nand2_1 _08953_ (.Y(_01965_),
    .A(_00573_),
    .B(_00577_));
 sg13g2_nor2b_1 _08954_ (.A(_01964_),
    .B_N(_01965_),
    .Y(_01966_));
 sg13g2_xnor2_1 _08955_ (.Y(_01967_),
    .A(_01963_),
    .B(_01966_));
 sg13g2_or2_1 _08956_ (.X(_01968_),
    .B(_01967_),
    .A(_00575_));
 sg13g2_xnor2_1 _08957_ (.Y(_01969_),
    .A(_00575_),
    .B(_01967_));
 sg13g2_or2_1 _08958_ (.X(_01970_),
    .B(_01969_),
    .A(_01933_));
 sg13g2_a21oi_1 _08959_ (.A1(_01933_),
    .A2(_01969_),
    .Y(_01971_),
    .B1(net1676));
 sg13g2_a21o_1 _08960_ (.A2(_01971_),
    .A1(_01970_),
    .B1(_01962_),
    .X(_00053_));
 sg13g2_nor2_1 _08961_ (.A(_01855_),
    .B(_01883_),
    .Y(_01972_));
 sg13g2_nand2_2 _08962_ (.Y(_01973_),
    .A(net1496),
    .B(_01856_));
 sg13g2_a21oi_2 _08963_ (.B1(_01890_),
    .Y(_01974_),
    .A2(_01972_),
    .A1(_01901_));
 sg13g2_o21ai_1 _08964_ (.B1(_01891_),
    .Y(_01975_),
    .A1(_01973_),
    .A2(_01902_));
 sg13g2_nand2_1 _08965_ (.Y(_01976_),
    .A(net1500),
    .B(_01879_));
 sg13g2_nand2_1 _08966_ (.Y(_01977_),
    .A(net1526),
    .B(_01860_));
 sg13g2_a22oi_1 _08967_ (.Y(_01978_),
    .B1(_01874_),
    .B2(net1505),
    .A2(_01870_),
    .A1(net1503));
 sg13g2_a22oi_1 _08968_ (.Y(_01979_),
    .B1(net1497),
    .B2(_01797_),
    .A2(net1498),
    .A1(_01857_));
 sg13g2_and4_2 _08969_ (.A(_01976_),
    .B(_01977_),
    .C(_01978_),
    .D(_01979_),
    .X(_01980_));
 sg13g2_nand2_1 _08970_ (.Y(_01981_),
    .A(_01975_),
    .B(_01980_));
 sg13g2_a22oi_1 _08971_ (.Y(_01982_),
    .B1(_01975_),
    .B2(_01980_),
    .A2(_01904_),
    .A1(_01887_));
 sg13g2_and4_1 _08972_ (.A(_01887_),
    .B(_01904_),
    .C(_01975_),
    .D(_01980_),
    .X(_01983_));
 sg13g2_or3_1 _08973_ (.A(_00624_),
    .B(_01982_),
    .C(_01983_),
    .X(_01984_));
 sg13g2_o21ai_1 _08974_ (.B1(_00624_),
    .Y(_01985_),
    .A1(_01982_),
    .A2(_01983_));
 sg13g2_a21o_1 _08975_ (.A2(_01956_),
    .A1(\vgadonut.donut.donuthit.cordicxy.xin[1] ),
    .B1(_01954_),
    .X(_01986_));
 sg13g2_and3_1 _08976_ (.X(_01987_),
    .A(_01984_),
    .B(_01985_),
    .C(_01986_));
 sg13g2_a21o_1 _08977_ (.A2(_01985_),
    .A1(_01984_),
    .B1(_01986_),
    .X(_01988_));
 sg13g2_nor2b_1 _08978_ (.A(_01987_),
    .B_N(_01988_),
    .Y(_01989_));
 sg13g2_and2_1 _08979_ (.A(_01959_),
    .B(_01989_),
    .X(_01990_));
 sg13g2_o21ai_1 _08980_ (.B1(net1677),
    .Y(_01991_),
    .A1(_01959_),
    .A2(_01989_));
 sg13g2_nand2_1 _08981_ (.Y(_01992_),
    .A(net1883),
    .B(\vgadonut.donut.donuthit.cordicxy.x2in[6] ));
 sg13g2_xor2_1 _08982_ (.B(net1882),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[4] ),
    .X(_01993_));
 sg13g2_and2_1 _08983_ (.A(_01963_),
    .B(_01965_),
    .X(_01994_));
 sg13g2_nor2_1 _08984_ (.A(_01964_),
    .B(_01994_),
    .Y(_01995_));
 sg13g2_o21ai_1 _08985_ (.B1(_01993_),
    .Y(_01996_),
    .A1(_01964_),
    .A2(_01994_));
 sg13g2_xnor2_1 _08986_ (.Y(_01997_),
    .A(_01993_),
    .B(_01995_));
 sg13g2_xnor2_1 _08987_ (.Y(_01998_),
    .A(\vgadonut.donut.donuthit.rxin[7] ),
    .B(_01997_));
 sg13g2_a21oi_1 _08988_ (.A1(_01968_),
    .A2(_01970_),
    .Y(_01999_),
    .B1(_01998_));
 sg13g2_nand3_1 _08989_ (.B(_01970_),
    .C(_01998_),
    .A(_01968_),
    .Y(_02000_));
 sg13g2_nand3b_1 _08990_ (.B(_02000_),
    .C(net1691),
    .Y(_02001_),
    .A_N(_01999_));
 sg13g2_o21ai_1 _08991_ (.B1(_02001_),
    .Y(_00054_),
    .A1(_01990_),
    .A2(_01991_));
 sg13g2_nand2b_1 _08992_ (.Y(_02002_),
    .B(_01984_),
    .A_N(_01982_));
 sg13g2_and2_1 _08993_ (.A(net1526),
    .B(_01870_),
    .X(_02003_));
 sg13g2_nand2_1 _08994_ (.Y(_02004_),
    .A(net1497),
    .B(_01891_));
 sg13g2_a221oi_1 _08995_ (.B2(net1505),
    .C1(_02003_),
    .B1(_01879_),
    .A1(net1503),
    .Y(_02005_),
    .A2(_01874_));
 sg13g2_a22oi_1 _08996_ (.Y(_02006_),
    .B1(net1498),
    .B2(_01797_),
    .A2(net1500),
    .A1(_01857_));
 sg13g2_and4_2 _08997_ (.A(_02004_),
    .B(_01975_),
    .C(_02005_),
    .D(_02006_),
    .X(_02007_));
 sg13g2_nor2_1 _08998_ (.A(_01945_),
    .B(_02007_),
    .Y(_02008_));
 sg13g2_xor2_1 _08999_ (.B(_02007_),
    .A(_01945_),
    .X(_02009_));
 sg13g2_xor2_1 _09000_ (.B(_02009_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[3] ),
    .X(_02010_));
 sg13g2_nor2_1 _09001_ (.A(_02002_),
    .B(_02010_),
    .Y(_02011_));
 sg13g2_xnor2_1 _09002_ (.Y(_02012_),
    .A(_02002_),
    .B(_02010_));
 sg13g2_nor2_1 _09003_ (.A(_01987_),
    .B(_01990_),
    .Y(_02013_));
 sg13g2_xnor2_1 _09004_ (.Y(_02014_),
    .A(_02012_),
    .B(_02013_));
 sg13g2_a21oi_1 _09005_ (.A1(\vgadonut.donut.donuthit.rxin[7] ),
    .A2(_01997_),
    .Y(_02015_),
    .B1(_01999_));
 sg13g2_xnor2_1 _09006_ (.Y(_02016_),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[5] ),
    .B(net1881));
 sg13g2_a21oi_1 _09007_ (.A1(_01992_),
    .A2(_01996_),
    .Y(_02017_),
    .B1(_02016_));
 sg13g2_nand3_1 _09008_ (.B(_01996_),
    .C(_02016_),
    .A(_01992_),
    .Y(_02018_));
 sg13g2_nor2b_1 _09009_ (.A(_02017_),
    .B_N(_02018_),
    .Y(_02019_));
 sg13g2_nand2_1 _09010_ (.Y(_02020_),
    .A(\vgadonut.donut.donuthit.rxin[8] ),
    .B(_02019_));
 sg13g2_xnor2_1 _09011_ (.Y(_02021_),
    .A(\vgadonut.donut.donuthit.rxin[8] ),
    .B(_02019_));
 sg13g2_a21oi_1 _09012_ (.A1(_02015_),
    .A2(_02021_),
    .Y(_02022_),
    .B1(net1676));
 sg13g2_o21ai_1 _09013_ (.B1(_02022_),
    .Y(_02023_),
    .A1(_02015_),
    .A2(_02021_));
 sg13g2_o21ai_1 _09014_ (.B1(_02023_),
    .Y(_00055_),
    .A1(net1692),
    .A2(_02014_));
 sg13g2_nand2b_1 _09015_ (.Y(_02024_),
    .B(_01891_),
    .A_N(_01852_));
 sg13g2_nand2_1 _09016_ (.Y(_02025_),
    .A(_01797_),
    .B(net1500));
 sg13g2_nand2_1 _09017_ (.Y(_02026_),
    .A(_01857_),
    .B(net1505));
 sg13g2_a22oi_1 _09018_ (.Y(_02027_),
    .B1(_01879_),
    .B2(net1502),
    .A2(_01874_),
    .A1(net1526));
 sg13g2_nand4_1 _09019_ (.B(_02025_),
    .C(_02026_),
    .A(_02024_),
    .Y(_02028_),
    .D(_02027_));
 sg13g2_nor2_2 _09020_ (.A(_01974_),
    .B(_02028_),
    .Y(_02029_));
 sg13g2_a21oi_1 _09021_ (.A1(_01975_),
    .A2(_01980_),
    .Y(_02030_),
    .B1(_02029_));
 sg13g2_xnor2_1 _09022_ (.Y(_02031_),
    .A(_01981_),
    .B(_02029_));
 sg13g2_xnor2_1 _09023_ (.Y(_02032_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[4] ),
    .B(_02031_));
 sg13g2_a21oi_1 _09024_ (.A1(\vgadonut.donut.donuthit.cordicxy.xin[3] ),
    .A2(_02009_),
    .Y(_02033_),
    .B1(_02008_));
 sg13g2_nor2_1 _09025_ (.A(_02032_),
    .B(_02033_),
    .Y(_02034_));
 sg13g2_xnor2_1 _09026_ (.Y(_02035_),
    .A(_02032_),
    .B(_02033_));
 sg13g2_a221oi_1 _09027_ (.B2(_02002_),
    .C1(_01987_),
    .B1(_02010_),
    .A1(_01959_),
    .Y(_02036_),
    .A2(_01988_));
 sg13g2_o21ai_1 _09028_ (.B1(_02035_),
    .Y(_02037_),
    .A1(_02011_),
    .A2(_02036_));
 sg13g2_nor3_2 _09029_ (.A(_02011_),
    .B(_02036_),
    .C(_02035_),
    .Y(_02038_));
 sg13g2_nor2_1 _09030_ (.A(net1692),
    .B(_02038_),
    .Y(_02039_));
 sg13g2_o21ai_1 _09031_ (.B1(_02020_),
    .Y(_02040_),
    .A1(_02015_),
    .A2(_02021_));
 sg13g2_xor2_1 _09032_ (.B(net1879),
    .A(net1882),
    .X(_02041_));
 sg13g2_a21oi_1 _09033_ (.A1(\vgadonut.donut.donuthit.cordicxy.x2in[5] ),
    .A2(net1881),
    .Y(_02042_),
    .B1(_02017_));
 sg13g2_nand2b_1 _09034_ (.Y(_02043_),
    .B(_02041_),
    .A_N(_02042_));
 sg13g2_xnor2_1 _09035_ (.Y(_02044_),
    .A(_02041_),
    .B(_02042_));
 sg13g2_nand2_1 _09036_ (.Y(_02045_),
    .A(\vgadonut.donut.donuthit.rxin[9] ),
    .B(_02044_));
 sg13g2_xnor2_1 _09037_ (.Y(_02046_),
    .A(\vgadonut.donut.donuthit.rxin[9] ),
    .B(_02044_));
 sg13g2_nand2b_1 _09038_ (.Y(_02047_),
    .B(_02040_),
    .A_N(_02046_));
 sg13g2_nand2b_1 _09039_ (.Y(_02048_),
    .B(_02046_),
    .A_N(_02040_));
 sg13g2_and3_1 _09040_ (.X(_02049_),
    .A(net1690),
    .B(_02047_),
    .C(_02048_));
 sg13g2_a21o_1 _09041_ (.A2(_02039_),
    .A1(_02037_),
    .B1(_02049_),
    .X(_00056_));
 sg13g2_nand2_1 _09042_ (.Y(_02050_),
    .A(_02045_),
    .B(_02047_));
 sg13g2_o21ai_1 _09043_ (.B1(_02043_),
    .Y(_02051_),
    .A1(_00579_),
    .A2(_00583_));
 sg13g2_xnor2_1 _09044_ (.Y(_02052_),
    .A(net1881),
    .B(net1878));
 sg13g2_xnor2_1 _09045_ (.Y(_02053_),
    .A(_02051_),
    .B(_02052_));
 sg13g2_nand2_1 _09046_ (.Y(_02054_),
    .A(\vgadonut.donut.donuthit.rxin[10] ),
    .B(_02053_));
 sg13g2_xnor2_1 _09047_ (.Y(_02055_),
    .A(_00584_),
    .B(_02053_));
 sg13g2_nor2_1 _09048_ (.A(_02050_),
    .B(_02055_),
    .Y(_02056_));
 sg13g2_nand2_1 _09049_ (.Y(_02057_),
    .A(_02050_),
    .B(_02055_));
 sg13g2_nand2_1 _09050_ (.Y(_02058_),
    .A(net1694),
    .B(_02057_));
 sg13g2_a21oi_2 _09051_ (.B1(_02030_),
    .Y(_02059_),
    .A2(_02031_),
    .A1(\vgadonut.donut.donuthit.cordicxy.xin[4] ));
 sg13g2_a22oi_1 _09052_ (.Y(_02060_),
    .B1(net1499),
    .B2(_01891_),
    .A2(net1502),
    .A1(_01857_));
 sg13g2_a22oi_1 _09053_ (.Y(_02061_),
    .B1(_01879_),
    .B2(net1526),
    .A2(net1504),
    .A1(_01797_));
 sg13g2_and4_2 _09054_ (.A(_01975_),
    .B(_02024_),
    .C(_02060_),
    .D(_02061_),
    .X(_02062_));
 sg13g2_nor2_1 _09055_ (.A(_02007_),
    .B(_02062_),
    .Y(_02063_));
 sg13g2_xor2_1 _09056_ (.B(_02062_),
    .A(_02007_),
    .X(_02064_));
 sg13g2_xnor2_1 _09057_ (.Y(_02065_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[5] ),
    .B(_02064_));
 sg13g2_nand2_1 _09058_ (.Y(_02066_),
    .A(_02059_),
    .B(_02065_));
 sg13g2_nor2_1 _09059_ (.A(_02059_),
    .B(_02065_),
    .Y(_02067_));
 sg13g2_xnor2_1 _09060_ (.Y(_02068_),
    .A(_02059_),
    .B(_02065_));
 sg13g2_nor2_1 _09061_ (.A(_02034_),
    .B(_02038_),
    .Y(_02069_));
 sg13g2_a21oi_1 _09062_ (.A1(_02068_),
    .A2(_02069_),
    .Y(_02070_),
    .B1(net1695));
 sg13g2_o21ai_1 _09063_ (.B1(_02070_),
    .Y(_02071_),
    .A1(_02068_),
    .A2(_02069_));
 sg13g2_o21ai_1 _09064_ (.B1(_02071_),
    .Y(_00057_),
    .A1(_02056_),
    .A2(_02058_));
 sg13g2_nand2_1 _09065_ (.Y(_02072_),
    .A(net1879),
    .B(net1876));
 sg13g2_nor2_1 _09066_ (.A(net1879),
    .B(net1875),
    .Y(_02073_));
 sg13g2_xor2_1 _09067_ (.B(net1875),
    .A(net1879),
    .X(_02074_));
 sg13g2_a21o_1 _09068_ (.A2(net1878),
    .A1(net1881),
    .B1(_02051_),
    .X(_02075_));
 sg13g2_o21ai_1 _09069_ (.B1(_02075_),
    .Y(_02076_),
    .A1(net1880),
    .A2(net1878));
 sg13g2_xnor2_1 _09070_ (.Y(_02077_),
    .A(_02074_),
    .B(_02076_));
 sg13g2_nand2_1 _09071_ (.Y(_02078_),
    .A(\vgadonut.donut.donuthit.rxin[11] ),
    .B(_02077_));
 sg13g2_xnor2_1 _09072_ (.Y(_02079_),
    .A(\vgadonut.donut.donuthit.rxin[11] ),
    .B(_02077_));
 sg13g2_nand3_1 _09073_ (.B(_02057_),
    .C(_02079_),
    .A(_02054_),
    .Y(_02080_));
 sg13g2_a21o_1 _09074_ (.A2(_02057_),
    .A1(_02054_),
    .B1(_02079_),
    .X(_02081_));
 sg13g2_and2_1 _09075_ (.A(_02080_),
    .B(_02081_),
    .X(_02082_));
 sg13g2_o21ai_1 _09076_ (.B1(_01891_),
    .Y(_02083_),
    .A1(net1504),
    .A2(net1499));
 sg13g2_nand2_2 _09077_ (.Y(_02084_),
    .A(_02024_),
    .B(_02083_));
 sg13g2_nand2b_2 _09078_ (.Y(_02085_),
    .B(_01975_),
    .A_N(_02084_));
 sg13g2_nand2_1 _09079_ (.Y(_02086_),
    .A(net1526),
    .B(_01857_));
 sg13g2_o21ai_1 _09080_ (.B1(_02086_),
    .Y(_02087_),
    .A1(_01798_),
    .A2(_01863_));
 sg13g2_nor3_2 _09081_ (.A(_01974_),
    .B(_02084_),
    .C(_02087_),
    .Y(_02088_));
 sg13g2_or2_1 _09082_ (.X(_02089_),
    .B(_02088_),
    .A(_02029_));
 sg13g2_xnor2_1 _09083_ (.Y(_02090_),
    .A(_02029_),
    .B(_02088_));
 sg13g2_xnor2_1 _09084_ (.Y(_02091_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[6] ),
    .B(_02090_));
 sg13g2_xnor2_1 _09085_ (.Y(_02092_),
    .A(_00623_),
    .B(_02090_));
 sg13g2_a21oi_2 _09086_ (.B1(_02063_),
    .Y(_02093_),
    .A2(_02064_),
    .A1(\vgadonut.donut.donuthit.cordicxy.xin[5] ));
 sg13g2_nor2_1 _09087_ (.A(_02092_),
    .B(_02093_),
    .Y(_02094_));
 sg13g2_nand2b_1 _09088_ (.Y(_02095_),
    .B(_02091_),
    .A_N(_02093_));
 sg13g2_xnor2_1 _09089_ (.Y(_02096_),
    .A(_02091_),
    .B(_02093_));
 sg13g2_xnor2_1 _09090_ (.Y(_02097_),
    .A(_02092_),
    .B(_02093_));
 sg13g2_or3_1 _09091_ (.A(_02034_),
    .B(_02038_),
    .C(_02067_),
    .X(_02098_));
 sg13g2_a21o_1 _09092_ (.A2(_02066_),
    .A1(_02034_),
    .B1(_02067_),
    .X(_02099_));
 sg13g2_a21o_1 _09093_ (.A2(_02098_),
    .A1(_02066_),
    .B1(_02096_),
    .X(_02100_));
 sg13g2_and3_1 _09094_ (.X(_02101_),
    .A(_02066_),
    .B(_02096_),
    .C(_02098_));
 sg13g2_nor2_1 _09095_ (.A(net1695),
    .B(_02101_),
    .Y(_02102_));
 sg13g2_a22oi_1 _09096_ (.Y(_02103_),
    .B1(_02100_),
    .B2(_02102_),
    .A2(_02082_),
    .A1(net1695));
 sg13g2_inv_1 _09097_ (.Y(_00058_),
    .A(_02103_));
 sg13g2_o21ai_1 _09098_ (.B1(_02072_),
    .Y(_02104_),
    .A1(_02073_),
    .A2(_02076_));
 sg13g2_xnor2_1 _09099_ (.Y(_02105_),
    .A(net1878),
    .B(net1874));
 sg13g2_xnor2_1 _09100_ (.Y(_02106_),
    .A(_02104_),
    .B(_02105_));
 sg13g2_nand2_1 _09101_ (.Y(_02107_),
    .A(\vgadonut.donut.donuthit.rxin[12] ),
    .B(_02106_));
 sg13g2_xnor2_1 _09102_ (.Y(_02108_),
    .A(\vgadonut.donut.donuthit.rxin[12] ),
    .B(_02106_));
 sg13g2_nand3_1 _09103_ (.B(_02081_),
    .C(_02108_),
    .A(_02078_),
    .Y(_02109_));
 sg13g2_a21o_1 _09104_ (.A2(_02081_),
    .A1(_02078_),
    .B1(_02108_),
    .X(_02110_));
 sg13g2_nand3_1 _09105_ (.B(_02109_),
    .C(_02110_),
    .A(net1694),
    .Y(_02111_));
 sg13g2_nor2_1 _09106_ (.A(_02094_),
    .B(_02101_),
    .Y(_02112_));
 sg13g2_o21ai_1 _09107_ (.B1(_02089_),
    .Y(_02113_),
    .A1(_00623_),
    .A2(_02090_));
 sg13g2_nand2_1 _09108_ (.Y(_02114_),
    .A(_01797_),
    .B(net1526));
 sg13g2_o21ai_1 _09109_ (.B1(_02114_),
    .Y(_02115_),
    .A1(_01863_),
    .A2(_01890_));
 sg13g2_nor3_2 _09110_ (.A(_01974_),
    .B(_02084_),
    .C(_02115_),
    .Y(_02116_));
 sg13g2_or2_1 _09111_ (.X(_02117_),
    .B(_02116_),
    .A(_02062_));
 sg13g2_xnor2_1 _09112_ (.Y(_02118_),
    .A(_02062_),
    .B(_02116_));
 sg13g2_xnor2_1 _09113_ (.Y(_02119_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[7] ),
    .B(_02118_));
 sg13g2_nor2_1 _09114_ (.A(_02113_),
    .B(_02119_),
    .Y(_02120_));
 sg13g2_nand2_1 _09115_ (.Y(_02121_),
    .A(_02113_),
    .B(_02119_));
 sg13g2_xnor2_1 _09116_ (.Y(_02122_),
    .A(_02113_),
    .B(_02119_));
 sg13g2_xnor2_1 _09117_ (.Y(_02123_),
    .A(_02112_),
    .B(_02122_));
 sg13g2_o21ai_1 _09118_ (.B1(_02111_),
    .Y(_00059_),
    .A1(net1695),
    .A2(_02123_));
 sg13g2_nand2_1 _09119_ (.Y(_02124_),
    .A(net1875),
    .B(net1872));
 sg13g2_nor2_1 _09120_ (.A(net1875),
    .B(net1872),
    .Y(_02125_));
 sg13g2_xor2_1 _09121_ (.B(net1872),
    .A(net1875),
    .X(_02126_));
 sg13g2_a21o_1 _09122_ (.A2(net1874),
    .A1(net1877),
    .B1(_02104_),
    .X(_02127_));
 sg13g2_o21ai_1 _09123_ (.B1(_02127_),
    .Y(_02128_),
    .A1(net1877),
    .A2(net1874));
 sg13g2_xnor2_1 _09124_ (.Y(_02129_),
    .A(_02126_),
    .B(_02128_));
 sg13g2_xnor2_1 _09125_ (.Y(_02130_),
    .A(\vgadonut.donut.donuthit.rxin[13] ),
    .B(_02129_));
 sg13g2_nand3_1 _09126_ (.B(_02110_),
    .C(_02130_),
    .A(_02107_),
    .Y(_02131_));
 sg13g2_a21o_1 _09127_ (.A2(_02110_),
    .A1(_02107_),
    .B1(_02130_),
    .X(_02132_));
 sg13g2_inv_1 _09128_ (.Y(_02133_),
    .A(_02132_));
 sg13g2_nand3_1 _09129_ (.B(_02131_),
    .C(_02132_),
    .A(net1694),
    .Y(_02134_));
 sg13g2_nor2_1 _09130_ (.A(_02097_),
    .B(_02122_),
    .Y(_02135_));
 sg13g2_nor3_1 _09131_ (.A(_02068_),
    .B(_02097_),
    .C(_02122_),
    .Y(_02136_));
 sg13g2_a21oi_1 _09132_ (.A1(_02095_),
    .A2(_02121_),
    .Y(_02137_),
    .B1(_02120_));
 sg13g2_a221oi_1 _09133_ (.B2(_02136_),
    .C1(_02137_),
    .B1(_02038_),
    .A1(_02099_),
    .Y(_02138_),
    .A2(_02135_));
 sg13g2_nor2_2 _09134_ (.A(net1519),
    .B(_01890_),
    .Y(_02139_));
 sg13g2_nor2_2 _09135_ (.A(_02085_),
    .B(_02139_),
    .Y(_02140_));
 sg13g2_nor2_1 _09136_ (.A(_02088_),
    .B(_02140_),
    .Y(_02141_));
 sg13g2_xnor2_1 _09137_ (.Y(_02142_),
    .A(_02088_),
    .B(_02140_));
 sg13g2_inv_1 _09138_ (.Y(_02143_),
    .A(_02142_));
 sg13g2_xnor2_1 _09139_ (.Y(_02144_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[8] ),
    .B(_02142_));
 sg13g2_o21ai_1 _09140_ (.B1(_02117_),
    .Y(_02145_),
    .A1(_00622_),
    .A2(_02118_));
 sg13g2_nand2_1 _09141_ (.Y(_02146_),
    .A(_02144_),
    .B(_02145_));
 sg13g2_xor2_1 _09142_ (.B(_02145_),
    .A(_02144_),
    .X(_02147_));
 sg13g2_nand2b_1 _09143_ (.Y(_02148_),
    .B(_02147_),
    .A_N(_02138_));
 sg13g2_xnor2_1 _09144_ (.Y(_02149_),
    .A(_02138_),
    .B(_02147_));
 sg13g2_nand2_1 _09145_ (.Y(_02150_),
    .A(net1677),
    .B(_02149_));
 sg13g2_nand2_1 _09146_ (.Y(_00060_),
    .A(_02134_),
    .B(_02150_));
 sg13g2_a21oi_1 _09147_ (.A1(\vgadonut.donut.donuthit.cordicxy.xin[8] ),
    .A2(_02143_),
    .Y(_02151_),
    .B1(_02141_));
 sg13g2_a21oi_1 _09148_ (.A1(_02115_),
    .A2(_02139_),
    .Y(_02152_),
    .B1(_02085_));
 sg13g2_xnor2_1 _09149_ (.Y(_02153_),
    .A(_02116_),
    .B(_02140_));
 sg13g2_xnor2_1 _09150_ (.Y(_02154_),
    .A(_00621_),
    .B(_02153_));
 sg13g2_nor2_1 _09151_ (.A(_02151_),
    .B(_02154_),
    .Y(_02155_));
 sg13g2_inv_1 _09152_ (.Y(_02156_),
    .A(_02155_));
 sg13g2_xnor2_1 _09153_ (.Y(_02157_),
    .A(_02151_),
    .B(_02154_));
 sg13g2_nand3_1 _09154_ (.B(_02148_),
    .C(_02157_),
    .A(_02146_),
    .Y(_02158_));
 sg13g2_a21o_1 _09155_ (.A2(_02148_),
    .A1(_02146_),
    .B1(_02157_),
    .X(_02159_));
 sg13g2_nand2_1 _09156_ (.Y(_02160_),
    .A(_02158_),
    .B(_02159_));
 sg13g2_a21oi_1 _09157_ (.A1(\vgadonut.donut.donuthit.rxin[13] ),
    .A2(_02129_),
    .Y(_02161_),
    .B1(_02133_));
 sg13g2_xnor2_1 _09158_ (.Y(_02162_),
    .A(net1874),
    .B(net1870));
 sg13g2_o21ai_1 _09159_ (.B1(_02124_),
    .Y(_02163_),
    .A1(_02125_),
    .A2(_02128_));
 sg13g2_xnor2_1 _09160_ (.Y(_02164_),
    .A(_02162_),
    .B(_02163_));
 sg13g2_xnor2_1 _09161_ (.Y(_02165_),
    .A(\vgadonut.donut.donuthit.rxin[14] ),
    .B(_02164_));
 sg13g2_nor2_1 _09162_ (.A(_02161_),
    .B(_02165_),
    .Y(_02166_));
 sg13g2_a21oi_1 _09163_ (.A1(_02161_),
    .A2(_02165_),
    .Y(_02167_),
    .B1(net1677));
 sg13g2_nand2b_1 _09164_ (.Y(_02168_),
    .B(_02167_),
    .A_N(_02166_));
 sg13g2_o21ai_1 _09165_ (.B1(_02168_),
    .Y(_00061_),
    .A1(net1697),
    .A2(_02160_));
 sg13g2_o21ai_1 _09166_ (.B1(_02152_),
    .Y(_02169_),
    .A1(_00621_),
    .A2(_02153_));
 sg13g2_nand2_1 _09167_ (.Y(_02170_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[10] ),
    .B(_02169_));
 sg13g2_xnor2_1 _09168_ (.Y(_02171_),
    .A(\vgadonut.donut.donuthit.cordicxy.xin[10] ),
    .B(_02169_));
 sg13g2_nand3_1 _09169_ (.B(_02159_),
    .C(_02171_),
    .A(_02156_),
    .Y(_02172_));
 sg13g2_a21o_1 _09170_ (.A2(_02159_),
    .A1(_02156_),
    .B1(_02171_),
    .X(_02173_));
 sg13g2_nand3_1 _09171_ (.B(_02172_),
    .C(_02173_),
    .A(net1677),
    .Y(_02174_));
 sg13g2_a21o_1 _09172_ (.A2(_02164_),
    .A1(\vgadonut.donut.donuthit.rxin[14] ),
    .B1(_02166_),
    .X(_02175_));
 sg13g2_nand2_1 _09173_ (.Y(_02176_),
    .A(net1872),
    .B(net1869));
 sg13g2_nor2_1 _09174_ (.A(net1871),
    .B(net1869),
    .Y(_02177_));
 sg13g2_xor2_1 _09175_ (.B(net1869),
    .A(net1871),
    .X(_02178_));
 sg13g2_a21o_1 _09176_ (.A2(net1869),
    .A1(net1873),
    .B1(_02163_),
    .X(_02179_));
 sg13g2_o21ai_1 _09177_ (.B1(_02179_),
    .Y(_02180_),
    .A1(net1873),
    .A2(net1869));
 sg13g2_xnor2_1 _09178_ (.Y(_02181_),
    .A(_02178_),
    .B(_02180_));
 sg13g2_inv_1 _09179_ (.Y(_02182_),
    .A(_02181_));
 sg13g2_xnor2_1 _09180_ (.Y(_02183_),
    .A(\vgadonut.donut.donuthit.rxin[15] ),
    .B(_02181_));
 sg13g2_nand2b_1 _09181_ (.Y(_02184_),
    .B(_02175_),
    .A_N(_02183_));
 sg13g2_nand2b_1 _09182_ (.Y(_02185_),
    .B(_02183_),
    .A_N(_02175_));
 sg13g2_nand3_1 _09183_ (.B(_02184_),
    .C(_02185_),
    .A(net1696),
    .Y(_02186_));
 sg13g2_nand2_1 _09184_ (.Y(_00047_),
    .A(_02174_),
    .B(_02186_));
 sg13g2_o21ai_1 _09185_ (.B1(_02184_),
    .Y(_02187_),
    .A1(net2182),
    .A2(_02182_));
 sg13g2_o21ai_1 _09186_ (.B1(_02176_),
    .Y(_02188_),
    .A1(_02177_),
    .A2(_02180_));
 sg13g2_nand2_1 _09187_ (.Y(_02189_),
    .A(\vgadonut.donut.donuthit.rxin[15] ),
    .B(_02188_));
 sg13g2_xnor2_1 _09188_ (.Y(_02190_),
    .A(_00593_),
    .B(_02188_));
 sg13g2_xnor2_1 _09189_ (.Y(_02191_),
    .A(_02187_),
    .B(_02190_));
 sg13g2_o21ai_1 _09190_ (.B1(_00159_),
    .Y(_02192_),
    .A1(_02085_),
    .A2(_02139_));
 sg13g2_xnor2_1 _09191_ (.Y(_02193_),
    .A(_00159_),
    .B(_02140_));
 sg13g2_a21oi_2 _09192_ (.B1(_02193_),
    .Y(_02194_),
    .A2(_02173_),
    .A1(_02170_));
 sg13g2_a21o_1 _09193_ (.A2(_02173_),
    .A1(_02170_),
    .B1(_02193_),
    .X(_02195_));
 sg13g2_nand3_1 _09194_ (.B(_02173_),
    .C(_02193_),
    .A(_02170_),
    .Y(_02196_));
 sg13g2_nand3_1 _09195_ (.B(_02195_),
    .C(_02196_),
    .A(net1677),
    .Y(_02197_));
 sg13g2_o21ai_1 _09196_ (.B1(_02197_),
    .Y(_00048_),
    .A1(net1677),
    .A2(_02191_));
 sg13g2_nand2b_1 _09197_ (.Y(_02198_),
    .B(_02188_),
    .A_N(_00160_));
 sg13g2_nand3b_1 _09198_ (.B(_02190_),
    .C(_02198_),
    .Y(_02199_),
    .A_N(_02187_));
 sg13g2_o21ai_1 _09199_ (.B1(_02199_),
    .Y(_02200_),
    .A1(net2182),
    .A2(_02189_));
 sg13g2_nand2_2 _09200_ (.Y(_02201_),
    .A(net1697),
    .B(net2183));
 sg13g2_xnor2_1 _09201_ (.Y(_02202_),
    .A(net2202),
    .B(_02192_));
 sg13g2_nand2b_1 _09202_ (.Y(_02203_),
    .B(_02194_),
    .A_N(_02202_));
 sg13g2_xnor2_1 _09203_ (.Y(_02204_),
    .A(_02195_),
    .B(_02202_));
 sg13g2_o21ai_1 _09204_ (.B1(_02201_),
    .Y(_00049_),
    .A1(net1697),
    .A2(_02204_));
 sg13g2_o21ai_1 _09205_ (.B1(net2361),
    .Y(_02205_),
    .A1(_02085_),
    .A2(_02139_));
 sg13g2_o21ai_1 _09206_ (.B1(_02203_),
    .Y(_02206_),
    .A1(net2353),
    .A2(_02205_));
 sg13g2_nor2b_1 _09207_ (.A(_02140_),
    .B_N(_00162_),
    .Y(_02207_));
 sg13g2_xnor2_1 _09208_ (.Y(_02208_),
    .A(net2197),
    .B(_02205_));
 sg13g2_xor2_1 _09209_ (.B(_02208_),
    .A(_02206_),
    .X(_02209_));
 sg13g2_o21ai_1 _09210_ (.B1(_02201_),
    .Y(_00050_),
    .A1(net1697),
    .A2(_02209_));
 sg13g2_nor2_1 _09211_ (.A(_02202_),
    .B(_02208_),
    .Y(_02210_));
 sg13g2_nand2_1 _09212_ (.Y(_02211_),
    .A(_00159_),
    .B(net2361));
 sg13g2_a22oi_1 _09213_ (.Y(_02212_),
    .B1(_02211_),
    .B2(_02207_),
    .A2(_02194_),
    .A1(_02210_));
 sg13g2_nor2b_1 _09214_ (.A(_02140_),
    .B_N(net2362),
    .Y(_02213_));
 sg13g2_nand2b_1 _09215_ (.Y(_02214_),
    .B(_02213_),
    .A_N(net2197));
 sg13g2_xor2_1 _09216_ (.B(_02207_),
    .A(net2352),
    .X(_02215_));
 sg13g2_xnor2_1 _09217_ (.Y(_02216_),
    .A(_02212_),
    .B(_02215_));
 sg13g2_o21ai_1 _09218_ (.B1(_02201_),
    .Y(_00051_),
    .A1(net1697),
    .A2(_02216_));
 sg13g2_o21ai_1 _09219_ (.B1(_02214_),
    .Y(_02217_),
    .A1(_02212_),
    .A2(_02215_));
 sg13g2_xor2_1 _09220_ (.B(_02213_),
    .A(net2186),
    .X(_02218_));
 sg13g2_xnor2_1 _09221_ (.Y(_02219_),
    .A(_02217_),
    .B(_02218_));
 sg13g2_o21ai_1 _09222_ (.B1(_02201_),
    .Y(_00052_),
    .A1(net1697),
    .A2(_02219_));
 sg13g2_xnor2_1 _09223_ (.Y(_02220_),
    .A(\vgadonut.donut.donuthit.ry[14] ),
    .B(net1532));
 sg13g2_xor2_1 _09224_ (.B(net1532),
    .A(\vgadonut.donut.donuthit.ry[14] ),
    .X(_02221_));
 sg13g2_xnor2_1 _09225_ (.Y(_02222_),
    .A(\vgadonut.donut.donuthit.ry[13] ),
    .B(net1532));
 sg13g2_inv_1 _09226_ (.Y(_02223_),
    .A(_02222_));
 sg13g2_xnor2_1 _09227_ (.Y(_02224_),
    .A(\vgadonut.donut.donuthit.ry[9] ),
    .B(net1532));
 sg13g2_nand3_1 _09228_ (.B(net1513),
    .C(_02224_),
    .A(net1515),
    .Y(_02225_));
 sg13g2_xnor2_1 _09229_ (.Y(_02226_),
    .A(\vgadonut.donut.donuthit.ry[7] ),
    .B(net1534));
 sg13g2_nand2_1 _09230_ (.Y(_02227_),
    .A(net1527),
    .B(_02226_));
 sg13g2_xnor2_1 _09231_ (.Y(_02228_),
    .A(\vgadonut.donut.donuthit.ry[8] ),
    .B(net1532));
 sg13g2_nand3_1 _09232_ (.B(net1524),
    .C(_02228_),
    .A(net1530),
    .Y(_02229_));
 sg13g2_xnor2_1 _09233_ (.Y(_02230_),
    .A(\vgadonut.donut.donuthit.ry[10] ),
    .B(net1532));
 sg13g2_inv_1 _09234_ (.Y(_02231_),
    .A(_02230_));
 sg13g2_nand3_1 _09235_ (.B(net1509),
    .C(_02230_),
    .A(net1515),
    .Y(_02232_));
 sg13g2_nand4_1 _09236_ (.B(_02227_),
    .C(_02229_),
    .A(_02225_),
    .Y(_02233_),
    .D(_02232_));
 sg13g2_xnor2_1 _09237_ (.Y(_02234_),
    .A(\vgadonut.donut.donuthit.ry[11] ),
    .B(net1532));
 sg13g2_nand4_1 _09238_ (.B(net1510),
    .C(_01845_),
    .A(net1516),
    .Y(_02235_),
    .D(_02234_));
 sg13g2_xnor2_1 _09239_ (.Y(_02236_),
    .A(\vgadonut.donut.donuthit.ry[12] ),
    .B(net1532));
 sg13g2_inv_1 _09240_ (.Y(_02237_),
    .A(_02236_));
 sg13g2_nand4_1 _09241_ (.B(net1510),
    .C(_01876_),
    .A(net1516),
    .Y(_02238_),
    .D(_02236_));
 sg13g2_o21ai_1 _09242_ (.B1(_02235_),
    .Y(_02239_),
    .A1(net1496),
    .A2(_02221_));
 sg13g2_o21ai_1 _09243_ (.B1(_02238_),
    .Y(_02240_),
    .A1(_01856_),
    .A2(_02223_));
 sg13g2_nand2_1 _09244_ (.Y(_02241_),
    .A(\vgadonut.donut.donuthit.ry[15] ),
    .B(net1533));
 sg13g2_or2_1 _09245_ (.X(_02242_),
    .B(net1533),
    .A(\vgadonut.donut.donuthit.ry[15] ));
 sg13g2_and2_1 _09246_ (.A(_02241_),
    .B(_02242_),
    .X(_02243_));
 sg13g2_nand2_2 _09247_ (.Y(_02244_),
    .A(_02241_),
    .B(_02242_));
 sg13g2_a221oi_1 _09248_ (.B2(_02242_),
    .C1(net1507),
    .B1(_02241_),
    .A1(net1495),
    .Y(_02245_),
    .A2(_01900_));
 sg13g2_nor4_2 _09249_ (.A(_02233_),
    .B(_02239_),
    .C(_02240_),
    .Y(_02246_),
    .D(_02245_));
 sg13g2_nand4_1 _09250_ (.B(net1510),
    .C(_01845_),
    .A(net1515),
    .Y(_02247_),
    .D(_02224_));
 sg13g2_o21ai_1 _09251_ (.B1(_02247_),
    .Y(_02248_),
    .A1(_01878_),
    .A2(_02231_));
 sg13g2_nand3_1 _09252_ (.B(net1513),
    .C(_02226_),
    .A(net1515),
    .Y(_02249_));
 sg13g2_nand3_1 _09253_ (.B(net1509),
    .C(_02228_),
    .A(net1515),
    .Y(_02250_));
 sg13g2_nand2_1 _09254_ (.Y(_02251_),
    .A(\vgadonut.donut.donuthit.ry[5] ),
    .B(_01818_));
 sg13g2_o21ai_1 _09255_ (.B1(_02251_),
    .Y(_02252_),
    .A1(\vgadonut.donut.donuthit.ry[5] ),
    .A2(_01815_));
 sg13g2_xnor2_1 _09256_ (.Y(_02253_),
    .A(\vgadonut.donut.donuthit.ry[6] ),
    .B(net1533));
 sg13g2_nand3_1 _09257_ (.B(net1524),
    .C(_02253_),
    .A(net1530),
    .Y(_02254_));
 sg13g2_nand4_1 _09258_ (.B(_02250_),
    .C(_02252_),
    .A(_02249_),
    .Y(_02255_),
    .D(_02254_));
 sg13g2_nor3_1 _09259_ (.A(net1507),
    .B(net1495),
    .C(_02221_),
    .Y(_02256_));
 sg13g2_and2_1 _09260_ (.A(_01855_),
    .B(_02234_),
    .X(_02257_));
 sg13g2_nor4_2 _09261_ (.A(_02248_),
    .B(_02255_),
    .C(_02256_),
    .Y(_02258_),
    .D(_02257_));
 sg13g2_a22oi_1 _09262_ (.Y(_02259_),
    .B1(_02236_),
    .B2(_01854_),
    .A2(_02222_),
    .A1(_01899_));
 sg13g2_a21oi_1 _09263_ (.A1(_02258_),
    .A2(_02259_),
    .Y(_02260_),
    .B1(_02246_));
 sg13g2_nand3_1 _09264_ (.B(_02258_),
    .C(_02259_),
    .A(_02246_),
    .Y(_02261_));
 sg13g2_nand2b_1 _09265_ (.Y(_02262_),
    .B(_02261_),
    .A_N(_02260_));
 sg13g2_a21oi_1 _09266_ (.A1(_00625_),
    .A2(_02262_),
    .Y(_02263_),
    .B1(net1684));
 sg13g2_o21ai_1 _09267_ (.B1(_02263_),
    .Y(_02264_),
    .A1(_00625_),
    .A2(_02262_));
 sg13g2_xor2_1 _09268_ (.B(net1931),
    .A(net1934),
    .X(_02265_));
 sg13g2_o21ai_1 _09269_ (.B1(\vgadonut.donut.sAcB[1] ),
    .Y(_02266_),
    .A1(\vgadonut.donut.sAcB[2] ),
    .A2(net1934));
 sg13g2_nand2b_1 _09270_ (.Y(_02267_),
    .B(_02266_),
    .A_N(net1932));
 sg13g2_o21ai_1 _09271_ (.B1(net1932),
    .Y(_02268_),
    .A1(\vgadonut.donut.sAcB[1] ),
    .A2(net1934));
 sg13g2_nor2_1 _09272_ (.A(\vgadonut.donut.sAcB[0] ),
    .B(net1934),
    .Y(_02269_));
 sg13g2_a21oi_1 _09273_ (.A1(_06898_),
    .A2(_02268_),
    .Y(_02270_),
    .B1(_02269_));
 sg13g2_a22oi_1 _09274_ (.Y(_02271_),
    .B1(_02270_),
    .B2(\vgadonut.donut.sAcB[2] ),
    .A2(_02267_),
    .A1(\vgadonut.donut.sAcB[3] ));
 sg13g2_nor2b_1 _09275_ (.A(_02271_),
    .B_N(_02265_),
    .Y(_02272_));
 sg13g2_xnor2_1 _09276_ (.Y(_02273_),
    .A(_02265_),
    .B(_02271_));
 sg13g2_and2_2 _09277_ (.A(\vgadonut.donut.donuthit.ryin[5] ),
    .B(_02273_),
    .X(_02274_));
 sg13g2_o21ai_1 _09278_ (.B1(net1682),
    .Y(_02275_),
    .A1(net2338),
    .A2(_02273_));
 sg13g2_o21ai_1 _09279_ (.B1(_02264_),
    .Y(_00062_),
    .A1(_02274_),
    .A2(_02275_));
 sg13g2_a21oi_1 _09280_ (.A1(\vgadonut.donut.donuthit.cordicxy.yin[0] ),
    .A2(_02261_),
    .Y(_02276_),
    .B1(_02260_));
 sg13g2_nand3_1 _09281_ (.B(net1513),
    .C(_02230_),
    .A(net1515),
    .Y(_02277_));
 sg13g2_nand3_1 _09282_ (.B(net1524),
    .C(_02224_),
    .A(net1530),
    .Y(_02278_));
 sg13g2_nand2_1 _09283_ (.Y(_02279_),
    .A(net1527),
    .B(_02228_));
 sg13g2_nand3_1 _09284_ (.B(net1509),
    .C(_02234_),
    .A(net1515),
    .Y(_02280_));
 sg13g2_nand4_1 _09285_ (.B(_02278_),
    .C(_02279_),
    .A(_02277_),
    .Y(_02281_),
    .D(_02280_));
 sg13g2_nand4_1 _09286_ (.B(net1510),
    .C(_01845_),
    .A(net1516),
    .Y(_02282_),
    .D(_02236_));
 sg13g2_nand4_1 _09287_ (.B(net1510),
    .C(_01876_),
    .A(net1515),
    .Y(_02283_),
    .D(_02222_));
 sg13g2_o21ai_1 _09288_ (.B1(_02282_),
    .Y(_02284_),
    .A1(net1496),
    .A2(_02243_));
 sg13g2_o21ai_1 _09289_ (.B1(_02283_),
    .Y(_02285_),
    .A1(_01856_),
    .A2(_02221_));
 sg13g2_nor4_2 _09290_ (.A(_02245_),
    .B(_02281_),
    .C(_02284_),
    .Y(_02286_),
    .D(_02285_));
 sg13g2_nand2_1 _09291_ (.Y(_02287_),
    .A(net1527),
    .B(_02253_));
 sg13g2_nand2_1 _09292_ (.Y(_02288_),
    .A(net1499),
    .B(_02224_));
 sg13g2_a22oi_1 _09293_ (.Y(_02289_),
    .B1(_02228_),
    .B2(net1504),
    .A2(_02226_),
    .A1(net1502));
 sg13g2_nand4_1 _09294_ (.B(net1510),
    .C(_01876_),
    .A(net1516),
    .Y(_02290_),
    .D(_02234_));
 sg13g2_a22oi_1 _09295_ (.Y(_02291_),
    .B1(_02230_),
    .B2(net1498),
    .A2(_02222_),
    .A1(_01883_));
 sg13g2_and4_1 _09296_ (.A(_02287_),
    .B(_02288_),
    .C(_02289_),
    .D(_02291_),
    .X(_02292_));
 sg13g2_o21ai_1 _09297_ (.B1(_02290_),
    .Y(_02293_),
    .A1(_01856_),
    .A2(_02237_));
 sg13g2_a221oi_1 _09298_ (.B2(_01897_),
    .C1(_02293_),
    .B1(_02244_),
    .A1(_01899_),
    .Y(_02294_),
    .A2(_02220_));
 sg13g2_a21oi_1 _09299_ (.A1(_02292_),
    .A2(_02294_),
    .Y(_02295_),
    .B1(_02286_));
 sg13g2_a21o_1 _09300_ (.A2(_02294_),
    .A1(_02292_),
    .B1(_02286_),
    .X(_02296_));
 sg13g2_nand3_1 _09301_ (.B(_02292_),
    .C(_02294_),
    .A(_02286_),
    .Y(_02297_));
 sg13g2_and3_1 _09302_ (.X(_02298_),
    .A(net291),
    .B(_02296_),
    .C(_02297_));
 sg13g2_a21oi_2 _09303_ (.B1(net300),
    .Y(_02299_),
    .A2(_02297_),
    .A1(_02296_));
 sg13g2_or2_1 _09304_ (.X(_02300_),
    .B(_02299_),
    .A(_02298_));
 sg13g2_nor3_2 _09305_ (.A(_02276_),
    .B(_02299_),
    .C(_02298_),
    .Y(_02301_));
 sg13g2_a21o_1 _09306_ (.A2(_02300_),
    .A1(_02276_),
    .B1(net1684),
    .X(_02302_));
 sg13g2_a21o_1 _09307_ (.A2(\vgadonut.donut.sAcB[6] ),
    .A1(\vgadonut.donut.sAcB[4] ),
    .B1(_02272_),
    .X(_02303_));
 sg13g2_xnor2_1 _09308_ (.Y(_02304_),
    .A(net1933),
    .B(\vgadonut.donut.sAcB[7] ));
 sg13g2_xnor2_1 _09309_ (.Y(_02305_),
    .A(_02303_),
    .B(_02304_));
 sg13g2_xnor2_1 _09310_ (.Y(_02306_),
    .A(net2326),
    .B(_02305_));
 sg13g2_a21oi_1 _09311_ (.A1(_02274_),
    .A2(_02306_),
    .Y(_02307_),
    .B1(net1675));
 sg13g2_o21ai_1 _09312_ (.B1(_02307_),
    .Y(_02308_),
    .A1(_02274_),
    .A2(_02306_));
 sg13g2_o21ai_1 _09313_ (.B1(_02308_),
    .Y(_00069_),
    .A1(_02301_),
    .A2(_02302_));
 sg13g2_a22oi_1 _09314_ (.Y(_02309_),
    .B1(_02306_),
    .B2(_02274_),
    .A2(_02305_),
    .A1(net2041));
 sg13g2_nand2_1 _09315_ (.Y(_02310_),
    .A(net1931),
    .B(net1929));
 sg13g2_xor2_1 _09316_ (.B(net1929),
    .A(net1931),
    .X(_02311_));
 sg13g2_a21o_1 _09317_ (.A2(\vgadonut.donut.sAcB[7] ),
    .A1(net1933),
    .B1(_02303_),
    .X(_02312_));
 sg13g2_o21ai_1 _09318_ (.B1(_02312_),
    .Y(_02313_),
    .A1(net1933),
    .A2(\vgadonut.donut.sAcB[7] ));
 sg13g2_inv_1 _09319_ (.Y(_02314_),
    .A(_02313_));
 sg13g2_nand2_1 _09320_ (.Y(_02315_),
    .A(_02311_),
    .B(_02314_));
 sg13g2_xnor2_1 _09321_ (.Y(_02316_),
    .A(_02311_),
    .B(_02313_));
 sg13g2_xnor2_1 _09322_ (.Y(_02317_),
    .A(\vgadonut.donut.donuthit.ryin[7] ),
    .B(_02316_));
 sg13g2_nor2_1 _09323_ (.A(_02309_),
    .B(_02317_),
    .Y(_02318_));
 sg13g2_xnor2_1 _09324_ (.Y(_02319_),
    .A(_02309_),
    .B(_02317_));
 sg13g2_o21ai_1 _09325_ (.B1(_02244_),
    .Y(_02320_),
    .A1(_01902_),
    .A2(_01973_));
 sg13g2_a22oi_1 _09326_ (.Y(_02321_),
    .B1(_02234_),
    .B2(net1504),
    .A2(_02224_),
    .A1(net1527));
 sg13g2_a22oi_1 _09327_ (.Y(_02322_),
    .B1(_02236_),
    .B2(net1499),
    .A2(_02230_),
    .A1(net1502));
 sg13g2_a22oi_1 _09328_ (.Y(_02323_),
    .B1(_02222_),
    .B2(net1498),
    .A2(_02220_),
    .A1(net1497));
 sg13g2_and3_1 _09329_ (.X(_02324_),
    .A(_02321_),
    .B(_02322_),
    .C(_02323_));
 sg13g2_and2_1 _09330_ (.A(net1494),
    .B(_02324_),
    .X(_02325_));
 sg13g2_nor2_1 _09331_ (.A(_02246_),
    .B(_02325_),
    .Y(_02326_));
 sg13g2_a21o_1 _09332_ (.A2(_02324_),
    .A1(net1494),
    .B1(_02246_),
    .X(_02327_));
 sg13g2_nand3_1 _09333_ (.B(net1494),
    .C(_02324_),
    .A(_02246_),
    .Y(_02328_));
 sg13g2_and3_1 _09334_ (.X(_02329_),
    .A(net296),
    .B(_02327_),
    .C(_02328_));
 sg13g2_a21oi_1 _09335_ (.A1(_02327_),
    .A2(_02328_),
    .Y(_02330_),
    .B1(\vgadonut.donut.donuthit.cordicxy.yin[2] ));
 sg13g2_a21oi_1 _09336_ (.A1(net292),
    .A2(_02297_),
    .Y(_02331_),
    .B1(_02295_));
 sg13g2_nor3_1 _09337_ (.A(_02329_),
    .B(_02330_),
    .C(_02331_),
    .Y(_02332_));
 sg13g2_o21ai_1 _09338_ (.B1(_02331_),
    .Y(_02333_),
    .A1(_02329_),
    .A2(_02330_));
 sg13g2_nor2b_1 _09339_ (.A(_02332_),
    .B_N(_02333_),
    .Y(_02334_));
 sg13g2_a21oi_1 _09340_ (.A1(_02301_),
    .A2(_02334_),
    .Y(_02335_),
    .B1(net1683));
 sg13g2_o21ai_1 _09341_ (.B1(_02335_),
    .Y(_02336_),
    .A1(_02301_),
    .A2(_02334_));
 sg13g2_o21ai_1 _09342_ (.B1(_02336_),
    .Y(_00070_),
    .A1(net1675),
    .A2(_02319_));
 sg13g2_a21oi_1 _09343_ (.A1(\vgadonut.donut.donuthit.ryin[7] ),
    .A2(_02316_),
    .Y(_02337_),
    .B1(_02318_));
 sg13g2_xnor2_1 _09344_ (.Y(_02338_),
    .A(net1930),
    .B(\vgadonut.donut.sAcB[9] ));
 sg13g2_a21oi_1 _09345_ (.A1(_02310_),
    .A2(_02315_),
    .Y(_02339_),
    .B1(_02338_));
 sg13g2_nand3_1 _09346_ (.B(_02315_),
    .C(_02338_),
    .A(_02310_),
    .Y(_02340_));
 sg13g2_nor2b_2 _09347_ (.A(_02339_),
    .B_N(_02340_),
    .Y(_02341_));
 sg13g2_nand2_1 _09348_ (.Y(_02342_),
    .A(\vgadonut.donut.donuthit.ryin[8] ),
    .B(_02341_));
 sg13g2_xnor2_1 _09349_ (.Y(_02343_),
    .A(net2327),
    .B(_02341_));
 sg13g2_or2_1 _09350_ (.X(_02344_),
    .B(_02343_),
    .A(_02337_));
 sg13g2_a21oi_1 _09351_ (.A1(_02337_),
    .A2(_02343_),
    .Y(_02345_),
    .B1(net1675));
 sg13g2_nand2_1 _09352_ (.Y(_02346_),
    .A(_02344_),
    .B(_02345_));
 sg13g2_or2_1 _09353_ (.X(_02347_),
    .B(_02329_),
    .A(_02326_));
 sg13g2_nand2_1 _09354_ (.Y(_02348_),
    .A(net1504),
    .B(_02236_));
 sg13g2_nor2_1 _09355_ (.A(net1530),
    .B(_02231_),
    .Y(_02349_));
 sg13g2_a221oi_1 _09356_ (.B2(net1502),
    .C1(_02349_),
    .B1(_02234_),
    .A1(net1499),
    .Y(_02350_),
    .A2(_02222_));
 sg13g2_a22oi_1 _09357_ (.Y(_02351_),
    .B1(_02244_),
    .B2(net1497),
    .A2(_02220_),
    .A1(net1498));
 sg13g2_and4_2 _09358_ (.A(net1494),
    .B(_02348_),
    .C(_02350_),
    .D(_02351_),
    .X(_02352_));
 sg13g2_nor2_1 _09359_ (.A(_02286_),
    .B(_02352_),
    .Y(_02353_));
 sg13g2_xor2_1 _09360_ (.B(_02352_),
    .A(_02286_),
    .X(_02354_));
 sg13g2_xor2_1 _09361_ (.B(_02354_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[3] ),
    .X(_02355_));
 sg13g2_nor2_1 _09362_ (.A(_02347_),
    .B(_02355_),
    .Y(_02356_));
 sg13g2_xnor2_1 _09363_ (.Y(_02357_),
    .A(_02347_),
    .B(_02355_));
 sg13g2_a21oi_1 _09364_ (.A1(_02301_),
    .A2(_02333_),
    .Y(_02358_),
    .B1(_02332_));
 sg13g2_xnor2_1 _09365_ (.Y(_02359_),
    .A(_02357_),
    .B(_02358_));
 sg13g2_o21ai_1 _09366_ (.B1(_02346_),
    .Y(_00071_),
    .A1(net1683),
    .A2(_02359_));
 sg13g2_nand2b_2 _09367_ (.Y(_02360_),
    .B(_02244_),
    .A_N(_01852_));
 sg13g2_nand2_1 _09368_ (.Y(_02361_),
    .A(net1499),
    .B(_02220_));
 sg13g2_nand2_1 _09369_ (.Y(_02362_),
    .A(net1504),
    .B(_02222_));
 sg13g2_a22oi_1 _09370_ (.Y(_02363_),
    .B1(_02236_),
    .B2(net1502),
    .A2(_02234_),
    .A1(net1527));
 sg13g2_nand4_1 _09371_ (.B(_02361_),
    .C(_02362_),
    .A(_02360_),
    .Y(_02364_),
    .D(_02363_));
 sg13g2_nor2b_2 _09372_ (.A(_02364_),
    .B_N(net1494),
    .Y(_02365_));
 sg13g2_nor2_1 _09373_ (.A(_02325_),
    .B(_02365_),
    .Y(_02366_));
 sg13g2_xor2_1 _09374_ (.B(_02365_),
    .A(_02325_),
    .X(_02367_));
 sg13g2_xnor2_1 _09375_ (.Y(_02368_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[4] ),
    .B(_02367_));
 sg13g2_a21oi_1 _09376_ (.A1(\vgadonut.donut.donuthit.cordicxy.yin[3] ),
    .A2(_02354_),
    .Y(_02369_),
    .B1(_02353_));
 sg13g2_nor2_1 _09377_ (.A(_02368_),
    .B(_02369_),
    .Y(_02370_));
 sg13g2_xnor2_1 _09378_ (.Y(_02371_),
    .A(_02368_),
    .B(_02369_));
 sg13g2_a221oi_1 _09379_ (.B2(_02355_),
    .C1(_02332_),
    .B1(_02347_),
    .A1(_02333_),
    .Y(_02372_),
    .A2(_02301_));
 sg13g2_or2_1 _09380_ (.X(_02373_),
    .B(_02372_),
    .A(_02356_));
 sg13g2_nor2_2 _09381_ (.A(_02372_),
    .B(_02356_),
    .Y(_02374_));
 sg13g2_nand2b_1 _09382_ (.Y(_02375_),
    .B(_02374_),
    .A_N(_02371_));
 sg13g2_a21oi_1 _09383_ (.A1(_02371_),
    .A2(_02373_),
    .Y(_02376_),
    .B1(net1684));
 sg13g2_xor2_1 _09384_ (.B(net1926),
    .A(net1929),
    .X(_02377_));
 sg13g2_a21oi_1 _09385_ (.A1(net1930),
    .A2(\vgadonut.donut.sAcB[9] ),
    .Y(_02378_),
    .B1(_02339_));
 sg13g2_nand2b_1 _09386_ (.Y(_02379_),
    .B(_02377_),
    .A_N(_02378_));
 sg13g2_xnor2_1 _09387_ (.Y(_02380_),
    .A(_02377_),
    .B(_02378_));
 sg13g2_xnor2_1 _09388_ (.Y(_02381_),
    .A(\vgadonut.donut.donuthit.ryin[9] ),
    .B(_02380_));
 sg13g2_a21oi_1 _09389_ (.A1(_02342_),
    .A2(_02344_),
    .Y(_02382_),
    .B1(_02381_));
 sg13g2_and3_1 _09390_ (.X(_02383_),
    .A(_02342_),
    .B(_02344_),
    .C(_02381_));
 sg13g2_nor3_1 _09391_ (.A(net1675),
    .B(_02382_),
    .C(_02383_),
    .Y(_02384_));
 sg13g2_a21o_1 _09392_ (.A2(_02376_),
    .A1(_02375_),
    .B1(_02384_),
    .X(_00072_));
 sg13g2_a21oi_1 _09393_ (.A1(net2187),
    .A2(_02380_),
    .Y(_02385_),
    .B1(_02382_));
 sg13g2_o21ai_1 _09394_ (.B1(_02379_),
    .Y(_02386_),
    .A1(_06910_),
    .A2(_00548_));
 sg13g2_xnor2_1 _09395_ (.Y(_02387_),
    .A(\vgadonut.donut.sAcB[9] ),
    .B(net1925));
 sg13g2_xnor2_1 _09396_ (.Y(_02388_),
    .A(_02386_),
    .B(_02387_));
 sg13g2_nand2_1 _09397_ (.Y(_02389_),
    .A(net2274),
    .B(_02388_));
 sg13g2_xnor2_1 _09398_ (.Y(_02390_),
    .A(net2274),
    .B(_02388_));
 sg13g2_or2_1 _09399_ (.X(_02391_),
    .B(_02390_),
    .A(_02385_));
 sg13g2_a21oi_1 _09400_ (.A1(_02385_),
    .A2(_02390_),
    .Y(_02392_),
    .B1(net1675));
 sg13g2_nand2_1 _09401_ (.Y(_02393_),
    .A(_02391_),
    .B(_02392_));
 sg13g2_a21oi_2 _09402_ (.B1(_02366_),
    .Y(_02394_),
    .A2(_02367_),
    .A1(\vgadonut.donut.donuthit.cordicxy.yin[4] ));
 sg13g2_nand2_1 _09403_ (.Y(_02395_),
    .A(net1527),
    .B(_02236_));
 sg13g2_o21ai_1 _09404_ (.B1(_02395_),
    .Y(_02396_),
    .A1(_01863_),
    .A2(_02223_));
 sg13g2_a221oi_1 _09405_ (.B2(net1499),
    .C1(_02396_),
    .B1(_02244_),
    .A1(net1504),
    .Y(_02397_),
    .A2(_02220_));
 sg13g2_and3_2 _09406_ (.X(_02398_),
    .A(_02320_),
    .B(_02360_),
    .C(_02397_));
 sg13g2_nor2_1 _09407_ (.A(_02352_),
    .B(_02398_),
    .Y(_02399_));
 sg13g2_xor2_1 _09408_ (.B(_02352_),
    .A(_02398_),
    .X(_02400_));
 sg13g2_xnor2_1 _09409_ (.Y(_02401_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[5] ),
    .B(_02400_));
 sg13g2_nand2_1 _09410_ (.Y(_02402_),
    .A(_02394_),
    .B(_02401_));
 sg13g2_nor2_1 _09411_ (.A(_02394_),
    .B(_02401_),
    .Y(_02403_));
 sg13g2_xnor2_1 _09412_ (.Y(_02404_),
    .A(_02394_),
    .B(_02401_));
 sg13g2_nor2b_1 _09413_ (.A(_02370_),
    .B_N(_02375_),
    .Y(_02405_));
 sg13g2_a21oi_1 _09414_ (.A1(_02404_),
    .A2(_02405_),
    .Y(_02406_),
    .B1(net1681));
 sg13g2_o21ai_1 _09415_ (.B1(_02406_),
    .Y(_02407_),
    .A1(_02404_),
    .A2(_02405_));
 sg13g2_nand2_1 _09416_ (.Y(_00073_),
    .A(_02393_),
    .B(_02407_));
 sg13g2_nand2_1 _09417_ (.Y(_02408_),
    .A(net1926),
    .B(net1923));
 sg13g2_nor2_1 _09418_ (.A(net1926),
    .B(net1923),
    .Y(_02409_));
 sg13g2_xor2_1 _09419_ (.B(net1923),
    .A(net1926),
    .X(_02410_));
 sg13g2_a21o_1 _09420_ (.A2(net1924),
    .A1(net1928),
    .B1(_02386_),
    .X(_02411_));
 sg13g2_o21ai_1 _09421_ (.B1(_02411_),
    .Y(_02412_),
    .A1(net1928),
    .A2(net1924));
 sg13g2_xnor2_1 _09422_ (.Y(_02413_),
    .A(_02410_),
    .B(_02412_));
 sg13g2_nand2_1 _09423_ (.Y(_02414_),
    .A(net2234),
    .B(_02413_));
 sg13g2_xnor2_1 _09424_ (.Y(_02415_),
    .A(\vgadonut.donut.donuthit.ryin[11] ),
    .B(_02413_));
 sg13g2_nand3_1 _09425_ (.B(_02391_),
    .C(_02415_),
    .A(_02389_),
    .Y(_02416_));
 sg13g2_a21o_1 _09426_ (.A2(_02391_),
    .A1(_02389_),
    .B1(_02415_),
    .X(_02417_));
 sg13g2_nand3_1 _09427_ (.B(_02416_),
    .C(_02417_),
    .A(net1682),
    .Y(_02418_));
 sg13g2_o21ai_1 _09428_ (.B1(_02244_),
    .Y(_02419_),
    .A1(net1504),
    .A2(net1499));
 sg13g2_nand3_1 _09429_ (.B(_02360_),
    .C(_02419_),
    .A(net1494),
    .Y(_02420_));
 sg13g2_a22oi_1 _09430_ (.Y(_02421_),
    .B1(_02222_),
    .B2(net1527),
    .A2(_02220_),
    .A1(net1502));
 sg13g2_and4_2 _09431_ (.A(net1494),
    .B(_02360_),
    .C(_02419_),
    .D(_02421_),
    .X(_02422_));
 sg13g2_nor2_1 _09432_ (.A(_02365_),
    .B(_02422_),
    .Y(_02423_));
 sg13g2_nand2_1 _09433_ (.Y(_02424_),
    .A(_02365_),
    .B(_02422_));
 sg13g2_xor2_1 _09434_ (.B(_02422_),
    .A(_02365_),
    .X(_02425_));
 sg13g2_xnor2_1 _09435_ (.Y(_02426_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[6] ),
    .B(_02425_));
 sg13g2_a21oi_2 _09436_ (.B1(_02399_),
    .Y(_02427_),
    .A2(_02400_),
    .A1(net294));
 sg13g2_nor2_1 _09437_ (.A(_02426_),
    .B(_02427_),
    .Y(_02428_));
 sg13g2_or2_1 _09438_ (.X(_02429_),
    .B(_02427_),
    .A(_02426_));
 sg13g2_xnor2_1 _09439_ (.Y(_02430_),
    .A(_02426_),
    .B(_02427_));
 sg13g2_nor2_1 _09440_ (.A(_02375_),
    .B(_02404_),
    .Y(_02431_));
 sg13g2_a21o_1 _09441_ (.A2(_02402_),
    .A1(_02370_),
    .B1(_02403_),
    .X(_02432_));
 sg13g2_or2_1 _09442_ (.X(_02433_),
    .B(_02432_),
    .A(_02431_));
 sg13g2_nand2b_1 _09443_ (.Y(_02434_),
    .B(_02430_),
    .A_N(_02433_));
 sg13g2_nor2b_1 _09444_ (.A(_02430_),
    .B_N(_02433_),
    .Y(_02435_));
 sg13g2_nand2_1 _09445_ (.Y(_02436_),
    .A(net1676),
    .B(_02434_));
 sg13g2_o21ai_1 _09446_ (.B1(_02418_),
    .Y(_00074_),
    .A1(_02435_),
    .A2(_02436_));
 sg13g2_o21ai_1 _09447_ (.B1(_02408_),
    .Y(_02437_),
    .A1(_02409_),
    .A2(_02412_));
 sg13g2_xor2_1 _09448_ (.B(net1920),
    .A(net1924),
    .X(_02438_));
 sg13g2_xnor2_1 _09449_ (.Y(_02439_),
    .A(_02437_),
    .B(_02438_));
 sg13g2_nand2b_1 _09450_ (.Y(_02440_),
    .B(net2020),
    .A_N(_02439_));
 sg13g2_xnor2_1 _09451_ (.Y(_02441_),
    .A(_00551_),
    .B(_02439_));
 sg13g2_nand3_1 _09452_ (.B(_02417_),
    .C(_02441_),
    .A(_02414_),
    .Y(_02442_));
 sg13g2_a21o_1 _09453_ (.A2(_02417_),
    .A1(_02414_),
    .B1(_02441_),
    .X(_02443_));
 sg13g2_nand3_1 _09454_ (.B(_02442_),
    .C(_02443_),
    .A(net1681),
    .Y(_02444_));
 sg13g2_nor2_1 _09455_ (.A(_02428_),
    .B(_02435_),
    .Y(_02445_));
 sg13g2_a21oi_2 _09456_ (.B1(_02423_),
    .Y(_02446_),
    .A2(_02424_),
    .A1(\vgadonut.donut.donuthit.cordicxy.yin[6] ));
 sg13g2_a22oi_1 _09457_ (.Y(_02447_),
    .B1(_02244_),
    .B2(net1502),
    .A2(_02220_),
    .A1(net1527));
 sg13g2_and4_2 _09458_ (.A(net1494),
    .B(_02360_),
    .C(_02419_),
    .D(_02447_),
    .X(_02448_));
 sg13g2_nor2_1 _09459_ (.A(_02398_),
    .B(_02448_),
    .Y(_02449_));
 sg13g2_xnor2_1 _09460_ (.Y(_02450_),
    .A(_02398_),
    .B(_02448_));
 sg13g2_inv_1 _09461_ (.Y(_02451_),
    .A(_02450_));
 sg13g2_xnor2_1 _09462_ (.Y(_02452_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[7] ),
    .B(_02450_));
 sg13g2_nand2b_1 _09463_ (.Y(_02453_),
    .B(_02452_),
    .A_N(_02446_));
 sg13g2_nor2b_1 _09464_ (.A(_02452_),
    .B_N(_02446_),
    .Y(_02454_));
 sg13g2_xor2_1 _09465_ (.B(_02452_),
    .A(_02446_),
    .X(_02455_));
 sg13g2_xnor2_1 _09466_ (.Y(_02456_),
    .A(_02445_),
    .B(_02455_));
 sg13g2_o21ai_1 _09467_ (.B1(_02444_),
    .Y(_00075_),
    .A1(net1693),
    .A2(_02456_));
 sg13g2_nand2_1 _09468_ (.Y(_02457_),
    .A(net1922),
    .B(\vgadonut.donut.sAcB[14] ));
 sg13g2_nor2_1 _09469_ (.A(net1922),
    .B(\vgadonut.donut.sAcB[14] ),
    .Y(_02458_));
 sg13g2_xor2_1 _09470_ (.B(net1919),
    .A(net1922),
    .X(_02459_));
 sg13g2_a21o_1 _09471_ (.A2(net1920),
    .A1(net1924),
    .B1(_02437_),
    .X(_02460_));
 sg13g2_o21ai_1 _09472_ (.B1(_02460_),
    .Y(_02461_),
    .A1(net1924),
    .A2(net1920));
 sg13g2_xnor2_1 _09473_ (.Y(_02462_),
    .A(_02459_),
    .B(_02461_));
 sg13g2_xnor2_1 _09474_ (.Y(_02463_),
    .A(\vgadonut.donut.donuthit.ryin[13] ),
    .B(_02462_));
 sg13g2_nand3_1 _09475_ (.B(_02443_),
    .C(_02463_),
    .A(_02440_),
    .Y(_02464_));
 sg13g2_a21oi_1 _09476_ (.A1(_02440_),
    .A2(_02443_),
    .Y(_02465_),
    .B1(_02463_));
 sg13g2_nor2_1 _09477_ (.A(net1676),
    .B(_02465_),
    .Y(_02466_));
 sg13g2_nor2_1 _09478_ (.A(_02430_),
    .B(_02455_),
    .Y(_02467_));
 sg13g2_nor4_1 _09479_ (.A(_02371_),
    .B(_02404_),
    .C(_02430_),
    .D(_02455_),
    .Y(_02468_));
 sg13g2_o21ai_1 _09480_ (.B1(_02453_),
    .Y(_02469_),
    .A1(_02429_),
    .A2(_02454_));
 sg13g2_a221oi_1 _09481_ (.B2(_02468_),
    .C1(_02469_),
    .B1(_02374_),
    .A1(_02432_),
    .Y(_02470_),
    .A2(_02467_));
 sg13g2_nor2_2 _09482_ (.A(net1522),
    .B(_02243_),
    .Y(_02471_));
 sg13g2_nor2_2 _09483_ (.A(_02420_),
    .B(_02471_),
    .Y(_02472_));
 sg13g2_or2_1 _09484_ (.X(_02473_),
    .B(_02472_),
    .A(_02422_));
 sg13g2_xnor2_1 _09485_ (.Y(_02474_),
    .A(_02422_),
    .B(_02472_));
 sg13g2_inv_1 _09486_ (.Y(_02475_),
    .A(_02474_));
 sg13g2_nand2_1 _09487_ (.Y(_02476_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[8] ),
    .B(_02475_));
 sg13g2_xor2_1 _09488_ (.B(_02474_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[8] ),
    .X(_02477_));
 sg13g2_a21oi_1 _09489_ (.A1(\vgadonut.donut.donuthit.cordicxy.yin[7] ),
    .A2(_02451_),
    .Y(_02478_),
    .B1(_02449_));
 sg13g2_nor2_1 _09490_ (.A(_02477_),
    .B(_02478_),
    .Y(_02479_));
 sg13g2_xnor2_1 _09491_ (.Y(_02480_),
    .A(_02477_),
    .B(_02478_));
 sg13g2_or2_1 _09492_ (.X(_02481_),
    .B(_02470_),
    .A(_02480_));
 sg13g2_a21oi_1 _09493_ (.A1(_02470_),
    .A2(_02480_),
    .Y(_02482_),
    .B1(net1693));
 sg13g2_a22oi_1 _09494_ (.Y(_02483_),
    .B1(_02481_),
    .B2(_02482_),
    .A2(_02466_),
    .A1(_02464_));
 sg13g2_inv_1 _09495_ (.Y(_00076_),
    .A(_02483_));
 sg13g2_nor2_1 _09496_ (.A(_02448_),
    .B(_02472_),
    .Y(_02484_));
 sg13g2_xnor2_1 _09497_ (.Y(_02485_),
    .A(_02448_),
    .B(_02472_));
 sg13g2_inv_1 _09498_ (.Y(_02486_),
    .A(_02485_));
 sg13g2_xor2_1 _09499_ (.B(_02485_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[9] ),
    .X(_02487_));
 sg13g2_a21oi_1 _09500_ (.A1(_02473_),
    .A2(_02476_),
    .Y(_02488_),
    .B1(_02487_));
 sg13g2_nand3_1 _09501_ (.B(_02476_),
    .C(_02487_),
    .A(_02473_),
    .Y(_02489_));
 sg13g2_inv_1 _09502_ (.Y(_02490_),
    .A(_02489_));
 sg13g2_nor2_1 _09503_ (.A(_02488_),
    .B(_02490_),
    .Y(_02491_));
 sg13g2_nor2b_1 _09504_ (.A(_02479_),
    .B_N(_02481_),
    .Y(_02492_));
 sg13g2_xor2_1 _09505_ (.B(_02492_),
    .A(_02491_),
    .X(_02493_));
 sg13g2_a21oi_1 _09506_ (.A1(_00556_),
    .A2(_02462_),
    .Y(_02494_),
    .B1(_02465_));
 sg13g2_xnor2_1 _09507_ (.Y(_02495_),
    .A(net1921),
    .B(\vgadonut.donut.sAcB[15] ));
 sg13g2_o21ai_1 _09508_ (.B1(_02457_),
    .Y(_02496_),
    .A1(_02458_),
    .A2(_02461_));
 sg13g2_xnor2_1 _09509_ (.Y(_02497_),
    .A(_02495_),
    .B(_02496_));
 sg13g2_nand2_1 _09510_ (.Y(_02498_),
    .A(\vgadonut.donut.donuthit.ryin[14] ),
    .B(_02497_));
 sg13g2_nor2_1 _09511_ (.A(\vgadonut.donut.donuthit.ryin[14] ),
    .B(_02497_),
    .Y(_02499_));
 sg13g2_xnor2_1 _09512_ (.Y(_02500_),
    .A(\vgadonut.donut.donuthit.ryin[14] ),
    .B(_02497_));
 sg13g2_a21oi_1 _09513_ (.A1(_02494_),
    .A2(_02500_),
    .Y(_02501_),
    .B1(net1676));
 sg13g2_o21ai_1 _09514_ (.B1(_02501_),
    .Y(_02502_),
    .A1(_02494_),
    .A2(_02500_));
 sg13g2_o21ai_1 _09515_ (.B1(_02502_),
    .Y(_00077_),
    .A1(net1693),
    .A2(_02493_));
 sg13g2_a21oi_1 _09516_ (.A1(\vgadonut.donut.donuthit.cordicxy.yin[9] ),
    .A2(_02486_),
    .Y(_02503_),
    .B1(_02484_));
 sg13g2_nor2b_1 _09517_ (.A(_02503_),
    .B_N(\vgadonut.donut.donuthit.cordicxy.yin[10] ),
    .Y(_02504_));
 sg13g2_xnor2_1 _09518_ (.Y(_02505_),
    .A(\vgadonut.donut.donuthit.cordicxy.yin[10] ),
    .B(_02503_));
 sg13g2_nor2_1 _09519_ (.A(_02479_),
    .B(_02488_),
    .Y(_02506_));
 sg13g2_a21oi_2 _09520_ (.B1(_02490_),
    .Y(_02507_),
    .A2(_02481_),
    .A1(_02506_));
 sg13g2_xnor2_1 _09521_ (.Y(_02508_),
    .A(_02505_),
    .B(_02507_));
 sg13g2_nand2_1 _09522_ (.Y(_02509_),
    .A(net1919),
    .B(net1918));
 sg13g2_nor2_1 _09523_ (.A(net1919),
    .B(net1918),
    .Y(_02510_));
 sg13g2_xor2_1 _09524_ (.B(net1918),
    .A(net1919),
    .X(_02511_));
 sg13g2_a21o_1 _09525_ (.A2(net1918),
    .A1(net1920),
    .B1(_02496_),
    .X(_02512_));
 sg13g2_o21ai_1 _09526_ (.B1(_02512_),
    .Y(_02513_),
    .A1(net1920),
    .A2(net1918));
 sg13g2_xnor2_1 _09527_ (.Y(_02514_),
    .A(_02511_),
    .B(_02513_));
 sg13g2_xnor2_1 _09528_ (.Y(_02515_),
    .A(_00559_),
    .B(_02514_));
 sg13g2_o21ai_1 _09529_ (.B1(_02498_),
    .Y(_02516_),
    .A1(_02494_),
    .A2(_02499_));
 sg13g2_and2_1 _09530_ (.A(_02515_),
    .B(_02516_),
    .X(_02517_));
 sg13g2_o21ai_1 _09531_ (.B1(net1693),
    .Y(_02518_),
    .A1(_02515_),
    .A2(_02516_));
 sg13g2_or2_1 _09532_ (.X(_02519_),
    .B(_02518_),
    .A(_02517_));
 sg13g2_o21ai_1 _09533_ (.B1(_02519_),
    .Y(_00063_),
    .A1(_02508_),
    .A2(net1692));
 sg13g2_a21o_1 _09534_ (.A2(_02514_),
    .A1(_00637_),
    .B1(_02517_),
    .X(_02520_));
 sg13g2_o21ai_1 _09535_ (.B1(_02509_),
    .Y(_02521_),
    .A1(_02510_),
    .A2(_02513_));
 sg13g2_xnor2_1 _09536_ (.Y(_02522_),
    .A(\vgadonut.donut.donuthit.ryin[15] ),
    .B(_02521_));
 sg13g2_or2_1 _09537_ (.X(_02523_),
    .B(_02522_),
    .A(_02520_));
 sg13g2_a21oi_1 _09538_ (.A1(_02520_),
    .A2(_02522_),
    .Y(_02524_),
    .B1(net1676));
 sg13g2_nor2b_1 _09539_ (.A(_02472_),
    .B_N(_00164_),
    .Y(_02525_));
 sg13g2_xor2_1 _09540_ (.B(_02472_),
    .A(_00164_),
    .X(_02526_));
 sg13g2_inv_2 _09541_ (.Y(_02527_),
    .A(_02526_));
 sg13g2_a21oi_2 _09542_ (.B1(_02504_),
    .Y(_02528_),
    .A2(_02505_),
    .A1(_02507_));
 sg13g2_nor2_1 _09543_ (.A(_02527_),
    .B(_02528_),
    .Y(_02529_));
 sg13g2_xnor2_1 _09544_ (.Y(_02530_),
    .A(_02527_),
    .B(_02528_));
 sg13g2_a22oi_1 _09545_ (.Y(_00064_),
    .B1(net1676),
    .B2(_02530_),
    .A2(_02524_),
    .A1(_02523_));
 sg13g2_and2_1 _09546_ (.A(_00637_),
    .B(_02521_),
    .X(_02531_));
 sg13g2_nor3_1 _09547_ (.A(_02520_),
    .B(_02522_),
    .C(_02531_),
    .Y(_02532_));
 sg13g2_and3_1 _09548_ (.X(_02533_),
    .A(\vgadonut.donut.donuthit.ryin[15] ),
    .B(_00637_),
    .C(_02521_));
 sg13g2_o21ai_1 _09549_ (.B1(net1692),
    .Y(_02534_),
    .A1(_02532_),
    .A2(_02533_));
 sg13g2_xnor2_1 _09550_ (.Y(_02535_),
    .A(net2329),
    .B(_02525_));
 sg13g2_inv_1 _09551_ (.Y(_02536_),
    .A(_02535_));
 sg13g2_nor2_1 _09552_ (.A(_02529_),
    .B(_02535_),
    .Y(_02537_));
 sg13g2_nand2_1 _09553_ (.Y(_02538_),
    .A(_02529_),
    .B(_02535_));
 sg13g2_nand2_1 _09554_ (.Y(_02539_),
    .A(net1680),
    .B(_02538_));
 sg13g2_o21ai_1 _09555_ (.B1(_02534_),
    .Y(_00065_),
    .A1(_02537_),
    .A2(_02539_));
 sg13g2_o21ai_1 _09556_ (.B1(_00166_),
    .Y(_02540_),
    .A1(_02420_),
    .A2(_02471_));
 sg13g2_o21ai_1 _09557_ (.B1(_02538_),
    .Y(_02541_),
    .A1(net2359),
    .A2(_02540_));
 sg13g2_xnor2_1 _09558_ (.Y(_02542_),
    .A(net2307),
    .B(_02540_));
 sg13g2_xor2_1 _09559_ (.B(_02542_),
    .A(_02541_),
    .X(_02543_));
 sg13g2_o21ai_1 _09560_ (.B1(_02534_),
    .Y(_00066_),
    .A1(net1698),
    .A2(_02543_));
 sg13g2_or4_1 _09561_ (.A(_02527_),
    .B(_02528_),
    .C(_02536_),
    .D(_02542_),
    .X(_02544_));
 sg13g2_nand2_1 _09562_ (.Y(_02545_),
    .A(_00164_),
    .B(net2357));
 sg13g2_nor2_1 _09563_ (.A(_00638_),
    .B(_02472_),
    .Y(_02546_));
 sg13g2_nand2_1 _09564_ (.Y(_02547_),
    .A(_02545_),
    .B(_02546_));
 sg13g2_nor2b_1 _09565_ (.A(_02472_),
    .B_N(_00168_),
    .Y(_02548_));
 sg13g2_xor2_1 _09566_ (.B(_02546_),
    .A(net2253),
    .X(_02549_));
 sg13g2_nand3_1 _09567_ (.B(_02547_),
    .C(_02549_),
    .A(_02544_),
    .Y(_02550_));
 sg13g2_a21oi_1 _09568_ (.A1(_02544_),
    .A2(_02547_),
    .Y(_02551_),
    .B1(_02549_));
 sg13g2_nand2_1 _09569_ (.Y(_02552_),
    .A(net1680),
    .B(_02550_));
 sg13g2_o21ai_1 _09570_ (.B1(_02534_),
    .Y(_00067_),
    .A1(_02551_),
    .A2(_02552_));
 sg13g2_a21oi_1 _09571_ (.A1(_00638_),
    .A2(_02548_),
    .Y(_02553_),
    .B1(_02551_));
 sg13g2_xor2_1 _09572_ (.B(_02548_),
    .A(net2321),
    .X(_02554_));
 sg13g2_xnor2_1 _09573_ (.Y(_02555_),
    .A(_02553_),
    .B(_02554_));
 sg13g2_o21ai_1 _09574_ (.B1(_02534_),
    .Y(_00068_),
    .A1(net1698),
    .A2(_02555_));
 sg13g2_xnor2_1 _09575_ (.Y(_02556_),
    .A(\vgadonut.donut.cAcB[1] ),
    .B(\vgadonut.donut.cAcB[3] ));
 sg13g2_nor2_1 _09576_ (.A(\vgadonut.donut.cAcB[2] ),
    .B(net1953),
    .Y(_02557_));
 sg13g2_nor2_1 _09577_ (.A(\vgadonut.donut.cAcB[0] ),
    .B(net1955),
    .Y(_02558_));
 sg13g2_nand3_1 _09578_ (.B(_02557_),
    .C(_02558_),
    .A(_02556_),
    .Y(_02559_));
 sg13g2_nor2_2 _09579_ (.A(net1957),
    .B(net1954),
    .Y(_02560_));
 sg13g2_nand2_1 _09580_ (.Y(_02561_),
    .A(\vgadonut.donut.cAcB[0] ),
    .B(net1955));
 sg13g2_nand2_1 _09581_ (.Y(_02562_),
    .A(\vgadonut.donut.cAcB[2] ),
    .B(net1955));
 sg13g2_o21ai_1 _09582_ (.B1(net1957),
    .Y(_02563_),
    .A1(\vgadonut.donut.cAcB[1] ),
    .A2(net1953));
 sg13g2_a22oi_1 _09583_ (.Y(_02564_),
    .B1(_02562_),
    .B2(_02563_),
    .A2(_02561_),
    .A1(_02557_));
 sg13g2_o21ai_1 _09584_ (.B1(_02559_),
    .Y(_02565_),
    .A1(_02560_),
    .A2(_02564_));
 sg13g2_xor2_1 _09585_ (.B(net1951),
    .A(net1955),
    .X(_02566_));
 sg13g2_xnor2_1 _09586_ (.Y(_02567_),
    .A(_02560_),
    .B(_02566_));
 sg13g2_nor2b_1 _09587_ (.A(_02567_),
    .B_N(_02565_),
    .Y(_02568_));
 sg13g2_xnor2_1 _09588_ (.Y(_02569_),
    .A(_02565_),
    .B(_02567_));
 sg13g2_nand2_1 _09589_ (.Y(_02570_),
    .A(\vgadonut.donut.donuthit.rzin[5] ),
    .B(_02569_));
 sg13g2_or2_1 _09590_ (.X(_02571_),
    .B(_02569_),
    .A(\vgadonut.donut.donuthit.rzin[5] ));
 sg13g2_a21oi_2 _09591_ (.B1(net1673),
    .Y(_02572_),
    .A2(_02571_),
    .A1(_02570_));
 sg13g2_xor2_1 _09592_ (.B(net1538),
    .A(\vgadonut.donut.donuthit.rz[14] ),
    .X(_02573_));
 sg13g2_xnor2_1 _09593_ (.Y(_02574_),
    .A(\vgadonut.donut.donuthit.rz[14] ),
    .B(net1538));
 sg13g2_xnor2_1 _09594_ (.Y(_02575_),
    .A(\vgadonut.donut.donuthit.rz[13] ),
    .B(net1538));
 sg13g2_xor2_1 _09595_ (.B(net1538),
    .A(\vgadonut.donut.donuthit.rz[13] ),
    .X(_02576_));
 sg13g2_xnor2_1 _09596_ (.Y(_02577_),
    .A(\vgadonut.donut.donuthit.rz[10] ),
    .B(net1538));
 sg13g2_nand3_1 _09597_ (.B(net1509),
    .C(_02577_),
    .A(net1518),
    .Y(_02578_));
 sg13g2_xnor2_1 _09598_ (.Y(_02579_),
    .A(\vgadonut.donut.donuthit.rz[7] ),
    .B(net1534));
 sg13g2_nand2_1 _09599_ (.Y(_02580_),
    .A(net1528),
    .B(_02579_));
 sg13g2_xnor2_1 _09600_ (.Y(_02581_),
    .A(\vgadonut.donut.donuthit.rz[8] ),
    .B(net1534));
 sg13g2_nand3_1 _09601_ (.B(net1524),
    .C(_02581_),
    .A(net1531),
    .Y(_02582_));
 sg13g2_xnor2_1 _09602_ (.Y(_02583_),
    .A(\vgadonut.donut.donuthit.rz[9] ),
    .B(net1538));
 sg13g2_nand3_1 _09603_ (.B(net1513),
    .C(_02583_),
    .A(net1517),
    .Y(_02584_));
 sg13g2_nand4_1 _09604_ (.B(_02580_),
    .C(_02582_),
    .A(_02578_),
    .Y(_02585_),
    .D(_02584_));
 sg13g2_xnor2_1 _09605_ (.Y(_02586_),
    .A(\vgadonut.donut.donuthit.rz[12] ),
    .B(net1538));
 sg13g2_nand4_1 _09606_ (.B(net1511),
    .C(_01876_),
    .A(net1518),
    .Y(_02587_),
    .D(_02586_));
 sg13g2_xnor2_1 _09607_ (.Y(_02588_),
    .A(\vgadonut.donut.donuthit.rz[11] ),
    .B(net1538));
 sg13g2_xor2_1 _09608_ (.B(net1534),
    .A(\vgadonut.donut.donuthit.rz[11] ),
    .X(_02589_));
 sg13g2_nand4_1 _09609_ (.B(net1511),
    .C(_01845_),
    .A(net1517),
    .Y(_02590_),
    .D(_02588_));
 sg13g2_o21ai_1 _09610_ (.B1(_02587_),
    .Y(_02591_),
    .A1(_01856_),
    .A2(_02576_));
 sg13g2_o21ai_1 _09611_ (.B1(_02590_),
    .Y(_02592_),
    .A1(_01884_),
    .A2(_02573_));
 sg13g2_nand2_1 _09612_ (.Y(_02593_),
    .A(\vgadonut.donut.donuthit.rz[15] ),
    .B(net1539));
 sg13g2_or2_1 _09613_ (.X(_02594_),
    .B(net1539),
    .A(\vgadonut.donut.donuthit.rz[15] ));
 sg13g2_and2_2 _09614_ (.A(_02593_),
    .B(_02594_),
    .X(_02595_));
 sg13g2_nand2_2 _09615_ (.Y(_02596_),
    .A(_02593_),
    .B(_02594_));
 sg13g2_o21ai_1 _09616_ (.B1(_02596_),
    .Y(_02597_),
    .A1(_01897_),
    .A2(_01899_));
 sg13g2_a221oi_1 _09617_ (.B2(_02594_),
    .C1(net1508),
    .B1(_02593_),
    .A1(_01896_),
    .Y(_02598_),
    .A2(_01900_));
 sg13g2_nor4_2 _09618_ (.A(_02585_),
    .B(_02591_),
    .C(_02592_),
    .Y(_02599_),
    .D(_02598_));
 sg13g2_nand3_1 _09619_ (.B(net1513),
    .C(_02579_),
    .A(net1517),
    .Y(_02600_));
 sg13g2_nand3_1 _09620_ (.B(net1509),
    .C(_02581_),
    .A(net1517),
    .Y(_02601_));
 sg13g2_nor2_1 _09621_ (.A(\vgadonut.donut.donuthit.rz[5] ),
    .B(_01816_),
    .Y(_02602_));
 sg13g2_a21oi_1 _09622_ (.A1(\vgadonut.donut.donuthit.rz[5] ),
    .A2(_01817_),
    .Y(_02603_),
    .B1(_02602_));
 sg13g2_xnor2_1 _09623_ (.Y(_02604_),
    .A(\vgadonut.donut.donuthit.rz[6] ),
    .B(net1534));
 sg13g2_nand3_1 _09624_ (.B(net1524),
    .C(_02604_),
    .A(net1530),
    .Y(_02605_));
 sg13g2_nand4_1 _09625_ (.B(_02601_),
    .C(_02603_),
    .A(_02600_),
    .Y(_02606_),
    .D(_02605_));
 sg13g2_nor3_1 _09626_ (.A(net1508),
    .B(_01896_),
    .C(_02573_),
    .Y(_02607_));
 sg13g2_nor2_1 _09627_ (.A(_01856_),
    .B(_02589_),
    .Y(_02608_));
 sg13g2_nor4_1 _09628_ (.A(_01807_),
    .B(net1508),
    .C(_01898_),
    .D(_02576_),
    .Y(_02609_));
 sg13g2_a221oi_1 _09629_ (.B2(_01873_),
    .C1(_02608_),
    .B1(_02583_),
    .A1(_01877_),
    .Y(_02610_),
    .A2(_02577_));
 sg13g2_nor2b_1 _09630_ (.A(_01884_),
    .B_N(_02586_),
    .Y(_02611_));
 sg13g2_nor4_1 _09631_ (.A(_02606_),
    .B(_02607_),
    .C(_02609_),
    .D(_02611_),
    .Y(_02612_));
 sg13g2_a21oi_1 _09632_ (.A1(_02610_),
    .A2(_02612_),
    .Y(_02613_),
    .B1(_02599_));
 sg13g2_nand3_1 _09633_ (.B(_02610_),
    .C(_02612_),
    .A(_02599_),
    .Y(_02614_));
 sg13g2_nand2b_1 _09634_ (.Y(_02615_),
    .B(_02614_),
    .A_N(_02613_));
 sg13g2_xnor2_1 _09635_ (.Y(_02616_),
    .A(net2094),
    .B(_02615_));
 sg13g2_a21oi_1 _09636_ (.A1(net1679),
    .A2(_02616_),
    .Y(_00078_),
    .B1(_02572_));
 sg13g2_nand2_1 _09637_ (.Y(_02617_),
    .A(_01855_),
    .B(_02574_));
 sg13g2_nand3_1 _09638_ (.B(net1513),
    .C(_02577_),
    .A(net1518),
    .Y(_02618_));
 sg13g2_nand3_1 _09639_ (.B(net1509),
    .C(_02588_),
    .A(net1518),
    .Y(_02619_));
 sg13g2_nand2_1 _09640_ (.Y(_02620_),
    .A(net1529),
    .B(_02581_));
 sg13g2_nand3_1 _09641_ (.B(net1524),
    .C(_02583_),
    .A(net1530),
    .Y(_02621_));
 sg13g2_and4_1 _09642_ (.A(_02618_),
    .B(_02619_),
    .C(_02620_),
    .D(_02621_),
    .X(_02622_));
 sg13g2_a22oi_1 _09643_ (.Y(_02623_),
    .B1(_02586_),
    .B2(_01873_),
    .A2(_02575_),
    .A1(net1497));
 sg13g2_nand2b_1 _09644_ (.Y(_02624_),
    .B(_02596_),
    .A_N(_01884_));
 sg13g2_and4_2 _09645_ (.A(_02617_),
    .B(_02622_),
    .C(_02623_),
    .D(_02624_),
    .X(_02625_));
 sg13g2_nand2_1 _09646_ (.Y(_02626_),
    .A(_02597_),
    .B(_02625_));
 sg13g2_nand3_1 _09647_ (.B(net1509),
    .C(_02583_),
    .A(net1517),
    .Y(_02627_));
 sg13g2_nand3_1 _09648_ (.B(net1513),
    .C(_02581_),
    .A(net1517),
    .Y(_02628_));
 sg13g2_nand3_1 _09649_ (.B(net1524),
    .C(_02579_),
    .A(net1530),
    .Y(_02629_));
 sg13g2_nand2_1 _09650_ (.Y(_02630_),
    .A(net1528),
    .B(_02604_));
 sg13g2_nand4_1 _09651_ (.B(_02628_),
    .C(_02629_),
    .A(_02627_),
    .Y(_02631_),
    .D(_02630_));
 sg13g2_nor2_1 _09652_ (.A(_01878_),
    .B(_02589_),
    .Y(_02632_));
 sg13g2_nor3_1 _09653_ (.A(net1508),
    .B(net1495),
    .C(_02595_),
    .Y(_02633_));
 sg13g2_nor4_1 _09654_ (.A(_01807_),
    .B(net1508),
    .C(_01898_),
    .D(_02573_),
    .Y(_02634_));
 sg13g2_nor2_1 _09655_ (.A(net1496),
    .B(_02576_),
    .Y(_02635_));
 sg13g2_a221oi_1 _09656_ (.B2(_01855_),
    .C1(_02635_),
    .B1(_02586_),
    .A1(_01873_),
    .Y(_02636_),
    .A2(_02577_));
 sg13g2_nor4_2 _09657_ (.A(_02631_),
    .B(_02632_),
    .C(_02633_),
    .Y(_02637_),
    .D(_02634_));
 sg13g2_and4_1 _09658_ (.A(_02597_),
    .B(_02625_),
    .C(_02636_),
    .D(_02637_),
    .X(_02638_));
 sg13g2_nand4_1 _09659_ (.B(_02625_),
    .C(_02636_),
    .A(_02597_),
    .Y(_02639_),
    .D(_02637_));
 sg13g2_a22oi_1 _09660_ (.Y(_02640_),
    .B1(_02636_),
    .B2(_02637_),
    .A2(_02625_),
    .A1(_02597_));
 sg13g2_o21ai_1 _09661_ (.B1(_00635_),
    .Y(_02641_),
    .A1(_02638_),
    .A2(_02640_));
 sg13g2_nand3b_1 _09662_ (.B(_00153_),
    .C(_02639_),
    .Y(_02642_),
    .A_N(_02640_));
 sg13g2_o21ai_1 _09663_ (.B1(_02614_),
    .Y(_02643_),
    .A1(net2290),
    .A2(_02613_));
 sg13g2_a21oi_2 _09664_ (.B1(_02643_),
    .Y(_02644_),
    .A2(_02642_),
    .A1(_02641_));
 sg13g2_nand3_1 _09665_ (.B(_02642_),
    .C(_02643_),
    .A(_02641_),
    .Y(_02645_));
 sg13g2_nand2b_1 _09666_ (.Y(_02646_),
    .B(_02645_),
    .A_N(_02644_));
 sg13g2_a21oi_2 _09667_ (.B1(_02568_),
    .Y(_02647_),
    .A2(_02566_),
    .A1(_02560_));
 sg13g2_nor2_1 _09668_ (.A(net1953),
    .B(net1950),
    .Y(_02648_));
 sg13g2_xnor2_1 _09669_ (.Y(_02649_),
    .A(net1953),
    .B(net1949));
 sg13g2_or3_1 _09670_ (.A(net1956),
    .B(net1951),
    .C(_02649_),
    .X(_02650_));
 sg13g2_o21ai_1 _09671_ (.B1(_02649_),
    .Y(_02651_),
    .A1(net1956),
    .A2(net1951));
 sg13g2_nand2_1 _09672_ (.Y(_02652_),
    .A(_02650_),
    .B(_02651_));
 sg13g2_xor2_1 _09673_ (.B(_02652_),
    .A(_02647_),
    .X(_02653_));
 sg13g2_nand2_1 _09674_ (.Y(_02654_),
    .A(\vgadonut.donut.donuthit.rzin[6] ),
    .B(_02653_));
 sg13g2_xnor2_1 _09675_ (.Y(_02655_),
    .A(\vgadonut.donut.donuthit.rzin[6] ),
    .B(_02653_));
 sg13g2_or2_1 _09676_ (.X(_02656_),
    .B(_02655_),
    .A(_02570_));
 sg13g2_a21oi_1 _09677_ (.A1(_02570_),
    .A2(_02655_),
    .Y(_02657_),
    .B1(net1673));
 sg13g2_nand2_2 _09678_ (.Y(_02658_),
    .A(_02656_),
    .B(_02657_));
 sg13g2_o21ai_1 _09679_ (.B1(_02658_),
    .Y(_00085_),
    .A1(net1700),
    .A2(net2292));
 sg13g2_a21oi_2 _09680_ (.B1(_02595_),
    .Y(_02659_),
    .A2(_01972_),
    .A1(_01901_));
 sg13g2_o21ai_1 _09681_ (.B1(_02596_),
    .Y(_02660_),
    .A1(_01973_),
    .A2(_01902_));
 sg13g2_nand3_1 _09682_ (.B(net1513),
    .C(_02588_),
    .A(net1517),
    .Y(_02661_));
 sg13g2_nand2_1 _09683_ (.Y(_02662_),
    .A(net1528),
    .B(_02583_));
 sg13g2_nand3_1 _09684_ (.B(net1524),
    .C(_02577_),
    .A(net1530),
    .Y(_02663_));
 sg13g2_nand3_1 _09685_ (.B(_02662_),
    .C(_02663_),
    .A(_02661_),
    .Y(_02664_));
 sg13g2_and2_1 _09686_ (.A(net1501),
    .B(_02586_),
    .X(_02665_));
 sg13g2_nor2_1 _09687_ (.A(_01878_),
    .B(_02573_),
    .Y(_02666_));
 sg13g2_and2_1 _09688_ (.A(net1498),
    .B(_02575_),
    .X(_02667_));
 sg13g2_nor4_2 _09689_ (.A(_02664_),
    .B(_02665_),
    .C(_02666_),
    .Y(_02668_),
    .D(_02667_));
 sg13g2_or4_1 _09690_ (.A(_02664_),
    .B(_02665_),
    .C(_02666_),
    .D(_02667_),
    .X(_02669_));
 sg13g2_a21oi_1 _09691_ (.A1(net1493),
    .A2(_02668_),
    .Y(_02670_),
    .B1(_02599_));
 sg13g2_a21o_1 _09692_ (.A2(_02668_),
    .A1(net1493),
    .B1(_02599_),
    .X(_02671_));
 sg13g2_nand3_1 _09693_ (.B(net1493),
    .C(_02668_),
    .A(_02599_),
    .Y(_02672_));
 sg13g2_and3_1 _09694_ (.X(_02673_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[2] ),
    .B(_02671_),
    .C(_02672_));
 sg13g2_a21oi_1 _09695_ (.A1(_02671_),
    .A2(_02672_),
    .Y(_02674_),
    .B1(\vgadonut.donut.donuthit.cordicxz.xin[2] ));
 sg13g2_a21oi_1 _09696_ (.A1(\vgadonut.donut.donuthit.cordicxz.xin[1] ),
    .A2(_02639_),
    .Y(_02675_),
    .B1(_02640_));
 sg13g2_nor3_2 _09697_ (.A(_02673_),
    .B(_02674_),
    .C(_02675_),
    .Y(_02676_));
 sg13g2_o21ai_1 _09698_ (.B1(_02675_),
    .Y(_02677_),
    .A1(_02674_),
    .A2(_02673_));
 sg13g2_nor2b_1 _09699_ (.A(_02676_),
    .B_N(_02677_),
    .Y(_02678_));
 sg13g2_nand3b_1 _09700_ (.B(_02644_),
    .C(_02677_),
    .Y(_02679_),
    .A_N(_02676_));
 sg13g2_xnor2_1 _09701_ (.Y(_02680_),
    .A(net2291),
    .B(_02678_));
 sg13g2_o21ai_1 _09702_ (.B1(_02650_),
    .Y(_02681_),
    .A1(_02647_),
    .A2(_02652_));
 sg13g2_nor2_1 _09703_ (.A(net1951),
    .B(\vgadonut.donut.cAcB[8] ),
    .Y(_02682_));
 sg13g2_xor2_1 _09704_ (.B(\vgadonut.donut.cAcB[8] ),
    .A(net1951),
    .X(_02683_));
 sg13g2_nand2_1 _09705_ (.Y(_02684_),
    .A(_02648_),
    .B(_02683_));
 sg13g2_xnor2_1 _09706_ (.Y(_02685_),
    .A(_02648_),
    .B(_02683_));
 sg13g2_nand2b_1 _09707_ (.Y(_02686_),
    .B(_02681_),
    .A_N(_02685_));
 sg13g2_xnor2_1 _09708_ (.Y(_02687_),
    .A(_02681_),
    .B(_02685_));
 sg13g2_nand2_1 _09709_ (.Y(_02688_),
    .A(\vgadonut.donut.donuthit.rzin[7] ),
    .B(_02687_));
 sg13g2_xnor2_1 _09710_ (.Y(_02689_),
    .A(\vgadonut.donut.donuthit.rzin[7] ),
    .B(_02687_));
 sg13g2_a21o_1 _09711_ (.A2(_02656_),
    .A1(_02654_),
    .B1(_02689_),
    .X(_02690_));
 sg13g2_nand3_1 _09712_ (.B(_02656_),
    .C(_02689_),
    .A(_02654_),
    .Y(_02691_));
 sg13g2_nand3_1 _09713_ (.B(_02690_),
    .C(_02691_),
    .A(net1689),
    .Y(_02692_));
 sg13g2_o21ai_1 _09714_ (.B1(_02692_),
    .Y(_00086_),
    .A1(net1700),
    .A2(_02680_));
 sg13g2_xor2_1 _09715_ (.B(net1946),
    .A(net1949),
    .X(_02693_));
 sg13g2_xnor2_1 _09716_ (.Y(_02694_),
    .A(_02682_),
    .B(_02693_));
 sg13g2_a21oi_1 _09717_ (.A1(_02684_),
    .A2(_02686_),
    .Y(_02695_),
    .B1(_02694_));
 sg13g2_nand3_1 _09718_ (.B(_02686_),
    .C(_02694_),
    .A(_02684_),
    .Y(_02696_));
 sg13g2_nor2b_1 _09719_ (.A(_02695_),
    .B_N(_02696_),
    .Y(_02697_));
 sg13g2_nand2_1 _09720_ (.Y(_02698_),
    .A(\vgadonut.donut.donuthit.rzin[8] ),
    .B(_02697_));
 sg13g2_xnor2_1 _09721_ (.Y(_02699_),
    .A(\vgadonut.donut.donuthit.rzin[8] ),
    .B(_02697_));
 sg13g2_a21o_1 _09722_ (.A2(_02690_),
    .A1(_02688_),
    .B1(_02699_),
    .X(_02700_));
 sg13g2_nand3_1 _09723_ (.B(_02690_),
    .C(_02699_),
    .A(_02688_),
    .Y(_02701_));
 sg13g2_a21oi_2 _09724_ (.B1(net1673),
    .Y(_02702_),
    .A2(_02701_),
    .A1(_02700_));
 sg13g2_or2_1 _09725_ (.X(_02703_),
    .B(_02673_),
    .A(_02670_));
 sg13g2_nand2_1 _09726_ (.Y(_02704_),
    .A(net1506),
    .B(_02586_));
 sg13g2_a22oi_1 _09727_ (.Y(_02705_),
    .B1(_02588_),
    .B2(net1503),
    .A2(_02577_),
    .A1(net1528));
 sg13g2_nand2_1 _09728_ (.Y(_02706_),
    .A(net1497),
    .B(_02596_));
 sg13g2_a22oi_1 _09729_ (.Y(_02707_),
    .B1(_02575_),
    .B2(net1501),
    .A2(_02574_),
    .A1(net1498));
 sg13g2_and4_2 _09730_ (.A(_02704_),
    .B(_02705_),
    .C(_02706_),
    .D(_02707_),
    .X(_02708_));
 sg13g2_nand2_1 _09731_ (.Y(_02709_),
    .A(net1493),
    .B(_02708_));
 sg13g2_nand4_1 _09732_ (.B(_02625_),
    .C(net1493),
    .A(_02597_),
    .Y(_02710_),
    .D(_02708_));
 sg13g2_a22oi_1 _09733_ (.Y(_02711_),
    .B1(net1493),
    .B2(_02708_),
    .A2(_02625_),
    .A1(_02597_));
 sg13g2_xor2_1 _09734_ (.B(_02709_),
    .A(_02626_),
    .X(_02712_));
 sg13g2_xnor2_1 _09735_ (.Y(_02713_),
    .A(_00151_),
    .B(_02712_));
 sg13g2_nor2_1 _09736_ (.A(_02703_),
    .B(_02713_),
    .Y(_02714_));
 sg13g2_xnor2_1 _09737_ (.Y(_02715_),
    .A(_02703_),
    .B(_02713_));
 sg13g2_a21oi_1 _09738_ (.A1(_02644_),
    .A2(_02677_),
    .Y(_02716_),
    .B1(_02676_));
 sg13g2_xnor2_1 _09739_ (.Y(_02717_),
    .A(_02715_),
    .B(_02716_));
 sg13g2_a21oi_1 _09740_ (.A1(net1679),
    .A2(_02717_),
    .Y(_00087_),
    .B1(_02702_));
 sg13g2_nand2b_2 _09741_ (.Y(_02718_),
    .B(_02596_),
    .A_N(_01852_));
 sg13g2_nand2_1 _09742_ (.Y(_02719_),
    .A(net1501),
    .B(_02574_));
 sg13g2_nand2_1 _09743_ (.Y(_02720_),
    .A(net1528),
    .B(_02588_));
 sg13g2_a22oi_1 _09744_ (.Y(_02721_),
    .B1(_02586_),
    .B2(net1503),
    .A2(_02575_),
    .A1(net1506));
 sg13g2_and4_1 _09745_ (.A(_02718_),
    .B(_02719_),
    .C(_02720_),
    .D(_02721_),
    .X(_02722_));
 sg13g2_nand4_1 _09746_ (.B(_02719_),
    .C(_02720_),
    .A(_02718_),
    .Y(_02723_),
    .D(_02721_));
 sg13g2_nor2_1 _09747_ (.A(_02659_),
    .B(_02723_),
    .Y(_02724_));
 sg13g2_o21ai_1 _09748_ (.B1(net1493),
    .Y(_02725_),
    .A1(_02668_),
    .A2(_02722_));
 sg13g2_a21oi_1 _09749_ (.A1(_02669_),
    .A2(_02723_),
    .Y(_02726_),
    .B1(_02659_));
 sg13g2_nand2_1 _09750_ (.Y(_02727_),
    .A(_02668_),
    .B(_02722_));
 sg13g2_nor3_1 _09751_ (.A(_02659_),
    .B(_02669_),
    .C(_02723_),
    .Y(_02728_));
 sg13g2_nor3_1 _09752_ (.A(_00631_),
    .B(_02725_),
    .C(_02728_),
    .Y(_02729_));
 sg13g2_a21oi_1 _09753_ (.A1(_02726_),
    .A2(_02727_),
    .Y(_02730_),
    .B1(\vgadonut.donut.donuthit.cordicxz.xin[4] ));
 sg13g2_a21oi_1 _09754_ (.A1(\vgadonut.donut.donuthit.cordicxz.xin[3] ),
    .A2(_02710_),
    .Y(_02731_),
    .B1(_02711_));
 sg13g2_nor3_1 _09755_ (.A(_02729_),
    .B(_02730_),
    .C(_02731_),
    .Y(_02732_));
 sg13g2_o21ai_1 _09756_ (.B1(_02731_),
    .Y(_02733_),
    .A1(_02729_),
    .A2(_02730_));
 sg13g2_nand2b_1 _09757_ (.Y(_02734_),
    .B(_02733_),
    .A_N(_02732_));
 sg13g2_a21oi_1 _09758_ (.A1(_02703_),
    .A2(_02713_),
    .Y(_02735_),
    .B1(_02676_));
 sg13g2_a21o_1 _09759_ (.A2(_02735_),
    .A1(_02679_),
    .B1(_02714_),
    .X(_02736_));
 sg13g2_a21oi_2 _09760_ (.B1(_02714_),
    .Y(_02737_),
    .A2(_02735_),
    .A1(_02679_));
 sg13g2_xnor2_1 _09761_ (.Y(_02738_),
    .A(_02734_),
    .B(_02736_));
 sg13g2_nor2_1 _09762_ (.A(net1948),
    .B(net1944),
    .Y(_02739_));
 sg13g2_xnor2_1 _09763_ (.Y(_02740_),
    .A(net1948),
    .B(net1944));
 sg13g2_nor3_1 _09764_ (.A(net1949),
    .B(net1946),
    .C(_02740_),
    .Y(_02741_));
 sg13g2_o21ai_1 _09765_ (.B1(_02740_),
    .Y(_02742_),
    .A1(net1949),
    .A2(net1946));
 sg13g2_nand2b_1 _09766_ (.Y(_02743_),
    .B(_02742_),
    .A_N(_02741_));
 sg13g2_a21o_1 _09767_ (.A2(_02693_),
    .A1(_02682_),
    .B1(_02695_),
    .X(_02744_));
 sg13g2_nand2b_1 _09768_ (.Y(_02745_),
    .B(_02744_),
    .A_N(_02743_));
 sg13g2_xor2_1 _09769_ (.B(_02744_),
    .A(_02743_),
    .X(_02746_));
 sg13g2_inv_1 _09770_ (.Y(_02747_),
    .A(_02746_));
 sg13g2_xor2_1 _09771_ (.B(_02746_),
    .A(\vgadonut.donut.donuthit.rzin[9] ),
    .X(_02748_));
 sg13g2_a21o_1 _09772_ (.A2(_02700_),
    .A1(_02698_),
    .B1(_02748_),
    .X(_02749_));
 sg13g2_inv_1 _09773_ (.Y(_02750_),
    .A(_02749_));
 sg13g2_nand3_1 _09774_ (.B(_02700_),
    .C(_02748_),
    .A(_02698_),
    .Y(_02751_));
 sg13g2_nand3_1 _09775_ (.B(_02749_),
    .C(_02751_),
    .A(net1689),
    .Y(_02752_));
 sg13g2_o21ai_1 _09776_ (.B1(_02752_),
    .Y(_00088_),
    .A1(net1687),
    .A2(_02738_));
 sg13g2_a21oi_1 _09777_ (.A1(_02733_),
    .A2(_02737_),
    .Y(_02753_),
    .B1(_02732_));
 sg13g2_nor2_1 _09778_ (.A(_02725_),
    .B(_02729_),
    .Y(_02754_));
 sg13g2_o21ai_1 _09779_ (.B1(_02726_),
    .Y(_02755_),
    .A1(_00631_),
    .A2(_02728_));
 sg13g2_nand2_1 _09780_ (.Y(_02756_),
    .A(net1501),
    .B(_02596_));
 sg13g2_nand2_1 _09781_ (.Y(_02757_),
    .A(net1506),
    .B(_02574_));
 sg13g2_a22oi_1 _09782_ (.Y(_02758_),
    .B1(_02586_),
    .B2(net1528),
    .A2(_02575_),
    .A1(net1503));
 sg13g2_and4_1 _09783_ (.A(_02718_),
    .B(_02756_),
    .C(_02757_),
    .D(_02758_),
    .X(_02759_));
 sg13g2_and2_1 _09784_ (.A(_02660_),
    .B(_02759_),
    .X(_02760_));
 sg13g2_o21ai_1 _09785_ (.B1(_02660_),
    .Y(_02761_),
    .A1(_02708_),
    .A2(_02759_));
 sg13g2_nand3_1 _09786_ (.B(_02708_),
    .C(_02759_),
    .A(_02660_),
    .Y(_02762_));
 sg13g2_nor2b_1 _09787_ (.A(_02761_),
    .B_N(_02762_),
    .Y(_02763_));
 sg13g2_xor2_1 _09788_ (.B(_02763_),
    .A(_00149_),
    .X(_02764_));
 sg13g2_xnor2_1 _09789_ (.Y(_02765_),
    .A(_00149_),
    .B(_02763_));
 sg13g2_xnor2_1 _09790_ (.Y(_02766_),
    .A(_02754_),
    .B(_02764_));
 sg13g2_a21oi_1 _09791_ (.A1(_02753_),
    .A2(_02766_),
    .Y(_02767_),
    .B1(net1687));
 sg13g2_o21ai_1 _09792_ (.B1(_02767_),
    .Y(_02768_),
    .A1(_02753_),
    .A2(_02766_));
 sg13g2_nand2_1 _09793_ (.Y(_02769_),
    .A(net1942),
    .B(_02741_));
 sg13g2_xor2_1 _09794_ (.B(net1942),
    .A(net1946),
    .X(_02770_));
 sg13g2_xnor2_1 _09795_ (.Y(_02771_),
    .A(_02739_),
    .B(_02770_));
 sg13g2_xor2_1 _09796_ (.B(_02771_),
    .A(_02745_),
    .X(_02772_));
 sg13g2_o21ai_1 _09797_ (.B1(_02769_),
    .Y(_02773_),
    .A1(_02741_),
    .A2(_02772_));
 sg13g2_xnor2_1 _09798_ (.Y(_02774_),
    .A(_06876_),
    .B(_02773_));
 sg13g2_a21oi_1 _09799_ (.A1(\vgadonut.donut.donuthit.rzin[9] ),
    .A2(_02747_),
    .Y(_02775_),
    .B1(_02750_));
 sg13g2_or2_1 _09800_ (.X(_02776_),
    .B(_02775_),
    .A(_02774_));
 sg13g2_a21oi_1 _09801_ (.A1(_02774_),
    .A2(_02775_),
    .Y(_02777_),
    .B1(net1673));
 sg13g2_nand2_1 _09802_ (.Y(_02778_),
    .A(_02776_),
    .B(_02777_));
 sg13g2_nand2_1 _09803_ (.Y(_00089_),
    .A(_02768_),
    .B(_02778_));
 sg13g2_o21ai_1 _09804_ (.B1(_02596_),
    .Y(_02779_),
    .A1(net1506),
    .A2(net1501));
 sg13g2_nand2_1 _09805_ (.Y(_02780_),
    .A(_02718_),
    .B(_02779_));
 sg13g2_a22oi_1 _09806_ (.Y(_02781_),
    .B1(_02575_),
    .B2(net1528),
    .A2(_02574_),
    .A1(net1503));
 sg13g2_and4_2 _09807_ (.A(net1493),
    .B(_02718_),
    .C(_02779_),
    .D(_02781_),
    .X(_02782_));
 sg13g2_nor2_1 _09808_ (.A(_02724_),
    .B(_02782_),
    .Y(_02783_));
 sg13g2_nand2_1 _09809_ (.Y(_02784_),
    .A(_02724_),
    .B(_02782_));
 sg13g2_xor2_1 _09810_ (.B(_02782_),
    .A(_02724_),
    .X(_02785_));
 sg13g2_xnor2_1 _09811_ (.Y(_02786_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[6] ),
    .B(_02785_));
 sg13g2_o21ai_1 _09812_ (.B1(_02762_),
    .Y(_02787_),
    .A1(\vgadonut.donut.donuthit.cordicxz.xin[5] ),
    .A2(_02761_));
 sg13g2_nor2_1 _09813_ (.A(_02786_),
    .B(_02787_),
    .Y(_02788_));
 sg13g2_or2_1 _09814_ (.X(_02789_),
    .B(_02787_),
    .A(_02786_));
 sg13g2_xnor2_1 _09815_ (.Y(_02790_),
    .A(_02787_),
    .B(_02786_));
 sg13g2_or3_1 _09816_ (.A(_02734_),
    .B(_02736_),
    .C(_02766_),
    .X(_02791_));
 sg13g2_o21ai_1 _09817_ (.B1(_02732_),
    .Y(_02792_),
    .A1(_02755_),
    .A2(_02765_));
 sg13g2_o21ai_1 _09818_ (.B1(_02792_),
    .Y(_02793_),
    .A1(_02754_),
    .A2(_02764_));
 sg13g2_nor2b_1 _09819_ (.A(_02793_),
    .B_N(_02791_),
    .Y(_02794_));
 sg13g2_nor2_1 _09820_ (.A(_02790_),
    .B(_02794_),
    .Y(_02795_));
 sg13g2_a21o_1 _09821_ (.A2(_02794_),
    .A1(_02790_),
    .B1(net1687),
    .X(_02796_));
 sg13g2_o21ai_1 _09822_ (.B1(_02776_),
    .Y(_02797_),
    .A1(_06876_),
    .A2(_02773_));
 sg13g2_xnor2_1 _09823_ (.Y(_02798_),
    .A(net1944),
    .B(net1941));
 sg13g2_nor3_1 _09824_ (.A(net1947),
    .B(net1942),
    .C(_02798_),
    .Y(_02799_));
 sg13g2_o21ai_1 _09825_ (.B1(_02798_),
    .Y(_02800_),
    .A1(net1947),
    .A2(net1942));
 sg13g2_nand2b_1 _09826_ (.Y(_02801_),
    .B(_02800_),
    .A_N(_02799_));
 sg13g2_o21ai_1 _09827_ (.B1(_02769_),
    .Y(_02802_),
    .A1(_02745_),
    .A2(_02771_));
 sg13g2_a21oi_1 _09828_ (.A1(_02739_),
    .A2(_02770_),
    .Y(_02803_),
    .B1(_02802_));
 sg13g2_or2_1 _09829_ (.X(_02804_),
    .B(_02803_),
    .A(_02801_));
 sg13g2_xor2_1 _09830_ (.B(_02803_),
    .A(_02801_),
    .X(_02805_));
 sg13g2_nand2_1 _09831_ (.Y(_02806_),
    .A(\vgadonut.donut.donuthit.rzin[11] ),
    .B(_02805_));
 sg13g2_xnor2_1 _09832_ (.Y(_02807_),
    .A(\vgadonut.donut.donuthit.rzin[11] ),
    .B(_02805_));
 sg13g2_nand2b_1 _09833_ (.Y(_02808_),
    .B(_02797_),
    .A_N(_02807_));
 sg13g2_nand2b_1 _09834_ (.Y(_02809_),
    .B(_02807_),
    .A_N(_02797_));
 sg13g2_nand3_1 _09835_ (.B(_02808_),
    .C(_02809_),
    .A(net1687),
    .Y(_02810_));
 sg13g2_o21ai_1 _09836_ (.B1(_02810_),
    .Y(_00090_),
    .A1(_02795_),
    .A2(_02796_));
 sg13g2_a21o_1 _09837_ (.A2(_02784_),
    .A1(\vgadonut.donut.donuthit.cordicxz.xin[6] ),
    .B1(_02783_),
    .X(_02811_));
 sg13g2_nand2_1 _09838_ (.Y(_02812_),
    .A(net1528),
    .B(_02574_));
 sg13g2_o21ai_1 _09839_ (.B1(_02812_),
    .Y(_02813_),
    .A1(_01863_),
    .A2(_02595_));
 sg13g2_nor3_2 _09840_ (.A(_02659_),
    .B(_02780_),
    .C(_02813_),
    .Y(_02814_));
 sg13g2_and2_1 _09841_ (.A(_02760_),
    .B(_02814_),
    .X(_02815_));
 sg13g2_nor2_1 _09842_ (.A(_02760_),
    .B(_02814_),
    .Y(_02816_));
 sg13g2_xnor2_1 _09843_ (.Y(_02817_),
    .A(_02760_),
    .B(_02814_));
 sg13g2_xor2_1 _09844_ (.B(_02817_),
    .A(_00147_),
    .X(_02818_));
 sg13g2_nor2_1 _09845_ (.A(_02811_),
    .B(_02818_),
    .Y(_02819_));
 sg13g2_nand2_1 _09846_ (.Y(_02820_),
    .A(_02811_),
    .B(_02818_));
 sg13g2_xnor2_1 _09847_ (.Y(_02821_),
    .A(_02811_),
    .B(_02818_));
 sg13g2_nor2_1 _09848_ (.A(_02788_),
    .B(_02795_),
    .Y(_02822_));
 sg13g2_a21oi_1 _09849_ (.A1(_02821_),
    .A2(_02822_),
    .Y(_02823_),
    .B1(net1687));
 sg13g2_o21ai_1 _09850_ (.B1(_02823_),
    .Y(_02824_),
    .A1(_02821_),
    .A2(_02822_));
 sg13g2_nand2_1 _09851_ (.Y(_02825_),
    .A(net1939),
    .B(_02799_));
 sg13g2_xnor2_1 _09852_ (.Y(_02826_),
    .A(net1943),
    .B(net1938));
 sg13g2_nor3_1 _09853_ (.A(net1945),
    .B(net1940),
    .C(_02826_),
    .Y(_02827_));
 sg13g2_o21ai_1 _09854_ (.B1(_02826_),
    .Y(_02828_),
    .A1(net1944),
    .A2(net1940));
 sg13g2_nand2b_1 _09855_ (.Y(_02829_),
    .B(_02828_),
    .A_N(_02827_));
 sg13g2_xnor2_1 _09856_ (.Y(_02830_),
    .A(_02804_),
    .B(_02829_));
 sg13g2_nand2b_1 _09857_ (.Y(_02831_),
    .B(_02830_),
    .A_N(_02799_));
 sg13g2_nand2_1 _09858_ (.Y(_02832_),
    .A(_02825_),
    .B(_02831_));
 sg13g2_nand3_1 _09859_ (.B(_02825_),
    .C(_02831_),
    .A(net2356),
    .Y(_02833_));
 sg13g2_xnor2_1 _09860_ (.Y(_02834_),
    .A(_06878_),
    .B(_02832_));
 sg13g2_a21o_1 _09861_ (.A2(_02808_),
    .A1(_02806_),
    .B1(_02834_),
    .X(_02835_));
 sg13g2_nand3_1 _09862_ (.B(_02808_),
    .C(_02834_),
    .A(_02806_),
    .Y(_02836_));
 sg13g2_nand3_1 _09863_ (.B(_02835_),
    .C(_02836_),
    .A(net1687),
    .Y(_02837_));
 sg13g2_nand2_1 _09864_ (.Y(_00091_),
    .A(_02824_),
    .B(_02837_));
 sg13g2_nor2_1 _09865_ (.A(net1940),
    .B(net1937),
    .Y(_02838_));
 sg13g2_xnor2_1 _09866_ (.Y(_02839_),
    .A(net1940),
    .B(net1936));
 sg13g2_nor3_2 _09867_ (.A(net1943),
    .B(net1939),
    .C(_02839_),
    .Y(_02840_));
 sg13g2_o21ai_1 _09868_ (.B1(_02839_),
    .Y(_02841_),
    .A1(net1943),
    .A2(net1939));
 sg13g2_nand2b_1 _09869_ (.Y(_02842_),
    .B(_02841_),
    .A_N(_02840_));
 sg13g2_o21ai_1 _09870_ (.B1(_02825_),
    .Y(_02843_),
    .A1(_02804_),
    .A2(_02829_));
 sg13g2_nor2_1 _09871_ (.A(_02827_),
    .B(_02843_),
    .Y(_02844_));
 sg13g2_nor2_1 _09872_ (.A(_02842_),
    .B(_02844_),
    .Y(_02845_));
 sg13g2_xor2_1 _09873_ (.B(_02844_),
    .A(_02842_),
    .X(_02846_));
 sg13g2_nand2_1 _09874_ (.Y(_02847_),
    .A(\vgadonut.donut.donuthit.rzin[13] ),
    .B(_02846_));
 sg13g2_xnor2_1 _09875_ (.Y(_02848_),
    .A(\vgadonut.donut.donuthit.rzin[13] ),
    .B(_02846_));
 sg13g2_nand3_1 _09876_ (.B(_02835_),
    .C(_02848_),
    .A(_02833_),
    .Y(_02849_));
 sg13g2_a21o_1 _09877_ (.A2(_02835_),
    .A1(_02833_),
    .B1(_02848_),
    .X(_02850_));
 sg13g2_nand3_1 _09878_ (.B(_02849_),
    .C(_02850_),
    .A(net1686),
    .Y(_02851_));
 sg13g2_nor2_1 _09879_ (.A(_02790_),
    .B(_02821_),
    .Y(_02852_));
 sg13g2_nor4_2 _09880_ (.A(_02734_),
    .B(_02766_),
    .C(_02790_),
    .Y(_02853_),
    .D(_02821_));
 sg13g2_nand2_1 _09881_ (.Y(_02854_),
    .A(_02737_),
    .B(_02853_));
 sg13g2_nand2_1 _09882_ (.Y(_02855_),
    .A(_02793_),
    .B(_02852_));
 sg13g2_o21ai_1 _09883_ (.B1(_02820_),
    .Y(_02856_),
    .A1(_02789_),
    .A2(_02819_));
 sg13g2_a221oi_1 _09884_ (.B2(_02737_),
    .C1(_02856_),
    .B1(_02853_),
    .A1(_02793_),
    .Y(_02857_),
    .A2(_02852_));
 sg13g2_nand3b_1 _09885_ (.B(_02855_),
    .C(_02854_),
    .Y(_02858_),
    .A_N(_02856_));
 sg13g2_nor2_1 _09886_ (.A(net1517),
    .B(_02595_),
    .Y(_02859_));
 sg13g2_nor3_2 _09887_ (.A(_02659_),
    .B(_02780_),
    .C(_02859_),
    .Y(_02860_));
 sg13g2_nor2_1 _09888_ (.A(_02782_),
    .B(net1492),
    .Y(_02861_));
 sg13g2_xnor2_1 _09889_ (.Y(_02862_),
    .A(_02782_),
    .B(net1492));
 sg13g2_inv_1 _09890_ (.Y(_02863_),
    .A(_02862_));
 sg13g2_xor2_1 _09891_ (.B(_02862_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[8] ),
    .X(_02864_));
 sg13g2_nor2_1 _09892_ (.A(\vgadonut.donut.donuthit.cordicxz.xin[7] ),
    .B(_02816_),
    .Y(_02865_));
 sg13g2_nor2_1 _09893_ (.A(_02815_),
    .B(_02865_),
    .Y(_02866_));
 sg13g2_nor3_1 _09894_ (.A(_02815_),
    .B(_02864_),
    .C(_02865_),
    .Y(_02867_));
 sg13g2_xnor2_1 _09895_ (.Y(_02868_),
    .A(_02864_),
    .B(_02866_));
 sg13g2_nor2b_2 _09896_ (.A(_02857_),
    .B_N(_02868_),
    .Y(_02869_));
 sg13g2_o21ai_1 _09897_ (.B1(net1673),
    .Y(_02870_),
    .A1(_02858_),
    .A2(_02868_));
 sg13g2_o21ai_1 _09898_ (.B1(_02851_),
    .Y(_00092_),
    .A1(_02869_),
    .A2(_02870_));
 sg13g2_nor2_1 _09899_ (.A(_02867_),
    .B(_02869_),
    .Y(_02871_));
 sg13g2_a21oi_1 _09900_ (.A1(\vgadonut.donut.donuthit.cordicxz.xin[8] ),
    .A2(_02863_),
    .Y(_02872_),
    .B1(_02861_));
 sg13g2_xnor2_1 _09901_ (.Y(_02873_),
    .A(_02814_),
    .B(net1492));
 sg13g2_xnor2_1 _09902_ (.Y(_02874_),
    .A(_00145_),
    .B(_02873_));
 sg13g2_nand2_1 _09903_ (.Y(_02875_),
    .A(_02872_),
    .B(_02874_));
 sg13g2_inv_1 _09904_ (.Y(_02876_),
    .A(_02875_));
 sg13g2_nor2_1 _09905_ (.A(_02872_),
    .B(_02874_),
    .Y(_02877_));
 sg13g2_or2_1 _09906_ (.X(_02878_),
    .B(_02877_),
    .A(_02876_));
 sg13g2_a21oi_1 _09907_ (.A1(_02871_),
    .A2(_02878_),
    .Y(_02879_),
    .B1(net1689));
 sg13g2_o21ai_1 _09908_ (.B1(_02879_),
    .Y(_02880_),
    .A1(_02871_),
    .A2(_02878_));
 sg13g2_xor2_1 _09909_ (.B(\vgadonut.donut.cAcB[15] ),
    .A(net1938),
    .X(_02881_));
 sg13g2_xnor2_1 _09910_ (.Y(_02882_),
    .A(_02838_),
    .B(_02881_));
 sg13g2_nor3_1 _09911_ (.A(_02842_),
    .B(_02844_),
    .C(_02882_),
    .Y(_02883_));
 sg13g2_xor2_1 _09912_ (.B(_02882_),
    .A(_02845_),
    .X(_02884_));
 sg13g2_mux2_1 _09913_ (.A0(_02884_),
    .A1(\vgadonut.donut.cAcB[15] ),
    .S(_02840_),
    .X(_02885_));
 sg13g2_nor2_1 _09914_ (.A(_06881_),
    .B(_02885_),
    .Y(_02886_));
 sg13g2_xnor2_1 _09915_ (.Y(_02887_),
    .A(_06881_),
    .B(_02885_));
 sg13g2_a21o_1 _09916_ (.A2(_02850_),
    .A1(_02847_),
    .B1(_02887_),
    .X(_02888_));
 sg13g2_nand3_1 _09917_ (.B(_02850_),
    .C(_02887_),
    .A(_02847_),
    .Y(_02889_));
 sg13g2_nand3_1 _09918_ (.B(_02888_),
    .C(_02889_),
    .A(net1686),
    .Y(_02890_));
 sg13g2_nand2_1 _09919_ (.Y(_00093_),
    .A(_02880_),
    .B(_02890_));
 sg13g2_or2_1 _09920_ (.X(_02891_),
    .B(_02877_),
    .A(_02867_));
 sg13g2_o21ai_1 _09921_ (.B1(_02875_),
    .Y(_02892_),
    .A1(_02891_),
    .A2(_02869_));
 sg13g2_a21o_1 _09922_ (.A2(net1492),
    .A1(_02814_),
    .B1(_00628_),
    .X(_02893_));
 sg13g2_o21ai_1 _09923_ (.B1(_02893_),
    .Y(_02894_),
    .A1(_02814_),
    .A2(net1492));
 sg13g2_xnor2_1 _09924_ (.Y(_02895_),
    .A(\vgadonut.donut.donuthit.cordicxz.xin[10] ),
    .B(_02894_));
 sg13g2_a21oi_1 _09925_ (.A1(_02892_),
    .A2(_02895_),
    .Y(_02896_),
    .B1(net1700));
 sg13g2_o21ai_1 _09926_ (.B1(_02896_),
    .Y(_02897_),
    .A1(_02892_),
    .A2(_02895_));
 sg13g2_nor2b_1 _09927_ (.A(_02886_),
    .B_N(_02888_),
    .Y(_02898_));
 sg13g2_a221oi_1 _09928_ (.B2(_02838_),
    .C1(_02883_),
    .B1(_02881_),
    .A1(net1935),
    .Y(_02899_),
    .A2(_02840_));
 sg13g2_nor2b_1 _09929_ (.A(net1935),
    .B_N(net1938),
    .Y(_02900_));
 sg13g2_xnor2_1 _09930_ (.Y(_02901_),
    .A(net1936),
    .B(_02900_));
 sg13g2_nand2b_1 _09931_ (.Y(_02902_),
    .B(_02901_),
    .A_N(_02899_));
 sg13g2_xnor2_1 _09932_ (.Y(_02903_),
    .A(_02899_),
    .B(_02901_));
 sg13g2_xnor2_1 _09933_ (.Y(_02904_),
    .A(\vgadonut.donut.donuthit.rzin[15] ),
    .B(_02903_));
 sg13g2_nor2_1 _09934_ (.A(_02898_),
    .B(_02904_),
    .Y(_02905_));
 sg13g2_a21o_1 _09935_ (.A2(_02904_),
    .A1(_02898_),
    .B1(net1673),
    .X(_02906_));
 sg13g2_o21ai_1 _09936_ (.B1(_02897_),
    .Y(_00079_),
    .A1(_02905_),
    .A2(_02906_));
 sg13g2_nand2_1 _09937_ (.Y(_02907_),
    .A(_00627_),
    .B(_02894_));
 sg13g2_o21ai_1 _09938_ (.B1(_02907_),
    .Y(_02908_),
    .A1(_02892_),
    .A2(_02895_));
 sg13g2_nor2_1 _09939_ (.A(_00626_),
    .B(_02860_),
    .Y(_02909_));
 sg13g2_xnor2_1 _09940_ (.Y(_02910_),
    .A(_00626_),
    .B(_02860_));
 sg13g2_and2_2 _09941_ (.A(_02908_),
    .B(_02910_),
    .X(_02911_));
 sg13g2_o21ai_1 _09942_ (.B1(net1673),
    .Y(_02912_),
    .A1(_02908_),
    .A2(_02910_));
 sg13g2_a21o_1 _09943_ (.A2(_02903_),
    .A1(_00639_),
    .B1(_02905_),
    .X(_02913_));
 sg13g2_nor3_1 _09944_ (.A(net1936),
    .B(net1935),
    .C(_02902_),
    .Y(_02914_));
 sg13g2_a21o_1 _09945_ (.A2(net1936),
    .A1(net1938),
    .B1(net1935),
    .X(_02915_));
 sg13g2_a21oi_2 _09946_ (.B1(_02914_),
    .Y(_02916_),
    .A2(_02915_),
    .A1(_02902_));
 sg13g2_xnor2_1 _09947_ (.Y(_02917_),
    .A(_06882_),
    .B(_02916_));
 sg13g2_nand2b_1 _09948_ (.Y(_02918_),
    .B(_02917_),
    .A_N(_02913_));
 sg13g2_xor2_1 _09949_ (.B(_02917_),
    .A(_02913_),
    .X(_02919_));
 sg13g2_nand2_1 _09950_ (.Y(_02920_),
    .A(net1688),
    .B(_02919_));
 sg13g2_o21ai_1 _09951_ (.B1(_02920_),
    .Y(_00080_),
    .A1(_02911_),
    .A2(_02912_));
 sg13g2_nand2_1 _09952_ (.Y(_02921_),
    .A(_00639_),
    .B(_02916_));
 sg13g2_o21ai_1 _09953_ (.B1(net1686),
    .Y(_02922_),
    .A1(\vgadonut.donut.donuthit.rzin[15] ),
    .A2(_02921_));
 sg13g2_a21o_2 _09954_ (.A2(_02921_),
    .A1(_02918_),
    .B1(_02922_),
    .X(_02923_));
 sg13g2_nand2_1 _09955_ (.Y(_02924_),
    .A(_00143_),
    .B(_00155_));
 sg13g2_xnor2_1 _09956_ (.Y(_02925_),
    .A(_00155_),
    .B(_02909_));
 sg13g2_nand2_1 _09957_ (.Y(_02926_),
    .A(_02911_),
    .B(_02925_));
 sg13g2_xnor2_1 _09958_ (.Y(_02927_),
    .A(_02911_),
    .B(_02925_));
 sg13g2_o21ai_1 _09959_ (.B1(_02923_),
    .Y(_00081_),
    .A1(net1688),
    .A2(_02927_));
 sg13g2_nand2b_1 _09960_ (.Y(_02928_),
    .B(_00155_),
    .A_N(net1492));
 sg13g2_o21ai_1 _09961_ (.B1(_02926_),
    .Y(_02929_),
    .A1(net2354),
    .A2(_02928_));
 sg13g2_nor2_1 _09962_ (.A(_00636_),
    .B(net1492),
    .Y(_02930_));
 sg13g2_xnor2_1 _09963_ (.Y(_02931_),
    .A(_00636_),
    .B(_02928_));
 sg13g2_xnor2_1 _09964_ (.Y(_02932_),
    .A(_02929_),
    .B(_02931_));
 sg13g2_o21ai_1 _09965_ (.B1(_02923_),
    .Y(_00082_),
    .A1(net1688),
    .A2(_02932_));
 sg13g2_and2_1 _09966_ (.A(_02925_),
    .B(_02931_),
    .X(_02933_));
 sg13g2_a22oi_1 _09967_ (.Y(_02934_),
    .B1(_02933_),
    .B2(_02911_),
    .A2(_02930_),
    .A1(_02924_));
 sg13g2_nor2b_1 _09968_ (.A(net1492),
    .B_N(_00158_),
    .Y(_02935_));
 sg13g2_nand2_1 _09969_ (.Y(_02936_),
    .A(_00636_),
    .B(_02935_));
 sg13g2_xnor2_1 _09970_ (.Y(_02937_),
    .A(_00158_),
    .B(_02930_));
 sg13g2_inv_1 _09971_ (.Y(_02938_),
    .A(_02937_));
 sg13g2_xnor2_1 _09972_ (.Y(_02939_),
    .A(_02934_),
    .B(_02938_));
 sg13g2_o21ai_1 _09973_ (.B1(_02923_),
    .Y(_00083_),
    .A1(net1688),
    .A2(_02939_));
 sg13g2_o21ai_1 _09974_ (.B1(_02936_),
    .Y(_02940_),
    .A1(_02934_),
    .A2(_02938_));
 sg13g2_xnor2_1 _09975_ (.Y(_02941_),
    .A(net2286),
    .B(_02935_));
 sg13g2_xnor2_1 _09976_ (.Y(_02942_),
    .A(_02940_),
    .B(_02941_));
 sg13g2_o21ai_1 _09977_ (.B1(_02923_),
    .Y(_00084_),
    .A1(net1688),
    .A2(_02942_));
 sg13g2_nand2b_2 _09978_ (.Y(_02943_),
    .B(net1801),
    .A_N(\vgadonut.donut.h_count[3] ));
 sg13g2_nand3_1 _09979_ (.B(\vgadonut.donut.h_count[7] ),
    .C(\vgadonut.donut.h_count[6] ),
    .A(\vgadonut.donut.h_count[5] ),
    .Y(_02944_));
 sg13g2_nor2b_1 _09980_ (.A(net2062),
    .B_N(\vgadonut.donut.h_count[10] ),
    .Y(_02945_));
 sg13g2_and2_2 _09981_ (.A(\vgadonut.donut.h_count[8] ),
    .B(_02945_),
    .X(_02946_));
 sg13g2_nor2_1 _09982_ (.A(net1802),
    .B(net1803),
    .Y(_02947_));
 sg13g2_nand3_1 _09983_ (.B(_02946_),
    .C(_02947_),
    .A(net1800),
    .Y(_02948_));
 sg13g2_nor3_1 _09984_ (.A(_02943_),
    .B(_02944_),
    .C(_02948_),
    .Y(_02949_));
 sg13g2_inv_1 _09985_ (.Y(_02950_),
    .A(net1740));
 sg13g2_nor2_1 _09986_ (.A(net1803),
    .B(net1741),
    .Y(_00014_));
 sg13g2_nand2b_2 _09987_ (.Y(_02951_),
    .B(net1802),
    .A_N(net1803));
 sg13g2_xor2_1 _09988_ (.B(\vgadonut.donut.h_count[0] ),
    .A(net2002),
    .X(_00016_));
 sg13g2_nand2_1 _09989_ (.Y(_02952_),
    .A(net1802),
    .B(net1803));
 sg13g2_nor2_1 _09990_ (.A(net1991),
    .B(_02952_),
    .Y(_02953_));
 sg13g2_and2_1 _09991_ (.A(net1991),
    .B(_02952_),
    .X(_02954_));
 sg13g2_nor3_1 _09992_ (.A(net1741),
    .B(_02953_),
    .C(_02954_),
    .Y(_00017_));
 sg13g2_xor2_1 _09993_ (.B(_02953_),
    .A(net2025),
    .X(_02955_));
 sg13g2_nor2_1 _09994_ (.A(net1741),
    .B(_02955_),
    .Y(_00018_));
 sg13g2_and3_1 _09995_ (.X(_02956_),
    .A(net1802),
    .B(net1803),
    .C(_00649_));
 sg13g2_nor2_1 _09996_ (.A(net2108),
    .B(_02956_),
    .Y(_02957_));
 sg13g2_and2_1 _09997_ (.A(net1800),
    .B(_02956_),
    .X(_02958_));
 sg13g2_nor3_1 _09998_ (.A(net1740),
    .B(_02957_),
    .C(_02958_),
    .Y(_00019_));
 sg13g2_nor2_1 _09999_ (.A(net2181),
    .B(_02958_),
    .Y(_02959_));
 sg13g2_and2_1 _10000_ (.A(net2181),
    .B(_02958_),
    .X(_02960_));
 sg13g2_nor3_1 _10001_ (.A(net1740),
    .B(_02959_),
    .C(_02960_),
    .Y(_00020_));
 sg13g2_nor2_1 _10002_ (.A(net2142),
    .B(_02960_),
    .Y(_02961_));
 sg13g2_and2_1 _10003_ (.A(net2142),
    .B(_02960_),
    .X(_02962_));
 sg13g2_nor3_1 _10004_ (.A(net1740),
    .B(net2143),
    .C(_02962_),
    .Y(_00021_));
 sg13g2_nor2b_1 _10005_ (.A(_00651_),
    .B_N(_02960_),
    .Y(_02963_));
 sg13g2_o21ai_1 _10006_ (.B1(_02950_),
    .Y(_02964_),
    .A1(net2076),
    .A2(_02962_));
 sg13g2_nor2_1 _10007_ (.A(_02963_),
    .B(_02964_),
    .Y(_00022_));
 sg13g2_nor2_1 _10008_ (.A(net2161),
    .B(_02963_),
    .Y(_02965_));
 sg13g2_and2_1 _10009_ (.A(net2161),
    .B(_02963_),
    .X(_02966_));
 sg13g2_nor3_1 _10010_ (.A(net1740),
    .B(_02965_),
    .C(_02966_),
    .Y(_00023_));
 sg13g2_nand2_1 _10011_ (.Y(_02967_),
    .A(\vgadonut.donut.h_count[9] ),
    .B(_02966_));
 sg13g2_xor2_1 _10012_ (.B(_02966_),
    .A(net2062),
    .X(_00024_));
 sg13g2_o21ai_1 _10013_ (.B1(_02950_),
    .Y(_02968_),
    .A1(net1445),
    .A2(_02967_));
 sg13g2_a21oi_1 _10014_ (.A1(net1445),
    .A2(_02967_),
    .Y(_00015_),
    .B1(_02968_));
 sg13g2_nand2_1 _10015_ (.Y(_02969_),
    .A(\vgadonut.donut.v_count[7] ),
    .B(\vgadonut.donut.v_count[6] ));
 sg13g2_nor2_1 _10016_ (.A(net2146),
    .B(_02969_),
    .Y(_02970_));
 sg13g2_and2_1 _10017_ (.A(\vgadonut.bayer_j[1] ),
    .B(net1915),
    .X(_02971_));
 sg13g2_o21ai_1 _10018_ (.B1(_02970_),
    .Y(_02972_),
    .A1(net2218),
    .A2(_02971_));
 sg13g2_o21ai_1 _10019_ (.B1(_02972_),
    .Y(_02973_),
    .A1(net1915),
    .A2(net2218));
 sg13g2_nand2_1 _10020_ (.Y(_02974_),
    .A(\vgadonut.donut.v_count[3] ),
    .B(net1914));
 sg13g2_nand3_1 _10021_ (.B(net1914),
    .C(_02970_),
    .A(net1913),
    .Y(_02975_));
 sg13g2_nor2b_1 _10022_ (.A(\vgadonut.donut.v_count[9] ),
    .B_N(\vgadonut.donut.v_count[8] ),
    .Y(_02976_));
 sg13g2_nand3_1 _10023_ (.B(net2026),
    .C(\vgadonut.donut.v_count[6] ),
    .A(\vgadonut.donut.v_count[5] ),
    .Y(_02977_));
 sg13g2_nor2_1 _10024_ (.A(\vgadonut.donut.v_count[4] ),
    .B(_02977_),
    .Y(_02978_));
 sg13g2_and4_1 _10025_ (.A(net2190),
    .B(net1913),
    .C(_02976_),
    .D(_02978_),
    .X(_02979_));
 sg13g2_or2_1 _10026_ (.X(_02980_),
    .B(net1915),
    .A(\vgadonut.bayer_j[1] ));
 sg13g2_nand3_1 _10027_ (.B(_02975_),
    .C(_02979_),
    .A(_02973_),
    .Y(_00026_));
 sg13g2_nor3_1 _10028_ (.A(net1801),
    .B(\vgadonut.donut.h_count[3] ),
    .C(net1800),
    .Y(_02981_));
 sg13g2_a21oi_1 _10029_ (.A1(_02952_),
    .A2(_02981_),
    .Y(_02982_),
    .B1(_02944_));
 sg13g2_nor2_1 _10030_ (.A(net1802),
    .B(net1801),
    .Y(_02983_));
 sg13g2_nor2_1 _10031_ (.A(\vgadonut.donut.h_count[5] ),
    .B(\vgadonut.donut.h_count[6] ),
    .Y(_02984_));
 sg13g2_o21ai_1 _10032_ (.B1(_02984_),
    .Y(_02985_),
    .A1(_00648_),
    .A2(_02983_));
 sg13g2_nand3_1 _10033_ (.B(\vgadonut.donut.h_count[8] ),
    .C(_02985_),
    .A(net2076),
    .Y(_02986_));
 sg13g2_o21ai_1 _10034_ (.B1(_02945_),
    .Y(_02987_),
    .A1(\vgadonut.donut.h_count[8] ),
    .A2(_02982_));
 sg13g2_nand2b_1 _10035_ (.Y(_00025_),
    .B(net2077),
    .A_N(_02987_));
 sg13g2_nor2b_1 _10036_ (.A(net1818),
    .B_N(net1922),
    .Y(_02988_));
 sg13g2_nand2b_1 _10037_ (.Y(_02989_),
    .B(net1818),
    .A_N(net1923));
 sg13g2_nand2b_1 _10038_ (.Y(_02990_),
    .B(_02989_),
    .A_N(_02988_));
 sg13g2_nor2b_1 _10039_ (.A(net1924),
    .B_N(net1820),
    .Y(_02991_));
 sg13g2_nand2b_1 _10040_ (.Y(_02992_),
    .B(net1924),
    .A_N(net1820));
 sg13g2_nor2b_1 _10041_ (.A(\vgadonut.donut.cA[10] ),
    .B_N(net1927),
    .Y(_02993_));
 sg13g2_nand2b_1 _10042_ (.Y(_02994_),
    .B(net1821),
    .A_N(net1927));
 sg13g2_nand2b_1 _10043_ (.Y(_02995_),
    .B(_02994_),
    .A_N(_02993_));
 sg13g2_xnor2_1 _10044_ (.Y(_02996_),
    .A(net1931),
    .B(\vgadonut.donut.cA[6] ));
 sg13g2_xor2_1 _10045_ (.B(\vgadonut.donut.cA[5] ),
    .A(net1932),
    .X(_02997_));
 sg13g2_xor2_1 _10046_ (.B(\vgadonut.donut.cA[4] ),
    .A(net1934),
    .X(_02998_));
 sg13g2_nor2b_1 _10047_ (.A(net1825),
    .B_N(\vgadonut.donut.sAcB[2] ),
    .Y(_02999_));
 sg13g2_xnor2_1 _10048_ (.Y(_03000_),
    .A(\vgadonut.donut.sAcB[2] ),
    .B(net1825));
 sg13g2_nor2b_1 _10049_ (.A(\vgadonut.donut.sAcB[1] ),
    .B_N(\vgadonut.donut.cA[1] ),
    .Y(_03001_));
 sg13g2_nand2b_1 _10050_ (.Y(_03002_),
    .B(\vgadonut.donut.sAcB[1] ),
    .A_N(\vgadonut.donut.cA[1] ));
 sg13g2_nor2b_1 _10051_ (.A(\vgadonut.donut.sAcB[0] ),
    .B_N(\vgadonut.donut.cA[0] ),
    .Y(_03003_));
 sg13g2_a21oi_1 _10052_ (.A1(_03002_),
    .A2(_03003_),
    .Y(_03004_),
    .B1(_03001_));
 sg13g2_a21oi_1 _10053_ (.A1(_03000_),
    .A2(_03004_),
    .Y(_03005_),
    .B1(_02999_));
 sg13g2_xnor2_1 _10054_ (.Y(_03006_),
    .A(\vgadonut.donut.sAcB[3] ),
    .B(\vgadonut.donut.cA[3] ));
 sg13g2_nor2b_1 _10055_ (.A(_03005_),
    .B_N(_03006_),
    .Y(_03007_));
 sg13g2_a21oi_1 _10056_ (.A1(\vgadonut.donut.sAcB[3] ),
    .A2(_00603_),
    .Y(_03008_),
    .B1(_03007_));
 sg13g2_nor2_1 _10057_ (.A(_02998_),
    .B(_03008_),
    .Y(_03009_));
 sg13g2_a21oi_1 _10058_ (.A1(net1934),
    .A2(_00602_),
    .Y(_03010_),
    .B1(_03009_));
 sg13g2_nor2_1 _10059_ (.A(_02997_),
    .B(_03010_),
    .Y(_03011_));
 sg13g2_a21oi_1 _10060_ (.A1(net1932),
    .A2(_00601_),
    .Y(_03012_),
    .B1(_03011_));
 sg13g2_nor2b_1 _10061_ (.A(_03012_),
    .B_N(_02996_),
    .Y(_03013_));
 sg13g2_a21oi_1 _10062_ (.A1(net1931),
    .A2(_00600_),
    .Y(_03014_),
    .B1(_03013_));
 sg13g2_xnor2_1 _10063_ (.Y(_03015_),
    .A(net1930),
    .B(net1824));
 sg13g2_nor2b_1 _10064_ (.A(_03014_),
    .B_N(_03015_),
    .Y(_03016_));
 sg13g2_a21oi_2 _10065_ (.B1(_03016_),
    .Y(_03017_),
    .A2(_00604_),
    .A1(net1930));
 sg13g2_xnor2_1 _10066_ (.Y(_03018_),
    .A(net1929),
    .B(net1823));
 sg13g2_nand2b_1 _10067_ (.Y(_03019_),
    .B(_03018_),
    .A_N(_03017_));
 sg13g2_o21ai_1 _10068_ (.B1(_03019_),
    .Y(_03020_),
    .A1(_06910_),
    .A2(net1823));
 sg13g2_a21oi_1 _10069_ (.A1(net1928),
    .A2(_00605_),
    .Y(_03021_),
    .B1(_03020_));
 sg13g2_a21oi_2 _10070_ (.B1(_03021_),
    .Y(_03022_),
    .A2(net1822),
    .A1(_06913_));
 sg13g2_a21oi_2 _10071_ (.B1(_02993_),
    .Y(_03023_),
    .A2(_03022_),
    .A1(_02994_));
 sg13g2_o21ai_1 _10072_ (.B1(_02992_),
    .Y(_03024_),
    .A1(_02991_),
    .A2(_03023_));
 sg13g2_a21oi_1 _10073_ (.A1(_02989_),
    .A2(_03024_),
    .Y(_03025_),
    .B1(_02988_));
 sg13g2_nand2b_1 _10074_ (.Y(_03026_),
    .B(net1920),
    .A_N(net1816));
 sg13g2_nor2b_1 _10075_ (.A(net1920),
    .B_N(net1816),
    .Y(_03027_));
 sg13g2_xnor2_1 _10076_ (.Y(_03028_),
    .A(net1920),
    .B(net1816));
 sg13g2_xnor2_1 _10077_ (.Y(_03029_),
    .A(_03025_),
    .B(_03028_));
 sg13g2_nand2b_1 _10078_ (.Y(_03030_),
    .B(_03029_),
    .A_N(_00127_));
 sg13g2_xnor2_1 _10079_ (.Y(_03031_),
    .A(_00127_),
    .B(_03029_));
 sg13g2_xnor2_1 _10080_ (.Y(_03032_),
    .A(_02990_),
    .B(_03024_));
 sg13g2_nand2_1 _10081_ (.Y(_03033_),
    .A(_00128_),
    .B(_03032_));
 sg13g2_nor2b_1 _10082_ (.A(_02991_),
    .B_N(_02992_),
    .Y(_03034_));
 sg13g2_xnor2_1 _10083_ (.Y(_03035_),
    .A(_03023_),
    .B(_03034_));
 sg13g2_inv_1 _10084_ (.Y(_03036_),
    .A(_03035_));
 sg13g2_nor2_1 _10085_ (.A(net1877),
    .B(_03036_),
    .Y(_03037_));
 sg13g2_xnor2_1 _10086_ (.Y(_03038_),
    .A(_02995_),
    .B(_03022_));
 sg13g2_xnor2_1 _10087_ (.Y(_03039_),
    .A(net1928),
    .B(net1822));
 sg13g2_xnor2_1 _10088_ (.Y(_03040_),
    .A(_03020_),
    .B(_03039_));
 sg13g2_or2_1 _10089_ (.X(_03041_),
    .B(_03040_),
    .A(net1880));
 sg13g2_nor2_1 _10090_ (.A(_00131_),
    .B(_03040_),
    .Y(_03042_));
 sg13g2_xnor2_1 _10091_ (.Y(_03043_),
    .A(_00131_),
    .B(_03040_));
 sg13g2_xnor2_1 _10092_ (.Y(_03044_),
    .A(_03017_),
    .B(_03018_));
 sg13g2_and2_1 _10093_ (.A(_00132_),
    .B(_03044_),
    .X(_03045_));
 sg13g2_xnor2_1 _10094_ (.Y(_03046_),
    .A(_03014_),
    .B(_03015_));
 sg13g2_xnor2_1 _10095_ (.Y(_03047_),
    .A(_02996_),
    .B(_03012_));
 sg13g2_nand2_1 _10096_ (.Y(_03048_),
    .A(_00134_),
    .B(_03047_));
 sg13g2_xor2_1 _10097_ (.B(_03010_),
    .A(_02997_),
    .X(_03049_));
 sg13g2_xnor2_1 _10098_ (.Y(_03050_),
    .A(_00135_),
    .B(_03049_));
 sg13g2_xor2_1 _10099_ (.B(_03008_),
    .A(_02998_),
    .X(_03051_));
 sg13g2_xor2_1 _10100_ (.B(_03006_),
    .A(_03005_),
    .X(_03052_));
 sg13g2_xnor2_1 _10101_ (.Y(_03053_),
    .A(_00569_),
    .B(_03052_));
 sg13g2_xor2_1 _10102_ (.B(_03004_),
    .A(_03000_),
    .X(_03054_));
 sg13g2_nor2_1 _10103_ (.A(_00138_),
    .B(_03054_),
    .Y(_03055_));
 sg13g2_nand2b_1 _10104_ (.Y(_03056_),
    .B(_03053_),
    .A_N(_03055_));
 sg13g2_o21ai_1 _10105_ (.B1(_03056_),
    .Y(_03057_),
    .A1(\vgadonut.donut.donuthit.cordicxy.x2in[1] ),
    .A2(_03052_));
 sg13g2_xnor2_1 _10106_ (.Y(_03058_),
    .A(_00136_),
    .B(_03051_));
 sg13g2_nor2b_1 _10107_ (.A(_03058_),
    .B_N(_03057_),
    .Y(_03059_));
 sg13g2_a21o_1 _10108_ (.A2(_03051_),
    .A1(_00136_),
    .B1(_03059_),
    .X(_03060_));
 sg13g2_nor2b_1 _10109_ (.A(_03050_),
    .B_N(_03060_),
    .Y(_03061_));
 sg13g2_a21oi_1 _10110_ (.A1(_00573_),
    .A2(_03049_),
    .Y(_03062_),
    .B1(_03061_));
 sg13g2_xnor2_1 _10111_ (.Y(_03063_),
    .A(_00134_),
    .B(_03047_));
 sg13g2_or2_1 _10112_ (.X(_03064_),
    .B(_03063_),
    .A(_03062_));
 sg13g2_xnor2_1 _10113_ (.Y(_03065_),
    .A(_00133_),
    .B(_03046_));
 sg13g2_a21oi_1 _10114_ (.A1(_03048_),
    .A2(_03064_),
    .Y(_03066_),
    .B1(_03065_));
 sg13g2_a21oi_1 _10115_ (.A1(_00577_),
    .A2(_03046_),
    .Y(_03067_),
    .B1(_03066_));
 sg13g2_xnor2_1 _10116_ (.Y(_03068_),
    .A(_00132_),
    .B(_03044_));
 sg13g2_nor2_1 _10117_ (.A(_03067_),
    .B(_03068_),
    .Y(_03069_));
 sg13g2_o21ai_1 _10118_ (.B1(_03043_),
    .Y(_03070_),
    .A1(_03045_),
    .A2(_03069_));
 sg13g2_nor2b_1 _10119_ (.A(_00130_),
    .B_N(_03038_),
    .Y(_03071_));
 sg13g2_xnor2_1 _10120_ (.Y(_03072_),
    .A(_00130_),
    .B(_03038_));
 sg13g2_a21oi_1 _10121_ (.A1(_03041_),
    .A2(_03070_),
    .Y(_03073_),
    .B1(_03072_));
 sg13g2_a21oi_1 _10122_ (.A1(_00130_),
    .A2(_03038_),
    .Y(_03074_),
    .B1(_03073_));
 sg13g2_xnor2_1 _10123_ (.Y(_03075_),
    .A(_00610_),
    .B(_03035_));
 sg13g2_nor2b_1 _10124_ (.A(_03074_),
    .B_N(_03075_),
    .Y(_03076_));
 sg13g2_and2_1 _10125_ (.A(_00609_),
    .B(_03032_),
    .X(_03077_));
 sg13g2_xnor2_1 _10126_ (.Y(_03078_),
    .A(_00128_),
    .B(_03032_));
 sg13g2_inv_1 _10127_ (.Y(_03079_),
    .A(_03078_));
 sg13g2_o21ai_1 _10128_ (.B1(_03079_),
    .Y(_03080_),
    .A1(_03037_),
    .A2(_03076_));
 sg13g2_a21oi_1 _10129_ (.A1(_03033_),
    .A2(_03080_),
    .Y(_03081_),
    .B1(_03031_));
 sg13g2_nand3_1 _10130_ (.B(_03033_),
    .C(_03080_),
    .A(_03031_),
    .Y(_03082_));
 sg13g2_nor2b_2 _10131_ (.A(_03081_),
    .B_N(_03082_),
    .Y(_03083_));
 sg13g2_nor2_1 _10132_ (.A(_00137_),
    .B(_03052_),
    .Y(_03084_));
 sg13g2_nand2_1 _10133_ (.Y(_03085_),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[0] ),
    .B(_03054_));
 sg13g2_nor2_1 _10134_ (.A(_03053_),
    .B(_03085_),
    .Y(_03086_));
 sg13g2_nor2_1 _10135_ (.A(_03084_),
    .B(_03086_),
    .Y(_03087_));
 sg13g2_xnor2_1 _10136_ (.Y(_03088_),
    .A(net1884),
    .B(_03051_));
 sg13g2_nor2_1 _10137_ (.A(_03087_),
    .B(_03088_),
    .Y(_03089_));
 sg13g2_a21oi_1 _10138_ (.A1(_00616_),
    .A2(_03051_),
    .Y(_03090_),
    .B1(_03089_));
 sg13g2_nor2b_1 _10139_ (.A(_03090_),
    .B_N(_03050_),
    .Y(_03091_));
 sg13g2_a21oi_1 _10140_ (.A1(_00615_),
    .A2(_03049_),
    .Y(_03092_),
    .B1(_03091_));
 sg13g2_xnor2_1 _10141_ (.Y(_03093_),
    .A(net1883),
    .B(_03047_));
 sg13g2_nor2_1 _10142_ (.A(_03092_),
    .B(_03093_),
    .Y(_03094_));
 sg13g2_a21oi_1 _10143_ (.A1(_00614_),
    .A2(_03047_),
    .Y(_03095_),
    .B1(_03094_));
 sg13g2_xnor2_1 _10144_ (.Y(_03096_),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[5] ),
    .B(_03046_));
 sg13g2_nor2_1 _10145_ (.A(_03095_),
    .B(_03096_),
    .Y(_03097_));
 sg13g2_a21oi_1 _10146_ (.A1(_00613_),
    .A2(_03046_),
    .Y(_03098_),
    .B1(_03097_));
 sg13g2_xnor2_1 _10147_ (.Y(_03099_),
    .A(net1882),
    .B(_03044_));
 sg13g2_nor2_1 _10148_ (.A(_03098_),
    .B(_03099_),
    .Y(_03100_));
 sg13g2_a21oi_1 _10149_ (.A1(_00612_),
    .A2(_03044_),
    .Y(_03101_),
    .B1(_03100_));
 sg13g2_nor2_1 _10150_ (.A(_03043_),
    .B(_03101_),
    .Y(_03102_));
 sg13g2_nor2_1 _10151_ (.A(_03042_),
    .B(_03102_),
    .Y(_03103_));
 sg13g2_xnor2_1 _10152_ (.Y(_03104_),
    .A(net1879),
    .B(_03038_));
 sg13g2_nor2_1 _10153_ (.A(_03103_),
    .B(_03104_),
    .Y(_03105_));
 sg13g2_xnor2_1 _10154_ (.Y(_03106_),
    .A(_00585_),
    .B(_03035_));
 sg13g2_o21ai_1 _10155_ (.B1(_03106_),
    .Y(_03107_),
    .A1(_03071_),
    .A2(_03105_));
 sg13g2_o21ai_1 _10156_ (.B1(_03107_),
    .Y(_03108_),
    .A1(_00129_),
    .A2(_03036_));
 sg13g2_xnor2_1 _10157_ (.Y(_03109_),
    .A(_00587_),
    .B(_03032_));
 sg13g2_and2_1 _10158_ (.A(_03108_),
    .B(_03109_),
    .X(_03110_));
 sg13g2_o21ai_1 _10159_ (.B1(_03031_),
    .Y(_03111_),
    .A1(_03077_),
    .A2(_03110_));
 sg13g2_or3_1 _10160_ (.A(_03031_),
    .B(_03077_),
    .C(_03110_),
    .X(_03112_));
 sg13g2_nand2_2 _10161_ (.Y(_03113_),
    .A(_03111_),
    .B(_03112_));
 sg13g2_nor2_1 _10162_ (.A(net1786),
    .B(_03113_),
    .Y(_03114_));
 sg13g2_a21oi_1 _10163_ (.A1(net1781),
    .A2(_03083_),
    .Y(_03115_),
    .B1(_03114_));
 sg13g2_xnor2_1 _10164_ (.Y(_03116_),
    .A(net1805),
    .B(_03115_));
 sg13g2_nor2_1 _10165_ (.A(_00553_),
    .B(\vgadonut.donut.cA[14] ),
    .Y(_03117_));
 sg13g2_nand2_1 _10166_ (.Y(_03118_),
    .A(_00553_),
    .B(\vgadonut.donut.cA[14] ));
 sg13g2_nand2b_1 _10167_ (.Y(_03119_),
    .B(_03118_),
    .A_N(_03117_));
 sg13g2_o21ai_1 _10168_ (.B1(_03026_),
    .Y(_03120_),
    .A1(_03025_),
    .A2(_03027_));
 sg13g2_xnor2_1 _10169_ (.Y(_03121_),
    .A(_03119_),
    .B(_03120_));
 sg13g2_xnor2_1 _10170_ (.Y(_03122_),
    .A(net1871),
    .B(_03121_));
 sg13g2_a21oi_1 _10171_ (.A1(_03030_),
    .A2(_03111_),
    .Y(_03123_),
    .B1(_03122_));
 sg13g2_nand3_1 _10172_ (.B(_03111_),
    .C(_03122_),
    .A(_03030_),
    .Y(_03124_));
 sg13g2_nand2b_2 _10173_ (.Y(_03125_),
    .B(_03124_),
    .A_N(_03123_));
 sg13g2_a21oi_1 _10174_ (.A1(_00589_),
    .A2(_03029_),
    .Y(_03126_),
    .B1(_03081_));
 sg13g2_and2_1 _10175_ (.A(_00126_),
    .B(_03121_),
    .X(_03127_));
 sg13g2_xnor2_1 _10176_ (.Y(_03128_),
    .A(_00126_),
    .B(_03121_));
 sg13g2_nor2_1 _10177_ (.A(_03126_),
    .B(_03128_),
    .Y(_03129_));
 sg13g2_xor2_1 _10178_ (.B(_03128_),
    .A(_03126_),
    .X(_03130_));
 sg13g2_nand2_1 _10179_ (.Y(_03131_),
    .A(net1796),
    .B(_03130_));
 sg13g2_o21ai_1 _10180_ (.B1(_03131_),
    .Y(_03132_),
    .A1(net1790),
    .A2(_03125_));
 sg13g2_xnor2_1 _10181_ (.Y(_03133_),
    .A(net1622),
    .B(_03132_));
 sg13g2_nand2_1 _10182_ (.Y(_03134_),
    .A(_03116_),
    .B(_03133_));
 sg13g2_xnor2_1 _10183_ (.Y(_03135_),
    .A(_03116_),
    .B(_03133_));
 sg13g2_a21oi_1 _10184_ (.A1(_03118_),
    .A2(_03120_),
    .Y(_03136_),
    .B1(_03117_));
 sg13g2_xor2_1 _10185_ (.B(net1809),
    .A(net1918),
    .X(_03137_));
 sg13g2_xnor2_1 _10186_ (.Y(_03138_),
    .A(_03136_),
    .B(_03137_));
 sg13g2_xor2_1 _10187_ (.B(_03138_),
    .A(_00176_),
    .X(_03139_));
 sg13g2_nor3_1 _10188_ (.A(_03127_),
    .B(_03129_),
    .C(_03139_),
    .Y(_03140_));
 sg13g2_o21ai_1 _10189_ (.B1(_03139_),
    .Y(_03141_),
    .A1(_03127_),
    .A2(_03129_));
 sg13g2_nor2b_2 _10190_ (.A(_03140_),
    .B_N(_03141_),
    .Y(_03142_));
 sg13g2_nor2_1 _10191_ (.A(net1790),
    .B(_03142_),
    .Y(_03143_));
 sg13g2_a21oi_1 _10192_ (.A1(_00608_),
    .A2(_03121_),
    .Y(_03144_),
    .B1(_03123_));
 sg13g2_nor2b_1 _10193_ (.A(_03144_),
    .B_N(_03139_),
    .Y(_03145_));
 sg13g2_xnor2_1 _10194_ (.Y(_03146_),
    .A(_03139_),
    .B(_03144_));
 sg13g2_a21oi_2 _10195_ (.B1(_03143_),
    .Y(_03147_),
    .A2(_03146_),
    .A1(net1790));
 sg13g2_xnor2_1 _10196_ (.Y(_03148_),
    .A(net1805),
    .B(_03147_));
 sg13g2_xnor2_1 _10197_ (.Y(_03149_),
    .A(net1616),
    .B(_03147_));
 sg13g2_inv_1 _10198_ (.Y(_03150_),
    .A(_03149_));
 sg13g2_nor2_1 _10199_ (.A(net1781),
    .B(_03125_),
    .Y(_03151_));
 sg13g2_a21oi_2 _10200_ (.B1(_03151_),
    .Y(_03152_),
    .A2(_03130_),
    .A1(net1781));
 sg13g2_xnor2_1 _10201_ (.Y(_03153_),
    .A(net1805),
    .B(_03152_));
 sg13g2_xnor2_1 _10202_ (.Y(_03154_),
    .A(net1616),
    .B(_03152_));
 sg13g2_nor2_1 _10203_ (.A(net1796),
    .B(_03113_),
    .Y(_03155_));
 sg13g2_a21oi_2 _10204_ (.B1(_03155_),
    .Y(_03156_),
    .A2(_03083_),
    .A1(net1790));
 sg13g2_nor2_1 _10205_ (.A(_03154_),
    .B(_03156_),
    .Y(_03157_));
 sg13g2_xnor2_1 _10206_ (.Y(_03158_),
    .A(net1617),
    .B(_03115_));
 sg13g2_xor2_1 _10207_ (.B(_03109_),
    .A(_03108_),
    .X(_03159_));
 sg13g2_or3_1 _10208_ (.A(_03037_),
    .B(_03076_),
    .C(_03079_),
    .X(_03160_));
 sg13g2_and2_1 _10209_ (.A(_03080_),
    .B(_03160_),
    .X(_03161_));
 sg13g2_mux2_2 _10210_ (.A0(_03159_),
    .A1(_03161_),
    .S(net1790),
    .X(_03162_));
 sg13g2_inv_1 _10211_ (.Y(_03163_),
    .A(_03162_));
 sg13g2_mux2_1 _10212_ (.A0(_03159_),
    .A1(_03161_),
    .S(net1781),
    .X(_03164_));
 sg13g2_xor2_1 _10213_ (.B(_03164_),
    .A(\vgadonut.donut.donuthit.cordicxy.xinvert ),
    .X(_03165_));
 sg13g2_xor2_1 _10214_ (.B(_03164_),
    .A(net1617),
    .X(_03166_));
 sg13g2_or3_1 _10215_ (.A(_03071_),
    .B(_03105_),
    .C(_03106_),
    .X(_03167_));
 sg13g2_nand2_2 _10216_ (.Y(_03168_),
    .A(_03107_),
    .B(_03167_));
 sg13g2_xor2_1 _10217_ (.B(_03075_),
    .A(_03074_),
    .X(_03169_));
 sg13g2_mux2_2 _10218_ (.A0(_03168_),
    .A1(_03169_),
    .S(net1789),
    .X(_03170_));
 sg13g2_nor2_1 _10219_ (.A(_03166_),
    .B(_03170_),
    .Y(_03171_));
 sg13g2_mux2_1 _10220_ (.A0(_03168_),
    .A1(_03169_),
    .S(net1780),
    .X(_03172_));
 sg13g2_xnor2_1 _10221_ (.Y(_03173_),
    .A(net1805),
    .B(_03172_));
 sg13g2_xnor2_1 _10222_ (.Y(_03174_),
    .A(net1617),
    .B(_03172_));
 sg13g2_xor2_1 _10223_ (.B(_03104_),
    .A(_03103_),
    .X(_03175_));
 sg13g2_nand3_1 _10224_ (.B(_03070_),
    .C(_03072_),
    .A(_03041_),
    .Y(_03176_));
 sg13g2_nand2b_2 _10225_ (.Y(_03177_),
    .B(_03176_),
    .A_N(_03073_));
 sg13g2_nor2_1 _10226_ (.A(net1780),
    .B(_03177_),
    .Y(_03178_));
 sg13g2_a21oi_2 _10227_ (.B1(_03178_),
    .Y(_03179_),
    .A2(_03175_),
    .A1(net1780));
 sg13g2_nor2_1 _10228_ (.A(_03174_),
    .B(_03179_),
    .Y(_03180_));
 sg13g2_nor2_1 _10229_ (.A(net1789),
    .B(_03177_),
    .Y(_03181_));
 sg13g2_a21oi_2 _10230_ (.B1(_03181_),
    .Y(_03182_),
    .A2(_03175_),
    .A1(net1789));
 sg13g2_xnor2_1 _10231_ (.Y(_03183_),
    .A(net1804),
    .B(_03182_));
 sg13g2_xnor2_1 _10232_ (.Y(_03184_),
    .A(net1617),
    .B(_03182_));
 sg13g2_xnor2_1 _10233_ (.Y(_03185_),
    .A(_03043_),
    .B(_03101_));
 sg13g2_nor2_1 _10234_ (.A(net1789),
    .B(_03185_),
    .Y(_03186_));
 sg13g2_or3_1 _10235_ (.A(_03043_),
    .B(_03045_),
    .C(_03069_),
    .X(_03187_));
 sg13g2_and2_2 _10236_ (.A(_03070_),
    .B(_03187_),
    .X(_03188_));
 sg13g2_a21oi_2 _10237_ (.B1(_03186_),
    .Y(_03189_),
    .A2(_03188_),
    .A1(net1789));
 sg13g2_nor2_1 _10238_ (.A(_03184_),
    .B(_03189_),
    .Y(_03190_));
 sg13g2_nor2_1 _10239_ (.A(net1780),
    .B(_03185_),
    .Y(_03191_));
 sg13g2_a21oi_2 _10240_ (.B1(_03191_),
    .Y(_03192_),
    .A2(_03188_),
    .A1(net1780));
 sg13g2_xnor2_1 _10241_ (.Y(_03193_),
    .A(net1804),
    .B(_03192_));
 sg13g2_xnor2_1 _10242_ (.Y(_03194_),
    .A(net1616),
    .B(_03192_));
 sg13g2_xnor2_1 _10243_ (.Y(_03195_),
    .A(_03098_),
    .B(_03099_));
 sg13g2_xor2_1 _10244_ (.B(_03068_),
    .A(_03067_),
    .X(_03196_));
 sg13g2_nand2_1 _10245_ (.Y(_03197_),
    .A(net1788),
    .B(_03196_));
 sg13g2_o21ai_1 _10246_ (.B1(_03197_),
    .Y(_03198_),
    .A1(net1788),
    .A2(_03195_));
 sg13g2_nor2b_1 _10247_ (.A(_03194_),
    .B_N(_03198_),
    .Y(_03199_));
 sg13g2_nor2_1 _10248_ (.A(net1779),
    .B(_03195_),
    .Y(_03200_));
 sg13g2_a21oi_2 _10249_ (.B1(_03200_),
    .Y(_03201_),
    .A2(_03196_),
    .A1(net1779));
 sg13g2_xnor2_1 _10250_ (.Y(_03202_),
    .A(net1805),
    .B(_03201_));
 sg13g2_xnor2_1 _10251_ (.Y(_03203_),
    .A(net1616),
    .B(_03201_));
 sg13g2_xnor2_1 _10252_ (.Y(_03204_),
    .A(_03095_),
    .B(_03096_));
 sg13g2_nand3_1 _10253_ (.B(_03064_),
    .C(_03065_),
    .A(_03048_),
    .Y(_03205_));
 sg13g2_nor2b_2 _10254_ (.A(_03066_),
    .B_N(_03205_),
    .Y(_03206_));
 sg13g2_nand2_1 _10255_ (.Y(_03207_),
    .A(net1788),
    .B(_03206_));
 sg13g2_o21ai_1 _10256_ (.B1(_03207_),
    .Y(_03208_),
    .A1(net1787),
    .A2(_03204_));
 sg13g2_nand2b_1 _10257_ (.Y(_03209_),
    .B(_03208_),
    .A_N(_03203_));
 sg13g2_nor2_1 _10258_ (.A(net1779),
    .B(_03204_),
    .Y(_03210_));
 sg13g2_a21oi_2 _10259_ (.B1(_03210_),
    .Y(_03211_),
    .A2(_03206_),
    .A1(net1779));
 sg13g2_xnor2_1 _10260_ (.Y(_03212_),
    .A(net1804),
    .B(_03211_));
 sg13g2_xnor2_1 _10261_ (.Y(_03213_),
    .A(net1616),
    .B(_03211_));
 sg13g2_xnor2_1 _10262_ (.Y(_03214_),
    .A(_03092_),
    .B(_03093_));
 sg13g2_xor2_1 _10263_ (.B(_03063_),
    .A(_03062_),
    .X(_03215_));
 sg13g2_nand2_1 _10264_ (.Y(_03216_),
    .A(net1788),
    .B(_03215_));
 sg13g2_o21ai_1 _10265_ (.B1(_03216_),
    .Y(_03217_),
    .A1(net1787),
    .A2(_03214_));
 sg13g2_nand2b_1 _10266_ (.Y(_03218_),
    .B(_03217_),
    .A_N(_03213_));
 sg13g2_nor2_1 _10267_ (.A(net1778),
    .B(_03214_),
    .Y(_03219_));
 sg13g2_a21oi_2 _10268_ (.B1(_03219_),
    .Y(_03220_),
    .A2(_03215_),
    .A1(net1778));
 sg13g2_xnor2_1 _10269_ (.Y(_03221_),
    .A(net1804),
    .B(_03220_));
 sg13g2_xnor2_1 _10270_ (.Y(_03222_),
    .A(net1616),
    .B(_03220_));
 sg13g2_xnor2_1 _10271_ (.Y(_03223_),
    .A(_03050_),
    .B(_03090_));
 sg13g2_xor2_1 _10272_ (.B(_03060_),
    .A(_03050_),
    .X(_03224_));
 sg13g2_nor2_1 _10273_ (.A(net1778),
    .B(_03224_),
    .Y(_03225_));
 sg13g2_a21oi_2 _10274_ (.B1(_03225_),
    .Y(_03226_),
    .A2(_03223_),
    .A1(net1778));
 sg13g2_or2_1 _10275_ (.X(_03227_),
    .B(_03226_),
    .A(_03222_));
 sg13g2_nor2_1 _10276_ (.A(net1787),
    .B(_03224_),
    .Y(_03228_));
 sg13g2_a21oi_2 _10277_ (.B1(_03228_),
    .Y(_03229_),
    .A2(_03223_),
    .A1(net1787));
 sg13g2_xnor2_1 _10278_ (.Y(_03230_),
    .A(net1804),
    .B(_03229_));
 sg13g2_xnor2_1 _10279_ (.Y(_03231_),
    .A(net1616),
    .B(_03229_));
 sg13g2_xnor2_1 _10280_ (.Y(_03232_),
    .A(_03087_),
    .B(_03088_));
 sg13g2_nor2_1 _10281_ (.A(net1787),
    .B(_03232_),
    .Y(_03233_));
 sg13g2_xnor2_1 _10282_ (.Y(_03234_),
    .A(_03057_),
    .B(_03058_));
 sg13g2_a21oi_2 _10283_ (.B1(_03233_),
    .Y(_03235_),
    .A2(_03234_),
    .A1(net1787));
 sg13g2_nor2_1 _10284_ (.A(_03231_),
    .B(_03235_),
    .Y(_03236_));
 sg13g2_xor2_1 _10285_ (.B(_03235_),
    .A(_03231_),
    .X(_03237_));
 sg13g2_nor2_1 _10286_ (.A(net1778),
    .B(_03232_),
    .Y(_03238_));
 sg13g2_a21oi_1 _10287_ (.A1(net1778),
    .A2(_03234_),
    .Y(_03239_),
    .B1(_03238_));
 sg13g2_xnor2_1 _10288_ (.Y(_03240_),
    .A(net1804),
    .B(_03239_));
 sg13g2_inv_1 _10289_ (.Y(_03241_),
    .A(_03240_));
 sg13g2_xor2_1 _10290_ (.B(_03240_),
    .A(net1620),
    .X(_03242_));
 sg13g2_xnor2_1 _10291_ (.Y(_03243_),
    .A(_03053_),
    .B(_03085_));
 sg13g2_xnor2_1 _10292_ (.Y(_03244_),
    .A(_03053_),
    .B(_03055_));
 sg13g2_nand2_1 _10293_ (.Y(_03245_),
    .A(net1787),
    .B(_03244_));
 sg13g2_o21ai_1 _10294_ (.B1(_03245_),
    .Y(_03246_),
    .A1(net1787),
    .A2(_03243_));
 sg13g2_nor2_1 _10295_ (.A(_03242_),
    .B(_03246_),
    .Y(_03247_));
 sg13g2_nor2_1 _10296_ (.A(net1778),
    .B(_03243_),
    .Y(_03248_));
 sg13g2_a21oi_1 _10297_ (.A1(net1778),
    .A2(_03244_),
    .Y(_03249_),
    .B1(_03248_));
 sg13g2_xnor2_1 _10298_ (.Y(_03250_),
    .A(net1804),
    .B(_03249_));
 sg13g2_inv_1 _10299_ (.Y(_03251_),
    .A(_03250_));
 sg13g2_or2_1 _10300_ (.X(_03252_),
    .B(_03250_),
    .A(net1620));
 sg13g2_xnor2_1 _10301_ (.Y(_03253_),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[0] ),
    .B(_03054_));
 sg13g2_a21oi_1 _10302_ (.A1(net1620),
    .A2(_03250_),
    .Y(_03254_),
    .B1(_03253_));
 sg13g2_a22oi_1 _10303_ (.Y(_03255_),
    .B1(_03252_),
    .B2(_03254_),
    .A2(_03246_),
    .A1(_03242_));
 sg13g2_nor2_1 _10304_ (.A(_03247_),
    .B(_03255_),
    .Y(_03256_));
 sg13g2_a21oi_1 _10305_ (.A1(_03237_),
    .A2(_03256_),
    .Y(_03257_),
    .B1(_03236_));
 sg13g2_xnor2_1 _10306_ (.Y(_03258_),
    .A(_03222_),
    .B(_03226_));
 sg13g2_o21ai_1 _10307_ (.B1(_03227_),
    .Y(_03259_),
    .A1(_03257_),
    .A2(_03258_));
 sg13g2_xor2_1 _10308_ (.B(_03217_),
    .A(_03213_),
    .X(_03260_));
 sg13g2_nand2b_1 _10309_ (.Y(_03261_),
    .B(_03259_),
    .A_N(_03260_));
 sg13g2_nand2_1 _10310_ (.Y(_03262_),
    .A(_03218_),
    .B(_03261_));
 sg13g2_xor2_1 _10311_ (.B(_03208_),
    .A(_03203_),
    .X(_03263_));
 sg13g2_nand2b_1 _10312_ (.Y(_03264_),
    .B(_03262_),
    .A_N(_03263_));
 sg13g2_nand2_1 _10313_ (.Y(_03265_),
    .A(_03209_),
    .B(_03264_));
 sg13g2_xor2_1 _10314_ (.B(_03198_),
    .A(_03194_),
    .X(_03266_));
 sg13g2_inv_1 _10315_ (.Y(_03267_),
    .A(_03266_));
 sg13g2_a21oi_1 _10316_ (.A1(_03265_),
    .A2(_03267_),
    .Y(_03268_),
    .B1(_03199_));
 sg13g2_xnor2_1 _10317_ (.Y(_03269_),
    .A(_03184_),
    .B(_03189_));
 sg13g2_nor2_1 _10318_ (.A(_03268_),
    .B(_03269_),
    .Y(_03270_));
 sg13g2_nor2_1 _10319_ (.A(_03190_),
    .B(_03270_),
    .Y(_03271_));
 sg13g2_xnor2_1 _10320_ (.Y(_03272_),
    .A(_03174_),
    .B(_03179_));
 sg13g2_nor2_1 _10321_ (.A(_03271_),
    .B(_03272_),
    .Y(_03273_));
 sg13g2_nor2_1 _10322_ (.A(_03180_),
    .B(_03273_),
    .Y(_03274_));
 sg13g2_xnor2_1 _10323_ (.Y(_03275_),
    .A(_03166_),
    .B(_03170_));
 sg13g2_nor2_1 _10324_ (.A(_03274_),
    .B(_03275_),
    .Y(_03276_));
 sg13g2_xnor2_1 _10325_ (.Y(_03277_),
    .A(_03158_),
    .B(_03162_));
 sg13g2_o21ai_1 _10326_ (.B1(_03277_),
    .Y(_03278_),
    .A1(_03171_),
    .A2(_03276_));
 sg13g2_o21ai_1 _10327_ (.B1(_03278_),
    .Y(_03279_),
    .A1(_03158_),
    .A2(_03163_));
 sg13g2_xnor2_1 _10328_ (.Y(_03280_),
    .A(_03154_),
    .B(_03156_));
 sg13g2_inv_1 _10329_ (.Y(_03281_),
    .A(_03280_));
 sg13g2_a21oi_1 _10330_ (.A1(_03279_),
    .A2(_03281_),
    .Y(_03282_),
    .B1(_03157_));
 sg13g2_xor2_1 _10331_ (.B(_03149_),
    .A(_03132_),
    .X(_03283_));
 sg13g2_nor2_1 _10332_ (.A(_03282_),
    .B(_03283_),
    .Y(_03284_));
 sg13g2_a21oi_1 _10333_ (.A1(_03132_),
    .A2(_03150_),
    .Y(_03285_),
    .B1(_03284_));
 sg13g2_nor2_1 _10334_ (.A(net1870),
    .B(_03138_),
    .Y(_03286_));
 sg13g2_mux2_1 _10335_ (.A0(_03140_),
    .A1(_00176_),
    .S(_03286_),
    .X(_03287_));
 sg13g2_nand2_1 _10336_ (.Y(_03288_),
    .A(net1781),
    .B(_03287_));
 sg13g2_a21o_1 _10337_ (.A2(_03138_),
    .A1(_00176_),
    .B1(_03145_),
    .X(_03289_));
 sg13g2_o21ai_1 _10338_ (.B1(_03288_),
    .Y(_03290_),
    .A1(net1781),
    .A2(_03289_));
 sg13g2_xor2_1 _10339_ (.B(_03290_),
    .A(net1616),
    .X(_03291_));
 sg13g2_nor2_1 _10340_ (.A(net1781),
    .B(_03142_),
    .Y(_03292_));
 sg13g2_a21oi_2 _10341_ (.B1(_03292_),
    .Y(_03293_),
    .A2(_03146_),
    .A1(net1781));
 sg13g2_nor2_1 _10342_ (.A(_03291_),
    .B(_03293_),
    .Y(_03294_));
 sg13g2_xnor2_1 _10343_ (.Y(_03295_),
    .A(_03291_),
    .B(_03293_));
 sg13g2_nor2_1 _10344_ (.A(_03285_),
    .B(_03295_),
    .Y(_03296_));
 sg13g2_xor2_1 _10345_ (.B(_03295_),
    .A(_03285_),
    .X(_03297_));
 sg13g2_xnor2_1 _10346_ (.Y(_03298_),
    .A(net1609),
    .B(_03297_));
 sg13g2_o21ai_1 _10347_ (.B1(_03134_),
    .Y(_03299_),
    .A1(_03135_),
    .A2(_03298_));
 sg13g2_xor2_1 _10348_ (.B(_03293_),
    .A(net1622),
    .X(_03300_));
 sg13g2_xnor2_1 _10349_ (.Y(_03301_),
    .A(_03153_),
    .B(_03300_));
 sg13g2_nand2_1 _10350_ (.Y(_03302_),
    .A(net1790),
    .B(_03287_));
 sg13g2_o21ai_1 _10351_ (.B1(_03302_),
    .Y(_03303_),
    .A1(net1790),
    .A2(_03289_));
 sg13g2_inv_1 _10352_ (.Y(_03304_),
    .A(_03303_));
 sg13g2_xnor2_1 _10353_ (.Y(_03305_),
    .A(_03291_),
    .B(_03304_));
 sg13g2_nor2_1 _10354_ (.A(_03294_),
    .B(_03296_),
    .Y(_03306_));
 sg13g2_nand2b_1 _10355_ (.Y(_03307_),
    .B(_03306_),
    .A_N(_03305_));
 sg13g2_xnor2_1 _10356_ (.Y(_03308_),
    .A(_03305_),
    .B(_03306_));
 sg13g2_xnor2_1 _10357_ (.Y(_03309_),
    .A(net1609),
    .B(_03308_));
 sg13g2_nor2b_1 _10358_ (.A(_03301_),
    .B_N(_03309_),
    .Y(_03310_));
 sg13g2_xnor2_1 _10359_ (.Y(_03311_),
    .A(_03301_),
    .B(_03309_));
 sg13g2_nand2_1 _10360_ (.Y(_03312_),
    .A(_03299_),
    .B(_03311_));
 sg13g2_xor2_1 _10361_ (.B(_03156_),
    .A(net1628),
    .X(_03313_));
 sg13g2_nand2_1 _10362_ (.Y(_03314_),
    .A(_03165_),
    .B(_03313_));
 sg13g2_xnor2_1 _10363_ (.Y(_03315_),
    .A(_03165_),
    .B(_03313_));
 sg13g2_xor2_1 _10364_ (.B(_03283_),
    .A(_03282_),
    .X(_03316_));
 sg13g2_xnor2_1 _10365_ (.Y(_03317_),
    .A(net1609),
    .B(_03316_));
 sg13g2_o21ai_1 _10366_ (.B1(_03314_),
    .Y(_03318_),
    .A1(_03315_),
    .A2(_03317_));
 sg13g2_xor2_1 _10367_ (.B(_03298_),
    .A(_03135_),
    .X(_03319_));
 sg13g2_xnor2_1 _10368_ (.Y(_03320_),
    .A(net1628),
    .B(_03162_));
 sg13g2_nand2_1 _10369_ (.Y(_03321_),
    .A(_03173_),
    .B(_03320_));
 sg13g2_xnor2_1 _10370_ (.Y(_03322_),
    .A(_03173_),
    .B(_03320_));
 sg13g2_xnor2_1 _10371_ (.Y(_03323_),
    .A(_03279_),
    .B(_03280_));
 sg13g2_xnor2_1 _10372_ (.Y(_03324_),
    .A(net1609),
    .B(_03323_));
 sg13g2_o21ai_1 _10373_ (.B1(_03321_),
    .Y(_03325_),
    .A1(_03322_),
    .A2(_03324_));
 sg13g2_xor2_1 _10374_ (.B(_03317_),
    .A(_03315_),
    .X(_03326_));
 sg13g2_nand2_1 _10375_ (.Y(_03327_),
    .A(_03325_),
    .B(_03326_));
 sg13g2_xor2_1 _10376_ (.B(_03170_),
    .A(net1621),
    .X(_03328_));
 sg13g2_nand2_1 _10377_ (.Y(_03329_),
    .A(_03183_),
    .B(_03328_));
 sg13g2_xnor2_1 _10378_ (.Y(_03330_),
    .A(_03183_),
    .B(_03328_));
 sg13g2_or3_1 _10379_ (.A(_03171_),
    .B(_03276_),
    .C(_03277_),
    .X(_03331_));
 sg13g2_and2_1 _10380_ (.A(_03278_),
    .B(_03331_),
    .X(_03332_));
 sg13g2_xnor2_1 _10381_ (.Y(_03333_),
    .A(net1609),
    .B(_03332_));
 sg13g2_o21ai_1 _10382_ (.B1(_03329_),
    .Y(_03334_),
    .A1(_03330_),
    .A2(_03333_));
 sg13g2_xor2_1 _10383_ (.B(_03324_),
    .A(_03322_),
    .X(_03335_));
 sg13g2_and2_1 _10384_ (.A(_03334_),
    .B(_03335_),
    .X(_03336_));
 sg13g2_xor2_1 _10385_ (.B(_03179_),
    .A(net1621),
    .X(_03337_));
 sg13g2_nand2_1 _10386_ (.Y(_03338_),
    .A(_03193_),
    .B(_03337_));
 sg13g2_xnor2_1 _10387_ (.Y(_03339_),
    .A(_03193_),
    .B(_03337_));
 sg13g2_xor2_1 _10388_ (.B(_03275_),
    .A(_03274_),
    .X(_03340_));
 sg13g2_xnor2_1 _10389_ (.Y(_03341_),
    .A(net1608),
    .B(_03340_));
 sg13g2_o21ai_1 _10390_ (.B1(_03338_),
    .Y(_03342_),
    .A1(_03339_),
    .A2(_03341_));
 sg13g2_xor2_1 _10391_ (.B(_03333_),
    .A(_03330_),
    .X(_03343_));
 sg13g2_nand2_1 _10392_ (.Y(_03344_),
    .A(_03342_),
    .B(_03343_));
 sg13g2_xor2_1 _10393_ (.B(_03189_),
    .A(net1621),
    .X(_03345_));
 sg13g2_nand2_1 _10394_ (.Y(_03346_),
    .A(_03202_),
    .B(_03345_));
 sg13g2_xnor2_1 _10395_ (.Y(_03347_),
    .A(_03202_),
    .B(_03345_));
 sg13g2_xor2_1 _10396_ (.B(_03272_),
    .A(_03271_),
    .X(_03348_));
 sg13g2_xnor2_1 _10397_ (.Y(_03349_),
    .A(net1608),
    .B(_03348_));
 sg13g2_o21ai_1 _10398_ (.B1(_03346_),
    .Y(_03350_),
    .A1(_03347_),
    .A2(_03349_));
 sg13g2_xor2_1 _10399_ (.B(_03341_),
    .A(_03339_),
    .X(_03351_));
 sg13g2_xnor2_1 _10400_ (.Y(_03352_),
    .A(net1620),
    .B(_03198_));
 sg13g2_nand2_1 _10401_ (.Y(_03353_),
    .A(_03212_),
    .B(_03352_));
 sg13g2_xnor2_1 _10402_ (.Y(_03354_),
    .A(_03212_),
    .B(_03352_));
 sg13g2_xor2_1 _10403_ (.B(_03269_),
    .A(_03268_),
    .X(_03355_));
 sg13g2_xnor2_1 _10404_ (.Y(_03356_),
    .A(net1608),
    .B(_03355_));
 sg13g2_o21ai_1 _10405_ (.B1(_03353_),
    .Y(_03357_),
    .A1(_03354_),
    .A2(_03356_));
 sg13g2_xor2_1 _10406_ (.B(_03349_),
    .A(_03347_),
    .X(_03358_));
 sg13g2_xnor2_1 _10407_ (.Y(_03359_),
    .A(net1621),
    .B(_03208_));
 sg13g2_nand2_1 _10408_ (.Y(_03360_),
    .A(_03221_),
    .B(_03359_));
 sg13g2_xnor2_1 _10409_ (.Y(_03361_),
    .A(_03221_),
    .B(_03359_));
 sg13g2_xnor2_1 _10410_ (.Y(_03362_),
    .A(_03265_),
    .B(_03266_));
 sg13g2_xnor2_1 _10411_ (.Y(_03363_),
    .A(net1608),
    .B(_03362_));
 sg13g2_o21ai_1 _10412_ (.B1(_03360_),
    .Y(_03364_),
    .A1(_03361_),
    .A2(_03363_));
 sg13g2_xor2_1 _10413_ (.B(_03356_),
    .A(_03354_),
    .X(_03365_));
 sg13g2_xnor2_1 _10414_ (.Y(_03366_),
    .A(net1620),
    .B(_03217_));
 sg13g2_nand2_1 _10415_ (.Y(_03367_),
    .A(_03230_),
    .B(_03366_));
 sg13g2_xnor2_1 _10416_ (.Y(_03368_),
    .A(_03230_),
    .B(_03366_));
 sg13g2_xnor2_1 _10417_ (.Y(_03369_),
    .A(_03262_),
    .B(_03263_));
 sg13g2_xnor2_1 _10418_ (.Y(_03370_),
    .A(net1608),
    .B(_03369_));
 sg13g2_o21ai_1 _10419_ (.B1(_03367_),
    .Y(_03371_),
    .A1(_03368_),
    .A2(_03370_));
 sg13g2_xor2_1 _10420_ (.B(_03363_),
    .A(_03361_),
    .X(_03372_));
 sg13g2_and2_1 _10421_ (.A(_03371_),
    .B(_03372_),
    .X(_03373_));
 sg13g2_xnor2_1 _10422_ (.Y(_03374_),
    .A(net1620),
    .B(_03226_));
 sg13g2_xnor2_1 _10423_ (.Y(_03375_),
    .A(_03240_),
    .B(_03374_));
 sg13g2_xnor2_1 _10424_ (.Y(_03376_),
    .A(_03259_),
    .B(_03260_));
 sg13g2_xnor2_1 _10425_ (.Y(_03377_),
    .A(net1608),
    .B(_03376_));
 sg13g2_nand2b_1 _10426_ (.Y(_03378_),
    .B(_03375_),
    .A_N(_03377_));
 sg13g2_o21ai_1 _10427_ (.B1(_03378_),
    .Y(_03379_),
    .A1(_03241_),
    .A2(_03374_));
 sg13g2_xor2_1 _10428_ (.B(_03370_),
    .A(_03368_),
    .X(_03380_));
 sg13g2_nand2_1 _10429_ (.Y(_03381_),
    .A(_03379_),
    .B(_03380_));
 sg13g2_xnor2_1 _10430_ (.Y(_03382_),
    .A(net1620),
    .B(_03235_));
 sg13g2_xnor2_1 _10431_ (.Y(_03383_),
    .A(_03250_),
    .B(_03382_));
 sg13g2_xor2_1 _10432_ (.B(_03258_),
    .A(_03257_),
    .X(_03384_));
 sg13g2_xnor2_1 _10433_ (.Y(_03385_),
    .A(net1608),
    .B(_03384_));
 sg13g2_nand2b_1 _10434_ (.Y(_03386_),
    .B(_03383_),
    .A_N(_03385_));
 sg13g2_o21ai_1 _10435_ (.B1(_03386_),
    .Y(_03387_),
    .A1(_03251_),
    .A2(_03382_));
 sg13g2_xnor2_1 _10436_ (.Y(_03388_),
    .A(_03375_),
    .B(_03377_));
 sg13g2_and2_1 _10437_ (.A(_03387_),
    .B(_03388_),
    .X(_03389_));
 sg13g2_xor2_1 _10438_ (.B(_03385_),
    .A(_03383_),
    .X(_03390_));
 sg13g2_xor2_1 _10439_ (.B(_03253_),
    .A(net1804),
    .X(_03391_));
 sg13g2_xor2_1 _10440_ (.B(_03246_),
    .A(net1620),
    .X(_03392_));
 sg13g2_nor2_1 _10441_ (.A(_03391_),
    .B(_03392_),
    .Y(_03393_));
 sg13g2_and2_1 _10442_ (.A(_03391_),
    .B(_03392_),
    .X(_03394_));
 sg13g2_xnor2_1 _10443_ (.Y(_03395_),
    .A(_03237_),
    .B(_03256_));
 sg13g2_xnor2_1 _10444_ (.Y(_03396_),
    .A(net1608),
    .B(_03395_));
 sg13g2_nor2_1 _10445_ (.A(_03393_),
    .B(_03396_),
    .Y(_03397_));
 sg13g2_nor3_2 _10446_ (.A(_03390_),
    .B(_03394_),
    .C(_03397_),
    .Y(_03398_));
 sg13g2_xor2_1 _10447_ (.B(_03388_),
    .A(_03387_),
    .X(_03399_));
 sg13g2_a21oi_1 _10448_ (.A1(_03398_),
    .A2(_03399_),
    .Y(_03400_),
    .B1(_03389_));
 sg13g2_xnor2_1 _10449_ (.Y(_03401_),
    .A(_03379_),
    .B(_03380_));
 sg13g2_o21ai_1 _10450_ (.B1(_03381_),
    .Y(_03402_),
    .A1(_03400_),
    .A2(_03401_));
 sg13g2_xor2_1 _10451_ (.B(_03372_),
    .A(_03371_),
    .X(_03403_));
 sg13g2_a21o_1 _10452_ (.A2(_03403_),
    .A1(_03402_),
    .B1(_03373_),
    .X(_03404_));
 sg13g2_xnor2_1 _10453_ (.Y(_03405_),
    .A(_03364_),
    .B(_03365_));
 sg13g2_nor2b_1 _10454_ (.A(_03405_),
    .B_N(_03404_),
    .Y(_03406_));
 sg13g2_a21o_1 _10455_ (.A2(_03365_),
    .A1(_03364_),
    .B1(_03406_),
    .X(_03407_));
 sg13g2_xnor2_1 _10456_ (.Y(_03408_),
    .A(_03357_),
    .B(_03358_));
 sg13g2_nor2b_1 _10457_ (.A(_03408_),
    .B_N(_03407_),
    .Y(_03409_));
 sg13g2_a21o_1 _10458_ (.A2(_03358_),
    .A1(_03357_),
    .B1(_03409_),
    .X(_03410_));
 sg13g2_xnor2_1 _10459_ (.Y(_03411_),
    .A(_03350_),
    .B(_03351_));
 sg13g2_nor2b_1 _10460_ (.A(_03411_),
    .B_N(_03410_),
    .Y(_03412_));
 sg13g2_a21oi_1 _10461_ (.A1(_03350_),
    .A2(_03351_),
    .Y(_03413_),
    .B1(_03412_));
 sg13g2_xnor2_1 _10462_ (.Y(_03414_),
    .A(_03342_),
    .B(_03343_));
 sg13g2_o21ai_1 _10463_ (.B1(_03344_),
    .Y(_03415_),
    .A1(_03413_),
    .A2(_03414_));
 sg13g2_xor2_1 _10464_ (.B(_03335_),
    .A(_03334_),
    .X(_03416_));
 sg13g2_a21oi_2 _10465_ (.B1(_03336_),
    .Y(_03417_),
    .A2(_03416_),
    .A1(_03415_));
 sg13g2_xnor2_1 _10466_ (.Y(_03418_),
    .A(_03325_),
    .B(_03326_));
 sg13g2_o21ai_1 _10467_ (.B1(_03327_),
    .Y(_03419_),
    .A1(_03417_),
    .A2(_03418_));
 sg13g2_xnor2_1 _10468_ (.Y(_03420_),
    .A(_03318_),
    .B(_03319_));
 sg13g2_nor2b_1 _10469_ (.A(_03420_),
    .B_N(_03419_),
    .Y(_03421_));
 sg13g2_a21oi_1 _10470_ (.A1(_03318_),
    .A2(_03319_),
    .Y(_03422_),
    .B1(_03421_));
 sg13g2_xnor2_1 _10471_ (.Y(_03423_),
    .A(_03299_),
    .B(_03311_));
 sg13g2_o21ai_1 _10472_ (.B1(_03312_),
    .Y(_03424_),
    .A1(_03422_),
    .A2(_03423_));
 sg13g2_a21o_1 _10473_ (.A2(_03300_),
    .A1(_03153_),
    .B1(_03310_),
    .X(_03425_));
 sg13g2_inv_1 _10474_ (.Y(_03426_),
    .A(_03425_));
 sg13g2_xnor2_1 _10475_ (.Y(_03427_),
    .A(net1622),
    .B(_03303_));
 sg13g2_and2_1 _10476_ (.A(_03148_),
    .B(_03427_),
    .X(_03428_));
 sg13g2_xor2_1 _10477_ (.B(_03427_),
    .A(_03148_),
    .X(_03429_));
 sg13g2_o21ai_1 _10478_ (.B1(_03307_),
    .Y(_03430_),
    .A1(_03291_),
    .A2(_03304_));
 sg13g2_xor2_1 _10479_ (.B(_03430_),
    .A(net1609),
    .X(_03431_));
 sg13g2_xnor2_1 _10480_ (.Y(_03432_),
    .A(_03429_),
    .B(_03431_));
 sg13g2_xor2_1 _10481_ (.B(_03432_),
    .A(_03425_),
    .X(_03433_));
 sg13g2_nand2b_1 _10482_ (.Y(_03434_),
    .B(_03424_),
    .A_N(_03433_));
 sg13g2_xor2_1 _10483_ (.B(_03433_),
    .A(_03424_),
    .X(_03435_));
 sg13g2_xor2_1 _10484_ (.B(_03420_),
    .A(_03419_),
    .X(_03436_));
 sg13g2_nor2_1 _10485_ (.A(_03435_),
    .B(_03436_),
    .Y(_03437_));
 sg13g2_xor2_1 _10486_ (.B(_03436_),
    .A(_03435_),
    .X(_03438_));
 sg13g2_xor2_1 _10487_ (.B(_03423_),
    .A(_03422_),
    .X(_03439_));
 sg13g2_inv_1 _10488_ (.Y(_03440_),
    .A(_03439_));
 sg13g2_xor2_1 _10489_ (.B(_03418_),
    .A(_03417_),
    .X(_03441_));
 sg13g2_nand2_1 _10490_ (.Y(_03442_),
    .A(_03439_),
    .B(_03441_));
 sg13g2_xnor2_1 _10491_ (.Y(_03443_),
    .A(_03415_),
    .B(_03416_));
 sg13g2_nor2_1 _10492_ (.A(_03436_),
    .B(_03443_),
    .Y(_03444_));
 sg13g2_xor2_1 _10493_ (.B(_03443_),
    .A(_03436_),
    .X(_03445_));
 sg13g2_xor2_1 _10494_ (.B(_03414_),
    .A(_03413_),
    .X(_03446_));
 sg13g2_nand2_1 _10495_ (.Y(_03447_),
    .A(_03441_),
    .B(_03446_));
 sg13g2_xor2_1 _10496_ (.B(_03411_),
    .A(_03410_),
    .X(_03448_));
 sg13g2_nor2_1 _10497_ (.A(_03443_),
    .B(_03448_),
    .Y(_03449_));
 sg13g2_xor2_1 _10498_ (.B(_03448_),
    .A(_03443_),
    .X(_03450_));
 sg13g2_xor2_1 _10499_ (.B(_03408_),
    .A(_03407_),
    .X(_03451_));
 sg13g2_inv_1 _10500_ (.Y(_03452_),
    .A(_03451_));
 sg13g2_nand2_1 _10501_ (.Y(_03453_),
    .A(_03446_),
    .B(_03452_));
 sg13g2_xor2_1 _10502_ (.B(_03405_),
    .A(_03404_),
    .X(_03454_));
 sg13g2_nor2_1 _10503_ (.A(_03448_),
    .B(_03454_),
    .Y(_03455_));
 sg13g2_xor2_1 _10504_ (.B(_03454_),
    .A(_03448_),
    .X(_03456_));
 sg13g2_xnor2_1 _10505_ (.Y(_03457_),
    .A(_03402_),
    .B(_03403_));
 sg13g2_nor2_1 _10506_ (.A(_03451_),
    .B(_03457_),
    .Y(_03458_));
 sg13g2_xor2_1 _10507_ (.B(_03401_),
    .A(_03400_),
    .X(_03459_));
 sg13g2_nor2b_1 _10508_ (.A(_03454_),
    .B_N(_03459_),
    .Y(_03460_));
 sg13g2_xnor2_1 _10509_ (.Y(_03461_),
    .A(_03454_),
    .B(_03459_));
 sg13g2_xnor2_1 _10510_ (.Y(_03462_),
    .A(_03398_),
    .B(_03399_));
 sg13g2_nor2_1 _10511_ (.A(_03457_),
    .B(_03462_),
    .Y(_03463_));
 sg13g2_o21ai_1 _10512_ (.B1(_03390_),
    .Y(_03464_),
    .A1(_03394_),
    .A2(_03397_));
 sg13g2_nor2b_1 _10513_ (.A(_03398_),
    .B_N(_03464_),
    .Y(_03465_));
 sg13g2_nand2_1 _10514_ (.Y(_03466_),
    .A(_03459_),
    .B(_03465_));
 sg13g2_xor2_1 _10515_ (.B(_03462_),
    .A(_03457_),
    .X(_03467_));
 sg13g2_nor2b_1 _10516_ (.A(_03466_),
    .B_N(_03467_),
    .Y(_03468_));
 sg13g2_nor2_1 _10517_ (.A(_03463_),
    .B(_03468_),
    .Y(_03469_));
 sg13g2_nor2b_1 _10518_ (.A(_03469_),
    .B_N(_03461_),
    .Y(_03470_));
 sg13g2_nor2_1 _10519_ (.A(_03460_),
    .B(_03470_),
    .Y(_03471_));
 sg13g2_xor2_1 _10520_ (.B(_03457_),
    .A(_03451_),
    .X(_03472_));
 sg13g2_nor2b_1 _10521_ (.A(_03471_),
    .B_N(_03472_),
    .Y(_03473_));
 sg13g2_nor2_1 _10522_ (.A(_03458_),
    .B(_03473_),
    .Y(_03474_));
 sg13g2_nor2b_1 _10523_ (.A(_03474_),
    .B_N(_03456_),
    .Y(_03475_));
 sg13g2_nor2_2 _10524_ (.A(_03455_),
    .B(_03475_),
    .Y(_03476_));
 sg13g2_xnor2_1 _10525_ (.Y(_03477_),
    .A(_03446_),
    .B(_03452_));
 sg13g2_o21ai_1 _10526_ (.B1(_03453_),
    .Y(_03478_),
    .A1(_03476_),
    .A2(_03477_));
 sg13g2_a21oi_1 _10527_ (.A1(_03450_),
    .A2(_03478_),
    .Y(_03479_),
    .B1(_03449_));
 sg13g2_xnor2_1 _10528_ (.Y(_03480_),
    .A(_03441_),
    .B(_03446_));
 sg13g2_o21ai_1 _10529_ (.B1(_03447_),
    .Y(_03481_),
    .A1(_03479_),
    .A2(_03480_));
 sg13g2_a21oi_2 _10530_ (.B1(_03444_),
    .Y(_03482_),
    .A2(_03481_),
    .A1(_03445_));
 sg13g2_xnor2_1 _10531_ (.Y(_03483_),
    .A(_03439_),
    .B(_03441_));
 sg13g2_o21ai_1 _10532_ (.B1(_03442_),
    .Y(_03484_),
    .A1(_03482_),
    .A2(_03483_));
 sg13g2_a21oi_1 _10533_ (.A1(_03438_),
    .A2(_03484_),
    .Y(_03485_),
    .B1(_03437_));
 sg13g2_xor2_1 _10534_ (.B(_03431_),
    .A(_03305_),
    .X(_03486_));
 sg13g2_a21o_1 _10535_ (.A2(_03431_),
    .A1(_03429_),
    .B1(_03428_),
    .X(_03487_));
 sg13g2_xnor2_1 _10536_ (.Y(_03488_),
    .A(_03486_),
    .B(_03487_));
 sg13g2_o21ai_1 _10537_ (.B1(_03434_),
    .Y(_03489_),
    .A1(_03426_),
    .A2(_03432_));
 sg13g2_nand2b_1 _10538_ (.Y(_03490_),
    .B(_03489_),
    .A_N(_03488_));
 sg13g2_xor2_1 _10539_ (.B(_03489_),
    .A(_03488_),
    .X(_03491_));
 sg13g2_or2_1 _10540_ (.X(_03492_),
    .B(_03491_),
    .A(_03440_));
 sg13g2_xnor2_1 _10541_ (.Y(_03493_),
    .A(_03440_),
    .B(_03491_));
 sg13g2_xor2_1 _10542_ (.B(_03493_),
    .A(_03485_),
    .X(_03494_));
 sg13g2_nor2_1 _10543_ (.A(net1942),
    .B(net1839),
    .Y(_03495_));
 sg13g2_nor2_1 _10544_ (.A(net1940),
    .B(net1836),
    .Y(_03496_));
 sg13g2_xor2_1 _10545_ (.B(net1836),
    .A(net1940),
    .X(_03497_));
 sg13g2_xnor2_1 _10546_ (.Y(_03498_),
    .A(_03495_),
    .B(_03497_));
 sg13g2_inv_1 _10547_ (.Y(_03499_),
    .A(_03498_));
 sg13g2_xor2_1 _10548_ (.B(net1839),
    .A(net1942),
    .X(_03500_));
 sg13g2_inv_1 _10549_ (.Y(_03501_),
    .A(_03500_));
 sg13g2_nor2_1 _10550_ (.A(net1946),
    .B(net1842),
    .Y(_03502_));
 sg13g2_nor2_1 _10551_ (.A(net1944),
    .B(net1841),
    .Y(_03503_));
 sg13g2_xor2_1 _10552_ (.B(net1841),
    .A(net1944),
    .X(_03504_));
 sg13g2_xnor2_1 _10553_ (.Y(_03505_),
    .A(_03502_),
    .B(_03504_));
 sg13g2_xor2_1 _10554_ (.B(net1842),
    .A(net1946),
    .X(_03506_));
 sg13g2_nor2_1 _10555_ (.A(net1949),
    .B(net1847),
    .Y(_03507_));
 sg13g2_nor2_1 _10556_ (.A(net1948),
    .B(net1844),
    .Y(_03508_));
 sg13g2_xor2_1 _10557_ (.B(net1844),
    .A(net1948),
    .X(_03509_));
 sg13g2_xnor2_1 _10558_ (.Y(_03510_),
    .A(net1949),
    .B(net1847));
 sg13g2_nor2_1 _10559_ (.A(net1952),
    .B(net1848),
    .Y(_03511_));
 sg13g2_nor2b_1 _10560_ (.A(_03510_),
    .B_N(_03511_),
    .Y(_03512_));
 sg13g2_xnor2_1 _10561_ (.Y(_03513_),
    .A(net1951),
    .B(net1849));
 sg13g2_or2_1 _10562_ (.X(_03514_),
    .B(net1851),
    .A(net1953));
 sg13g2_xnor2_1 _10563_ (.Y(_03515_),
    .A(net1953),
    .B(net1851));
 sg13g2_nor2_1 _10564_ (.A(net1955),
    .B(net1852),
    .Y(_03516_));
 sg13g2_nor2b_1 _10565_ (.A(_03515_),
    .B_N(_03516_),
    .Y(_03517_));
 sg13g2_xnor2_1 _10566_ (.Y(_03518_),
    .A(net1955),
    .B(net1852));
 sg13g2_or2_1 _10567_ (.X(_03519_),
    .B(\vgadonut.donut.sA[3] ),
    .A(net1957));
 sg13g2_xnor2_1 _10568_ (.Y(_03520_),
    .A(net1957),
    .B(net1853));
 sg13g2_nor2_1 _10569_ (.A(\vgadonut.donut.cAcB[2] ),
    .B(\vgadonut.donut.sA[2] ),
    .Y(_03521_));
 sg13g2_nor2b_1 _10570_ (.A(_03520_),
    .B_N(_03521_),
    .Y(_03522_));
 sg13g2_xor2_1 _10571_ (.B(net1854),
    .A(\vgadonut.donut.cAcB[2] ),
    .X(_03523_));
 sg13g2_nand2_1 _10572_ (.Y(_03524_),
    .A(\vgadonut.donut.cAcB[1] ),
    .B(\vgadonut.donut.sA[1] ));
 sg13g2_xor2_1 _10573_ (.B(\vgadonut.donut.sA[1] ),
    .A(\vgadonut.donut.cAcB[1] ),
    .X(_03525_));
 sg13g2_nor3_1 _10574_ (.A(\vgadonut.donut.cAcB[0] ),
    .B(\vgadonut.donut.sA[0] ),
    .C(_03525_),
    .Y(_03526_));
 sg13g2_xnor2_1 _10575_ (.Y(_03527_),
    .A(_03523_),
    .B(_03524_));
 sg13g2_nor4_1 _10576_ (.A(\vgadonut.donut.cAcB[0] ),
    .B(\vgadonut.donut.sA[0] ),
    .C(_03525_),
    .D(_03527_),
    .Y(_03528_));
 sg13g2_a21o_1 _10577_ (.A2(_03524_),
    .A1(_03523_),
    .B1(_03528_),
    .X(_03529_));
 sg13g2_xnor2_1 _10578_ (.Y(_03530_),
    .A(_03520_),
    .B(_03521_));
 sg13g2_a21oi_1 _10579_ (.A1(_03529_),
    .A2(_03530_),
    .Y(_03531_),
    .B1(_03522_));
 sg13g2_xor2_1 _10580_ (.B(_03519_),
    .A(_03518_),
    .X(_03532_));
 sg13g2_nand2b_1 _10581_ (.Y(_03533_),
    .B(_03532_),
    .A_N(_03531_));
 sg13g2_o21ai_1 _10582_ (.B1(_03533_),
    .Y(_03534_),
    .A1(_03518_),
    .A2(_03519_));
 sg13g2_xnor2_1 _10583_ (.Y(_03535_),
    .A(_03515_),
    .B(_03516_));
 sg13g2_a21oi_1 _10584_ (.A1(_03534_),
    .A2(_03535_),
    .Y(_03536_),
    .B1(_03517_));
 sg13g2_xor2_1 _10585_ (.B(_03514_),
    .A(_03513_),
    .X(_03537_));
 sg13g2_nand2b_1 _10586_ (.Y(_03538_),
    .B(_03537_),
    .A_N(_03536_));
 sg13g2_o21ai_1 _10587_ (.B1(_03538_),
    .Y(_03539_),
    .A1(_03513_),
    .A2(_03514_));
 sg13g2_xnor2_1 _10588_ (.Y(_03540_),
    .A(_03510_),
    .B(_03511_));
 sg13g2_a21o_1 _10589_ (.A2(_03540_),
    .A1(_03539_),
    .B1(_03512_),
    .X(_03541_));
 sg13g2_xnor2_1 _10590_ (.Y(_03542_),
    .A(_03507_),
    .B(_03509_));
 sg13g2_nor2b_1 _10591_ (.A(_03542_),
    .B_N(_03541_),
    .Y(_03543_));
 sg13g2_a21o_1 _10592_ (.A2(_03509_),
    .A1(_03507_),
    .B1(_03543_),
    .X(_03544_));
 sg13g2_nand2_1 _10593_ (.Y(_03545_),
    .A(_03506_),
    .B(_03544_));
 sg13g2_o21ai_1 _10594_ (.B1(_03508_),
    .Y(_03546_),
    .A1(_03506_),
    .A2(_03543_));
 sg13g2_nand2_1 _10595_ (.Y(_03547_),
    .A(_03545_),
    .B(_03546_));
 sg13g2_a21oi_1 _10596_ (.A1(_03545_),
    .A2(_03546_),
    .Y(_03548_),
    .B1(_03505_));
 sg13g2_a21oi_1 _10597_ (.A1(_03502_),
    .A2(_03504_),
    .Y(_03549_),
    .B1(_03548_));
 sg13g2_o21ai_1 _10598_ (.B1(_03503_),
    .Y(_03550_),
    .A1(_03500_),
    .A2(_03548_));
 sg13g2_o21ai_1 _10599_ (.B1(_03550_),
    .Y(_03551_),
    .A1(_03501_),
    .A2(_03549_));
 sg13g2_and2_1 _10600_ (.A(_03499_),
    .B(_03551_),
    .X(_03552_));
 sg13g2_a21oi_1 _10601_ (.A1(_03495_),
    .A2(_03497_),
    .Y(_03553_),
    .B1(_03552_));
 sg13g2_nor2_1 _10602_ (.A(net1938),
    .B(net1833),
    .Y(_03554_));
 sg13g2_xor2_1 _10603_ (.B(net1833),
    .A(net1938),
    .X(_03555_));
 sg13g2_nor2_1 _10604_ (.A(_03496_),
    .B(_03555_),
    .Y(_03556_));
 sg13g2_xor2_1 _10605_ (.B(_03555_),
    .A(_03496_),
    .X(_03557_));
 sg13g2_nor2_1 _10606_ (.A(_03553_),
    .B(_03556_),
    .Y(_03558_));
 sg13g2_xnor2_1 _10607_ (.Y(_03559_),
    .A(_03553_),
    .B(_03557_));
 sg13g2_inv_1 _10608_ (.Y(_03560_),
    .A(_03559_));
 sg13g2_and2_1 _10609_ (.A(_03494_),
    .B(_03559_),
    .X(_03561_));
 sg13g2_nand2_1 _10610_ (.Y(_03562_),
    .A(_03494_),
    .B(_03560_));
 sg13g2_xnor2_1 _10611_ (.Y(_03563_),
    .A(_03494_),
    .B(_03560_));
 sg13g2_xor2_1 _10612_ (.B(_03484_),
    .A(_03438_),
    .X(_03564_));
 sg13g2_xnor2_1 _10613_ (.Y(_03565_),
    .A(_03499_),
    .B(_03551_));
 sg13g2_inv_1 _10614_ (.Y(_03566_),
    .A(_03565_));
 sg13g2_and2_1 _10615_ (.A(_03564_),
    .B(_03566_),
    .X(_03567_));
 sg13g2_nand2_1 _10616_ (.Y(_03568_),
    .A(_03564_),
    .B(_03565_));
 sg13g2_xnor2_1 _10617_ (.Y(_03569_),
    .A(_03564_),
    .B(_03566_));
 sg13g2_inv_1 _10618_ (.Y(_03570_),
    .A(_03569_));
 sg13g2_xor2_1 _10619_ (.B(_03483_),
    .A(_03482_),
    .X(_03571_));
 sg13g2_xor2_1 _10620_ (.B(_03503_),
    .A(_03500_),
    .X(_03572_));
 sg13g2_xnor2_1 _10621_ (.Y(_03573_),
    .A(_03549_),
    .B(_03572_));
 sg13g2_nand2b_1 _10622_ (.Y(_03574_),
    .B(_03571_),
    .A_N(_03573_));
 sg13g2_xnor2_1 _10623_ (.Y(_03575_),
    .A(_03571_),
    .B(_03573_));
 sg13g2_xor2_1 _10624_ (.B(_03547_),
    .A(_03505_),
    .X(_03576_));
 sg13g2_xor2_1 _10625_ (.B(_03481_),
    .A(_03445_),
    .X(_03577_));
 sg13g2_nand2b_1 _10626_ (.Y(_03578_),
    .B(_03577_),
    .A_N(_03576_));
 sg13g2_and2_1 _10627_ (.A(_03576_),
    .B(_03577_),
    .X(_03579_));
 sg13g2_xnor2_1 _10628_ (.Y(_03580_),
    .A(_03576_),
    .B(_03577_));
 sg13g2_xor2_1 _10629_ (.B(_03480_),
    .A(_03479_),
    .X(_03581_));
 sg13g2_inv_1 _10630_ (.Y(_03582_),
    .A(_03581_));
 sg13g2_xor2_1 _10631_ (.B(_03508_),
    .A(_03506_),
    .X(_03583_));
 sg13g2_xnor2_1 _10632_ (.Y(_03584_),
    .A(_03544_),
    .B(_03583_));
 sg13g2_nand2_1 _10633_ (.Y(_03585_),
    .A(_03581_),
    .B(_03584_));
 sg13g2_xor2_1 _10634_ (.B(_03584_),
    .A(_03581_),
    .X(_03586_));
 sg13g2_xor2_1 _10635_ (.B(_03542_),
    .A(_03541_),
    .X(_03587_));
 sg13g2_xor2_1 _10636_ (.B(_03478_),
    .A(_03450_),
    .X(_03588_));
 sg13g2_nand2b_1 _10637_ (.Y(_03589_),
    .B(_03588_),
    .A_N(_03587_));
 sg13g2_and2_1 _10638_ (.A(_03587_),
    .B(_03588_),
    .X(_03590_));
 sg13g2_xnor2_1 _10639_ (.Y(_03591_),
    .A(_03587_),
    .B(_03588_));
 sg13g2_xor2_1 _10640_ (.B(_03477_),
    .A(_03476_),
    .X(_03592_));
 sg13g2_xnor2_1 _10641_ (.Y(_03593_),
    .A(_03539_),
    .B(_03540_));
 sg13g2_inv_1 _10642_ (.Y(_03594_),
    .A(_03593_));
 sg13g2_nand2_1 _10643_ (.Y(_03595_),
    .A(_03592_),
    .B(_03593_));
 sg13g2_xnor2_1 _10644_ (.Y(_03596_),
    .A(_03592_),
    .B(_03594_));
 sg13g2_xnor2_1 _10645_ (.Y(_03597_),
    .A(_03456_),
    .B(_03474_));
 sg13g2_xnor2_1 _10646_ (.Y(_03598_),
    .A(_03536_),
    .B(_03537_));
 sg13g2_nand2_1 _10647_ (.Y(_03599_),
    .A(_03597_),
    .B(_03598_));
 sg13g2_nand2b_1 _10648_ (.Y(_03600_),
    .B(_03597_),
    .A_N(_03598_));
 sg13g2_xnor2_1 _10649_ (.Y(_03601_),
    .A(_03597_),
    .B(_03598_));
 sg13g2_xnor2_1 _10650_ (.Y(_03602_),
    .A(_03471_),
    .B(_03472_));
 sg13g2_xnor2_1 _10651_ (.Y(_03603_),
    .A(_03534_),
    .B(_03535_));
 sg13g2_inv_1 _10652_ (.Y(_03604_),
    .A(_03603_));
 sg13g2_and2_1 _10653_ (.A(_03602_),
    .B(_03603_),
    .X(_03605_));
 sg13g2_xnor2_1 _10654_ (.Y(_03606_),
    .A(_03602_),
    .B(_03604_));
 sg13g2_xnor2_1 _10655_ (.Y(_03607_),
    .A(_03461_),
    .B(_03469_));
 sg13g2_xnor2_1 _10656_ (.Y(_03608_),
    .A(_03531_),
    .B(_03532_));
 sg13g2_nand2b_1 _10657_ (.Y(_03609_),
    .B(_03607_),
    .A_N(_03608_));
 sg13g2_xnor2_1 _10658_ (.Y(_03610_),
    .A(_03607_),
    .B(_03608_));
 sg13g2_xnor2_1 _10659_ (.Y(_03611_),
    .A(_03466_),
    .B(_03467_));
 sg13g2_xor2_1 _10660_ (.B(_03530_),
    .A(_03529_),
    .X(_03612_));
 sg13g2_nand2_1 _10661_ (.Y(_03613_),
    .A(_03611_),
    .B(_03612_));
 sg13g2_nor2b_1 _10662_ (.A(_03612_),
    .B_N(_03611_),
    .Y(_03614_));
 sg13g2_xnor2_1 _10663_ (.Y(_03615_),
    .A(_03611_),
    .B(_03612_));
 sg13g2_xnor2_1 _10664_ (.Y(_03616_),
    .A(_03459_),
    .B(_03465_));
 sg13g2_xnor2_1 _10665_ (.Y(_03617_),
    .A(_03526_),
    .B(_03527_));
 sg13g2_nand2b_1 _10666_ (.Y(_03618_),
    .B(_03617_),
    .A_N(_03616_));
 sg13g2_o21ai_1 _10667_ (.B1(_03613_),
    .Y(_03619_),
    .A1(_03615_),
    .A2(_03618_));
 sg13g2_nor2b_1 _10668_ (.A(_03610_),
    .B_N(_03619_),
    .Y(_03620_));
 sg13g2_a21o_1 _10669_ (.A2(_03608_),
    .A1(_03607_),
    .B1(_03620_),
    .X(_03621_));
 sg13g2_nor2b_1 _10670_ (.A(_03606_),
    .B_N(_03621_),
    .Y(_03622_));
 sg13g2_a21oi_1 _10671_ (.A1(_03602_),
    .A2(_03604_),
    .Y(_03623_),
    .B1(_03622_));
 sg13g2_o21ai_1 _10672_ (.B1(_03599_),
    .Y(_03624_),
    .A1(_03601_),
    .A2(_03623_));
 sg13g2_nor2b_1 _10673_ (.A(_03596_),
    .B_N(_03624_),
    .Y(_03625_));
 sg13g2_a21oi_1 _10674_ (.A1(_03592_),
    .A2(_03594_),
    .Y(_03626_),
    .B1(_03625_));
 sg13g2_nand2b_1 _10675_ (.Y(_03627_),
    .B(_03591_),
    .A_N(_03626_));
 sg13g2_a21o_1 _10676_ (.A2(_03627_),
    .A1(_03589_),
    .B1(_03586_),
    .X(_03628_));
 sg13g2_o21ai_1 _10677_ (.B1(_03628_),
    .Y(_03629_),
    .A1(_03582_),
    .A2(_03584_));
 sg13g2_nand2_1 _10678_ (.Y(_03630_),
    .A(_03580_),
    .B(_03629_));
 sg13g2_a21oi_1 _10679_ (.A1(_03578_),
    .A2(_03630_),
    .Y(_03631_),
    .B1(_03575_));
 sg13g2_a21o_1 _10680_ (.A2(_03573_),
    .A1(_03571_),
    .B1(_03631_),
    .X(_03632_));
 sg13g2_a21oi_2 _10681_ (.B1(_03567_),
    .Y(_03633_),
    .A2(_03632_),
    .A1(_03570_));
 sg13g2_nor2b_1 _10682_ (.A(_03633_),
    .B_N(_03563_),
    .Y(_03634_));
 sg13g2_xor2_1 _10683_ (.B(_03633_),
    .A(_03563_),
    .X(_03635_));
 sg13g2_nand2_1 _10684_ (.Y(_03636_),
    .A(_03616_),
    .B(_03617_));
 sg13g2_and2_1 _10685_ (.A(_03615_),
    .B(_03636_),
    .X(_03637_));
 sg13g2_o21ai_1 _10686_ (.B1(_03610_),
    .Y(_03638_),
    .A1(_03614_),
    .A2(_03637_));
 sg13g2_nand2_1 _10687_ (.Y(_03639_),
    .A(_03609_),
    .B(_03638_));
 sg13g2_and2_1 _10688_ (.A(_03606_),
    .B(_03639_),
    .X(_03640_));
 sg13g2_nor2_1 _10689_ (.A(_03605_),
    .B(_03640_),
    .Y(_03641_));
 sg13g2_o21ai_1 _10690_ (.B1(_03601_),
    .Y(_03642_),
    .A1(_03605_),
    .A2(_03640_));
 sg13g2_nand2_1 _10691_ (.Y(_03643_),
    .A(_03600_),
    .B(_03642_));
 sg13g2_nand2_1 _10692_ (.Y(_03644_),
    .A(_03596_),
    .B(_03643_));
 sg13g2_nand2_1 _10693_ (.Y(_03645_),
    .A(_03595_),
    .B(_03644_));
 sg13g2_a21oi_1 _10694_ (.A1(_03595_),
    .A2(_03644_),
    .Y(_03646_),
    .B1(_03591_));
 sg13g2_nor2_1 _10695_ (.A(_03590_),
    .B(_03646_),
    .Y(_03647_));
 sg13g2_o21ai_1 _10696_ (.B1(_03586_),
    .Y(_03648_),
    .A1(_03590_),
    .A2(_03646_));
 sg13g2_and2_1 _10697_ (.A(_03585_),
    .B(_03648_),
    .X(_03649_));
 sg13g2_nor2_1 _10698_ (.A(_03580_),
    .B(_03649_),
    .Y(_03650_));
 sg13g2_o21ai_1 _10699_ (.B1(_03575_),
    .Y(_03651_),
    .A1(_03579_),
    .A2(_03650_));
 sg13g2_and2_1 _10700_ (.A(_03574_),
    .B(_03651_),
    .X(_03652_));
 sg13g2_o21ai_1 _10701_ (.B1(_03568_),
    .Y(_03653_),
    .A1(_03570_),
    .A2(_03652_));
 sg13g2_nand2b_1 _10702_ (.Y(_03654_),
    .B(_03653_),
    .A_N(_03563_));
 sg13g2_xor2_1 _10703_ (.B(_03653_),
    .A(_03563_),
    .X(_03655_));
 sg13g2_mux2_1 _10704_ (.A0(_03635_),
    .A1(_03655_),
    .S(net1573),
    .X(_03656_));
 sg13g2_xnor2_1 _10705_ (.Y(_03657_),
    .A(net1548),
    .B(_03656_));
 sg13g2_xnor2_1 _10706_ (.Y(_03658_),
    .A(_03570_),
    .B(_03652_));
 sg13g2_xnor2_1 _10707_ (.Y(_03659_),
    .A(_03570_),
    .B(_03632_));
 sg13g2_mux2_1 _10708_ (.A0(_03658_),
    .A1(_03659_),
    .S(net1572),
    .X(_03660_));
 sg13g2_xor2_1 _10709_ (.B(_03660_),
    .A(net1591),
    .X(_03661_));
 sg13g2_mux2_1 _10710_ (.A0(_03658_),
    .A1(_03659_),
    .S(net1581),
    .X(_03662_));
 sg13g2_xnor2_1 _10711_ (.Y(_03663_),
    .A(net1548),
    .B(_03662_));
 sg13g2_or3_1 _10712_ (.A(_03575_),
    .B(_03579_),
    .C(_03650_),
    .X(_03664_));
 sg13g2_and2_1 _10713_ (.A(_03651_),
    .B(_03664_),
    .X(_03665_));
 sg13g2_nand2_1 _10714_ (.Y(_03666_),
    .A(net1581),
    .B(_03665_));
 sg13g2_nand3_1 _10715_ (.B(_03578_),
    .C(_03630_),
    .A(_03575_),
    .Y(_03667_));
 sg13g2_nand2b_1 _10716_ (.Y(_03668_),
    .B(_03667_),
    .A_N(_03631_));
 sg13g2_o21ai_1 _10717_ (.B1(_03666_),
    .Y(_03669_),
    .A1(net1581),
    .A2(_03668_));
 sg13g2_xnor2_1 _10718_ (.Y(_03670_),
    .A(net1591),
    .B(_03669_));
 sg13g2_nor2_1 _10719_ (.A(net1572),
    .B(_03668_),
    .Y(_03671_));
 sg13g2_a21oi_1 _10720_ (.A1(net1572),
    .A2(_03665_),
    .Y(_03672_),
    .B1(_03671_));
 sg13g2_xnor2_1 _10721_ (.Y(_03673_),
    .A(net1548),
    .B(_03672_));
 sg13g2_xor2_1 _10722_ (.B(_03629_),
    .A(_03580_),
    .X(_03674_));
 sg13g2_xnor2_1 _10723_ (.Y(_03675_),
    .A(_03580_),
    .B(_03649_));
 sg13g2_nor2_1 _10724_ (.A(net1572),
    .B(_03675_),
    .Y(_03676_));
 sg13g2_a21oi_1 _10725_ (.A1(net1572),
    .A2(_03674_),
    .Y(_03677_),
    .B1(_03676_));
 sg13g2_xor2_1 _10726_ (.B(_03677_),
    .A(net1591),
    .X(_03678_));
 sg13g2_nor2_1 _10727_ (.A(net1581),
    .B(_03675_),
    .Y(_03679_));
 sg13g2_a21oi_1 _10728_ (.A1(net1581),
    .A2(_03674_),
    .Y(_03680_),
    .B1(_03679_));
 sg13g2_xnor2_1 _10729_ (.Y(_03681_),
    .A(net1548),
    .B(_03680_));
 sg13g2_nand3_1 _10730_ (.B(_03589_),
    .C(_03627_),
    .A(_03586_),
    .Y(_03682_));
 sg13g2_nand2_1 _10731_ (.Y(_03683_),
    .A(_03628_),
    .B(_03682_));
 sg13g2_xnor2_1 _10732_ (.Y(_03684_),
    .A(_03586_),
    .B(_03647_));
 sg13g2_nand2_1 _10733_ (.Y(_03685_),
    .A(net1581),
    .B(_03684_));
 sg13g2_o21ai_1 _10734_ (.B1(_03685_),
    .Y(_03686_),
    .A1(net1581),
    .A2(_03683_));
 sg13g2_xor2_1 _10735_ (.B(_03686_),
    .A(net1591),
    .X(_03687_));
 sg13g2_inv_1 _10736_ (.Y(_03688_),
    .A(_03687_));
 sg13g2_nand2_1 _10737_ (.Y(_03689_),
    .A(_03681_),
    .B(_03688_));
 sg13g2_nand2_1 _10738_ (.Y(_03690_),
    .A(net1572),
    .B(_03684_));
 sg13g2_o21ai_1 _10739_ (.B1(_03690_),
    .Y(_03691_),
    .A1(net1572),
    .A2(_03683_));
 sg13g2_xnor2_1 _10740_ (.Y(_03692_),
    .A(net1548),
    .B(_03691_));
 sg13g2_xor2_1 _10741_ (.B(_03645_),
    .A(_03591_),
    .X(_03693_));
 sg13g2_xor2_1 _10742_ (.B(_03626_),
    .A(_03591_),
    .X(_03694_));
 sg13g2_mux2_1 _10743_ (.A0(_03693_),
    .A1(_03694_),
    .S(net1572),
    .X(_03695_));
 sg13g2_xnor2_1 _10744_ (.Y(_03696_),
    .A(net1591),
    .B(_03695_));
 sg13g2_nor2_1 _10745_ (.A(_03692_),
    .B(_03696_),
    .Y(_03697_));
 sg13g2_mux2_1 _10746_ (.A0(_03693_),
    .A1(_03694_),
    .S(net1581),
    .X(_03698_));
 sg13g2_xnor2_1 _10747_ (.Y(_03699_),
    .A(net1548),
    .B(_03698_));
 sg13g2_xor2_1 _10748_ (.B(_03643_),
    .A(_03596_),
    .X(_03700_));
 sg13g2_nand2_1 _10749_ (.Y(_03701_),
    .A(net1582),
    .B(_03700_));
 sg13g2_xor2_1 _10750_ (.B(_03624_),
    .A(_03596_),
    .X(_03702_));
 sg13g2_o21ai_1 _10751_ (.B1(_03701_),
    .Y(_03703_),
    .A1(net1582),
    .A2(_03702_));
 sg13g2_xnor2_1 _10752_ (.Y(_03704_),
    .A(net1591),
    .B(_03703_));
 sg13g2_nor2_1 _10753_ (.A(net1573),
    .B(_03702_),
    .Y(_03705_));
 sg13g2_a21oi_1 _10754_ (.A1(net1573),
    .A2(_03700_),
    .Y(_03706_),
    .B1(_03705_));
 sg13g2_xnor2_1 _10755_ (.Y(_03707_),
    .A(net1549),
    .B(_03706_));
 sg13g2_xnor2_1 _10756_ (.Y(_03708_),
    .A(_03601_),
    .B(_03623_));
 sg13g2_xnor2_1 _10757_ (.Y(_03709_),
    .A(_03601_),
    .B(_03641_));
 sg13g2_nand2_1 _10758_ (.Y(_03710_),
    .A(net1582),
    .B(_03709_));
 sg13g2_o21ai_1 _10759_ (.B1(_03710_),
    .Y(_03711_),
    .A1(net1582),
    .A2(_03708_));
 sg13g2_xnor2_1 _10760_ (.Y(_03712_),
    .A(net1592),
    .B(_03711_));
 sg13g2_nor2_1 _10761_ (.A(net1573),
    .B(_03708_),
    .Y(_03713_));
 sg13g2_a21oi_1 _10762_ (.A1(net1573),
    .A2(_03709_),
    .Y(_03714_),
    .B1(_03713_));
 sg13g2_xnor2_1 _10763_ (.Y(_03715_),
    .A(net1548),
    .B(_03714_));
 sg13g2_xnor2_1 _10764_ (.Y(_03716_),
    .A(_03606_),
    .B(_03639_));
 sg13g2_xnor2_1 _10765_ (.Y(_03717_),
    .A(_03606_),
    .B(_03621_));
 sg13g2_nand2_1 _10766_ (.Y(_03718_),
    .A(net1575),
    .B(_03717_));
 sg13g2_o21ai_1 _10767_ (.B1(_03718_),
    .Y(_03719_),
    .A1(net1575),
    .A2(_03716_));
 sg13g2_xnor2_1 _10768_ (.Y(_03720_),
    .A(net1591),
    .B(_03719_));
 sg13g2_nand2_1 _10769_ (.Y(_03721_),
    .A(net1584),
    .B(_03717_));
 sg13g2_o21ai_1 _10770_ (.B1(_03721_),
    .Y(_03722_),
    .A1(net1584),
    .A2(_03716_));
 sg13g2_xnor2_1 _10771_ (.Y(_03723_),
    .A(net1548),
    .B(_03722_));
 sg13g2_or3_1 _10772_ (.A(_03610_),
    .B(_03614_),
    .C(_03637_),
    .X(_03724_));
 sg13g2_and2_1 _10773_ (.A(_03638_),
    .B(_03724_),
    .X(_03725_));
 sg13g2_xor2_1 _10774_ (.B(_03619_),
    .A(_03610_),
    .X(_03726_));
 sg13g2_nor2_1 _10775_ (.A(net1584),
    .B(_03726_),
    .Y(_03727_));
 sg13g2_a21oi_1 _10776_ (.A1(net1584),
    .A2(_03725_),
    .Y(_03728_),
    .B1(_03727_));
 sg13g2_xnor2_1 _10777_ (.Y(_03729_),
    .A(net1592),
    .B(_03728_));
 sg13g2_or2_1 _10778_ (.X(_03730_),
    .B(_03729_),
    .A(_03723_));
 sg13g2_nand2_1 _10779_ (.Y(_03731_),
    .A(net1575),
    .B(_03725_));
 sg13g2_o21ai_1 _10780_ (.B1(_03731_),
    .Y(_03732_),
    .A1(net1575),
    .A2(_03726_));
 sg13g2_xnor2_1 _10781_ (.Y(_03733_),
    .A(_01529_),
    .B(_03732_));
 sg13g2_xor2_1 _10782_ (.B(_03636_),
    .A(_03615_),
    .X(_03734_));
 sg13g2_xor2_1 _10783_ (.B(_03618_),
    .A(_03615_),
    .X(_03735_));
 sg13g2_mux2_1 _10784_ (.A0(_03734_),
    .A1(_03735_),
    .S(net1575),
    .X(_03736_));
 sg13g2_xnor2_1 _10785_ (.Y(_03737_),
    .A(net1592),
    .B(_03736_));
 sg13g2_and2_1 _10786_ (.A(_03733_),
    .B(_03737_),
    .X(_03738_));
 sg13g2_and2_1 _10787_ (.A(net1584),
    .B(_03735_),
    .X(_03739_));
 sg13g2_a21oi_1 _10788_ (.A1(net1575),
    .A2(_03734_),
    .Y(_03740_),
    .B1(_03739_));
 sg13g2_xor2_1 _10789_ (.B(_03617_),
    .A(_03616_),
    .X(_03741_));
 sg13g2_xnor2_1 _10790_ (.Y(_03742_),
    .A(net1592),
    .B(_03741_));
 sg13g2_xnor2_1 _10791_ (.Y(_03743_),
    .A(_01529_),
    .B(_03740_));
 sg13g2_nor2_1 _10792_ (.A(_03742_),
    .B(_03743_),
    .Y(_03744_));
 sg13g2_xnor2_1 _10793_ (.Y(_03745_),
    .A(_03733_),
    .B(_03737_));
 sg13g2_nor3_1 _10794_ (.A(_03742_),
    .B(_03743_),
    .C(_03745_),
    .Y(_03746_));
 sg13g2_nor2_1 _10795_ (.A(_03738_),
    .B(_03746_),
    .Y(_03747_));
 sg13g2_xor2_1 _10796_ (.B(_03729_),
    .A(_03723_),
    .X(_03748_));
 sg13g2_o21ai_1 _10797_ (.B1(_03748_),
    .Y(_03749_),
    .A1(_03738_),
    .A2(_03746_));
 sg13g2_xnor2_1 _10798_ (.Y(_03750_),
    .A(_03715_),
    .B(_03720_));
 sg13g2_a21oi_1 _10799_ (.A1(_03730_),
    .A2(_03749_),
    .Y(_03751_),
    .B1(_03750_));
 sg13g2_a21oi_1 _10800_ (.A1(_03715_),
    .A2(_03720_),
    .Y(_03752_),
    .B1(_03751_));
 sg13g2_xnor2_1 _10801_ (.Y(_03753_),
    .A(_03707_),
    .B(_03712_));
 sg13g2_nor2_1 _10802_ (.A(_03752_),
    .B(_03753_),
    .Y(_03754_));
 sg13g2_a21oi_1 _10803_ (.A1(_03707_),
    .A2(_03712_),
    .Y(_03755_),
    .B1(_03754_));
 sg13g2_xnor2_1 _10804_ (.Y(_03756_),
    .A(_03699_),
    .B(_03704_));
 sg13g2_nor2_1 _10805_ (.A(_03755_),
    .B(_03756_),
    .Y(_03757_));
 sg13g2_a21oi_1 _10806_ (.A1(_03699_),
    .A2(_03704_),
    .Y(_03758_),
    .B1(_03757_));
 sg13g2_xnor2_1 _10807_ (.Y(_03759_),
    .A(_03692_),
    .B(_03696_));
 sg13g2_nor2_1 _10808_ (.A(_03758_),
    .B(_03759_),
    .Y(_03760_));
 sg13g2_nor2_1 _10809_ (.A(_03697_),
    .B(_03760_),
    .Y(_03761_));
 sg13g2_xor2_1 _10810_ (.B(_03687_),
    .A(_03681_),
    .X(_03762_));
 sg13g2_inv_1 _10811_ (.Y(_03763_),
    .A(_03762_));
 sg13g2_o21ai_1 _10812_ (.B1(_03763_),
    .Y(_03764_),
    .A1(_03697_),
    .A2(_03760_));
 sg13g2_xnor2_1 _10813_ (.Y(_03765_),
    .A(_03673_),
    .B(_03678_));
 sg13g2_a21oi_1 _10814_ (.A1(_03689_),
    .A2(_03764_),
    .Y(_03766_),
    .B1(_03765_));
 sg13g2_a21oi_1 _10815_ (.A1(_03673_),
    .A2(_03678_),
    .Y(_03767_),
    .B1(_03766_));
 sg13g2_xnor2_1 _10816_ (.Y(_03768_),
    .A(_03663_),
    .B(_03670_));
 sg13g2_nor2_1 _10817_ (.A(_03767_),
    .B(_03768_),
    .Y(_03769_));
 sg13g2_a21oi_1 _10818_ (.A1(_03663_),
    .A2(_03670_),
    .Y(_03770_),
    .B1(_03769_));
 sg13g2_xnor2_1 _10819_ (.Y(_03771_),
    .A(_03657_),
    .B(_03661_));
 sg13g2_nor2_1 _10820_ (.A(_03770_),
    .B(_03771_),
    .Y(_03772_));
 sg13g2_a21oi_1 _10821_ (.A1(_03657_),
    .A2(_03661_),
    .Y(_03773_),
    .B1(_03772_));
 sg13g2_xor2_1 _10822_ (.B(_03290_),
    .A(net1805),
    .X(_03774_));
 sg13g2_and2_1 _10823_ (.A(_03427_),
    .B(_03774_),
    .X(_03775_));
 sg13g2_nor3_1 _10824_ (.A(_03305_),
    .B(_03431_),
    .C(_03775_),
    .Y(_03776_));
 sg13g2_a21oi_1 _10825_ (.A1(_03486_),
    .A2(_03487_),
    .Y(_03777_),
    .B1(_03776_));
 sg13g2_a22oi_1 _10826_ (.Y(_03778_),
    .B1(_03777_),
    .B2(_03490_),
    .A2(_03775_),
    .A1(_03486_));
 sg13g2_nor2_1 _10827_ (.A(_03435_),
    .B(_03778_),
    .Y(_03779_));
 sg13g2_nand2_1 _10828_ (.Y(_03780_),
    .A(_03435_),
    .B(_03778_));
 sg13g2_nand2b_1 _10829_ (.Y(_03781_),
    .B(_03780_),
    .A_N(_03779_));
 sg13g2_o21ai_1 _10830_ (.B1(_03492_),
    .Y(_03782_),
    .A1(_03485_),
    .A2(_03493_));
 sg13g2_xor2_1 _10831_ (.B(_03782_),
    .A(_03781_),
    .X(_03783_));
 sg13g2_nor2_1 _10832_ (.A(net1936),
    .B(\vgadonut.donut.sA[14] ),
    .Y(_03784_));
 sg13g2_xor2_1 _10833_ (.B(\vgadonut.donut.sA[14] ),
    .A(net1936),
    .X(_03785_));
 sg13g2_nand2_1 _10834_ (.Y(_03786_),
    .A(_03554_),
    .B(_03785_));
 sg13g2_xnor2_1 _10835_ (.Y(_03787_),
    .A(_03554_),
    .B(_03785_));
 sg13g2_a21oi_1 _10836_ (.A1(_03496_),
    .A2(_03555_),
    .Y(_03788_),
    .B1(_03558_));
 sg13g2_xnor2_1 _10837_ (.Y(_03789_),
    .A(_03787_),
    .B(_03788_));
 sg13g2_nor2_1 _10838_ (.A(_03783_),
    .B(_03789_),
    .Y(_03790_));
 sg13g2_nor2b_1 _10839_ (.A(_03783_),
    .B_N(_03789_),
    .Y(_03791_));
 sg13g2_xor2_1 _10840_ (.B(_03789_),
    .A(_03783_),
    .X(_03792_));
 sg13g2_a21oi_1 _10841_ (.A1(_03562_),
    .A2(_03654_),
    .Y(_03793_),
    .B1(_03792_));
 sg13g2_nand3_1 _10842_ (.B(_03654_),
    .C(_03792_),
    .A(_03562_),
    .Y(_03794_));
 sg13g2_nor2b_1 _10843_ (.A(_03793_),
    .B_N(_03794_),
    .Y(_03795_));
 sg13g2_o21ai_1 _10844_ (.B1(_03792_),
    .Y(_03796_),
    .A1(_03561_),
    .A2(_03634_));
 sg13g2_or3_1 _10845_ (.A(_03561_),
    .B(_03634_),
    .C(_03792_),
    .X(_03797_));
 sg13g2_and2_1 _10846_ (.A(_03796_),
    .B(_03797_),
    .X(_03798_));
 sg13g2_mux2_1 _10847_ (.A0(_03795_),
    .A1(_03798_),
    .S(net1583),
    .X(_03799_));
 sg13g2_xnor2_1 _10848_ (.Y(_03800_),
    .A(_01529_),
    .B(_03799_));
 sg13g2_mux2_1 _10849_ (.A0(_03635_),
    .A1(_03655_),
    .S(net1582),
    .X(_03801_));
 sg13g2_xor2_1 _10850_ (.B(_03801_),
    .A(net1591),
    .X(_03802_));
 sg13g2_xnor2_1 _10851_ (.Y(_03803_),
    .A(_03800_),
    .B(_03802_));
 sg13g2_nor2_1 _10852_ (.A(_03773_),
    .B(_03803_),
    .Y(_03804_));
 sg13g2_xor2_1 _10853_ (.B(_03803_),
    .A(_03773_),
    .X(_03805_));
 sg13g2_xor2_1 _10854_ (.B(_03768_),
    .A(_03767_),
    .X(_03806_));
 sg13g2_xnor2_1 _10855_ (.Y(_03807_),
    .A(_03805_),
    .B(_03806_));
 sg13g2_xnor2_1 _10856_ (.Y(_03808_),
    .A(_03761_),
    .B(_03763_));
 sg13g2_nand3_1 _10857_ (.B(_03764_),
    .C(_03765_),
    .A(_03689_),
    .Y(_03809_));
 sg13g2_nor2b_1 _10858_ (.A(_03766_),
    .B_N(_03809_),
    .Y(_03810_));
 sg13g2_xor2_1 _10859_ (.B(_03759_),
    .A(_03758_),
    .X(_03811_));
 sg13g2_xor2_1 _10860_ (.B(_03756_),
    .A(_03755_),
    .X(_03812_));
 sg13g2_or3_1 _10861_ (.A(_03806_),
    .B(_03811_),
    .C(_03812_),
    .X(_03813_));
 sg13g2_xor2_1 _10862_ (.B(_03771_),
    .A(_03770_),
    .X(_03814_));
 sg13g2_a21o_1 _10863_ (.A2(_03812_),
    .A1(_03811_),
    .B1(_03806_),
    .X(_03815_));
 sg13g2_a22oi_1 _10864_ (.Y(_03816_),
    .B1(_03814_),
    .B2(_03815_),
    .A2(_03813_),
    .A1(_03810_));
 sg13g2_nand2b_1 _10865_ (.Y(_03817_),
    .B(_03808_),
    .A_N(_03816_));
 sg13g2_a21oi_1 _10866_ (.A1(_03811_),
    .A2(_03814_),
    .Y(_03818_),
    .B1(_03810_));
 sg13g2_a21o_1 _10867_ (.A2(_03811_),
    .A1(_03806_),
    .B1(_03814_),
    .X(_03819_));
 sg13g2_xor2_1 _10868_ (.B(_03753_),
    .A(_03752_),
    .X(_03820_));
 sg13g2_xnor2_1 _10869_ (.Y(_03821_),
    .A(_03747_),
    .B(_03748_));
 sg13g2_and2_1 _10870_ (.A(_03812_),
    .B(_03821_),
    .X(_03822_));
 sg13g2_o21ai_1 _10871_ (.B1(_03820_),
    .Y(_03823_),
    .A1(_03811_),
    .A2(_03822_));
 sg13g2_and3_1 _10872_ (.X(_03824_),
    .A(_03730_),
    .B(_03749_),
    .C(_03750_));
 sg13g2_or2_1 _10873_ (.X(_03825_),
    .B(_03824_),
    .A(_03751_));
 sg13g2_xnor2_1 _10874_ (.Y(_03826_),
    .A(_03744_),
    .B(_03745_));
 sg13g2_a21o_1 _10875_ (.A2(_03826_),
    .A1(_03821_),
    .B1(_03812_),
    .X(_03827_));
 sg13g2_or3_1 _10876_ (.A(_03812_),
    .B(_03821_),
    .C(_03826_),
    .X(_03828_));
 sg13g2_a22oi_1 _10877_ (.Y(_03829_),
    .B1(_03828_),
    .B2(_03820_),
    .A2(_03827_),
    .A1(_03811_));
 sg13g2_o21ai_1 _10878_ (.B1(_03823_),
    .Y(_03830_),
    .A1(_03825_),
    .A2(_03829_));
 sg13g2_a21o_1 _10879_ (.A2(_03812_),
    .A1(_03806_),
    .B1(_03808_),
    .X(_03831_));
 sg13g2_a22oi_1 _10880_ (.Y(_03832_),
    .B1(_03830_),
    .B2(_03831_),
    .A2(_03819_),
    .A1(_03810_));
 sg13g2_o21ai_1 _10881_ (.B1(_03817_),
    .Y(_03833_),
    .A1(_03818_),
    .A2(_03832_));
 sg13g2_nor2b_1 _10882_ (.A(_03807_),
    .B_N(_03833_),
    .Y(_03834_));
 sg13g2_xnor2_1 _10883_ (.Y(\vgadonut.donut.donuthit.cordicxz.x2out[8] ),
    .A(_03807_),
    .B(_03833_));
 sg13g2_a21oi_1 _10884_ (.A1(_03800_),
    .A2(_03802_),
    .Y(_03835_),
    .B1(_03804_));
 sg13g2_a21oi_1 _10885_ (.A1(_03780_),
    .A2(_03782_),
    .Y(_03836_),
    .B1(_03779_));
 sg13g2_or2_1 _10886_ (.X(_03837_),
    .B(_03778_),
    .A(_03491_));
 sg13g2_xnor2_1 _10887_ (.Y(_03838_),
    .A(_03491_),
    .B(_03778_));
 sg13g2_xor2_1 _10888_ (.B(_03838_),
    .A(_03836_),
    .X(_03839_));
 sg13g2_inv_1 _10889_ (.Y(_03840_),
    .A(_03839_));
 sg13g2_o21ai_1 _10890_ (.B1(_03786_),
    .Y(_03841_),
    .A1(_03787_),
    .A2(_03788_));
 sg13g2_xor2_1 _10891_ (.B(net1830),
    .A(net1935),
    .X(_03842_));
 sg13g2_xnor2_1 _10892_ (.Y(_03843_),
    .A(_03784_),
    .B(_03842_));
 sg13g2_xnor2_1 _10893_ (.Y(_03844_),
    .A(_03841_),
    .B(_03843_));
 sg13g2_nand2_1 _10894_ (.Y(_03845_),
    .A(_03839_),
    .B(_03844_));
 sg13g2_xnor2_1 _10895_ (.Y(_03846_),
    .A(_03839_),
    .B(_03844_));
 sg13g2_nor2b_1 _10896_ (.A(_03790_),
    .B_N(_03796_),
    .Y(_03847_));
 sg13g2_xnor2_1 _10897_ (.Y(_03848_),
    .A(_03846_),
    .B(_03847_));
 sg13g2_nor2_1 _10898_ (.A(_03791_),
    .B(_03793_),
    .Y(_03849_));
 sg13g2_nand2b_1 _10899_ (.Y(_03850_),
    .B(_03846_),
    .A_N(_03849_));
 sg13g2_xor2_1 _10900_ (.B(_03849_),
    .A(_03846_),
    .X(_03851_));
 sg13g2_mux2_1 _10901_ (.A0(_03848_),
    .A1(_03851_),
    .S(net1574),
    .X(_03852_));
 sg13g2_xnor2_1 _10902_ (.Y(_03853_),
    .A(_01529_),
    .B(_03852_));
 sg13g2_mux2_1 _10903_ (.A0(_03795_),
    .A1(_03798_),
    .S(net1574),
    .X(_03854_));
 sg13g2_xor2_1 _10904_ (.B(_03854_),
    .A(net1593),
    .X(_03855_));
 sg13g2_nor2_1 _10905_ (.A(_03853_),
    .B(_03855_),
    .Y(_03856_));
 sg13g2_xnor2_1 _10906_ (.Y(_03857_),
    .A(_03853_),
    .B(_03855_));
 sg13g2_nor2_1 _10907_ (.A(_03835_),
    .B(_03857_),
    .Y(_03858_));
 sg13g2_xor2_1 _10908_ (.B(_03857_),
    .A(_03835_),
    .X(_03859_));
 sg13g2_xnor2_1 _10909_ (.Y(_03860_),
    .A(_03814_),
    .B(_03859_));
 sg13g2_a21oi_1 _10910_ (.A1(_03805_),
    .A2(_03806_),
    .Y(_03861_),
    .B1(_03834_));
 sg13g2_nor2_1 _10911_ (.A(_03860_),
    .B(_03861_),
    .Y(_03862_));
 sg13g2_xor2_1 _10912_ (.B(_03861_),
    .A(_03860_),
    .X(\vgadonut.donut.donuthit.cordicxz.x2out[9] ));
 sg13g2_nor2_1 _10913_ (.A(_03856_),
    .B(_03858_),
    .Y(_03863_));
 sg13g2_o21ai_1 _10914_ (.B1(_03837_),
    .Y(_03864_),
    .A1(_03836_),
    .A2(_03838_));
 sg13g2_and2_1 _10915_ (.A(_03844_),
    .B(_03864_),
    .X(_03865_));
 sg13g2_nand2b_1 _10916_ (.Y(_03866_),
    .B(_03864_),
    .A_N(_03844_));
 sg13g2_xor2_1 _10917_ (.B(_03864_),
    .A(_03844_),
    .X(_03867_));
 sg13g2_o21ai_1 _10918_ (.B1(_03845_),
    .Y(_03868_),
    .A1(_03846_),
    .A2(_03847_));
 sg13g2_xor2_1 _10919_ (.B(_03868_),
    .A(_03867_),
    .X(_03869_));
 sg13g2_nand2_1 _10920_ (.Y(_03870_),
    .A(net1583),
    .B(_03869_));
 sg13g2_o21ai_1 _10921_ (.B1(_03850_),
    .Y(_03871_),
    .A1(_03840_),
    .A2(_03844_));
 sg13g2_nand2b_1 _10922_ (.Y(_03872_),
    .B(_03871_),
    .A_N(_03867_));
 sg13g2_xor2_1 _10923_ (.B(_03871_),
    .A(_03867_),
    .X(_03873_));
 sg13g2_o21ai_1 _10924_ (.B1(_03870_),
    .Y(_03874_),
    .A1(net1583),
    .A2(_03873_));
 sg13g2_xnor2_1 _10925_ (.Y(_03875_),
    .A(net1549),
    .B(_03874_));
 sg13g2_mux2_1 _10926_ (.A0(_03848_),
    .A1(_03851_),
    .S(net1583),
    .X(_03876_));
 sg13g2_xnor2_1 _10927_ (.Y(_03877_),
    .A(net1593),
    .B(_03876_));
 sg13g2_nor2_1 _10928_ (.A(_03875_),
    .B(_03877_),
    .Y(_03878_));
 sg13g2_xnor2_1 _10929_ (.Y(_03879_),
    .A(_03875_),
    .B(_03877_));
 sg13g2_nor2_1 _10930_ (.A(_03863_),
    .B(_03879_),
    .Y(_03880_));
 sg13g2_xor2_1 _10931_ (.B(_03879_),
    .A(_03863_),
    .X(_03881_));
 sg13g2_nand2_1 _10932_ (.Y(_03882_),
    .A(_03805_),
    .B(_03881_));
 sg13g2_xnor2_1 _10933_ (.Y(_03883_),
    .A(_03805_),
    .B(_03881_));
 sg13g2_a21oi_1 _10934_ (.A1(_03814_),
    .A2(_03859_),
    .Y(_03884_),
    .B1(_03862_));
 sg13g2_xor2_1 _10935_ (.B(_03884_),
    .A(_03883_),
    .X(\vgadonut.donut.donuthit.cordicxz.x2out[10] ));
 sg13g2_nor2_1 _10936_ (.A(_03878_),
    .B(_03880_),
    .Y(_03885_));
 sg13g2_xnor2_1 _10937_ (.Y(_03886_),
    .A(_03778_),
    .B(_03844_));
 sg13g2_a21oi_1 _10938_ (.A1(_03866_),
    .A2(_03872_),
    .Y(_03887_),
    .B1(_03886_));
 sg13g2_a21oi_1 _10939_ (.A1(_03778_),
    .A2(_03844_),
    .Y(_03888_),
    .B1(_03887_));
 sg13g2_a21oi_1 _10940_ (.A1(_03867_),
    .A2(_03868_),
    .Y(_03889_),
    .B1(_03865_));
 sg13g2_xnor2_1 _10941_ (.Y(_03890_),
    .A(_03886_),
    .B(_03889_));
 sg13g2_mux2_1 _10942_ (.A0(_03888_),
    .A1(_03890_),
    .S(net1583),
    .X(_03891_));
 sg13g2_xnor2_1 _10943_ (.Y(_03892_),
    .A(net1549),
    .B(_03891_));
 sg13g2_nand2_1 _10944_ (.Y(_03893_),
    .A(net1574),
    .B(_03869_));
 sg13g2_o21ai_1 _10945_ (.B1(_03893_),
    .Y(_03894_),
    .A1(net1574),
    .A2(_03873_));
 sg13g2_xnor2_1 _10946_ (.Y(_03895_),
    .A(net1593),
    .B(_03894_));
 sg13g2_nand2b_1 _10947_ (.Y(_03896_),
    .B(_03895_),
    .A_N(_03892_));
 sg13g2_xnor2_1 _10948_ (.Y(_03897_),
    .A(_03892_),
    .B(_03895_));
 sg13g2_o21ai_1 _10949_ (.B1(_03897_),
    .Y(_03898_),
    .A1(_03878_),
    .A2(_03880_));
 sg13g2_xnor2_1 _10950_ (.Y(_03899_),
    .A(_03885_),
    .B(_03897_));
 sg13g2_xnor2_1 _10951_ (.Y(_03900_),
    .A(_03859_),
    .B(_03899_));
 sg13g2_o21ai_1 _10952_ (.B1(_03882_),
    .Y(_03901_),
    .A1(_03883_),
    .A2(_03884_));
 sg13g2_nor2b_1 _10953_ (.A(_03900_),
    .B_N(_03901_),
    .Y(_03902_));
 sg13g2_xnor2_1 _10954_ (.Y(\vgadonut.donut.donuthit.cordicxz.x2out[11] ),
    .A(_03900_),
    .B(_03901_));
 sg13g2_mux2_1 _10955_ (.A0(_03888_),
    .A1(_03890_),
    .S(net1574),
    .X(_03903_));
 sg13g2_xnor2_1 _10956_ (.Y(_03904_),
    .A(net1593),
    .B(_03903_));
 sg13g2_xor2_1 _10957_ (.B(_03904_),
    .A(_03892_),
    .X(_03905_));
 sg13g2_a21oi_1 _10958_ (.A1(_03896_),
    .A2(_03898_),
    .Y(_03906_),
    .B1(_03905_));
 sg13g2_nand3_1 _10959_ (.B(_03898_),
    .C(_03905_),
    .A(_03896_),
    .Y(_03907_));
 sg13g2_nand2b_2 _10960_ (.Y(_03908_),
    .B(_03907_),
    .A_N(_03906_));
 sg13g2_nor2b_1 _10961_ (.A(_03908_),
    .B_N(_03881_),
    .Y(_03909_));
 sg13g2_xnor2_1 _10962_ (.Y(_03910_),
    .A(_03881_),
    .B(_03908_));
 sg13g2_a21o_1 _10963_ (.A2(_03899_),
    .A1(_03859_),
    .B1(_03902_),
    .X(_03911_));
 sg13g2_xor2_1 _10964_ (.B(_03911_),
    .A(_03910_),
    .X(\vgadonut.donut.donuthit.cordicxz.x2out[12] ));
 sg13g2_a21o_1 _10965_ (.A2(_03911_),
    .A1(_03910_),
    .B1(_03909_),
    .X(_03912_));
 sg13g2_xor2_1 _10966_ (.B(_03908_),
    .A(_03899_),
    .X(_03913_));
 sg13g2_xnor2_1 _10967_ (.Y(\vgadonut.donut.donuthit.cordicxz.x2out[13] ),
    .A(_03912_),
    .B(_03913_));
 sg13g2_nor4_2 _10968_ (.A(net1800),
    .B(_02943_),
    .C(_02944_),
    .Y(_03914_),
    .D(_02951_));
 sg13g2_nor4_2 _10969_ (.A(net1800),
    .B(_02943_),
    .C(_02944_),
    .Y(_03915_),
    .D(_02951_));
 sg13g2_nor4_2 _10970_ (.A(net1800),
    .B(_02943_),
    .C(_02944_),
    .Y(_03916_),
    .D(_02951_));
 sg13g2_or2_1 _10971_ (.X(_03917_),
    .B(_03914_),
    .A(_00654_));
 sg13g2_or2_1 _10972_ (.X(_03918_),
    .B(_02953_),
    .A(_02946_));
 sg13g2_nor3_1 _10973_ (.A(\vgadonut.donut.v_count[7] ),
    .B(\vgadonut.donut.v_count[6] ),
    .C(\vgadonut.donut.v_count[8] ),
    .Y(_03919_));
 sg13g2_nand2_1 _10974_ (.Y(_03920_),
    .A(\vgadonut.donut.v_count[9] ),
    .B(_03919_));
 sg13g2_nor4_1 _10975_ (.A(\vgadonut.donut.v_count[5] ),
    .B(\vgadonut.donut.v_count[4] ),
    .C(_02974_),
    .D(_02980_),
    .Y(_03921_));
 sg13g2_nor2b_1 _10976_ (.A(_03920_),
    .B_N(_03921_),
    .Y(_03922_));
 sg13g2_nand2b_1 _10977_ (.Y(_03923_),
    .B(_03921_),
    .A_N(_03920_));
 sg13g2_and2_1 _10978_ (.A(_02946_),
    .B(_03914_),
    .X(_03924_));
 sg13g2_nand2_2 _10979_ (.Y(_03925_),
    .A(net1774),
    .B(net1761));
 sg13g2_nand3_1 _10980_ (.B(\vgadonut.donut.v_count[9] ),
    .C(_03919_),
    .A(_06848_),
    .Y(_03926_));
 sg13g2_nor4_2 _10981_ (.A(\vgadonut.donut.v_count[4] ),
    .B(_02974_),
    .C(_02980_),
    .Y(_03927_),
    .D(_03926_));
 sg13g2_and2_1 _10982_ (.A(_02946_),
    .B(_03915_),
    .X(_03928_));
 sg13g2_nand2_2 _10983_ (.Y(_03929_),
    .A(_02946_),
    .B(_03915_));
 sg13g2_nand2_2 _10984_ (.Y(_03930_),
    .A(net1760),
    .B(net1757));
 sg13g2_and2_2 _10985_ (.A(_02946_),
    .B(_03916_),
    .X(_03931_));
 sg13g2_nand2_1 _10986_ (.Y(_03932_),
    .A(_02946_),
    .B(_03916_));
 sg13g2_nand2_1 _10987_ (.Y(_03933_),
    .A(net1777),
    .B(_03931_));
 sg13g2_and4_2 _10988_ (.A(net1974),
    .B(_03917_),
    .C(_03918_),
    .D(net1726),
    .X(_03934_));
 sg13g2_nand4_1 _10989_ (.B(_03917_),
    .C(_03918_),
    .A(net1974),
    .Y(_03935_),
    .D(net1726));
 sg13g2_a21oi_1 _10990_ (.A1(net1867),
    .A2(net1670),
    .Y(_03936_),
    .B1(net1987));
 sg13g2_nand2_1 _10991_ (.Y(_03937_),
    .A(net1987),
    .B(net1867));
 sg13g2_a21oi_1 _10992_ (.A1(net1755),
    .A2(_03937_),
    .Y(_03938_),
    .B1(net1658));
 sg13g2_nor2_1 _10993_ (.A(net1988),
    .B(_03938_),
    .Y(_00223_));
 sg13g2_nand2_1 _10994_ (.Y(_03939_),
    .A(\vgadonut.donut.rx6[1] ),
    .B(net1866));
 sg13g2_xor2_1 _10995_ (.B(net1866),
    .A(\vgadonut.donut.rx6[1] ),
    .X(_03940_));
 sg13g2_nand2b_1 _10996_ (.Y(_03941_),
    .B(_03940_),
    .A_N(_03937_));
 sg13g2_xor2_1 _10997_ (.B(_03940_),
    .A(_03937_),
    .X(_03942_));
 sg13g2_nor3_1 _10998_ (.A(net1763),
    .B(net1658),
    .C(_03942_),
    .Y(_03943_));
 sg13g2_a21o_1 _10999_ (.A2(net1658),
    .A1(net2073),
    .B1(_03943_),
    .X(_00224_));
 sg13g2_nor2_1 _11000_ (.A(net2017),
    .B(_01892_),
    .Y(_03944_));
 sg13g2_and2_1 _11001_ (.A(net2017),
    .B(_01892_),
    .X(_03945_));
 sg13g2_nor3_1 _11002_ (.A(net1699),
    .B(_03944_),
    .C(_03945_),
    .Y(_00226_));
 sg13g2_nor2_1 _11003_ (.A(_00640_),
    .B(_01894_),
    .Y(_03946_));
 sg13g2_xnor2_1 _11004_ (.Y(_03947_),
    .A(net2252),
    .B(_01894_));
 sg13g2_and2_1 _11005_ (.A(_03945_),
    .B(_03947_),
    .X(_03948_));
 sg13g2_o21ai_1 _11006_ (.B1(net1678),
    .Y(_03949_),
    .A1(_03945_),
    .A2(_03947_));
 sg13g2_nor2_1 _11007_ (.A(_03948_),
    .B(_03949_),
    .Y(_00227_));
 sg13g2_nor2_1 _11008_ (.A(_03946_),
    .B(_03948_),
    .Y(_03950_));
 sg13g2_nand2_1 _11009_ (.Y(_03951_),
    .A(net2249),
    .B(_01799_));
 sg13g2_xnor2_1 _11010_ (.Y(_03952_),
    .A(net2249),
    .B(_01799_));
 sg13g2_o21ai_1 _11011_ (.B1(net1678),
    .Y(_03953_),
    .A1(_03950_),
    .A2(_03952_));
 sg13g2_a21oi_1 _11012_ (.A1(_03950_),
    .A2(_03952_),
    .Y(_00228_),
    .B1(_03953_));
 sg13g2_o21ai_1 _11013_ (.B1(_03951_),
    .Y(_03954_),
    .A1(_03950_),
    .A2(_03952_));
 sg13g2_nor2_1 _11014_ (.A(_00641_),
    .B(_01804_),
    .Y(_03955_));
 sg13g2_nand2_1 _11015_ (.Y(_03956_),
    .A(_00641_),
    .B(_01804_));
 sg13g2_nor2b_1 _11016_ (.A(_03955_),
    .B_N(_03956_),
    .Y(_03957_));
 sg13g2_o21ai_1 _11017_ (.B1(net1679),
    .Y(_03958_),
    .A1(_03954_),
    .A2(_03957_));
 sg13g2_a21oi_1 _11018_ (.A1(_03954_),
    .A2(_03957_),
    .Y(_00229_),
    .B1(_03958_));
 sg13g2_a21o_1 _11019_ (.A2(_03956_),
    .A1(_03954_),
    .B1(_03955_),
    .X(_03959_));
 sg13g2_xor2_1 _11020_ (.B(_01846_),
    .A(net2207),
    .X(_03960_));
 sg13g2_and2_1 _11021_ (.A(_03959_),
    .B(_03960_),
    .X(_03961_));
 sg13g2_o21ai_1 _11022_ (.B1(net1678),
    .Y(_03962_),
    .A1(_03959_),
    .A2(_03960_));
 sg13g2_nor2_1 _11023_ (.A(_03961_),
    .B(_03962_),
    .Y(_00230_));
 sg13g2_a21oi_1 _11024_ (.A1(net2207),
    .A2(_01846_),
    .Y(_03963_),
    .B1(_03961_));
 sg13g2_nor2_1 _11025_ (.A(\vgadonut.donut.donuthit.t[5] ),
    .B(_01842_),
    .Y(_03964_));
 sg13g2_xnor2_1 _11026_ (.Y(_03965_),
    .A(\vgadonut.donut.donuthit.t[5] ),
    .B(_01842_));
 sg13g2_o21ai_1 _11027_ (.B1(net1678),
    .Y(_03966_),
    .A1(_03963_),
    .A2(_03965_));
 sg13g2_a21oi_1 _11028_ (.A1(_03963_),
    .A2(_03965_),
    .Y(_00231_),
    .B1(_03966_));
 sg13g2_xnor2_1 _11029_ (.Y(_03967_),
    .A(net2295),
    .B(_01828_));
 sg13g2_a221oi_1 _11030_ (.B2(\vgadonut.donut.donuthit.t[4] ),
    .C1(_03961_),
    .B1(_01846_),
    .A1(\vgadonut.donut.donuthit.t[5] ),
    .Y(_03968_),
    .A2(_01842_));
 sg13g2_o21ai_1 _11031_ (.B1(_03967_),
    .Y(_03969_),
    .A1(_03964_),
    .A2(_03968_));
 sg13g2_nor3_1 _11032_ (.A(_03964_),
    .B(_03967_),
    .C(_03968_),
    .Y(_03970_));
 sg13g2_or2_1 _11033_ (.X(_03971_),
    .B(_03970_),
    .A(net1699));
 sg13g2_nor2b_1 _11034_ (.A(_03971_),
    .B_N(net2296),
    .Y(_00232_));
 sg13g2_a21o_1 _11035_ (.A2(_01828_),
    .A1(net2295),
    .B1(_03970_),
    .X(_03972_));
 sg13g2_nand2_1 _11036_ (.Y(_03973_),
    .A(\vgadonut.donut.donuthit.t[7] ),
    .B(_01836_));
 sg13g2_xnor2_1 _11037_ (.Y(_03974_),
    .A(net2314),
    .B(_01835_));
 sg13g2_nand2_1 _11038_ (.Y(_03975_),
    .A(_03972_),
    .B(_03974_));
 sg13g2_o21ai_1 _11039_ (.B1(net1678),
    .Y(_03976_),
    .A1(_03972_),
    .A2(_03974_));
 sg13g2_nor2b_1 _11040_ (.A(_03976_),
    .B_N(_03975_),
    .Y(_00233_));
 sg13g2_nand2_1 _11041_ (.Y(_03977_),
    .A(net2257),
    .B(_01822_));
 sg13g2_xnor2_1 _11042_ (.Y(_03978_),
    .A(net2257),
    .B(_01822_));
 sg13g2_and2_1 _11043_ (.A(_03973_),
    .B(_03975_),
    .X(_03979_));
 sg13g2_o21ai_1 _11044_ (.B1(net1679),
    .Y(_03980_),
    .A1(_03978_),
    .A2(_03979_));
 sg13g2_a21oi_1 _11045_ (.A1(_03978_),
    .A2(_03979_),
    .Y(_00234_),
    .B1(_03980_));
 sg13g2_o21ai_1 _11046_ (.B1(_03977_),
    .Y(_03981_),
    .A1(_03978_),
    .A2(_03979_));
 sg13g2_nor2_1 _11047_ (.A(_00642_),
    .B(_01814_),
    .Y(_03982_));
 sg13g2_xnor2_1 _11048_ (.Y(_03983_),
    .A(_00642_),
    .B(_01814_));
 sg13g2_inv_1 _11049_ (.Y(_03984_),
    .A(_03983_));
 sg13g2_xnor2_1 _11050_ (.Y(_03985_),
    .A(_03981_),
    .B(_03984_));
 sg13g2_nand2_1 _11051_ (.Y(_00235_),
    .A(net1678),
    .B(_03985_));
 sg13g2_a21oi_1 _11052_ (.A1(_03981_),
    .A2(_03984_),
    .Y(_03986_),
    .B1(_03982_));
 sg13g2_nand3_1 _11053_ (.B(net1544),
    .C(net1541),
    .A(net2300),
    .Y(_03987_));
 sg13g2_xor2_1 _11054_ (.B(net1539),
    .A(net2300),
    .X(_03988_));
 sg13g2_o21ai_1 _11055_ (.B1(net1678),
    .Y(_03989_),
    .A1(_03986_),
    .A2(_03988_));
 sg13g2_a21oi_1 _11056_ (.A1(_03986_),
    .A2(_03988_),
    .Y(_00236_),
    .B1(_03989_));
 sg13g2_o21ai_1 _11057_ (.B1(_03987_),
    .Y(_03990_),
    .A1(_03986_),
    .A2(_03988_));
 sg13g2_mux2_1 _11058_ (.A0(_01700_),
    .A1(_01701_),
    .S(net1578),
    .X(_03991_));
 sg13g2_xnor2_1 _11059_ (.Y(_03992_),
    .A(net1595),
    .B(_03991_));
 sg13g2_a21oi_2 _11060_ (.B1(_03992_),
    .Y(_03993_),
    .A2(_01706_),
    .A1(_01704_));
 sg13g2_nand3_1 _11061_ (.B(_01706_),
    .C(_03992_),
    .A(_01704_),
    .Y(_03994_));
 sg13g2_nor2b_2 _11062_ (.A(_03993_),
    .B_N(_03994_),
    .Y(_03995_));
 sg13g2_nor2_1 _11063_ (.A(_01694_),
    .B(_03995_),
    .Y(_03996_));
 sg13g2_xor2_1 _11064_ (.B(_03995_),
    .A(_01694_),
    .X(_03997_));
 sg13g2_nor2_1 _11065_ (.A(_01710_),
    .B(_03997_),
    .Y(_03998_));
 sg13g2_xor2_1 _11066_ (.B(_03997_),
    .A(_01710_),
    .X(_03999_));
 sg13g2_nor2_1 _11067_ (.A(_01712_),
    .B(net1545),
    .Y(_04000_));
 sg13g2_nor2b_1 _11068_ (.A(_04000_),
    .B_N(_03999_),
    .Y(_04001_));
 sg13g2_xnor2_1 _11069_ (.Y(_04002_),
    .A(_03999_),
    .B(_04000_));
 sg13g2_and2_1 _11070_ (.A(\vgadonut.donut.donuthit.t[11] ),
    .B(_04002_),
    .X(_04003_));
 sg13g2_xor2_1 _11071_ (.B(_04002_),
    .A(net2328),
    .X(_04004_));
 sg13g2_xnor2_1 _11072_ (.Y(_04005_),
    .A(_03990_),
    .B(_04004_));
 sg13g2_nor2_1 _11073_ (.A(net1699),
    .B(_04005_),
    .Y(_00237_));
 sg13g2_a21oi_1 _11074_ (.A1(_03990_),
    .A2(_04004_),
    .Y(_04006_),
    .B1(_04003_));
 sg13g2_nor3_1 _11075_ (.A(net1579),
    .B(_01523_),
    .C(_01525_),
    .Y(_04007_));
 sg13g2_a21oi_1 _11076_ (.A1(net1578),
    .A2(_01506_),
    .Y(_04008_),
    .B1(_04007_));
 sg13g2_xnor2_1 _11077_ (.Y(_04009_),
    .A(net1594),
    .B(_04008_));
 sg13g2_xor2_1 _11078_ (.B(_04009_),
    .A(_03993_),
    .X(_04010_));
 sg13g2_inv_1 _11079_ (.Y(_04011_),
    .A(_04010_));
 sg13g2_nand2b_1 _11080_ (.Y(_04012_),
    .B(_04010_),
    .A_N(_01707_));
 sg13g2_xor2_1 _11081_ (.B(_04010_),
    .A(_01707_),
    .X(_04013_));
 sg13g2_nor2b_1 _11082_ (.A(_03996_),
    .B_N(_04013_),
    .Y(_04014_));
 sg13g2_xor2_1 _11083_ (.B(_04013_),
    .A(_03996_),
    .X(_04015_));
 sg13g2_nor2_1 _11084_ (.A(_03998_),
    .B(_04001_),
    .Y(_04016_));
 sg13g2_nor2_1 _11085_ (.A(_04015_),
    .B(_04016_),
    .Y(_04017_));
 sg13g2_xnor2_1 _11086_ (.Y(_04018_),
    .A(_04015_),
    .B(_04016_));
 sg13g2_xnor2_1 _11087_ (.Y(_04019_),
    .A(\vgadonut.donut.donuthit.t[12] ),
    .B(_04018_));
 sg13g2_nand2b_1 _11088_ (.Y(_04020_),
    .B(_04019_),
    .A_N(_04006_));
 sg13g2_xnor2_1 _11089_ (.Y(_04021_),
    .A(_04006_),
    .B(_04019_));
 sg13g2_and2_1 _11090_ (.A(net1678),
    .B(_04021_),
    .X(_00238_));
 sg13g2_o21ai_1 _11091_ (.B1(_04020_),
    .Y(_04022_),
    .A1(_00643_),
    .A2(_04018_));
 sg13g2_nor2_1 _11092_ (.A(_04014_),
    .B(_04017_),
    .Y(_04023_));
 sg13g2_nor2_1 _11093_ (.A(_03995_),
    .B(_04011_),
    .Y(_04024_));
 sg13g2_mux2_1 _11094_ (.A0(_04011_),
    .A1(_04009_),
    .S(_03995_),
    .X(_04025_));
 sg13g2_inv_1 _11095_ (.Y(_04026_),
    .A(_04025_));
 sg13g2_xnor2_1 _11096_ (.Y(_04027_),
    .A(_04012_),
    .B(_04025_));
 sg13g2_nor2b_1 _11097_ (.A(_04023_),
    .B_N(_04027_),
    .Y(_04028_));
 sg13g2_xnor2_1 _11098_ (.Y(_04029_),
    .A(_04023_),
    .B(_04027_));
 sg13g2_and2_1 _11099_ (.A(\vgadonut.donut.donuthit.t[13] ),
    .B(_04029_),
    .X(_04030_));
 sg13g2_xor2_1 _11100_ (.B(_04029_),
    .A(net2315),
    .X(_04031_));
 sg13g2_xnor2_1 _11101_ (.Y(_04032_),
    .A(_04022_),
    .B(_04031_));
 sg13g2_nor2_1 _11102_ (.A(net1699),
    .B(net2316),
    .Y(_00239_));
 sg13g2_a21oi_1 _11103_ (.A1(_04022_),
    .A2(_04031_),
    .Y(_04033_),
    .B1(_04030_));
 sg13g2_a21oi_1 _11104_ (.A1(_04012_),
    .A2(_04026_),
    .Y(_04034_),
    .B1(_04028_));
 sg13g2_xor2_1 _11105_ (.B(_04034_),
    .A(_04024_),
    .X(_04035_));
 sg13g2_xnor2_1 _11106_ (.Y(_04036_),
    .A(net2346),
    .B(_04035_));
 sg13g2_nand2b_1 _11107_ (.Y(_04037_),
    .B(_04036_),
    .A_N(_04033_));
 sg13g2_xor2_1 _11108_ (.B(_04036_),
    .A(_04033_),
    .X(_04038_));
 sg13g2_nor2_1 _11109_ (.A(net1699),
    .B(_04038_),
    .Y(_00240_));
 sg13g2_o21ai_1 _11110_ (.B1(_04037_),
    .Y(_04039_),
    .A1(_00644_),
    .A2(_04035_));
 sg13g2_a21o_1 _11111_ (.A2(_04034_),
    .A1(_04024_),
    .B1(_04011_),
    .X(_04040_));
 sg13g2_xor2_1 _11112_ (.B(_04040_),
    .A(net2323),
    .X(_04041_));
 sg13g2_nor2b_1 _11113_ (.A(_04039_),
    .B_N(_04041_),
    .Y(_04042_));
 sg13g2_xnor2_1 _11114_ (.Y(_04043_),
    .A(_04039_),
    .B(_04041_));
 sg13g2_nor2_1 _11115_ (.A(net1699),
    .B(_04043_),
    .Y(_00241_));
 sg13g2_nor2_1 _11116_ (.A(net1642),
    .B(_00742_),
    .Y(_00242_));
 sg13g2_and2_1 _11117_ (.A(net1958),
    .B(net1761),
    .X(_04044_));
 sg13g2_nand2_2 _11118_ (.Y(_04045_),
    .A(net1959),
    .B(net1762));
 sg13g2_nand2_1 _11119_ (.Y(_04046_),
    .A(net1969),
    .B(net1749));
 sg13g2_nand2_1 _11120_ (.Y(_04047_),
    .A(\vgadonut.donut.ysA[3] ),
    .B(net1850));
 sg13g2_xnor2_1 _11121_ (.Y(_04048_),
    .A(\vgadonut.donut.ysA[3] ),
    .B(net1850));
 sg13g2_nand2_1 _11122_ (.Y(_04049_),
    .A(net2363),
    .B(net1852));
 sg13g2_nand2_1 _11123_ (.Y(_04050_),
    .A(\vgadonut.donut.ysA[1] ),
    .B(net1853));
 sg13g2_nand2_1 _11124_ (.Y(_04051_),
    .A(net2018),
    .B(net1854));
 sg13g2_xnor2_1 _11125_ (.Y(_04052_),
    .A(\vgadonut.donut.ysA[1] ),
    .B(net1853));
 sg13g2_o21ai_1 _11126_ (.B1(_04050_),
    .Y(_04053_),
    .A1(_04051_),
    .A2(_04052_));
 sg13g2_xnor2_1 _11127_ (.Y(_04054_),
    .A(net2363),
    .B(net1852));
 sg13g2_nand2b_1 _11128_ (.Y(_04055_),
    .B(_04053_),
    .A_N(_04054_));
 sg13g2_a21o_1 _11129_ (.A2(_04055_),
    .A1(_04049_),
    .B1(_04048_),
    .X(_04056_));
 sg13g2_xnor2_1 _11130_ (.Y(_04057_),
    .A(\vgadonut.donut.ysA[4] ),
    .B(net1849));
 sg13g2_a21oi_1 _11131_ (.A1(_04047_),
    .A2(_04056_),
    .Y(_04058_),
    .B1(_04057_));
 sg13g2_nand3_1 _11132_ (.B(_04056_),
    .C(_04057_),
    .A(_04047_),
    .Y(_04059_));
 sg13g2_nand2b_1 _11133_ (.Y(_04060_),
    .B(_04059_),
    .A_N(_04058_));
 sg13g2_nand2_2 _11134_ (.Y(_04061_),
    .A(net1765),
    .B(net1710));
 sg13g2_nand2_1 _11135_ (.Y(_04062_),
    .A(net1854),
    .B(net1712));
 sg13g2_a22oi_1 _11136_ (.Y(_04063_),
    .B1(_04061_),
    .B2(_04062_),
    .A2(_04060_),
    .A1(net1767));
 sg13g2_nor2_1 _11137_ (.A(net1776),
    .B(net1704),
    .Y(_04064_));
 sg13g2_a21o_1 _11138_ (.A2(net1703),
    .A1(net2097),
    .B1(_04063_),
    .X(_00243_));
 sg13g2_a21o_1 _11139_ (.A2(net1849),
    .A1(\vgadonut.donut.ysA[4] ),
    .B1(_04058_),
    .X(_04065_));
 sg13g2_nand2_1 _11140_ (.Y(_04066_),
    .A(\vgadonut.donut.ysA[5] ),
    .B(net1846));
 sg13g2_xor2_1 _11141_ (.B(net1846),
    .A(\vgadonut.donut.ysA[5] ),
    .X(_04067_));
 sg13g2_o21ai_1 _11142_ (.B1(net1767),
    .Y(_04068_),
    .A1(_04065_),
    .A2(_04067_));
 sg13g2_a21o_1 _11143_ (.A2(_04067_),
    .A1(_04065_),
    .B1(_04068_),
    .X(_04069_));
 sg13g2_a21oi_1 _11144_ (.A1(net1853),
    .A2(net1774),
    .Y(_04070_),
    .B1(net1707));
 sg13g2_a22oi_1 _11145_ (.Y(_00244_),
    .B1(_04069_),
    .B2(_04070_),
    .A2(net1706),
    .A1(_06854_));
 sg13g2_xnor2_1 _11146_ (.Y(_04071_),
    .A(\vgadonut.donut.ysA[6] ),
    .B(net1844));
 sg13g2_o21ai_1 _11147_ (.B1(_04065_),
    .Y(_04072_),
    .A1(\vgadonut.donut.ysA[5] ),
    .A2(net1846));
 sg13g2_a21oi_1 _11148_ (.A1(_04066_),
    .A2(_04072_),
    .Y(_04073_),
    .B1(_04071_));
 sg13g2_nand3_1 _11149_ (.B(_04071_),
    .C(_04072_),
    .A(_04066_),
    .Y(_04074_));
 sg13g2_nand2b_1 _11150_ (.Y(_04075_),
    .B(_04074_),
    .A_N(_04073_));
 sg13g2_o21ai_1 _11151_ (.B1(net1712),
    .Y(_04076_),
    .A1(net1852),
    .A2(net1767));
 sg13g2_a21oi_1 _11152_ (.A1(net1767),
    .A2(_04075_),
    .Y(_04077_),
    .B1(_04076_));
 sg13g2_a21o_1 _11153_ (.A2(net1702),
    .A1(net2167),
    .B1(_04077_),
    .X(_00245_));
 sg13g2_a21oi_1 _11154_ (.A1(\vgadonut.donut.ysA[6] ),
    .A2(net1844),
    .Y(_04078_),
    .B1(_04073_));
 sg13g2_xnor2_1 _11155_ (.Y(_04079_),
    .A(\vgadonut.donut.ysA[7] ),
    .B(net1842));
 sg13g2_nor2_1 _11156_ (.A(_04078_),
    .B(_04079_),
    .Y(_04080_));
 sg13g2_xnor2_1 _11157_ (.Y(_04081_),
    .A(_04078_),
    .B(_04079_));
 sg13g2_o21ai_1 _11158_ (.B1(net1714),
    .Y(_04082_),
    .A1(net1851),
    .A2(net1767));
 sg13g2_a21oi_1 _11159_ (.A1(net1767),
    .A2(_04081_),
    .Y(_04083_),
    .B1(_04082_));
 sg13g2_a21o_1 _11160_ (.A2(net1702),
    .A1(net2172),
    .B1(_04083_),
    .X(_00246_));
 sg13g2_xnor2_1 _11161_ (.Y(_04084_),
    .A(\vgadonut.donut.ysA[8] ),
    .B(net1840));
 sg13g2_a21oi_1 _11162_ (.A1(\vgadonut.donut.ysA[7] ),
    .A2(net1842),
    .Y(_04085_),
    .B1(_04080_));
 sg13g2_or2_1 _11163_ (.X(_04086_),
    .B(_04085_),
    .A(_04084_));
 sg13g2_a21oi_1 _11164_ (.A1(_04084_),
    .A2(_04085_),
    .Y(_04087_),
    .B1(net1760));
 sg13g2_nand2b_1 _11165_ (.Y(_04088_),
    .B(net1854),
    .A_N(net1848));
 sg13g2_xor2_1 _11166_ (.B(net1854),
    .A(net1848),
    .X(_04089_));
 sg13g2_a221oi_1 _11167_ (.B2(net1774),
    .C1(net1709),
    .B1(_04089_),
    .A1(_04086_),
    .Y(_04090_),
    .A2(_04087_));
 sg13g2_a21oi_1 _11168_ (.A1(_06861_),
    .A2(net1704),
    .Y(_00247_),
    .B1(_04090_));
 sg13g2_o21ai_1 _11169_ (.B1(_04086_),
    .Y(_04091_),
    .A1(_06861_),
    .A2(_00596_));
 sg13g2_nor2_1 _11170_ (.A(\vgadonut.donut.ysA[9] ),
    .B(net1837),
    .Y(_04092_));
 sg13g2_xnor2_1 _11171_ (.Y(_04093_),
    .A(\vgadonut.donut.ysA[9] ),
    .B(net1837));
 sg13g2_xnor2_1 _11172_ (.Y(_04094_),
    .A(_04091_),
    .B(_04093_));
 sg13g2_nor2_1 _11173_ (.A(net1853),
    .B(_00594_),
    .Y(_04095_));
 sg13g2_xnor2_1 _11174_ (.Y(_04096_),
    .A(net1853),
    .B(net1847));
 sg13g2_xnor2_1 _11175_ (.Y(_04097_),
    .A(_04088_),
    .B(_04096_));
 sg13g2_o21ai_1 _11176_ (.B1(net1714),
    .Y(_04098_),
    .A1(net1768),
    .A2(_04097_));
 sg13g2_a21oi_1 _11177_ (.A1(net1768),
    .A2(_04094_),
    .Y(_04099_),
    .B1(_04098_));
 sg13g2_a21oi_1 _11178_ (.A1(_06863_),
    .A2(net1704),
    .Y(_00248_),
    .B1(_04099_));
 sg13g2_xnor2_1 _11179_ (.Y(_04100_),
    .A(\vgadonut.donut.ysA[10] ),
    .B(net1834));
 sg13g2_a21oi_1 _11180_ (.A1(\vgadonut.donut.ysA[9] ),
    .A2(net1837),
    .Y(_04101_),
    .B1(_04091_));
 sg13g2_nor3_1 _11181_ (.A(_04092_),
    .B(_04100_),
    .C(_04101_),
    .Y(_04102_));
 sg13g2_o21ai_1 _11182_ (.B1(_04100_),
    .Y(_04103_),
    .A1(_04092_),
    .A2(_04101_));
 sg13g2_nand2_1 _11183_ (.Y(_04104_),
    .A(net1768),
    .B(_04103_));
 sg13g2_nand2b_1 _11184_ (.Y(_04105_),
    .B(net1845),
    .A_N(\vgadonut.donut.sA[4] ));
 sg13g2_xor2_1 _11185_ (.B(net1845),
    .A(net1852),
    .X(_04106_));
 sg13g2_a21oi_1 _11186_ (.A1(_04088_),
    .A2(_04096_),
    .Y(_04107_),
    .B1(_04095_));
 sg13g2_or2_1 _11187_ (.X(_04108_),
    .B(_04107_),
    .A(_04106_));
 sg13g2_a21oi_1 _11188_ (.A1(_04106_),
    .A2(_04107_),
    .Y(_04109_),
    .B1(net1772));
 sg13g2_a21oi_1 _11189_ (.A1(_04108_),
    .A2(_04109_),
    .Y(_04110_),
    .B1(net1709));
 sg13g2_o21ai_1 _11190_ (.B1(_04110_),
    .Y(_04111_),
    .A1(_04102_),
    .A2(_04104_));
 sg13g2_o21ai_1 _11191_ (.B1(_04111_),
    .Y(_04112_),
    .A1(net2283),
    .A2(net1714));
 sg13g2_inv_1 _11192_ (.Y(_00249_),
    .A(_04112_));
 sg13g2_a21o_1 _11193_ (.A2(net1834),
    .A1(\vgadonut.donut.ysA[10] ),
    .B1(_04102_),
    .X(_04113_));
 sg13g2_nor2_1 _11194_ (.A(\vgadonut.donut.ysA[11] ),
    .B(net1832),
    .Y(_04114_));
 sg13g2_xnor2_1 _11195_ (.Y(_04115_),
    .A(\vgadonut.donut.ysA[11] ),
    .B(net1832));
 sg13g2_xnor2_1 _11196_ (.Y(_04116_),
    .A(_04113_),
    .B(_04115_));
 sg13g2_nand2b_1 _11197_ (.Y(_04117_),
    .B(net1843),
    .A_N(net1851));
 sg13g2_xor2_1 _11198_ (.B(net1843),
    .A(net1850),
    .X(_04118_));
 sg13g2_a21o_1 _11199_ (.A2(_04108_),
    .A1(_04105_),
    .B1(_04118_),
    .X(_04119_));
 sg13g2_nand3_1 _11200_ (.B(_04108_),
    .C(_04118_),
    .A(_04105_),
    .Y(_04120_));
 sg13g2_and2_1 _11201_ (.A(net1777),
    .B(_04120_),
    .X(_04121_));
 sg13g2_a221oi_1 _11202_ (.B2(_04121_),
    .C1(net1709),
    .B1(_04119_),
    .A1(net1772),
    .Y(_04122_),
    .A2(_04116_));
 sg13g2_a21oi_1 _11203_ (.A1(_06866_),
    .A2(net1704),
    .Y(_00250_),
    .B1(_04122_));
 sg13g2_xnor2_1 _11204_ (.Y(_04123_),
    .A(\vgadonut.donut.ysA[12] ),
    .B(net1831));
 sg13g2_a21oi_1 _11205_ (.A1(\vgadonut.donut.ysA[11] ),
    .A2(net1832),
    .Y(_04124_),
    .B1(_04113_));
 sg13g2_o21ai_1 _11206_ (.B1(_04123_),
    .Y(_04125_),
    .A1(_04114_),
    .A2(_04124_));
 sg13g2_nor3_1 _11207_ (.A(_04114_),
    .B(_04123_),
    .C(_04124_),
    .Y(_04126_));
 sg13g2_nand2_1 _11208_ (.Y(_04127_),
    .A(net1772),
    .B(_04125_));
 sg13g2_nand2b_1 _11209_ (.Y(_04128_),
    .B(net1840),
    .A_N(net1848));
 sg13g2_xor2_1 _11210_ (.B(net1840),
    .A(net1848),
    .X(_04129_));
 sg13g2_a21o_1 _11211_ (.A2(_04119_),
    .A1(_04117_),
    .B1(_04129_),
    .X(_04130_));
 sg13g2_nand3_1 _11212_ (.B(_04119_),
    .C(_04129_),
    .A(_04117_),
    .Y(_04131_));
 sg13g2_nand3_1 _11213_ (.B(_04130_),
    .C(_04131_),
    .A(net1776),
    .Y(_04132_));
 sg13g2_and2_1 _11214_ (.A(net1714),
    .B(_04132_),
    .X(_04133_));
 sg13g2_o21ai_1 _11215_ (.B1(_04133_),
    .Y(_04134_),
    .A1(_04126_),
    .A2(_04127_));
 sg13g2_o21ai_1 _11216_ (.B1(_04134_),
    .Y(_04135_),
    .A1(net2280),
    .A2(net1714));
 sg13g2_inv_1 _11217_ (.Y(_00251_),
    .A(_04135_));
 sg13g2_xor2_1 _11218_ (.B(net1826),
    .A(\vgadonut.donut.ysA[13] ),
    .X(_04136_));
 sg13g2_a21o_1 _11219_ (.A2(net1831),
    .A1(\vgadonut.donut.ysA[12] ),
    .B1(_04126_),
    .X(_04137_));
 sg13g2_xnor2_1 _11220_ (.Y(_04138_),
    .A(_04136_),
    .B(_04137_));
 sg13g2_nor2_1 _11221_ (.A(_00594_),
    .B(net1837),
    .Y(_04139_));
 sg13g2_nor2b_1 _11222_ (.A(net1847),
    .B_N(net1837),
    .Y(_04140_));
 sg13g2_or2_1 _11223_ (.X(_04141_),
    .B(_04140_),
    .A(_04139_));
 sg13g2_and2_1 _11224_ (.A(_04128_),
    .B(_04130_),
    .X(_04142_));
 sg13g2_or2_1 _11225_ (.X(_04143_),
    .B(_04142_),
    .A(_04141_));
 sg13g2_a21oi_1 _11226_ (.A1(_04141_),
    .A2(_04142_),
    .Y(_04144_),
    .B1(net1772));
 sg13g2_a21oi_1 _11227_ (.A1(_04143_),
    .A2(_04144_),
    .Y(_04145_),
    .B1(_04045_));
 sg13g2_o21ai_1 _11228_ (.B1(_04145_),
    .Y(_04146_),
    .A1(_03927_),
    .A2(_04138_));
 sg13g2_o21ai_1 _11229_ (.B1(_04146_),
    .Y(_04147_),
    .A1(net2239),
    .A2(net1715));
 sg13g2_inv_1 _11230_ (.Y(_00252_),
    .A(_04147_));
 sg13g2_xnor2_1 _11231_ (.Y(_04148_),
    .A(\vgadonut.donut.ysA[14] ),
    .B(net1827));
 sg13g2_o21ai_1 _11232_ (.B1(_04137_),
    .Y(_04149_),
    .A1(\vgadonut.donut.ysA[13] ),
    .A2(net1826));
 sg13g2_o21ai_1 _11233_ (.B1(_04149_),
    .Y(_04150_),
    .A1(_06870_),
    .A2(net1797));
 sg13g2_nand2b_1 _11234_ (.Y(_04151_),
    .B(_04150_),
    .A_N(_04148_));
 sg13g2_xor2_1 _11235_ (.B(_04150_),
    .A(_04148_),
    .X(_04152_));
 sg13g2_nor2_1 _11236_ (.A(_03927_),
    .B(_04152_),
    .Y(_04153_));
 sg13g2_nand2b_1 _11237_ (.Y(_04154_),
    .B(net1835),
    .A_N(net1845));
 sg13g2_xor2_1 _11238_ (.B(net1835),
    .A(net1845),
    .X(_04155_));
 sg13g2_nor2_1 _11239_ (.A(_04139_),
    .B(_04142_),
    .Y(_04156_));
 sg13g2_nor2_1 _11240_ (.A(_04140_),
    .B(_04156_),
    .Y(_04157_));
 sg13g2_nor2_1 _11241_ (.A(_04155_),
    .B(_04157_),
    .Y(_04158_));
 sg13g2_and2_1 _11242_ (.A(_04155_),
    .B(_04157_),
    .X(_04159_));
 sg13g2_nor3_1 _11243_ (.A(net1772),
    .B(_04158_),
    .C(_04159_),
    .Y(_04160_));
 sg13g2_nor3_1 _11244_ (.A(net1709),
    .B(_04153_),
    .C(_04160_),
    .Y(_04161_));
 sg13g2_a21oi_1 _11245_ (.A1(_06871_),
    .A2(net1705),
    .Y(_00253_),
    .B1(_04161_));
 sg13g2_nand2_1 _11246_ (.Y(_04162_),
    .A(\vgadonut.donut.ysA[15] ),
    .B(net1827));
 sg13g2_xor2_1 _11247_ (.B(net1827),
    .A(\vgadonut.donut.ysA[15] ),
    .X(_04163_));
 sg13g2_o21ai_1 _11248_ (.B1(_04151_),
    .Y(_04164_),
    .A1(_06871_),
    .A2(net1798));
 sg13g2_o21ai_1 _11249_ (.B1(net1772),
    .Y(_04165_),
    .A1(_04163_),
    .A2(_04164_));
 sg13g2_a21oi_1 _11250_ (.A1(_04163_),
    .A2(_04164_),
    .Y(_04166_),
    .B1(_04165_));
 sg13g2_nor2_1 _11251_ (.A(net1842),
    .B(_00597_),
    .Y(_04167_));
 sg13g2_xnor2_1 _11252_ (.Y(_04168_),
    .A(net1843),
    .B(net1832));
 sg13g2_o21ai_1 _11253_ (.B1(_04154_),
    .Y(_04169_),
    .A1(_04155_),
    .A2(_04157_));
 sg13g2_and2_1 _11254_ (.A(_04168_),
    .B(_04169_),
    .X(_04170_));
 sg13g2_o21ai_1 _11255_ (.B1(net1776),
    .Y(_04171_),
    .A1(_04168_),
    .A2(_04169_));
 sg13g2_o21ai_1 _11256_ (.B1(net1715),
    .Y(_04172_),
    .A1(_04170_),
    .A2(_04171_));
 sg13g2_nor2_1 _11257_ (.A(_04166_),
    .B(_04172_),
    .Y(_04173_));
 sg13g2_a21oi_1 _11258_ (.A1(_06874_),
    .A2(net1705),
    .Y(_00254_),
    .B1(_04173_));
 sg13g2_nor2_1 _11259_ (.A(net2201),
    .B(net1715),
    .Y(_04174_));
 sg13g2_nand2_1 _11260_ (.Y(_04175_),
    .A(\vgadonut.donut.ysA[16] ),
    .B(net1828));
 sg13g2_xnor2_1 _11261_ (.Y(_04176_),
    .A(\vgadonut.donut.ysA[16] ),
    .B(net1827));
 sg13g2_o21ai_1 _11262_ (.B1(_04164_),
    .Y(_04177_),
    .A1(\vgadonut.donut.ysA[15] ),
    .A2(net1827));
 sg13g2_a21o_1 _11263_ (.A2(_04177_),
    .A1(_04162_),
    .B1(_04176_),
    .X(_04178_));
 sg13g2_nand3_1 _11264_ (.B(_04176_),
    .C(_04177_),
    .A(_04162_),
    .Y(_04179_));
 sg13g2_nand3_1 _11265_ (.B(_04178_),
    .C(_04179_),
    .A(net1772),
    .Y(_04180_));
 sg13g2_xnor2_1 _11266_ (.Y(_04181_),
    .A(net1841),
    .B(net1831));
 sg13g2_o21ai_1 _11267_ (.B1(_04181_),
    .Y(_04182_),
    .A1(_04167_),
    .A2(_04170_));
 sg13g2_or3_1 _11268_ (.A(_04167_),
    .B(_04170_),
    .C(_04181_),
    .X(_04183_));
 sg13g2_and2_1 _11269_ (.A(net1776),
    .B(_04183_),
    .X(_04184_));
 sg13g2_a21oi_1 _11270_ (.A1(_04182_),
    .A2(_04184_),
    .Y(_04185_),
    .B1(net1709));
 sg13g2_a21oi_1 _11271_ (.A1(_04180_),
    .A2(_04185_),
    .Y(_00255_),
    .B1(_04174_));
 sg13g2_xnor2_1 _11272_ (.Y(_04186_),
    .A(\vgadonut.donut.ysA[17] ),
    .B(net1828));
 sg13g2_nand3_1 _11273_ (.B(_04178_),
    .C(_04186_),
    .A(_04175_),
    .Y(_04187_));
 sg13g2_a21o_1 _11274_ (.A2(_04178_),
    .A1(_04175_),
    .B1(_04186_),
    .X(_04188_));
 sg13g2_nand3_1 _11275_ (.B(_04187_),
    .C(_04188_),
    .A(net1771),
    .Y(_04189_));
 sg13g2_nand2_1 _11276_ (.Y(_04190_),
    .A(net1838),
    .B(net1798));
 sg13g2_nor2_1 _11277_ (.A(net1837),
    .B(net1798),
    .Y(_04191_));
 sg13g2_xnor2_1 _11278_ (.Y(_04192_),
    .A(net1838),
    .B(net1828));
 sg13g2_o21ai_1 _11279_ (.B1(_04182_),
    .Y(_04193_),
    .A1(net1841),
    .A2(_00598_));
 sg13g2_a21oi_1 _11280_ (.A1(_04192_),
    .A2(_04193_),
    .Y(_04194_),
    .B1(net1771));
 sg13g2_o21ai_1 _11281_ (.B1(_04194_),
    .Y(_04195_),
    .A1(_04192_),
    .A2(_04193_));
 sg13g2_nand3_1 _11282_ (.B(_04189_),
    .C(_04195_),
    .A(net1715),
    .Y(_04196_));
 sg13g2_o21ai_1 _11283_ (.B1(_04196_),
    .Y(_04197_),
    .A1(net2216),
    .A2(net1714));
 sg13g2_inv_1 _11284_ (.Y(_00256_),
    .A(_04197_));
 sg13g2_and2_1 _11285_ (.A(\vgadonut.donut.ysA[18] ),
    .B(net1828),
    .X(_04198_));
 sg13g2_xor2_1 _11286_ (.B(net1828),
    .A(\vgadonut.donut.ysA[18] ),
    .X(_04199_));
 sg13g2_o21ai_1 _11287_ (.B1(net1830),
    .Y(_04200_),
    .A1(\vgadonut.donut.ysA[16] ),
    .A2(\vgadonut.donut.ysA[17] ));
 sg13g2_nor2_1 _11288_ (.A(_04178_),
    .B(_04186_),
    .Y(_04201_));
 sg13g2_o21ai_1 _11289_ (.B1(_04200_),
    .Y(_04202_),
    .A1(_04178_),
    .A2(_04186_));
 sg13g2_xnor2_1 _11290_ (.Y(_04203_),
    .A(_04199_),
    .B(_04202_));
 sg13g2_xor2_1 _11291_ (.B(net1828),
    .A(net1834),
    .X(_04204_));
 sg13g2_a21oi_1 _11292_ (.A1(_04190_),
    .A2(_04193_),
    .Y(_04205_),
    .B1(_04191_));
 sg13g2_or2_1 _11293_ (.X(_04206_),
    .B(_04205_),
    .A(_04204_));
 sg13g2_a21oi_1 _11294_ (.A1(_04204_),
    .A2(_04205_),
    .Y(_04207_),
    .B1(net1771));
 sg13g2_a21oi_1 _11295_ (.A1(_04206_),
    .A2(_04207_),
    .Y(_04208_),
    .B1(net1709));
 sg13g2_o21ai_1 _11296_ (.B1(_04208_),
    .Y(_04209_),
    .A1(net1760),
    .A2(_04203_));
 sg13g2_o21ai_1 _11297_ (.B1(_04209_),
    .Y(_04210_),
    .A1(net2260),
    .A2(net1714));
 sg13g2_inv_1 _11298_ (.Y(_00257_),
    .A(_04210_));
 sg13g2_xor2_1 _11299_ (.B(net1828),
    .A(\vgadonut.donut.ysA[19] ),
    .X(_04211_));
 sg13g2_a21o_1 _11300_ (.A2(_04202_),
    .A1(_04199_),
    .B1(_04198_),
    .X(_04212_));
 sg13g2_o21ai_1 _11301_ (.B1(net1771),
    .Y(_04213_),
    .A1(_04211_),
    .A2(_04212_));
 sg13g2_a21oi_1 _11302_ (.A1(_04211_),
    .A2(_04212_),
    .Y(_04214_),
    .B1(_04213_));
 sg13g2_xnor2_1 _11303_ (.Y(_04215_),
    .A(net1832),
    .B(net1829));
 sg13g2_o21ai_1 _11304_ (.B1(_04206_),
    .Y(_04216_),
    .A1(net1834),
    .A2(net1798));
 sg13g2_o21ai_1 _11305_ (.B1(net1776),
    .Y(_04217_),
    .A1(_04215_),
    .A2(_04216_));
 sg13g2_a21oi_1 _11306_ (.A1(_04215_),
    .A2(_04216_),
    .Y(_04218_),
    .B1(_04217_));
 sg13g2_nor3_1 _11307_ (.A(net1704),
    .B(_04214_),
    .C(_04218_),
    .Y(_04219_));
 sg13g2_a21oi_1 _11308_ (.A1(_06879_),
    .A2(net1704),
    .Y(_00258_),
    .B1(_04219_));
 sg13g2_xnor2_1 _11309_ (.Y(_04220_),
    .A(\vgadonut.donut.ysA[20] ),
    .B(net1830));
 sg13g2_nand3_1 _11310_ (.B(_04201_),
    .C(_04211_),
    .A(_04199_),
    .Y(_04221_));
 sg13g2_o21ai_1 _11311_ (.B1(net1830),
    .Y(_04222_),
    .A1(\vgadonut.donut.ysA[18] ),
    .A2(\vgadonut.donut.ysA[19] ));
 sg13g2_nand3_1 _11312_ (.B(_04221_),
    .C(_04222_),
    .A(_04200_),
    .Y(_04223_));
 sg13g2_nand2b_1 _11313_ (.Y(_04224_),
    .B(_04220_),
    .A_N(_04223_));
 sg13g2_nand2b_1 _11314_ (.Y(_04225_),
    .B(_04223_),
    .A_N(_04220_));
 sg13g2_and2_1 _11315_ (.A(net1771),
    .B(_04225_),
    .X(_04226_));
 sg13g2_xnor2_1 _11316_ (.Y(_04227_),
    .A(net1831),
    .B(net1829));
 sg13g2_o21ai_1 _11317_ (.B1(_04216_),
    .Y(_04228_),
    .A1(_00597_),
    .A2(net1828));
 sg13g2_o21ai_1 _11318_ (.B1(_04228_),
    .Y(_04229_),
    .A1(net1832),
    .A2(net1798));
 sg13g2_a21o_1 _11319_ (.A2(_04229_),
    .A1(_04227_),
    .B1(net1771),
    .X(_04230_));
 sg13g2_nor2_1 _11320_ (.A(_04227_),
    .B(_04229_),
    .Y(_04231_));
 sg13g2_o21ai_1 _11321_ (.B1(net1714),
    .Y(_04232_),
    .A1(_04230_),
    .A2(_04231_));
 sg13g2_a21oi_1 _11322_ (.A1(_04224_),
    .A2(_04226_),
    .Y(_04233_),
    .B1(_04232_));
 sg13g2_a21oi_1 _11323_ (.A1(_06880_),
    .A2(net1704),
    .Y(_00259_),
    .B1(_04233_));
 sg13g2_nor3_1 _11324_ (.A(net2124),
    .B(net1709),
    .C(_04230_),
    .Y(_04234_));
 sg13g2_a21oi_1 _11325_ (.A1(\vgadonut.donut.ysA[21] ),
    .A2(net1704),
    .Y(_04235_),
    .B1(_04234_));
 sg13g2_o21ai_1 _11326_ (.B1(_04225_),
    .Y(_04236_),
    .A1(_06880_),
    .A2(net1797));
 sg13g2_xor2_1 _11327_ (.B(net1830),
    .A(\vgadonut.donut.ysA[21] ),
    .X(_04237_));
 sg13g2_and2_1 _11328_ (.A(_04236_),
    .B(_04237_),
    .X(_04238_));
 sg13g2_o21ai_1 _11329_ (.B1(_04064_),
    .Y(_04239_),
    .A1(_04236_),
    .A2(_04237_));
 sg13g2_o21ai_1 _11330_ (.B1(net2125),
    .Y(_00260_),
    .A1(_04238_),
    .A2(_04239_));
 sg13g2_nand2_1 _11331_ (.Y(_04240_),
    .A(\vgadonut.donut.ycA[3] ),
    .B(\vgadonut.donut.cA[5] ));
 sg13g2_xor2_1 _11332_ (.B(\vgadonut.donut.cA[5] ),
    .A(\vgadonut.donut.ycA[3] ),
    .X(_04241_));
 sg13g2_xnor2_1 _11333_ (.Y(_04242_),
    .A(\vgadonut.donut.ycA[2] ),
    .B(\vgadonut.donut.cA[4] ));
 sg13g2_nand2_1 _11334_ (.Y(_04243_),
    .A(net2091),
    .B(\vgadonut.donut.cA[3] ));
 sg13g2_nand2_1 _11335_ (.Y(_04244_),
    .A(net1993),
    .B(net1825));
 sg13g2_xor2_1 _11336_ (.B(\vgadonut.donut.cA[3] ),
    .A(\vgadonut.donut.ycA[1] ),
    .X(_04245_));
 sg13g2_nand2b_1 _11337_ (.Y(_04246_),
    .B(_04245_),
    .A_N(_04244_));
 sg13g2_a21oi_1 _11338_ (.A1(_04243_),
    .A2(_04246_),
    .Y(_04247_),
    .B1(_04242_));
 sg13g2_a21oi_1 _11339_ (.A1(\vgadonut.donut.ycA[2] ),
    .A2(\vgadonut.donut.cA[4] ),
    .Y(_04248_),
    .B1(_04247_));
 sg13g2_nand2b_1 _11340_ (.Y(_04249_),
    .B(_04241_),
    .A_N(_04248_));
 sg13g2_xnor2_1 _11341_ (.Y(_04250_),
    .A(\vgadonut.donut.ycA[4] ),
    .B(\vgadonut.donut.cA[6] ));
 sg13g2_a21oi_1 _11342_ (.A1(_04240_),
    .A2(_04249_),
    .Y(_04251_),
    .B1(_04250_));
 sg13g2_nand3_1 _11343_ (.B(_04249_),
    .C(_04250_),
    .A(_04240_),
    .Y(_04252_));
 sg13g2_nand2b_1 _11344_ (.Y(_04253_),
    .B(_04252_),
    .A_N(_04251_));
 sg13g2_nand2_1 _11345_ (.Y(_04254_),
    .A(net1825),
    .B(net1710));
 sg13g2_a22oi_1 _11346_ (.Y(_04255_),
    .B1(_04254_),
    .B2(_04061_),
    .A2(_04253_),
    .A1(net1765));
 sg13g2_a21o_1 _11347_ (.A2(net1702),
    .A1(net2184),
    .B1(_04255_),
    .X(_00261_));
 sg13g2_a21o_1 _11348_ (.A2(\vgadonut.donut.cA[6] ),
    .A1(\vgadonut.donut.ycA[4] ),
    .B1(_04251_),
    .X(_04256_));
 sg13g2_nor2_1 _11349_ (.A(\vgadonut.donut.ycA[5] ),
    .B(net1824),
    .Y(_04257_));
 sg13g2_xor2_1 _11350_ (.B(net1824),
    .A(\vgadonut.donut.ycA[5] ),
    .X(_04258_));
 sg13g2_o21ai_1 _11351_ (.B1(net1765),
    .Y(_04259_),
    .A1(_04256_),
    .A2(_04258_));
 sg13g2_a21o_1 _11352_ (.A2(_04258_),
    .A1(_04256_),
    .B1(_04259_),
    .X(_04260_));
 sg13g2_a21oi_1 _11353_ (.A1(\vgadonut.donut.cA[3] ),
    .A2(net1774),
    .Y(_04261_),
    .B1(net1706));
 sg13g2_a22oi_1 _11354_ (.Y(_00262_),
    .B1(_04260_),
    .B2(_04261_),
    .A2(net1706),
    .A1(_06889_));
 sg13g2_xnor2_1 _11355_ (.Y(_04262_),
    .A(\vgadonut.donut.ycA[6] ),
    .B(net1823));
 sg13g2_a21oi_1 _11356_ (.A1(\vgadonut.donut.ycA[5] ),
    .A2(net1824),
    .Y(_04263_),
    .B1(_04256_));
 sg13g2_nor3_1 _11357_ (.A(_04257_),
    .B(_04262_),
    .C(_04263_),
    .Y(_04264_));
 sg13g2_o21ai_1 _11358_ (.B1(_04262_),
    .Y(_04265_),
    .A1(_04257_),
    .A2(_04263_));
 sg13g2_nand2b_1 _11359_ (.Y(_04266_),
    .B(_04265_),
    .A_N(_04264_));
 sg13g2_o21ai_1 _11360_ (.B1(net1710),
    .Y(_04267_),
    .A1(\vgadonut.donut.cA[4] ),
    .A2(net1766));
 sg13g2_a21oi_1 _11361_ (.A1(net1766),
    .A2(_04266_),
    .Y(_04268_),
    .B1(_04267_));
 sg13g2_a21o_1 _11362_ (.A2(net1702),
    .A1(net2191),
    .B1(_04268_),
    .X(_00263_));
 sg13g2_a21oi_1 _11363_ (.A1(\vgadonut.donut.ycA[6] ),
    .A2(net1823),
    .Y(_04269_),
    .B1(_04264_));
 sg13g2_xnor2_1 _11364_ (.Y(_04270_),
    .A(\vgadonut.donut.ycA[7] ),
    .B(net1822));
 sg13g2_nor2_1 _11365_ (.A(_04269_),
    .B(_04270_),
    .Y(_04271_));
 sg13g2_xnor2_1 _11366_ (.Y(_04272_),
    .A(_04269_),
    .B(_04270_));
 sg13g2_o21ai_1 _11367_ (.B1(net1711),
    .Y(_04273_),
    .A1(\vgadonut.donut.cA[5] ),
    .A2(net1765));
 sg13g2_a21oi_1 _11368_ (.A1(net1765),
    .A2(_04272_),
    .Y(_04274_),
    .B1(_04273_));
 sg13g2_a21o_1 _11369_ (.A2(net1702),
    .A1(net2137),
    .B1(_04274_),
    .X(_00264_));
 sg13g2_xnor2_1 _11370_ (.Y(_04275_),
    .A(\vgadonut.donut.ycA[8] ),
    .B(net1821));
 sg13g2_a21oi_1 _11371_ (.A1(\vgadonut.donut.ycA[7] ),
    .A2(net1822),
    .Y(_04276_),
    .B1(_04271_));
 sg13g2_or2_1 _11372_ (.X(_04277_),
    .B(_04276_),
    .A(_04275_));
 sg13g2_a21oi_1 _11373_ (.A1(_04275_),
    .A2(_04276_),
    .Y(_04278_),
    .B1(net1760));
 sg13g2_nand2_1 _11374_ (.Y(_04279_),
    .A(_00600_),
    .B(net1825));
 sg13g2_xor2_1 _11375_ (.B(net2194),
    .A(\vgadonut.donut.cA[6] ),
    .X(_04280_));
 sg13g2_a221oi_1 _11376_ (.B2(net1774),
    .C1(net1706),
    .B1(_04280_),
    .A1(_04277_),
    .Y(_04281_),
    .A2(_04278_));
 sg13g2_a21oi_1 _11377_ (.A1(_06895_),
    .A2(net1702),
    .Y(_00265_),
    .B1(_04281_));
 sg13g2_o21ai_1 _11378_ (.B1(_04277_),
    .Y(_04282_),
    .A1(_06895_),
    .A2(_00606_));
 sg13g2_nor2_1 _11379_ (.A(\vgadonut.donut.ycA[9] ),
    .B(net1819),
    .Y(_04283_));
 sg13g2_xnor2_1 _11380_ (.Y(_04284_),
    .A(\vgadonut.donut.ycA[9] ),
    .B(net1819));
 sg13g2_xnor2_1 _11381_ (.Y(_04285_),
    .A(_04282_),
    .B(_04284_));
 sg13g2_nor2_1 _11382_ (.A(\vgadonut.donut.cA[3] ),
    .B(_00604_),
    .Y(_04286_));
 sg13g2_xnor2_1 _11383_ (.Y(_04287_),
    .A(\vgadonut.donut.cA[3] ),
    .B(net1824));
 sg13g2_xnor2_1 _11384_ (.Y(_04288_),
    .A(_04279_),
    .B(_04287_));
 sg13g2_o21ai_1 _11385_ (.B1(net1711),
    .Y(_04289_),
    .A1(net1766),
    .A2(_04288_));
 sg13g2_a21oi_1 _11386_ (.A1(net1769),
    .A2(_04285_),
    .Y(_04290_),
    .B1(_04289_));
 sg13g2_a21oi_1 _11387_ (.A1(_06899_),
    .A2(net1702),
    .Y(_00266_),
    .B1(_04290_));
 sg13g2_xnor2_1 _11388_ (.Y(_04291_),
    .A(\vgadonut.donut.ycA[10] ),
    .B(net1817));
 sg13g2_a21oi_1 _11389_ (.A1(\vgadonut.donut.ycA[9] ),
    .A2(net1819),
    .Y(_04292_),
    .B1(_04282_));
 sg13g2_nor3_1 _11390_ (.A(_04283_),
    .B(_04291_),
    .C(_04292_),
    .Y(_04293_));
 sg13g2_o21ai_1 _11391_ (.B1(_04291_),
    .Y(_04294_),
    .A1(_04283_),
    .A2(_04292_));
 sg13g2_nand2_1 _11392_ (.Y(_04295_),
    .A(net1766),
    .B(_04294_));
 sg13g2_nand2_1 _11393_ (.Y(_04296_),
    .A(_00602_),
    .B(net1823));
 sg13g2_xor2_1 _11394_ (.B(net1823),
    .A(\vgadonut.donut.cA[4] ),
    .X(_04297_));
 sg13g2_a21oi_1 _11395_ (.A1(_04279_),
    .A2(_04287_),
    .Y(_04298_),
    .B1(_04286_));
 sg13g2_or2_1 _11396_ (.X(_04299_),
    .B(_04298_),
    .A(_04297_));
 sg13g2_a21oi_1 _11397_ (.A1(_04297_),
    .A2(_04298_),
    .Y(_04300_),
    .B1(net1769));
 sg13g2_a21oi_1 _11398_ (.A1(_04299_),
    .A2(_04300_),
    .Y(_04301_),
    .B1(net1706));
 sg13g2_o21ai_1 _11399_ (.B1(_04301_),
    .Y(_04302_),
    .A1(_04293_),
    .A2(_04295_));
 sg13g2_o21ai_1 _11400_ (.B1(_04302_),
    .Y(_04303_),
    .A1(net2287),
    .A2(net1711));
 sg13g2_inv_1 _11401_ (.Y(_00267_),
    .A(_04303_));
 sg13g2_a21o_1 _11402_ (.A2(net1817),
    .A1(\vgadonut.donut.ycA[10] ),
    .B1(_04293_),
    .X(_04304_));
 sg13g2_nor2_1 _11403_ (.A(\vgadonut.donut.ycA[11] ),
    .B(net1815),
    .Y(_04305_));
 sg13g2_xnor2_1 _11404_ (.Y(_04306_),
    .A(\vgadonut.donut.ycA[11] ),
    .B(net1815));
 sg13g2_xnor2_1 _11405_ (.Y(_04307_),
    .A(_04304_),
    .B(_04306_));
 sg13g2_nand2_1 _11406_ (.Y(_04308_),
    .A(_00601_),
    .B(net1822));
 sg13g2_xor2_1 _11407_ (.B(net1822),
    .A(\vgadonut.donut.cA[5] ),
    .X(_04309_));
 sg13g2_a21o_1 _11408_ (.A2(_04299_),
    .A1(_04296_),
    .B1(_04309_),
    .X(_04310_));
 sg13g2_nand3_1 _11409_ (.B(_04299_),
    .C(_04309_),
    .A(_04296_),
    .Y(_04311_));
 sg13g2_and2_1 _11410_ (.A(net1774),
    .B(_04311_),
    .X(_04312_));
 sg13g2_a221oi_1 _11411_ (.B2(_04312_),
    .C1(net1706),
    .B1(_04310_),
    .A1(net1766),
    .Y(_04313_),
    .A2(_04307_));
 sg13g2_a21oi_1 _11412_ (.A1(_06905_),
    .A2(net1702),
    .Y(_00268_),
    .B1(_04313_));
 sg13g2_xnor2_1 _11413_ (.Y(_04314_),
    .A(\vgadonut.donut.ycA[12] ),
    .B(net1814));
 sg13g2_a21oi_1 _11414_ (.A1(\vgadonut.donut.ycA[11] ),
    .A2(net1815),
    .Y(_04315_),
    .B1(_04304_));
 sg13g2_o21ai_1 _11415_ (.B1(_04314_),
    .Y(_04316_),
    .A1(_04305_),
    .A2(_04315_));
 sg13g2_nor3_1 _11416_ (.A(_04305_),
    .B(_04314_),
    .C(_04315_),
    .Y(_04317_));
 sg13g2_nand2_1 _11417_ (.Y(_04318_),
    .A(net1766),
    .B(_04316_));
 sg13g2_nand2_1 _11418_ (.Y(_04319_),
    .A(_00600_),
    .B(net1821));
 sg13g2_xor2_1 _11419_ (.B(net1821),
    .A(\vgadonut.donut.cA[6] ),
    .X(_04320_));
 sg13g2_a21o_1 _11420_ (.A2(_04310_),
    .A1(_04308_),
    .B1(_04320_),
    .X(_04321_));
 sg13g2_nand3_1 _11421_ (.B(_04310_),
    .C(_04320_),
    .A(_04308_),
    .Y(_04322_));
 sg13g2_nand3_1 _11422_ (.B(_04321_),
    .C(_04322_),
    .A(net1774),
    .Y(_04323_));
 sg13g2_and2_1 _11423_ (.A(net1711),
    .B(_04323_),
    .X(_04324_));
 sg13g2_o21ai_1 _11424_ (.B1(_04324_),
    .Y(_04325_),
    .A1(_04317_),
    .A2(_04318_));
 sg13g2_o21ai_1 _11425_ (.B1(_04325_),
    .Y(_04326_),
    .A1(net2309),
    .A2(net1711));
 sg13g2_inv_1 _11426_ (.Y(_00269_),
    .A(_04326_));
 sg13g2_nand2_1 _11427_ (.Y(_04327_),
    .A(\vgadonut.donut.ycA[13] ),
    .B(net1813));
 sg13g2_xor2_1 _11428_ (.B(net1813),
    .A(\vgadonut.donut.ycA[13] ),
    .X(_04328_));
 sg13g2_a21o_1 _11429_ (.A2(net1814),
    .A1(\vgadonut.donut.ycA[12] ),
    .B1(_04317_),
    .X(_04329_));
 sg13g2_xnor2_1 _11430_ (.Y(_04330_),
    .A(_04328_),
    .B(_04329_));
 sg13g2_nor2_1 _11431_ (.A(_00604_),
    .B(net1819),
    .Y(_04331_));
 sg13g2_nor2b_1 _11432_ (.A(net1824),
    .B_N(net1819),
    .Y(_04332_));
 sg13g2_or2_1 _11433_ (.X(_04333_),
    .B(_04332_),
    .A(_04331_));
 sg13g2_and2_1 _11434_ (.A(_04319_),
    .B(_04321_),
    .X(_04334_));
 sg13g2_or2_1 _11435_ (.X(_04335_),
    .B(_04334_),
    .A(_04333_));
 sg13g2_a21oi_1 _11436_ (.A1(_04333_),
    .A2(_04334_),
    .Y(_04336_),
    .B1(net1766));
 sg13g2_a21oi_1 _11437_ (.A1(_04335_),
    .A2(_04336_),
    .Y(_04337_),
    .B1(net1708));
 sg13g2_o21ai_1 _11438_ (.B1(_04337_),
    .Y(_04338_),
    .A1(net1760),
    .A2(_04330_));
 sg13g2_o21ai_1 _11439_ (.B1(_04338_),
    .Y(_04339_),
    .A1(net2337),
    .A2(net1713));
 sg13g2_inv_1 _11440_ (.Y(_00270_),
    .A(_04339_));
 sg13g2_xnor2_1 _11441_ (.Y(_04340_),
    .A(\vgadonut.donut.ycA[14] ),
    .B(net1813));
 sg13g2_o21ai_1 _11442_ (.B1(_04329_),
    .Y(_04341_),
    .A1(\vgadonut.donut.ycA[13] ),
    .A2(net1813));
 sg13g2_nand3_1 _11443_ (.B(_04340_),
    .C(_04341_),
    .A(_04327_),
    .Y(_04342_));
 sg13g2_a21o_1 _11444_ (.A2(_04341_),
    .A1(_04327_),
    .B1(_04340_),
    .X(_04343_));
 sg13g2_and3_1 _11445_ (.X(_04344_),
    .A(net1770),
    .B(_04342_),
    .C(_04343_));
 sg13g2_nand2b_1 _11446_ (.Y(_04345_),
    .B(net1817),
    .A_N(net1823));
 sg13g2_xor2_1 _11447_ (.B(net1817),
    .A(net1823),
    .X(_04346_));
 sg13g2_nor2_1 _11448_ (.A(_04331_),
    .B(_04334_),
    .Y(_04347_));
 sg13g2_nor2_2 _11449_ (.A(_04332_),
    .B(_04347_),
    .Y(_04348_));
 sg13g2_nor2_1 _11450_ (.A(_04346_),
    .B(_04348_),
    .Y(_04349_));
 sg13g2_and2_1 _11451_ (.A(_04346_),
    .B(_04348_),
    .X(_04350_));
 sg13g2_nor3_1 _11452_ (.A(net1770),
    .B(_04349_),
    .C(_04350_),
    .Y(_04351_));
 sg13g2_nor3_1 _11453_ (.A(net1708),
    .B(_04344_),
    .C(_04351_),
    .Y(_04352_));
 sg13g2_a21oi_1 _11454_ (.A1(_06911_),
    .A2(net1703),
    .Y(_00271_),
    .B1(_04352_));
 sg13g2_nand2_1 _11455_ (.Y(_04353_),
    .A(net2150),
    .B(net1809));
 sg13g2_xor2_1 _11456_ (.B(net1809),
    .A(\vgadonut.donut.ycA[15] ),
    .X(_04354_));
 sg13g2_o21ai_1 _11457_ (.B1(_04343_),
    .Y(_04355_),
    .A1(_06911_),
    .A2(_00607_));
 sg13g2_o21ai_1 _11458_ (.B1(net1770),
    .Y(_04356_),
    .A1(_04354_),
    .A2(_04355_));
 sg13g2_a21oi_1 _11459_ (.A1(_04354_),
    .A2(_04355_),
    .Y(_04357_),
    .B1(_04356_));
 sg13g2_xnor2_1 _11460_ (.Y(_04358_),
    .A(net1822),
    .B(net1815));
 sg13g2_o21ai_1 _11461_ (.B1(_04345_),
    .Y(_04359_),
    .A1(_04346_),
    .A2(_04348_));
 sg13g2_and2_1 _11462_ (.A(_04358_),
    .B(_04359_),
    .X(_04360_));
 sg13g2_o21ai_1 _11463_ (.B1(net1775),
    .Y(_04361_),
    .A1(_04358_),
    .A2(_04359_));
 sg13g2_o21ai_1 _11464_ (.B1(net1713),
    .Y(_04362_),
    .A1(_04360_),
    .A2(_04361_));
 sg13g2_nor2_1 _11465_ (.A(_04357_),
    .B(_04362_),
    .Y(_04363_));
 sg13g2_a21oi_1 _11466_ (.A1(_06914_),
    .A2(net1703),
    .Y(_00272_),
    .B1(_04363_));
 sg13g2_nor2_1 _11467_ (.A(net2158),
    .B(net1713),
    .Y(_04364_));
 sg13g2_nand2_1 _11468_ (.Y(_04365_),
    .A(\vgadonut.donut.ycA[16] ),
    .B(net1812));
 sg13g2_xnor2_1 _11469_ (.Y(_04366_),
    .A(\vgadonut.donut.ycA[16] ),
    .B(net1809));
 sg13g2_o21ai_1 _11470_ (.B1(_04355_),
    .Y(_04367_),
    .A1(\vgadonut.donut.ycA[15] ),
    .A2(net1809));
 sg13g2_a21o_2 _11471_ (.A2(_04367_),
    .A1(_04353_),
    .B1(_04366_),
    .X(_04368_));
 sg13g2_nand3_1 _11472_ (.B(_04366_),
    .C(_04367_),
    .A(_04353_),
    .Y(_04369_));
 sg13g2_nand3_1 _11473_ (.B(_04368_),
    .C(_04369_),
    .A(net1770),
    .Y(_04370_));
 sg13g2_xnor2_1 _11474_ (.Y(_04371_),
    .A(net1821),
    .B(net1814));
 sg13g2_a21o_1 _11475_ (.A2(net1815),
    .A1(_00605_),
    .B1(_04360_),
    .X(_04372_));
 sg13g2_and2_1 _11476_ (.A(_04371_),
    .B(_04372_),
    .X(_04373_));
 sg13g2_o21ai_1 _11477_ (.B1(net1775),
    .Y(_04374_),
    .A1(_04371_),
    .A2(_04372_));
 sg13g2_nor2_1 _11478_ (.A(_04373_),
    .B(_04374_),
    .Y(_04375_));
 sg13g2_nor2_1 _11479_ (.A(net1708),
    .B(_04375_),
    .Y(_04376_));
 sg13g2_a21oi_1 _11480_ (.A1(_04370_),
    .A2(_04376_),
    .Y(_00273_),
    .B1(_04364_));
 sg13g2_xnor2_1 _11481_ (.Y(_04377_),
    .A(\vgadonut.donut.ycA[17] ),
    .B(net1809));
 sg13g2_nand3_1 _11482_ (.B(_04368_),
    .C(_04377_),
    .A(_04365_),
    .Y(_04378_));
 sg13g2_a21o_1 _11483_ (.A2(_04368_),
    .A1(_04365_),
    .B1(_04377_),
    .X(_04379_));
 sg13g2_nand3_1 _11484_ (.B(_04378_),
    .C(_04379_),
    .A(net1770),
    .Y(_04380_));
 sg13g2_nand2b_1 _11485_ (.Y(_04381_),
    .B(net1820),
    .A_N(net1811));
 sg13g2_nor2b_1 _11486_ (.A(net1820),
    .B_N(net1811),
    .Y(_04382_));
 sg13g2_xnor2_1 _11487_ (.Y(_04383_),
    .A(net1820),
    .B(net1809));
 sg13g2_a21o_1 _11488_ (.A2(net1814),
    .A1(_00606_),
    .B1(_04373_),
    .X(_04384_));
 sg13g2_a21oi_1 _11489_ (.A1(_04383_),
    .A2(_04384_),
    .Y(_04385_),
    .B1(net1770));
 sg13g2_o21ai_1 _11490_ (.B1(_04385_),
    .Y(_04386_),
    .A1(_04383_),
    .A2(_04384_));
 sg13g2_nand3_1 _11491_ (.B(_04380_),
    .C(_04386_),
    .A(net1713),
    .Y(_04387_));
 sg13g2_o21ai_1 _11492_ (.B1(_04387_),
    .Y(_04388_),
    .A1(net2223),
    .A2(net1713));
 sg13g2_inv_1 _11493_ (.Y(_00274_),
    .A(_04388_));
 sg13g2_and2_1 _11494_ (.A(\vgadonut.donut.ycA[18] ),
    .B(net1810),
    .X(_04389_));
 sg13g2_xor2_1 _11495_ (.B(net1810),
    .A(\vgadonut.donut.ycA[18] ),
    .X(_04390_));
 sg13g2_o21ai_1 _11496_ (.B1(net1809),
    .Y(_04391_),
    .A1(\vgadonut.donut.ycA[16] ),
    .A2(\vgadonut.donut.ycA[17] ));
 sg13g2_nor2_1 _11497_ (.A(_04368_),
    .B(_04377_),
    .Y(_04392_));
 sg13g2_o21ai_1 _11498_ (.B1(_04391_),
    .Y(_04393_),
    .A1(_04368_),
    .A2(_04377_));
 sg13g2_xnor2_1 _11499_ (.Y(_04394_),
    .A(_04390_),
    .B(_04393_));
 sg13g2_nand2b_1 _11500_ (.Y(_04395_),
    .B(net1811),
    .A_N(net1818));
 sg13g2_xor2_1 _11501_ (.B(net1811),
    .A(net1818),
    .X(_04396_));
 sg13g2_a21oi_1 _11502_ (.A1(_04381_),
    .A2(_04384_),
    .Y(_04397_),
    .B1(_04382_));
 sg13g2_or2_1 _11503_ (.X(_04398_),
    .B(_04397_),
    .A(_04396_));
 sg13g2_a21oi_1 _11504_ (.A1(_04396_),
    .A2(_04397_),
    .Y(_04399_),
    .B1(net1773));
 sg13g2_a21oi_1 _11505_ (.A1(_04398_),
    .A2(_04399_),
    .Y(_04400_),
    .B1(net1708));
 sg13g2_o21ai_1 _11506_ (.B1(_04400_),
    .Y(_04401_),
    .A1(net1760),
    .A2(_04394_));
 sg13g2_o21ai_1 _11507_ (.B1(_04401_),
    .Y(_04402_),
    .A1(net2262),
    .A2(net1713));
 sg13g2_inv_1 _11508_ (.Y(_00275_),
    .A(_04402_));
 sg13g2_xor2_1 _11509_ (.B(net1810),
    .A(\vgadonut.donut.ycA[19] ),
    .X(_04403_));
 sg13g2_a21oi_1 _11510_ (.A1(_04390_),
    .A2(_04393_),
    .Y(_04404_),
    .B1(_04389_));
 sg13g2_xor2_1 _11511_ (.B(_04404_),
    .A(_04403_),
    .X(_04405_));
 sg13g2_nand2b_1 _11512_ (.Y(_04406_),
    .B(net1811),
    .A_N(net1816));
 sg13g2_nor2b_1 _11513_ (.A(net1811),
    .B_N(net1816),
    .Y(_04407_));
 sg13g2_xor2_1 _11514_ (.B(net1810),
    .A(net1816),
    .X(_04408_));
 sg13g2_and2_1 _11515_ (.A(_04395_),
    .B(_04398_),
    .X(_04409_));
 sg13g2_o21ai_1 _11516_ (.B1(net1777),
    .Y(_04410_),
    .A1(_04408_),
    .A2(_04409_));
 sg13g2_a21o_1 _11517_ (.A2(_04409_),
    .A1(_04408_),
    .B1(_04410_),
    .X(_04411_));
 sg13g2_o21ai_1 _11518_ (.B1(_04411_),
    .Y(_04412_),
    .A1(net1760),
    .A2(_04405_));
 sg13g2_mux2_1 _11519_ (.A0(_04412_),
    .A1(net2175),
    .S(net1703),
    .X(_00276_));
 sg13g2_xnor2_1 _11520_ (.Y(_04413_),
    .A(\vgadonut.donut.ycA[20] ),
    .B(net1812));
 sg13g2_nand3_1 _11521_ (.B(_04392_),
    .C(_04403_),
    .A(_04390_),
    .Y(_04414_));
 sg13g2_o21ai_1 _11522_ (.B1(net1810),
    .Y(_04415_),
    .A1(\vgadonut.donut.ycA[18] ),
    .A2(\vgadonut.donut.ycA[19] ));
 sg13g2_nand3_1 _11523_ (.B(_04414_),
    .C(_04415_),
    .A(_04391_),
    .Y(_04416_));
 sg13g2_nor2b_1 _11524_ (.A(_04416_),
    .B_N(_04413_),
    .Y(_04417_));
 sg13g2_nor2b_1 _11525_ (.A(_04413_),
    .B_N(_04416_),
    .Y(_04418_));
 sg13g2_nor3_1 _11526_ (.A(net1777),
    .B(_04417_),
    .C(_04418_),
    .Y(_04419_));
 sg13g2_xnor2_1 _11527_ (.Y(_04420_),
    .A(net1814),
    .B(net1811));
 sg13g2_o21ai_1 _11528_ (.B1(_04406_),
    .Y(_04421_),
    .A1(_04407_),
    .A2(_04409_));
 sg13g2_a21o_1 _11529_ (.A2(_04421_),
    .A1(_04420_),
    .B1(net1770),
    .X(_04422_));
 sg13g2_nor2_1 _11530_ (.A(_04420_),
    .B(_04421_),
    .Y(_04423_));
 sg13g2_o21ai_1 _11531_ (.B1(net1716),
    .Y(_04424_),
    .A1(_04422_),
    .A2(_04423_));
 sg13g2_nor2_1 _11532_ (.A(_04419_),
    .B(_04424_),
    .Y(_04425_));
 sg13g2_a21oi_1 _11533_ (.A1(_00554_),
    .A2(net1703),
    .Y(_00277_),
    .B1(_04425_));
 sg13g2_a21oi_1 _11534_ (.A1(\vgadonut.donut.ycA[20] ),
    .A2(net1810),
    .Y(_04426_),
    .B1(_04418_));
 sg13g2_xnor2_1 _11535_ (.Y(_04427_),
    .A(\vgadonut.donut.ycA[21] ),
    .B(net1810));
 sg13g2_o21ai_1 _11536_ (.B1(net1770),
    .Y(_04428_),
    .A1(_04426_),
    .A2(_04427_));
 sg13g2_a21oi_1 _11537_ (.A1(_04426_),
    .A2(_04427_),
    .Y(_04429_),
    .B1(_04428_));
 sg13g2_o21ai_1 _11538_ (.B1(net1716),
    .Y(_04430_),
    .A1(net1810),
    .A2(_04422_));
 sg13g2_nor2_1 _11539_ (.A(_04429_),
    .B(_04430_),
    .Y(_04431_));
 sg13g2_a21oi_1 _11540_ (.A1(_00558_),
    .A2(net1703),
    .Y(_00278_),
    .B1(_04431_));
 sg13g2_a21oi_1 _11541_ (.A1(net1825),
    .A2(net1710),
    .Y(_04432_),
    .B1(net1993));
 sg13g2_a21oi_1 _11542_ (.A1(net1765),
    .A2(_04244_),
    .Y(_04433_),
    .B1(net1706));
 sg13g2_nor2_1 _11543_ (.A(net1994),
    .B(_04433_),
    .Y(_00279_));
 sg13g2_xnor2_1 _11544_ (.Y(_04434_),
    .A(_04244_),
    .B(_04245_));
 sg13g2_nand3_1 _11545_ (.B(net1710),
    .C(_04434_),
    .A(net1765),
    .Y(_04435_));
 sg13g2_o21ai_1 _11546_ (.B1(_04435_),
    .Y(_00280_),
    .A1(_06883_),
    .A2(net1710));
 sg13g2_nand2_1 _11547_ (.Y(_04436_),
    .A(net2136),
    .B(net1706));
 sg13g2_nand3_1 _11548_ (.B(_04243_),
    .C(_04246_),
    .A(_04242_),
    .Y(_04437_));
 sg13g2_nand2b_1 _11549_ (.Y(_04438_),
    .B(_04437_),
    .A_N(_04247_));
 sg13g2_o21ai_1 _11550_ (.B1(_04436_),
    .Y(_00281_),
    .A1(_04061_),
    .A2(_04438_));
 sg13g2_nand2b_1 _11551_ (.Y(_04439_),
    .B(_04248_),
    .A_N(_04241_));
 sg13g2_nand4_1 _11552_ (.B(net1710),
    .C(_04249_),
    .A(net1765),
    .Y(_04440_),
    .D(_04439_));
 sg13g2_o21ai_1 _11553_ (.B1(_04440_),
    .Y(_00282_),
    .A1(_06885_),
    .A2(net1710));
 sg13g2_o21ai_1 _11554_ (.B1(net1642),
    .Y(_00283_),
    .A1(net1646),
    .A2(_00755_));
 sg13g2_a21oi_1 _11555_ (.A1(net1854),
    .A2(net1712),
    .Y(_04441_),
    .B1(net2018));
 sg13g2_a21oi_1 _11556_ (.A1(net1767),
    .A2(_04051_),
    .Y(_04442_),
    .B1(net1707));
 sg13g2_nor2_1 _11557_ (.A(net2019),
    .B(_04442_),
    .Y(_00284_));
 sg13g2_nand2_1 _11558_ (.Y(_04443_),
    .A(net2038),
    .B(net1707));
 sg13g2_xnor2_1 _11559_ (.Y(_04444_),
    .A(_04051_),
    .B(_04052_));
 sg13g2_o21ai_1 _11560_ (.B1(_04443_),
    .Y(_00285_),
    .A1(_04061_),
    .A2(_04444_));
 sg13g2_nand2_1 _11561_ (.Y(_04445_),
    .A(net2053),
    .B(net1707));
 sg13g2_xor2_1 _11562_ (.B(_04054_),
    .A(_04053_),
    .X(_04446_));
 sg13g2_o21ai_1 _11563_ (.B1(_04445_),
    .Y(_00286_),
    .A1(_04061_),
    .A2(_04446_));
 sg13g2_nand3_1 _11564_ (.B(_04049_),
    .C(_04055_),
    .A(_04048_),
    .Y(_04447_));
 sg13g2_nand4_1 _11565_ (.B(net1712),
    .C(_04056_),
    .A(net1767),
    .Y(_04448_),
    .D(_04447_));
 sg13g2_o21ai_1 _11566_ (.B1(_04448_),
    .Y(_00287_),
    .A1(_06850_),
    .A2(net1712));
 sg13g2_nand2_1 _11567_ (.Y(_04449_),
    .A(net1456),
    .B(net1718));
 sg13g2_nand2b_1 _11568_ (.Y(_04450_),
    .B(net1932),
    .A_N(\vgadonut.donut.cAcB[0] ));
 sg13g2_xnor2_1 _11569_ (.Y(_04451_),
    .A(\vgadonut.donut.cAcB[0] ),
    .B(net1932));
 sg13g2_nor2b_1 _11570_ (.A(\vgadonut.donut.sAsB[11] ),
    .B_N(\vgadonut.donut.cAsB[6] ),
    .Y(_04452_));
 sg13g2_nand2b_1 _11571_ (.Y(_04453_),
    .B(net1888),
    .A_N(net1906));
 sg13g2_nand2b_1 _11572_ (.Y(_04454_),
    .B(_04453_),
    .A_N(_04452_));
 sg13g2_nor2_1 _11573_ (.A(net1907),
    .B(_06903_),
    .Y(_04455_));
 sg13g2_nand2_1 _11574_ (.Y(_04456_),
    .A(\vgadonut.donut.cAsB[5] ),
    .B(_06903_));
 sg13g2_nor2b_1 _11575_ (.A(\vgadonut.donut.sAsB[7] ),
    .B_N(\vgadonut.donut.cAsB[2] ),
    .Y(_04457_));
 sg13g2_xnor2_1 _11576_ (.Y(_04458_),
    .A(\vgadonut.donut.cAsB[2] ),
    .B(\vgadonut.donut.sAsB[7] ));
 sg13g2_nor2b_1 _11577_ (.A(\vgadonut.donut.sAsB[6] ),
    .B_N(\vgadonut.donut.cAsB[1] ),
    .Y(_04459_));
 sg13g2_nand2b_1 _11578_ (.Y(_04460_),
    .B(\vgadonut.donut.sAsB[5] ),
    .A_N(net1912));
 sg13g2_xnor2_1 _11579_ (.Y(_04461_),
    .A(\vgadonut.donut.cAsB[1] ),
    .B(\vgadonut.donut.sAsB[6] ));
 sg13g2_a21oi_1 _11580_ (.A1(_04460_),
    .A2(_04461_),
    .Y(_04462_),
    .B1(_04459_));
 sg13g2_inv_1 _11581_ (.Y(_04463_),
    .A(_04462_));
 sg13g2_a21oi_1 _11582_ (.A1(_04458_),
    .A2(_04463_),
    .Y(_04464_),
    .B1(_04457_));
 sg13g2_xnor2_1 _11583_ (.Y(_04465_),
    .A(net1909),
    .B(\vgadonut.donut.sAsB[8] ));
 sg13g2_nor2b_1 _11584_ (.A(_04464_),
    .B_N(_04465_),
    .Y(_04466_));
 sg13g2_a21oi_1 _11585_ (.A1(\vgadonut.donut.cAsB[3] ),
    .A2(_06896_),
    .Y(_04467_),
    .B1(_04466_));
 sg13g2_xnor2_1 _11586_ (.Y(_04468_),
    .A(\vgadonut.donut.cAsB[4] ),
    .B(\vgadonut.donut.sAsB[9] ));
 sg13g2_nor2b_1 _11587_ (.A(_04467_),
    .B_N(_04468_),
    .Y(_04469_));
 sg13g2_a21oi_1 _11588_ (.A1(net1908),
    .A2(_06900_),
    .Y(_04470_),
    .B1(_04469_));
 sg13g2_o21ai_1 _11589_ (.B1(_04456_),
    .Y(_04471_),
    .A1(_04455_),
    .A2(_04470_));
 sg13g2_xnor2_1 _11590_ (.Y(_04472_),
    .A(_04454_),
    .B(_04471_));
 sg13g2_nand2_1 _11591_ (.Y(_04473_),
    .A(_04451_),
    .B(_04472_));
 sg13g2_xnor2_1 _11592_ (.Y(_04474_),
    .A(_04451_),
    .B(_04472_));
 sg13g2_nor2b_1 _11593_ (.A(net1869),
    .B_N(net1862),
    .Y(_04475_));
 sg13g2_nand2b_1 _11594_ (.Y(_04476_),
    .B(net1869),
    .A_N(net1862));
 sg13g2_nand2b_1 _11595_ (.Y(_04477_),
    .B(_04476_),
    .A_N(_04475_));
 sg13g2_nor2_1 _11596_ (.A(\vgadonut.donut.cB[13] ),
    .B(_00592_),
    .Y(_04478_));
 sg13g2_nand2_1 _11597_ (.Y(_04479_),
    .A(\vgadonut.donut.cB[13] ),
    .B(_00592_));
 sg13g2_xor2_1 _11598_ (.B(net1868),
    .A(\vgadonut.donut.cB[12] ),
    .X(_04480_));
 sg13g2_nor2b_1 _11599_ (.A(net1868),
    .B_N(\vgadonut.donut.cB[11] ),
    .Y(_04481_));
 sg13g2_nand2b_1 _11600_ (.Y(_04482_),
    .B(net1868),
    .A_N(\vgadonut.donut.cB[11] ));
 sg13g2_xnor2_1 _11601_ (.Y(_04483_),
    .A(\vgadonut.donut.cB[10] ),
    .B(net1868));
 sg13g2_nor2b_1 _11602_ (.A(net1868),
    .B_N(\vgadonut.donut.cB[9] ),
    .Y(_04484_));
 sg13g2_nand2b_1 _11603_ (.Y(_04485_),
    .B(net1868),
    .A_N(\vgadonut.donut.cB[9] ));
 sg13g2_xnor2_1 _11604_ (.Y(_04486_),
    .A(\vgadonut.donut.cB[7] ),
    .B(net1873));
 sg13g2_xor2_1 _11605_ (.B(net1876),
    .A(\vgadonut.donut.cB[6] ),
    .X(_04487_));
 sg13g2_xor2_1 _11606_ (.B(net1877),
    .A(\vgadonut.donut.cB[5] ),
    .X(_04488_));
 sg13g2_xor2_1 _11607_ (.B(net1879),
    .A(\vgadonut.donut.cB[4] ),
    .X(_04489_));
 sg13g2_nor2_1 _11608_ (.A(_00561_),
    .B(net1880),
    .Y(_04490_));
 sg13g2_nand2b_1 _11609_ (.Y(_04491_),
    .B(net1864),
    .A_N(net1882));
 sg13g2_xor2_1 _11610_ (.B(net1882),
    .A(net1864),
    .X(_04492_));
 sg13g2_nor2b_1 _11611_ (.A(net1867),
    .B_N(net1883),
    .Y(_04493_));
 sg13g2_xor2_1 _11612_ (.B(\vgadonut.donut.donuthit.cordicxy.x2in[5] ),
    .A(net1866),
    .X(_04494_));
 sg13g2_nor2_1 _11613_ (.A(_04493_),
    .B(_04494_),
    .Y(_04495_));
 sg13g2_a21oi_1 _11614_ (.A1(net1866),
    .A2(_00577_),
    .Y(_04496_),
    .B1(_04495_));
 sg13g2_o21ai_1 _11615_ (.B1(_04491_),
    .Y(_04497_),
    .A1(_04492_),
    .A2(_04496_));
 sg13g2_xnor2_1 _11616_ (.Y(_04498_),
    .A(net1863),
    .B(net1880));
 sg13g2_a21oi_1 _11617_ (.A1(_04497_),
    .A2(_04498_),
    .Y(_04499_),
    .B1(_04490_));
 sg13g2_nor2_1 _11618_ (.A(_04489_),
    .B(_04499_),
    .Y(_04500_));
 sg13g2_a21oi_1 _11619_ (.A1(\vgadonut.donut.cB[4] ),
    .A2(_00583_),
    .Y(_04501_),
    .B1(_04500_));
 sg13g2_nor2_1 _11620_ (.A(_04488_),
    .B(_04501_),
    .Y(_04502_));
 sg13g2_a21oi_1 _11621_ (.A1(\vgadonut.donut.cB[5] ),
    .A2(_00585_),
    .Y(_04503_),
    .B1(_04502_));
 sg13g2_nor2_1 _11622_ (.A(_04487_),
    .B(_04503_),
    .Y(_04504_));
 sg13g2_a21oi_1 _11623_ (.A1(\vgadonut.donut.cB[6] ),
    .A2(_00587_),
    .Y(_04505_),
    .B1(_04504_));
 sg13g2_nand2b_1 _11624_ (.Y(_04506_),
    .B(_04486_),
    .A_N(_04505_));
 sg13g2_o21ai_1 _11625_ (.B1(_04506_),
    .Y(_04507_),
    .A1(_00566_),
    .A2(net1873));
 sg13g2_xnor2_1 _11626_ (.Y(_04508_),
    .A(\vgadonut.donut.cB[8] ),
    .B(net1871));
 sg13g2_nand2_1 _11627_ (.Y(_04509_),
    .A(_04507_),
    .B(_04508_));
 sg13g2_o21ai_1 _11628_ (.B1(_04509_),
    .Y(_04510_),
    .A1(_00568_),
    .A2(net1871));
 sg13g2_nor2b_1 _11629_ (.A(_04484_),
    .B_N(_04485_),
    .Y(_04511_));
 sg13g2_a21oi_1 _11630_ (.A1(_04485_),
    .A2(_04510_),
    .Y(_04512_),
    .B1(_04484_));
 sg13g2_nand2b_1 _11631_ (.Y(_04513_),
    .B(_04483_),
    .A_N(_04512_));
 sg13g2_o21ai_1 _11632_ (.B1(_04513_),
    .Y(_04514_),
    .A1(_00572_),
    .A2(net1868));
 sg13g2_nor2b_1 _11633_ (.A(_04481_),
    .B_N(_04482_),
    .Y(_04515_));
 sg13g2_a21oi_1 _11634_ (.A1(_04482_),
    .A2(_04514_),
    .Y(_04516_),
    .B1(_04481_));
 sg13g2_nor2_1 _11635_ (.A(_04480_),
    .B(_04516_),
    .Y(_04517_));
 sg13g2_a21oi_1 _11636_ (.A1(\vgadonut.donut.cB[12] ),
    .A2(_00592_),
    .Y(_04518_),
    .B1(_04517_));
 sg13g2_o21ai_1 _11637_ (.B1(_04479_),
    .Y(_04519_),
    .A1(_04478_),
    .A2(_04518_));
 sg13g2_a21oi_2 _11638_ (.B1(_04475_),
    .Y(_04520_),
    .A2(_04519_),
    .A1(_04476_));
 sg13g2_xnor2_1 _11639_ (.Y(_04521_),
    .A(net1861),
    .B(_04520_));
 sg13g2_xnor2_1 _11640_ (.Y(_04522_),
    .A(net1861),
    .B(net1868));
 sg13g2_xnor2_1 _11641_ (.Y(_04523_),
    .A(_04520_),
    .B(_04522_));
 sg13g2_inv_1 _11642_ (.Y(_04524_),
    .A(net1601));
 sg13g2_nor2_1 _11643_ (.A(_00126_),
    .B(_04524_),
    .Y(_04525_));
 sg13g2_xnor2_1 _11644_ (.Y(_04526_),
    .A(_00126_),
    .B(net1601));
 sg13g2_nor2b_1 _11645_ (.A(net1601),
    .B_N(_00127_),
    .Y(_04527_));
 sg13g2_nand2b_1 _11646_ (.Y(_04528_),
    .B(net1600),
    .A_N(_00127_));
 sg13g2_nand2_1 _11647_ (.Y(_04529_),
    .A(_00610_),
    .B(net1600));
 sg13g2_xnor2_1 _11648_ (.Y(_04530_),
    .A(_04477_),
    .B(_04519_));
 sg13g2_nand2_1 _11649_ (.Y(_04531_),
    .A(_00612_),
    .B(_04530_));
 sg13g2_nor2b_1 _11650_ (.A(_04478_),
    .B_N(_04479_),
    .Y(_04532_));
 sg13g2_xnor2_1 _11651_ (.Y(_04533_),
    .A(_04518_),
    .B(_04532_));
 sg13g2_and2_1 _11652_ (.A(_00613_),
    .B(_04533_),
    .X(_04534_));
 sg13g2_xnor2_1 _11653_ (.Y(_04535_),
    .A(_04480_),
    .B(_04516_));
 sg13g2_nand2b_1 _11654_ (.Y(_04536_),
    .B(_00614_),
    .A_N(_04535_));
 sg13g2_xnor2_1 _11655_ (.Y(_04537_),
    .A(_04514_),
    .B(_04515_));
 sg13g2_nor2_1 _11656_ (.A(_00135_),
    .B(_04537_),
    .Y(_04538_));
 sg13g2_xnor2_1 _11657_ (.Y(_04539_),
    .A(_04483_),
    .B(_04512_));
 sg13g2_inv_1 _11658_ (.Y(_04540_),
    .A(_04539_));
 sg13g2_xnor2_1 _11659_ (.Y(_04541_),
    .A(_04510_),
    .B(_04511_));
 sg13g2_nor2_1 _11660_ (.A(_00137_),
    .B(_04541_),
    .Y(_04542_));
 sg13g2_xor2_1 _11661_ (.B(_04508_),
    .A(_04507_),
    .X(_04543_));
 sg13g2_xnor2_1 _11662_ (.Y(_04544_),
    .A(_04486_),
    .B(_04505_));
 sg13g2_inv_1 _11663_ (.Y(_04545_),
    .A(_04544_));
 sg13g2_nand2_1 _11664_ (.Y(_04546_),
    .A(\vgadonut.donut.sB[1] ),
    .B(_04544_));
 sg13g2_xor2_1 _11665_ (.B(_04503_),
    .A(_04487_),
    .X(_04547_));
 sg13g2_inv_1 _11666_ (.Y(_04548_),
    .A(_04547_));
 sg13g2_nand2_1 _11667_ (.Y(_04549_),
    .A(\vgadonut.donut.sB[0] ),
    .B(_04547_));
 sg13g2_xnor2_1 _11668_ (.Y(_04550_),
    .A(\vgadonut.donut.sB[1] ),
    .B(_04544_));
 sg13g2_o21ai_1 _11669_ (.B1(_04546_),
    .Y(_04551_),
    .A1(_04549_),
    .A2(_04550_));
 sg13g2_xnor2_1 _11670_ (.Y(_04552_),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[0] ),
    .B(_04543_));
 sg13g2_inv_1 _11671_ (.Y(_04553_),
    .A(_04552_));
 sg13g2_a22oi_1 _11672_ (.Y(_04554_),
    .B1(_04551_),
    .B2(_04553_),
    .A2(_04543_),
    .A1(_00617_));
 sg13g2_xnor2_1 _11673_ (.Y(_04555_),
    .A(_00137_),
    .B(_04541_));
 sg13g2_nor2_1 _11674_ (.A(_04554_),
    .B(_04555_),
    .Y(_04556_));
 sg13g2_nor2_1 _11675_ (.A(_04542_),
    .B(_04556_),
    .Y(_04557_));
 sg13g2_xnor2_1 _11676_ (.Y(_04558_),
    .A(net1884),
    .B(_04539_));
 sg13g2_nor2_1 _11677_ (.A(_04557_),
    .B(_04558_),
    .Y(_04559_));
 sg13g2_a21oi_1 _11678_ (.A1(_00616_),
    .A2(_04539_),
    .Y(_04560_),
    .B1(_04559_));
 sg13g2_inv_1 _11679_ (.Y(_04561_),
    .A(_04560_));
 sg13g2_xnor2_1 _11680_ (.Y(_04562_),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[3] ),
    .B(_04537_));
 sg13g2_a21oi_1 _11681_ (.A1(_04561_),
    .A2(_04562_),
    .Y(_04563_),
    .B1(_04538_));
 sg13g2_xor2_1 _11682_ (.B(_04535_),
    .A(net1883),
    .X(_04564_));
 sg13g2_o21ai_1 _11683_ (.B1(_04536_),
    .Y(_04565_),
    .A1(_04563_),
    .A2(_04564_));
 sg13g2_xnor2_1 _11684_ (.Y(_04566_),
    .A(_00133_),
    .B(_04533_));
 sg13g2_a21oi_1 _11685_ (.A1(_04565_),
    .A2(_04566_),
    .Y(_04567_),
    .B1(_04534_));
 sg13g2_xnor2_1 _11686_ (.Y(_04568_),
    .A(net1882),
    .B(_04530_));
 sg13g2_or2_1 _11687_ (.X(_04569_),
    .B(_04568_),
    .A(_04567_));
 sg13g2_xnor2_1 _11688_ (.Y(_04570_),
    .A(net1880),
    .B(net1600));
 sg13g2_a21oi_1 _11689_ (.A1(_04531_),
    .A2(_04569_),
    .Y(_04571_),
    .B1(_04570_));
 sg13g2_a21oi_1 _11690_ (.A1(_00611_),
    .A2(net1600),
    .Y(_04572_),
    .B1(_04571_));
 sg13g2_xnor2_1 _11691_ (.Y(_04573_),
    .A(_00583_),
    .B(net1600));
 sg13g2_nand2b_1 _11692_ (.Y(_04574_),
    .B(_04573_),
    .A_N(_04572_));
 sg13g2_o21ai_1 _11693_ (.B1(_04574_),
    .Y(_04575_),
    .A1(_00130_),
    .A2(_04524_));
 sg13g2_o21ai_1 _11694_ (.B1(_04575_),
    .Y(_04576_),
    .A1(_00610_),
    .A2(net1600));
 sg13g2_xnor2_1 _11695_ (.Y(_04577_),
    .A(net1876),
    .B(net1601));
 sg13g2_a21oi_1 _11696_ (.A1(_04529_),
    .A2(_04576_),
    .Y(_04578_),
    .B1(_04577_));
 sg13g2_a21oi_1 _11697_ (.A1(_00609_),
    .A2(net1600),
    .Y(_04579_),
    .B1(_04578_));
 sg13g2_o21ai_1 _11698_ (.B1(_04528_),
    .Y(_04580_),
    .A1(_04527_),
    .A2(_04579_));
 sg13g2_a21oi_1 _11699_ (.A1(_04526_),
    .A2(_04580_),
    .Y(_04581_),
    .B1(_04525_));
 sg13g2_xnor2_1 _11700_ (.Y(_04582_),
    .A(_04521_),
    .B(_04581_));
 sg13g2_and2_2 _11701_ (.A(net1870),
    .B(_04582_),
    .X(_04583_));
 sg13g2_nor2_1 _11702_ (.A(net1732),
    .B(_04583_),
    .Y(_04584_));
 sg13g2_or2_1 _11703_ (.X(_04585_),
    .B(_04583_),
    .A(net1731));
 sg13g2_or2_2 _11704_ (.X(_04586_),
    .B(_04583_),
    .A(_03930_));
 sg13g2_nor2_2 _11705_ (.A(_03933_),
    .B(_04583_),
    .Y(_04587_));
 sg13g2_o21ai_1 _11706_ (.B1(_04449_),
    .Y(_00294_),
    .A1(_04474_),
    .A2(net1552));
 sg13g2_nand2_1 _11707_ (.Y(_04588_),
    .A(net1455),
    .B(net1717));
 sg13g2_a21oi_1 _11708_ (.A1(_04453_),
    .A2(_04471_),
    .Y(_04589_),
    .B1(_04452_));
 sg13g2_xnor2_1 _11709_ (.Y(_04590_),
    .A(net1905),
    .B(\vgadonut.donut.sAsB[12] ));
 sg13g2_nand2b_1 _11710_ (.Y(_04591_),
    .B(_04590_),
    .A_N(_04589_));
 sg13g2_xnor2_1 _11711_ (.Y(_04592_),
    .A(_04589_),
    .B(_04590_));
 sg13g2_nor2b_1 _11712_ (.A(net1931),
    .B_N(\vgadonut.donut.cAcB[1] ),
    .Y(_04593_));
 sg13g2_xnor2_1 _11713_ (.Y(_04594_),
    .A(\vgadonut.donut.cAcB[1] ),
    .B(net1931));
 sg13g2_xor2_1 _11714_ (.B(_04594_),
    .A(_04450_),
    .X(_04595_));
 sg13g2_nor2b_1 _11715_ (.A(_04592_),
    .B_N(_04595_),
    .Y(_04596_));
 sg13g2_xnor2_1 _11716_ (.Y(_04597_),
    .A(_04592_),
    .B(_04595_));
 sg13g2_xor2_1 _11717_ (.B(_04597_),
    .A(_04473_),
    .X(_04598_));
 sg13g2_o21ai_1 _11718_ (.B1(_04588_),
    .Y(_00295_),
    .A1(net1551),
    .A2(_04598_));
 sg13g2_nand2_1 _11719_ (.Y(_04599_),
    .A(net1474),
    .B(net1717));
 sg13g2_a21oi_1 _11720_ (.A1(_04473_),
    .A2(_04597_),
    .Y(_04600_),
    .B1(_04596_));
 sg13g2_nor2b_1 _11721_ (.A(\vgadonut.donut.sAsB[13] ),
    .B_N(net1904),
    .Y(_04601_));
 sg13g2_xnor2_1 _11722_ (.Y(_04602_),
    .A(net1904),
    .B(\vgadonut.donut.sAsB[13] ));
 sg13g2_o21ai_1 _11723_ (.B1(_04591_),
    .Y(_04603_),
    .A1(_06859_),
    .A2(net1887));
 sg13g2_and2_1 _11724_ (.A(_04602_),
    .B(_04603_),
    .X(_04604_));
 sg13g2_xnor2_1 _11725_ (.Y(_04605_),
    .A(_04602_),
    .B(_04603_));
 sg13g2_a21oi_1 _11726_ (.A1(_04450_),
    .A2(_04594_),
    .Y(_04606_),
    .B1(_04593_));
 sg13g2_xnor2_1 _11727_ (.Y(_04607_),
    .A(\vgadonut.donut.cAcB[2] ),
    .B(net1930));
 sg13g2_nand2b_1 _11728_ (.Y(_04608_),
    .B(_04607_),
    .A_N(_04606_));
 sg13g2_xnor2_1 _11729_ (.Y(_04609_),
    .A(_04606_),
    .B(_04607_));
 sg13g2_nand2_1 _11730_ (.Y(_04610_),
    .A(_04605_),
    .B(_04609_));
 sg13g2_xnor2_1 _11731_ (.Y(_04611_),
    .A(_04605_),
    .B(_04609_));
 sg13g2_or2_1 _11732_ (.X(_04612_),
    .B(_04611_),
    .A(_04600_));
 sg13g2_xor2_1 _11733_ (.B(_04611_),
    .A(_04600_),
    .X(_04613_));
 sg13g2_o21ai_1 _11734_ (.B1(_04599_),
    .Y(_00296_),
    .A1(net1551),
    .A2(_04613_));
 sg13g2_nand2_1 _11735_ (.Y(_04614_),
    .A(net1479),
    .B(net1717));
 sg13g2_o21ai_1 _11736_ (.B1(_04608_),
    .Y(_04615_),
    .A1(_06860_),
    .A2(net1930));
 sg13g2_nor2b_1 _11737_ (.A(net1929),
    .B_N(net1957),
    .Y(_04616_));
 sg13g2_xnor2_1 _11738_ (.Y(_04617_),
    .A(net1957),
    .B(net1929));
 sg13g2_xor2_1 _11739_ (.B(_04617_),
    .A(_04615_),
    .X(_04618_));
 sg13g2_nor2b_1 _11740_ (.A(\vgadonut.donut.sAsB[14] ),
    .B_N(net1903),
    .Y(_04619_));
 sg13g2_nand2b_1 _11741_ (.Y(_04620_),
    .B(\vgadonut.donut.sAsB[14] ),
    .A_N(net1903));
 sg13g2_nor2b_1 _11742_ (.A(_04619_),
    .B_N(_04620_),
    .Y(_04621_));
 sg13g2_nor2_1 _11743_ (.A(_04601_),
    .B(_04604_),
    .Y(_04622_));
 sg13g2_xor2_1 _11744_ (.B(_04622_),
    .A(_04621_),
    .X(_04623_));
 sg13g2_and2_1 _11745_ (.A(_04618_),
    .B(_04623_),
    .X(_04624_));
 sg13g2_xnor2_1 _11746_ (.Y(_04625_),
    .A(_04618_),
    .B(_04623_));
 sg13g2_a21oi_1 _11747_ (.A1(_04610_),
    .A2(_04612_),
    .Y(_04626_),
    .B1(_04625_));
 sg13g2_nand3_1 _11748_ (.B(_04612_),
    .C(_04625_),
    .A(_04610_),
    .Y(_04627_));
 sg13g2_nor2b_1 _11749_ (.A(_04626_),
    .B_N(_04627_),
    .Y(_04628_));
 sg13g2_o21ai_1 _11750_ (.B1(_04614_),
    .Y(_00297_),
    .A1(net1551),
    .A2(_04628_));
 sg13g2_nand2_1 _11751_ (.Y(_04629_),
    .A(net1489),
    .B(net1721));
 sg13g2_xnor2_1 _11752_ (.Y(_04630_),
    .A(net1902),
    .B(net1885));
 sg13g2_nand2_1 _11753_ (.Y(_04631_),
    .A(_04604_),
    .B(_04621_));
 sg13g2_o21ai_1 _11754_ (.B1(_04620_),
    .Y(_04632_),
    .A1(_04601_),
    .A2(_04619_));
 sg13g2_and2_1 _11755_ (.A(_04631_),
    .B(_04632_),
    .X(_04633_));
 sg13g2_nand2b_1 _11756_ (.Y(_04634_),
    .B(_04630_),
    .A_N(_04633_));
 sg13g2_xnor2_1 _11757_ (.Y(_04635_),
    .A(_04630_),
    .B(_04633_));
 sg13g2_xnor2_1 _11758_ (.Y(_04636_),
    .A(net1956),
    .B(net1928));
 sg13g2_a21oi_1 _11759_ (.A1(_04615_),
    .A2(_04617_),
    .Y(_04637_),
    .B1(_04616_));
 sg13g2_nor2b_1 _11760_ (.A(_04637_),
    .B_N(_04636_),
    .Y(_04638_));
 sg13g2_xnor2_1 _11761_ (.Y(_04639_),
    .A(_04636_),
    .B(_04637_));
 sg13g2_nand2b_1 _11762_ (.Y(_04640_),
    .B(_04639_),
    .A_N(_04635_));
 sg13g2_xnor2_1 _11763_ (.Y(_04641_),
    .A(_04635_),
    .B(_04639_));
 sg13g2_o21ai_1 _11764_ (.B1(_04641_),
    .Y(_04642_),
    .A1(_04624_),
    .A2(_04626_));
 sg13g2_or3_1 _11765_ (.A(_04624_),
    .B(_04626_),
    .C(_04641_),
    .X(_04643_));
 sg13g2_and2_1 _11766_ (.A(_04642_),
    .B(_04643_),
    .X(_04644_));
 sg13g2_o21ai_1 _11767_ (.B1(_04629_),
    .Y(_00298_),
    .A1(net1554),
    .A2(_04644_));
 sg13g2_nand2_1 _11768_ (.Y(_04645_),
    .A(net1477),
    .B(net1721));
 sg13g2_and2_1 _11769_ (.A(_04640_),
    .B(_04642_),
    .X(_04646_));
 sg13g2_xnor2_1 _11770_ (.Y(_04647_),
    .A(net1901),
    .B(net1885));
 sg13g2_o21ai_1 _11771_ (.B1(_04634_),
    .Y(_04648_),
    .A1(_06865_),
    .A2(net1885));
 sg13g2_xor2_1 _11772_ (.B(_04648_),
    .A(_04647_),
    .X(_04649_));
 sg13g2_a21oi_1 _11773_ (.A1(net1956),
    .A2(_06913_),
    .Y(_04650_),
    .B1(_04638_));
 sg13g2_nand2b_1 _11774_ (.Y(_04651_),
    .B(net1954),
    .A_N(net1927));
 sg13g2_nor2b_1 _11775_ (.A(net1954),
    .B_N(net1927),
    .Y(_04652_));
 sg13g2_xnor2_1 _11776_ (.Y(_04653_),
    .A(net1954),
    .B(net1927));
 sg13g2_xnor2_1 _11777_ (.Y(_04654_),
    .A(_04650_),
    .B(_04653_));
 sg13g2_nor2b_1 _11778_ (.A(_04654_),
    .B_N(_04649_),
    .Y(_04655_));
 sg13g2_nand2b_1 _11779_ (.Y(_04656_),
    .B(_04654_),
    .A_N(_04649_));
 sg13g2_nor2b_1 _11780_ (.A(_04655_),
    .B_N(_04656_),
    .Y(_04657_));
 sg13g2_xnor2_1 _11781_ (.Y(_04658_),
    .A(_04646_),
    .B(_04657_));
 sg13g2_o21ai_1 _11782_ (.B1(_04645_),
    .Y(_00299_),
    .A1(net1554),
    .A2(_04658_));
 sg13g2_nand2_1 _11783_ (.Y(_04659_),
    .A(net1952),
    .B(net1721));
 sg13g2_nor2b_1 _11784_ (.A(net1885),
    .B_N(net1900),
    .Y(_04660_));
 sg13g2_nand2b_1 _11785_ (.Y(_04661_),
    .B(net1885),
    .A_N(net1900));
 sg13g2_nand2b_1 _11786_ (.Y(_04662_),
    .B(_04661_),
    .A_N(_04660_));
 sg13g2_nand2_1 _11787_ (.Y(_04663_),
    .A(_04630_),
    .B(_04647_));
 sg13g2_o21ai_1 _11788_ (.B1(_00546_),
    .Y(_04664_),
    .A1(net1902),
    .A2(net1901));
 sg13g2_o21ai_1 _11789_ (.B1(_04664_),
    .Y(_04665_),
    .A1(_04632_),
    .A2(_04663_));
 sg13g2_inv_1 _11790_ (.Y(_04666_),
    .A(_04665_));
 sg13g2_o21ai_1 _11791_ (.B1(_04666_),
    .Y(_04667_),
    .A1(_04631_),
    .A2(_04663_));
 sg13g2_xnor2_1 _11792_ (.Y(_04668_),
    .A(_04662_),
    .B(_04667_));
 sg13g2_nor2b_1 _11793_ (.A(net1925),
    .B_N(net1952),
    .Y(_04669_));
 sg13g2_nand2b_1 _11794_ (.Y(_04670_),
    .B(net1925),
    .A_N(net1952));
 sg13g2_nand2b_1 _11795_ (.Y(_04671_),
    .B(_04670_),
    .A_N(_04669_));
 sg13g2_o21ai_1 _11796_ (.B1(_04651_),
    .Y(_04672_),
    .A1(_04650_),
    .A2(_04652_));
 sg13g2_xnor2_1 _11797_ (.Y(_04673_),
    .A(_04671_),
    .B(_04672_));
 sg13g2_nor2b_1 _11798_ (.A(_04668_),
    .B_N(_04673_),
    .Y(_04674_));
 sg13g2_xnor2_1 _11799_ (.Y(_04675_),
    .A(_04668_),
    .B(_04673_));
 sg13g2_o21ai_1 _11800_ (.B1(_04656_),
    .Y(_04676_),
    .A1(_04646_),
    .A2(_04655_));
 sg13g2_xnor2_1 _11801_ (.Y(_04677_),
    .A(_04675_),
    .B(_04676_));
 sg13g2_o21ai_1 _11802_ (.B1(_04659_),
    .Y(_00300_),
    .A1(net1554),
    .A2(_04677_));
 sg13g2_nand2_1 _11803_ (.Y(_04678_),
    .A(net1950),
    .B(net1722));
 sg13g2_a21oi_1 _11804_ (.A1(_04675_),
    .A2(_04676_),
    .Y(_04679_),
    .B1(_04674_));
 sg13g2_a21oi_1 _11805_ (.A1(_04670_),
    .A2(_04672_),
    .Y(_04680_),
    .B1(_04669_));
 sg13g2_xnor2_1 _11806_ (.Y(_04681_),
    .A(net1950),
    .B(net1922));
 sg13g2_nand2b_1 _11807_ (.Y(_04682_),
    .B(_04681_),
    .A_N(_04680_));
 sg13g2_xnor2_1 _11808_ (.Y(_04683_),
    .A(_04680_),
    .B(_04681_));
 sg13g2_inv_1 _11809_ (.Y(_04684_),
    .A(_04683_));
 sg13g2_a21oi_1 _11810_ (.A1(_04661_),
    .A2(_04667_),
    .Y(_04685_),
    .B1(_04660_));
 sg13g2_nand2_1 _11811_ (.Y(_04686_),
    .A(net1899),
    .B(_00546_));
 sg13g2_nor2_1 _11812_ (.A(net1899),
    .B(_00546_),
    .Y(_04687_));
 sg13g2_xnor2_1 _11813_ (.Y(_04688_),
    .A(net1899),
    .B(net1885));
 sg13g2_xnor2_1 _11814_ (.Y(_04689_),
    .A(_04685_),
    .B(_04688_));
 sg13g2_xnor2_1 _11815_ (.Y(_04690_),
    .A(_04683_),
    .B(_04689_));
 sg13g2_nand2b_1 _11816_ (.Y(_04691_),
    .B(_04690_),
    .A_N(_04679_));
 sg13g2_xnor2_1 _11817_ (.Y(_04692_),
    .A(_04679_),
    .B(_04690_));
 sg13g2_inv_1 _11818_ (.Y(_04693_),
    .A(_04692_));
 sg13g2_o21ai_1 _11819_ (.B1(_04678_),
    .Y(_00301_),
    .A1(net1555),
    .A2(_04693_));
 sg13g2_nand2_1 _11820_ (.Y(_04694_),
    .A(net1469),
    .B(net1722));
 sg13g2_o21ai_1 _11821_ (.B1(_04691_),
    .Y(_04695_),
    .A1(_04684_),
    .A2(_04689_));
 sg13g2_nor2b_1 _11822_ (.A(net1885),
    .B_N(net1897),
    .Y(_04696_));
 sg13g2_nand2b_1 _11823_ (.Y(_04697_),
    .B(net1885),
    .A_N(net1897));
 sg13g2_nand2b_1 _11824_ (.Y(_04698_),
    .B(_04697_),
    .A_N(_04696_));
 sg13g2_o21ai_1 _11825_ (.B1(_04686_),
    .Y(_04699_),
    .A1(_04685_),
    .A2(_04687_));
 sg13g2_xnor2_1 _11826_ (.Y(_04700_),
    .A(_04698_),
    .B(_04699_));
 sg13g2_nor2b_1 _11827_ (.A(net1921),
    .B_N(net1948),
    .Y(_04701_));
 sg13g2_xnor2_1 _11828_ (.Y(_04702_),
    .A(net1948),
    .B(net1921));
 sg13g2_o21ai_1 _11829_ (.B1(_04682_),
    .Y(_04703_),
    .A1(_06869_),
    .A2(net1922));
 sg13g2_xor2_1 _11830_ (.B(_04703_),
    .A(_04702_),
    .X(_04704_));
 sg13g2_nor2b_1 _11831_ (.A(_04700_),
    .B_N(_04704_),
    .Y(_04705_));
 sg13g2_xnor2_1 _11832_ (.Y(_04706_),
    .A(_04700_),
    .B(_04704_));
 sg13g2_xor2_1 _11833_ (.B(_04706_),
    .A(_04695_),
    .X(_04707_));
 sg13g2_o21ai_1 _11834_ (.B1(_04694_),
    .Y(_00302_),
    .A1(net1555),
    .A2(_04707_));
 sg13g2_nand2_1 _11835_ (.Y(_04708_),
    .A(net1947),
    .B(net1722));
 sg13g2_a21oi_1 _11836_ (.A1(_04695_),
    .A2(_04706_),
    .Y(_04709_),
    .B1(_04705_));
 sg13g2_a21oi_1 _11837_ (.A1(_04697_),
    .A2(_04699_),
    .Y(_04710_),
    .B1(_04696_));
 sg13g2_xnor2_1 _11838_ (.Y(_04711_),
    .A(net1894),
    .B(_04710_));
 sg13g2_xnor2_1 _11839_ (.Y(_04712_),
    .A(_00546_),
    .B(_04711_));
 sg13g2_xnor2_1 _11840_ (.Y(_04713_),
    .A(net1947),
    .B(net1919));
 sg13g2_a21oi_1 _11841_ (.A1(_04702_),
    .A2(_04703_),
    .Y(_04714_),
    .B1(_04701_));
 sg13g2_xnor2_1 _11842_ (.Y(_04715_),
    .A(_04713_),
    .B(_04714_));
 sg13g2_nor2_1 _11843_ (.A(net1606),
    .B(_04715_),
    .Y(_04716_));
 sg13g2_nand2_1 _11844_ (.Y(_04717_),
    .A(net1606),
    .B(_04715_));
 sg13g2_nand2b_1 _11845_ (.Y(_04718_),
    .B(_04717_),
    .A_N(_04716_));
 sg13g2_xnor2_1 _11846_ (.Y(_04719_),
    .A(_04709_),
    .B(_04718_));
 sg13g2_o21ai_1 _11847_ (.B1(_04708_),
    .Y(_00303_),
    .A1(net1555),
    .A2(_04719_));
 sg13g2_nand2_1 _11848_ (.Y(_04720_),
    .A(net1449),
    .B(net1721));
 sg13g2_nand2_1 _11849_ (.Y(_04721_),
    .A(net1945),
    .B(_00557_));
 sg13g2_xor2_1 _11850_ (.B(net1916),
    .A(net1945),
    .X(_04722_));
 sg13g2_a21oi_1 _11851_ (.A1(_06873_),
    .A2(net1919),
    .Y(_04723_),
    .B1(_04714_));
 sg13g2_a21oi_2 _11852_ (.B1(_04723_),
    .Y(_04724_),
    .A2(_00553_),
    .A1(net1947));
 sg13g2_xnor2_1 _11853_ (.Y(_04725_),
    .A(_04722_),
    .B(_04724_));
 sg13g2_inv_2 _11854_ (.Y(_04726_),
    .A(_04725_));
 sg13g2_xnor2_1 _11855_ (.Y(_04727_),
    .A(net1606),
    .B(_04726_));
 sg13g2_o21ai_1 _11856_ (.B1(_04717_),
    .Y(_04728_),
    .A1(_04709_),
    .A2(_04716_));
 sg13g2_nor2b_1 _11857_ (.A(_04727_),
    .B_N(_04728_),
    .Y(_04729_));
 sg13g2_xnor2_1 _11858_ (.Y(_04730_),
    .A(_04727_),
    .B(_04728_));
 sg13g2_o21ai_1 _11859_ (.B1(_04720_),
    .Y(_00304_),
    .A1(net1554),
    .A2(_04730_));
 sg13g2_nand2_1 _11860_ (.Y(_04731_),
    .A(net1468),
    .B(net1722));
 sg13g2_a21oi_1 _11861_ (.A1(net1606),
    .A2(_04726_),
    .Y(_04732_),
    .B1(_04729_));
 sg13g2_xor2_1 _11862_ (.B(net1917),
    .A(net1943),
    .X(_04733_));
 sg13g2_o21ai_1 _11863_ (.B1(_04721_),
    .Y(_04734_),
    .A1(_04722_),
    .A2(_04724_));
 sg13g2_xnor2_1 _11864_ (.Y(_04735_),
    .A(_04733_),
    .B(_04734_));
 sg13g2_nand2_1 _11865_ (.Y(_04736_),
    .A(net1605),
    .B(_04735_));
 sg13g2_nor2_1 _11866_ (.A(net1605),
    .B(_04735_),
    .Y(_04737_));
 sg13g2_xor2_1 _11867_ (.B(_04735_),
    .A(net1605),
    .X(_04738_));
 sg13g2_xnor2_1 _11868_ (.Y(_04739_),
    .A(_04732_),
    .B(_04738_));
 sg13g2_o21ai_1 _11869_ (.B1(_04731_),
    .Y(_00305_),
    .A1(net1555),
    .A2(_04739_));
 sg13g2_nand2_1 _11870_ (.Y(_04740_),
    .A(net1941),
    .B(net1729));
 sg13g2_nor2b_1 _11871_ (.A(net1916),
    .B_N(net1941),
    .Y(_04741_));
 sg13g2_nand2b_1 _11872_ (.Y(_04742_),
    .B(net1916),
    .A_N(net1941));
 sg13g2_nand2b_1 _11873_ (.Y(_04743_),
    .B(_04742_),
    .A_N(_04741_));
 sg13g2_o21ai_1 _11874_ (.B1(_04734_),
    .Y(_04744_),
    .A1(net1943),
    .A2(_00557_));
 sg13g2_o21ai_1 _11875_ (.B1(_04744_),
    .Y(_04745_),
    .A1(_06877_),
    .A2(net1916));
 sg13g2_xnor2_1 _11876_ (.Y(_04746_),
    .A(_04743_),
    .B(_04745_));
 sg13g2_xnor2_1 _11877_ (.Y(_04747_),
    .A(net1605),
    .B(_04746_));
 sg13g2_o21ai_1 _11878_ (.B1(_04736_),
    .Y(_04748_),
    .A1(_04732_),
    .A2(_04737_));
 sg13g2_nor2b_1 _11879_ (.A(_04747_),
    .B_N(_04748_),
    .Y(_04749_));
 sg13g2_xnor2_1 _11880_ (.Y(_04750_),
    .A(_04747_),
    .B(_04748_));
 sg13g2_inv_1 _11881_ (.Y(_04751_),
    .A(_04750_));
 sg13g2_o21ai_1 _11882_ (.B1(_04740_),
    .Y(_00306_),
    .A1(net1562),
    .A2(_04751_));
 sg13g2_nand2_1 _11883_ (.Y(_04752_),
    .A(net1458),
    .B(net1729));
 sg13g2_a21oi_1 _11884_ (.A1(net1605),
    .A2(_04746_),
    .Y(_04753_),
    .B1(_04749_));
 sg13g2_a21oi_1 _11885_ (.A1(_04742_),
    .A2(_04745_),
    .Y(_04754_),
    .B1(_04741_));
 sg13g2_nand2_1 _11886_ (.Y(_04755_),
    .A(net1939),
    .B(_00557_));
 sg13g2_nor2_1 _11887_ (.A(net1939),
    .B(_00557_),
    .Y(_04756_));
 sg13g2_xnor2_1 _11888_ (.Y(_04757_),
    .A(net1939),
    .B(net1916));
 sg13g2_xnor2_1 _11889_ (.Y(_04758_),
    .A(_04754_),
    .B(_04757_));
 sg13g2_nand2_1 _11890_ (.Y(_04759_),
    .A(net1606),
    .B(_04758_));
 sg13g2_nor2_1 _11891_ (.A(net1606),
    .B(_04758_),
    .Y(_04760_));
 sg13g2_xor2_1 _11892_ (.B(_04758_),
    .A(net1605),
    .X(_04761_));
 sg13g2_xnor2_1 _11893_ (.Y(_04762_),
    .A(_04753_),
    .B(_04761_));
 sg13g2_o21ai_1 _11894_ (.B1(_04752_),
    .Y(_00307_),
    .A1(net1562),
    .A2(_04762_));
 sg13g2_nand2_1 _11895_ (.Y(_04763_),
    .A(net1937),
    .B(net1729));
 sg13g2_nor2b_1 _11896_ (.A(net1916),
    .B_N(net1937),
    .Y(_04764_));
 sg13g2_nand2b_1 _11897_ (.Y(_04765_),
    .B(net1916),
    .A_N(net1937));
 sg13g2_nand2b_1 _11898_ (.Y(_04766_),
    .B(_04765_),
    .A_N(_04764_));
 sg13g2_o21ai_1 _11899_ (.B1(_04755_),
    .Y(_04767_),
    .A1(_04754_),
    .A2(_04756_));
 sg13g2_xnor2_1 _11900_ (.Y(_04768_),
    .A(_04766_),
    .B(_04767_));
 sg13g2_xnor2_1 _11901_ (.Y(_04769_),
    .A(net1606),
    .B(_04768_));
 sg13g2_o21ai_1 _11902_ (.B1(_04759_),
    .Y(_04770_),
    .A1(_04753_),
    .A2(_04760_));
 sg13g2_nor2b_1 _11903_ (.A(_04769_),
    .B_N(_04770_),
    .Y(_04771_));
 sg13g2_xnor2_1 _11904_ (.Y(_04772_),
    .A(_04769_),
    .B(_04770_));
 sg13g2_inv_1 _11905_ (.Y(_04773_),
    .A(_04772_));
 sg13g2_o21ai_1 _11906_ (.B1(_04763_),
    .Y(_00308_),
    .A1(net1562),
    .A2(_04773_));
 sg13g2_nand2_1 _11907_ (.Y(_04774_),
    .A(net1935),
    .B(net1729));
 sg13g2_a21oi_1 _11908_ (.A1(net1605),
    .A2(_04768_),
    .Y(_04775_),
    .B1(_04771_));
 sg13g2_a21oi_1 _11909_ (.A1(_04765_),
    .A2(_04767_),
    .Y(_04776_),
    .B1(_04764_));
 sg13g2_xnor2_1 _11910_ (.Y(_04777_),
    .A(net1935),
    .B(_04776_));
 sg13g2_xnor2_1 _11911_ (.Y(_04778_),
    .A(net1917),
    .B(_04777_));
 sg13g2_inv_2 _11912_ (.Y(_04779_),
    .A(_04778_));
 sg13g2_xnor2_1 _11913_ (.Y(_04780_),
    .A(_04775_),
    .B(_04778_));
 sg13g2_xnor2_1 _11914_ (.Y(_04781_),
    .A(net1605),
    .B(_04780_));
 sg13g2_inv_2 _11915_ (.Y(_04782_),
    .A(_04781_));
 sg13g2_o21ai_1 _11916_ (.B1(_04774_),
    .Y(_00309_),
    .A1(net1561),
    .A2(net1597));
 sg13g2_nand2_1 _11917_ (.Y(_04783_),
    .A(net1475),
    .B(net1719));
 sg13g2_and2_1 _11918_ (.A(\vgadonut.donut.sAsB[6] ),
    .B(_04649_),
    .X(_04784_));
 sg13g2_xor2_1 _11919_ (.B(_04649_),
    .A(\vgadonut.donut.sAsB[6] ),
    .X(_04785_));
 sg13g2_nor2_1 _11920_ (.A(net1889),
    .B(_04635_),
    .Y(_04786_));
 sg13g2_nor2_1 _11921_ (.A(_06888_),
    .B(_04623_),
    .Y(_04787_));
 sg13g2_xnor2_1 _11922_ (.Y(_04788_),
    .A(net1890),
    .B(_04592_));
 sg13g2_xnor2_1 _11923_ (.Y(_04789_),
    .A(\vgadonut.donut.sAsB[1] ),
    .B(_04472_));
 sg13g2_nor2b_1 _11924_ (.A(_04455_),
    .B_N(_04456_),
    .Y(_04790_));
 sg13g2_xnor2_1 _11925_ (.Y(_04791_),
    .A(_04470_),
    .B(_04790_));
 sg13g2_nand2_1 _11926_ (.Y(_04792_),
    .A(net1893),
    .B(_04791_));
 sg13g2_nor2_1 _11927_ (.A(_04789_),
    .B(_04792_),
    .Y(_04793_));
 sg13g2_a21oi_1 _11928_ (.A1(net1891),
    .A2(_04472_),
    .Y(_04794_),
    .B1(_04793_));
 sg13g2_nor2_1 _11929_ (.A(_04788_),
    .B(_04794_),
    .Y(_04795_));
 sg13g2_a21oi_1 _11930_ (.A1(net1890),
    .A2(_04592_),
    .Y(_04796_),
    .B1(_04795_));
 sg13g2_xor2_1 _11931_ (.B(_04605_),
    .A(_00139_),
    .X(_04797_));
 sg13g2_nand2b_1 _11932_ (.Y(_04798_),
    .B(_04797_),
    .A_N(_04796_));
 sg13g2_o21ai_1 _11933_ (.B1(_04798_),
    .Y(_04799_),
    .A1(_00139_),
    .A2(_04605_));
 sg13g2_nand2_1 _11934_ (.Y(_04800_),
    .A(_06888_),
    .B(_04623_));
 sg13g2_nand2b_1 _11935_ (.Y(_04801_),
    .B(_04800_),
    .A_N(_04787_));
 sg13g2_a21o_1 _11936_ (.A2(_04800_),
    .A1(_04799_),
    .B1(_04787_),
    .X(_04802_));
 sg13g2_a21oi_1 _11937_ (.A1(net1889),
    .A2(_04635_),
    .Y(_04803_),
    .B1(_04802_));
 sg13g2_nor2_1 _11938_ (.A(_04786_),
    .B(_04803_),
    .Y(_04804_));
 sg13g2_xnor2_1 _11939_ (.Y(_04805_),
    .A(_04785_),
    .B(_04804_));
 sg13g2_nor2_1 _11940_ (.A(_04654_),
    .B(_04805_),
    .Y(_04806_));
 sg13g2_xnor2_1 _11941_ (.Y(_04807_),
    .A(_04654_),
    .B(_04805_));
 sg13g2_nand2_1 _11942_ (.Y(_04808_),
    .A(\vgadonut.donut.sAcB[0] ),
    .B(_04807_));
 sg13g2_xor2_1 _11943_ (.B(_04807_),
    .A(\vgadonut.donut.sAcB[0] ),
    .X(_04809_));
 sg13g2_o21ai_1 _11944_ (.B1(_04783_),
    .Y(_00310_),
    .A1(net1553),
    .A2(_04809_));
 sg13g2_nand2_1 _11945_ (.Y(_04810_),
    .A(net1453),
    .B(net1719));
 sg13g2_xnor2_1 _11946_ (.Y(_04811_),
    .A(\vgadonut.donut.sAsB[7] ),
    .B(_04668_));
 sg13g2_a21o_1 _11947_ (.A2(_04804_),
    .A1(_04785_),
    .B1(_04784_),
    .X(_04812_));
 sg13g2_nor2b_1 _11948_ (.A(_04811_),
    .B_N(_04812_),
    .Y(_04813_));
 sg13g2_xor2_1 _11949_ (.B(_04812_),
    .A(_04811_),
    .X(_04814_));
 sg13g2_and2_1 _11950_ (.A(\vgadonut.donut.sAcB[1] ),
    .B(_04814_),
    .X(_04815_));
 sg13g2_xor2_1 _11951_ (.B(_04814_),
    .A(\vgadonut.donut.sAcB[1] ),
    .X(_04816_));
 sg13g2_xor2_1 _11952_ (.B(_04816_),
    .A(_04673_),
    .X(_04817_));
 sg13g2_nand2b_1 _11953_ (.Y(_04818_),
    .B(_04817_),
    .A_N(_04806_));
 sg13g2_xnor2_1 _11954_ (.Y(_04819_),
    .A(_04806_),
    .B(_04817_));
 sg13g2_nand2b_1 _11955_ (.Y(_04820_),
    .B(_04819_),
    .A_N(_04808_));
 sg13g2_xnor2_1 _11956_ (.Y(_04821_),
    .A(_04808_),
    .B(_04819_));
 sg13g2_o21ai_1 _11957_ (.B1(_04810_),
    .Y(_00311_),
    .A1(net1553),
    .A2(_04821_));
 sg13g2_nand2_1 _11958_ (.Y(_04822_),
    .A(net1450),
    .B(net1719));
 sg13g2_nand2_1 _11959_ (.Y(_04823_),
    .A(_04818_),
    .B(_04820_));
 sg13g2_a21o_1 _11960_ (.A2(_04816_),
    .A1(_04673_),
    .B1(_04815_),
    .X(_04824_));
 sg13g2_xnor2_1 _11961_ (.Y(_04825_),
    .A(\vgadonut.donut.sAsB[8] ),
    .B(_04689_));
 sg13g2_a21oi_1 _11962_ (.A1(\vgadonut.donut.sAsB[7] ),
    .A2(_04668_),
    .Y(_04826_),
    .B1(_04813_));
 sg13g2_nor2_1 _11963_ (.A(_04825_),
    .B(_04826_),
    .Y(_04827_));
 sg13g2_xnor2_1 _11964_ (.Y(_04828_),
    .A(_04825_),
    .B(_04826_));
 sg13g2_and2_1 _11965_ (.A(\vgadonut.donut.sAcB[2] ),
    .B(_04828_),
    .X(_04829_));
 sg13g2_xor2_1 _11966_ (.B(_04828_),
    .A(\vgadonut.donut.sAcB[2] ),
    .X(_04830_));
 sg13g2_xnor2_1 _11967_ (.Y(_04831_),
    .A(_04683_),
    .B(_04830_));
 sg13g2_nor2b_1 _11968_ (.A(_04831_),
    .B_N(_04824_),
    .Y(_04832_));
 sg13g2_xor2_1 _11969_ (.B(_04831_),
    .A(_04824_),
    .X(_04833_));
 sg13g2_nor2b_1 _11970_ (.A(_04833_),
    .B_N(_04823_),
    .Y(_04834_));
 sg13g2_xnor2_1 _11971_ (.Y(_04835_),
    .A(_04823_),
    .B(_04833_));
 sg13g2_o21ai_1 _11972_ (.B1(_04822_),
    .Y(_00312_),
    .A1(net1553),
    .A2(_04835_));
 sg13g2_nand2_1 _11973_ (.Y(_04836_),
    .A(net1480),
    .B(net1720));
 sg13g2_nor2_1 _11974_ (.A(_04832_),
    .B(_04834_),
    .Y(_04837_));
 sg13g2_a21o_1 _11975_ (.A2(_04830_),
    .A1(_04683_),
    .B1(_04829_),
    .X(_04838_));
 sg13g2_a21oi_1 _11976_ (.A1(\vgadonut.donut.sAsB[8] ),
    .A2(_04689_),
    .Y(_04839_),
    .B1(_04827_));
 sg13g2_nand2_1 _11977_ (.Y(_04840_),
    .A(\vgadonut.donut.sAsB[9] ),
    .B(_04700_));
 sg13g2_nor2_1 _11978_ (.A(\vgadonut.donut.sAsB[9] ),
    .B(_04700_),
    .Y(_04841_));
 sg13g2_xnor2_1 _11979_ (.Y(_04842_),
    .A(\vgadonut.donut.sAsB[9] ),
    .B(_04700_));
 sg13g2_xnor2_1 _11980_ (.Y(_04843_),
    .A(_04839_),
    .B(_04842_));
 sg13g2_and2_1 _11981_ (.A(\vgadonut.donut.sAcB[3] ),
    .B(_04843_),
    .X(_04844_));
 sg13g2_xnor2_1 _11982_ (.Y(_04845_),
    .A(_06898_),
    .B(_04843_));
 sg13g2_xor2_1 _11983_ (.B(_04845_),
    .A(_04704_),
    .X(_04846_));
 sg13g2_nand2_1 _11984_ (.Y(_04847_),
    .A(_04838_),
    .B(_04846_));
 sg13g2_xnor2_1 _11985_ (.Y(_04848_),
    .A(_04838_),
    .B(_04846_));
 sg13g2_or2_1 _11986_ (.X(_04849_),
    .B(_04848_),
    .A(_04837_));
 sg13g2_xor2_1 _11987_ (.B(_04848_),
    .A(_04837_),
    .X(_04850_));
 sg13g2_o21ai_1 _11988_ (.B1(_04836_),
    .Y(_00313_),
    .A1(net1553),
    .A2(_04850_));
 sg13g2_nand2_1 _11989_ (.Y(_04851_),
    .A(net1457),
    .B(net1731));
 sg13g2_a21o_1 _11990_ (.A2(_04845_),
    .A1(_04704_),
    .B1(_04844_),
    .X(_04852_));
 sg13g2_xnor2_1 _11991_ (.Y(_04853_),
    .A(\vgadonut.donut.sAsB[10] ),
    .B(net1604));
 sg13g2_o21ai_1 _11992_ (.B1(_04840_),
    .Y(_04854_),
    .A1(_04839_),
    .A2(_04841_));
 sg13g2_nand2_1 _11993_ (.Y(_04855_),
    .A(_04853_),
    .B(_04854_));
 sg13g2_xnor2_1 _11994_ (.Y(_04856_),
    .A(_04853_),
    .B(_04854_));
 sg13g2_and2_1 _11995_ (.A(\vgadonut.donut.sAcB[4] ),
    .B(_04856_),
    .X(_04857_));
 sg13g2_xor2_1 _11996_ (.B(_04856_),
    .A(\vgadonut.donut.sAcB[4] ),
    .X(_04858_));
 sg13g2_xor2_1 _11997_ (.B(_04858_),
    .A(_04715_),
    .X(_04859_));
 sg13g2_and2_1 _11998_ (.A(_04852_),
    .B(_04859_),
    .X(_04860_));
 sg13g2_xnor2_1 _11999_ (.Y(_04861_),
    .A(_04852_),
    .B(_04859_));
 sg13g2_a21oi_1 _12000_ (.A1(_04847_),
    .A2(_04849_),
    .Y(_04862_),
    .B1(_04861_));
 sg13g2_nand3_1 _12001_ (.B(_04849_),
    .C(_04861_),
    .A(_04847_),
    .Y(_04863_));
 sg13g2_nor2b_1 _12002_ (.A(_04862_),
    .B_N(_04863_),
    .Y(_04864_));
 sg13g2_o21ai_1 _12003_ (.B1(_04851_),
    .Y(_00314_),
    .A1(net1564),
    .A2(_04864_));
 sg13g2_nand2_1 _12004_ (.Y(_04865_),
    .A(net1472),
    .B(net1731));
 sg13g2_a21oi_1 _12005_ (.A1(_04715_),
    .A2(_04858_),
    .Y(_04866_),
    .B1(_04857_));
 sg13g2_o21ai_1 _12006_ (.B1(_04855_),
    .Y(_04867_),
    .A1(_06903_),
    .A2(net1604));
 sg13g2_nor2b_1 _12007_ (.A(net1604),
    .B_N(net1888),
    .Y(_04868_));
 sg13g2_nand2b_1 _12008_ (.Y(_04869_),
    .B(net1604),
    .A_N(net1888));
 sg13g2_nor2b_1 _12009_ (.A(_04868_),
    .B_N(_04869_),
    .Y(_04870_));
 sg13g2_xnor2_1 _12010_ (.Y(_04871_),
    .A(_04867_),
    .B(_04870_));
 sg13g2_and2_1 _12011_ (.A(net1933),
    .B(_04871_),
    .X(_04872_));
 sg13g2_xor2_1 _12012_ (.B(_04871_),
    .A(net1933),
    .X(_04873_));
 sg13g2_xnor2_1 _12013_ (.Y(_04874_),
    .A(_04725_),
    .B(_04873_));
 sg13g2_inv_1 _12014_ (.Y(_04875_),
    .A(_04874_));
 sg13g2_xnor2_1 _12015_ (.Y(_04876_),
    .A(_04866_),
    .B(_04874_));
 sg13g2_o21ai_1 _12016_ (.B1(_04876_),
    .Y(_04877_),
    .A1(_04860_),
    .A2(_04862_));
 sg13g2_or3_1 _12017_ (.A(_04860_),
    .B(_04862_),
    .C(_04876_),
    .X(_04878_));
 sg13g2_and2_1 _12018_ (.A(_04877_),
    .B(_04878_),
    .X(_04879_));
 sg13g2_o21ai_1 _12019_ (.B1(_04865_),
    .Y(_00315_),
    .A1(net1564),
    .A2(_04879_));
 sg13g2_nand2_1 _12020_ (.Y(_04880_),
    .A(net1931),
    .B(net1720));
 sg13g2_o21ai_1 _12021_ (.B1(_04877_),
    .Y(_04881_),
    .A1(_04866_),
    .A2(_04875_));
 sg13g2_a21o_1 _12022_ (.A2(_04873_),
    .A1(_04726_),
    .B1(_04872_),
    .X(_04882_));
 sg13g2_nand2b_1 _12023_ (.Y(_04883_),
    .B(net1887),
    .A_N(net1604));
 sg13g2_nor2b_1 _12024_ (.A(net1887),
    .B_N(net1604),
    .Y(_04884_));
 sg13g2_xnor2_1 _12025_ (.Y(_04885_),
    .A(net1887),
    .B(net1604));
 sg13g2_a21oi_1 _12026_ (.A1(_04867_),
    .A2(_04869_),
    .Y(_04886_),
    .B1(_04868_));
 sg13g2_xor2_1 _12027_ (.B(_04886_),
    .A(_04885_),
    .X(_04887_));
 sg13g2_xor2_1 _12028_ (.B(_04887_),
    .A(_00108_),
    .X(_04888_));
 sg13g2_nor2b_1 _12029_ (.A(_04888_),
    .B_N(_04735_),
    .Y(_04889_));
 sg13g2_xnor2_1 _12030_ (.Y(_04890_),
    .A(_04735_),
    .B(_04888_));
 sg13g2_xnor2_1 _12031_ (.Y(_04891_),
    .A(_04882_),
    .B(_04890_));
 sg13g2_nor2b_1 _12032_ (.A(_04891_),
    .B_N(_04881_),
    .Y(_04892_));
 sg13g2_xnor2_1 _12033_ (.Y(_04893_),
    .A(_04881_),
    .B(_04891_));
 sg13g2_inv_1 _12034_ (.Y(_04894_),
    .A(_04893_));
 sg13g2_o21ai_1 _12035_ (.B1(_04880_),
    .Y(_00316_),
    .A1(net1556),
    .A2(_04894_));
 sg13g2_nand2_1 _12036_ (.Y(_04895_),
    .A(net1930),
    .B(net1720));
 sg13g2_a21o_1 _12037_ (.A2(_04890_),
    .A1(_04882_),
    .B1(_04892_),
    .X(_04896_));
 sg13g2_o21ai_1 _12038_ (.B1(_04883_),
    .Y(_04897_),
    .A1(_04884_),
    .A2(_04886_));
 sg13g2_nor2_1 _12039_ (.A(_06908_),
    .B(net1604),
    .Y(_04898_));
 sg13g2_nand2_1 _12040_ (.Y(_04899_),
    .A(_06908_),
    .B(net1607));
 sg13g2_nor2b_1 _12041_ (.A(_04898_),
    .B_N(_04899_),
    .Y(_04900_));
 sg13g2_xnor2_1 _12042_ (.Y(_04901_),
    .A(_04897_),
    .B(_04900_));
 sg13g2_xnor2_1 _12043_ (.Y(_04902_),
    .A(_00109_),
    .B(_04901_));
 sg13g2_xor2_1 _12044_ (.B(_04902_),
    .A(_04746_),
    .X(_04903_));
 sg13g2_a21o_1 _12045_ (.A2(_04887_),
    .A1(\vgadonut.donut.sAcB[6] ),
    .B1(_04889_),
    .X(_04904_));
 sg13g2_nand2_1 _12046_ (.Y(_04905_),
    .A(_04903_),
    .B(_04904_));
 sg13g2_xor2_1 _12047_ (.B(_04904_),
    .A(_04903_),
    .X(_04906_));
 sg13g2_nand2_1 _12048_ (.Y(_04907_),
    .A(_04896_),
    .B(_04906_));
 sg13g2_xnor2_1 _12049_ (.Y(_04908_),
    .A(_04896_),
    .B(_04906_));
 sg13g2_o21ai_1 _12050_ (.B1(_04895_),
    .Y(_00317_),
    .A1(net1556),
    .A2(_04908_));
 sg13g2_nand2_1 _12051_ (.Y(_04909_),
    .A(net1454),
    .B(net1719));
 sg13g2_and2_1 _12052_ (.A(net1930),
    .B(_04901_),
    .X(_04910_));
 sg13g2_a21o_1 _12053_ (.A2(_04902_),
    .A1(_04746_),
    .B1(_04910_),
    .X(_04911_));
 sg13g2_or2_1 _12054_ (.X(_04912_),
    .B(net1607),
    .A(_00140_));
 sg13g2_xnor2_1 _12055_ (.Y(_04913_),
    .A(_00140_),
    .B(net1607));
 sg13g2_a21oi_1 _12056_ (.A1(_04897_),
    .A2(_04899_),
    .Y(_04914_),
    .B1(_04898_));
 sg13g2_xor2_1 _12057_ (.B(_04914_),
    .A(_04913_),
    .X(_04915_));
 sg13g2_xnor2_1 _12058_ (.Y(_04916_),
    .A(net1929),
    .B(_04915_));
 sg13g2_nand2_1 _12059_ (.Y(_04917_),
    .A(_04758_),
    .B(_04916_));
 sg13g2_xor2_1 _12060_ (.B(_04916_),
    .A(_04758_),
    .X(_04918_));
 sg13g2_and2_1 _12061_ (.A(_04911_),
    .B(_04918_),
    .X(_04919_));
 sg13g2_xnor2_1 _12062_ (.Y(_04920_),
    .A(_04911_),
    .B(_04918_));
 sg13g2_a21oi_2 _12063_ (.B1(_04920_),
    .Y(_04921_),
    .A2(_04907_),
    .A1(_04905_));
 sg13g2_nand3_1 _12064_ (.B(_04907_),
    .C(_04920_),
    .A(_04905_),
    .Y(_04922_));
 sg13g2_nor2b_2 _12065_ (.A(_04921_),
    .B_N(_04922_),
    .Y(_04923_));
 sg13g2_o21ai_1 _12066_ (.B1(_04909_),
    .Y(_00318_),
    .A1(net1553),
    .A2(_04923_));
 sg13g2_nand2_1 _12067_ (.Y(_04924_),
    .A(net1928),
    .B(net1719));
 sg13g2_o21ai_1 _12068_ (.B1(_04912_),
    .Y(_04925_),
    .A1(_04913_),
    .A2(_04914_));
 sg13g2_xor2_1 _12069_ (.B(_04925_),
    .A(_04711_),
    .X(_04926_));
 sg13g2_xnor2_1 _12070_ (.Y(_04927_),
    .A(_00111_),
    .B(net1599));
 sg13g2_xor2_1 _12071_ (.B(_04927_),
    .A(_04768_),
    .X(_04928_));
 sg13g2_o21ai_1 _12072_ (.B1(_04917_),
    .Y(_04929_),
    .A1(_06910_),
    .A2(_04915_));
 sg13g2_nand2_1 _12073_ (.Y(_04930_),
    .A(_04928_),
    .B(_04929_));
 sg13g2_xor2_1 _12074_ (.B(_04929_),
    .A(_04928_),
    .X(_04931_));
 sg13g2_o21ai_1 _12075_ (.B1(_04931_),
    .Y(_04932_),
    .A1(_04919_),
    .A2(_04921_));
 sg13g2_or3_1 _12076_ (.A(_04919_),
    .B(_04921_),
    .C(_04931_),
    .X(_04933_));
 sg13g2_nand2_2 _12077_ (.Y(_04934_),
    .A(_04932_),
    .B(_04933_));
 sg13g2_o21ai_1 _12078_ (.B1(_04924_),
    .Y(_00319_),
    .A1(net1553),
    .A2(_04934_));
 sg13g2_nand2_1 _12079_ (.Y(_04935_),
    .A(net1452),
    .B(net1719));
 sg13g2_and2_1 _12080_ (.A(net1928),
    .B(net1599),
    .X(_04936_));
 sg13g2_a21o_1 _12081_ (.A2(_04927_),
    .A1(_04768_),
    .B1(_04936_),
    .X(_04937_));
 sg13g2_nand2_1 _12082_ (.Y(_04938_),
    .A(net1926),
    .B(net1599));
 sg13g2_xnor2_1 _12083_ (.Y(_04939_),
    .A(net1927),
    .B(net1599));
 sg13g2_xnor2_1 _12084_ (.Y(_04940_),
    .A(_04778_),
    .B(_04939_));
 sg13g2_nand2_1 _12085_ (.Y(_04941_),
    .A(_04937_),
    .B(_04940_));
 sg13g2_xnor2_1 _12086_ (.Y(_04942_),
    .A(_04937_),
    .B(_04940_));
 sg13g2_a21o_1 _12087_ (.A2(_04932_),
    .A1(_04930_),
    .B1(_04942_),
    .X(_04943_));
 sg13g2_nand3_1 _12088_ (.B(_04932_),
    .C(_04942_),
    .A(_04930_),
    .Y(_04944_));
 sg13g2_and2_2 _12089_ (.A(_04943_),
    .B(_04944_),
    .X(_04945_));
 sg13g2_o21ai_1 _12090_ (.B1(_04935_),
    .Y(_00320_),
    .A1(net1553),
    .A2(_04945_));
 sg13g2_and2_1 _12091_ (.A(net2119),
    .B(net1731),
    .X(_04946_));
 sg13g2_o21ai_1 _12092_ (.B1(_04938_),
    .Y(_04947_),
    .A1(_04779_),
    .A2(_04939_));
 sg13g2_nand2_1 _12093_ (.Y(_04948_),
    .A(net1925),
    .B(net1598));
 sg13g2_xnor2_1 _12094_ (.Y(_04949_),
    .A(net1925),
    .B(net1598));
 sg13g2_xnor2_1 _12095_ (.Y(_04950_),
    .A(_04778_),
    .B(_04949_));
 sg13g2_nand2_1 _12096_ (.Y(_04951_),
    .A(_04947_),
    .B(_04950_));
 sg13g2_xnor2_1 _12097_ (.Y(_04952_),
    .A(_04947_),
    .B(_04950_));
 sg13g2_a21o_1 _12098_ (.A2(_04943_),
    .A1(_04941_),
    .B1(_04952_),
    .X(_04953_));
 sg13g2_nand3_1 _12099_ (.B(_04943_),
    .C(_04952_),
    .A(_04941_),
    .Y(_04954_));
 sg13g2_nand2_2 _12100_ (.Y(_04955_),
    .A(_04953_),
    .B(_04954_));
 sg13g2_a21o_1 _12101_ (.A2(_04955_),
    .A1(net1571),
    .B1(_04946_),
    .X(_00321_));
 sg13g2_and2_1 _12102_ (.A(net1922),
    .B(net1731),
    .X(_04956_));
 sg13g2_xnor2_1 _12103_ (.Y(_04957_),
    .A(_00112_),
    .B(net1598));
 sg13g2_xnor2_1 _12104_ (.Y(_04958_),
    .A(_04779_),
    .B(_04957_));
 sg13g2_o21ai_1 _12105_ (.B1(_04948_),
    .Y(_04959_),
    .A1(_04779_),
    .A2(_04949_));
 sg13g2_xnor2_1 _12106_ (.Y(_04960_),
    .A(_04958_),
    .B(_04959_));
 sg13g2_a21oi_1 _12107_ (.A1(_04951_),
    .A2(_04953_),
    .Y(_04961_),
    .B1(_04960_));
 sg13g2_nand3_1 _12108_ (.B(_04953_),
    .C(_04960_),
    .A(_04951_),
    .Y(_04962_));
 sg13g2_nor2b_2 _12109_ (.A(_04961_),
    .B_N(_04962_),
    .Y(_04963_));
 sg13g2_a21o_1 _12110_ (.A2(_04963_),
    .A1(net1571),
    .B1(_04956_),
    .X(_00322_));
 sg13g2_and2_1 _12111_ (.A(net2127),
    .B(net1732),
    .X(_04964_));
 sg13g2_a21oi_1 _12112_ (.A1(_04958_),
    .A2(_04959_),
    .Y(_04965_),
    .B1(_04961_));
 sg13g2_and2_1 _12113_ (.A(net1922),
    .B(net1598),
    .X(_04966_));
 sg13g2_a21o_1 _12114_ (.A2(_04957_),
    .A1(_04778_),
    .B1(_04966_),
    .X(_04967_));
 sg13g2_nand2_1 _12115_ (.Y(_04968_),
    .A(net1921),
    .B(net1598));
 sg13g2_xnor2_1 _12116_ (.Y(_04969_),
    .A(net1921),
    .B(net1598));
 sg13g2_xnor2_1 _12117_ (.Y(_04970_),
    .A(_04779_),
    .B(_04969_));
 sg13g2_nand2b_1 _12118_ (.Y(_04971_),
    .B(_04967_),
    .A_N(_04970_));
 sg13g2_xor2_1 _12119_ (.B(_04970_),
    .A(_04967_),
    .X(_04972_));
 sg13g2_xnor2_1 _12120_ (.Y(_04973_),
    .A(_04965_),
    .B(_04972_));
 sg13g2_a21o_1 _12121_ (.A2(_04973_),
    .A1(net1571),
    .B1(_04964_),
    .X(_00323_));
 sg13g2_nand2_1 _12122_ (.Y(_04974_),
    .A(net1919),
    .B(net1733));
 sg13g2_o21ai_1 _12123_ (.B1(_04971_),
    .Y(_04975_),
    .A1(_04965_),
    .A2(_04972_));
 sg13g2_o21ai_1 _12124_ (.B1(_04968_),
    .Y(_04976_),
    .A1(_04779_),
    .A2(_04969_));
 sg13g2_xnor2_1 _12125_ (.Y(_04977_),
    .A(_00113_),
    .B(net1598));
 sg13g2_nand2_1 _12126_ (.Y(_04978_),
    .A(_04778_),
    .B(_04977_));
 sg13g2_xnor2_1 _12127_ (.Y(_04979_),
    .A(_04779_),
    .B(_04977_));
 sg13g2_xnor2_1 _12128_ (.Y(_04980_),
    .A(_04976_),
    .B(_04979_));
 sg13g2_nor2b_1 _12129_ (.A(_04980_),
    .B_N(_04975_),
    .Y(_04981_));
 sg13g2_xor2_1 _12130_ (.B(_04980_),
    .A(_04975_),
    .X(_04982_));
 sg13g2_o21ai_1 _12131_ (.B1(_04974_),
    .Y(_00324_),
    .A1(net1569),
    .A2(_04982_));
 sg13g2_nand2_1 _12132_ (.Y(_04983_),
    .A(net1918),
    .B(net1733));
 sg13g2_a21oi_1 _12133_ (.A1(_04976_),
    .A2(_04979_),
    .Y(_04984_),
    .B1(_04981_));
 sg13g2_nand2_1 _12134_ (.Y(_04985_),
    .A(_00553_),
    .B(net1598));
 sg13g2_mux2_1 _12135_ (.A0(net1599),
    .A1(_04985_),
    .S(_04978_),
    .X(_04986_));
 sg13g2_xnor2_1 _12136_ (.Y(_04987_),
    .A(_04777_),
    .B(_04986_));
 sg13g2_xnor2_1 _12137_ (.Y(_04988_),
    .A(_04984_),
    .B(_04987_));
 sg13g2_inv_1 _12138_ (.Y(_04989_),
    .A(net1547));
 sg13g2_o21ai_1 _12139_ (.B1(_04983_),
    .Y(_00325_),
    .A1(net1564),
    .A2(_04988_));
 sg13g2_nand2_1 _12140_ (.Y(_04990_),
    .A(net1915),
    .B(net1741));
 sg13g2_a21oi_1 _12141_ (.A1(net1741),
    .A2(net1773),
    .Y(_04991_),
    .B1(net1478));
 sg13g2_a21oi_1 _12142_ (.A1(net1915),
    .A2(net1741),
    .Y(_00326_),
    .B1(_04991_));
 sg13g2_xnor2_1 _12143_ (.Y(_00327_),
    .A(net2190),
    .B(_04990_));
 sg13g2_xnor2_1 _12144_ (.Y(_04992_),
    .A(_06847_),
    .B(_02971_));
 sg13g2_nand3_1 _12145_ (.B(net1771),
    .C(_04992_),
    .A(net1738),
    .Y(_04993_));
 sg13g2_o21ai_1 _12146_ (.B1(_04993_),
    .Y(_00328_),
    .A1(_06847_),
    .A2(net1738));
 sg13g2_nand3_1 _12147_ (.B(net1739),
    .C(_02971_),
    .A(net1914),
    .Y(_04994_));
 sg13g2_nand4_1 _12148_ (.B(net1914),
    .C(net1739),
    .A(net1913),
    .Y(_04995_),
    .D(_02971_));
 sg13g2_and2_1 _12149_ (.A(net1739),
    .B(net1760),
    .X(_04996_));
 sg13g2_xor2_1 _12150_ (.B(_04994_),
    .A(net1913),
    .X(_04997_));
 sg13g2_nor2_1 _12151_ (.A(_04996_),
    .B(_04997_),
    .Y(_00329_));
 sg13g2_and4_2 _12152_ (.A(net1913),
    .B(net1914),
    .C(\vgadonut.donut.v_count[4] ),
    .D(_02971_),
    .X(_04998_));
 sg13g2_nand2_1 _12153_ (.Y(_04999_),
    .A(net1738),
    .B(_04998_));
 sg13g2_a22oi_1 _12154_ (.Y(_00330_),
    .B1(_04998_),
    .B2(net1738),
    .A2(_04995_),
    .A1(_06849_));
 sg13g2_xnor2_1 _12155_ (.Y(_05000_),
    .A(net2146),
    .B(_04998_));
 sg13g2_nand3_1 _12156_ (.B(net1771),
    .C(_05000_),
    .A(net1738),
    .Y(_05001_));
 sg13g2_o21ai_1 _12157_ (.B1(_05001_),
    .Y(_00331_),
    .A1(_06848_),
    .A2(net1738));
 sg13g2_nand3_1 _12158_ (.B(net1738),
    .C(_04998_),
    .A(\vgadonut.donut.v_count[5] ),
    .Y(_05002_));
 sg13g2_nand4_1 _12159_ (.B(\vgadonut.donut.v_count[6] ),
    .C(net1738),
    .A(\vgadonut.donut.v_count[5] ),
    .Y(_05003_),
    .D(_04998_));
 sg13g2_xnor2_1 _12160_ (.Y(_00332_),
    .A(net2112),
    .B(_05002_));
 sg13g2_nor2_1 _12161_ (.A(_02977_),
    .B(_04999_),
    .Y(_05004_));
 sg13g2_xnor2_1 _12162_ (.Y(_00333_),
    .A(net2026),
    .B(_05003_));
 sg13g2_nand2_1 _12163_ (.Y(_05005_),
    .A(net2069),
    .B(_05004_));
 sg13g2_xor2_1 _12164_ (.B(_05004_),
    .A(net2069),
    .X(_00334_));
 sg13g2_xor2_1 _12165_ (.B(_05005_),
    .A(net2166),
    .X(_05006_));
 sg13g2_nor2_1 _12166_ (.A(_04996_),
    .B(_05006_),
    .Y(_00335_));
 sg13g2_nand2_1 _12167_ (.Y(_05007_),
    .A(net1986),
    .B(net1718));
 sg13g2_xnor2_1 _12168_ (.Y(_05008_),
    .A(net1912),
    .B(net1889));
 sg13g2_xnor2_1 _12169_ (.Y(_05009_),
    .A(_04677_),
    .B(_05008_));
 sg13g2_o21ai_1 _12170_ (.B1(_05007_),
    .Y(_00336_),
    .A1(net1552),
    .A2(_05009_));
 sg13g2_nand2_1 _12171_ (.Y(_05010_),
    .A(net1911),
    .B(net1718));
 sg13g2_xor2_1 _12172_ (.B(_04461_),
    .A(_04460_),
    .X(_05011_));
 sg13g2_xnor2_1 _12173_ (.Y(_05012_),
    .A(_04692_),
    .B(_05011_));
 sg13g2_nor3_1 _12174_ (.A(_04677_),
    .B(_05008_),
    .C(_05012_),
    .Y(_05013_));
 sg13g2_o21ai_1 _12175_ (.B1(_05012_),
    .Y(_05014_),
    .A1(_04677_),
    .A2(_05008_));
 sg13g2_nand2b_1 _12176_ (.Y(_05015_),
    .B(_05014_),
    .A_N(_05013_));
 sg13g2_o21ai_1 _12177_ (.B1(_05010_),
    .Y(_00337_),
    .A1(net1554),
    .A2(_05015_));
 sg13g2_nand2_1 _12178_ (.Y(_05016_),
    .A(net2028),
    .B(net1721));
 sg13g2_a21oi_1 _12179_ (.A1(_04692_),
    .A2(_05011_),
    .Y(_05017_),
    .B1(_05013_));
 sg13g2_xnor2_1 _12180_ (.Y(_05018_),
    .A(_04458_),
    .B(_04462_));
 sg13g2_nand2_1 _12181_ (.Y(_05019_),
    .A(_04707_),
    .B(_05018_));
 sg13g2_xnor2_1 _12182_ (.Y(_05020_),
    .A(_04707_),
    .B(_05018_));
 sg13g2_xnor2_1 _12183_ (.Y(_05021_),
    .A(_05017_),
    .B(_05020_));
 sg13g2_o21ai_1 _12184_ (.B1(_05016_),
    .Y(_00338_),
    .A1(net1554),
    .A2(_05021_));
 sg13g2_nand2_1 _12185_ (.Y(_05022_),
    .A(net2006),
    .B(net1721));
 sg13g2_o21ai_1 _12186_ (.B1(_05019_),
    .Y(_05023_),
    .A1(_05017_),
    .A2(_05020_));
 sg13g2_xor2_1 _12187_ (.B(_04465_),
    .A(_04464_),
    .X(_05024_));
 sg13g2_nor2_1 _12188_ (.A(_04719_),
    .B(_05024_),
    .Y(_05025_));
 sg13g2_xor2_1 _12189_ (.B(_05024_),
    .A(_04719_),
    .X(_05026_));
 sg13g2_xnor2_1 _12190_ (.Y(_05027_),
    .A(_05023_),
    .B(_05026_));
 sg13g2_o21ai_1 _12191_ (.B1(_05022_),
    .Y(_00339_),
    .A1(net1554),
    .A2(_05027_));
 sg13g2_nand2_1 _12192_ (.Y(_05028_),
    .A(net1908),
    .B(net1728));
 sg13g2_a21oi_1 _12193_ (.A1(_05023_),
    .A2(_05026_),
    .Y(_05029_),
    .B1(_05025_));
 sg13g2_xnor2_1 _12194_ (.Y(_05030_),
    .A(_04467_),
    .B(_04468_));
 sg13g2_xnor2_1 _12195_ (.Y(_05031_),
    .A(_04730_),
    .B(_05030_));
 sg13g2_nor2_1 _12196_ (.A(_05029_),
    .B(_05031_),
    .Y(_05032_));
 sg13g2_xnor2_1 _12197_ (.Y(_05033_),
    .A(_05029_),
    .B(_05031_));
 sg13g2_o21ai_1 _12198_ (.B1(_05028_),
    .Y(_00340_),
    .A1(net1561),
    .A2(_05033_));
 sg13g2_nand2_1 _12199_ (.Y(_05034_),
    .A(net1997),
    .B(net1728));
 sg13g2_a21oi_1 _12200_ (.A1(_04730_),
    .A2(_05030_),
    .Y(_05035_),
    .B1(_05032_));
 sg13g2_nor2_1 _12201_ (.A(_04739_),
    .B(_04791_),
    .Y(_05036_));
 sg13g2_nand2_1 _12202_ (.Y(_05037_),
    .A(_04739_),
    .B(_04791_));
 sg13g2_nand2b_1 _12203_ (.Y(_05038_),
    .B(_05037_),
    .A_N(_05036_));
 sg13g2_xnor2_1 _12204_ (.Y(_05039_),
    .A(_05035_),
    .B(_05038_));
 sg13g2_o21ai_1 _12205_ (.B1(_05034_),
    .Y(_00341_),
    .A1(net1561),
    .A2(_05039_));
 sg13g2_nand2_1 _12206_ (.Y(_05040_),
    .A(net1906),
    .B(net1728));
 sg13g2_and2_1 _12207_ (.A(_04472_),
    .B(_04750_),
    .X(_05041_));
 sg13g2_xor2_1 _12208_ (.B(_04750_),
    .A(_04472_),
    .X(_05042_));
 sg13g2_a21oi_1 _12209_ (.A1(_05035_),
    .A2(_05037_),
    .Y(_05043_),
    .B1(_05036_));
 sg13g2_xnor2_1 _12210_ (.Y(_05044_),
    .A(_05042_),
    .B(_05043_));
 sg13g2_o21ai_1 _12211_ (.B1(_05040_),
    .Y(_00342_),
    .A1(net1561),
    .A2(_05044_));
 sg13g2_nand2_1 _12212_ (.Y(_05045_),
    .A(net1905),
    .B(net1728));
 sg13g2_and2_1 _12213_ (.A(_04592_),
    .B(_04762_),
    .X(_05046_));
 sg13g2_xor2_1 _12214_ (.B(_04762_),
    .A(_04592_),
    .X(_05047_));
 sg13g2_a21o_1 _12215_ (.A2(_05043_),
    .A1(_05042_),
    .B1(_05041_),
    .X(_05048_));
 sg13g2_xnor2_1 _12216_ (.Y(_05049_),
    .A(_05047_),
    .B(_05048_));
 sg13g2_o21ai_1 _12217_ (.B1(_05045_),
    .Y(_00343_),
    .A1(net1561),
    .A2(_05049_));
 sg13g2_nand2_1 _12218_ (.Y(_05050_),
    .A(net1992),
    .B(net1728));
 sg13g2_a21o_1 _12219_ (.A2(_05048_),
    .A1(_05047_),
    .B1(_05046_),
    .X(_05051_));
 sg13g2_nor2_1 _12220_ (.A(_04605_),
    .B(_04773_),
    .Y(_05052_));
 sg13g2_xnor2_1 _12221_ (.Y(_05053_),
    .A(_04605_),
    .B(_04772_));
 sg13g2_xnor2_1 _12222_ (.Y(_05054_),
    .A(_05051_),
    .B(_05053_));
 sg13g2_o21ai_1 _12223_ (.B1(_05050_),
    .Y(_00344_),
    .A1(net1561),
    .A2(_05054_));
 sg13g2_nand2_1 _12224_ (.Y(_05055_),
    .A(net1995),
    .B(net1728));
 sg13g2_nor2_1 _12225_ (.A(_04623_),
    .B(net1597),
    .Y(_05056_));
 sg13g2_a21oi_1 _12226_ (.A1(_05051_),
    .A2(_05053_),
    .Y(_05057_),
    .B1(_05052_));
 sg13g2_a21oi_1 _12227_ (.A1(_04623_),
    .A2(net1597),
    .Y(_05058_),
    .B1(_05057_));
 sg13g2_xnor2_1 _12228_ (.Y(_05059_),
    .A(_04623_),
    .B(net1597));
 sg13g2_a21oi_1 _12229_ (.A1(_05057_),
    .A2(_05059_),
    .Y(_05060_),
    .B1(net1561));
 sg13g2_o21ai_1 _12230_ (.B1(_05060_),
    .Y(_05061_),
    .A1(_05057_),
    .A2(_05059_));
 sg13g2_nand2_1 _12231_ (.Y(_00345_),
    .A(_05055_),
    .B(_05061_));
 sg13g2_a21oi_1 _12232_ (.A1(net1775),
    .A2(net1764),
    .Y(_05062_),
    .B1(_06865_));
 sg13g2_nand2_1 _12233_ (.Y(_05063_),
    .A(_04635_),
    .B(_04782_));
 sg13g2_xor2_1 _12234_ (.B(net1597),
    .A(_04635_),
    .X(_05064_));
 sg13g2_nor2_1 _12235_ (.A(_05056_),
    .B(_05058_),
    .Y(_05065_));
 sg13g2_or2_1 _12236_ (.X(_05066_),
    .B(_05065_),
    .A(_05064_));
 sg13g2_a21oi_1 _12237_ (.A1(_05064_),
    .A2(_05065_),
    .Y(_05067_),
    .B1(net1562));
 sg13g2_a21o_1 _12238_ (.A2(_05067_),
    .A1(_05066_),
    .B1(_05062_),
    .X(_00346_));
 sg13g2_nand2_1 _12239_ (.Y(_05068_),
    .A(net1901),
    .B(net1728));
 sg13g2_xor2_1 _12240_ (.B(net1597),
    .A(_04649_),
    .X(_05069_));
 sg13g2_nand3_1 _12241_ (.B(_05066_),
    .C(_05069_),
    .A(_05063_),
    .Y(_05070_));
 sg13g2_a21oi_1 _12242_ (.A1(_05063_),
    .A2(_05066_),
    .Y(_05071_),
    .B1(_05069_));
 sg13g2_nand2_1 _12243_ (.Y(_05072_),
    .A(_04587_),
    .B(_05070_));
 sg13g2_o21ai_1 _12244_ (.B1(_05068_),
    .Y(_00347_),
    .A1(_05071_),
    .A2(_05072_));
 sg13g2_nand2_1 _12245_ (.Y(_05073_),
    .A(net1900),
    .B(net1729));
 sg13g2_xor2_1 _12246_ (.B(net1597),
    .A(_04668_),
    .X(_05074_));
 sg13g2_a21oi_1 _12247_ (.A1(_04649_),
    .A2(_04782_),
    .Y(_05075_),
    .B1(_05071_));
 sg13g2_nor2_1 _12248_ (.A(_05074_),
    .B(_05075_),
    .Y(_05076_));
 sg13g2_a21o_1 _12249_ (.A2(_05075_),
    .A1(_05074_),
    .B1(net1561),
    .X(_05077_));
 sg13g2_o21ai_1 _12250_ (.B1(_05073_),
    .Y(_00348_),
    .A1(_05076_),
    .A2(_05077_));
 sg13g2_nand2_1 _12251_ (.Y(_05078_),
    .A(net1899),
    .B(net1729));
 sg13g2_a21oi_1 _12252_ (.A1(_04668_),
    .A2(_04782_),
    .Y(_05079_),
    .B1(_05076_));
 sg13g2_nor2_1 _12253_ (.A(_04689_),
    .B(_04782_),
    .Y(_05080_));
 sg13g2_xor2_1 _12254_ (.B(_04781_),
    .A(_04689_),
    .X(_05081_));
 sg13g2_xnor2_1 _12255_ (.Y(_05082_),
    .A(_05079_),
    .B(_05081_));
 sg13g2_o21ai_1 _12256_ (.B1(_05078_),
    .Y(_00349_),
    .A1(_04586_),
    .A2(_05082_));
 sg13g2_nand2_1 _12257_ (.Y(_05083_),
    .A(net1897),
    .B(net1728));
 sg13g2_xor2_1 _12258_ (.B(net1597),
    .A(_04700_),
    .X(_05084_));
 sg13g2_nor2_1 _12259_ (.A(_05079_),
    .B(_05080_),
    .Y(_05085_));
 sg13g2_a21oi_1 _12260_ (.A1(_04689_),
    .A2(_04782_),
    .Y(_05086_),
    .B1(_05085_));
 sg13g2_nor2_1 _12261_ (.A(_05084_),
    .B(_05086_),
    .Y(_05087_));
 sg13g2_a21o_1 _12262_ (.A2(_05086_),
    .A1(_05084_),
    .B1(net1562),
    .X(_05088_));
 sg13g2_o21ai_1 _12263_ (.B1(_05083_),
    .Y(_00350_),
    .A1(_05087_),
    .A2(_05088_));
 sg13g2_a21oi_1 _12264_ (.A1(_04700_),
    .A2(_04782_),
    .Y(_05089_),
    .B1(_05087_));
 sg13g2_o21ai_1 _12265_ (.B1(net1571),
    .Y(_05090_),
    .A1(_04780_),
    .A2(_05089_));
 sg13g2_a21oi_1 _12266_ (.A1(_04780_),
    .A2(_05089_),
    .Y(_05091_),
    .B1(_05090_));
 sg13g2_a21o_1 _12267_ (.A2(_03930_),
    .A1(net1894),
    .B1(_05091_),
    .X(_00351_));
 sg13g2_nand2_1 _12268_ (.Y(_05092_),
    .A(net1892),
    .B(net1718));
 sg13g2_xor2_1 _12269_ (.B(_04791_),
    .A(net1893),
    .X(_05093_));
 sg13g2_xnor2_1 _12270_ (.Y(_05094_),
    .A(_04893_),
    .B(_05093_));
 sg13g2_o21ai_1 _12271_ (.B1(_05092_),
    .Y(_00352_),
    .A1(net1552),
    .A2(_05094_));
 sg13g2_nand2_1 _12272_ (.Y(_05095_),
    .A(net1891),
    .B(net1718));
 sg13g2_xor2_1 _12273_ (.B(_04792_),
    .A(_04789_),
    .X(_05096_));
 sg13g2_nand2b_1 _12274_ (.Y(_05097_),
    .B(_05096_),
    .A_N(_04908_));
 sg13g2_xnor2_1 _12275_ (.Y(_05098_),
    .A(_04908_),
    .B(_05096_));
 sg13g2_nand3_1 _12276_ (.B(_05093_),
    .C(_05098_),
    .A(_04893_),
    .Y(_05099_));
 sg13g2_a21o_1 _12277_ (.A2(_05093_),
    .A1(_04893_),
    .B1(_05098_),
    .X(_05100_));
 sg13g2_nand3_1 _12278_ (.B(_05099_),
    .C(_05100_),
    .A(net1570),
    .Y(_05101_));
 sg13g2_nand2_1 _12279_ (.Y(_00353_),
    .A(_05095_),
    .B(_05101_));
 sg13g2_nand2_1 _12280_ (.Y(_05102_),
    .A(net1989),
    .B(net1718));
 sg13g2_nand2_1 _12281_ (.Y(_05103_),
    .A(_05097_),
    .B(_05099_));
 sg13g2_xor2_1 _12282_ (.B(_04794_),
    .A(_04788_),
    .X(_05104_));
 sg13g2_nand2_1 _12283_ (.Y(_05105_),
    .A(_04923_),
    .B(_05104_));
 sg13g2_xnor2_1 _12284_ (.Y(_05106_),
    .A(_04923_),
    .B(_05104_));
 sg13g2_nand2b_1 _12285_ (.Y(_05107_),
    .B(_05103_),
    .A_N(_05106_));
 sg13g2_nand2b_1 _12286_ (.Y(_05108_),
    .B(_05106_),
    .A_N(_05103_));
 sg13g2_nand3_1 _12287_ (.B(_05107_),
    .C(_05108_),
    .A(net1570),
    .Y(_05109_));
 sg13g2_nand2_1 _12288_ (.Y(_00354_),
    .A(_05102_),
    .B(_05109_));
 sg13g2_nand2_1 _12289_ (.Y(_05110_),
    .A(net2022),
    .B(net1718));
 sg13g2_nand2_1 _12290_ (.Y(_05111_),
    .A(_05105_),
    .B(_05107_));
 sg13g2_xor2_1 _12291_ (.B(_04797_),
    .A(_04796_),
    .X(_05112_));
 sg13g2_nor2_1 _12292_ (.A(_04934_),
    .B(_05112_),
    .Y(_05113_));
 sg13g2_xor2_1 _12293_ (.B(_05112_),
    .A(_04934_),
    .X(_05114_));
 sg13g2_and2_1 _12294_ (.A(_05111_),
    .B(_05114_),
    .X(_05115_));
 sg13g2_o21ai_1 _12295_ (.B1(net1570),
    .Y(_05116_),
    .A1(_05111_),
    .A2(_05114_));
 sg13g2_o21ai_1 _12296_ (.B1(_05110_),
    .Y(_00355_),
    .A1(_05115_),
    .A2(_05116_));
 sg13g2_a21oi_1 _12297_ (.A1(net1774),
    .A2(net1761),
    .Y(_05117_),
    .B1(_06888_));
 sg13g2_nor2_1 _12298_ (.A(_05113_),
    .B(_05115_),
    .Y(_05118_));
 sg13g2_xnor2_1 _12299_ (.Y(_05119_),
    .A(_04799_),
    .B(_04801_));
 sg13g2_nand2_1 _12300_ (.Y(_05120_),
    .A(_04945_),
    .B(_05119_));
 sg13g2_xnor2_1 _12301_ (.Y(_05121_),
    .A(_04945_),
    .B(_05119_));
 sg13g2_or2_1 _12302_ (.X(_05122_),
    .B(_05121_),
    .A(_05118_));
 sg13g2_a21oi_1 _12303_ (.A1(_05118_),
    .A2(_05121_),
    .Y(_05123_),
    .B1(net1552));
 sg13g2_a21o_1 _12304_ (.A2(_05123_),
    .A1(_05122_),
    .B1(_05117_),
    .X(_00356_));
 sg13g2_and2_1 _12305_ (.A(_05120_),
    .B(_05122_),
    .X(_05124_));
 sg13g2_xor2_1 _12306_ (.B(_04635_),
    .A(net1889),
    .X(_05125_));
 sg13g2_xnor2_1 _12307_ (.Y(_05126_),
    .A(_04802_),
    .B(_05125_));
 sg13g2_nor2_1 _12308_ (.A(_04955_),
    .B(_05126_),
    .Y(_05127_));
 sg13g2_xnor2_1 _12309_ (.Y(_05128_),
    .A(_04955_),
    .B(_05126_));
 sg13g2_nor2_1 _12310_ (.A(_05124_),
    .B(_05128_),
    .Y(_05129_));
 sg13g2_a21oi_1 _12311_ (.A1(_05124_),
    .A2(_05128_),
    .Y(_05130_),
    .B1(net1553));
 sg13g2_nor2b_1 _12312_ (.A(_05129_),
    .B_N(_05130_),
    .Y(_05131_));
 sg13g2_a21o_1 _12313_ (.A2(_03930_),
    .A1(net1889),
    .B1(_05131_),
    .X(_00357_));
 sg13g2_or2_1 _12314_ (.X(_05132_),
    .B(_05129_),
    .A(_05127_));
 sg13g2_nand2b_1 _12315_ (.Y(_05133_),
    .B(_04963_),
    .A_N(_04805_));
 sg13g2_xnor2_1 _12316_ (.Y(_05134_),
    .A(_04805_),
    .B(_04963_));
 sg13g2_nand2_1 _12317_ (.Y(_05135_),
    .A(_05132_),
    .B(_05134_));
 sg13g2_o21ai_1 _12318_ (.B1(net1570),
    .Y(_05136_),
    .A1(_05132_),
    .A2(_05134_));
 sg13g2_nor2b_1 _12319_ (.A(_05136_),
    .B_N(_05135_),
    .Y(_05137_));
 sg13g2_a21o_1 _12320_ (.A2(_03930_),
    .A1(net2320),
    .B1(_05137_),
    .X(_00358_));
 sg13g2_nand2_1 _12321_ (.Y(_05138_),
    .A(net2237),
    .B(net1719));
 sg13g2_nor2_1 _12322_ (.A(_04814_),
    .B(_04973_),
    .Y(_05139_));
 sg13g2_xnor2_1 _12323_ (.Y(_05140_),
    .A(_04814_),
    .B(_04973_));
 sg13g2_a21o_1 _12324_ (.A2(_05135_),
    .A1(_05133_),
    .B1(_05140_),
    .X(_05141_));
 sg13g2_nand3_1 _12325_ (.B(_05135_),
    .C(_05140_),
    .A(_05133_),
    .Y(_05142_));
 sg13g2_nand3_1 _12326_ (.B(_05141_),
    .C(_05142_),
    .A(net1570),
    .Y(_05143_));
 sg13g2_nand2_1 _12327_ (.Y(_00359_),
    .A(_05138_),
    .B(_05143_));
 sg13g2_nand2_1 _12328_ (.Y(_05144_),
    .A(net2246),
    .B(net1720));
 sg13g2_xnor2_1 _12329_ (.Y(_05145_),
    .A(_04828_),
    .B(_04982_));
 sg13g2_nor2b_1 _12330_ (.A(_05139_),
    .B_N(_05141_),
    .Y(_05146_));
 sg13g2_nor2_1 _12331_ (.A(_05145_),
    .B(_05146_),
    .Y(_05147_));
 sg13g2_inv_1 _12332_ (.Y(_05148_),
    .A(_05147_));
 sg13g2_a21o_1 _12333_ (.A2(_05146_),
    .A1(_05145_),
    .B1(net1556),
    .X(_05149_));
 sg13g2_o21ai_1 _12334_ (.B1(_05144_),
    .Y(_00360_),
    .A1(_05147_),
    .A2(_05149_));
 sg13g2_nand2_1 _12335_ (.Y(_05150_),
    .A(net2276),
    .B(net1719));
 sg13g2_nand2_1 _12336_ (.Y(_05151_),
    .A(_04843_),
    .B(net1546));
 sg13g2_or2_1 _12337_ (.X(_05152_),
    .B(net1546),
    .A(_04843_));
 sg13g2_nand2_1 _12338_ (.Y(_05153_),
    .A(_05151_),
    .B(_05152_));
 sg13g2_o21ai_1 _12339_ (.B1(_05148_),
    .Y(_05154_),
    .A1(_04828_),
    .A2(_04982_));
 sg13g2_xor2_1 _12340_ (.B(_05154_),
    .A(_05153_),
    .X(_05155_));
 sg13g2_o21ai_1 _12341_ (.B1(_05150_),
    .Y(_00361_),
    .A1(_04586_),
    .A2(_05155_));
 sg13g2_nand2_1 _12342_ (.Y(_05156_),
    .A(net2153),
    .B(net1731));
 sg13g2_nor2_1 _12343_ (.A(_04856_),
    .B(net1546),
    .Y(_05157_));
 sg13g2_xnor2_1 _12344_ (.Y(_05158_),
    .A(_04856_),
    .B(net1546));
 sg13g2_nand2b_1 _12345_ (.Y(_05159_),
    .B(_05152_),
    .A_N(_05154_));
 sg13g2_nand2_1 _12346_ (.Y(_05160_),
    .A(_05151_),
    .B(_05159_));
 sg13g2_nor2_1 _12347_ (.A(_05158_),
    .B(_05160_),
    .Y(_05161_));
 sg13g2_a21o_1 _12348_ (.A2(_05160_),
    .A1(_05158_),
    .B1(net1564),
    .X(_05162_));
 sg13g2_o21ai_1 _12349_ (.B1(_05156_),
    .Y(_00362_),
    .A1(_05161_),
    .A2(_05162_));
 sg13g2_nand2_1 _12350_ (.Y(_05163_),
    .A(net1888),
    .B(net1731));
 sg13g2_nor2_1 _12351_ (.A(_04871_),
    .B(net1546),
    .Y(_05164_));
 sg13g2_xor2_1 _12352_ (.B(net1546),
    .A(_04871_),
    .X(_05165_));
 sg13g2_o21ai_1 _12353_ (.B1(_05165_),
    .Y(_05166_),
    .A1(_05157_),
    .A2(_05161_));
 sg13g2_or3_1 _12354_ (.A(_05157_),
    .B(_05161_),
    .C(_05165_),
    .X(_05167_));
 sg13g2_nand3_1 _12355_ (.B(_05166_),
    .C(_05167_),
    .A(net1571),
    .Y(_05168_));
 sg13g2_nand2_1 _12356_ (.Y(_00363_),
    .A(_05163_),
    .B(_05168_));
 sg13g2_nand2_1 _12357_ (.Y(_05169_),
    .A(net1887),
    .B(net1731));
 sg13g2_nor2_1 _12358_ (.A(_04887_),
    .B(net1546),
    .Y(_05170_));
 sg13g2_xor2_1 _12359_ (.B(net1546),
    .A(_04887_),
    .X(_05171_));
 sg13g2_nor2b_1 _12360_ (.A(_05164_),
    .B_N(_05166_),
    .Y(_05172_));
 sg13g2_nand2b_1 _12361_ (.Y(_05173_),
    .B(_05171_),
    .A_N(_05172_));
 sg13g2_nand2b_1 _12362_ (.Y(_05174_),
    .B(_05172_),
    .A_N(_05171_));
 sg13g2_nand3_1 _12363_ (.B(_05173_),
    .C(_05174_),
    .A(net1571),
    .Y(_05175_));
 sg13g2_nand2_1 _12364_ (.Y(_00364_),
    .A(_05169_),
    .B(_05175_));
 sg13g2_nand2_1 _12365_ (.Y(_05176_),
    .A(net2196),
    .B(net1721));
 sg13g2_nor2b_1 _12366_ (.A(_05170_),
    .B_N(_05173_),
    .Y(_05177_));
 sg13g2_nor2_1 _12367_ (.A(_04901_),
    .B(net1547),
    .Y(_05178_));
 sg13g2_xor2_1 _12368_ (.B(net1547),
    .A(_04901_),
    .X(_05179_));
 sg13g2_nand2b_1 _12369_ (.Y(_05180_),
    .B(_05179_),
    .A_N(_05177_));
 sg13g2_nand2b_1 _12370_ (.Y(_05181_),
    .B(_05177_),
    .A_N(_05179_));
 sg13g2_nand3_1 _12371_ (.B(_05180_),
    .C(_05181_),
    .A(net1570),
    .Y(_05182_));
 sg13g2_nand2_1 _12372_ (.Y(_00365_),
    .A(_05176_),
    .B(_05182_));
 sg13g2_nand2_1 _12373_ (.Y(_05183_),
    .A(net2241),
    .B(net1721));
 sg13g2_nor2b_1 _12374_ (.A(_05178_),
    .B_N(_05180_),
    .Y(_05184_));
 sg13g2_xor2_1 _12375_ (.B(net1547),
    .A(_04915_),
    .X(_05185_));
 sg13g2_or2_1 _12376_ (.X(_05186_),
    .B(_05185_),
    .A(_05184_));
 sg13g2_inv_1 _12377_ (.Y(_05187_),
    .A(_05186_));
 sg13g2_a21o_1 _12378_ (.A2(_05185_),
    .A1(_05184_),
    .B1(net1554),
    .X(_05188_));
 sg13g2_o21ai_1 _12379_ (.B1(_05183_),
    .Y(_00366_),
    .A1(_05187_),
    .A2(_05188_));
 sg13g2_a21oi_2 _12380_ (.B1(_05187_),
    .Y(_05189_),
    .A2(_04989_),
    .A1(_04915_));
 sg13g2_xnor2_1 _12381_ (.Y(_05190_),
    .A(net1599),
    .B(net1547));
 sg13g2_o21ai_1 _12382_ (.B1(net1570),
    .Y(_05191_),
    .A1(_05189_),
    .A2(_05190_));
 sg13g2_a21oi_2 _12383_ (.B1(_05191_),
    .Y(_05192_),
    .A2(_05190_),
    .A1(_05189_));
 sg13g2_a21o_1 _12384_ (.A2(_03930_),
    .A1(net1886),
    .B1(_05192_),
    .X(_00367_));
 sg13g2_nand2_1 _12385_ (.Y(_05193_),
    .A(net2005),
    .B(net1892));
 sg13g2_or2_1 _12386_ (.X(_05194_),
    .B(net1892),
    .A(\vgadonut.donut.ry6[0] ));
 sg13g2_and3_1 _12387_ (.X(_05195_),
    .A(net1742),
    .B(_05193_),
    .C(_05194_));
 sg13g2_a21oi_1 _12388_ (.A1(net1993),
    .A2(net1761),
    .Y(_05196_),
    .B1(_05195_));
 sg13g2_nand2_1 _12389_ (.Y(_05197_),
    .A(net2005),
    .B(net1649));
 sg13g2_o21ai_1 _12390_ (.B1(_05197_),
    .Y(_00368_),
    .A1(net1649),
    .A2(_05196_));
 sg13g2_xnor2_1 _12391_ (.Y(_05198_),
    .A(net1892),
    .B(net1891));
 sg13g2_inv_1 _12392_ (.Y(_05199_),
    .A(_05198_));
 sg13g2_nand2_1 _12393_ (.Y(_05200_),
    .A(net2009),
    .B(_05199_));
 sg13g2_xor2_1 _12394_ (.B(_05198_),
    .A(\vgadonut.donut.ry6[1] ),
    .X(_05201_));
 sg13g2_nand2_1 _12395_ (.Y(_05202_),
    .A(_05193_),
    .B(_05201_));
 sg13g2_or2_1 _12396_ (.X(_05203_),
    .B(_05201_),
    .A(_05193_));
 sg13g2_nor2b_1 _12397_ (.A(net1761),
    .B_N(_05203_),
    .Y(_05204_));
 sg13g2_a22oi_1 _12398_ (.Y(_05205_),
    .B1(_05202_),
    .B2(_05204_),
    .A2(net1761),
    .A1(\vgadonut.donut.ycA[1] ));
 sg13g2_nand2_1 _12399_ (.Y(_05206_),
    .A(net2009),
    .B(net1648));
 sg13g2_o21ai_1 _12400_ (.B1(_05206_),
    .Y(_00369_),
    .A1(net1648),
    .A2(_05205_));
 sg13g2_nor3_2 _12401_ (.A(net1893),
    .B(net1891),
    .C(net1890),
    .Y(_05207_));
 sg13g2_o21ai_1 _12402_ (.B1(net1890),
    .Y(_05208_),
    .A1(net1892),
    .A2(\vgadonut.donut.sAsB[1] ));
 sg13g2_nor2b_2 _12403_ (.A(_05207_),
    .B_N(_05208_),
    .Y(_05209_));
 sg13g2_nand2_1 _12404_ (.Y(_05210_),
    .A(\vgadonut.donut.ry6[2] ),
    .B(_05209_));
 sg13g2_xnor2_1 _12405_ (.Y(_05211_),
    .A(\vgadonut.donut.ry6[2] ),
    .B(_05209_));
 sg13g2_a21o_1 _12406_ (.A2(_05203_),
    .A1(_05200_),
    .B1(_05211_),
    .X(_05212_));
 sg13g2_nand3_1 _12407_ (.B(_05203_),
    .C(_05211_),
    .A(_05200_),
    .Y(_05213_));
 sg13g2_nand3_1 _12408_ (.B(_05212_),
    .C(_05213_),
    .A(net1742),
    .Y(_05214_));
 sg13g2_nor2b_1 _12409_ (.A(\vgadonut.donut.ycA[2] ),
    .B_N(net1892),
    .Y(_05215_));
 sg13g2_xor2_1 _12410_ (.B(net1892),
    .A(\vgadonut.donut.ycA[2] ),
    .X(_05216_));
 sg13g2_a21oi_1 _12411_ (.A1(net1761),
    .A2(_05216_),
    .Y(_05217_),
    .B1(net1648));
 sg13g2_a22oi_1 _12412_ (.Y(_00370_),
    .B1(_05214_),
    .B2(_05217_),
    .A2(net1648),
    .A1(_06884_));
 sg13g2_and2_1 _12413_ (.A(_06886_),
    .B(_05207_),
    .X(_05218_));
 sg13g2_xnor2_1 _12414_ (.Y(_05219_),
    .A(\vgadonut.donut.sAsB[3] ),
    .B(_05207_));
 sg13g2_inv_1 _12415_ (.Y(_05220_),
    .A(_05219_));
 sg13g2_nand2_1 _12416_ (.Y(_05221_),
    .A(\vgadonut.donut.ry6[3] ),
    .B(_05219_));
 sg13g2_xnor2_1 _12417_ (.Y(_05222_),
    .A(\vgadonut.donut.ry6[3] ),
    .B(_05219_));
 sg13g2_nand3_1 _12418_ (.B(_05212_),
    .C(_05222_),
    .A(_05210_),
    .Y(_05223_));
 sg13g2_a21o_1 _12419_ (.A2(_05212_),
    .A1(_05210_),
    .B1(_05222_),
    .X(_05224_));
 sg13g2_and2_1 _12420_ (.A(net1742),
    .B(_05223_),
    .X(_05225_));
 sg13g2_nand2_1 _12421_ (.Y(_05226_),
    .A(net1891),
    .B(_00106_));
 sg13g2_xor2_1 _12422_ (.B(_00106_),
    .A(net1891),
    .X(_05227_));
 sg13g2_xnor2_1 _12423_ (.Y(_05228_),
    .A(_05215_),
    .B(_05227_));
 sg13g2_a221oi_1 _12424_ (.B2(net1757),
    .C1(net1648),
    .B1(_05228_),
    .A1(_05224_),
    .Y(_05229_),
    .A2(_05225_));
 sg13g2_a21oi_1 _12425_ (.A1(_06887_),
    .A2(net1648),
    .Y(_00371_),
    .B1(_05229_));
 sg13g2_and2_1 _12426_ (.A(_06888_),
    .B(_05218_),
    .X(_05230_));
 sg13g2_xnor2_1 _12427_ (.Y(_05231_),
    .A(\vgadonut.donut.sAsB[4] ),
    .B(_05218_));
 sg13g2_xnor2_1 _12428_ (.Y(_05232_),
    .A(\vgadonut.donut.ry6[4] ),
    .B(_05231_));
 sg13g2_a21oi_1 _12429_ (.A1(_05221_),
    .A2(_05224_),
    .Y(_05233_),
    .B1(_05232_));
 sg13g2_and3_1 _12430_ (.X(_05234_),
    .A(_05221_),
    .B(_05224_),
    .C(_05232_));
 sg13g2_o21ai_1 _12431_ (.B1(net1742),
    .Y(_05235_),
    .A1(_05233_),
    .A2(_05234_));
 sg13g2_nand2_1 _12432_ (.Y(_05236_),
    .A(net1893),
    .B(net1890));
 sg13g2_nor2_1 _12433_ (.A(\vgadonut.donut.sAsB[1] ),
    .B(_05236_),
    .Y(_05237_));
 sg13g2_xnor2_1 _12434_ (.Y(_05238_),
    .A(net1893),
    .B(net1890));
 sg13g2_nor2_1 _12435_ (.A(\vgadonut.donut.ycA[4] ),
    .B(_05238_),
    .Y(_05239_));
 sg13g2_xor2_1 _12436_ (.B(_05238_),
    .A(\vgadonut.donut.ycA[4] ),
    .X(_05240_));
 sg13g2_nor2b_1 _12437_ (.A(_00107_),
    .B_N(\vgadonut.donut.ycA[2] ),
    .Y(_05241_));
 sg13g2_o21ai_1 _12438_ (.B1(net1892),
    .Y(_05242_),
    .A1(net1891),
    .A2(_00106_));
 sg13g2_o21ai_1 _12439_ (.B1(_05226_),
    .Y(_05243_),
    .A1(_05241_),
    .A2(_05242_));
 sg13g2_nand2_1 _12440_ (.Y(_05244_),
    .A(_05240_),
    .B(_05243_));
 sg13g2_a21oi_1 _12441_ (.A1(net1891),
    .A2(_00106_),
    .Y(_05245_),
    .B1(_05240_));
 sg13g2_xnor2_1 _12442_ (.Y(_05246_),
    .A(_05240_),
    .B(_05243_));
 sg13g2_o21ai_1 _12443_ (.B1(_05235_),
    .Y(_05247_),
    .A1(net1742),
    .A2(_05246_));
 sg13g2_nand2_1 _12444_ (.Y(_05248_),
    .A(net1998),
    .B(net1648));
 sg13g2_o21ai_1 _12445_ (.B1(_05248_),
    .Y(_00372_),
    .A1(net1648),
    .A2(_05247_));
 sg13g2_a21o_1 _12446_ (.A2(_05231_),
    .A1(\vgadonut.donut.ry6[4] ),
    .B1(_05233_),
    .X(_05249_));
 sg13g2_nor2b_1 _12447_ (.A(net1889),
    .B_N(_05230_),
    .Y(_05250_));
 sg13g2_xnor2_1 _12448_ (.Y(_05251_),
    .A(net1889),
    .B(_05230_));
 sg13g2_nand2_1 _12449_ (.Y(_05252_),
    .A(\vgadonut.donut.ry6[5] ),
    .B(net1701));
 sg13g2_xnor2_1 _12450_ (.Y(_05253_),
    .A(_06890_),
    .B(net1701));
 sg13g2_a21oi_1 _12451_ (.A1(_05249_),
    .A2(_05253_),
    .Y(_05254_),
    .B1(net1757));
 sg13g2_o21ai_1 _12452_ (.B1(_05254_),
    .Y(_05255_),
    .A1(_05249_),
    .A2(_05253_));
 sg13g2_o21ai_1 _12453_ (.B1(_05208_),
    .Y(_05256_),
    .A1(net1890),
    .A2(_05198_));
 sg13g2_xnor2_1 _12454_ (.Y(_05257_),
    .A(_06886_),
    .B(_05256_));
 sg13g2_nor2_1 _12455_ (.A(_05237_),
    .B(_05257_),
    .Y(_05258_));
 sg13g2_a21oi_1 _12456_ (.A1(_06886_),
    .A2(_05237_),
    .Y(_05259_),
    .B1(_05258_));
 sg13g2_xnor2_1 _12457_ (.Y(_05260_),
    .A(\vgadonut.donut.ycA[5] ),
    .B(_05259_));
 sg13g2_nor2_1 _12458_ (.A(_05239_),
    .B(_05260_),
    .Y(_05261_));
 sg13g2_nand2_1 _12459_ (.Y(_05262_),
    .A(_05239_),
    .B(_05260_));
 sg13g2_nand2b_1 _12460_ (.Y(_05263_),
    .B(_05262_),
    .A_N(_05261_));
 sg13g2_xnor2_1 _12461_ (.Y(_05264_),
    .A(_05244_),
    .B(_05263_));
 sg13g2_a21oi_1 _12462_ (.A1(net1761),
    .A2(_05264_),
    .Y(_05265_),
    .B1(net1649));
 sg13g2_a22oi_1 _12463_ (.Y(_00373_),
    .B1(_05255_),
    .B2(_05265_),
    .A2(net1649),
    .A1(_06890_));
 sg13g2_nor2b_1 _12464_ (.A(\vgadonut.donut.sAsB[6] ),
    .B_N(_05250_),
    .Y(_05266_));
 sg13g2_xnor2_1 _12465_ (.Y(_05267_),
    .A(\vgadonut.donut.sAsB[6] ),
    .B(_05250_));
 sg13g2_nand2_1 _12466_ (.Y(_05268_),
    .A(\vgadonut.donut.donuthit.ryin[0] ),
    .B(_05267_));
 sg13g2_xnor2_1 _12467_ (.Y(_05269_),
    .A(\vgadonut.donut.donuthit.ryin[0] ),
    .B(_05267_));
 sg13g2_o21ai_1 _12468_ (.B1(_05249_),
    .Y(_05270_),
    .A1(\vgadonut.donut.ry6[5] ),
    .A2(net1701));
 sg13g2_a21o_1 _12469_ (.A2(_05270_),
    .A1(_05252_),
    .B1(_05269_),
    .X(_05271_));
 sg13g2_nand3_1 _12470_ (.B(_05269_),
    .C(_05270_),
    .A(_05252_),
    .Y(_05272_));
 sg13g2_nand3_1 _12471_ (.B(_05271_),
    .C(_05272_),
    .A(net1742),
    .Y(_05273_));
 sg13g2_a21oi_1 _12472_ (.A1(_05245_),
    .A2(_05262_),
    .Y(_05274_),
    .B1(_05261_));
 sg13g2_nand2_1 _12473_ (.Y(_05275_),
    .A(_05264_),
    .B(_05274_));
 sg13g2_or3_1 _12474_ (.A(net1890),
    .B(_06886_),
    .C(_05198_),
    .X(_05276_));
 sg13g2_and2_1 _12475_ (.A(_06886_),
    .B(_05209_),
    .X(_05277_));
 sg13g2_nor2_1 _12476_ (.A(_05219_),
    .B(_05231_),
    .Y(_05278_));
 sg13g2_a21oi_1 _12477_ (.A1(_06888_),
    .A2(_05219_),
    .Y(_05279_),
    .B1(_05278_));
 sg13g2_xnor2_1 _12478_ (.Y(_05280_),
    .A(_00107_),
    .B(_05279_));
 sg13g2_or2_1 _12479_ (.X(_05281_),
    .B(_05280_),
    .A(_05277_));
 sg13g2_xnor2_1 _12480_ (.Y(_05282_),
    .A(_05277_),
    .B(_05280_));
 sg13g2_xor2_1 _12481_ (.B(_05282_),
    .A(\vgadonut.donut.sAcB[0] ),
    .X(_05283_));
 sg13g2_and2_1 _12482_ (.A(_05276_),
    .B(_05283_),
    .X(_05284_));
 sg13g2_xor2_1 _12483_ (.B(_05283_),
    .A(_05276_),
    .X(_05285_));
 sg13g2_xnor2_1 _12484_ (.Y(_05286_),
    .A(\vgadonut.donut.ycA[6] ),
    .B(_05285_));
 sg13g2_a21oi_1 _12485_ (.A1(\vgadonut.donut.ycA[5] ),
    .A2(_05259_),
    .Y(_05287_),
    .B1(_05258_));
 sg13g2_nor2_1 _12486_ (.A(_05286_),
    .B(_05287_),
    .Y(_05288_));
 sg13g2_xnor2_1 _12487_ (.Y(_05289_),
    .A(_05286_),
    .B(_05287_));
 sg13g2_nor2b_1 _12488_ (.A(_05289_),
    .B_N(_05275_),
    .Y(_05290_));
 sg13g2_nor2b_1 _12489_ (.A(_05275_),
    .B_N(_05289_),
    .Y(_05291_));
 sg13g2_nor3_1 _12490_ (.A(net1752),
    .B(_05290_),
    .C(_05291_),
    .Y(_05292_));
 sg13g2_nor2_1 _12491_ (.A(net1650),
    .B(_05292_),
    .Y(_05293_));
 sg13g2_a22oi_1 _12492_ (.Y(_00374_),
    .B1(_05273_),
    .B2(_05293_),
    .A2(net1650),
    .A1(_06891_));
 sg13g2_nand2_2 _12493_ (.Y(_05294_),
    .A(_06893_),
    .B(_05266_));
 sg13g2_xnor2_1 _12494_ (.Y(_05295_),
    .A(\vgadonut.donut.sAsB[7] ),
    .B(_05266_));
 sg13g2_nand2_1 _12495_ (.Y(_05296_),
    .A(\vgadonut.donut.donuthit.ryin[1] ),
    .B(_05295_));
 sg13g2_xnor2_1 _12496_ (.Y(_05297_),
    .A(\vgadonut.donut.donuthit.ryin[1] ),
    .B(_05295_));
 sg13g2_nand3_1 _12497_ (.B(_05271_),
    .C(_05297_),
    .A(_05268_),
    .Y(_05298_));
 sg13g2_a21o_1 _12498_ (.A2(_05271_),
    .A1(_05268_),
    .B1(_05297_),
    .X(_05299_));
 sg13g2_and2_1 _12499_ (.A(_05298_),
    .B(_05299_),
    .X(_05300_));
 sg13g2_a21oi_1 _12500_ (.A1(net1752),
    .A2(_05300_),
    .Y(_05301_),
    .B1(net1650));
 sg13g2_nor2_1 _12501_ (.A(_05288_),
    .B(_05290_),
    .Y(_05302_));
 sg13g2_o21ai_1 _12502_ (.B1(_05281_),
    .Y(_05303_),
    .A1(\vgadonut.donut.sAcB[0] ),
    .A2(_05282_));
 sg13g2_a21oi_1 _12503_ (.A1(_00107_),
    .A2(_05279_),
    .Y(_05304_),
    .B1(_05278_));
 sg13g2_mux2_1 _12504_ (.A0(net1701),
    .A1(net1889),
    .S(_05231_),
    .X(_05305_));
 sg13g2_nand2_1 _12505_ (.Y(_05306_),
    .A(_05198_),
    .B(_05305_));
 sg13g2_xnor2_1 _12506_ (.Y(_05307_),
    .A(_05199_),
    .B(_05305_));
 sg13g2_nand2b_1 _12507_ (.Y(_05308_),
    .B(_05307_),
    .A_N(_05304_));
 sg13g2_xnor2_1 _12508_ (.Y(_05309_),
    .A(_05304_),
    .B(_05307_));
 sg13g2_inv_1 _12509_ (.Y(_05310_),
    .A(_05309_));
 sg13g2_xnor2_1 _12510_ (.Y(_05311_),
    .A(\vgadonut.donut.sAcB[1] ),
    .B(_05309_));
 sg13g2_nand2_1 _12511_ (.Y(_05312_),
    .A(_05303_),
    .B(_05311_));
 sg13g2_xnor2_1 _12512_ (.Y(_05313_),
    .A(_05303_),
    .B(_05311_));
 sg13g2_xnor2_1 _12513_ (.Y(_05314_),
    .A(_06892_),
    .B(_05313_));
 sg13g2_a21oi_1 _12514_ (.A1(\vgadonut.donut.ycA[6] ),
    .A2(_05285_),
    .Y(_05315_),
    .B1(_05284_));
 sg13g2_and2_1 _12515_ (.A(_05314_),
    .B(_05315_),
    .X(_05316_));
 sg13g2_nor2_1 _12516_ (.A(_05314_),
    .B(_05315_),
    .Y(_05317_));
 sg13g2_or2_1 _12517_ (.X(_05318_),
    .B(_05317_),
    .A(_05316_));
 sg13g2_o21ai_1 _12518_ (.B1(net1748),
    .Y(_05319_),
    .A1(_05302_),
    .A2(_05318_));
 sg13g2_a21o_1 _12519_ (.A2(_05318_),
    .A1(_05302_),
    .B1(_05319_),
    .X(_05320_));
 sg13g2_a22oi_1 _12520_ (.Y(_00375_),
    .B1(_05301_),
    .B2(_05320_),
    .A2(net1650),
    .A1(_06894_));
 sg13g2_xnor2_1 _12521_ (.Y(_05321_),
    .A(_06896_),
    .B(_05294_));
 sg13g2_nand2_1 _12522_ (.Y(_05322_),
    .A(\vgadonut.donut.donuthit.ryin[2] ),
    .B(_05321_));
 sg13g2_xnor2_1 _12523_ (.Y(_05323_),
    .A(\vgadonut.donut.donuthit.ryin[2] ),
    .B(_05321_));
 sg13g2_a21o_1 _12524_ (.A2(_05299_),
    .A1(_05296_),
    .B1(_05323_),
    .X(_05324_));
 sg13g2_nand3_1 _12525_ (.B(_05299_),
    .C(_05323_),
    .A(_05296_),
    .Y(_05325_));
 sg13g2_nand3_1 _12526_ (.B(_05324_),
    .C(_05325_),
    .A(net1743),
    .Y(_05326_));
 sg13g2_and2_1 _12527_ (.A(net1670),
    .B(_05326_),
    .X(_05327_));
 sg13g2_o21ai_1 _12528_ (.B1(_05308_),
    .Y(_05328_),
    .A1(\vgadonut.donut.sAcB[1] ),
    .A2(_05310_));
 sg13g2_o21ai_1 _12529_ (.B1(_05306_),
    .Y(_05329_),
    .A1(_05231_),
    .A2(net1701));
 sg13g2_mux2_1 _12530_ (.A0(_05267_),
    .A1(\vgadonut.donut.sAsB[6] ),
    .S(net1701),
    .X(_05330_));
 sg13g2_nand2b_1 _12531_ (.Y(_05331_),
    .B(_05330_),
    .A_N(_05209_));
 sg13g2_xnor2_1 _12532_ (.Y(_05332_),
    .A(_05209_),
    .B(_05330_));
 sg13g2_nand2_1 _12533_ (.Y(_05333_),
    .A(_05329_),
    .B(_05332_));
 sg13g2_xnor2_1 _12534_ (.Y(_05334_),
    .A(_05329_),
    .B(_05332_));
 sg13g2_xor2_1 _12535_ (.B(_05334_),
    .A(\vgadonut.donut.sAcB[2] ),
    .X(_05335_));
 sg13g2_and2_1 _12536_ (.A(_05328_),
    .B(_05335_),
    .X(_05336_));
 sg13g2_xor2_1 _12537_ (.B(_05335_),
    .A(_05328_),
    .X(_05337_));
 sg13g2_xnor2_1 _12538_ (.Y(_05338_),
    .A(\vgadonut.donut.ycA[8] ),
    .B(_05337_));
 sg13g2_inv_1 _12539_ (.Y(_05339_),
    .A(_05338_));
 sg13g2_o21ai_1 _12540_ (.B1(_05312_),
    .Y(_05340_),
    .A1(_06892_),
    .A2(_05313_));
 sg13g2_xor2_1 _12541_ (.B(_05340_),
    .A(_05338_),
    .X(_05341_));
 sg13g2_nor3_1 _12542_ (.A(_05288_),
    .B(_05290_),
    .C(_05317_),
    .Y(_05342_));
 sg13g2_nor3_1 _12543_ (.A(_05316_),
    .B(_05341_),
    .C(_05342_),
    .Y(_05343_));
 sg13g2_o21ai_1 _12544_ (.B1(_05341_),
    .Y(_05344_),
    .A1(_05316_),
    .A2(_05342_));
 sg13g2_nand3b_1 _12545_ (.B(_05344_),
    .C(net1748),
    .Y(_05345_),
    .A_N(_05343_));
 sg13g2_a22oi_1 _12546_ (.Y(_00376_),
    .B1(_05327_),
    .B2(_05345_),
    .A2(net1653),
    .A1(_06897_));
 sg13g2_nor3_2 _12547_ (.A(\vgadonut.donut.sAsB[8] ),
    .B(\vgadonut.donut.sAsB[9] ),
    .C(_05294_),
    .Y(_05346_));
 sg13g2_o21ai_1 _12548_ (.B1(\vgadonut.donut.sAsB[9] ),
    .Y(_05347_),
    .A1(\vgadonut.donut.sAsB[8] ),
    .A2(_05294_));
 sg13g2_nor2b_2 _12549_ (.A(_05346_),
    .B_N(_05347_),
    .Y(_05348_));
 sg13g2_inv_1 _12550_ (.Y(_05349_),
    .A(_05348_));
 sg13g2_nand2_1 _12551_ (.Y(_05350_),
    .A(\vgadonut.donut.donuthit.ryin[3] ),
    .B(_05348_));
 sg13g2_xnor2_1 _12552_ (.Y(_05351_),
    .A(\vgadonut.donut.donuthit.ryin[3] ),
    .B(_05348_));
 sg13g2_a21o_1 _12553_ (.A2(_05324_),
    .A1(_05322_),
    .B1(_05351_),
    .X(_05352_));
 sg13g2_nand3_1 _12554_ (.B(_05324_),
    .C(_05351_),
    .A(_05322_),
    .Y(_05353_));
 sg13g2_nand3_1 _12555_ (.B(_05352_),
    .C(_05353_),
    .A(net1743),
    .Y(_05354_));
 sg13g2_and2_1 _12556_ (.A(net1670),
    .B(_05354_),
    .X(_05355_));
 sg13g2_a21oi_1 _12557_ (.A1(_05339_),
    .A2(_05340_),
    .Y(_05356_),
    .B1(_05343_));
 sg13g2_o21ai_1 _12558_ (.B1(_05333_),
    .Y(_05357_),
    .A1(\vgadonut.donut.sAcB[2] ),
    .A2(_05334_));
 sg13g2_o21ai_1 _12559_ (.B1(_05331_),
    .Y(_05358_),
    .A1(net1701),
    .A2(_05267_));
 sg13g2_nor2_1 _12560_ (.A(_05267_),
    .B(_05295_),
    .Y(_05359_));
 sg13g2_a21oi_1 _12561_ (.A1(_06893_),
    .A2(_05267_),
    .Y(_05360_),
    .B1(_05359_));
 sg13g2_xnor2_1 _12562_ (.Y(_05361_),
    .A(_05219_),
    .B(_05360_));
 sg13g2_nand2_1 _12563_ (.Y(_05362_),
    .A(_05358_),
    .B(_05361_));
 sg13g2_xnor2_1 _12564_ (.Y(_05363_),
    .A(_05358_),
    .B(_05361_));
 sg13g2_xnor2_1 _12565_ (.Y(_05364_),
    .A(_06898_),
    .B(_05363_));
 sg13g2_and2_1 _12566_ (.A(_05357_),
    .B(_05364_),
    .X(_05365_));
 sg13g2_xor2_1 _12567_ (.B(_05364_),
    .A(_05357_),
    .X(_05366_));
 sg13g2_xnor2_1 _12568_ (.Y(_05367_),
    .A(\vgadonut.donut.ycA[9] ),
    .B(_05366_));
 sg13g2_a21o_1 _12569_ (.A2(_05337_),
    .A1(\vgadonut.donut.ycA[8] ),
    .B1(_05336_),
    .X(_05368_));
 sg13g2_nor2b_1 _12570_ (.A(_05367_),
    .B_N(_05368_),
    .Y(_05369_));
 sg13g2_xor2_1 _12571_ (.B(_05368_),
    .A(_05367_),
    .X(_05370_));
 sg13g2_nor2_1 _12572_ (.A(_05356_),
    .B(_05370_),
    .Y(_05371_));
 sg13g2_a21oi_1 _12573_ (.A1(_05356_),
    .A2(_05370_),
    .Y(_05372_),
    .B1(net1742));
 sg13g2_nand2b_1 _12574_ (.Y(_05373_),
    .B(_05372_),
    .A_N(_05371_));
 sg13g2_a22oi_1 _12575_ (.Y(_00377_),
    .B1(_05355_),
    .B2(_05373_),
    .A2(net1653),
    .A1(_06901_));
 sg13g2_nand2_2 _12576_ (.Y(_05374_),
    .A(_06903_),
    .B(_05346_));
 sg13g2_xnor2_1 _12577_ (.Y(_05375_),
    .A(\vgadonut.donut.sAsB[10] ),
    .B(_05346_));
 sg13g2_xnor2_1 _12578_ (.Y(_05376_),
    .A(\vgadonut.donut.donuthit.ryin[4] ),
    .B(_05375_));
 sg13g2_a21oi_1 _12579_ (.A1(_05350_),
    .A2(_05352_),
    .Y(_05377_),
    .B1(_05376_));
 sg13g2_and3_1 _12580_ (.X(_05378_),
    .A(_05350_),
    .B(_05352_),
    .C(_05376_));
 sg13g2_or3_1 _12581_ (.A(net1748),
    .B(_05377_),
    .C(_05378_),
    .X(_05379_));
 sg13g2_nor2_1 _12582_ (.A(_05369_),
    .B(_05371_),
    .Y(_05380_));
 sg13g2_o21ai_1 _12583_ (.B1(_05362_),
    .Y(_05381_),
    .A1(\vgadonut.donut.sAcB[3] ),
    .A2(_05363_));
 sg13g2_a21oi_1 _12584_ (.A1(_05220_),
    .A2(_05360_),
    .Y(_05382_),
    .B1(_05359_));
 sg13g2_nor2_1 _12585_ (.A(_05295_),
    .B(_05321_),
    .Y(_05383_));
 sg13g2_a21oi_1 _12586_ (.A1(_06896_),
    .A2(_05295_),
    .Y(_05384_),
    .B1(_05383_));
 sg13g2_nand2b_1 _12587_ (.Y(_05385_),
    .B(_05384_),
    .A_N(_05231_));
 sg13g2_xnor2_1 _12588_ (.Y(_05386_),
    .A(_05231_),
    .B(_05384_));
 sg13g2_nand2b_1 _12589_ (.Y(_05387_),
    .B(_05386_),
    .A_N(_05382_));
 sg13g2_xnor2_1 _12590_ (.Y(_05388_),
    .A(_05382_),
    .B(_05386_));
 sg13g2_inv_1 _12591_ (.Y(_05389_),
    .A(_05388_));
 sg13g2_xnor2_1 _12592_ (.Y(_05390_),
    .A(net1934),
    .B(_05388_));
 sg13g2_nand2_1 _12593_ (.Y(_05391_),
    .A(_05381_),
    .B(_05390_));
 sg13g2_xnor2_1 _12594_ (.Y(_05392_),
    .A(_05381_),
    .B(_05390_));
 sg13g2_xnor2_1 _12595_ (.Y(_05393_),
    .A(_06902_),
    .B(_05392_));
 sg13g2_a21o_1 _12596_ (.A2(_05366_),
    .A1(\vgadonut.donut.ycA[9] ),
    .B1(_05365_),
    .X(_05394_));
 sg13g2_nand2b_1 _12597_ (.Y(_05395_),
    .B(_05394_),
    .A_N(_05393_));
 sg13g2_xor2_1 _12598_ (.B(_05394_),
    .A(_05393_),
    .X(_05396_));
 sg13g2_or2_1 _12599_ (.X(_05397_),
    .B(_05396_),
    .A(_05380_));
 sg13g2_a21oi_1 _12600_ (.A1(_05380_),
    .A2(_05396_),
    .Y(_05398_),
    .B1(net1752));
 sg13g2_a21oi_1 _12601_ (.A1(_05397_),
    .A2(_05398_),
    .Y(_05399_),
    .B1(net1653));
 sg13g2_a22oi_1 _12602_ (.Y(_00378_),
    .B1(_05379_),
    .B2(_05399_),
    .A2(net1653),
    .A1(_06904_));
 sg13g2_o21ai_1 _12603_ (.B1(_05391_),
    .Y(_05400_),
    .A1(_06902_),
    .A2(_05392_));
 sg13g2_o21ai_1 _12604_ (.B1(_05387_),
    .Y(_05401_),
    .A1(net1934),
    .A2(_05389_));
 sg13g2_nand2b_1 _12605_ (.Y(_05402_),
    .B(_05385_),
    .A_N(_05383_));
 sg13g2_or2_1 _12606_ (.X(_05403_),
    .B(_05348_),
    .A(_05321_));
 sg13g2_nand2_1 _12607_ (.Y(_05404_),
    .A(_06900_),
    .B(_05321_));
 sg13g2_nand2_1 _12608_ (.Y(_05405_),
    .A(_05403_),
    .B(_05404_));
 sg13g2_xor2_1 _12609_ (.B(_05405_),
    .A(_05251_),
    .X(_05406_));
 sg13g2_nand2_1 _12610_ (.Y(_05407_),
    .A(_05402_),
    .B(_05406_));
 sg13g2_xnor2_1 _12611_ (.Y(_05408_),
    .A(_05402_),
    .B(_05406_));
 sg13g2_xor2_1 _12612_ (.B(_05408_),
    .A(net1932),
    .X(_05409_));
 sg13g2_and2_1 _12613_ (.A(_05401_),
    .B(_05409_),
    .X(_05410_));
 sg13g2_xor2_1 _12614_ (.B(_05409_),
    .A(_05401_),
    .X(_05411_));
 sg13g2_xnor2_1 _12615_ (.Y(_05412_),
    .A(\vgadonut.donut.ycA[11] ),
    .B(_05411_));
 sg13g2_inv_1 _12616_ (.Y(_05413_),
    .A(_05412_));
 sg13g2_xor2_1 _12617_ (.B(_05412_),
    .A(_05400_),
    .X(_05414_));
 sg13g2_and3_1 _12618_ (.X(_05415_),
    .A(_05395_),
    .B(_05397_),
    .C(_05414_));
 sg13g2_a21oi_1 _12619_ (.A1(_05395_),
    .A2(_05397_),
    .Y(_05416_),
    .B1(_05414_));
 sg13g2_a21o_1 _12620_ (.A2(_05375_),
    .A1(\vgadonut.donut.donuthit.ryin[4] ),
    .B1(_05377_),
    .X(_05417_));
 sg13g2_xor2_1 _12621_ (.B(_05374_),
    .A(net1888),
    .X(_05418_));
 sg13g2_nand2_1 _12622_ (.Y(_05419_),
    .A(\vgadonut.donut.donuthit.ryin[5] ),
    .B(net1619));
 sg13g2_xnor2_1 _12623_ (.Y(_05420_),
    .A(_06906_),
    .B(net1619));
 sg13g2_o21ai_1 _12624_ (.B1(net1757),
    .Y(_05421_),
    .A1(_05415_),
    .A2(_05416_));
 sg13g2_xnor2_1 _12625_ (.Y(_05422_),
    .A(_05417_),
    .B(_05420_));
 sg13g2_a21oi_1 _12626_ (.A1(net1745),
    .A2(_05422_),
    .Y(_05423_),
    .B1(net1653));
 sg13g2_nand2_1 _12627_ (.Y(_05424_),
    .A(_05421_),
    .B(_05423_));
 sg13g2_o21ai_1 _12628_ (.B1(_05424_),
    .Y(_00379_),
    .A1(_06906_),
    .A2(net1670));
 sg13g2_o21ai_1 _12629_ (.B1(_05417_),
    .Y(_05425_),
    .A1(\vgadonut.donut.donuthit.ryin[5] ),
    .A2(net1619));
 sg13g2_nor3_2 _12630_ (.A(net1888),
    .B(net1887),
    .C(_05374_),
    .Y(_05426_));
 sg13g2_o21ai_1 _12631_ (.B1(net1887),
    .Y(_05427_),
    .A1(net1888),
    .A2(_05374_));
 sg13g2_nor2b_2 _12632_ (.A(_05426_),
    .B_N(_05427_),
    .Y(_05428_));
 sg13g2_xnor2_1 _12633_ (.Y(_05429_),
    .A(\vgadonut.donut.donuthit.ryin[6] ),
    .B(_05428_));
 sg13g2_a21oi_1 _12634_ (.A1(_05419_),
    .A2(_05425_),
    .Y(_05430_),
    .B1(_05429_));
 sg13g2_nand3_1 _12635_ (.B(_05425_),
    .C(_05429_),
    .A(_05419_),
    .Y(_05431_));
 sg13g2_nor2b_1 _12636_ (.A(_05430_),
    .B_N(_05431_),
    .Y(_05432_));
 sg13g2_a21oi_1 _12637_ (.A1(net1752),
    .A2(_05432_),
    .Y(_05433_),
    .B1(net1660));
 sg13g2_a21oi_1 _12638_ (.A1(_05400_),
    .A2(_05413_),
    .Y(_05434_),
    .B1(_05416_));
 sg13g2_o21ai_1 _12639_ (.B1(_05407_),
    .Y(_05435_),
    .A1(net1932),
    .A2(_05408_));
 sg13g2_o21ai_1 _12640_ (.B1(_05403_),
    .Y(_05436_),
    .A1(net1701),
    .A2(_05405_));
 sg13g2_nor2_1 _12641_ (.A(_05348_),
    .B(_05375_),
    .Y(_05437_));
 sg13g2_a21oi_1 _12642_ (.A1(_06903_),
    .A2(_05348_),
    .Y(_05438_),
    .B1(_05437_));
 sg13g2_nand2b_1 _12643_ (.Y(_05439_),
    .B(_05438_),
    .A_N(_05267_));
 sg13g2_xnor2_1 _12644_ (.Y(_05440_),
    .A(_05267_),
    .B(_05438_));
 sg13g2_and2_1 _12645_ (.A(_05436_),
    .B(_05440_),
    .X(_05441_));
 sg13g2_xor2_1 _12646_ (.B(_05440_),
    .A(_05436_),
    .X(_05442_));
 sg13g2_xnor2_1 _12647_ (.Y(_05443_),
    .A(_00108_),
    .B(_05442_));
 sg13g2_nand2b_1 _12648_ (.Y(_05444_),
    .B(_05435_),
    .A_N(_05443_));
 sg13g2_xor2_1 _12649_ (.B(_05443_),
    .A(_05435_),
    .X(_05445_));
 sg13g2_inv_1 _12650_ (.Y(_05446_),
    .A(_05445_));
 sg13g2_nand2_1 _12651_ (.Y(_05447_),
    .A(\vgadonut.donut.ycA[12] ),
    .B(_05446_));
 sg13g2_xor2_1 _12652_ (.B(_05445_),
    .A(\vgadonut.donut.ycA[12] ),
    .X(_05448_));
 sg13g2_a21o_1 _12653_ (.A2(_05411_),
    .A1(\vgadonut.donut.ycA[11] ),
    .B1(_05410_),
    .X(_05449_));
 sg13g2_inv_1 _12654_ (.Y(_05450_),
    .A(_05449_));
 sg13g2_xor2_1 _12655_ (.B(_05449_),
    .A(_05448_),
    .X(_05451_));
 sg13g2_or2_1 _12656_ (.X(_05452_),
    .B(_05451_),
    .A(_05434_));
 sg13g2_a21oi_1 _12657_ (.A1(_05434_),
    .A2(_05451_),
    .Y(_05453_),
    .B1(net1743));
 sg13g2_nand2_2 _12658_ (.Y(_05454_),
    .A(_05452_),
    .B(_05453_));
 sg13g2_a22oi_1 _12659_ (.Y(_00380_),
    .B1(_05433_),
    .B2(_05454_),
    .A2(net1660),
    .A1(_06907_));
 sg13g2_o21ai_1 _12660_ (.B1(_05452_),
    .Y(_05455_),
    .A1(_05448_),
    .A2(_05450_));
 sg13g2_a21o_1 _12661_ (.A2(_05442_),
    .A1(_00108_),
    .B1(_05441_),
    .X(_05456_));
 sg13g2_nand2b_1 _12662_ (.Y(_05457_),
    .B(_05439_),
    .A_N(_05437_));
 sg13g2_mux2_1 _12663_ (.A0(net1619),
    .A1(net1888),
    .S(_05375_),
    .X(_05458_));
 sg13g2_nand2b_1 _12664_ (.Y(_05459_),
    .B(_05458_),
    .A_N(_05295_));
 sg13g2_xnor2_1 _12665_ (.Y(_05460_),
    .A(_05295_),
    .B(_05458_));
 sg13g2_xor2_1 _12666_ (.B(_05460_),
    .A(_05457_),
    .X(_05461_));
 sg13g2_and2_1 _12667_ (.A(_00109_),
    .B(_05461_),
    .X(_05462_));
 sg13g2_xnor2_1 _12668_ (.Y(_05463_),
    .A(_00109_),
    .B(_05461_));
 sg13g2_nor2b_1 _12669_ (.A(_05463_),
    .B_N(_05456_),
    .Y(_05464_));
 sg13g2_xnor2_1 _12670_ (.Y(_05465_),
    .A(_05456_),
    .B(_05463_));
 sg13g2_xnor2_1 _12671_ (.Y(_05466_),
    .A(\vgadonut.donut.ycA[13] ),
    .B(_05465_));
 sg13g2_nand3_1 _12672_ (.B(_05447_),
    .C(_05466_),
    .A(_05444_),
    .Y(_05467_));
 sg13g2_inv_1 _12673_ (.Y(_05468_),
    .A(_05467_));
 sg13g2_a21oi_1 _12674_ (.A1(_05444_),
    .A2(_05447_),
    .Y(_05469_),
    .B1(_05466_));
 sg13g2_nor2_1 _12675_ (.A(_05468_),
    .B(_05469_),
    .Y(_05470_));
 sg13g2_a21oi_1 _12676_ (.A1(_06909_),
    .A2(_05428_),
    .Y(_05471_),
    .B1(_05430_));
 sg13g2_nand2_1 _12677_ (.Y(_05472_),
    .A(_06908_),
    .B(_05426_));
 sg13g2_xnor2_1 _12678_ (.Y(_05473_),
    .A(\vgadonut.donut.sAsB[13] ),
    .B(_05426_));
 sg13g2_nor2_1 _12679_ (.A(\vgadonut.donut.donuthit.ryin[7] ),
    .B(_05473_),
    .Y(_05474_));
 sg13g2_nand2_1 _12680_ (.Y(_05475_),
    .A(\vgadonut.donut.donuthit.ryin[7] ),
    .B(_05473_));
 sg13g2_nand2b_1 _12681_ (.Y(_05476_),
    .B(_05475_),
    .A_N(_05474_));
 sg13g2_xnor2_1 _12682_ (.Y(_05477_),
    .A(_05471_),
    .B(_05476_));
 sg13g2_xnor2_1 _12683_ (.Y(_05478_),
    .A(_05455_),
    .B(_05470_));
 sg13g2_a221oi_1 _12684_ (.B2(net1759),
    .C1(net1659),
    .B1(_05478_),
    .A1(net1745),
    .Y(_05479_),
    .A2(_05477_));
 sg13g2_a21o_1 _12685_ (.A2(net1658),
    .A1(net2282),
    .B1(_05479_),
    .X(_00381_));
 sg13g2_nor2_1 _12686_ (.A(\vgadonut.donut.sAsB[14] ),
    .B(_05472_),
    .Y(_05480_));
 sg13g2_xor2_1 _12687_ (.B(_05472_),
    .A(\vgadonut.donut.sAsB[14] ),
    .X(_05481_));
 sg13g2_xnor2_1 _12688_ (.Y(_05482_),
    .A(\vgadonut.donut.donuthit.ryin[8] ),
    .B(_05481_));
 sg13g2_or2_1 _12689_ (.X(_05483_),
    .B(_05474_),
    .A(_05471_));
 sg13g2_a21oi_1 _12690_ (.A1(_05475_),
    .A2(_05483_),
    .Y(_05484_),
    .B1(_05482_));
 sg13g2_and3_1 _12691_ (.X(_05485_),
    .A(_05475_),
    .B(_05482_),
    .C(_05483_));
 sg13g2_nor3_1 _12692_ (.A(_03931_),
    .B(_05484_),
    .C(_05485_),
    .Y(_05486_));
 sg13g2_nor2_1 _12693_ (.A(net1660),
    .B(_05486_),
    .Y(_05487_));
 sg13g2_a21oi_2 _12694_ (.B1(_05462_),
    .Y(_05488_),
    .A2(_05460_),
    .A1(_05457_));
 sg13g2_o21ai_1 _12695_ (.B1(_05459_),
    .Y(_05489_),
    .A1(_05375_),
    .A2(net1619));
 sg13g2_nor2_1 _12696_ (.A(net1619),
    .B(_05428_),
    .Y(_05490_));
 sg13g2_or2_1 _12697_ (.X(_05491_),
    .B(_05428_),
    .A(net1619));
 sg13g2_nor2b_1 _12698_ (.A(net1887),
    .B_N(net1619),
    .Y(_05492_));
 sg13g2_nor2_1 _12699_ (.A(_05490_),
    .B(_05492_),
    .Y(_05493_));
 sg13g2_xnor2_1 _12700_ (.Y(_05494_),
    .A(_05321_),
    .B(_05493_));
 sg13g2_nand2_1 _12701_ (.Y(_05495_),
    .A(_05489_),
    .B(_05494_));
 sg13g2_xnor2_1 _12702_ (.Y(_05496_),
    .A(_05489_),
    .B(_05494_));
 sg13g2_xnor2_1 _12703_ (.Y(_05497_),
    .A(_06910_),
    .B(_05496_));
 sg13g2_nor2b_1 _12704_ (.A(_05488_),
    .B_N(_05497_),
    .Y(_05498_));
 sg13g2_xnor2_1 _12705_ (.Y(_05499_),
    .A(_05488_),
    .B(_05497_));
 sg13g2_xnor2_1 _12706_ (.Y(_05500_),
    .A(\vgadonut.donut.ycA[14] ),
    .B(_05499_));
 sg13g2_a21oi_2 _12707_ (.B1(_05464_),
    .Y(_05501_),
    .A2(_05465_),
    .A1(\vgadonut.donut.ycA[13] ));
 sg13g2_nor2_1 _12708_ (.A(_05500_),
    .B(_05501_),
    .Y(_05502_));
 sg13g2_xnor2_1 _12709_ (.Y(_05503_),
    .A(_05500_),
    .B(_05501_));
 sg13g2_a21oi_2 _12710_ (.B1(_05469_),
    .Y(_05504_),
    .A2(_05467_),
    .A1(_05455_));
 sg13g2_nor2_1 _12711_ (.A(_05503_),
    .B(_05504_),
    .Y(_05505_));
 sg13g2_a21oi_1 _12712_ (.A1(_05503_),
    .A2(_05504_),
    .Y(_05506_),
    .B1(net1743));
 sg13g2_nand2b_1 _12713_ (.Y(_05507_),
    .B(_05506_),
    .A_N(_05505_));
 sg13g2_a22oi_1 _12714_ (.Y(_00382_),
    .B1(_05487_),
    .B2(_05507_),
    .A2(net1660),
    .A1(_06912_));
 sg13g2_xnor2_1 _12715_ (.Y(_05508_),
    .A(net1886),
    .B(_05480_));
 sg13g2_xnor2_1 _12716_ (.Y(_05509_),
    .A(\vgadonut.donut.donuthit.ryin[9] ),
    .B(net1614));
 sg13g2_a21oi_2 _12717_ (.B1(_05484_),
    .Y(_05510_),
    .A2(_05481_),
    .A1(\vgadonut.donut.donuthit.ryin[8] ));
 sg13g2_nor2_1 _12718_ (.A(_05509_),
    .B(_05510_),
    .Y(_05511_));
 sg13g2_a221oi_1 _12719_ (.B2(_05510_),
    .C1(_05511_),
    .B1(_05509_),
    .A1(_02946_),
    .Y(_05512_),
    .A2(_03914_));
 sg13g2_nor2_1 _12720_ (.A(net1656),
    .B(_05512_),
    .Y(_05513_));
 sg13g2_nor2_1 _12721_ (.A(_05502_),
    .B(_05505_),
    .Y(_05514_));
 sg13g2_o21ai_1 _12722_ (.B1(_05495_),
    .Y(_05515_),
    .A1(\vgadonut.donut.sAcB[8] ),
    .A2(_05496_));
 sg13g2_o21ai_1 _12723_ (.B1(_05491_),
    .Y(_05516_),
    .A1(_05321_),
    .A2(_05492_));
 sg13g2_nor2_1 _12724_ (.A(_05428_),
    .B(_05473_),
    .Y(_05517_));
 sg13g2_a21oi_1 _12725_ (.A1(_06908_),
    .A2(_05428_),
    .Y(_05518_),
    .B1(_05517_));
 sg13g2_xnor2_1 _12726_ (.Y(_05519_),
    .A(_05348_),
    .B(_05518_));
 sg13g2_and2_1 _12727_ (.A(_05516_),
    .B(_05519_),
    .X(_05520_));
 sg13g2_xor2_1 _12728_ (.B(_05519_),
    .A(_05516_),
    .X(_05521_));
 sg13g2_xnor2_1 _12729_ (.Y(_05522_),
    .A(_00111_),
    .B(_05521_));
 sg13g2_nor2b_1 _12730_ (.A(_05522_),
    .B_N(_05515_),
    .Y(_05523_));
 sg13g2_xor2_1 _12731_ (.B(_05522_),
    .A(_05515_),
    .X(_05524_));
 sg13g2_inv_1 _12732_ (.Y(_05525_),
    .A(_05524_));
 sg13g2_xnor2_1 _12733_ (.Y(_05526_),
    .A(_06914_),
    .B(_05524_));
 sg13g2_a21oi_1 _12734_ (.A1(\vgadonut.donut.ycA[14] ),
    .A2(_05499_),
    .Y(_05527_),
    .B1(_05498_));
 sg13g2_nor2_1 _12735_ (.A(_05526_),
    .B(_05527_),
    .Y(_05528_));
 sg13g2_xnor2_1 _12736_ (.Y(_05529_),
    .A(_05526_),
    .B(_05527_));
 sg13g2_nor2_1 _12737_ (.A(_05514_),
    .B(_05529_),
    .Y(_05530_));
 sg13g2_a21oi_1 _12738_ (.A1(_05514_),
    .A2(_05529_),
    .Y(_05531_),
    .B1(net1745));
 sg13g2_nand2b_1 _12739_ (.Y(_05532_),
    .B(_05531_),
    .A_N(_05530_));
 sg13g2_a22oi_1 _12740_ (.Y(_00383_),
    .B1(_05513_),
    .B2(_05532_),
    .A2(net1656),
    .A1(_00547_));
 sg13g2_xnor2_1 _12741_ (.Y(_05533_),
    .A(_00549_),
    .B(net1614));
 sg13g2_a21oi_1 _12742_ (.A1(\vgadonut.donut.donuthit.ryin[9] ),
    .A2(net1614),
    .Y(_05534_),
    .B1(_05511_));
 sg13g2_nor2b_1 _12743_ (.A(_05534_),
    .B_N(_05533_),
    .Y(_05535_));
 sg13g2_xnor2_1 _12744_ (.Y(_05536_),
    .A(_05533_),
    .B(_05534_));
 sg13g2_a21oi_1 _12745_ (.A1(net1756),
    .A2(_05536_),
    .Y(_05537_),
    .B1(net1668));
 sg13g2_nor2_1 _12746_ (.A(_05528_),
    .B(_05530_),
    .Y(_05538_));
 sg13g2_a21oi_1 _12747_ (.A1(_00111_),
    .A2(_05521_),
    .Y(_05539_),
    .B1(_05520_));
 sg13g2_a21oi_1 _12748_ (.A1(_05349_),
    .A2(_05518_),
    .Y(_05540_),
    .B1(_05517_));
 sg13g2_mux2_1 _12749_ (.A0(_05481_),
    .A1(\vgadonut.donut.sAsB[14] ),
    .S(_05473_),
    .X(_05541_));
 sg13g2_nand2b_1 _12750_ (.Y(_05542_),
    .B(_05541_),
    .A_N(_05375_));
 sg13g2_xnor2_1 _12751_ (.Y(_05543_),
    .A(_05375_),
    .B(_05541_));
 sg13g2_nand2b_1 _12752_ (.Y(_05544_),
    .B(_05543_),
    .A_N(_05540_));
 sg13g2_xnor2_1 _12753_ (.Y(_05545_),
    .A(_05540_),
    .B(_05543_));
 sg13g2_inv_1 _12754_ (.Y(_05546_),
    .A(_05545_));
 sg13g2_xnor2_1 _12755_ (.Y(_05547_),
    .A(net1926),
    .B(_05545_));
 sg13g2_nor2b_1 _12756_ (.A(_05539_),
    .B_N(_05547_),
    .Y(_05548_));
 sg13g2_xnor2_1 _12757_ (.Y(_05549_),
    .A(_05539_),
    .B(_05547_));
 sg13g2_xnor2_1 _12758_ (.Y(_05550_),
    .A(\vgadonut.donut.ycA[16] ),
    .B(_05549_));
 sg13g2_a21oi_1 _12759_ (.A1(\vgadonut.donut.ycA[15] ),
    .A2(_05525_),
    .Y(_05551_),
    .B1(_05523_));
 sg13g2_xnor2_1 _12760_ (.Y(_05552_),
    .A(_05550_),
    .B(_05551_));
 sg13g2_or2_1 _12761_ (.X(_05553_),
    .B(_05552_),
    .A(_05538_));
 sg13g2_a21oi_1 _12762_ (.A1(_05538_),
    .A2(_05552_),
    .Y(_05554_),
    .B1(net1746));
 sg13g2_nand2_1 _12763_ (.Y(_05555_),
    .A(_05553_),
    .B(_05554_));
 sg13g2_a22oi_1 _12764_ (.Y(_00384_),
    .B1(_05537_),
    .B2(_05555_),
    .A2(net1668),
    .A1(_00549_));
 sg13g2_o21ai_1 _12765_ (.B1(_05553_),
    .Y(_05556_),
    .A1(_05550_),
    .A2(_05551_));
 sg13g2_a21oi_1 _12766_ (.A1(\vgadonut.donut.ycA[16] ),
    .A2(_05549_),
    .Y(_05557_),
    .B1(_05548_));
 sg13g2_o21ai_1 _12767_ (.B1(_05544_),
    .Y(_05558_),
    .A1(net1926),
    .A2(_05546_));
 sg13g2_nor2_1 _12768_ (.A(_05481_),
    .B(net1614),
    .Y(_05559_));
 sg13g2_a21oi_2 _12769_ (.B1(_05559_),
    .Y(_05560_),
    .A2(_05481_),
    .A1(_00546_));
 sg13g2_nand2b_1 _12770_ (.Y(_05561_),
    .B(_05560_),
    .A_N(_05418_));
 sg13g2_xnor2_1 _12771_ (.Y(_05562_),
    .A(_05418_),
    .B(_05560_));
 sg13g2_o21ai_1 _12772_ (.B1(_05542_),
    .Y(_05563_),
    .A1(_05473_),
    .A2(_05481_));
 sg13g2_nand2_1 _12773_ (.Y(_05564_),
    .A(_05562_),
    .B(_05563_));
 sg13g2_xor2_1 _12774_ (.B(_05563_),
    .A(_05562_),
    .X(_05565_));
 sg13g2_inv_1 _12775_ (.Y(_05566_),
    .A(_05565_));
 sg13g2_xnor2_1 _12776_ (.Y(_05567_),
    .A(net1925),
    .B(_05565_));
 sg13g2_and2_1 _12777_ (.A(_05558_),
    .B(_05567_),
    .X(_05568_));
 sg13g2_xor2_1 _12778_ (.B(_05567_),
    .A(_05558_),
    .X(_05569_));
 sg13g2_xnor2_1 _12779_ (.Y(_05570_),
    .A(\vgadonut.donut.ycA[17] ),
    .B(_05569_));
 sg13g2_nor2_1 _12780_ (.A(_05557_),
    .B(_05570_),
    .Y(_05571_));
 sg13g2_nand2_1 _12781_ (.Y(_05572_),
    .A(_05557_),
    .B(_05570_));
 sg13g2_nand2b_1 _12782_ (.Y(_05573_),
    .B(_05572_),
    .A_N(_05571_));
 sg13g2_a21o_1 _12783_ (.A2(net1613),
    .A1(\vgadonut.donut.donuthit.ryin[10] ),
    .B1(_05535_),
    .X(_05574_));
 sg13g2_nor2_1 _12784_ (.A(\vgadonut.donut.donuthit.ryin[11] ),
    .B(_05508_),
    .Y(_05575_));
 sg13g2_xnor2_1 _12785_ (.Y(_05576_),
    .A(_00550_),
    .B(net1613));
 sg13g2_xnor2_1 _12786_ (.Y(_05577_),
    .A(_05556_),
    .B(_05573_));
 sg13g2_xnor2_1 _12787_ (.Y(_05578_),
    .A(_05574_),
    .B(_05576_));
 sg13g2_a21oi_1 _12788_ (.A1(net1745),
    .A2(_05578_),
    .Y(_05579_),
    .B1(net1660));
 sg13g2_o21ai_1 _12789_ (.B1(_05579_),
    .Y(_05580_),
    .A1(net1755),
    .A2(_05577_));
 sg13g2_o21ai_1 _12790_ (.B1(_05580_),
    .Y(_00385_),
    .A1(_00550_),
    .A2(net1670));
 sg13g2_xnor2_1 _12791_ (.Y(_05581_),
    .A(\vgadonut.donut.donuthit.ryin[12] ),
    .B(net1614));
 sg13g2_a21oi_1 _12792_ (.A1(\vgadonut.donut.donuthit.ryin[11] ),
    .A2(net1613),
    .Y(_05582_),
    .B1(_05574_));
 sg13g2_nor3_1 _12793_ (.A(_05575_),
    .B(_05581_),
    .C(_05582_),
    .Y(_05583_));
 sg13g2_o21ai_1 _12794_ (.B1(_05581_),
    .Y(_05584_),
    .A1(_05575_),
    .A2(_05582_));
 sg13g2_nor2b_1 _12795_ (.A(_05583_),
    .B_N(_05584_),
    .Y(_05585_));
 sg13g2_a21oi_1 _12796_ (.A1(net1755),
    .A2(_05585_),
    .Y(_05586_),
    .B1(net1661));
 sg13g2_a21oi_1 _12797_ (.A1(_05556_),
    .A2(_05572_),
    .Y(_05587_),
    .B1(_05571_));
 sg13g2_o21ai_1 _12798_ (.B1(_05564_),
    .Y(_05588_),
    .A1(net1924),
    .A2(_05566_));
 sg13g2_nand2b_1 _12799_ (.Y(_05589_),
    .B(_05561_),
    .A_N(_05559_));
 sg13g2_nor2b_1 _12800_ (.A(_05428_),
    .B_N(_05589_),
    .Y(_05590_));
 sg13g2_xnor2_1 _12801_ (.Y(_05591_),
    .A(_05428_),
    .B(_05589_));
 sg13g2_xnor2_1 _12802_ (.Y(_05592_),
    .A(_00112_),
    .B(_05591_));
 sg13g2_nor2b_1 _12803_ (.A(_05592_),
    .B_N(_05588_),
    .Y(_05593_));
 sg13g2_xnor2_1 _12804_ (.Y(_05594_),
    .A(_05588_),
    .B(_05592_));
 sg13g2_xnor2_1 _12805_ (.Y(_05595_),
    .A(\vgadonut.donut.ycA[18] ),
    .B(_05594_));
 sg13g2_inv_1 _12806_ (.Y(_05596_),
    .A(_05595_));
 sg13g2_a21o_1 _12807_ (.A2(_05569_),
    .A1(\vgadonut.donut.ycA[17] ),
    .B1(_05568_),
    .X(_05597_));
 sg13g2_xor2_1 _12808_ (.B(_05597_),
    .A(_05595_),
    .X(_05598_));
 sg13g2_nor2_1 _12809_ (.A(_05587_),
    .B(_05598_),
    .Y(_05599_));
 sg13g2_a21oi_1 _12810_ (.A1(_05587_),
    .A2(_05598_),
    .Y(_05600_),
    .B1(net1745));
 sg13g2_nand2b_1 _12811_ (.Y(_05601_),
    .B(_05600_),
    .A_N(_05599_));
 sg13g2_a22oi_1 _12812_ (.Y(_00386_),
    .B1(_05586_),
    .B2(_05601_),
    .A2(net1661),
    .A1(_00551_));
 sg13g2_a21o_1 _12813_ (.A2(_05508_),
    .A1(\vgadonut.donut.donuthit.ryin[12] ),
    .B1(_05583_),
    .X(_05602_));
 sg13g2_xnor2_1 _12814_ (.Y(_05603_),
    .A(_00552_),
    .B(net1613));
 sg13g2_xor2_1 _12815_ (.B(_05603_),
    .A(_05602_),
    .X(_05604_));
 sg13g2_a21oi_1 _12816_ (.A1(net1755),
    .A2(_05604_),
    .Y(_05605_),
    .B1(net1660));
 sg13g2_a21oi_1 _12817_ (.A1(_05596_),
    .A2(_05597_),
    .Y(_05606_),
    .B1(_05599_));
 sg13g2_a21oi_1 _12818_ (.A1(_00112_),
    .A2(_05591_),
    .Y(_05607_),
    .B1(_05590_));
 sg13g2_nor2_1 _12819_ (.A(_05473_),
    .B(net1614),
    .Y(_05608_));
 sg13g2_a21oi_1 _12820_ (.A1(_00546_),
    .A2(_05473_),
    .Y(_05609_),
    .B1(_05608_));
 sg13g2_nand2b_1 _12821_ (.Y(_05610_),
    .B(_05609_),
    .A_N(net1921));
 sg13g2_xnor2_1 _12822_ (.Y(_05611_),
    .A(net1921),
    .B(_05609_));
 sg13g2_nor2b_1 _12823_ (.A(_05607_),
    .B_N(_05611_),
    .Y(_05612_));
 sg13g2_xnor2_1 _12824_ (.Y(_05613_),
    .A(_05607_),
    .B(_05611_));
 sg13g2_xnor2_1 _12825_ (.Y(_05614_),
    .A(\vgadonut.donut.ycA[19] ),
    .B(_05613_));
 sg13g2_a21oi_1 _12826_ (.A1(\vgadonut.donut.ycA[18] ),
    .A2(_05594_),
    .Y(_05615_),
    .B1(_05593_));
 sg13g2_nor2_1 _12827_ (.A(_05614_),
    .B(_05615_),
    .Y(_05616_));
 sg13g2_xnor2_1 _12828_ (.Y(_05617_),
    .A(_05614_),
    .B(_05615_));
 sg13g2_nor2_1 _12829_ (.A(_05606_),
    .B(_05617_),
    .Y(_05618_));
 sg13g2_a21oi_1 _12830_ (.A1(_05606_),
    .A2(_05617_),
    .Y(_05619_),
    .B1(net1745));
 sg13g2_nand2b_1 _12831_ (.Y(_05620_),
    .B(_05619_),
    .A_N(_05618_));
 sg13g2_a22oi_1 _12832_ (.Y(_00387_),
    .B1(_05605_),
    .B2(_05620_),
    .A2(net1660),
    .A1(_00552_));
 sg13g2_xnor2_1 _12833_ (.Y(_05621_),
    .A(\vgadonut.donut.donuthit.ryin[14] ),
    .B(net1613));
 sg13g2_nand2_1 _12834_ (.Y(_05622_),
    .A(_05583_),
    .B(_05603_));
 sg13g2_o21ai_1 _12835_ (.B1(_00114_),
    .Y(_05623_),
    .A1(_00551_),
    .A2(\vgadonut.donut.donuthit.ryin[13] ));
 sg13g2_nand2_1 _12836_ (.Y(_05624_),
    .A(net1613),
    .B(_05623_));
 sg13g2_a21oi_1 _12837_ (.A1(_05622_),
    .A2(_05624_),
    .Y(_05625_),
    .B1(_05621_));
 sg13g2_nand3_1 _12838_ (.B(_05622_),
    .C(_05624_),
    .A(_05621_),
    .Y(_05626_));
 sg13g2_nand2_1 _12839_ (.Y(_05627_),
    .A(net1745),
    .B(_05626_));
 sg13g2_o21ai_1 _12840_ (.B1(net1670),
    .Y(_05628_),
    .A1(_05625_),
    .A2(_05627_));
 sg13g2_nor2_1 _12841_ (.A(_05616_),
    .B(_05618_),
    .Y(_05629_));
 sg13g2_xnor2_1 _12842_ (.Y(_05630_),
    .A(_00113_),
    .B(_05560_));
 sg13g2_o21ai_1 _12843_ (.B1(_05610_),
    .Y(_05631_),
    .A1(_05473_),
    .A2(net1614));
 sg13g2_nor2b_1 _12844_ (.A(_05630_),
    .B_N(_05631_),
    .Y(_05632_));
 sg13g2_xnor2_1 _12845_ (.Y(_05633_),
    .A(_05630_),
    .B(_05631_));
 sg13g2_xnor2_1 _12846_ (.Y(_05634_),
    .A(\vgadonut.donut.ycA[20] ),
    .B(_05633_));
 sg13g2_a21oi_1 _12847_ (.A1(\vgadonut.donut.ycA[19] ),
    .A2(_05613_),
    .Y(_05635_),
    .B1(_05612_));
 sg13g2_nor2_1 _12848_ (.A(_05634_),
    .B(_05635_),
    .Y(_05636_));
 sg13g2_xnor2_1 _12849_ (.Y(_05637_),
    .A(_05634_),
    .B(_05635_));
 sg13g2_or2_1 _12850_ (.X(_05638_),
    .B(_05637_),
    .A(_05629_));
 sg13g2_a21oi_1 _12851_ (.A1(_05629_),
    .A2(_05637_),
    .Y(_05639_),
    .B1(net1745));
 sg13g2_a21oi_1 _12852_ (.A1(_05638_),
    .A2(_05639_),
    .Y(_05640_),
    .B1(_05628_));
 sg13g2_a21oi_1 _12853_ (.A1(_00555_),
    .A2(net1668),
    .Y(_00388_),
    .B1(_05640_));
 sg13g2_a21oi_1 _12854_ (.A1(\vgadonut.donut.donuthit.ryin[14] ),
    .A2(net1613),
    .Y(_05641_),
    .B1(_05625_));
 sg13g2_xnor2_1 _12855_ (.Y(_05642_),
    .A(_00559_),
    .B(net1613));
 sg13g2_xnor2_1 _12856_ (.Y(_05643_),
    .A(_05641_),
    .B(_05642_));
 sg13g2_a21oi_1 _12857_ (.A1(net1755),
    .A2(_05643_),
    .Y(_05644_),
    .B1(net1661));
 sg13g2_nor2b_1 _12858_ (.A(_05636_),
    .B_N(_05638_),
    .Y(_05645_));
 sg13g2_a21oi_1 _12859_ (.A1(\vgadonut.donut.ycA[20] ),
    .A2(_05633_),
    .Y(_05646_),
    .B1(_05632_));
 sg13g2_a21oi_1 _12860_ (.A1(_00113_),
    .A2(_05560_),
    .Y(_05647_),
    .B1(_05559_));
 sg13g2_xor2_1 _12861_ (.B(\vgadonut.donut.ycA[21] ),
    .A(net1917),
    .X(_05648_));
 sg13g2_xnor2_1 _12862_ (.Y(_05649_),
    .A(_05647_),
    .B(_05648_));
 sg13g2_xnor2_1 _12863_ (.Y(_05650_),
    .A(_05646_),
    .B(_05649_));
 sg13g2_o21ai_1 _12864_ (.B1(net1749),
    .Y(_05651_),
    .A1(_05645_),
    .A2(_05650_));
 sg13g2_a21o_1 _12865_ (.A2(_05650_),
    .A1(_05645_),
    .B1(_05651_),
    .X(_05652_));
 sg13g2_a22oi_1 _12866_ (.Y(_00389_),
    .B1(_05644_),
    .B2(_05652_),
    .A2(net1660),
    .A1(_00559_));
 sg13g2_xnor2_1 _12867_ (.Y(_05653_),
    .A(\vgadonut.donut.rx6[2] ),
    .B(net1864));
 sg13g2_and3_1 _12868_ (.X(_05654_),
    .A(_03939_),
    .B(_03941_),
    .C(_05653_));
 sg13g2_a21oi_1 _12869_ (.A1(_03939_),
    .A2(_03941_),
    .Y(_05655_),
    .B1(_05653_));
 sg13g2_nor3_1 _12870_ (.A(net1763),
    .B(_05654_),
    .C(_05655_),
    .Y(_05656_));
 sg13g2_a21oi_1 _12871_ (.A1(net1867),
    .A2(net1763),
    .Y(_05657_),
    .B1(_05656_));
 sg13g2_nand2_1 _12872_ (.Y(_05658_),
    .A(net2012),
    .B(net1658));
 sg13g2_o21ai_1 _12873_ (.B1(_05658_),
    .Y(_00390_),
    .A1(net1658),
    .A2(_05657_));
 sg13g2_a21oi_1 _12874_ (.A1(\vgadonut.donut.rx6[2] ),
    .A2(net1864),
    .Y(_05659_),
    .B1(_05655_));
 sg13g2_xnor2_1 _12875_ (.Y(_05660_),
    .A(\vgadonut.donut.rx6[3] ),
    .B(net1863));
 sg13g2_nand2_1 _12876_ (.Y(_05661_),
    .A(_05659_),
    .B(_05660_));
 sg13g2_nor2_1 _12877_ (.A(_05659_),
    .B(_05660_),
    .Y(_05662_));
 sg13g2_nor2_1 _12878_ (.A(net1763),
    .B(_05662_),
    .Y(_05663_));
 sg13g2_a221oi_1 _12879_ (.B2(_05663_),
    .C1(net1658),
    .B1(_05661_),
    .A1(net1866),
    .Y(_05664_),
    .A2(net1763));
 sg13g2_a21oi_1 _12880_ (.A1(_00560_),
    .A2(net1658),
    .Y(_00391_),
    .B1(_05664_));
 sg13g2_a21oi_1 _12881_ (.A1(\vgadonut.donut.rx6[3] ),
    .A2(net1863),
    .Y(_05665_),
    .B1(_05662_));
 sg13g2_nand2_1 _12882_ (.Y(_05666_),
    .A(\vgadonut.donut.rx6[4] ),
    .B(\vgadonut.donut.cB[4] ));
 sg13g2_xnor2_1 _12883_ (.Y(_05667_),
    .A(\vgadonut.donut.rx6[4] ),
    .B(\vgadonut.donut.cB[4] ));
 sg13g2_xnor2_1 _12884_ (.Y(_05668_),
    .A(_05665_),
    .B(_05667_));
 sg13g2_nor2b_1 _12885_ (.A(net1865),
    .B_N(\vgadonut.donut.cB[0] ),
    .Y(_05669_));
 sg13g2_xnor2_1 _12886_ (.Y(_05670_),
    .A(net1864),
    .B(\vgadonut.donut.cB[0] ));
 sg13g2_a221oi_1 _12887_ (.B2(net1763),
    .C1(net1659),
    .B1(_05670_),
    .A1(net1755),
    .Y(_05671_),
    .A2(_05668_));
 sg13g2_a21o_1 _12888_ (.A2(net1659),
    .A1(net2060),
    .B1(_05671_),
    .X(_00392_));
 sg13g2_o21ai_1 _12889_ (.B1(_05666_),
    .Y(_05672_),
    .A1(_05665_),
    .A2(_05667_));
 sg13g2_xnor2_1 _12890_ (.Y(_05673_),
    .A(\vgadonut.donut.rx6[5] ),
    .B(\vgadonut.donut.cB[5] ));
 sg13g2_xnor2_1 _12891_ (.Y(_05674_),
    .A(_05672_),
    .B(_05673_));
 sg13g2_nand2b_1 _12892_ (.Y(_05675_),
    .B(\vgadonut.donut.cB[3] ),
    .A_N(\vgadonut.donut.cB[1] ));
 sg13g2_xnor2_1 _12893_ (.Y(_05676_),
    .A(\vgadonut.donut.cB[1] ),
    .B(\vgadonut.donut.cB[3] ));
 sg13g2_nand2b_1 _12894_ (.Y(_05677_),
    .B(_05676_),
    .A_N(_05669_));
 sg13g2_xnor2_1 _12895_ (.Y(_05678_),
    .A(_05669_),
    .B(_05676_));
 sg13g2_a221oi_1 _12896_ (.B2(_03931_),
    .C1(net1659),
    .B1(_05678_),
    .A1(net1755),
    .Y(_05679_),
    .A2(_05674_));
 sg13g2_a21oi_1 _12897_ (.A1(_00562_),
    .A2(net1659),
    .Y(_00393_),
    .B1(_05679_));
 sg13g2_nand2_1 _12898_ (.Y(_05680_),
    .A(net2043),
    .B(\vgadonut.donut.cB[6] ));
 sg13g2_xnor2_1 _12899_ (.Y(_05681_),
    .A(\vgadonut.donut.donuthit.rxin[0] ),
    .B(\vgadonut.donut.cB[6] ));
 sg13g2_a21oi_1 _12900_ (.A1(\vgadonut.donut.rx6[5] ),
    .A2(\vgadonut.donut.cB[5] ),
    .Y(_05682_),
    .B1(_05672_));
 sg13g2_a21oi_2 _12901_ (.B1(_05682_),
    .Y(_05683_),
    .A2(_00563_),
    .A1(_00562_));
 sg13g2_nand2b_1 _12902_ (.Y(_05684_),
    .B(_05683_),
    .A_N(_05681_));
 sg13g2_xnor2_1 _12903_ (.Y(_05685_),
    .A(_05681_),
    .B(_05683_));
 sg13g2_o21ai_1 _12904_ (.B1(_05677_),
    .Y(_05686_),
    .A1(net1865),
    .A2(_05675_));
 sg13g2_nand2_1 _12905_ (.Y(_05687_),
    .A(net1865),
    .B(_05675_));
 sg13g2_nor2_1 _12906_ (.A(net1867),
    .B(\vgadonut.donut.sB[0] ),
    .Y(_05688_));
 sg13g2_xor2_1 _12907_ (.B(\vgadonut.donut.sB[0] ),
    .A(net1867),
    .X(_05689_));
 sg13g2_xnor2_1 _12908_ (.Y(_05690_),
    .A(_00115_),
    .B(_05689_));
 sg13g2_xor2_1 _12909_ (.B(_05690_),
    .A(_05687_),
    .X(_05691_));
 sg13g2_a21oi_1 _12910_ (.A1(_05686_),
    .A2(_05691_),
    .Y(_05692_),
    .B1(net1753));
 sg13g2_o21ai_1 _12911_ (.B1(_05692_),
    .Y(_05693_),
    .A1(_05686_),
    .A2(_05691_));
 sg13g2_a21oi_1 _12912_ (.A1(net1753),
    .A2(_05685_),
    .Y(_05694_),
    .B1(net1663));
 sg13g2_a22oi_1 _12913_ (.Y(_00394_),
    .B1(_05693_),
    .B2(_05694_),
    .A2(net1663),
    .A1(_00564_));
 sg13g2_nand2_1 _12914_ (.Y(_05695_),
    .A(net2084),
    .B(\vgadonut.donut.cB[7] ));
 sg13g2_xnor2_1 _12915_ (.Y(_05696_),
    .A(\vgadonut.donut.donuthit.rxin[1] ),
    .B(\vgadonut.donut.cB[7] ));
 sg13g2_nand3_1 _12916_ (.B(_05684_),
    .C(_05696_),
    .A(_05680_),
    .Y(_05697_));
 sg13g2_a21o_1 _12917_ (.A2(_05684_),
    .A1(_05680_),
    .B1(_05696_),
    .X(_05698_));
 sg13g2_nand3_1 _12918_ (.B(_05697_),
    .C(_05698_),
    .A(net1746),
    .Y(_05699_));
 sg13g2_o21ai_1 _12919_ (.B1(_05690_),
    .Y(_05700_),
    .A1(net1865),
    .A2(_00561_));
 sg13g2_nor2b_1 _12920_ (.A(_05700_),
    .B_N(_05687_),
    .Y(_05701_));
 sg13g2_a21o_1 _12921_ (.A2(_05691_),
    .A1(_05686_),
    .B1(_05701_),
    .X(_05702_));
 sg13g2_nand2_1 _12922_ (.Y(_05703_),
    .A(net1863),
    .B(_05690_));
 sg13g2_a21oi_1 _12923_ (.A1(_00115_),
    .A2(_05689_),
    .Y(_05704_),
    .B1(_05688_));
 sg13g2_nor2_1 _12924_ (.A(net1866),
    .B(\vgadonut.donut.sB[1] ),
    .Y(_05705_));
 sg13g2_xor2_1 _12925_ (.B(\vgadonut.donut.sB[1] ),
    .A(net1866),
    .X(_05706_));
 sg13g2_xnor2_1 _12926_ (.Y(_05707_),
    .A(_00116_),
    .B(_05706_));
 sg13g2_or2_1 _12927_ (.X(_05708_),
    .B(_05707_),
    .A(_05704_));
 sg13g2_xor2_1 _12928_ (.B(_05707_),
    .A(_05704_),
    .X(_05709_));
 sg13g2_nand2_1 _12929_ (.Y(_05710_),
    .A(_00115_),
    .B(_05709_));
 sg13g2_xnor2_1 _12930_ (.Y(_05711_),
    .A(_00115_),
    .B(_05709_));
 sg13g2_nand2b_1 _12931_ (.Y(_05712_),
    .B(_05703_),
    .A_N(_05711_));
 sg13g2_xor2_1 _12932_ (.B(_05711_),
    .A(_05703_),
    .X(_05713_));
 sg13g2_o21ai_1 _12933_ (.B1(_05700_),
    .Y(_05714_),
    .A1(_00561_),
    .A2(_05690_));
 sg13g2_nor2_1 _12934_ (.A(_05713_),
    .B(_05714_),
    .Y(_05715_));
 sg13g2_xor2_1 _12935_ (.B(_05714_),
    .A(_05713_),
    .X(_05716_));
 sg13g2_and2_1 _12936_ (.A(_05702_),
    .B(_05716_),
    .X(_05717_));
 sg13g2_o21ai_1 _12937_ (.B1(net1749),
    .Y(_05718_),
    .A1(_05702_),
    .A2(_05716_));
 sg13g2_nor2_1 _12938_ (.A(_05717_),
    .B(_05718_),
    .Y(_05719_));
 sg13g2_nor2_1 _12939_ (.A(net1663),
    .B(_05719_),
    .Y(_05720_));
 sg13g2_a22oi_1 _12940_ (.Y(_00395_),
    .B1(_05699_),
    .B2(_05720_),
    .A2(net1662),
    .A1(_00565_));
 sg13g2_xnor2_1 _12941_ (.Y(_05721_),
    .A(\vgadonut.donut.donuthit.rxin[2] ),
    .B(\vgadonut.donut.cB[8] ));
 sg13g2_a21o_1 _12942_ (.A2(_05698_),
    .A1(_05695_),
    .B1(_05721_),
    .X(_05722_));
 sg13g2_nand3_1 _12943_ (.B(_05698_),
    .C(_05721_),
    .A(_05695_),
    .Y(_05723_));
 sg13g2_nand3_1 _12944_ (.B(_05722_),
    .C(_05723_),
    .A(net1746),
    .Y(_05724_));
 sg13g2_nor2_1 _12945_ (.A(_05715_),
    .B(_05717_),
    .Y(_05725_));
 sg13g2_a21oi_1 _12946_ (.A1(_00116_),
    .A2(_05706_),
    .Y(_05726_),
    .B1(_05705_));
 sg13g2_nor2_1 _12947_ (.A(net1864),
    .B(\vgadonut.donut.donuthit.cordicxy.x2in[0] ),
    .Y(_05727_));
 sg13g2_xor2_1 _12948_ (.B(\vgadonut.donut.donuthit.cordicxy.x2in[0] ),
    .A(net1864),
    .X(_05728_));
 sg13g2_xnor2_1 _12949_ (.Y(_05729_),
    .A(_00117_),
    .B(_05728_));
 sg13g2_nor2_1 _12950_ (.A(_05726_),
    .B(_05729_),
    .Y(_05730_));
 sg13g2_xor2_1 _12951_ (.B(_05729_),
    .A(_05726_),
    .X(_05731_));
 sg13g2_xnor2_1 _12952_ (.Y(_05732_),
    .A(_00116_),
    .B(_05731_));
 sg13g2_and3_1 _12953_ (.X(_05733_),
    .A(_05708_),
    .B(_05710_),
    .C(_05732_));
 sg13g2_a21oi_2 _12954_ (.B1(_05732_),
    .Y(_05734_),
    .A2(_05710_),
    .A1(_05708_));
 sg13g2_or2_1 _12955_ (.X(_05735_),
    .B(_05734_),
    .A(_05733_));
 sg13g2_xnor2_1 _12956_ (.Y(_05736_),
    .A(_05712_),
    .B(_05735_));
 sg13g2_or2_1 _12957_ (.X(_05737_),
    .B(_05736_),
    .A(_05725_));
 sg13g2_a21oi_1 _12958_ (.A1(_05725_),
    .A2(_05736_),
    .Y(_05738_),
    .B1(net1746));
 sg13g2_a21oi_1 _12959_ (.A1(_05737_),
    .A2(_05738_),
    .Y(_05739_),
    .B1(net1663));
 sg13g2_a22oi_1 _12960_ (.Y(_00396_),
    .B1(_05724_),
    .B2(_05739_),
    .A2(net1662),
    .A1(_00567_));
 sg13g2_o21ai_1 _12961_ (.B1(_05722_),
    .Y(_05740_),
    .A1(_00567_),
    .A2(_00568_));
 sg13g2_nor2_1 _12962_ (.A(\vgadonut.donut.donuthit.rxin[3] ),
    .B(\vgadonut.donut.cB[9] ),
    .Y(_05741_));
 sg13g2_xnor2_1 _12963_ (.Y(_05742_),
    .A(\vgadonut.donut.donuthit.rxin[3] ),
    .B(\vgadonut.donut.cB[9] ));
 sg13g2_xnor2_1 _12964_ (.Y(_05743_),
    .A(_05740_),
    .B(_05742_));
 sg13g2_o21ai_1 _12965_ (.B1(_05737_),
    .Y(_05744_),
    .A1(_05712_),
    .A2(_05735_));
 sg13g2_a21oi_1 _12966_ (.A1(_00117_),
    .A2(_05728_),
    .Y(_05745_),
    .B1(_05727_));
 sg13g2_nor2_1 _12967_ (.A(net1863),
    .B(\vgadonut.donut.donuthit.cordicxy.x2in[1] ),
    .Y(_05746_));
 sg13g2_xor2_1 _12968_ (.B(\vgadonut.donut.donuthit.cordicxy.x2in[1] ),
    .A(net1863),
    .X(_05747_));
 sg13g2_xnor2_1 _12969_ (.Y(_05748_),
    .A(_00118_),
    .B(_05747_));
 sg13g2_nor2_1 _12970_ (.A(_05745_),
    .B(_05748_),
    .Y(_05749_));
 sg13g2_xor2_1 _12971_ (.B(_05748_),
    .A(_05745_),
    .X(_05750_));
 sg13g2_xnor2_1 _12972_ (.Y(_05751_),
    .A(_00117_),
    .B(_05750_));
 sg13g2_a21oi_1 _12973_ (.A1(_00116_),
    .A2(_05731_),
    .Y(_05752_),
    .B1(_05730_));
 sg13g2_nor2_1 _12974_ (.A(_05751_),
    .B(_05752_),
    .Y(_05753_));
 sg13g2_xnor2_1 _12975_ (.Y(_05754_),
    .A(_05751_),
    .B(_05752_));
 sg13g2_inv_1 _12976_ (.Y(_05755_),
    .A(_05754_));
 sg13g2_nand2_1 _12977_ (.Y(_05756_),
    .A(_05734_),
    .B(_05755_));
 sg13g2_xnor2_1 _12978_ (.Y(_05757_),
    .A(_05734_),
    .B(_05754_));
 sg13g2_or2_1 _12979_ (.X(_05758_),
    .B(_05757_),
    .A(_05744_));
 sg13g2_nand2_1 _12980_ (.Y(_05759_),
    .A(_05744_),
    .B(_05757_));
 sg13g2_nand3_1 _12981_ (.B(_05758_),
    .C(_05759_),
    .A(net1758),
    .Y(_05760_));
 sg13g2_a21oi_1 _12982_ (.A1(net1753),
    .A2(_05743_),
    .Y(_05761_),
    .B1(net1662));
 sg13g2_a22oi_1 _12983_ (.Y(_00397_),
    .B1(_05760_),
    .B2(_05761_),
    .A2(net1662),
    .A1(_00570_));
 sg13g2_xnor2_1 _12984_ (.Y(_05762_),
    .A(\vgadonut.donut.donuthit.rxin[4] ),
    .B(\vgadonut.donut.cB[10] ));
 sg13g2_a21oi_1 _12985_ (.A1(\vgadonut.donut.donuthit.rxin[3] ),
    .A2(\vgadonut.donut.cB[9] ),
    .Y(_05763_),
    .B1(_05740_));
 sg13g2_nor3_1 _12986_ (.A(_05741_),
    .B(_05762_),
    .C(_05763_),
    .Y(_05764_));
 sg13g2_o21ai_1 _12987_ (.B1(_05762_),
    .Y(_05765_),
    .A1(_05741_),
    .A2(_05763_));
 sg13g2_nor2b_1 _12988_ (.A(_05764_),
    .B_N(_05765_),
    .Y(_05766_));
 sg13g2_a21oi_1 _12989_ (.A1(_00118_),
    .A2(_05747_),
    .Y(_05767_),
    .B1(_05746_));
 sg13g2_nor2_1 _12990_ (.A(\vgadonut.donut.cB[4] ),
    .B(net1884),
    .Y(_05768_));
 sg13g2_xor2_1 _12991_ (.B(net1884),
    .A(\vgadonut.donut.cB[4] ),
    .X(_05769_));
 sg13g2_xnor2_1 _12992_ (.Y(_05770_),
    .A(_00119_),
    .B(_05769_));
 sg13g2_nor2_1 _12993_ (.A(_05767_),
    .B(_05770_),
    .Y(_05771_));
 sg13g2_xor2_1 _12994_ (.B(_05770_),
    .A(_05767_),
    .X(_05772_));
 sg13g2_xnor2_1 _12995_ (.Y(_05773_),
    .A(_00118_),
    .B(_05772_));
 sg13g2_a21oi_1 _12996_ (.A1(_00117_),
    .A2(_05750_),
    .Y(_05774_),
    .B1(_05749_));
 sg13g2_nor2_1 _12997_ (.A(_05773_),
    .B(_05774_),
    .Y(_05775_));
 sg13g2_xor2_1 _12998_ (.B(_05774_),
    .A(_05773_),
    .X(_05776_));
 sg13g2_nand2_1 _12999_ (.Y(_05777_),
    .A(_05753_),
    .B(_05776_));
 sg13g2_xnor2_1 _13000_ (.Y(_05778_),
    .A(_05753_),
    .B(_05776_));
 sg13g2_nand3_1 _13001_ (.B(_05759_),
    .C(_05778_),
    .A(_05756_),
    .Y(_05779_));
 sg13g2_a21o_1 _13002_ (.A2(_05759_),
    .A1(_05756_),
    .B1(_05778_),
    .X(_05780_));
 sg13g2_nand3_1 _13003_ (.B(_05779_),
    .C(_05780_),
    .A(net1758),
    .Y(_05781_));
 sg13g2_a21oi_1 _13004_ (.A1(net1753),
    .A2(_05766_),
    .Y(_05782_),
    .B1(net1662));
 sg13g2_a22oi_1 _13005_ (.Y(_00398_),
    .B1(_05781_),
    .B2(_05782_),
    .A2(net1662),
    .A1(_00571_));
 sg13g2_a21o_1 _13006_ (.A2(\vgadonut.donut.cB[10] ),
    .A1(\vgadonut.donut.donuthit.rxin[4] ),
    .B1(_05764_),
    .X(_05783_));
 sg13g2_nor2_1 _13007_ (.A(\vgadonut.donut.donuthit.rxin[5] ),
    .B(\vgadonut.donut.cB[11] ),
    .Y(_05784_));
 sg13g2_xnor2_1 _13008_ (.Y(_05785_),
    .A(\vgadonut.donut.donuthit.rxin[5] ),
    .B(\vgadonut.donut.cB[11] ));
 sg13g2_xnor2_1 _13009_ (.Y(_05786_),
    .A(_05783_),
    .B(_05785_));
 sg13g2_a21oi_1 _13010_ (.A1(_00119_),
    .A2(_05769_),
    .Y(_05787_),
    .B1(_05768_));
 sg13g2_nor2_1 _13011_ (.A(\vgadonut.donut.cB[5] ),
    .B(\vgadonut.donut.donuthit.cordicxy.x2in[3] ),
    .Y(_05788_));
 sg13g2_xor2_1 _13012_ (.B(\vgadonut.donut.donuthit.cordicxy.x2in[3] ),
    .A(\vgadonut.donut.cB[5] ),
    .X(_05789_));
 sg13g2_xnor2_1 _13013_ (.Y(_05790_),
    .A(_00120_),
    .B(_05789_));
 sg13g2_nor2_1 _13014_ (.A(_05787_),
    .B(_05790_),
    .Y(_05791_));
 sg13g2_xor2_1 _13015_ (.B(_05790_),
    .A(_05787_),
    .X(_05792_));
 sg13g2_xnor2_1 _13016_ (.Y(_05793_),
    .A(_00119_),
    .B(_05792_));
 sg13g2_a21oi_1 _13017_ (.A1(_00118_),
    .A2(_05772_),
    .Y(_05794_),
    .B1(_05771_));
 sg13g2_nor2_1 _13018_ (.A(_05793_),
    .B(_05794_),
    .Y(_05795_));
 sg13g2_xor2_1 _13019_ (.B(_05794_),
    .A(_05793_),
    .X(_05796_));
 sg13g2_nand2_1 _13020_ (.Y(_05797_),
    .A(_05775_),
    .B(_05796_));
 sg13g2_xnor2_1 _13021_ (.Y(_05798_),
    .A(_05775_),
    .B(_05796_));
 sg13g2_nand3_1 _13022_ (.B(_05780_),
    .C(_05798_),
    .A(_05777_),
    .Y(_05799_));
 sg13g2_a21o_1 _13023_ (.A2(_05780_),
    .A1(_05777_),
    .B1(_05798_),
    .X(_05800_));
 sg13g2_nand3_1 _13024_ (.B(_05799_),
    .C(_05800_),
    .A(net1758),
    .Y(_05801_));
 sg13g2_a21oi_1 _13025_ (.A1(net1753),
    .A2(_05786_),
    .Y(_05802_),
    .B1(net1662));
 sg13g2_a22oi_1 _13026_ (.Y(_00399_),
    .B1(_05801_),
    .B2(_05802_),
    .A2(net1662),
    .A1(_00574_));
 sg13g2_xnor2_1 _13027_ (.Y(_05803_),
    .A(\vgadonut.donut.donuthit.rxin[6] ),
    .B(\vgadonut.donut.cB[12] ));
 sg13g2_a21oi_1 _13028_ (.A1(\vgadonut.donut.donuthit.rxin[5] ),
    .A2(\vgadonut.donut.cB[11] ),
    .Y(_05804_),
    .B1(_05783_));
 sg13g2_or3_1 _13029_ (.A(_05784_),
    .B(_05803_),
    .C(_05804_),
    .X(_05805_));
 sg13g2_o21ai_1 _13030_ (.B1(_05803_),
    .Y(_05806_),
    .A1(_05784_),
    .A2(_05804_));
 sg13g2_and2_1 _13031_ (.A(_05805_),
    .B(_05806_),
    .X(_05807_));
 sg13g2_a21oi_1 _13032_ (.A1(_00120_),
    .A2(_05789_),
    .Y(_05808_),
    .B1(_05788_));
 sg13g2_nor2_1 _13033_ (.A(\vgadonut.donut.cB[6] ),
    .B(net1883),
    .Y(_05809_));
 sg13g2_xor2_1 _13034_ (.B(net1883),
    .A(\vgadonut.donut.cB[6] ),
    .X(_05810_));
 sg13g2_xnor2_1 _13035_ (.Y(_05811_),
    .A(_00121_),
    .B(_05810_));
 sg13g2_nor2_1 _13036_ (.A(_05808_),
    .B(_05811_),
    .Y(_05812_));
 sg13g2_xor2_1 _13037_ (.B(_05811_),
    .A(_05808_),
    .X(_05813_));
 sg13g2_xnor2_1 _13038_ (.Y(_05814_),
    .A(_00120_),
    .B(_05813_));
 sg13g2_a21oi_1 _13039_ (.A1(_00119_),
    .A2(_05792_),
    .Y(_05815_),
    .B1(_05791_));
 sg13g2_nor2_1 _13040_ (.A(_05814_),
    .B(_05815_),
    .Y(_05816_));
 sg13g2_xor2_1 _13041_ (.B(_05815_),
    .A(_05814_),
    .X(_05817_));
 sg13g2_nand2_1 _13042_ (.Y(_05818_),
    .A(_05795_),
    .B(_05817_));
 sg13g2_xnor2_1 _13043_ (.Y(_05819_),
    .A(_05795_),
    .B(_05817_));
 sg13g2_nand3_1 _13044_ (.B(_05800_),
    .C(_05819_),
    .A(_05797_),
    .Y(_05820_));
 sg13g2_a21o_1 _13045_ (.A2(_05800_),
    .A1(_05797_),
    .B1(_05819_),
    .X(_05821_));
 sg13g2_nand3_1 _13046_ (.B(_05820_),
    .C(_05821_),
    .A(net1758),
    .Y(_05822_));
 sg13g2_a21oi_1 _13047_ (.A1(net1753),
    .A2(_05807_),
    .Y(_05823_),
    .B1(net1667));
 sg13g2_a22oi_1 _13048_ (.Y(_00400_),
    .B1(_05822_),
    .B2(_05823_),
    .A2(net1663),
    .A1(_00575_));
 sg13g2_o21ai_1 _13049_ (.B1(_05805_),
    .Y(_05824_),
    .A1(_00575_),
    .A2(_00576_));
 sg13g2_nor2_1 _13050_ (.A(\vgadonut.donut.donuthit.rxin[7] ),
    .B(\vgadonut.donut.cB[13] ),
    .Y(_05825_));
 sg13g2_xnor2_1 _13051_ (.Y(_05826_),
    .A(\vgadonut.donut.donuthit.rxin[7] ),
    .B(\vgadonut.donut.cB[13] ));
 sg13g2_xnor2_1 _13052_ (.Y(_05827_),
    .A(_05824_),
    .B(_05826_));
 sg13g2_a21oi_1 _13053_ (.A1(_00121_),
    .A2(_05810_),
    .Y(_05828_),
    .B1(_05809_));
 sg13g2_nor2_1 _13054_ (.A(\vgadonut.donut.cB[7] ),
    .B(\vgadonut.donut.donuthit.cordicxy.x2in[5] ),
    .Y(_05829_));
 sg13g2_xor2_1 _13055_ (.B(\vgadonut.donut.donuthit.cordicxy.x2in[5] ),
    .A(\vgadonut.donut.cB[7] ),
    .X(_05830_));
 sg13g2_xnor2_1 _13056_ (.Y(_05831_),
    .A(_00122_),
    .B(_05830_));
 sg13g2_nor2_1 _13057_ (.A(_05828_),
    .B(_05831_),
    .Y(_05832_));
 sg13g2_xor2_1 _13058_ (.B(_05831_),
    .A(_05828_),
    .X(_05833_));
 sg13g2_xnor2_1 _13059_ (.Y(_05834_),
    .A(_00121_),
    .B(_05833_));
 sg13g2_a21oi_1 _13060_ (.A1(_00120_),
    .A2(_05813_),
    .Y(_05835_),
    .B1(_05812_));
 sg13g2_nor2_1 _13061_ (.A(_05834_),
    .B(_05835_),
    .Y(_05836_));
 sg13g2_xor2_1 _13062_ (.B(_05835_),
    .A(_05834_),
    .X(_05837_));
 sg13g2_nand2_1 _13063_ (.Y(_05838_),
    .A(_05816_),
    .B(_05837_));
 sg13g2_xnor2_1 _13064_ (.Y(_05839_),
    .A(_05816_),
    .B(_05837_));
 sg13g2_nand3_1 _13065_ (.B(_05821_),
    .C(_05839_),
    .A(_05818_),
    .Y(_05840_));
 sg13g2_a21o_1 _13066_ (.A2(_05821_),
    .A1(_05818_),
    .B1(_05839_),
    .X(_05841_));
 sg13g2_nand3_1 _13067_ (.B(_05840_),
    .C(_05841_),
    .A(net1759),
    .Y(_05842_));
 sg13g2_a21oi_1 _13068_ (.A1(net1753),
    .A2(_05827_),
    .Y(_05843_),
    .B1(net1663));
 sg13g2_a22oi_1 _13069_ (.Y(_00401_),
    .B1(_05842_),
    .B2(_05843_),
    .A2(net1663),
    .A1(_00578_));
 sg13g2_xnor2_1 _13070_ (.Y(_05844_),
    .A(\vgadonut.donut.donuthit.rxin[8] ),
    .B(net1862));
 sg13g2_a21oi_1 _13071_ (.A1(\vgadonut.donut.donuthit.rxin[7] ),
    .A2(\vgadonut.donut.cB[13] ),
    .Y(_05845_),
    .B1(_05824_));
 sg13g2_nor3_1 _13072_ (.A(_05825_),
    .B(_05844_),
    .C(_05845_),
    .Y(_05846_));
 sg13g2_o21ai_1 _13073_ (.B1(_05844_),
    .Y(_05847_),
    .A1(_05825_),
    .A2(_05845_));
 sg13g2_nor2b_1 _13074_ (.A(_05846_),
    .B_N(_05847_),
    .Y(_05848_));
 sg13g2_a21oi_1 _13075_ (.A1(_00122_),
    .A2(_05830_),
    .Y(_05849_),
    .B1(_05829_));
 sg13g2_nor2_1 _13076_ (.A(\vgadonut.donut.cB[8] ),
    .B(\vgadonut.donut.donuthit.cordicxy.x2in[6] ),
    .Y(_05850_));
 sg13g2_xor2_1 _13077_ (.B(\vgadonut.donut.donuthit.cordicxy.x2in[6] ),
    .A(\vgadonut.donut.cB[8] ),
    .X(_05851_));
 sg13g2_xnor2_1 _13078_ (.Y(_05852_),
    .A(_00123_),
    .B(_05851_));
 sg13g2_nor2_1 _13079_ (.A(_05849_),
    .B(_05852_),
    .Y(_05853_));
 sg13g2_xor2_1 _13080_ (.B(_05852_),
    .A(_05849_),
    .X(_05854_));
 sg13g2_xnor2_1 _13081_ (.Y(_05855_),
    .A(_00122_),
    .B(_05854_));
 sg13g2_a21oi_1 _13082_ (.A1(_00121_),
    .A2(_05833_),
    .Y(_05856_),
    .B1(_05832_));
 sg13g2_nor2_1 _13083_ (.A(_05855_),
    .B(_05856_),
    .Y(_05857_));
 sg13g2_xor2_1 _13084_ (.B(_05856_),
    .A(_05855_),
    .X(_05858_));
 sg13g2_nand2_1 _13085_ (.Y(_05859_),
    .A(_05836_),
    .B(_05858_));
 sg13g2_xnor2_1 _13086_ (.Y(_05860_),
    .A(_05836_),
    .B(_05858_));
 sg13g2_nand3_1 _13087_ (.B(_05841_),
    .C(_05860_),
    .A(_05838_),
    .Y(_05861_));
 sg13g2_a21o_1 _13088_ (.A2(_05841_),
    .A1(_05838_),
    .B1(_05860_),
    .X(_05862_));
 sg13g2_nand3_1 _13089_ (.B(_05861_),
    .C(_05862_),
    .A(net1758),
    .Y(_05863_));
 sg13g2_a21oi_1 _13090_ (.A1(net1754),
    .A2(_05848_),
    .Y(_05864_),
    .B1(net1666));
 sg13g2_a22oi_1 _13091_ (.Y(_00402_),
    .B1(_05863_),
    .B2(_05864_),
    .A2(net1666),
    .A1(_00580_));
 sg13g2_a21o_1 _13092_ (.A2(net1862),
    .A1(\vgadonut.donut.donuthit.rxin[8] ),
    .B1(_05846_),
    .X(_05865_));
 sg13g2_nor2_1 _13093_ (.A(\vgadonut.donut.donuthit.rxin[9] ),
    .B(net1860),
    .Y(_05866_));
 sg13g2_xnor2_1 _13094_ (.Y(_05867_),
    .A(\vgadonut.donut.donuthit.rxin[9] ),
    .B(net1861));
 sg13g2_xnor2_1 _13095_ (.Y(_05868_),
    .A(_05865_),
    .B(_05867_));
 sg13g2_a21oi_1 _13096_ (.A1(_00123_),
    .A2(_05851_),
    .Y(_05869_),
    .B1(_05850_));
 sg13g2_nor2_1 _13097_ (.A(\vgadonut.donut.cB[9] ),
    .B(net1880),
    .Y(_05870_));
 sg13g2_xor2_1 _13098_ (.B(net1880),
    .A(\vgadonut.donut.cB[9] ),
    .X(_05871_));
 sg13g2_xnor2_1 _13099_ (.Y(_05872_),
    .A(_00124_),
    .B(_05871_));
 sg13g2_or2_1 _13100_ (.X(_05873_),
    .B(_05872_),
    .A(_05869_));
 sg13g2_xor2_1 _13101_ (.B(_05872_),
    .A(_05869_),
    .X(_05874_));
 sg13g2_nand2_1 _13102_ (.Y(_05875_),
    .A(_00123_),
    .B(_05874_));
 sg13g2_xnor2_1 _13103_ (.Y(_05876_),
    .A(_00123_),
    .B(_05874_));
 sg13g2_a21oi_1 _13104_ (.A1(_00122_),
    .A2(_05854_),
    .Y(_05877_),
    .B1(_05853_));
 sg13g2_nor2_1 _13105_ (.A(_05876_),
    .B(_05877_),
    .Y(_05878_));
 sg13g2_xor2_1 _13106_ (.B(_05877_),
    .A(_05876_),
    .X(_05879_));
 sg13g2_nand2_1 _13107_ (.Y(_05880_),
    .A(_05857_),
    .B(_05879_));
 sg13g2_xnor2_1 _13108_ (.Y(_05881_),
    .A(_05857_),
    .B(_05879_));
 sg13g2_nand3_1 _13109_ (.B(_05862_),
    .C(_05881_),
    .A(_05859_),
    .Y(_05882_));
 sg13g2_a21o_1 _13110_ (.A2(_05862_),
    .A1(_05859_),
    .B1(_05881_),
    .X(_05883_));
 sg13g2_nand3_1 _13111_ (.B(_05882_),
    .C(_05883_),
    .A(net1758),
    .Y(_05884_));
 sg13g2_a21oi_1 _13112_ (.A1(net1754),
    .A2(_05868_),
    .Y(_05885_),
    .B1(net1666));
 sg13g2_a22oi_1 _13113_ (.Y(_00403_),
    .B1(_05884_),
    .B2(_05885_),
    .A2(net1666),
    .A1(_00581_));
 sg13g2_xnor2_1 _13114_ (.Y(_05886_),
    .A(net1860),
    .B(\vgadonut.donut.donuthit.rxin[10] ));
 sg13g2_a21oi_1 _13115_ (.A1(\vgadonut.donut.donuthit.rxin[9] ),
    .A2(net1861),
    .Y(_05887_),
    .B1(_05865_));
 sg13g2_o21ai_1 _13116_ (.B1(_05886_),
    .Y(_05888_),
    .A1(_05866_),
    .A2(_05887_));
 sg13g2_or3_1 _13117_ (.A(_05866_),
    .B(_05886_),
    .C(_05887_),
    .X(_05889_));
 sg13g2_and2_1 _13118_ (.A(_05888_),
    .B(_05889_),
    .X(_05890_));
 sg13g2_a21oi_1 _13119_ (.A1(_00124_),
    .A2(_05871_),
    .Y(_05891_),
    .B1(_05870_));
 sg13g2_xor2_1 _13120_ (.B(net1879),
    .A(\vgadonut.donut.cB[10] ),
    .X(_05892_));
 sg13g2_nand2b_1 _13121_ (.Y(_05893_),
    .B(_05892_),
    .A_N(\vgadonut.donut.cB[14] ));
 sg13g2_xnor2_1 _13122_ (.Y(_05894_),
    .A(\vgadonut.donut.cB[14] ),
    .B(_05892_));
 sg13g2_nor2b_1 _13123_ (.A(_05891_),
    .B_N(_05894_),
    .Y(_05895_));
 sg13g2_xnor2_1 _13124_ (.Y(_05896_),
    .A(_05891_),
    .B(_05894_));
 sg13g2_xnor2_1 _13125_ (.Y(_05897_),
    .A(_00124_),
    .B(_05896_));
 sg13g2_a21oi_2 _13126_ (.B1(_05897_),
    .Y(_05898_),
    .A2(_05875_),
    .A1(_05873_));
 sg13g2_nand3_1 _13127_ (.B(_05875_),
    .C(_05897_),
    .A(_05873_),
    .Y(_05899_));
 sg13g2_nor2b_1 _13128_ (.A(_05898_),
    .B_N(_05899_),
    .Y(_05900_));
 sg13g2_nand2_1 _13129_ (.Y(_05901_),
    .A(_05878_),
    .B(_05900_));
 sg13g2_xnor2_1 _13130_ (.Y(_05902_),
    .A(_05878_),
    .B(_05900_));
 sg13g2_nand3_1 _13131_ (.B(_05883_),
    .C(_05902_),
    .A(_05880_),
    .Y(_05903_));
 sg13g2_a21o_1 _13132_ (.A2(_05883_),
    .A1(_05880_),
    .B1(_05902_),
    .X(_05904_));
 sg13g2_nand3_1 _13133_ (.B(_05903_),
    .C(_05904_),
    .A(net1758),
    .Y(_05905_));
 sg13g2_a21oi_1 _13134_ (.A1(net1754),
    .A2(_05890_),
    .Y(_05906_),
    .B1(net1664));
 sg13g2_a22oi_1 _13135_ (.Y(_00404_),
    .B1(_05905_),
    .B2(_05906_),
    .A2(net1664),
    .A1(_00584_));
 sg13g2_xnor2_1 _13136_ (.Y(_05907_),
    .A(net1860),
    .B(\vgadonut.donut.donuthit.rxin[11] ));
 sg13g2_o21ai_1 _13137_ (.B1(_05889_),
    .Y(_05908_),
    .A1(_00582_),
    .A2(_00584_));
 sg13g2_xnor2_1 _13138_ (.Y(_05909_),
    .A(_05907_),
    .B(_05908_));
 sg13g2_nand2_1 _13139_ (.Y(_05910_),
    .A(_05901_),
    .B(_05904_));
 sg13g2_o21ai_1 _13140_ (.B1(_05893_),
    .Y(_05911_),
    .A1(\vgadonut.donut.cB[10] ),
    .A2(net1879));
 sg13g2_nor2_1 _13141_ (.A(\vgadonut.donut.cB[11] ),
    .B(net1877),
    .Y(_05912_));
 sg13g2_nand2_1 _13142_ (.Y(_05913_),
    .A(\vgadonut.donut.cB[11] ),
    .B(net1877));
 sg13g2_nor2_1 _13143_ (.A(net1858),
    .B(_05912_),
    .Y(_05914_));
 sg13g2_a21oi_1 _13144_ (.A1(net1858),
    .A2(_05913_),
    .Y(_05915_),
    .B1(_05912_));
 sg13g2_or2_1 _13145_ (.X(_05916_),
    .B(_05913_),
    .A(net1858));
 sg13g2_a22oi_1 _13146_ (.Y(_05917_),
    .B1(_05915_),
    .B2(_05916_),
    .A2(_05912_),
    .A1(net1858));
 sg13g2_nand2b_1 _13147_ (.Y(_05918_),
    .B(_05911_),
    .A_N(_05917_));
 sg13g2_xor2_1 _13148_ (.B(_05917_),
    .A(_05911_),
    .X(_05919_));
 sg13g2_or2_1 _13149_ (.X(_05920_),
    .B(_05919_),
    .A(net1862));
 sg13g2_xor2_1 _13150_ (.B(_05919_),
    .A(net1862),
    .X(_05921_));
 sg13g2_a21oi_1 _13151_ (.A1(_00124_),
    .A2(_05896_),
    .Y(_05922_),
    .B1(_05895_));
 sg13g2_nand2b_1 _13152_ (.Y(_05923_),
    .B(_05921_),
    .A_N(_05922_));
 sg13g2_xor2_1 _13153_ (.B(_05922_),
    .A(_05921_),
    .X(_05924_));
 sg13g2_inv_1 _13154_ (.Y(_05925_),
    .A(_05924_));
 sg13g2_nand2_1 _13155_ (.Y(_05926_),
    .A(_05904_),
    .B(_05924_));
 sg13g2_xnor2_1 _13156_ (.Y(_05927_),
    .A(_05910_),
    .B(_05924_));
 sg13g2_o21ai_1 _13157_ (.B1(net1758),
    .Y(_05928_),
    .A1(_05898_),
    .A2(_05927_));
 sg13g2_a21o_1 _13158_ (.A2(_05927_),
    .A1(_05898_),
    .B1(_05928_),
    .X(_05929_));
 sg13g2_a21oi_1 _13159_ (.A1(net1754),
    .A2(_05909_),
    .Y(_05930_),
    .B1(net1664));
 sg13g2_a22oi_1 _13160_ (.Y(_00405_),
    .B1(_05929_),
    .B2(_05930_),
    .A2(net1664),
    .A1(_00586_));
 sg13g2_xnor2_1 _13161_ (.Y(_05931_),
    .A(net1860),
    .B(\vgadonut.donut.donuthit.rxin[12] ));
 sg13g2_o21ai_1 _13162_ (.B1(net1860),
    .Y(_05932_),
    .A1(\vgadonut.donut.donuthit.rxin[10] ),
    .A2(\vgadonut.donut.donuthit.rxin[11] ));
 sg13g2_nor2_1 _13163_ (.A(_05889_),
    .B(_05907_),
    .Y(_05933_));
 sg13g2_nor2b_1 _13164_ (.A(_05933_),
    .B_N(_05932_),
    .Y(_05934_));
 sg13g2_or2_1 _13165_ (.X(_05935_),
    .B(_05934_),
    .A(_05931_));
 sg13g2_a21oi_1 _13166_ (.A1(_05931_),
    .A2(_05934_),
    .Y(_05936_),
    .B1(net1749));
 sg13g2_nor2_1 _13167_ (.A(\vgadonut.donut.cB[12] ),
    .B(net1875),
    .Y(_05937_));
 sg13g2_xor2_1 _13168_ (.B(net1875),
    .A(\vgadonut.donut.cB[12] ),
    .X(_05938_));
 sg13g2_xnor2_1 _13169_ (.Y(_05939_),
    .A(net1859),
    .B(_05938_));
 sg13g2_a21oi_1 _13170_ (.A1(net1858),
    .A2(_05913_),
    .Y(_05940_),
    .B1(_05914_));
 sg13g2_xnor2_1 _13171_ (.Y(_05941_),
    .A(_05939_),
    .B(_05940_));
 sg13g2_a21o_1 _13172_ (.A2(_05920_),
    .A1(_05918_),
    .B1(_05941_),
    .X(_05942_));
 sg13g2_nand3_1 _13173_ (.B(_05920_),
    .C(_05941_),
    .A(_05918_),
    .Y(_05943_));
 sg13g2_nand2_1 _13174_ (.Y(_05944_),
    .A(_05942_),
    .B(_05943_));
 sg13g2_nor2_1 _13175_ (.A(_05923_),
    .B(_05944_),
    .Y(_05945_));
 sg13g2_xnor2_1 _13176_ (.Y(_05946_),
    .A(_05923_),
    .B(_05944_));
 sg13g2_a22oi_1 _13177_ (.Y(_05947_),
    .B1(_05926_),
    .B2(_05898_),
    .A2(_05925_),
    .A1(_05910_));
 sg13g2_nor2_1 _13178_ (.A(_05946_),
    .B(_05947_),
    .Y(_05948_));
 sg13g2_nand2_1 _13179_ (.Y(_05949_),
    .A(_05946_),
    .B(_05947_));
 sg13g2_nor2_1 _13180_ (.A(net1753),
    .B(_05948_),
    .Y(_05950_));
 sg13g2_a221oi_1 _13181_ (.B2(_05950_),
    .C1(net1667),
    .B1(_05949_),
    .A1(_05935_),
    .Y(_05951_),
    .A2(_05936_));
 sg13g2_a21oi_1 _13182_ (.A1(_00588_),
    .A2(net1665),
    .Y(_00406_),
    .B1(_05951_));
 sg13g2_xor2_1 _13183_ (.B(\vgadonut.donut.donuthit.rxin[13] ),
    .A(net1859),
    .X(_05952_));
 sg13g2_o21ai_1 _13184_ (.B1(_05935_),
    .Y(_05953_),
    .A1(_00582_),
    .A2(_00588_));
 sg13g2_xor2_1 _13185_ (.B(_05953_),
    .A(_05952_),
    .X(_05954_));
 sg13g2_a21oi_1 _13186_ (.A1(net1754),
    .A2(_05954_),
    .Y(_05955_),
    .B1(net1665));
 sg13g2_nor2_1 _13187_ (.A(_05945_),
    .B(_05948_),
    .Y(_05956_));
 sg13g2_nand2_1 _13188_ (.Y(_05957_),
    .A(_05915_),
    .B(_05938_));
 sg13g2_o21ai_1 _13189_ (.B1(_05957_),
    .Y(_05958_),
    .A1(_00582_),
    .A2(_05938_));
 sg13g2_nor2_1 _13190_ (.A(\vgadonut.donut.cB[13] ),
    .B(net1873),
    .Y(_05959_));
 sg13g2_nand2_1 _13191_ (.Y(_05960_),
    .A(\vgadonut.donut.cB[13] ),
    .B(net1873));
 sg13g2_nand2b_1 _13192_ (.Y(_05961_),
    .B(_05960_),
    .A_N(_05959_));
 sg13g2_xnor2_1 _13193_ (.Y(_05962_),
    .A(net1859),
    .B(_05961_));
 sg13g2_o21ai_1 _13194_ (.B1(_00125_),
    .Y(_05963_),
    .A1(_00576_),
    .A2(_00587_));
 sg13g2_o21ai_1 _13195_ (.B1(_05963_),
    .Y(_05964_),
    .A1(net1858),
    .A2(_05937_));
 sg13g2_xnor2_1 _13196_ (.Y(_05965_),
    .A(_05962_),
    .B(_05964_));
 sg13g2_xnor2_1 _13197_ (.Y(_05966_),
    .A(_05958_),
    .B(_05965_));
 sg13g2_xnor2_1 _13198_ (.Y(_05967_),
    .A(_05956_),
    .B(_05966_));
 sg13g2_o21ai_1 _13199_ (.B1(net1764),
    .Y(_05968_),
    .A1(_05942_),
    .A2(_05967_));
 sg13g2_a21o_1 _13200_ (.A2(_05967_),
    .A1(_05942_),
    .B1(_05968_),
    .X(_05969_));
 sg13g2_a22oi_1 _13201_ (.Y(_00407_),
    .B1(_05955_),
    .B2(_05969_),
    .A2(net1665),
    .A1(_00590_));
 sg13g2_nor2_1 _13202_ (.A(_05937_),
    .B(_05961_),
    .Y(_05970_));
 sg13g2_a22oi_1 _13203_ (.Y(_05971_),
    .B1(_05963_),
    .B2(_05970_),
    .A2(_05961_),
    .A1(net1859));
 sg13g2_nand2_1 _13204_ (.Y(_05972_),
    .A(net1858),
    .B(_05960_));
 sg13g2_o21ai_1 _13205_ (.B1(_05972_),
    .Y(_05973_),
    .A1(net1858),
    .A2(_05959_));
 sg13g2_nor2_1 _13206_ (.A(net1862),
    .B(net1871),
    .Y(_05974_));
 sg13g2_nand2_1 _13207_ (.Y(_05975_),
    .A(net1862),
    .B(net1871));
 sg13g2_nor2b_1 _13208_ (.A(_05974_),
    .B_N(_05975_),
    .Y(_05976_));
 sg13g2_xnor2_1 _13209_ (.Y(_05977_),
    .A(_00582_),
    .B(_05976_));
 sg13g2_xnor2_1 _13210_ (.Y(_05978_),
    .A(_05973_),
    .B(_05977_));
 sg13g2_nand2b_1 _13211_ (.Y(_05979_),
    .B(_05971_),
    .A_N(_05978_));
 sg13g2_xor2_1 _13212_ (.B(_05978_),
    .A(_05971_),
    .X(_05980_));
 sg13g2_nor3_1 _13213_ (.A(_05958_),
    .B(_05965_),
    .C(_05980_),
    .Y(_05981_));
 sg13g2_o21ai_1 _13214_ (.B1(_05980_),
    .Y(_05982_),
    .A1(_05958_),
    .A2(_05965_));
 sg13g2_nor2b_1 _13215_ (.A(_05981_),
    .B_N(_05982_),
    .Y(_05983_));
 sg13g2_o21ai_1 _13216_ (.B1(_05966_),
    .Y(_05984_),
    .A1(_05946_),
    .A2(_05947_));
 sg13g2_nand2b_1 _13217_ (.Y(_05985_),
    .B(_05984_),
    .A_N(_05942_));
 sg13g2_o21ai_1 _13218_ (.B1(_05985_),
    .Y(_05986_),
    .A1(_05956_),
    .A2(_05966_));
 sg13g2_and2_1 _13219_ (.A(_05983_),
    .B(_05986_),
    .X(_05987_));
 sg13g2_nor2b_1 _13220_ (.A(_05987_),
    .B_N(net1763),
    .Y(_05988_));
 sg13g2_o21ai_1 _13221_ (.B1(_05988_),
    .Y(_05989_),
    .A1(_05983_),
    .A2(_05986_));
 sg13g2_xnor2_1 _13222_ (.Y(_05990_),
    .A(net1859),
    .B(\vgadonut.donut.donuthit.rxin[14] ));
 sg13g2_nand3b_1 _13223_ (.B(_05933_),
    .C(_05952_),
    .Y(_05991_),
    .A_N(_05931_));
 sg13g2_o21ai_1 _13224_ (.B1(net1859),
    .Y(_05992_),
    .A1(\vgadonut.donut.donuthit.rxin[12] ),
    .A2(\vgadonut.donut.donuthit.rxin[13] ));
 sg13g2_nand3_1 _13225_ (.B(_05991_),
    .C(_05992_),
    .A(_05932_),
    .Y(_05993_));
 sg13g2_nand2b_1 _13226_ (.Y(_05994_),
    .B(_05993_),
    .A_N(_05990_));
 sg13g2_xnor2_1 _13227_ (.Y(_05995_),
    .A(_05990_),
    .B(_05993_));
 sg13g2_a21oi_1 _13228_ (.A1(net1754),
    .A2(_05995_),
    .Y(_05996_),
    .B1(net1664));
 sg13g2_a22oi_1 _13229_ (.Y(_00408_),
    .B1(_05989_),
    .B2(_05996_),
    .A2(net1664),
    .A1(_00591_));
 sg13g2_o21ai_1 _13230_ (.B1(_05994_),
    .Y(_05997_),
    .A1(_00582_),
    .A2(_00591_));
 sg13g2_xnor2_1 _13231_ (.Y(_05998_),
    .A(net1859),
    .B(\vgadonut.donut.donuthit.rxin[15] ));
 sg13g2_xnor2_1 _13232_ (.Y(_05999_),
    .A(_05997_),
    .B(_05998_));
 sg13g2_a21oi_1 _13233_ (.A1(net1754),
    .A2(_05999_),
    .Y(_06000_),
    .B1(net1664));
 sg13g2_nor2_1 _13234_ (.A(_05981_),
    .B(_05987_),
    .Y(_06001_));
 sg13g2_nand3b_1 _13235_ (.B(_05972_),
    .C(_05976_),
    .Y(_06002_),
    .A_N(_05959_));
 sg13g2_o21ai_1 _13236_ (.B1(_06002_),
    .Y(_06003_),
    .A1(_00582_),
    .A2(_05976_));
 sg13g2_o21ai_1 _13237_ (.B1(_05975_),
    .Y(_06004_),
    .A1(_00125_),
    .A2(_05974_));
 sg13g2_xnor2_1 _13238_ (.Y(_06005_),
    .A(_04522_),
    .B(_06004_));
 sg13g2_xnor2_1 _13239_ (.Y(_06006_),
    .A(_06003_),
    .B(_06005_));
 sg13g2_xnor2_1 _13240_ (.Y(_06007_),
    .A(_05979_),
    .B(_06006_));
 sg13g2_o21ai_1 _13241_ (.B1(net1749),
    .Y(_06008_),
    .A1(_06001_),
    .A2(_06007_));
 sg13g2_a21o_1 _13242_ (.A2(_06007_),
    .A1(_06001_),
    .B1(_06008_),
    .X(_06009_));
 sg13g2_a22oi_1 _13243_ (.Y(_00409_),
    .B1(_06000_),
    .B2(_06009_),
    .A2(net1664),
    .A1(_00593_));
 sg13g2_nand2_1 _13244_ (.Y(_06010_),
    .A(net2141),
    .B(net1735));
 sg13g2_xnor2_1 _13245_ (.Y(_06011_),
    .A(net2141),
    .B(_04547_));
 sg13g2_o21ai_1 _13246_ (.B1(_06010_),
    .Y(_00410_),
    .A1(net1565),
    .A2(_06011_));
 sg13g2_nand2_1 _13247_ (.Y(_06012_),
    .A(net2168),
    .B(net1734));
 sg13g2_xnor2_1 _13248_ (.Y(_06013_),
    .A(_04549_),
    .B(_04550_));
 sg13g2_o21ai_1 _13249_ (.B1(_06012_),
    .Y(_00411_),
    .A1(net1565),
    .A2(_06013_));
 sg13g2_nand2_1 _13250_ (.Y(_06014_),
    .A(net2265),
    .B(net1732));
 sg13g2_xor2_1 _13251_ (.B(_04552_),
    .A(_04551_),
    .X(_06015_));
 sg13g2_o21ai_1 _13252_ (.B1(_06014_),
    .Y(_00412_),
    .A1(net1564),
    .A2(_06015_));
 sg13g2_nand2_1 _13253_ (.Y(_06016_),
    .A(net2148),
    .B(net1732));
 sg13g2_xnor2_1 _13254_ (.Y(_06017_),
    .A(_04554_),
    .B(_04555_));
 sg13g2_o21ai_1 _13255_ (.B1(_06016_),
    .Y(_00413_),
    .A1(net1564),
    .A2(_06017_));
 sg13g2_nand2_1 _13256_ (.Y(_06018_),
    .A(net1884),
    .B(net1732));
 sg13g2_xnor2_1 _13257_ (.Y(_06019_),
    .A(_04557_),
    .B(_04558_));
 sg13g2_o21ai_1 _13258_ (.B1(_06018_),
    .Y(_00414_),
    .A1(net1564),
    .A2(_06019_));
 sg13g2_nand2_1 _13259_ (.Y(_06020_),
    .A(net2180),
    .B(net1734));
 sg13g2_xor2_1 _13260_ (.B(_04562_),
    .A(_04560_),
    .X(_06021_));
 sg13g2_o21ai_1 _13261_ (.B1(_06020_),
    .Y(_00415_),
    .A1(net1565),
    .A2(_06021_));
 sg13g2_nand2_1 _13262_ (.Y(_06022_),
    .A(net1883),
    .B(net1734));
 sg13g2_xnor2_1 _13263_ (.Y(_06023_),
    .A(_04563_),
    .B(_04564_));
 sg13g2_o21ai_1 _13264_ (.B1(_06022_),
    .Y(_00416_),
    .A1(net1565),
    .A2(_06023_));
 sg13g2_nand2_1 _13265_ (.Y(_06024_),
    .A(net2302),
    .B(net1734));
 sg13g2_xnor2_1 _13266_ (.Y(_06025_),
    .A(_04565_),
    .B(_04566_));
 sg13g2_o21ai_1 _13267_ (.B1(_06024_),
    .Y(_00417_),
    .A1(net1565),
    .A2(_06025_));
 sg13g2_nand2_1 _13268_ (.Y(_06026_),
    .A(net1882),
    .B(net1734));
 sg13g2_xnor2_1 _13269_ (.Y(_06027_),
    .A(_04567_),
    .B(_04568_));
 sg13g2_o21ai_1 _13270_ (.B1(_06026_),
    .Y(_00418_),
    .A1(net1567),
    .A2(_06027_));
 sg13g2_nand2_1 _13271_ (.Y(_06028_),
    .A(net1880),
    .B(net1736));
 sg13g2_nand3_1 _13272_ (.B(_04569_),
    .C(_04570_),
    .A(_04531_),
    .Y(_06029_));
 sg13g2_nand2b_1 _13273_ (.Y(_06030_),
    .B(_06029_),
    .A_N(_04571_));
 sg13g2_o21ai_1 _13274_ (.B1(_06028_),
    .Y(_00419_),
    .A1(net1567),
    .A2(_06030_));
 sg13g2_a21oi_1 _13275_ (.A1(net1777),
    .A2(net1763),
    .Y(_06031_),
    .B1(_00583_));
 sg13g2_xnor2_1 _13276_ (.Y(_06032_),
    .A(_04572_),
    .B(_04573_));
 sg13g2_a21o_1 _13277_ (.A2(_06032_),
    .A1(net1571),
    .B1(_06031_),
    .X(_00420_));
 sg13g2_nand2_1 _13278_ (.Y(_06033_),
    .A(net1877),
    .B(net1736));
 sg13g2_xnor2_1 _13279_ (.Y(_06034_),
    .A(_00129_),
    .B(net1600));
 sg13g2_xnor2_1 _13280_ (.Y(_06035_),
    .A(_04575_),
    .B(_06034_));
 sg13g2_o21ai_1 _13281_ (.B1(_06033_),
    .Y(_00421_),
    .A1(net1567),
    .A2(_06035_));
 sg13g2_nand2_1 _13282_ (.Y(_06036_),
    .A(net1876),
    .B(net1737));
 sg13g2_nand3_1 _13283_ (.B(_04576_),
    .C(_04577_),
    .A(_04529_),
    .Y(_06037_));
 sg13g2_nand2b_1 _13284_ (.Y(_06038_),
    .B(_06037_),
    .A_N(_04578_));
 sg13g2_o21ai_1 _13285_ (.B1(_06036_),
    .Y(_00422_),
    .A1(net1568),
    .A2(_06038_));
 sg13g2_nand2_1 _13286_ (.Y(_06039_),
    .A(net1873),
    .B(net1737));
 sg13g2_nand2b_1 _13287_ (.Y(_06040_),
    .B(_04528_),
    .A_N(_04527_));
 sg13g2_xnor2_1 _13288_ (.Y(_06041_),
    .A(_04579_),
    .B(_06040_));
 sg13g2_o21ai_1 _13289_ (.B1(_06039_),
    .Y(_00423_),
    .A1(net1568),
    .A2(_06041_));
 sg13g2_nand2_1 _13290_ (.Y(_06042_),
    .A(net1871),
    .B(net1737));
 sg13g2_xnor2_1 _13291_ (.Y(_06043_),
    .A(_04526_),
    .B(_04580_));
 sg13g2_o21ai_1 _13292_ (.B1(_06042_),
    .Y(_00424_),
    .A1(net1568),
    .A2(_06043_));
 sg13g2_nand2_1 _13293_ (.Y(_06044_),
    .A(net1870),
    .B(net1737));
 sg13g2_o21ai_1 _13294_ (.B1(_06044_),
    .Y(_00425_),
    .A1(net1733),
    .A2(_04582_));
 sg13g2_xor2_1 _13295_ (.B(net1883),
    .A(net1867),
    .X(_06045_));
 sg13g2_a22oi_1 _13296_ (.Y(_06046_),
    .B1(_04587_),
    .B2(_06045_),
    .A2(_03933_),
    .A1(net1867));
 sg13g2_inv_1 _13297_ (.Y(_00426_),
    .A(_06046_));
 sg13g2_nand2_1 _13298_ (.Y(_06047_),
    .A(net1866),
    .B(net1732));
 sg13g2_xnor2_1 _13299_ (.Y(_06048_),
    .A(_04493_),
    .B(_04494_));
 sg13g2_o21ai_1 _13300_ (.B1(_06047_),
    .Y(_00427_),
    .A1(net1564),
    .A2(_06048_));
 sg13g2_nand2_1 _13301_ (.Y(_06049_),
    .A(net1864),
    .B(net1734));
 sg13g2_xnor2_1 _13302_ (.Y(_06050_),
    .A(_04492_),
    .B(_04496_));
 sg13g2_o21ai_1 _13303_ (.B1(_06049_),
    .Y(_00428_),
    .A1(net1565),
    .A2(_06050_));
 sg13g2_nand2_1 _13304_ (.Y(_06051_),
    .A(net1863),
    .B(net1734));
 sg13g2_xnor2_1 _13305_ (.Y(_06052_),
    .A(_04497_),
    .B(_04498_));
 sg13g2_o21ai_1 _13306_ (.B1(_06051_),
    .Y(_00429_),
    .A1(net1565),
    .A2(_06052_));
 sg13g2_nand2_1 _13307_ (.Y(_06053_),
    .A(net2259),
    .B(net1734));
 sg13g2_xnor2_1 _13308_ (.Y(_06054_),
    .A(_04489_),
    .B(_04499_));
 sg13g2_o21ai_1 _13309_ (.B1(_06053_),
    .Y(_00430_),
    .A1(net1565),
    .A2(_06054_));
 sg13g2_nand2_1 _13310_ (.Y(_06055_),
    .A(net2293),
    .B(net1735));
 sg13g2_xnor2_1 _13311_ (.Y(_06056_),
    .A(_04488_),
    .B(_04501_));
 sg13g2_o21ai_1 _13312_ (.B1(_06055_),
    .Y(_00431_),
    .A1(net1566),
    .A2(_06056_));
 sg13g2_nand2_1 _13313_ (.Y(_06057_),
    .A(net2261),
    .B(net1735));
 sg13g2_o21ai_1 _13314_ (.B1(_06057_),
    .Y(_00432_),
    .A1(_04548_),
    .A2(net1566));
 sg13g2_nand2_1 _13315_ (.Y(_06058_),
    .A(net2233),
    .B(net1735));
 sg13g2_o21ai_1 _13316_ (.B1(_06058_),
    .Y(_00433_),
    .A1(_04545_),
    .A2(net1566));
 sg13g2_a22oi_1 _13317_ (.Y(_06059_),
    .B1(_04543_),
    .B2(_04587_),
    .A2(_03930_),
    .A1(net2242));
 sg13g2_inv_1 _13318_ (.Y(_00434_),
    .A(_06059_));
 sg13g2_nand2_1 _13319_ (.Y(_06060_),
    .A(net2205),
    .B(net1735));
 sg13g2_o21ai_1 _13320_ (.B1(_06060_),
    .Y(_00435_),
    .A1(_04541_),
    .A2(net1566));
 sg13g2_nand2_1 _13321_ (.Y(_06061_),
    .A(net2224),
    .B(net1735));
 sg13g2_o21ai_1 _13322_ (.B1(_06061_),
    .Y(_00436_),
    .A1(_04540_),
    .A2(net1566));
 sg13g2_nand2_1 _13323_ (.Y(_06062_),
    .A(net2176),
    .B(net1735));
 sg13g2_o21ai_1 _13324_ (.B1(_06062_),
    .Y(_00437_),
    .A1(_04537_),
    .A2(net1566));
 sg13g2_nand2_1 _13325_ (.Y(_06063_),
    .A(net2248),
    .B(net1736));
 sg13g2_o21ai_1 _13326_ (.B1(_06063_),
    .Y(_00438_),
    .A1(_04535_),
    .A2(net1567));
 sg13g2_a22oi_1 _13327_ (.Y(_06064_),
    .B1(_04533_),
    .B2(_04587_),
    .A2(_03930_),
    .A1(net2268));
 sg13g2_inv_1 _13328_ (.Y(_00439_),
    .A(_06064_));
 sg13g2_nand2_1 _13329_ (.Y(_06065_),
    .A(net1451),
    .B(net1735));
 sg13g2_o21ai_1 _13330_ (.B1(_06065_),
    .Y(_00440_),
    .A1(_04530_),
    .A2(net1566));
 sg13g2_nand2_1 _13331_ (.Y(_06066_),
    .A(net1861),
    .B(net1736));
 sg13g2_o21ai_1 _13332_ (.B1(_06066_),
    .Y(_00441_),
    .A1(_04524_),
    .A2(net1566));
 sg13g2_nor2_1 _13333_ (.A(net2004),
    .B(net1672),
    .Y(_06067_));
 sg13g2_a21oi_1 _13334_ (.A1(_00645_),
    .A2(net1671),
    .Y(_00442_),
    .B1(_06067_));
 sg13g2_nand2_1 _13335_ (.Y(_06068_),
    .A(net1461),
    .B(net1727));
 sg13g2_xnor2_1 _13336_ (.Y(_06069_),
    .A(net1842),
    .B(\vgadonut.donut.cA[4] ));
 sg13g2_nor2_1 _13337_ (.A(net1844),
    .B(_00603_),
    .Y(_06070_));
 sg13g2_xnor2_1 _13338_ (.Y(_06071_),
    .A(net1844),
    .B(\vgadonut.donut.cA[3] ));
 sg13g2_xnor2_1 _13339_ (.Y(_06072_),
    .A(net1846),
    .B(net1825));
 sg13g2_nor2b_1 _13340_ (.A(net1849),
    .B_N(\vgadonut.donut.cA[1] ),
    .Y(_06073_));
 sg13g2_xnor2_1 _13341_ (.Y(_06074_),
    .A(net1849),
    .B(\vgadonut.donut.cA[1] ));
 sg13g2_nand2b_1 _13342_ (.Y(_06075_),
    .B(net1850),
    .A_N(\vgadonut.donut.cA[0] ));
 sg13g2_a21oi_1 _13343_ (.A1(_06074_),
    .A2(_06075_),
    .Y(_06076_),
    .B1(_06073_));
 sg13g2_nor2b_1 _13344_ (.A(_06076_),
    .B_N(_06072_),
    .Y(_06077_));
 sg13g2_a21oi_2 _13345_ (.B1(_06077_),
    .Y(_06078_),
    .A2(net1825),
    .A1(_00594_));
 sg13g2_nor2b_1 _13346_ (.A(_06078_),
    .B_N(_06071_),
    .Y(_06079_));
 sg13g2_o21ai_1 _13347_ (.B1(_06069_),
    .Y(_06080_),
    .A1(_06070_),
    .A2(_06079_));
 sg13g2_o21ai_1 _13348_ (.B1(_06080_),
    .Y(_06081_),
    .A1(net1842),
    .A2(_00602_));
 sg13g2_xor2_1 _13349_ (.B(\vgadonut.donut.cA[5] ),
    .A(net1840),
    .X(_06082_));
 sg13g2_xnor2_1 _13350_ (.Y(_06083_),
    .A(_06081_),
    .B(_06082_));
 sg13g2_nand2_1 _13351_ (.Y(_06084_),
    .A(\vgadonut.donut.sA[0] ),
    .B(_06083_));
 sg13g2_xor2_1 _13352_ (.B(_06083_),
    .A(\vgadonut.donut.sA[0] ),
    .X(_06085_));
 sg13g2_o21ai_1 _13353_ (.B1(_06068_),
    .Y(_00443_),
    .A1(net1560),
    .A2(_06085_));
 sg13g2_nand2_1 _13354_ (.Y(_06086_),
    .A(net1466),
    .B(net1727));
 sg13g2_nor2_1 _13355_ (.A(net1837),
    .B(_00600_),
    .Y(_06087_));
 sg13g2_nand2_1 _13356_ (.Y(_06088_),
    .A(net1837),
    .B(_00600_));
 sg13g2_nand2b_1 _13357_ (.Y(_06089_),
    .B(_06088_),
    .A_N(_06087_));
 sg13g2_a21oi_1 _13358_ (.A1(_00596_),
    .A2(\vgadonut.donut.cA[5] ),
    .Y(_06090_),
    .B1(_06081_));
 sg13g2_a21oi_1 _13359_ (.A1(net1840),
    .A2(_00601_),
    .Y(_06091_),
    .B1(_06090_));
 sg13g2_xnor2_1 _13360_ (.Y(_06092_),
    .A(_06089_),
    .B(_06091_));
 sg13g2_xnor2_1 _13361_ (.Y(_06093_),
    .A(\vgadonut.donut.sA[1] ),
    .B(_06092_));
 sg13g2_nor2_1 _13362_ (.A(_06084_),
    .B(_06093_),
    .Y(_06094_));
 sg13g2_xor2_1 _13363_ (.B(_06093_),
    .A(_06084_),
    .X(_06095_));
 sg13g2_o21ai_1 _13364_ (.B1(_06086_),
    .Y(_00444_),
    .A1(net1560),
    .A2(_06095_));
 sg13g2_nand2_1 _13365_ (.Y(_06096_),
    .A(net1459),
    .B(net1727));
 sg13g2_a21oi_1 _13366_ (.A1(\vgadonut.donut.sA[1] ),
    .A2(_06092_),
    .Y(_06097_),
    .B1(_06094_));
 sg13g2_xnor2_1 _13367_ (.Y(_06098_),
    .A(net1834),
    .B(net1824));
 sg13g2_a21oi_1 _13368_ (.A1(_06088_),
    .A2(_06091_),
    .Y(_06099_),
    .B1(_06087_));
 sg13g2_nand2b_1 _13369_ (.Y(_06100_),
    .B(_06098_),
    .A_N(_06099_));
 sg13g2_xnor2_1 _13370_ (.Y(_06101_),
    .A(_06098_),
    .B(_06099_));
 sg13g2_inv_1 _13371_ (.Y(_06102_),
    .A(_06101_));
 sg13g2_and2_1 _13372_ (.A(net1854),
    .B(_06101_),
    .X(_06103_));
 sg13g2_xnor2_1 _13373_ (.Y(_06104_),
    .A(net1854),
    .B(_06101_));
 sg13g2_nor2_1 _13374_ (.A(_06097_),
    .B(_06104_),
    .Y(_06105_));
 sg13g2_xor2_1 _13375_ (.B(_06104_),
    .A(_06097_),
    .X(_06106_));
 sg13g2_o21ai_1 _13376_ (.B1(_06096_),
    .Y(_00445_),
    .A1(net1560),
    .A2(_06106_));
 sg13g2_nor2b_1 _13377_ (.A(net1832),
    .B_N(\vgadonut.donut.cA[8] ),
    .Y(_06107_));
 sg13g2_xnor2_1 _13378_ (.Y(_06108_),
    .A(net1832),
    .B(\vgadonut.donut.cA[8] ));
 sg13g2_o21ai_1 _13379_ (.B1(_06100_),
    .Y(_06109_),
    .A1(net1834),
    .A2(_00604_));
 sg13g2_xor2_1 _13380_ (.B(_06109_),
    .A(_06108_),
    .X(_06110_));
 sg13g2_nand2_1 _13381_ (.Y(_06111_),
    .A(net1853),
    .B(_06110_));
 sg13g2_xor2_1 _13382_ (.B(_06110_),
    .A(net1853),
    .X(_06112_));
 sg13g2_o21ai_1 _13383_ (.B1(_06112_),
    .Y(_06113_),
    .A1(_06103_),
    .A2(_06105_));
 sg13g2_or3_1 _13384_ (.A(_06103_),
    .B(_06105_),
    .C(_06112_),
    .X(_06114_));
 sg13g2_a21oi_1 _13385_ (.A1(_06113_),
    .A2(_06114_),
    .Y(_06115_),
    .B1(net1560));
 sg13g2_a21o_1 _13386_ (.A2(_03930_),
    .A1(net1990),
    .B1(_06115_),
    .X(_00446_));
 sg13g2_nand2_1 _13387_ (.Y(_06116_),
    .A(net1482),
    .B(net1727));
 sg13g2_xnor2_1 _13388_ (.Y(_06117_),
    .A(net1831),
    .B(net1822));
 sg13g2_a21oi_2 _13389_ (.B1(_06107_),
    .Y(_06118_),
    .A2(_06109_),
    .A1(_06108_));
 sg13g2_xnor2_1 _13390_ (.Y(_06119_),
    .A(_06117_),
    .B(_06118_));
 sg13g2_inv_1 _13391_ (.Y(_06120_),
    .A(_06119_));
 sg13g2_xnor2_1 _13392_ (.Y(_06121_),
    .A(net1852),
    .B(_06119_));
 sg13g2_a21oi_1 _13393_ (.A1(_06111_),
    .A2(_06113_),
    .Y(_06122_),
    .B1(_06121_));
 sg13g2_nand3_1 _13394_ (.B(_06113_),
    .C(_06121_),
    .A(_06111_),
    .Y(_06123_));
 sg13g2_nor2b_1 _13395_ (.A(_06122_),
    .B_N(_06123_),
    .Y(_06124_));
 sg13g2_o21ai_1 _13396_ (.B1(_06116_),
    .Y(_00447_),
    .A1(net1560),
    .A2(_06124_));
 sg13g2_nand2_1 _13397_ (.Y(_06125_),
    .A(net1985),
    .B(net1725));
 sg13g2_a21o_1 _13398_ (.A2(_06119_),
    .A1(net1852),
    .B1(_06122_),
    .X(_06126_));
 sg13g2_xnor2_1 _13399_ (.Y(_06127_),
    .A(net1827),
    .B(net1821));
 sg13g2_a21oi_1 _13400_ (.A1(net1831),
    .A2(_00605_),
    .Y(_06128_),
    .B1(_06118_));
 sg13g2_a21oi_1 _13401_ (.A1(_00598_),
    .A2(\vgadonut.donut.cA[9] ),
    .Y(_06129_),
    .B1(_06128_));
 sg13g2_nand2b_1 _13402_ (.Y(_06130_),
    .B(_06127_),
    .A_N(_06129_));
 sg13g2_xnor2_1 _13403_ (.Y(_06131_),
    .A(_06127_),
    .B(_06129_));
 sg13g2_xnor2_1 _13404_ (.Y(_06132_),
    .A(net1850),
    .B(_06131_));
 sg13g2_xnor2_1 _13405_ (.Y(_06133_),
    .A(_06126_),
    .B(_06132_));
 sg13g2_o21ai_1 _13406_ (.B1(_06125_),
    .Y(_00448_),
    .A1(net1559),
    .A2(_06133_));
 sg13g2_nand2_1 _13407_ (.Y(_06134_),
    .A(net1848),
    .B(net1725));
 sg13g2_nor2_1 _13408_ (.A(net1797),
    .B(net1819),
    .Y(_06135_));
 sg13g2_xor2_1 _13409_ (.B(net1819),
    .A(net1826),
    .X(_06136_));
 sg13g2_o21ai_1 _13410_ (.B1(_06130_),
    .Y(_06137_),
    .A1(net1826),
    .A2(_00606_));
 sg13g2_xnor2_1 _13411_ (.Y(_06138_),
    .A(_06136_),
    .B(_06137_));
 sg13g2_xnor2_1 _13412_ (.Y(_06139_),
    .A(net1848),
    .B(_06138_));
 sg13g2_a21o_1 _13413_ (.A2(_06131_),
    .A1(net1850),
    .B1(_06126_),
    .X(_06140_));
 sg13g2_o21ai_1 _13414_ (.B1(_06140_),
    .Y(_06141_),
    .A1(net1850),
    .A2(_06131_));
 sg13g2_nor2_1 _13415_ (.A(_06139_),
    .B(_06141_),
    .Y(_06142_));
 sg13g2_xnor2_1 _13416_ (.Y(_06143_),
    .A(_06139_),
    .B(_06141_));
 sg13g2_o21ai_1 _13417_ (.B1(_06134_),
    .Y(_00449_),
    .A1(net1559),
    .A2(_06143_));
 sg13g2_nand2_1 _13418_ (.Y(_06144_),
    .A(net1846),
    .B(net1724));
 sg13g2_a21oi_1 _13419_ (.A1(net1848),
    .A2(_06138_),
    .Y(_06145_),
    .B1(_06142_));
 sg13g2_xnor2_1 _13420_ (.Y(_06146_),
    .A(net1826),
    .B(net1817));
 sg13g2_o21ai_1 _13421_ (.B1(net1797),
    .Y(_06147_),
    .A1(net1821),
    .A2(net1819));
 sg13g2_o21ai_1 _13422_ (.B1(_06147_),
    .Y(_06148_),
    .A1(_06130_),
    .A2(_06135_));
 sg13g2_and2_1 _13423_ (.A(_06146_),
    .B(_06148_),
    .X(_06149_));
 sg13g2_xor2_1 _13424_ (.B(_06148_),
    .A(_06146_),
    .X(_06150_));
 sg13g2_inv_1 _13425_ (.Y(_06151_),
    .A(_06150_));
 sg13g2_nand2_1 _13426_ (.Y(_06152_),
    .A(net1846),
    .B(_06150_));
 sg13g2_xnor2_1 _13427_ (.Y(_06153_),
    .A(net1846),
    .B(_06150_));
 sg13g2_or2_1 _13428_ (.X(_06154_),
    .B(_06153_),
    .A(_06145_));
 sg13g2_xnor2_1 _13429_ (.Y(_06155_),
    .A(_06145_),
    .B(_06153_));
 sg13g2_o21ai_1 _13430_ (.B1(_06144_),
    .Y(_00450_),
    .A1(net1557),
    .A2(_06155_));
 sg13g2_nand2_1 _13431_ (.Y(_06156_),
    .A(net1471),
    .B(net1725));
 sg13g2_xnor2_1 _13432_ (.Y(_06157_),
    .A(net1826),
    .B(net1815));
 sg13g2_a21oi_1 _13433_ (.A1(net1797),
    .A2(net1817),
    .Y(_06158_),
    .B1(_06149_));
 sg13g2_xnor2_1 _13434_ (.Y(_06159_),
    .A(_06157_),
    .B(_06158_));
 sg13g2_xnor2_1 _13435_ (.Y(_06160_),
    .A(net1844),
    .B(_06159_));
 sg13g2_a21oi_1 _13436_ (.A1(_06152_),
    .A2(_06154_),
    .Y(_06161_),
    .B1(_06160_));
 sg13g2_nand3_1 _13437_ (.B(_06154_),
    .C(_06160_),
    .A(_06152_),
    .Y(_06162_));
 sg13g2_nor2b_1 _13438_ (.A(_06161_),
    .B_N(_06162_),
    .Y(_06163_));
 sg13g2_o21ai_1 _13439_ (.B1(_06156_),
    .Y(_00451_),
    .A1(net1559),
    .A2(_06163_));
 sg13g2_nand2_1 _13440_ (.Y(_06164_),
    .A(net1843),
    .B(net1724));
 sg13g2_a21o_1 _13441_ (.A2(_06159_),
    .A1(net1844),
    .B1(_06161_),
    .X(_06165_));
 sg13g2_o21ai_1 _13442_ (.B1(_06149_),
    .Y(_06166_),
    .A1(net1797),
    .A2(net1815));
 sg13g2_o21ai_1 _13443_ (.B1(net1797),
    .Y(_06167_),
    .A1(net1817),
    .A2(net1815));
 sg13g2_nand2_1 _13444_ (.Y(_06168_),
    .A(_06166_),
    .B(_06167_));
 sg13g2_nor2b_1 _13445_ (.A(net1826),
    .B_N(net1814),
    .Y(_06169_));
 sg13g2_xnor2_1 _13446_ (.Y(_06170_),
    .A(net1826),
    .B(net1814));
 sg13g2_xnor2_1 _13447_ (.Y(_06171_),
    .A(_06168_),
    .B(_06170_));
 sg13g2_nor2_1 _13448_ (.A(_00595_),
    .B(_06171_),
    .Y(_06172_));
 sg13g2_nand2_1 _13449_ (.Y(_06173_),
    .A(_00595_),
    .B(_06171_));
 sg13g2_nor2b_1 _13450_ (.A(_06172_),
    .B_N(_06173_),
    .Y(_06174_));
 sg13g2_xnor2_1 _13451_ (.Y(_06175_),
    .A(_06165_),
    .B(_06174_));
 sg13g2_o21ai_1 _13452_ (.B1(_06164_),
    .Y(_00452_),
    .A1(net1557),
    .A2(_06175_));
 sg13g2_nand2_1 _13453_ (.Y(_06176_),
    .A(net1470),
    .B(net1724));
 sg13g2_a21oi_1 _13454_ (.A1(_06168_),
    .A2(_06170_),
    .Y(_06177_),
    .B1(_06169_));
 sg13g2_xnor2_1 _13455_ (.Y(_06178_),
    .A(net1813),
    .B(_06177_));
 sg13g2_xnor2_1 _13456_ (.Y(_06179_),
    .A(net1797),
    .B(_06178_));
 sg13g2_nor2b_1 _13457_ (.A(net1840),
    .B_N(net1602),
    .Y(_06180_));
 sg13g2_nand2b_1 _13458_ (.Y(_06181_),
    .B(net1840),
    .A_N(net1602));
 sg13g2_nor2b_1 _13459_ (.A(_06180_),
    .B_N(_06181_),
    .Y(_06182_));
 sg13g2_a21oi_1 _13460_ (.A1(_06165_),
    .A2(_06173_),
    .Y(_06183_),
    .B1(_06172_));
 sg13g2_xnor2_1 _13461_ (.Y(_06184_),
    .A(_06182_),
    .B(_06183_));
 sg13g2_o21ai_1 _13462_ (.B1(_06176_),
    .Y(_00453_),
    .A1(net1557),
    .A2(_06184_));
 sg13g2_nand2_1 _13463_ (.Y(_06185_),
    .A(net1491),
    .B(net1724));
 sg13g2_nand2b_1 _13464_ (.Y(_06186_),
    .B(net1602),
    .A_N(net1838));
 sg13g2_nor2b_1 _13465_ (.A(net1602),
    .B_N(net1838),
    .Y(_06187_));
 sg13g2_xor2_1 _13466_ (.B(net1602),
    .A(net1838),
    .X(_06188_));
 sg13g2_o21ai_1 _13467_ (.B1(_06181_),
    .Y(_06189_),
    .A1(_06180_),
    .A2(_06183_));
 sg13g2_xnor2_1 _13468_ (.Y(_06190_),
    .A(_06188_),
    .B(_06189_));
 sg13g2_o21ai_1 _13469_ (.B1(_06185_),
    .Y(_00454_),
    .A1(net1557),
    .A2(_06190_));
 sg13g2_nand2_1 _13470_ (.Y(_06191_),
    .A(net1835),
    .B(net1724));
 sg13g2_nand2b_1 _13471_ (.Y(_06192_),
    .B(net1835),
    .A_N(net1602));
 sg13g2_nor2b_1 _13472_ (.A(net1834),
    .B_N(net1602),
    .Y(_06193_));
 sg13g2_xnor2_1 _13473_ (.Y(_06194_),
    .A(net1834),
    .B(net1602));
 sg13g2_a21oi_1 _13474_ (.A1(_06186_),
    .A2(_06189_),
    .Y(_06195_),
    .B1(_06187_));
 sg13g2_xor2_1 _13475_ (.B(_06195_),
    .A(_06194_),
    .X(_06196_));
 sg13g2_o21ai_1 _13476_ (.B1(_06191_),
    .Y(_00455_),
    .A1(net1557),
    .A2(_06196_));
 sg13g2_nand2_1 _13477_ (.Y(_06197_),
    .A(net1490),
    .B(net1724));
 sg13g2_nand2_1 _13478_ (.Y(_06198_),
    .A(_00597_),
    .B(net1603));
 sg13g2_nor2_1 _13479_ (.A(_00597_),
    .B(net1603),
    .Y(_06199_));
 sg13g2_xnor2_1 _13480_ (.Y(_06200_),
    .A(_00597_),
    .B(net1603));
 sg13g2_o21ai_1 _13481_ (.B1(_06192_),
    .Y(_06201_),
    .A1(_06193_),
    .A2(_06195_));
 sg13g2_xnor2_1 _13482_ (.Y(_06202_),
    .A(_06200_),
    .B(_06201_));
 sg13g2_o21ai_1 _13483_ (.B1(_06197_),
    .Y(_00456_),
    .A1(net1557),
    .A2(_06202_));
 sg13g2_nand2_1 _13484_ (.Y(_06203_),
    .A(net1831),
    .B(net1724));
 sg13g2_or2_1 _13485_ (.X(_06204_),
    .B(net1603),
    .A(net2311));
 sg13g2_xnor2_1 _13486_ (.Y(_06205_),
    .A(net2311),
    .B(net1603));
 sg13g2_o21ai_1 _13487_ (.B1(_06198_),
    .Y(_06206_),
    .A1(_06199_),
    .A2(_06201_));
 sg13g2_xnor2_1 _13488_ (.Y(_06207_),
    .A(_06205_),
    .B(_06206_));
 sg13g2_o21ai_1 _13489_ (.B1(_06203_),
    .Y(_00457_),
    .A1(net1558),
    .A2(_06207_));
 sg13g2_nand2_1 _13490_ (.Y(_06208_),
    .A(net1829),
    .B(net1725));
 sg13g2_o21ai_1 _13491_ (.B1(_06204_),
    .Y(_06209_),
    .A1(_06205_),
    .A2(_06206_));
 sg13g2_xor2_1 _13492_ (.B(_06209_),
    .A(_06178_),
    .X(_06210_));
 sg13g2_o21ai_1 _13493_ (.B1(_06208_),
    .Y(_00458_),
    .A1(net1558),
    .A2(_06210_));
 sg13g2_nand2_1 _13494_ (.Y(_06211_),
    .A(net1483),
    .B(net1717));
 sg13g2_xor2_1 _13495_ (.B(\vgadonut.donut.cA[0] ),
    .A(net1850),
    .X(_06212_));
 sg13g2_o21ai_1 _13496_ (.B1(_06211_),
    .Y(_00459_),
    .A1(net1551),
    .A2(_06212_));
 sg13g2_nand2_1 _13497_ (.Y(_06213_),
    .A(net1488),
    .B(net1717));
 sg13g2_xor2_1 _13498_ (.B(_06075_),
    .A(_06074_),
    .X(_06214_));
 sg13g2_o21ai_1 _13499_ (.B1(_06213_),
    .Y(_00460_),
    .A1(net1551),
    .A2(_06214_));
 sg13g2_nand2_1 _13500_ (.Y(_06215_),
    .A(net1485),
    .B(net1717));
 sg13g2_xnor2_1 _13501_ (.Y(_06216_),
    .A(_06072_),
    .B(_06076_));
 sg13g2_o21ai_1 _13502_ (.B1(_06215_),
    .Y(_00461_),
    .A1(net1551),
    .A2(_06216_));
 sg13g2_nand2_1 _13503_ (.Y(_06217_),
    .A(net1486),
    .B(net1717));
 sg13g2_xnor2_1 _13504_ (.Y(_06218_),
    .A(_06071_),
    .B(_06078_));
 sg13g2_o21ai_1 _13505_ (.B1(_06217_),
    .Y(_00462_),
    .A1(net1551),
    .A2(_06218_));
 sg13g2_nand2_1 _13506_ (.Y(_06219_),
    .A(net1481),
    .B(net1717));
 sg13g2_or3_1 _13507_ (.A(_06069_),
    .B(_06070_),
    .C(_06079_),
    .X(_06220_));
 sg13g2_and2_1 _13508_ (.A(_06080_),
    .B(_06220_),
    .X(_06221_));
 sg13g2_o21ai_1 _13509_ (.B1(_06219_),
    .Y(_00463_),
    .A1(net1551),
    .A2(_06221_));
 sg13g2_nand2_1 _13510_ (.Y(_06222_),
    .A(net1463),
    .B(net1727));
 sg13g2_o21ai_1 _13511_ (.B1(_06222_),
    .Y(_00464_),
    .A1(net1560),
    .A2(_06083_));
 sg13g2_a21oi_1 _13512_ (.A1(net1775),
    .A2(net1762),
    .Y(_06223_),
    .B1(_00600_));
 sg13g2_a21o_1 _13513_ (.A2(_06092_),
    .A1(net1570),
    .B1(_06223_),
    .X(_00465_));
 sg13g2_nand2_1 _13514_ (.Y(_06224_),
    .A(net1824),
    .B(net1727));
 sg13g2_o21ai_1 _13515_ (.B1(_06224_),
    .Y(_00466_),
    .A1(net1560),
    .A2(_06102_));
 sg13g2_nand2_1 _13516_ (.Y(_06225_),
    .A(net1487),
    .B(net1727));
 sg13g2_o21ai_1 _13517_ (.B1(_06225_),
    .Y(_00467_),
    .A1(net1560),
    .A2(_06110_));
 sg13g2_nand2_1 _13518_ (.Y(_06226_),
    .A(net2039),
    .B(net1726));
 sg13g2_o21ai_1 _13519_ (.B1(_06226_),
    .Y(_00468_),
    .A1(net1563),
    .A2(_06120_));
 sg13g2_nand2_1 _13520_ (.Y(_06227_),
    .A(net1465),
    .B(net1726));
 sg13g2_o21ai_1 _13521_ (.B1(_06227_),
    .Y(_00469_),
    .A1(net1563),
    .A2(_06131_));
 sg13g2_nand2_1 _13522_ (.Y(_06228_),
    .A(net1473),
    .B(net1726));
 sg13g2_o21ai_1 _13523_ (.B1(_06228_),
    .Y(_00470_),
    .A1(net1559),
    .A2(_06138_));
 sg13g2_nand2_1 _13524_ (.Y(_06229_),
    .A(net1817),
    .B(net1725));
 sg13g2_o21ai_1 _13525_ (.B1(_06229_),
    .Y(_00471_),
    .A1(net1558),
    .A2(_06151_));
 sg13g2_nand2_1 _13526_ (.Y(_06230_),
    .A(net1464),
    .B(net1725));
 sg13g2_o21ai_1 _13527_ (.B1(_06230_),
    .Y(_00472_),
    .A1(net1557),
    .A2(_06159_));
 sg13g2_nand2_1 _13528_ (.Y(_06231_),
    .A(net1814),
    .B(net1724));
 sg13g2_o21ai_1 _13529_ (.B1(_06231_),
    .Y(_00473_),
    .A1(net1557),
    .A2(_06171_));
 sg13g2_nand2_1 _13530_ (.Y(_06232_),
    .A(net1813),
    .B(net1725));
 sg13g2_o21ai_1 _13531_ (.B1(_06232_),
    .Y(_00474_),
    .A1(net1558),
    .A2(net1603));
 sg13g2_a221oi_1 _13532_ (.B2(_00683_),
    .C1(net1642),
    .B1(_00740_),
    .A1(net1646),
    .Y(_00475_),
    .A2(_00734_));
 sg13g2_nor2b_1 _13533_ (.A(_04021_),
    .B_N(_04032_),
    .Y(_06233_));
 sg13g2_nand4_1 _13534_ (.B(_04038_),
    .C(_04043_),
    .A(_04005_),
    .Y(_06234_),
    .D(_06233_));
 sg13g2_a21oi_1 _13535_ (.A1(net2355),
    .A2(_04040_),
    .Y(_06235_),
    .B1(_04042_));
 sg13g2_nand2_2 _13536_ (.Y(_06236_),
    .A(_06234_),
    .B(_06235_));
 sg13g2_a21o_1 _13537_ (.A2(_06236_),
    .A1(net2004),
    .B1(net1689),
    .X(_00476_));
 sg13g2_nand2_1 _13538_ (.Y(_06237_),
    .A(\vgadonut.donut.rz6[0] ),
    .B(net1912));
 sg13g2_or2_1 _13539_ (.X(_06238_),
    .B(net1912),
    .A(\vgadonut.donut.rz6[0] ));
 sg13g2_nand3_1 _13540_ (.B(_06237_),
    .C(_06238_),
    .A(net1743),
    .Y(_06239_));
 sg13g2_nand2_1 _13541_ (.Y(_06240_),
    .A(\vgadonut.donut.ysA[0] ),
    .B(net1749));
 sg13g2_a21oi_1 _13542_ (.A1(_06239_),
    .A2(_06240_),
    .Y(_06241_),
    .B1(net1651));
 sg13g2_a21o_1 _13543_ (.A2(net1651),
    .A1(net2015),
    .B1(_06241_),
    .X(_00477_));
 sg13g2_nand2_1 _13544_ (.Y(_06242_),
    .A(\vgadonut.donut.rz6[1] ),
    .B(net1911));
 sg13g2_xnor2_1 _13545_ (.Y(_06243_),
    .A(\vgadonut.donut.rz6[1] ),
    .B(net1911));
 sg13g2_xnor2_1 _13546_ (.Y(_06244_),
    .A(_06237_),
    .B(_06243_));
 sg13g2_nor2_1 _13547_ (.A(net1762),
    .B(_06244_),
    .Y(_06245_));
 sg13g2_a21oi_1 _13548_ (.A1(\vgadonut.donut.ysA[1] ),
    .A2(net1762),
    .Y(_06246_),
    .B1(_06245_));
 sg13g2_nand2_1 _13549_ (.Y(_06247_),
    .A(net1999),
    .B(net1651));
 sg13g2_o21ai_1 _13550_ (.B1(_06247_),
    .Y(_00478_),
    .A1(net1651),
    .A2(_06246_));
 sg13g2_nand2_1 _13551_ (.Y(_06248_),
    .A(\vgadonut.donut.rz6[2] ),
    .B(net1910));
 sg13g2_xor2_1 _13552_ (.B(net1910),
    .A(\vgadonut.donut.rz6[2] ),
    .X(_06249_));
 sg13g2_o21ai_1 _13553_ (.B1(_06242_),
    .Y(_06250_),
    .A1(_06237_),
    .A2(_06243_));
 sg13g2_nand2_1 _13554_ (.Y(_06251_),
    .A(_06249_),
    .B(_06250_));
 sg13g2_xor2_1 _13555_ (.B(_06250_),
    .A(_06249_),
    .X(_06252_));
 sg13g2_nand2b_1 _13556_ (.Y(_06253_),
    .B(net2360),
    .A_N(net1912));
 sg13g2_nor2b_1 _13557_ (.A(\vgadonut.donut.ysA[2] ),
    .B_N(net1912),
    .Y(_06254_));
 sg13g2_nand3b_1 _13558_ (.B(net1762),
    .C(_06253_),
    .Y(_06255_),
    .A_N(_06254_));
 sg13g2_o21ai_1 _13559_ (.B1(_06255_),
    .Y(_06256_),
    .A1(net1757),
    .A2(_06252_));
 sg13g2_nand2_1 _13560_ (.Y(_06257_),
    .A(net1996),
    .B(net1651));
 sg13g2_o21ai_1 _13561_ (.B1(_06257_),
    .Y(_00479_),
    .A1(net1651),
    .A2(_06256_));
 sg13g2_xnor2_1 _13562_ (.Y(_06258_),
    .A(\vgadonut.donut.rz6[3] ),
    .B(net1909));
 sg13g2_a21oi_1 _13563_ (.A1(_06248_),
    .A2(_06251_),
    .Y(_06259_),
    .B1(_06258_));
 sg13g2_nand3_1 _13564_ (.B(_06251_),
    .C(_06258_),
    .A(_06248_),
    .Y(_06260_));
 sg13g2_nand2b_1 _13565_ (.Y(_06261_),
    .B(_06260_),
    .A_N(_06259_));
 sg13g2_nand2_1 _13566_ (.Y(_06262_),
    .A(net1912),
    .B(net1911));
 sg13g2_xnor2_1 _13567_ (.Y(_06263_),
    .A(net1912),
    .B(net1911));
 sg13g2_nor2_2 _13568_ (.A(\vgadonut.donut.ysA[3] ),
    .B(_06263_),
    .Y(_06264_));
 sg13g2_xnor2_1 _13569_ (.Y(_06265_),
    .A(_06850_),
    .B(_06263_));
 sg13g2_nor2_1 _13570_ (.A(_06254_),
    .B(_06265_),
    .Y(_06266_));
 sg13g2_nand2_1 _13571_ (.Y(_06267_),
    .A(_06254_),
    .B(_06265_));
 sg13g2_nor2_1 _13572_ (.A(net1742),
    .B(_06266_),
    .Y(_06268_));
 sg13g2_a22oi_1 _13573_ (.Y(_06269_),
    .B1(_06267_),
    .B2(_06268_),
    .A2(_06261_),
    .A1(net1752));
 sg13g2_mux2_1 _13574_ (.A0(net2037),
    .A1(_06269_),
    .S(net1670),
    .X(_00480_));
 sg13g2_xnor2_1 _13575_ (.Y(_06270_),
    .A(\vgadonut.donut.rz6[4] ),
    .B(net1908));
 sg13g2_a21oi_1 _13576_ (.A1(\vgadonut.donut.rz6[3] ),
    .A2(net1909),
    .Y(_06271_),
    .B1(_06259_));
 sg13g2_or2_1 _13577_ (.X(_06272_),
    .B(_06271_),
    .A(_06270_));
 sg13g2_a21oi_1 _13578_ (.A1(_06270_),
    .A2(_06271_),
    .Y(_06273_),
    .B1(net1762));
 sg13g2_xnor2_1 _13579_ (.Y(_06274_),
    .A(net1911),
    .B(net1910));
 sg13g2_nand2_1 _13580_ (.Y(_06275_),
    .A(_06262_),
    .B(_06274_));
 sg13g2_o21ai_1 _13581_ (.B1(_06275_),
    .Y(_06276_),
    .A1(net1910),
    .A2(_06262_));
 sg13g2_xnor2_1 _13582_ (.Y(_06277_),
    .A(_06851_),
    .B(_06276_));
 sg13g2_xor2_1 _13583_ (.B(_06277_),
    .A(_06264_),
    .X(_06278_));
 sg13g2_nand2_1 _13584_ (.Y(_06279_),
    .A(_06267_),
    .B(_06278_));
 sg13g2_or2_1 _13585_ (.X(_06280_),
    .B(_06278_),
    .A(_06267_));
 sg13g2_nand3_1 _13586_ (.B(_06279_),
    .C(_06280_),
    .A(net1748),
    .Y(_06281_));
 sg13g2_a21oi_1 _13587_ (.A1(_06272_),
    .A2(_06273_),
    .Y(_06282_),
    .B1(net1652));
 sg13g2_a22oi_1 _13588_ (.Y(_00481_),
    .B1(_06281_),
    .B2(_06282_),
    .A2(net1652),
    .A1(_06852_));
 sg13g2_o21ai_1 _13589_ (.B1(_06272_),
    .Y(_06283_),
    .A1(_06852_),
    .A2(_06853_));
 sg13g2_xnor2_1 _13590_ (.Y(_06284_),
    .A(\vgadonut.donut.rz6[5] ),
    .B(net1907));
 sg13g2_xnor2_1 _13591_ (.Y(_06285_),
    .A(_06283_),
    .B(_06284_));
 sg13g2_a21oi_1 _13592_ (.A1(net1752),
    .A2(_06285_),
    .Y(_06286_),
    .B1(net1651));
 sg13g2_nand2_1 _13593_ (.Y(_06287_),
    .A(net1910),
    .B(net1909));
 sg13g2_or2_1 _13594_ (.X(_06288_),
    .B(net1909),
    .A(net1910));
 sg13g2_a22oi_1 _13595_ (.Y(_06289_),
    .B1(_06287_),
    .B2(_06288_),
    .A2(net1910),
    .A1(net1911));
 sg13g2_nand3b_1 _13596_ (.B(net1910),
    .C(net1911),
    .Y(_06290_),
    .A_N(net1909));
 sg13g2_nor2b_1 _13597_ (.A(_06289_),
    .B_N(_06290_),
    .Y(_06291_));
 sg13g2_xnor2_1 _13598_ (.Y(_06292_),
    .A(\vgadonut.donut.ysA[5] ),
    .B(_06291_));
 sg13g2_o21ai_1 _13599_ (.B1(_06275_),
    .Y(_06293_),
    .A1(_06851_),
    .A2(_06276_));
 sg13g2_nand2b_1 _13600_ (.Y(_06294_),
    .B(_06293_),
    .A_N(_06292_));
 sg13g2_xor2_1 _13601_ (.B(_06293_),
    .A(_06292_),
    .X(_06295_));
 sg13g2_nor3_1 _13602_ (.A(_06264_),
    .B(_06277_),
    .C(_06295_),
    .Y(_06296_));
 sg13g2_o21ai_1 _13603_ (.B1(_06295_),
    .Y(_06297_),
    .A1(_06264_),
    .A2(_06277_));
 sg13g2_nand2b_1 _13604_ (.Y(_06298_),
    .B(_06297_),
    .A_N(_06296_));
 sg13g2_nor2_1 _13605_ (.A(_06279_),
    .B(_06298_),
    .Y(_06299_));
 sg13g2_a21oi_1 _13606_ (.A1(_06279_),
    .A2(_06298_),
    .Y(_06300_),
    .B1(net1750));
 sg13g2_nand2b_1 _13607_ (.Y(_06301_),
    .B(_06300_),
    .A_N(_06299_));
 sg13g2_a22oi_1 _13608_ (.Y(_00482_),
    .B1(_06286_),
    .B2(_06301_),
    .A2(net1651),
    .A1(_06855_));
 sg13g2_and2_1 _13609_ (.A(\vgadonut.donut.donuthit.rzin[0] ),
    .B(net1906),
    .X(_06302_));
 sg13g2_xor2_1 _13610_ (.B(net1906),
    .A(\vgadonut.donut.donuthit.rzin[0] ),
    .X(_06303_));
 sg13g2_a21oi_1 _13611_ (.A1(\vgadonut.donut.rz6[5] ),
    .A2(net1907),
    .Y(_06304_),
    .B1(_06283_));
 sg13g2_a21oi_1 _13612_ (.A1(_06855_),
    .A2(_06856_),
    .Y(_06305_),
    .B1(_06304_));
 sg13g2_xor2_1 _13613_ (.B(_06305_),
    .A(_06303_),
    .X(_06306_));
 sg13g2_a21oi_1 _13614_ (.A1(net1750),
    .A2(_06306_),
    .Y(_06307_),
    .B1(net1657));
 sg13g2_nor2_1 _13615_ (.A(_06296_),
    .B(_06299_),
    .Y(_06308_));
 sg13g2_a21o_1 _13616_ (.A2(_06291_),
    .A1(\vgadonut.donut.ysA[5] ),
    .B1(_06289_),
    .X(_06309_));
 sg13g2_nor2_1 _13617_ (.A(net1909),
    .B(net1908),
    .Y(_06310_));
 sg13g2_xor2_1 _13618_ (.B(net1908),
    .A(net1909),
    .X(_06311_));
 sg13g2_xnor2_1 _13619_ (.Y(_06312_),
    .A(_00094_),
    .B(_06311_));
 sg13g2_nor2b_1 _13620_ (.A(_06312_),
    .B_N(_06287_),
    .Y(_06313_));
 sg13g2_xnor2_1 _13621_ (.Y(_06314_),
    .A(_06287_),
    .B(_06312_));
 sg13g2_xnor2_1 _13622_ (.Y(_06315_),
    .A(\vgadonut.donut.cAcB[0] ),
    .B(_06314_));
 sg13g2_nor2b_1 _13623_ (.A(_06315_),
    .B_N(_06309_),
    .Y(_06316_));
 sg13g2_xnor2_1 _13624_ (.Y(_06317_),
    .A(_06309_),
    .B(_06315_));
 sg13g2_xnor2_1 _13625_ (.Y(_06318_),
    .A(\vgadonut.donut.ysA[6] ),
    .B(_06317_));
 sg13g2_or2_1 _13626_ (.X(_06319_),
    .B(_06318_),
    .A(_06294_));
 sg13g2_xnor2_1 _13627_ (.Y(_06320_),
    .A(_06294_),
    .B(_06318_));
 sg13g2_or2_1 _13628_ (.X(_06321_),
    .B(_06320_),
    .A(_06308_));
 sg13g2_a21oi_1 _13629_ (.A1(_06308_),
    .A2(_06320_),
    .Y(_06322_),
    .B1(net1744));
 sg13g2_nand2_1 _13630_ (.Y(_06323_),
    .A(_06321_),
    .B(_06322_));
 sg13g2_a22oi_1 _13631_ (.Y(_00483_),
    .B1(_06307_),
    .B2(_06323_),
    .A2(net1657),
    .A1(_06857_));
 sg13g2_xnor2_1 _13632_ (.Y(_06324_),
    .A(\vgadonut.donut.donuthit.rzin[1] ),
    .B(net1905));
 sg13g2_a21oi_1 _13633_ (.A1(_06303_),
    .A2(_06305_),
    .Y(_06325_),
    .B1(_06302_));
 sg13g2_nor2_1 _13634_ (.A(_06324_),
    .B(_06325_),
    .Y(_06326_));
 sg13g2_xor2_1 _13635_ (.B(_06325_),
    .A(_06324_),
    .X(_06327_));
 sg13g2_a21oi_1 _13636_ (.A1(net1750),
    .A2(_06327_),
    .Y(_06328_),
    .B1(net1657));
 sg13g2_a21oi_1 _13637_ (.A1(\vgadonut.donut.cAcB[0] ),
    .A2(_06314_),
    .Y(_06329_),
    .B1(_06313_));
 sg13g2_a21oi_1 _13638_ (.A1(_00094_),
    .A2(_06311_),
    .Y(_06330_),
    .B1(_06310_));
 sg13g2_nor2_1 _13639_ (.A(net1908),
    .B(net1907),
    .Y(_06331_));
 sg13g2_xor2_1 _13640_ (.B(net1907),
    .A(net1908),
    .X(_06332_));
 sg13g2_xnor2_1 _13641_ (.Y(_06333_),
    .A(_00095_),
    .B(_06332_));
 sg13g2_nor2_1 _13642_ (.A(_06330_),
    .B(_06333_),
    .Y(_06334_));
 sg13g2_xor2_1 _13643_ (.B(_06333_),
    .A(_06330_),
    .X(_06335_));
 sg13g2_xnor2_1 _13644_ (.Y(_06336_),
    .A(\vgadonut.donut.cAcB[1] ),
    .B(_06335_));
 sg13g2_nor2_1 _13645_ (.A(_06329_),
    .B(_06336_),
    .Y(_06337_));
 sg13g2_xor2_1 _13646_ (.B(_06336_),
    .A(_06329_),
    .X(_06338_));
 sg13g2_xnor2_1 _13647_ (.Y(_06339_),
    .A(\vgadonut.donut.ysA[7] ),
    .B(_06338_));
 sg13g2_a21oi_1 _13648_ (.A1(\vgadonut.donut.ysA[6] ),
    .A2(_06317_),
    .Y(_06340_),
    .B1(_06316_));
 sg13g2_nor2_1 _13649_ (.A(_06339_),
    .B(_06340_),
    .Y(_06341_));
 sg13g2_xnor2_1 _13650_ (.Y(_06342_),
    .A(_06339_),
    .B(_06340_));
 sg13g2_a21o_1 _13651_ (.A2(_06321_),
    .A1(_06319_),
    .B1(_06342_),
    .X(_06343_));
 sg13g2_nand3_1 _13652_ (.B(_06321_),
    .C(_06342_),
    .A(_06319_),
    .Y(_06344_));
 sg13g2_nand3_1 _13653_ (.B(_06343_),
    .C(_06344_),
    .A(net1749),
    .Y(_06345_));
 sg13g2_a22oi_1 _13654_ (.Y(_00484_),
    .B1(_06328_),
    .B2(_06345_),
    .A2(net1657),
    .A1(_06858_));
 sg13g2_xnor2_1 _13655_ (.Y(_06346_),
    .A(\vgadonut.donut.donuthit.rzin[2] ),
    .B(net1904));
 sg13g2_a21oi_1 _13656_ (.A1(\vgadonut.donut.donuthit.rzin[1] ),
    .A2(net1905),
    .Y(_06347_),
    .B1(_06326_));
 sg13g2_nor2_1 _13657_ (.A(_06346_),
    .B(_06347_),
    .Y(_06348_));
 sg13g2_xor2_1 _13658_ (.B(_06347_),
    .A(_06346_),
    .X(_06349_));
 sg13g2_a21oi_1 _13659_ (.A1(net1750),
    .A2(_06349_),
    .Y(_06350_),
    .B1(net1657));
 sg13g2_nor2b_1 _13660_ (.A(_06341_),
    .B_N(_06343_),
    .Y(_06351_));
 sg13g2_a21oi_1 _13661_ (.A1(\vgadonut.donut.cAcB[1] ),
    .A2(_06335_),
    .Y(_06352_),
    .B1(_06334_));
 sg13g2_a21oi_1 _13662_ (.A1(_00095_),
    .A2(_06332_),
    .Y(_06353_),
    .B1(_06331_));
 sg13g2_nor2_1 _13663_ (.A(net1907),
    .B(net1906),
    .Y(_06354_));
 sg13g2_xor2_1 _13664_ (.B(net1906),
    .A(net1907),
    .X(_06355_));
 sg13g2_xnor2_1 _13665_ (.Y(_06356_),
    .A(_00096_),
    .B(_06355_));
 sg13g2_nor2_1 _13666_ (.A(_06353_),
    .B(_06356_),
    .Y(_06357_));
 sg13g2_xor2_1 _13667_ (.B(_06356_),
    .A(_06353_),
    .X(_06358_));
 sg13g2_xnor2_1 _13668_ (.Y(_06359_),
    .A(\vgadonut.donut.cAcB[2] ),
    .B(_06358_));
 sg13g2_nor2_1 _13669_ (.A(_06352_),
    .B(_06359_),
    .Y(_06360_));
 sg13g2_xor2_1 _13670_ (.B(_06359_),
    .A(_06352_),
    .X(_06361_));
 sg13g2_xnor2_1 _13671_ (.Y(_06362_),
    .A(\vgadonut.donut.ysA[8] ),
    .B(_06361_));
 sg13g2_a21oi_1 _13672_ (.A1(\vgadonut.donut.ysA[7] ),
    .A2(_06338_),
    .Y(_06363_),
    .B1(_06337_));
 sg13g2_nor2_1 _13673_ (.A(_06362_),
    .B(_06363_),
    .Y(_06364_));
 sg13g2_xnor2_1 _13674_ (.Y(_06365_),
    .A(_06362_),
    .B(_06363_));
 sg13g2_nor2_1 _13675_ (.A(_06351_),
    .B(_06365_),
    .Y(_06366_));
 sg13g2_a21oi_1 _13676_ (.A1(_06351_),
    .A2(_06365_),
    .Y(_06367_),
    .B1(net1744));
 sg13g2_nand2b_1 _13677_ (.Y(_06368_),
    .B(_06367_),
    .A_N(_06366_));
 sg13g2_a22oi_1 _13678_ (.Y(_00485_),
    .B1(_06350_),
    .B2(_06368_),
    .A2(net1657),
    .A1(_06862_));
 sg13g2_a21oi_1 _13679_ (.A1(\vgadonut.donut.ysA[8] ),
    .A2(_06361_),
    .Y(_06369_),
    .B1(_06360_));
 sg13g2_a21oi_2 _13680_ (.B1(_06357_),
    .Y(_06370_),
    .A2(_06358_),
    .A1(\vgadonut.donut.cAcB[2] ));
 sg13g2_a21oi_2 _13681_ (.B1(_06354_),
    .Y(_06371_),
    .A2(_06355_),
    .A1(_00096_));
 sg13g2_nor2_1 _13682_ (.A(net1906),
    .B(net1905),
    .Y(_06372_));
 sg13g2_xor2_1 _13683_ (.B(net1905),
    .A(net1906),
    .X(_06373_));
 sg13g2_xnor2_1 _13684_ (.Y(_06374_),
    .A(_00097_),
    .B(_06373_));
 sg13g2_nor2_1 _13685_ (.A(_06371_),
    .B(_06374_),
    .Y(_06375_));
 sg13g2_xor2_1 _13686_ (.B(_06374_),
    .A(_06371_),
    .X(_06376_));
 sg13g2_xnor2_1 _13687_ (.Y(_06377_),
    .A(net1957),
    .B(_06376_));
 sg13g2_nor2_1 _13688_ (.A(_06370_),
    .B(_06377_),
    .Y(_06378_));
 sg13g2_xor2_1 _13689_ (.B(_06377_),
    .A(_06370_),
    .X(_06379_));
 sg13g2_xnor2_1 _13690_ (.Y(_06380_),
    .A(\vgadonut.donut.ysA[9] ),
    .B(_06379_));
 sg13g2_nor2_1 _13691_ (.A(_06369_),
    .B(_06380_),
    .Y(_06381_));
 sg13g2_xor2_1 _13692_ (.B(_06380_),
    .A(_06369_),
    .X(_06382_));
 sg13g2_nor3_1 _13693_ (.A(_06364_),
    .B(_06366_),
    .C(_06382_),
    .Y(_06383_));
 sg13g2_o21ai_1 _13694_ (.B1(_06382_),
    .Y(_06384_),
    .A1(_06364_),
    .A2(_06366_));
 sg13g2_a21oi_1 _13695_ (.A1(\vgadonut.donut.donuthit.rzin[2] ),
    .A2(net1904),
    .Y(_06385_),
    .B1(_06348_));
 sg13g2_nor2_1 _13696_ (.A(\vgadonut.donut.donuthit.rzin[3] ),
    .B(\vgadonut.donut.cAsB[9] ),
    .Y(_06386_));
 sg13g2_xnor2_1 _13697_ (.Y(_06387_),
    .A(\vgadonut.donut.donuthit.rzin[3] ),
    .B(net1903));
 sg13g2_xnor2_1 _13698_ (.Y(_06388_),
    .A(_06385_),
    .B(_06387_));
 sg13g2_nand2b_1 _13699_ (.Y(_06389_),
    .B(_06384_),
    .A_N(_06383_));
 sg13g2_a221oi_1 _13700_ (.B2(net1759),
    .C1(net1657),
    .B1(_06389_),
    .A1(net1744),
    .Y(_06390_),
    .A2(_06388_));
 sg13g2_a21o_1 _13701_ (.A2(net1657),
    .A1(net2130),
    .B1(_06390_),
    .X(_00486_));
 sg13g2_nand2_1 _13702_ (.Y(_06391_),
    .A(\vgadonut.donut.donuthit.rzin[4] ),
    .B(\vgadonut.donut.cAsB[10] ));
 sg13g2_nor2_1 _13703_ (.A(\vgadonut.donut.donuthit.rzin[4] ),
    .B(\vgadonut.donut.cAsB[10] ),
    .Y(_06392_));
 sg13g2_xor2_1 _13704_ (.B(net1902),
    .A(\vgadonut.donut.donuthit.rzin[4] ),
    .X(_06393_));
 sg13g2_nor2_1 _13705_ (.A(_06385_),
    .B(_06386_),
    .Y(_06394_));
 sg13g2_a21oi_2 _13706_ (.B1(_06394_),
    .Y(_06395_),
    .A2(net1903),
    .A1(\vgadonut.donut.donuthit.rzin[3] ));
 sg13g2_xnor2_1 _13707_ (.Y(_06396_),
    .A(_06393_),
    .B(_06395_));
 sg13g2_a21oi_1 _13708_ (.A1(net1750),
    .A2(_06396_),
    .Y(_06397_),
    .B1(net1656));
 sg13g2_nor2b_1 _13709_ (.A(_06381_),
    .B_N(_06384_),
    .Y(_06398_));
 sg13g2_a21oi_1 _13710_ (.A1(net1957),
    .A2(_06376_),
    .Y(_06399_),
    .B1(_06375_));
 sg13g2_a21oi_2 _13711_ (.B1(_06372_),
    .Y(_06400_),
    .A2(_06373_),
    .A1(_00097_));
 sg13g2_nor2_1 _13712_ (.A(net1905),
    .B(net1904),
    .Y(_06401_));
 sg13g2_xor2_1 _13713_ (.B(net1904),
    .A(net1905),
    .X(_06402_));
 sg13g2_xnor2_1 _13714_ (.Y(_06403_),
    .A(_00098_),
    .B(_06402_));
 sg13g2_nor2_1 _13715_ (.A(_06400_),
    .B(_06403_),
    .Y(_06404_));
 sg13g2_xor2_1 _13716_ (.B(_06403_),
    .A(_06400_),
    .X(_06405_));
 sg13g2_xnor2_1 _13717_ (.Y(_06406_),
    .A(net1955),
    .B(_06405_));
 sg13g2_or2_1 _13718_ (.X(_06407_),
    .B(_06406_),
    .A(_06399_));
 sg13g2_xor2_1 _13719_ (.B(_06406_),
    .A(_06399_),
    .X(_06408_));
 sg13g2_nand2_1 _13720_ (.Y(_06409_),
    .A(\vgadonut.donut.ysA[10] ),
    .B(_06408_));
 sg13g2_xnor2_1 _13721_ (.Y(_06410_),
    .A(\vgadonut.donut.ysA[10] ),
    .B(_06408_));
 sg13g2_a21oi_1 _13722_ (.A1(\vgadonut.donut.ysA[9] ),
    .A2(_06379_),
    .Y(_06411_),
    .B1(_06378_));
 sg13g2_or2_1 _13723_ (.X(_06412_),
    .B(_06411_),
    .A(_06410_));
 sg13g2_xnor2_1 _13724_ (.Y(_06413_),
    .A(_06410_),
    .B(_06411_));
 sg13g2_a21oi_1 _13725_ (.A1(_06398_),
    .A2(_06413_),
    .Y(_06414_),
    .B1(net1744));
 sg13g2_o21ai_1 _13726_ (.B1(_06414_),
    .Y(_06415_),
    .A1(_06398_),
    .A2(_06413_));
 sg13g2_a22oi_1 _13727_ (.Y(_00487_),
    .B1(_06397_),
    .B2(_06415_),
    .A2(net1656),
    .A1(_06864_));
 sg13g2_o21ai_1 _13728_ (.B1(_06412_),
    .Y(_06416_),
    .A1(_06398_),
    .A2(_06413_));
 sg13g2_a21oi_1 _13729_ (.A1(net1955),
    .A2(_06405_),
    .Y(_06417_),
    .B1(_06404_));
 sg13g2_a21oi_1 _13730_ (.A1(_00098_),
    .A2(_06402_),
    .Y(_06418_),
    .B1(_06401_));
 sg13g2_nor2_1 _13731_ (.A(net1904),
    .B(net1903),
    .Y(_06419_));
 sg13g2_xor2_1 _13732_ (.B(net1903),
    .A(net1904),
    .X(_06420_));
 sg13g2_xnor2_1 _13733_ (.Y(_06421_),
    .A(_00099_),
    .B(_06420_));
 sg13g2_nor2_1 _13734_ (.A(_06418_),
    .B(_06421_),
    .Y(_06422_));
 sg13g2_xor2_1 _13735_ (.B(_06421_),
    .A(_06418_),
    .X(_06423_));
 sg13g2_xnor2_1 _13736_ (.Y(_06424_),
    .A(net1953),
    .B(_06423_));
 sg13g2_nor2_1 _13737_ (.A(_06417_),
    .B(_06424_),
    .Y(_06425_));
 sg13g2_xor2_1 _13738_ (.B(_06424_),
    .A(_06417_),
    .X(_06426_));
 sg13g2_xnor2_1 _13739_ (.Y(_06427_),
    .A(\vgadonut.donut.ysA[11] ),
    .B(_06426_));
 sg13g2_nand3_1 _13740_ (.B(_06409_),
    .C(_06427_),
    .A(_06407_),
    .Y(_06428_));
 sg13g2_a21o_1 _13741_ (.A2(_06409_),
    .A1(_06407_),
    .B1(_06427_),
    .X(_06429_));
 sg13g2_nand2_1 _13742_ (.Y(_06430_),
    .A(_06428_),
    .B(_06429_));
 sg13g2_o21ai_1 _13743_ (.B1(_06391_),
    .Y(_06431_),
    .A1(_06392_),
    .A2(_06395_));
 sg13g2_nor2_1 _13744_ (.A(\vgadonut.donut.donuthit.rzin[5] ),
    .B(net1901),
    .Y(_06432_));
 sg13g2_xnor2_1 _13745_ (.Y(_06433_),
    .A(\vgadonut.donut.donuthit.rzin[5] ),
    .B(net1901));
 sg13g2_xnor2_1 _13746_ (.Y(_06434_),
    .A(_06431_),
    .B(_06433_));
 sg13g2_xnor2_1 _13747_ (.Y(_06435_),
    .A(_06416_),
    .B(_06430_));
 sg13g2_a221oi_1 _13748_ (.B2(net1748),
    .C1(net1655),
    .B1(_06435_),
    .A1(net1751),
    .Y(_06436_),
    .A2(_06434_));
 sg13g2_a21oi_1 _13749_ (.A1(_06867_),
    .A2(net1654),
    .Y(_00488_),
    .B1(_06436_));
 sg13g2_xnor2_1 _13750_ (.Y(_06437_),
    .A(\vgadonut.donut.donuthit.rzin[6] ),
    .B(net1900));
 sg13g2_a21oi_1 _13751_ (.A1(\vgadonut.donut.donuthit.rzin[5] ),
    .A2(net1901),
    .Y(_06438_),
    .B1(_06431_));
 sg13g2_nor3_1 _13752_ (.A(_06432_),
    .B(_06437_),
    .C(_06438_),
    .Y(_06439_));
 sg13g2_o21ai_1 _13753_ (.B1(_06437_),
    .Y(_06440_),
    .A1(_06432_),
    .A2(_06438_));
 sg13g2_nor2b_1 _13754_ (.A(_06439_),
    .B_N(_06440_),
    .Y(_06441_));
 sg13g2_a21oi_1 _13755_ (.A1(net1751),
    .A2(_06441_),
    .Y(_06442_),
    .B1(net1655));
 sg13g2_a21oi_1 _13756_ (.A1(net1953),
    .A2(_06423_),
    .Y(_06443_),
    .B1(_06422_));
 sg13g2_a21oi_1 _13757_ (.A1(_00099_),
    .A2(_06420_),
    .Y(_06444_),
    .B1(_06419_));
 sg13g2_nor2_1 _13758_ (.A(net1903),
    .B(net1902),
    .Y(_06445_));
 sg13g2_xor2_1 _13759_ (.B(net1902),
    .A(net1903),
    .X(_06446_));
 sg13g2_xnor2_1 _13760_ (.Y(_06447_),
    .A(_00100_),
    .B(_06446_));
 sg13g2_nor2_1 _13761_ (.A(_06444_),
    .B(_06447_),
    .Y(_06448_));
 sg13g2_xor2_1 _13762_ (.B(_06447_),
    .A(_06444_),
    .X(_06449_));
 sg13g2_xnor2_1 _13763_ (.Y(_06450_),
    .A(net1951),
    .B(_06449_));
 sg13g2_nor2_1 _13764_ (.A(_06443_),
    .B(_06450_),
    .Y(_06451_));
 sg13g2_xor2_1 _13765_ (.B(_06450_),
    .A(_06443_),
    .X(_06452_));
 sg13g2_xnor2_1 _13766_ (.Y(_06453_),
    .A(\vgadonut.donut.ysA[12] ),
    .B(_06452_));
 sg13g2_a21oi_1 _13767_ (.A1(\vgadonut.donut.ysA[11] ),
    .A2(_06426_),
    .Y(_06454_),
    .B1(_06425_));
 sg13g2_nor2_1 _13768_ (.A(_06453_),
    .B(_06454_),
    .Y(_06455_));
 sg13g2_xnor2_1 _13769_ (.Y(_06456_),
    .A(_06453_),
    .B(_06454_));
 sg13g2_nand2_1 _13770_ (.Y(_06457_),
    .A(_06416_),
    .B(_06428_));
 sg13g2_nand3_1 _13771_ (.B(_06456_),
    .C(_06457_),
    .A(_06429_),
    .Y(_06458_));
 sg13g2_a21oi_1 _13772_ (.A1(_06429_),
    .A2(_06457_),
    .Y(_06459_),
    .B1(_06456_));
 sg13g2_nand3b_1 _13773_ (.B(net1759),
    .C(_06458_),
    .Y(_06460_),
    .A_N(_06459_));
 sg13g2_a22oi_1 _13774_ (.Y(_00489_),
    .B1(_06442_),
    .B2(_06460_),
    .A2(net1655),
    .A1(_06868_));
 sg13g2_a21oi_1 _13775_ (.A1(\vgadonut.donut.ysA[12] ),
    .A2(_06452_),
    .Y(_06461_),
    .B1(_06451_));
 sg13g2_a21oi_1 _13776_ (.A1(net1951),
    .A2(_06449_),
    .Y(_06462_),
    .B1(_06448_));
 sg13g2_a21oi_1 _13777_ (.A1(_00100_),
    .A2(_06446_),
    .Y(_06463_),
    .B1(_06445_));
 sg13g2_nor2_1 _13778_ (.A(net1902),
    .B(\vgadonut.donut.cAsB[11] ),
    .Y(_06464_));
 sg13g2_xor2_1 _13779_ (.B(\vgadonut.donut.cAsB[11] ),
    .A(net1902),
    .X(_06465_));
 sg13g2_xnor2_1 _13780_ (.Y(_06466_),
    .A(_00101_),
    .B(_06465_));
 sg13g2_nor2_1 _13781_ (.A(_06463_),
    .B(_06466_),
    .Y(_06467_));
 sg13g2_xor2_1 _13782_ (.B(_06466_),
    .A(_06463_),
    .X(_06468_));
 sg13g2_xnor2_1 _13783_ (.Y(_06469_),
    .A(net1949),
    .B(_06468_));
 sg13g2_nor2_1 _13784_ (.A(_06462_),
    .B(_06469_),
    .Y(_06470_));
 sg13g2_xor2_1 _13785_ (.B(_06469_),
    .A(_06462_),
    .X(_06471_));
 sg13g2_xnor2_1 _13786_ (.Y(_06472_),
    .A(\vgadonut.donut.ysA[13] ),
    .B(_06471_));
 sg13g2_nor2_1 _13787_ (.A(_06461_),
    .B(_06472_),
    .Y(_06473_));
 sg13g2_xor2_1 _13788_ (.B(_06472_),
    .A(_06461_),
    .X(_06474_));
 sg13g2_nor3_1 _13789_ (.A(_06455_),
    .B(_06459_),
    .C(_06474_),
    .Y(_06475_));
 sg13g2_o21ai_1 _13790_ (.B1(_06474_),
    .Y(_06476_),
    .A1(_06455_),
    .A2(_06459_));
 sg13g2_a21o_1 _13791_ (.A2(net1900),
    .A1(\vgadonut.donut.donuthit.rzin[6] ),
    .B1(_06439_),
    .X(_06477_));
 sg13g2_nand2_1 _13792_ (.Y(_06478_),
    .A(\vgadonut.donut.donuthit.rzin[7] ),
    .B(net1898));
 sg13g2_xor2_1 _13793_ (.B(net1898),
    .A(\vgadonut.donut.donuthit.rzin[7] ),
    .X(_06479_));
 sg13g2_xnor2_1 _13794_ (.Y(_06480_),
    .A(_06477_),
    .B(_06479_));
 sg13g2_nand2b_1 _13795_ (.Y(_06481_),
    .B(_06476_),
    .A_N(_06475_));
 sg13g2_a221oi_1 _13796_ (.B2(net1759),
    .C1(net1655),
    .B1(_06481_),
    .A1(net1744),
    .Y(_06482_),
    .A2(_06480_));
 sg13g2_a21o_1 _13797_ (.A2(net1655),
    .A1(net2232),
    .B1(_06482_),
    .X(_00490_));
 sg13g2_xnor2_1 _13798_ (.Y(_06483_),
    .A(\vgadonut.donut.donuthit.rzin[8] ),
    .B(\vgadonut.donut.cAsB[14] ));
 sg13g2_o21ai_1 _13799_ (.B1(_06477_),
    .Y(_06484_),
    .A1(\vgadonut.donut.donuthit.rzin[7] ),
    .A2(net1898));
 sg13g2_a21oi_1 _13800_ (.A1(_06478_),
    .A2(_06484_),
    .Y(_06485_),
    .B1(_06483_));
 sg13g2_nand3_1 _13801_ (.B(_06483_),
    .C(_06484_),
    .A(_06478_),
    .Y(_06486_));
 sg13g2_nor2b_1 _13802_ (.A(_06485_),
    .B_N(_06486_),
    .Y(_06487_));
 sg13g2_a21oi_1 _13803_ (.A1(net1751),
    .A2(_06487_),
    .Y(_06488_),
    .B1(net1654));
 sg13g2_nor2b_1 _13804_ (.A(_06473_),
    .B_N(_06476_),
    .Y(_06489_));
 sg13g2_a21oi_1 _13805_ (.A1(net1949),
    .A2(_06468_),
    .Y(_06490_),
    .B1(_06467_));
 sg13g2_a21oi_1 _13806_ (.A1(_00101_),
    .A2(_06465_),
    .Y(_06491_),
    .B1(_06464_));
 sg13g2_nor2_1 _13807_ (.A(net1901),
    .B(net1900),
    .Y(_06492_));
 sg13g2_xor2_1 _13808_ (.B(net1900),
    .A(net1901),
    .X(_06493_));
 sg13g2_xnor2_1 _13809_ (.Y(_06494_),
    .A(_00102_),
    .B(_06493_));
 sg13g2_nor2_1 _13810_ (.A(_06491_),
    .B(_06494_),
    .Y(_06495_));
 sg13g2_xor2_1 _13811_ (.B(_06494_),
    .A(_06491_),
    .X(_06496_));
 sg13g2_xnor2_1 _13812_ (.Y(_06497_),
    .A(net1948),
    .B(_06496_));
 sg13g2_nor2_1 _13813_ (.A(_06490_),
    .B(_06497_),
    .Y(_06498_));
 sg13g2_xor2_1 _13814_ (.B(_06497_),
    .A(_06490_),
    .X(_06499_));
 sg13g2_xnor2_1 _13815_ (.Y(_06500_),
    .A(\vgadonut.donut.ysA[14] ),
    .B(_06499_));
 sg13g2_a21oi_1 _13816_ (.A1(\vgadonut.donut.ysA[13] ),
    .A2(_06471_),
    .Y(_06501_),
    .B1(_06470_));
 sg13g2_nor2_1 _13817_ (.A(_06500_),
    .B(_06501_),
    .Y(_06502_));
 sg13g2_xnor2_1 _13818_ (.Y(_06503_),
    .A(_06500_),
    .B(_06501_));
 sg13g2_nor2_1 _13819_ (.A(_06489_),
    .B(_06503_),
    .Y(_06504_));
 sg13g2_a21oi_1 _13820_ (.A1(_06489_),
    .A2(_06503_),
    .Y(_06505_),
    .B1(net1744));
 sg13g2_nand2b_1 _13821_ (.Y(_06506_),
    .B(_06505_),
    .A_N(_06504_));
 sg13g2_a22oi_1 _13822_ (.Y(_00491_),
    .B1(_06488_),
    .B2(_06506_),
    .A2(net1654),
    .A1(_06872_));
 sg13g2_a21oi_1 _13823_ (.A1(\vgadonut.donut.ysA[14] ),
    .A2(_06499_),
    .Y(_06507_),
    .B1(_06498_));
 sg13g2_a21oi_1 _13824_ (.A1(net1948),
    .A2(_06496_),
    .Y(_06508_),
    .B1(_06495_));
 sg13g2_a21oi_1 _13825_ (.A1(_00102_),
    .A2(_06493_),
    .Y(_06509_),
    .B1(_06492_));
 sg13g2_nor2_1 _13826_ (.A(\vgadonut.donut.cAsB[12] ),
    .B(net1898),
    .Y(_06510_));
 sg13g2_xor2_1 _13827_ (.B(net1898),
    .A(\vgadonut.donut.cAsB[12] ),
    .X(_06511_));
 sg13g2_xnor2_1 _13828_ (.Y(_06512_),
    .A(_00103_),
    .B(_06511_));
 sg13g2_nor2_1 _13829_ (.A(_06509_),
    .B(_06512_),
    .Y(_06513_));
 sg13g2_xor2_1 _13830_ (.B(_06512_),
    .A(_06509_),
    .X(_06514_));
 sg13g2_xnor2_1 _13831_ (.Y(_06515_),
    .A(net1946),
    .B(_06514_));
 sg13g2_nor2_1 _13832_ (.A(_06508_),
    .B(_06515_),
    .Y(_06516_));
 sg13g2_xor2_1 _13833_ (.B(_06515_),
    .A(_06508_),
    .X(_06517_));
 sg13g2_xnor2_1 _13834_ (.Y(_06518_),
    .A(\vgadonut.donut.ysA[15] ),
    .B(_06517_));
 sg13g2_nor2_1 _13835_ (.A(_06507_),
    .B(_06518_),
    .Y(_06519_));
 sg13g2_xor2_1 _13836_ (.B(_06518_),
    .A(_06507_),
    .X(_06520_));
 sg13g2_o21ai_1 _13837_ (.B1(_06520_),
    .Y(_06521_),
    .A1(_06502_),
    .A2(_06504_));
 sg13g2_or3_1 _13838_ (.A(_06502_),
    .B(_06504_),
    .C(_06520_),
    .X(_06522_));
 sg13g2_a21oi_1 _13839_ (.A1(\vgadonut.donut.donuthit.rzin[8] ),
    .A2(net1897),
    .Y(_06523_),
    .B1(_06485_));
 sg13g2_or2_1 _13840_ (.X(_06524_),
    .B(net1894),
    .A(\vgadonut.donut.donuthit.rzin[9] ));
 sg13g2_nand2_1 _13841_ (.Y(_06525_),
    .A(\vgadonut.donut.donuthit.rzin[9] ),
    .B(net1896));
 sg13g2_nand2_1 _13842_ (.Y(_06526_),
    .A(_06524_),
    .B(_06525_));
 sg13g2_xnor2_1 _13843_ (.Y(_06527_),
    .A(_06523_),
    .B(_06526_));
 sg13g2_nand2_1 _13844_ (.Y(_06528_),
    .A(_06521_),
    .B(_06522_));
 sg13g2_a221oi_1 _13845_ (.B2(net1757),
    .C1(net1655),
    .B1(_06528_),
    .A1(net1744),
    .Y(_06529_),
    .A2(_06527_));
 sg13g2_a21o_1 _13846_ (.A2(net1655),
    .A1(net2171),
    .B1(_06529_),
    .X(_00492_));
 sg13g2_nand2_1 _13847_ (.Y(_06530_),
    .A(_06875_),
    .B(_06876_));
 sg13g2_nand2_1 _13848_ (.Y(_06531_),
    .A(net1894),
    .B(\vgadonut.donut.donuthit.rzin[10] ));
 sg13g2_nand2_1 _13849_ (.Y(_06532_),
    .A(_06523_),
    .B(_06525_));
 sg13g2_and4_1 _13850_ (.A(_06524_),
    .B(_06530_),
    .C(_06531_),
    .D(_06532_),
    .X(_06533_));
 sg13g2_a22oi_1 _13851_ (.Y(_06534_),
    .B1(_06532_),
    .B2(_06524_),
    .A2(_06531_),
    .A1(_06530_));
 sg13g2_nor3_1 _13852_ (.A(net1748),
    .B(_06533_),
    .C(_06534_),
    .Y(_06535_));
 sg13g2_nor2_1 _13853_ (.A(net1656),
    .B(_06535_),
    .Y(_06536_));
 sg13g2_nor2b_1 _13854_ (.A(_06519_),
    .B_N(_06521_),
    .Y(_06537_));
 sg13g2_a21oi_1 _13855_ (.A1(net1946),
    .A2(_06514_),
    .Y(_06538_),
    .B1(_06513_));
 sg13g2_a21oi_1 _13856_ (.A1(_00103_),
    .A2(_06511_),
    .Y(_06539_),
    .B1(_06510_));
 sg13g2_nor2_1 _13857_ (.A(net1898),
    .B(net1897),
    .Y(_06540_));
 sg13g2_xor2_1 _13858_ (.B(net1897),
    .A(net1898),
    .X(_06541_));
 sg13g2_xnor2_1 _13859_ (.Y(_06542_),
    .A(_00104_),
    .B(_06541_));
 sg13g2_nor2_1 _13860_ (.A(_06539_),
    .B(_06542_),
    .Y(_06543_));
 sg13g2_xor2_1 _13861_ (.B(_06542_),
    .A(_06539_),
    .X(_06544_));
 sg13g2_xnor2_1 _13862_ (.Y(_06545_),
    .A(net1944),
    .B(_06544_));
 sg13g2_or2_1 _13863_ (.X(_06546_),
    .B(_06545_),
    .A(_06538_));
 sg13g2_xor2_1 _13864_ (.B(_06545_),
    .A(_06538_),
    .X(_06547_));
 sg13g2_nand2_1 _13865_ (.Y(_06548_),
    .A(\vgadonut.donut.ysA[16] ),
    .B(_06547_));
 sg13g2_xnor2_1 _13866_ (.Y(_06549_),
    .A(\vgadonut.donut.ysA[16] ),
    .B(_06547_));
 sg13g2_a21oi_1 _13867_ (.A1(\vgadonut.donut.ysA[15] ),
    .A2(_06517_),
    .Y(_06550_),
    .B1(_06516_));
 sg13g2_nor2_1 _13868_ (.A(_06549_),
    .B(_06550_),
    .Y(_06551_));
 sg13g2_xnor2_1 _13869_ (.Y(_06552_),
    .A(_06549_),
    .B(_06550_));
 sg13g2_nor2_1 _13870_ (.A(_06537_),
    .B(_06552_),
    .Y(_06553_));
 sg13g2_a21oi_1 _13871_ (.A1(_06537_),
    .A2(_06552_),
    .Y(_06554_),
    .B1(net1747));
 sg13g2_nand2b_1 _13872_ (.Y(_06555_),
    .B(_06554_),
    .A_N(_06553_));
 sg13g2_a22oi_1 _13873_ (.Y(_00493_),
    .B1(_06536_),
    .B2(_06555_),
    .A2(net1654),
    .A1(_06876_));
 sg13g2_nor2_1 _13874_ (.A(net2164),
    .B(_03934_),
    .Y(_06556_));
 sg13g2_nor2_1 _13875_ (.A(_06551_),
    .B(_06553_),
    .Y(_06557_));
 sg13g2_a21oi_2 _13876_ (.B1(_06543_),
    .Y(_06558_),
    .A2(_06544_),
    .A1(net1944));
 sg13g2_a21oi_1 _13877_ (.A1(_00104_),
    .A2(_06541_),
    .Y(_06559_),
    .B1(_06540_));
 sg13g2_nor2_1 _13878_ (.A(net1897),
    .B(net1894),
    .Y(_06560_));
 sg13g2_xor2_1 _13879_ (.B(net1894),
    .A(net1897),
    .X(_06561_));
 sg13g2_xnor2_1 _13880_ (.Y(_06562_),
    .A(_00105_),
    .B(_06561_));
 sg13g2_nor2_1 _13881_ (.A(_06559_),
    .B(_06562_),
    .Y(_06563_));
 sg13g2_xor2_1 _13882_ (.B(_06562_),
    .A(_06559_),
    .X(_06564_));
 sg13g2_xnor2_1 _13883_ (.Y(_06565_),
    .A(net1942),
    .B(_06564_));
 sg13g2_nor2_1 _13884_ (.A(_06558_),
    .B(_06565_),
    .Y(_06566_));
 sg13g2_xor2_1 _13885_ (.B(_06565_),
    .A(_06558_),
    .X(_06567_));
 sg13g2_xnor2_1 _13886_ (.Y(_06568_),
    .A(\vgadonut.donut.ysA[17] ),
    .B(_06567_));
 sg13g2_nand3_1 _13887_ (.B(_06548_),
    .C(_06568_),
    .A(_06546_),
    .Y(_06569_));
 sg13g2_a21o_1 _13888_ (.A2(_06548_),
    .A1(_06546_),
    .B1(_06568_),
    .X(_06570_));
 sg13g2_nand2_1 _13889_ (.Y(_06571_),
    .A(_06569_),
    .B(_06570_));
 sg13g2_xor2_1 _13890_ (.B(\vgadonut.donut.donuthit.rzin[11] ),
    .A(net1895),
    .X(_06572_));
 sg13g2_a21oi_1 _13891_ (.A1(net1895),
    .A2(\vgadonut.donut.donuthit.rzin[10] ),
    .Y(_06573_),
    .B1(_06533_));
 sg13g2_xnor2_1 _13892_ (.Y(_06574_),
    .A(_06572_),
    .B(_06573_));
 sg13g2_xor2_1 _13893_ (.B(_06571_),
    .A(_06557_),
    .X(_06575_));
 sg13g2_a22oi_1 _13894_ (.Y(_06576_),
    .B1(_06575_),
    .B2(net1748),
    .A2(_06574_),
    .A1(net1751));
 sg13g2_a21oi_1 _13895_ (.A1(_03934_),
    .A2(_06576_),
    .Y(_00494_),
    .B1(_06556_));
 sg13g2_nor2_1 _13896_ (.A(_06875_),
    .B(_06878_),
    .Y(_06577_));
 sg13g2_xor2_1 _13897_ (.B(\vgadonut.donut.donuthit.rzin[12] ),
    .A(net1896),
    .X(_06578_));
 sg13g2_nand2_1 _13898_ (.Y(_06579_),
    .A(_06533_),
    .B(_06572_));
 sg13g2_o21ai_1 _13899_ (.B1(net1895),
    .Y(_06580_),
    .A1(\vgadonut.donut.donuthit.rzin[10] ),
    .A2(\vgadonut.donut.donuthit.rzin[11] ));
 sg13g2_nand2_1 _13900_ (.Y(_06581_),
    .A(_06579_),
    .B(_06580_));
 sg13g2_xor2_1 _13901_ (.B(_06581_),
    .A(_06578_),
    .X(_06582_));
 sg13g2_a21oi_1 _13902_ (.A1(net1750),
    .A2(_06582_),
    .Y(_06583_),
    .B1(net1654));
 sg13g2_a21oi_1 _13903_ (.A1(net1942),
    .A2(_06564_),
    .Y(_06584_),
    .B1(_06563_));
 sg13g2_a21oi_1 _13904_ (.A1(_00105_),
    .A2(_06561_),
    .Y(_06585_),
    .B1(_06560_));
 sg13g2_nor2_1 _13905_ (.A(\vgadonut.donut.cAsB[12] ),
    .B(_06585_),
    .Y(_06586_));
 sg13g2_xor2_1 _13906_ (.B(_06585_),
    .A(net1900),
    .X(_06587_));
 sg13g2_xnor2_1 _13907_ (.Y(_06588_),
    .A(net1940),
    .B(_06587_));
 sg13g2_or2_1 _13908_ (.X(_06589_),
    .B(_06588_),
    .A(_06584_));
 sg13g2_xor2_1 _13909_ (.B(_06588_),
    .A(_06584_),
    .X(_06590_));
 sg13g2_nand2_1 _13910_ (.Y(_06591_),
    .A(\vgadonut.donut.ysA[18] ),
    .B(_06590_));
 sg13g2_xnor2_1 _13911_ (.Y(_06592_),
    .A(\vgadonut.donut.ysA[18] ),
    .B(_06590_));
 sg13g2_a21oi_1 _13912_ (.A1(\vgadonut.donut.ysA[17] ),
    .A2(_06567_),
    .Y(_06593_),
    .B1(_06566_));
 sg13g2_nor2_1 _13913_ (.A(_06592_),
    .B(_06593_),
    .Y(_06594_));
 sg13g2_xnor2_1 _13914_ (.Y(_06595_),
    .A(_06592_),
    .B(_06593_));
 sg13g2_o21ai_1 _13915_ (.B1(_06569_),
    .Y(_06596_),
    .A1(_06551_),
    .A2(_06553_));
 sg13g2_nand3_1 _13916_ (.B(_06595_),
    .C(_06596_),
    .A(_06570_),
    .Y(_06597_));
 sg13g2_a21oi_1 _13917_ (.A1(_06570_),
    .A2(_06596_),
    .Y(_06598_),
    .B1(_06595_));
 sg13g2_nand3b_1 _13918_ (.B(net1757),
    .C(_06597_),
    .Y(_06599_),
    .A_N(_06598_));
 sg13g2_a22oi_1 _13919_ (.Y(_00495_),
    .B1(_06583_),
    .B2(_06599_),
    .A2(net1654),
    .A1(_06878_));
 sg13g2_nor2_1 _13920_ (.A(net2189),
    .B(_03934_),
    .Y(_06600_));
 sg13g2_nor2_1 _13921_ (.A(_06594_),
    .B(_06598_),
    .Y(_06601_));
 sg13g2_a21oi_1 _13922_ (.A1(net1940),
    .A2(_06587_),
    .Y(_06602_),
    .B1(_06586_));
 sg13g2_nor2_1 _13923_ (.A(net1899),
    .B(net1894),
    .Y(_06603_));
 sg13g2_xor2_1 _13924_ (.B(net1894),
    .A(net1898),
    .X(_06604_));
 sg13g2_xnor2_1 _13925_ (.Y(_06605_),
    .A(net1938),
    .B(_06604_));
 sg13g2_nor2_1 _13926_ (.A(_06602_),
    .B(_06605_),
    .Y(_06606_));
 sg13g2_xor2_1 _13927_ (.B(_06605_),
    .A(_06602_),
    .X(_06607_));
 sg13g2_xnor2_1 _13928_ (.Y(_06608_),
    .A(\vgadonut.donut.ysA[19] ),
    .B(_06607_));
 sg13g2_nand3_1 _13929_ (.B(_06591_),
    .C(_06608_),
    .A(_06589_),
    .Y(_06609_));
 sg13g2_a21o_1 _13930_ (.A2(_06591_),
    .A1(_06589_),
    .B1(_06608_),
    .X(_06610_));
 sg13g2_nand2_1 _13931_ (.Y(_06611_),
    .A(_06609_),
    .B(_06610_));
 sg13g2_xnor2_1 _13932_ (.Y(_06612_),
    .A(net1895),
    .B(\vgadonut.donut.donuthit.rzin[13] ));
 sg13g2_a21oi_1 _13933_ (.A1(_06578_),
    .A2(_06581_),
    .Y(_06613_),
    .B1(_06577_));
 sg13g2_xor2_1 _13934_ (.B(_06613_),
    .A(_06612_),
    .X(_06614_));
 sg13g2_xor2_1 _13935_ (.B(_06611_),
    .A(_06601_),
    .X(_06615_));
 sg13g2_a22oi_1 _13936_ (.Y(_06616_),
    .B1(_06615_),
    .B2(net1748),
    .A2(_06614_),
    .A1(net1750));
 sg13g2_a21oi_1 _13937_ (.A1(net1670),
    .A2(_06616_),
    .Y(_00496_),
    .B1(_06600_));
 sg13g2_xor2_1 _13938_ (.B(\vgadonut.donut.donuthit.rzin[14] ),
    .A(net1895),
    .X(_06617_));
 sg13g2_nor2_1 _13939_ (.A(_06579_),
    .B(_06612_),
    .Y(_06618_));
 sg13g2_o21ai_1 _13940_ (.B1(net1895),
    .Y(_06619_),
    .A1(\vgadonut.donut.donuthit.rzin[12] ),
    .A2(\vgadonut.donut.donuthit.rzin[13] ));
 sg13g2_nand2_1 _13941_ (.Y(_06620_),
    .A(_06580_),
    .B(_06619_));
 sg13g2_a21oi_1 _13942_ (.A1(_06578_),
    .A2(_06618_),
    .Y(_06621_),
    .B1(_06620_));
 sg13g2_nand2b_1 _13943_ (.Y(_06622_),
    .B(_06617_),
    .A_N(_06621_));
 sg13g2_xnor2_1 _13944_ (.Y(_06623_),
    .A(_06617_),
    .B(_06621_));
 sg13g2_a21oi_1 _13945_ (.A1(net1750),
    .A2(_06623_),
    .Y(_06624_),
    .B1(net1654));
 sg13g2_a21oi_1 _13946_ (.A1(net1938),
    .A2(_06604_),
    .Y(_06625_),
    .B1(_06603_));
 sg13g2_xnor2_1 _13947_ (.Y(_06626_),
    .A(net1936),
    .B(_06561_));
 sg13g2_nor2_1 _13948_ (.A(_06625_),
    .B(_06626_),
    .Y(_06627_));
 sg13g2_xor2_1 _13949_ (.B(_06626_),
    .A(_06625_),
    .X(_06628_));
 sg13g2_xnor2_1 _13950_ (.Y(_06629_),
    .A(\vgadonut.donut.ysA[20] ),
    .B(_06628_));
 sg13g2_a21oi_1 _13951_ (.A1(\vgadonut.donut.ysA[19] ),
    .A2(_06607_),
    .Y(_06630_),
    .B1(_06606_));
 sg13g2_nor2_1 _13952_ (.A(_06629_),
    .B(_06630_),
    .Y(_06631_));
 sg13g2_xnor2_1 _13953_ (.Y(_06632_),
    .A(_06629_),
    .B(_06630_));
 sg13g2_o21ai_1 _13954_ (.B1(_06609_),
    .Y(_06633_),
    .A1(_06594_),
    .A2(_06598_));
 sg13g2_nand3_1 _13955_ (.B(_06632_),
    .C(_06633_),
    .A(_06610_),
    .Y(_06634_));
 sg13g2_a21oi_1 _13956_ (.A1(_06610_),
    .A2(_06633_),
    .Y(_06635_),
    .B1(_06632_));
 sg13g2_nand3b_1 _13957_ (.B(net1757),
    .C(_06634_),
    .Y(_06636_),
    .A_N(_06635_));
 sg13g2_a22oi_1 _13958_ (.Y(_00497_),
    .B1(_06624_),
    .B2(_06636_),
    .A2(net1654),
    .A1(_06881_));
 sg13g2_o21ai_1 _13959_ (.B1(_06622_),
    .Y(_06637_),
    .A1(_06875_),
    .A2(_06881_));
 sg13g2_xnor2_1 _13960_ (.Y(_06638_),
    .A(net1895),
    .B(\vgadonut.donut.donuthit.rzin[15] ));
 sg13g2_xnor2_1 _13961_ (.Y(_06639_),
    .A(_06637_),
    .B(_06638_));
 sg13g2_a21oi_1 _13962_ (.A1(net1756),
    .A2(_06639_),
    .Y(_06640_),
    .B1(net1668));
 sg13g2_nor2_1 _13963_ (.A(_06631_),
    .B(_06635_),
    .Y(_06641_));
 sg13g2_a21oi_1 _13964_ (.A1(\vgadonut.donut.ysA[20] ),
    .A2(_06628_),
    .Y(_06642_),
    .B1(_06627_));
 sg13g2_a21oi_1 _13965_ (.A1(net1936),
    .A2(_06561_),
    .Y(_06643_),
    .B1(_06560_));
 sg13g2_xnor2_1 _13966_ (.Y(_06644_),
    .A(net1935),
    .B(\vgadonut.donut.ysA[21] ));
 sg13g2_xnor2_1 _13967_ (.Y(_06645_),
    .A(_06643_),
    .B(_06644_));
 sg13g2_xnor2_1 _13968_ (.Y(_06646_),
    .A(_06642_),
    .B(_06645_));
 sg13g2_a21oi_1 _13969_ (.A1(_06641_),
    .A2(_06646_),
    .Y(_06647_),
    .B1(net1744));
 sg13g2_o21ai_1 _13970_ (.B1(_06647_),
    .Y(_06648_),
    .A1(_06641_),
    .A2(_06646_));
 sg13g2_a22oi_1 _13971_ (.Y(_00498_),
    .B1(_06640_),
    .B2(_06648_),
    .A2(net1668),
    .A1(_06882_));
 sg13g2_nor2_1 _13972_ (.A(net2156),
    .B(net1691),
    .Y(_06649_));
 sg13g2_a21oi_1 _13973_ (.A1(_00574_),
    .A2(net1694),
    .Y(_00499_),
    .B1(_06649_));
 sg13g2_nor2_1 _13974_ (.A(\vgadonut.donut.donuthit.rx[6] ),
    .B(net1691),
    .Y(_06650_));
 sg13g2_a21oi_1 _13975_ (.A1(_00575_),
    .A2(net1691),
    .Y(_00500_),
    .B1(_06650_));
 sg13g2_nor2_1 _13976_ (.A(net2110),
    .B(net1690),
    .Y(_06651_));
 sg13g2_a21oi_1 _13977_ (.A1(_00578_),
    .A2(net1690),
    .Y(_00501_),
    .B1(_06651_));
 sg13g2_nor2_1 _13978_ (.A(net2071),
    .B(net1690),
    .Y(_06652_));
 sg13g2_a21oi_1 _13979_ (.A1(_00580_),
    .A2(net1690),
    .Y(_00502_),
    .B1(_06652_));
 sg13g2_nor2_1 _13980_ (.A(net2092),
    .B(net1690),
    .Y(_06653_));
 sg13g2_a21oi_1 _13981_ (.A1(_00581_),
    .A2(net1690),
    .Y(_00503_),
    .B1(_06653_));
 sg13g2_nor2_1 _13982_ (.A(net2122),
    .B(net1694),
    .Y(_06654_));
 sg13g2_a21oi_1 _13983_ (.A1(_00584_),
    .A2(net1694),
    .Y(_00504_),
    .B1(_06654_));
 sg13g2_nor2_1 _13984_ (.A(net2120),
    .B(net1694),
    .Y(_06655_));
 sg13g2_a21oi_1 _13985_ (.A1(_00586_),
    .A2(net1694),
    .Y(_00505_),
    .B1(_06655_));
 sg13g2_nor2_1 _13986_ (.A(net2198),
    .B(net1696),
    .Y(_06656_));
 sg13g2_a21oi_1 _13987_ (.A1(_00588_),
    .A2(net1697),
    .Y(_00506_),
    .B1(_06656_));
 sg13g2_nor2_1 _13988_ (.A(\vgadonut.donut.donuthit.rx[13] ),
    .B(net1696),
    .Y(_06657_));
 sg13g2_a21oi_1 _13989_ (.A1(_00590_),
    .A2(net1696),
    .Y(_00507_),
    .B1(_06657_));
 sg13g2_nor2_1 _13990_ (.A(net2203),
    .B(net1696),
    .Y(_06658_));
 sg13g2_a21oi_1 _13991_ (.A1(_00591_),
    .A2(net1696),
    .Y(_00508_),
    .B1(_06658_));
 sg13g2_nor2_1 _13992_ (.A(net2144),
    .B(net1696),
    .Y(_06659_));
 sg13g2_a21oi_1 _13993_ (.A1(_00593_),
    .A2(net1696),
    .Y(_00509_),
    .B1(_06659_));
 sg13g2_nor2_1 _13994_ (.A(net2162),
    .B(net1685),
    .Y(_06660_));
 sg13g2_a21oi_1 _13995_ (.A1(_06906_),
    .A2(net1685),
    .Y(_00510_),
    .B1(_06660_));
 sg13g2_nor2_1 _13996_ (.A(\vgadonut.donut.donuthit.ry[6] ),
    .B(net1681),
    .Y(_06661_));
 sg13g2_a21oi_1 _13997_ (.A1(_06907_),
    .A2(net1681),
    .Y(_00511_),
    .B1(_06661_));
 sg13g2_mux2_1 _13998_ (.A0(\vgadonut.donut.donuthit.ryin[7] ),
    .A1(net2134),
    .S(net1675),
    .X(_00512_));
 sg13g2_nor2_1 _13999_ (.A(net2051),
    .B(net1683),
    .Y(_06662_));
 sg13g2_a21oi_1 _14000_ (.A1(_06912_),
    .A2(net1683),
    .Y(_00513_),
    .B1(_06662_));
 sg13g2_nor2_1 _14001_ (.A(net2087),
    .B(net1685),
    .Y(_06663_));
 sg13g2_a21oi_1 _14002_ (.A1(_00547_),
    .A2(net1685),
    .Y(_00514_),
    .B1(_06663_));
 sg13g2_nor2_1 _14003_ (.A(net2049),
    .B(net1683),
    .Y(_06664_));
 sg13g2_a21oi_1 _14004_ (.A1(_00549_),
    .A2(net1683),
    .Y(_00515_),
    .B1(_06664_));
 sg13g2_nor2_1 _14005_ (.A(net2056),
    .B(net1682),
    .Y(_06665_));
 sg13g2_a21oi_1 _14006_ (.A1(_00550_),
    .A2(net1682),
    .Y(_00516_),
    .B1(_06665_));
 sg13g2_nor2_1 _14007_ (.A(\vgadonut.donut.donuthit.ry[12] ),
    .B(net1681),
    .Y(_06666_));
 sg13g2_a21oi_1 _14008_ (.A1(_00551_),
    .A2(net1681),
    .Y(_00517_),
    .B1(_06666_));
 sg13g2_nor2_1 _14009_ (.A(net2035),
    .B(net1681),
    .Y(_06667_));
 sg13g2_a21oi_1 _14010_ (.A1(_00552_),
    .A2(net1681),
    .Y(_00518_),
    .B1(_06667_));
 sg13g2_nor2_1 _14011_ (.A(net2128),
    .B(net1683),
    .Y(_06668_));
 sg13g2_a21oi_1 _14012_ (.A1(_00555_),
    .A2(net1683),
    .Y(_00519_),
    .B1(_06668_));
 sg13g2_nor2_1 _14013_ (.A(net2116),
    .B(net1693),
    .Y(_06669_));
 sg13g2_a21oi_1 _14014_ (.A1(_00559_),
    .A2(net1693),
    .Y(_00520_),
    .B1(_06669_));
 sg13g2_nor2_1 _14015_ (.A(net2100),
    .B(net1689),
    .Y(_06670_));
 sg13g2_a21oi_1 _14016_ (.A1(_06867_),
    .A2(net1689),
    .Y(_00521_),
    .B1(_06670_));
 sg13g2_nor2_1 _14017_ (.A(net2014),
    .B(net1684),
    .Y(_06671_));
 sg13g2_a21oi_1 _14018_ (.A1(_06868_),
    .A2(net1684),
    .Y(_00522_),
    .B1(_06671_));
 sg13g2_mux2_1 _14019_ (.A0(\vgadonut.donut.donuthit.rzin[7] ),
    .A1(net2114),
    .S(net1675),
    .X(_00523_));
 sg13g2_nor2_1 _14020_ (.A(net2067),
    .B(net1688),
    .Y(_06672_));
 sg13g2_a21oi_1 _14021_ (.A1(_06872_),
    .A2(net1688),
    .Y(_00524_),
    .B1(_06672_));
 sg13g2_mux2_1 _14022_ (.A0(\vgadonut.donut.donuthit.rzin[9] ),
    .A1(net2046),
    .S(net1674),
    .X(_00525_));
 sg13g2_nor2_1 _14023_ (.A(net2054),
    .B(net1686),
    .Y(_06673_));
 sg13g2_a21oi_1 _14024_ (.A1(_06876_),
    .A2(net1686),
    .Y(_00526_),
    .B1(_06673_));
 sg13g2_mux2_1 _14025_ (.A0(\vgadonut.donut.donuthit.rzin[11] ),
    .A1(net2131),
    .S(net1674),
    .X(_00527_));
 sg13g2_nor2_1 _14026_ (.A(net2023),
    .B(net1687),
    .Y(_06674_));
 sg13g2_a21oi_1 _14027_ (.A1(_06878_),
    .A2(net1686),
    .Y(_00528_),
    .B1(_06674_));
 sg13g2_mux2_1 _14028_ (.A0(\vgadonut.donut.donuthit.rzin[13] ),
    .A1(net2138),
    .S(net1674),
    .X(_00529_));
 sg13g2_nor2_1 _14029_ (.A(net2074),
    .B(net1686),
    .Y(_06675_));
 sg13g2_a21oi_1 _14030_ (.A1(_06881_),
    .A2(net1686),
    .Y(_00530_),
    .B1(_06675_));
 sg13g2_nand2_1 _14031_ (.Y(_06676_),
    .A(net2029),
    .B(net1674));
 sg13g2_o21ai_1 _14032_ (.B1(_06676_),
    .Y(_00531_),
    .A1(_06882_),
    .A2(net1673));
 sg13g2_xnor2_1 _14033_ (.Y(_06677_),
    .A(net1799),
    .B(\vgadonut.donut.h_count[0] ));
 sg13g2_nor2_2 _14034_ (.A(_00645_),
    .B(_00030_),
    .Y(_06678_));
 sg13g2_nor2_1 _14035_ (.A(_06677_),
    .B(_06678_),
    .Y(_06679_));
 sg13g2_nand2_1 _14036_ (.Y(_06680_),
    .A(\vgadonut.donut.h_count[5] ),
    .B(\vgadonut.frame[5] ));
 sg13g2_or2_1 _14037_ (.X(_06681_),
    .B(\vgadonut.frame[3] ),
    .A(\vgadonut.donut.h_count[3] ));
 sg13g2_a22oi_1 _14038_ (.Y(_06682_),
    .B1(\vgadonut.frame[1] ),
    .B2(net1802),
    .A2(net1803),
    .A1(net1799));
 sg13g2_or2_1 _14039_ (.X(_06683_),
    .B(\vgadonut.frame[2] ),
    .A(net1801));
 sg13g2_o21ai_1 _14040_ (.B1(_06683_),
    .Y(_06684_),
    .A1(net1802),
    .A2(\vgadonut.frame[1] ));
 sg13g2_a22oi_1 _14041_ (.Y(_06685_),
    .B1(\vgadonut.frame[2] ),
    .B2(net1801),
    .A2(\vgadonut.frame[3] ),
    .A1(\vgadonut.donut.h_count[3] ));
 sg13g2_o21ai_1 _14042_ (.B1(_06685_),
    .Y(_06686_),
    .A1(_06682_),
    .A2(_06684_));
 sg13g2_a22oi_1 _14043_ (.Y(_06687_),
    .B1(_06681_),
    .B2(_06686_),
    .A2(\vgadonut.frame[4] ),
    .A1(\vgadonut.donut.h_count[4] ));
 sg13g2_or2_1 _14044_ (.X(_06688_),
    .B(\vgadonut.frame[5] ),
    .A(\vgadonut.donut.h_count[5] ));
 sg13g2_o21ai_1 _14045_ (.B1(_06688_),
    .Y(_06689_),
    .A1(\vgadonut.donut.h_count[4] ),
    .A2(\vgadonut.frame[4] ));
 sg13g2_o21ai_1 _14046_ (.B1(_06680_),
    .Y(_06690_),
    .A1(_06687_),
    .A2(_06689_));
 sg13g2_nor2_1 _14047_ (.A(\vgadonut.bayer_j[1] ),
    .B(\vgadonut.frame[3] ),
    .Y(_06691_));
 sg13g2_nand2_1 _14048_ (.Y(_06692_),
    .A(net1915),
    .B(\vgadonut.frame[2] ));
 sg13g2_nand2_1 _14049_ (.Y(_06693_),
    .A(net1913),
    .B(\vgadonut.frame[5] ));
 sg13g2_a22oi_1 _14050_ (.Y(_06694_),
    .B1(\vgadonut.frame[3] ),
    .B2(\vgadonut.bayer_j[1] ),
    .A2(\vgadonut.frame[4] ),
    .A1(net1914));
 sg13g2_o21ai_1 _14051_ (.B1(_06694_),
    .Y(_06695_),
    .A1(_06691_),
    .A2(_06692_));
 sg13g2_o21ai_1 _14052_ (.B1(_06695_),
    .Y(_06696_),
    .A1(\vgadonut.donut.v_count[2] ),
    .A2(\vgadonut.frame[4] ));
 sg13g2_nor2_1 _14053_ (.A(net1913),
    .B(\vgadonut.frame[5] ),
    .Y(_06697_));
 sg13g2_a221oi_1 _14054_ (.B2(_06696_),
    .C1(_06697_),
    .B1(_06693_),
    .A1(_06849_),
    .Y(_06698_),
    .A2(_00646_));
 sg13g2_a21oi_1 _14055_ (.A1(\vgadonut.donut.v_count[4] ),
    .A2(\vgadonut.frame[6] ),
    .Y(_06699_),
    .B1(_06698_));
 sg13g2_xor2_1 _14056_ (.B(\vgadonut.frame[7] ),
    .A(\vgadonut.frame[6] ),
    .X(_06700_));
 sg13g2_xor2_1 _14057_ (.B(\vgadonut.donut.v_count[5] ),
    .A(\vgadonut.donut.h_count[6] ),
    .X(_06701_));
 sg13g2_xnor2_1 _14058_ (.Y(_06702_),
    .A(_06700_),
    .B(_06701_));
 sg13g2_xnor2_1 _14059_ (.Y(_06703_),
    .A(_06699_),
    .B(_06702_));
 sg13g2_o21ai_1 _14060_ (.B1(_00645_),
    .Y(_06704_),
    .A1(_06690_),
    .A2(_06703_));
 sg13g2_a21oi_1 _14061_ (.A1(_06690_),
    .A2(_06703_),
    .Y(_06705_),
    .B1(_06704_));
 sg13g2_a21oi_2 _14062_ (.B1(net1641),
    .Y(_06706_),
    .A2(_00170_),
    .A1(net1855));
 sg13g2_inv_1 _14063_ (.Y(_06707_),
    .A(_06706_));
 sg13g2_xor2_1 _14064_ (.B(_06678_),
    .A(_06677_),
    .X(_06708_));
 sg13g2_a21oi_1 _14065_ (.A1(_06706_),
    .A2(_06708_),
    .Y(_06709_),
    .B1(_06679_));
 sg13g2_nor2_2 _14066_ (.A(net2344),
    .B(_00645_),
    .Y(_06710_));
 sg13g2_xor2_1 _14067_ (.B(_00655_),
    .A(net1803),
    .X(_06711_));
 sg13g2_xnor2_1 _14068_ (.Y(_06712_),
    .A(net1803),
    .B(_00655_));
 sg13g2_nand2_1 _14069_ (.Y(_06713_),
    .A(_06706_),
    .B(_06712_));
 sg13g2_xnor2_1 _14070_ (.Y(_06714_),
    .A(_06706_),
    .B(_06712_));
 sg13g2_xnor2_1 _14071_ (.Y(_06715_),
    .A(_06710_),
    .B(_06714_));
 sg13g2_or2_1 _14072_ (.X(_06716_),
    .B(_06715_),
    .A(_06709_));
 sg13g2_a21oi_2 _14073_ (.B1(net1640),
    .Y(_06717_),
    .A2(_00171_),
    .A1(net1855));
 sg13g2_inv_1 _14074_ (.Y(_06718_),
    .A(_06717_));
 sg13g2_xnor2_1 _14075_ (.Y(_06719_),
    .A(_00659_),
    .B(_06717_));
 sg13g2_nand2b_1 _14076_ (.Y(_06720_),
    .B(_06719_),
    .A_N(_06678_));
 sg13g2_o21ai_1 _14077_ (.B1(_06720_),
    .Y(_06721_),
    .A1(_00659_),
    .A2(_06718_));
 sg13g2_xor2_1 _14078_ (.B(_06708_),
    .A(_06706_),
    .X(_06722_));
 sg13g2_nor2_1 _14079_ (.A(_06721_),
    .B(_06722_),
    .Y(_06723_));
 sg13g2_a21oi_1 _14080_ (.A1(net1855),
    .A2(_00172_),
    .Y(_06724_),
    .B1(net1641));
 sg13g2_inv_1 _14081_ (.Y(_06725_),
    .A(_06724_));
 sg13g2_nor2_1 _14082_ (.A(_00645_),
    .B(_00028_),
    .Y(_06726_));
 sg13g2_nand2b_1 _14083_ (.Y(_06727_),
    .B(net1855),
    .A_N(_00028_));
 sg13g2_xnor2_1 _14084_ (.Y(_06728_),
    .A(_00658_),
    .B(_06724_));
 sg13g2_nand2_1 _14085_ (.Y(_06729_),
    .A(_06727_),
    .B(_06728_));
 sg13g2_o21ai_1 _14086_ (.B1(_06729_),
    .Y(_06730_),
    .A1(_00658_),
    .A2(_06725_));
 sg13g2_xnor2_1 _14087_ (.Y(_06731_),
    .A(_06678_),
    .B(_06719_));
 sg13g2_nand2_1 _14088_ (.Y(_06732_),
    .A(_06730_),
    .B(_06731_));
 sg13g2_o21ai_1 _14089_ (.B1(_06716_),
    .Y(_06733_),
    .A1(_06723_),
    .A2(_06732_));
 sg13g2_a21oi_1 _14090_ (.A1(_06721_),
    .A2(_06722_),
    .Y(_06734_),
    .B1(_06733_));
 sg13g2_xnor2_1 _14091_ (.Y(_06735_),
    .A(net1799),
    .B(net1801));
 sg13g2_xor2_1 _14092_ (.B(net1801),
    .A(net1799),
    .X(_06736_));
 sg13g2_o21ai_1 _14093_ (.B1(_06736_),
    .Y(_06737_),
    .A1(_00032_),
    .A2(_06727_));
 sg13g2_o21ai_1 _14094_ (.B1(_06737_),
    .Y(_06738_),
    .A1(_06710_),
    .A2(_06726_));
 sg13g2_o21ai_1 _14095_ (.B1(_06732_),
    .Y(_06739_),
    .A1(_06717_),
    .A2(_06738_));
 sg13g2_nand2b_1 _14096_ (.Y(_06740_),
    .B(_06726_),
    .A_N(_06728_));
 sg13g2_a22oi_1 _14097_ (.Y(_06741_),
    .B1(_06740_),
    .B2(_06729_),
    .A2(_06738_),
    .A1(_06717_));
 sg13g2_nor2_1 _14098_ (.A(_06730_),
    .B(_06731_),
    .Y(_06742_));
 sg13g2_or4_1 _14099_ (.A(_06723_),
    .B(_06739_),
    .C(_06741_),
    .D(_06742_),
    .X(_06743_));
 sg13g2_a22oi_1 _14100_ (.Y(_06744_),
    .B1(_06734_),
    .B2(_06743_),
    .A2(_06715_),
    .A1(_06709_));
 sg13g2_a21oi_1 _14101_ (.A1(_06707_),
    .A2(_06711_),
    .Y(_06745_),
    .B1(_06710_));
 sg13g2_a21oi_1 _14102_ (.A1(_06710_),
    .A2(_06713_),
    .Y(_06746_),
    .B1(_06745_));
 sg13g2_nand2_1 _14103_ (.Y(_06747_),
    .A(_06744_),
    .B(_06746_));
 sg13g2_inv_1 _14104_ (.Y(_06748_),
    .A(_06747_));
 sg13g2_nor2_1 _14105_ (.A(_06744_),
    .B(_06746_),
    .Y(_06749_));
 sg13g2_or2_1 _14106_ (.X(_06750_),
    .B(_02981_),
    .A(_00651_));
 sg13g2_nand3_1 _14107_ (.B(_02944_),
    .C(_06750_),
    .A(_00652_),
    .Y(_06751_));
 sg13g2_nand2b_1 _14108_ (.Y(_06752_),
    .B(_06751_),
    .A_N(_00179_));
 sg13g2_a21oi_1 _14109_ (.A1(net2351),
    .A2(_02970_),
    .Y(_06753_),
    .B1(net2166));
 sg13g2_nor3_1 _14110_ (.A(net1913),
    .B(net1914),
    .C(_02980_),
    .Y(_06754_));
 sg13g2_nand3_1 _14111_ (.B(_02978_),
    .C(_06754_),
    .A(_02976_),
    .Y(_06755_));
 sg13g2_nand3_1 _14112_ (.B(_06753_),
    .C(_06755_),
    .A(_06752_),
    .Y(_06756_));
 sg13g2_nor3_1 _14113_ (.A(_06748_),
    .B(_06749_),
    .C(_06756_),
    .Y(_00532_));
 sg13g2_nor2_1 _14114_ (.A(_06745_),
    .B(_06748_),
    .Y(_06757_));
 sg13g2_nor2_1 _14115_ (.A(_06756_),
    .B(_06757_),
    .Y(_00533_));
 sg13g2_a21oi_2 _14116_ (.B1(net1640),
    .Y(_06758_),
    .A2(_00036_),
    .A1(net1856));
 sg13g2_nor2_1 _14117_ (.A(_06677_),
    .B(_06758_),
    .Y(_06759_));
 sg13g2_a21oi_2 _14118_ (.B1(net1641),
    .Y(_06760_),
    .A2(_00173_),
    .A1(net1856));
 sg13g2_nand2_1 _14119_ (.Y(_06761_),
    .A(_06677_),
    .B(_06758_));
 sg13g2_nand2b_1 _14120_ (.Y(_06762_),
    .B(_06761_),
    .A_N(_06759_));
 sg13g2_a21oi_1 _14121_ (.A1(_06760_),
    .A2(_06761_),
    .Y(_06763_),
    .B1(_06759_));
 sg13g2_nand2_1 _14122_ (.Y(_06764_),
    .A(net1856),
    .B(_00038_));
 sg13g2_nor2b_2 _14123_ (.A(net1640),
    .B_N(_06764_),
    .Y(_06765_));
 sg13g2_nand2_1 _14124_ (.Y(_06766_),
    .A(_06712_),
    .B(_06760_));
 sg13g2_nand2b_1 _14125_ (.Y(_06767_),
    .B(_06711_),
    .A_N(_06760_));
 sg13g2_nand2_1 _14126_ (.Y(_06768_),
    .A(_06766_),
    .B(_06767_));
 sg13g2_xnor2_1 _14127_ (.Y(_06769_),
    .A(_06765_),
    .B(_06768_));
 sg13g2_nor2_1 _14128_ (.A(_06763_),
    .B(_06769_),
    .Y(_06770_));
 sg13g2_a21oi_1 _14129_ (.A1(net1856),
    .A2(_00175_),
    .Y(_06771_),
    .B1(net1640));
 sg13g2_nand2_1 _14130_ (.Y(_06772_),
    .A(_00657_),
    .B(_06771_));
 sg13g2_a21oi_2 _14131_ (.B1(net1640),
    .Y(_06773_),
    .A2(_00034_),
    .A1(net1856));
 sg13g2_xnor2_1 _14132_ (.Y(_06774_),
    .A(_00657_),
    .B(_06771_));
 sg13g2_o21ai_1 _14133_ (.B1(_06772_),
    .Y(_06775_),
    .A1(_06773_),
    .A2(_06774_));
 sg13g2_a21oi_2 _14134_ (.B1(net1640),
    .Y(_06776_),
    .A2(_00174_),
    .A1(net1856));
 sg13g2_inv_1 _14135_ (.Y(_06777_),
    .A(_06776_));
 sg13g2_xnor2_1 _14136_ (.Y(_06778_),
    .A(_00659_),
    .B(_06776_));
 sg13g2_nand2b_1 _14137_ (.Y(_06779_),
    .B(_06778_),
    .A_N(_06758_));
 sg13g2_xnor2_1 _14138_ (.Y(_06780_),
    .A(_06758_),
    .B(_06778_));
 sg13g2_o21ai_1 _14139_ (.B1(_06773_),
    .Y(_06781_),
    .A1(_06735_),
    .A2(_06764_));
 sg13g2_nand2_1 _14140_ (.Y(_06782_),
    .A(_06735_),
    .B(_06765_));
 sg13g2_nand3_1 _14141_ (.B(_06781_),
    .C(_06782_),
    .A(_06776_),
    .Y(_06783_));
 sg13g2_a21oi_1 _14142_ (.A1(_06781_),
    .A2(_06782_),
    .Y(_06784_),
    .B1(_06776_));
 sg13g2_xnor2_1 _14143_ (.Y(_06785_),
    .A(_06773_),
    .B(_06774_));
 sg13g2_a21oi_1 _14144_ (.A1(_06783_),
    .A2(_06785_),
    .Y(_06786_),
    .B1(_06784_));
 sg13g2_o21ai_1 _14145_ (.B1(_06786_),
    .Y(_06787_),
    .A1(_06775_),
    .A2(_06780_));
 sg13g2_xnor2_1 _14146_ (.Y(_06788_),
    .A(_06760_),
    .B(_06762_));
 sg13g2_o21ai_1 _14147_ (.B1(_06779_),
    .Y(_06789_),
    .A1(_00659_),
    .A2(_06777_));
 sg13g2_a22oi_1 _14148_ (.Y(_06790_),
    .B1(_06788_),
    .B2(_06789_),
    .A2(_06780_),
    .A1(_06775_));
 sg13g2_nor2_1 _14149_ (.A(_06788_),
    .B(_06789_),
    .Y(_06791_));
 sg13g2_a221oi_1 _14150_ (.B2(_06790_),
    .C1(_06791_),
    .B1(_06787_),
    .A1(_06763_),
    .Y(_06792_),
    .A2(_06769_));
 sg13g2_nor2b_1 _14151_ (.A(_06765_),
    .B_N(_06767_),
    .Y(_06793_));
 sg13g2_nand2b_1 _14152_ (.Y(_06794_),
    .B(_06767_),
    .A_N(_06765_));
 sg13g2_a21oi_1 _14153_ (.A1(_06765_),
    .A2(_06766_),
    .Y(_06795_),
    .B1(_06793_));
 sg13g2_nor3_1 _14154_ (.A(_06770_),
    .B(_06792_),
    .C(_06795_),
    .Y(_06796_));
 sg13g2_o21ai_1 _14155_ (.B1(_06795_),
    .Y(_06797_),
    .A1(_06770_),
    .A2(_06792_));
 sg13g2_inv_1 _14156_ (.Y(_06798_),
    .A(_06797_));
 sg13g2_nor3_1 _14157_ (.A(_06756_),
    .B(_06796_),
    .C(_06798_),
    .Y(_00534_));
 sg13g2_a21oi_1 _14158_ (.A1(_06794_),
    .A2(_06797_),
    .Y(_00535_),
    .B1(_06756_));
 sg13g2_a21oi_2 _14159_ (.B1(net1640),
    .Y(_06799_),
    .A2(_00042_),
    .A1(net1857));
 sg13g2_nor2_1 _14160_ (.A(_06677_),
    .B(_06799_),
    .Y(_06800_));
 sg13g2_nand2_2 _14161_ (.Y(_06801_),
    .A(net1857),
    .B(net2342));
 sg13g2_xnor2_1 _14162_ (.Y(_06802_),
    .A(_06677_),
    .B(_06799_));
 sg13g2_nor2_1 _14163_ (.A(_06801_),
    .B(_06802_),
    .Y(_06803_));
 sg13g2_nor2_1 _14164_ (.A(_06800_),
    .B(_06803_),
    .Y(_06804_));
 sg13g2_a21oi_2 _14165_ (.B1(net1641),
    .Y(_06805_),
    .A2(_00044_),
    .A1(net1856));
 sg13g2_xnor2_1 _14166_ (.Y(_06806_),
    .A(_06711_),
    .B(_06801_));
 sg13g2_xnor2_1 _14167_ (.Y(_06807_),
    .A(_06805_),
    .B(_06806_));
 sg13g2_nand2_2 _14168_ (.Y(_06808_),
    .A(net1855),
    .B(_00041_));
 sg13g2_a21oi_2 _14169_ (.B1(net1640),
    .Y(_06809_),
    .A2(_00040_),
    .A1(net1855));
 sg13g2_nand2_1 _14170_ (.Y(_06810_),
    .A(net1855),
    .B(_00039_));
 sg13g2_nor2_1 _14171_ (.A(_00658_),
    .B(_06810_),
    .Y(_06811_));
 sg13g2_xnor2_1 _14172_ (.Y(_06812_),
    .A(_00658_),
    .B(_06810_));
 sg13g2_nor2_1 _14173_ (.A(_06809_),
    .B(_06812_),
    .Y(_06813_));
 sg13g2_xnor2_1 _14174_ (.Y(_06814_),
    .A(_06809_),
    .B(_06812_));
 sg13g2_nor2_1 _14175_ (.A(_06808_),
    .B(_06814_),
    .Y(_06815_));
 sg13g2_nand3_1 _14176_ (.B(_00044_),
    .C(_06736_),
    .A(net1855),
    .Y(_06816_));
 sg13g2_a22oi_1 _14177_ (.Y(_06817_),
    .B1(_06809_),
    .B2(_06816_),
    .A2(_06805_),
    .A1(_06735_));
 sg13g2_nor2_1 _14178_ (.A(_06815_),
    .B(_06817_),
    .Y(_06818_));
 sg13g2_xor2_1 _14179_ (.B(_06808_),
    .A(_00659_),
    .X(_06819_));
 sg13g2_nand2b_1 _14180_ (.Y(_06820_),
    .B(_06819_),
    .A_N(_06799_));
 sg13g2_xor2_1 _14181_ (.B(_06819_),
    .A(_06799_),
    .X(_06821_));
 sg13g2_nor2_1 _14182_ (.A(_06811_),
    .B(_06813_),
    .Y(_06822_));
 sg13g2_a221oi_1 _14183_ (.B2(_06822_),
    .C1(_06818_),
    .B1(_06821_),
    .A1(_06808_),
    .Y(_06823_),
    .A2(_06814_));
 sg13g2_o21ai_1 _14184_ (.B1(_06820_),
    .Y(_06824_),
    .A1(_00659_),
    .A2(_06808_));
 sg13g2_xor2_1 _14185_ (.B(_06802_),
    .A(_06801_),
    .X(_06825_));
 sg13g2_nand2_1 _14186_ (.Y(_06826_),
    .A(_06824_),
    .B(_06825_));
 sg13g2_o21ai_1 _14187_ (.B1(_06826_),
    .Y(_06827_),
    .A1(_06821_),
    .A2(_06822_));
 sg13g2_nor2_1 _14188_ (.A(_06824_),
    .B(_06825_),
    .Y(_06828_));
 sg13g2_a21oi_1 _14189_ (.A1(_06804_),
    .A2(_06807_),
    .Y(_06829_),
    .B1(_06828_));
 sg13g2_o21ai_1 _14190_ (.B1(_06829_),
    .Y(_06830_),
    .A1(_06823_),
    .A2(_06827_));
 sg13g2_o21ai_1 _14191_ (.B1(_06830_),
    .Y(_06831_),
    .A1(_06804_),
    .A2(_06807_));
 sg13g2_a21oi_1 _14192_ (.A1(_06711_),
    .A2(_06801_),
    .Y(_06832_),
    .B1(_06805_));
 sg13g2_o21ai_1 _14193_ (.B1(_06805_),
    .Y(_06833_),
    .A1(_06711_),
    .A2(_06801_));
 sg13g2_nor2b_1 _14194_ (.A(_06832_),
    .B_N(_06833_),
    .Y(_06834_));
 sg13g2_nor2_1 _14195_ (.A(_06831_),
    .B(_06834_),
    .Y(_06835_));
 sg13g2_and2_1 _14196_ (.A(_06831_),
    .B(_06834_),
    .X(_06836_));
 sg13g2_nor3_1 _14197_ (.A(_06756_),
    .B(_06835_),
    .C(_06836_),
    .Y(_00536_));
 sg13g2_nor2_1 _14198_ (.A(net2343),
    .B(_06836_),
    .Y(_06837_));
 sg13g2_nor2_1 _14199_ (.A(_06756_),
    .B(_06837_),
    .Y(_00537_));
 sg13g2_nand3_1 _14200_ (.B(net1741),
    .C(net1776),
    .A(net1974),
    .Y(_06838_));
 sg13g2_mux2_1 _14201_ (.A0(net1447),
    .A1(\vgadonut.donut.frame ),
    .S(_06838_),
    .X(_00538_));
 sg13g2_nand4_1 _14202_ (.B(net1972),
    .C(net1740),
    .A(net1799),
    .Y(_06839_),
    .D(net1776));
 sg13g2_nand4_1 _14203_ (.B(net1972),
    .C(net2033),
    .A(net1799),
    .Y(_06840_),
    .D(_04996_));
 sg13g2_xnor2_1 _14204_ (.Y(_00539_),
    .A(net2033),
    .B(_06839_));
 sg13g2_nor2_1 _14205_ (.A(_00647_),
    .B(_06840_),
    .Y(_06841_));
 sg13g2_xnor2_1 _14206_ (.Y(_00540_),
    .A(net2082),
    .B(_06840_));
 sg13g2_and2_1 _14207_ (.A(net2126),
    .B(_06841_),
    .X(_06842_));
 sg13g2_xor2_1 _14208_ (.B(_06841_),
    .A(net2126),
    .X(_00541_));
 sg13g2_xor2_1 _14209_ (.B(_06842_),
    .A(net2160),
    .X(_00542_));
 sg13g2_a21oi_1 _14210_ (.A1(\vgadonut.frame[4] ),
    .A2(_06842_),
    .Y(_06843_),
    .B1(net2102));
 sg13g2_nand3_1 _14211_ (.B(\vgadonut.frame[4] ),
    .C(_06842_),
    .A(\vgadonut.frame[5] ),
    .Y(_06844_));
 sg13g2_nor2b_1 _14212_ (.A(net2103),
    .B_N(_06844_),
    .Y(_00543_));
 sg13g2_or2_1 _14213_ (.X(_06845_),
    .B(_06844_),
    .A(_00646_));
 sg13g2_xnor2_1 _14214_ (.Y(_00544_),
    .A(net2089),
    .B(_06844_));
 sg13g2_nor3_1 _14215_ (.A(_00646_),
    .B(net2044),
    .C(_06844_),
    .Y(_06846_));
 sg13g2_a21o_1 _14216_ (.A2(_06845_),
    .A1(net2044),
    .B1(_06846_),
    .X(_00545_));
 sg13g2_dfrbp_1 _14217_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net19),
    .D(_00223_),
    .Q_N(_07140_),
    .Q(\vgadonut.donut.rx6[0] ));
 sg13g2_dfrbp_1 _14218_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net20),
    .D(_00224_),
    .Q_N(_07141_),
    .Q(\vgadonut.donut.rx6[1] ));
 sg13g2_dfrbp_1 _14219_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net21),
    .D(_00009_),
    .Q_N(_07142_),
    .Q(_00039_));
 sg13g2_dfrbp_1 _14220_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net22),
    .D(_00010_),
    .Q_N(_07143_),
    .Q(_00040_));
 sg13g2_dfrbp_1 _14221_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net23),
    .D(_00011_),
    .Q_N(_07144_),
    .Q(_00041_));
 sg13g2_dfrbp_1 _14222_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net24),
    .D(_00012_),
    .Q_N(_07145_),
    .Q(_00042_));
 sg13g2_dfrbp_1 _14223_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net25),
    .D(_00013_),
    .Q_N(_07146_),
    .Q(_00043_));
 sg13g2_dfrbp_1 _14224_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net26),
    .D(_00004_),
    .Q_N(_00175_),
    .Q(_00033_));
 sg13g2_dfrbp_1 _14225_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net27),
    .D(_00005_),
    .Q_N(_07147_),
    .Q(_00034_));
 sg13g2_dfrbp_1 _14226_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net28),
    .D(_00006_),
    .Q_N(_00174_),
    .Q(_00035_));
 sg13g2_dfrbp_1 _14227_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net29),
    .D(_00007_),
    .Q_N(_07148_),
    .Q(_00036_));
 sg13g2_dfrbp_1 _14228_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net30),
    .D(_00008_),
    .Q_N(_00173_),
    .Q(_00037_));
 sg13g2_dfrbp_1 _14229_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net31),
    .D(_00000_),
    .Q_N(_00172_),
    .Q(_00027_));
 sg13g2_dfrbp_1 _14230_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net32),
    .D(_00001_),
    .Q_N(_07149_),
    .Q(_00028_));
 sg13g2_dfrbp_1 _14231_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net162),
    .D(_00002_),
    .Q_N(_00171_),
    .Q(_00029_));
 sg13g2_dfrbp_1 _14232_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net56),
    .D(_00003_),
    .Q_N(_07139_),
    .Q(_00030_));
 sg13g2_dfrbp_1 _14233_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net54),
    .D(_00225_),
    .Q_N(_07138_),
    .Q(_00032_));
 sg13g2_dfrbp_1 _14234_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net53),
    .D(_00226_),
    .Q_N(_07137_),
    .Q(\vgadonut.donut.donuthit.t[0] ));
 sg13g2_dfrbp_1 _14235_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net52),
    .D(_00227_),
    .Q_N(_07136_),
    .Q(\vgadonut.donut.donuthit.t[1] ));
 sg13g2_dfrbp_1 _14236_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net51),
    .D(_00228_),
    .Q_N(_07135_),
    .Q(\vgadonut.donut.donuthit.t[2] ));
 sg13g2_dfrbp_1 _14237_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net50),
    .D(net2250),
    .Q_N(_07134_),
    .Q(\vgadonut.donut.donuthit.t[3] ));
 sg13g2_dfrbp_1 _14238_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net49),
    .D(_00230_),
    .Q_N(_07133_),
    .Q(\vgadonut.donut.donuthit.t[4] ));
 sg13g2_dfrbp_1 _14239_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net48),
    .D(net2208),
    .Q_N(_07132_),
    .Q(\vgadonut.donut.donuthit.t[5] ));
 sg13g2_dfrbp_1 _14240_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net47),
    .D(_00232_),
    .Q_N(_07131_),
    .Q(\vgadonut.donut.donuthit.t[6] ));
 sg13g2_dfrbp_1 _14241_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net46),
    .D(_00233_),
    .Q_N(_07130_),
    .Q(\vgadonut.donut.donuthit.t[7] ));
 sg13g2_dfrbp_1 _14242_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net45),
    .D(net2258),
    .Q_N(_07129_),
    .Q(\vgadonut.donut.donuthit.t[8] ));
 sg13g2_dfrbp_1 _14243_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net44),
    .D(_00235_),
    .Q_N(_07128_),
    .Q(\vgadonut.donut.donuthit.t[9] ));
 sg13g2_dfrbp_1 _14244_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net43),
    .D(net2301),
    .Q_N(_07127_),
    .Q(\vgadonut.donut.donuthit.t[10] ));
 sg13g2_dfrbp_1 _14245_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net42),
    .D(_00237_),
    .Q_N(_07126_),
    .Q(\vgadonut.donut.donuthit.t[11] ));
 sg13g2_dfrbp_1 _14246_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net41),
    .D(_00238_),
    .Q_N(_07125_),
    .Q(\vgadonut.donut.donuthit.t[12] ));
 sg13g2_dfrbp_1 _14247_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net40),
    .D(_00239_),
    .Q_N(_07124_),
    .Q(\vgadonut.donut.donuthit.t[13] ));
 sg13g2_dfrbp_1 _14248_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net39),
    .D(_00240_),
    .Q_N(_07123_),
    .Q(\vgadonut.donut.donuthit.t[14] ));
 sg13g2_dfrbp_1 _14249_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net38),
    .D(_00241_),
    .Q_N(_07122_),
    .Q(\vgadonut.donut.donuthit.t[15] ));
 sg13g2_dfrbp_1 _14250_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net37),
    .D(_00242_),
    .Q_N(_07121_),
    .Q(_00038_));
 sg13g2_dfrbp_1 _14251_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net36),
    .D(_00243_),
    .Q_N(_07120_),
    .Q(\vgadonut.donut.ysA[4] ));
 sg13g2_dfrbp_1 _14252_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net35),
    .D(net2211),
    .Q_N(_07119_),
    .Q(\vgadonut.donut.ysA[5] ));
 sg13g2_dfrbp_1 _14253_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net34),
    .D(_00245_),
    .Q_N(_07118_),
    .Q(\vgadonut.donut.ysA[6] ));
 sg13g2_dfrbp_1 _14254_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net33),
    .D(_00246_),
    .Q_N(_07117_),
    .Q(\vgadonut.donut.ysA[7] ));
 sg13g2_dfrbp_1 _14255_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net18),
    .D(_00247_),
    .Q_N(_07116_),
    .Q(\vgadonut.donut.ysA[8] ));
 sg13g2_dfrbp_1 _14256_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net17),
    .D(_00248_),
    .Q_N(_07115_),
    .Q(\vgadonut.donut.ysA[9] ));
 sg13g2_dfrbp_1 _14257_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net271),
    .D(_00249_),
    .Q_N(_07114_),
    .Q(\vgadonut.donut.ysA[10] ));
 sg13g2_dfrbp_1 _14258_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net270),
    .D(_00250_),
    .Q_N(_07113_),
    .Q(\vgadonut.donut.ysA[11] ));
 sg13g2_dfrbp_1 _14259_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net269),
    .D(_00251_),
    .Q_N(_07112_),
    .Q(\vgadonut.donut.ysA[12] ));
 sg13g2_dfrbp_1 _14260_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net268),
    .D(_00252_),
    .Q_N(_07111_),
    .Q(\vgadonut.donut.ysA[13] ));
 sg13g2_dfrbp_1 _14261_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net267),
    .D(_00253_),
    .Q_N(_07110_),
    .Q(\vgadonut.donut.ysA[14] ));
 sg13g2_dfrbp_1 _14262_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net266),
    .D(_00254_),
    .Q_N(_07109_),
    .Q(\vgadonut.donut.ysA[15] ));
 sg13g2_dfrbp_1 _14263_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net265),
    .D(_00255_),
    .Q_N(_07108_),
    .Q(\vgadonut.donut.ysA[16] ));
 sg13g2_dfrbp_1 _14264_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net264),
    .D(_00256_),
    .Q_N(_07107_),
    .Q(\vgadonut.donut.ysA[17] ));
 sg13g2_dfrbp_1 _14265_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net262),
    .D(_00257_),
    .Q_N(_07106_),
    .Q(\vgadonut.donut.ysA[18] ));
 sg13g2_dfrbp_1 _14266_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net261),
    .D(_00258_),
    .Q_N(_07105_),
    .Q(\vgadonut.donut.ysA[19] ));
 sg13g2_dfrbp_1 _14267_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net260),
    .D(_00259_),
    .Q_N(_07104_),
    .Q(\vgadonut.donut.ysA[20] ));
 sg13g2_dfrbp_1 _14268_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net259),
    .D(_00260_),
    .Q_N(_07103_),
    .Q(\vgadonut.donut.ysA[21] ));
 sg13g2_dfrbp_1 _14269_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net256),
    .D(net2185),
    .Q_N(_07102_),
    .Q(\vgadonut.donut.ycA[4] ));
 sg13g2_dfrbp_1 _14270_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net255),
    .D(_00262_),
    .Q_N(_07101_),
    .Q(\vgadonut.donut.ycA[5] ));
 sg13g2_dfrbp_1 _14271_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net254),
    .D(_00263_),
    .Q_N(_07100_),
    .Q(\vgadonut.donut.ycA[6] ));
 sg13g2_dfrbp_1 _14272_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net253),
    .D(_00264_),
    .Q_N(_07099_),
    .Q(\vgadonut.donut.ycA[7] ));
 sg13g2_dfrbp_1 _14273_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net252),
    .D(net2195),
    .Q_N(_07098_),
    .Q(\vgadonut.donut.ycA[8] ));
 sg13g2_dfrbp_1 _14274_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net251),
    .D(_00266_),
    .Q_N(_07097_),
    .Q(\vgadonut.donut.ycA[9] ));
 sg13g2_dfrbp_1 _14275_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net250),
    .D(_00267_),
    .Q_N(_07096_),
    .Q(\vgadonut.donut.ycA[10] ));
 sg13g2_dfrbp_1 _14276_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net249),
    .D(_00268_),
    .Q_N(_07095_),
    .Q(\vgadonut.donut.ycA[11] ));
 sg13g2_dfrbp_1 _14277_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net248),
    .D(_00269_),
    .Q_N(_07094_),
    .Q(\vgadonut.donut.ycA[12] ));
 sg13g2_dfrbp_1 _14278_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net247),
    .D(_00270_),
    .Q_N(_07093_),
    .Q(\vgadonut.donut.ycA[13] ));
 sg13g2_dfrbp_1 _14279_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net246),
    .D(_00271_),
    .Q_N(_07092_),
    .Q(\vgadonut.donut.ycA[14] ));
 sg13g2_dfrbp_1 _14280_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net245),
    .D(_00272_),
    .Q_N(_07091_),
    .Q(\vgadonut.donut.ycA[15] ));
 sg13g2_dfrbp_1 _14281_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net244),
    .D(_00273_),
    .Q_N(_07090_),
    .Q(\vgadonut.donut.ycA[16] ));
 sg13g2_dfrbp_1 _14282_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net243),
    .D(_00274_),
    .Q_N(_07089_),
    .Q(\vgadonut.donut.ycA[17] ));
 sg13g2_dfrbp_1 _14283_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net242),
    .D(_00275_),
    .Q_N(_07088_),
    .Q(\vgadonut.donut.ycA[18] ));
 sg13g2_dfrbp_1 _14284_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net241),
    .D(_00276_),
    .Q_N(_07087_),
    .Q(\vgadonut.donut.ycA[19] ));
 sg13g2_dfrbp_1 _14285_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net240),
    .D(_00277_),
    .Q_N(_07086_),
    .Q(\vgadonut.donut.ycA[20] ));
 sg13g2_dfrbp_1 _14286_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net239),
    .D(_00278_),
    .Q_N(_07085_),
    .Q(\vgadonut.donut.ycA[21] ));
 sg13g2_dfrbp_1 _14287_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net238),
    .D(_00279_),
    .Q_N(_07084_),
    .Q(\vgadonut.donut.ycA[0] ));
 sg13g2_dfrbp_1 _14288_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net237),
    .D(_00280_),
    .Q_N(_07083_),
    .Q(\vgadonut.donut.ycA[1] ));
 sg13g2_dfrbp_1 _14289_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net236),
    .D(_00281_),
    .Q_N(_07082_),
    .Q(\vgadonut.donut.ycA[2] ));
 sg13g2_dfrbp_1 _14290_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net235),
    .D(_00282_),
    .Q_N(_00106_),
    .Q(\vgadonut.donut.ycA[3] ));
 sg13g2_dfrbp_1 _14291_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net233),
    .D(_00283_),
    .Q_N(_07081_),
    .Q(_00044_));
 sg13g2_dfrbp_1 _14292_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net232),
    .D(_00284_),
    .Q_N(_07080_),
    .Q(\vgadonut.donut.ysA[0] ));
 sg13g2_dfrbp_1 _14293_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net230),
    .D(_00285_),
    .Q_N(_07079_),
    .Q(\vgadonut.donut.ysA[1] ));
 sg13g2_dfrbp_1 _14294_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net229),
    .D(_00286_),
    .Q_N(_07078_),
    .Q(\vgadonut.donut.ysA[2] ));
 sg13g2_dfrbp_1 _14295_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net228),
    .D(_00287_),
    .Q_N(_07077_),
    .Q(\vgadonut.donut.ysA[3] ));
 sg13g2_dfrbp_1 _14296_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net178),
    .D(net2008),
    .Q_N(_07076_),
    .Q(\vgadonut.donut.donut_luma[0] ));
 sg13g2_dfrbp_1 _14297_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net177),
    .D(_00289_),
    .Q_N(_07075_),
    .Q(\vgadonut.donut.donut_luma[1] ));
 sg13g2_dfrbp_1 _14298_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net176),
    .D(_00290_),
    .Q_N(_07074_),
    .Q(\vgadonut.donut.donut_luma[2] ));
 sg13g2_dfrbp_1 _14299_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net175),
    .D(_00291_),
    .Q_N(_07073_),
    .Q(\vgadonut.donut.donut_luma[3] ));
 sg13g2_dfrbp_1 _14300_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net174),
    .D(net1639),
    .Q_N(_07072_),
    .Q(\vgadonut.donut.donut_luma[4] ));
 sg13g2_dfrbp_1 _14301_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net173),
    .D(net1631),
    .Q_N(_07071_),
    .Q(\vgadonut.donut.donut_luma[5] ));
 sg13g2_dfrbp_1 _14302_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1959),
    .D(_00294_),
    .Q_N(\vgadonut.donut.cAcB[0] ),
    .Q(_00182_));
 sg13g2_dfrbp_1 _14303_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1959),
    .D(_00295_),
    .Q_N(\vgadonut.donut.cAcB[1] ),
    .Q(_00183_));
 sg13g2_dfrbp_1 _14304_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1959),
    .D(_00296_),
    .Q_N(\vgadonut.donut.cAcB[2] ),
    .Q(_00184_));
 sg13g2_dfrbp_1 _14305_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1959),
    .D(_00297_),
    .Q_N(\vgadonut.donut.cAcB[3] ),
    .Q(_00185_));
 sg13g2_dfrbp_1 _14306_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1963),
    .D(_00298_),
    .Q_N(\vgadonut.donut.cAcB[4] ),
    .Q(_00186_));
 sg13g2_dfrbp_1 _14307_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1963),
    .D(_00299_),
    .Q_N(\vgadonut.donut.cAcB[5] ),
    .Q(_00187_));
 sg13g2_dfrbp_1 _14308_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1963),
    .D(_00300_),
    .Q_N(_07070_),
    .Q(\vgadonut.donut.cAcB[6] ));
 sg13g2_dfrbp_1 _14309_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1964),
    .D(_00301_),
    .Q_N(_07069_),
    .Q(\vgadonut.donut.cAcB[7] ));
 sg13g2_dfrbp_1 _14310_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1964),
    .D(_00302_),
    .Q_N(\vgadonut.donut.cAcB[8] ),
    .Q(_00188_));
 sg13g2_dfrbp_1 _14311_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1964),
    .D(_00303_),
    .Q_N(_07068_),
    .Q(\vgadonut.donut.cAcB[9] ));
 sg13g2_dfrbp_1 _14312_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1964),
    .D(_00304_),
    .Q_N(\vgadonut.donut.cAcB[10] ),
    .Q(_00189_));
 sg13g2_dfrbp_1 _14313_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1965),
    .D(_00305_),
    .Q_N(\vgadonut.donut.cAcB[11] ),
    .Q(_00190_));
 sg13g2_dfrbp_1 _14314_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1964),
    .D(_00306_),
    .Q_N(_07067_),
    .Q(\vgadonut.donut.cAcB[12] ));
 sg13g2_dfrbp_1 _14315_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1964),
    .D(_00307_),
    .Q_N(\vgadonut.donut.cAcB[13] ),
    .Q(_00191_));
 sg13g2_dfrbp_1 _14316_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1964),
    .D(_00308_),
    .Q_N(_07066_),
    .Q(\vgadonut.donut.cAcB[14] ));
 sg13g2_dfrbp_1 _14317_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1984),
    .D(_00309_),
    .Q_N(_07065_),
    .Q(\vgadonut.donut.cAcB[15] ));
 sg13g2_dfrbp_1 _14318_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1961),
    .D(net1476),
    .Q_N(\vgadonut.donut.sAcB[0] ),
    .Q(_00192_));
 sg13g2_dfrbp_1 _14319_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1961),
    .D(_00311_),
    .Q_N(\vgadonut.donut.sAcB[1] ),
    .Q(_00193_));
 sg13g2_dfrbp_1 _14320_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1961),
    .D(_00312_),
    .Q_N(\vgadonut.donut.sAcB[2] ),
    .Q(_00194_));
 sg13g2_dfrbp_1 _14321_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1962),
    .D(_00313_),
    .Q_N(\vgadonut.donut.sAcB[3] ),
    .Q(_00195_));
 sg13g2_dfrbp_1 _14322_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1977),
    .D(_00314_),
    .Q_N(\vgadonut.donut.sAcB[4] ),
    .Q(_00196_));
 sg13g2_dfrbp_1 _14323_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1977),
    .D(_00315_),
    .Q_N(\vgadonut.donut.sAcB[5] ),
    .Q(_00197_));
 sg13g2_dfrbp_1 _14324_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1962),
    .D(_00316_),
    .Q_N(_00108_),
    .Q(\vgadonut.donut.sAcB[6] ));
 sg13g2_dfrbp_1 _14325_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1962),
    .D(_00317_),
    .Q_N(_00109_),
    .Q(\vgadonut.donut.sAcB[7] ));
 sg13g2_dfrbp_1 _14326_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1961),
    .D(_00318_),
    .Q_N(\vgadonut.donut.sAcB[8] ),
    .Q(_00198_));
 sg13g2_dfrbp_1 _14327_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1962),
    .D(_00319_),
    .Q_N(_00111_),
    .Q(\vgadonut.donut.sAcB[9] ));
 sg13g2_dfrbp_1 _14328_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1961),
    .D(_00320_),
    .Q_N(\vgadonut.donut.sAcB[10] ),
    .Q(_00199_));
 sg13g2_dfrbp_1 _14329_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1977),
    .D(_00321_),
    .Q_N(\vgadonut.donut.sAcB[11] ),
    .Q(_00200_));
 sg13g2_dfrbp_1 _14330_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1978),
    .D(_00322_),
    .Q_N(_00112_),
    .Q(\vgadonut.donut.sAcB[12] ));
 sg13g2_dfrbp_1 _14331_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1977),
    .D(_00323_),
    .Q_N(\vgadonut.donut.sAcB[13] ),
    .Q(_00201_));
 sg13g2_dfrbp_1 _14332_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1977),
    .D(_00324_),
    .Q_N(_00113_),
    .Q(\vgadonut.donut.sAcB[14] ));
 sg13g2_dfrbp_1 _14333_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1978),
    .D(_00325_),
    .Q_N(_07064_),
    .Q(\vgadonut.donut.sAcB[15] ));
 sg13g2_dfrbp_1 _14334_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1974),
    .D(_00326_),
    .Q_N(_07063_),
    .Q(\vgadonut.bayer_j[0] ));
 sg13g2_dfrbp_1 _14335_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1975),
    .D(_00327_),
    .Q_N(_07062_),
    .Q(\vgadonut.bayer_j[1] ));
 sg13g2_dfrbp_1 _14336_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1972),
    .D(_00328_),
    .Q_N(_07061_),
    .Q(\vgadonut.donut.v_count[2] ));
 sg13g2_dfrbp_1 _14337_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1973),
    .D(_00329_),
    .Q_N(_07060_),
    .Q(\vgadonut.donut.v_count[3] ));
 sg13g2_dfrbp_1 _14338_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1973),
    .D(net2236),
    .Q_N(_07059_),
    .Q(\vgadonut.donut.v_count[4] ));
 sg13g2_dfrbp_1 _14339_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1972),
    .D(net2147),
    .Q_N(_00180_),
    .Q(\vgadonut.donut.v_count[5] ));
 sg13g2_dfrbp_1 _14340_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1971),
    .D(net2113),
    .Q_N(_07058_),
    .Q(\vgadonut.donut.v_count[6] ));
 sg13g2_dfrbp_1 _14341_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1973),
    .D(net2027),
    .Q_N(_07057_),
    .Q(\vgadonut.donut.v_count[7] ));
 sg13g2_dfrbp_1 _14342_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1973),
    .D(net2070),
    .Q_N(_07056_),
    .Q(\vgadonut.donut.v_count[8] ));
 sg13g2_dfrbp_1 _14343_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1972),
    .D(_00335_),
    .Q_N(_07055_),
    .Q(\vgadonut.donut.v_count[9] ));
 sg13g2_dfrbp_1 _14344_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1959),
    .D(_00336_),
    .Q_N(_00094_),
    .Q(\vgadonut.donut.cAsB[0] ));
 sg13g2_dfrbp_1 _14345_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1959),
    .D(_00337_),
    .Q_N(_00095_),
    .Q(\vgadonut.donut.cAsB[1] ));
 sg13g2_dfrbp_1 _14346_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1963),
    .D(_00338_),
    .Q_N(_00096_),
    .Q(\vgadonut.donut.cAsB[2] ));
 sg13g2_dfrbp_1 _14347_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1965),
    .D(_00339_),
    .Q_N(_00097_),
    .Q(\vgadonut.donut.cAsB[3] ));
 sg13g2_dfrbp_1 _14348_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1965),
    .D(_00340_),
    .Q_N(_00098_),
    .Q(\vgadonut.donut.cAsB[4] ));
 sg13g2_dfrbp_1 _14349_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1963),
    .D(_00341_),
    .Q_N(_00099_),
    .Q(\vgadonut.donut.cAsB[5] ));
 sg13g2_dfrbp_1 _14350_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1963),
    .D(_00342_),
    .Q_N(_00100_),
    .Q(\vgadonut.donut.cAsB[6] ));
 sg13g2_dfrbp_1 _14351_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1963),
    .D(_00343_),
    .Q_N(_00101_),
    .Q(\vgadonut.donut.cAsB[7] ));
 sg13g2_dfrbp_1 _14352_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1963),
    .D(_00344_),
    .Q_N(_00102_),
    .Q(\vgadonut.donut.cAsB[8] ));
 sg13g2_dfrbp_1 _14353_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1976),
    .D(_00345_),
    .Q_N(_00103_),
    .Q(\vgadonut.donut.cAsB[9] ));
 sg13g2_dfrbp_1 _14354_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1976),
    .D(_00346_),
    .Q_N(_00104_),
    .Q(\vgadonut.donut.cAsB[10] ));
 sg13g2_dfrbp_1 _14355_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1976),
    .D(_00347_),
    .Q_N(_00105_),
    .Q(\vgadonut.donut.cAsB[11] ));
 sg13g2_dfrbp_1 _14356_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1976),
    .D(_00348_),
    .Q_N(_07054_),
    .Q(\vgadonut.donut.cAsB[12] ));
 sg13g2_dfrbp_1 _14357_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1976),
    .D(_00349_),
    .Q_N(_07053_),
    .Q(\vgadonut.donut.cAsB[13] ));
 sg13g2_dfrbp_1 _14358_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1976),
    .D(_00350_),
    .Q_N(_07052_),
    .Q(\vgadonut.donut.cAsB[14] ));
 sg13g2_dfrbp_1 _14359_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1979),
    .D(_00351_),
    .Q_N(_07051_),
    .Q(\vgadonut.donut.cAsB[15] ));
 sg13g2_dfrbp_1 _14360_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1958),
    .D(_00352_),
    .Q_N(_00107_),
    .Q(\vgadonut.donut.sAsB[0] ));
 sg13g2_dfrbp_1 _14361_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1958),
    .D(_00353_),
    .Q_N(_07050_),
    .Q(\vgadonut.donut.sAsB[1] ));
 sg13g2_dfrbp_1 _14362_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1960),
    .D(_00354_),
    .Q_N(_07049_),
    .Q(\vgadonut.donut.sAsB[2] ));
 sg13g2_dfrbp_1 _14363_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1960),
    .D(_00355_),
    .Q_N(_00139_),
    .Q(\vgadonut.donut.sAsB[3] ));
 sg13g2_dfrbp_1 _14364_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1960),
    .D(_00356_),
    .Q_N(_07048_),
    .Q(\vgadonut.donut.sAsB[4] ));
 sg13g2_dfrbp_1 _14365_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1961),
    .D(_00357_),
    .Q_N(_07047_),
    .Q(\vgadonut.donut.sAsB[5] ));
 sg13g2_dfrbp_1 _14366_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1961),
    .D(_00358_),
    .Q_N(_07046_),
    .Q(\vgadonut.donut.sAsB[6] ));
 sg13g2_dfrbp_1 _14367_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1961),
    .D(_00359_),
    .Q_N(_07045_),
    .Q(\vgadonut.donut.sAsB[7] ));
 sg13g2_dfrbp_1 _14368_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1962),
    .D(_00360_),
    .Q_N(_07044_),
    .Q(\vgadonut.donut.sAsB[8] ));
 sg13g2_dfrbp_1 _14369_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1962),
    .D(_00361_),
    .Q_N(_07043_),
    .Q(\vgadonut.donut.sAsB[9] ));
 sg13g2_dfrbp_1 _14370_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1977),
    .D(_00362_),
    .Q_N(_07042_),
    .Q(\vgadonut.donut.sAsB[10] ));
 sg13g2_dfrbp_1 _14371_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1977),
    .D(_00363_),
    .Q_N(_07041_),
    .Q(\vgadonut.donut.sAsB[11] ));
 sg13g2_dfrbp_1 _14372_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1977),
    .D(_00364_),
    .Q_N(_07040_),
    .Q(\vgadonut.donut.sAsB[12] ));
 sg13g2_dfrbp_1 _14373_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1962),
    .D(_00365_),
    .Q_N(_07039_),
    .Q(\vgadonut.donut.sAsB[13] ));
 sg13g2_dfrbp_1 _14374_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1962),
    .D(_00366_),
    .Q_N(_00140_),
    .Q(\vgadonut.donut.sAsB[14] ));
 sg13g2_dfrbp_1 _14375_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1964),
    .D(_00367_),
    .Q_N(_07038_),
    .Q(\vgadonut.donut.sAsB[15] ));
 sg13g2_dfrbp_1 _14376_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net131),
    .D(_00368_),
    .Q_N(_07037_),
    .Q(\vgadonut.donut.ry6[0] ));
 sg13g2_dfrbp_1 _14377_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net130),
    .D(net2010),
    .Q_N(_07036_),
    .Q(\vgadonut.donut.ry6[1] ));
 sg13g2_dfrbp_1 _14378_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net129),
    .D(_00370_),
    .Q_N(_07035_),
    .Q(\vgadonut.donut.ry6[2] ));
 sg13g2_dfrbp_1 _14379_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net128),
    .D(_00371_),
    .Q_N(_07034_),
    .Q(\vgadonut.donut.ry6[3] ));
 sg13g2_dfrbp_1 _14380_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net127),
    .D(_00372_),
    .Q_N(_07033_),
    .Q(\vgadonut.donut.ry6[4] ));
 sg13g2_dfrbp_1 _14381_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net126),
    .D(_00373_),
    .Q_N(_07032_),
    .Q(\vgadonut.donut.ry6[5] ));
 sg13g2_dfrbp_1 _14382_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net125),
    .D(net2081),
    .Q_N(_07031_),
    .Q(\vgadonut.donut.donuthit.ryin[0] ));
 sg13g2_dfrbp_1 _14383_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net124),
    .D(_00375_),
    .Q_N(_07030_),
    .Q(\vgadonut.donut.donuthit.ryin[1] ));
 sg13g2_dfrbp_1 _14384_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net123),
    .D(_00376_),
    .Q_N(_07029_),
    .Q(\vgadonut.donut.donuthit.ryin[2] ));
 sg13g2_dfrbp_1 _14385_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net122),
    .D(_00377_),
    .Q_N(_07028_),
    .Q(\vgadonut.donut.donuthit.ryin[3] ));
 sg13g2_dfrbp_1 _14386_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net121),
    .D(_00378_),
    .Q_N(_07027_),
    .Q(\vgadonut.donut.donuthit.ryin[4] ));
 sg13g2_dfrbp_1 _14387_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net120),
    .D(_00379_),
    .Q_N(_07026_),
    .Q(\vgadonut.donut.donuthit.ryin[5] ));
 sg13g2_dfrbp_1 _14388_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net119),
    .D(_00380_),
    .Q_N(_00110_),
    .Q(\vgadonut.donut.donuthit.ryin[6] ));
 sg13g2_dfrbp_1 _14389_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net118),
    .D(_00381_),
    .Q_N(_07025_),
    .Q(\vgadonut.donut.donuthit.ryin[7] ));
 sg13g2_dfrbp_1 _14390_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net117),
    .D(_00382_),
    .Q_N(_07024_),
    .Q(\vgadonut.donut.donuthit.ryin[8] ));
 sg13g2_dfrbp_1 _14391_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net116),
    .D(_00383_),
    .Q_N(_07023_),
    .Q(\vgadonut.donut.donuthit.ryin[9] ));
 sg13g2_dfrbp_1 _14392_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net115),
    .D(_00384_),
    .Q_N(_07022_),
    .Q(\vgadonut.donut.donuthit.ryin[10] ));
 sg13g2_dfrbp_1 _14393_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net114),
    .D(_00385_),
    .Q_N(_07021_),
    .Q(\vgadonut.donut.donuthit.ryin[11] ));
 sg13g2_dfrbp_1 _14394_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net113),
    .D(_00386_),
    .Q_N(_07020_),
    .Q(\vgadonut.donut.donuthit.ryin[12] ));
 sg13g2_dfrbp_1 _14395_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net112),
    .D(_00387_),
    .Q_N(_00114_),
    .Q(\vgadonut.donut.donuthit.ryin[13] ));
 sg13g2_dfrbp_1 _14396_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net111),
    .D(_00388_),
    .Q_N(_07019_),
    .Q(\vgadonut.donut.donuthit.ryin[14] ));
 sg13g2_dfrbp_1 _14397_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net110),
    .D(_00389_),
    .Q_N(_00165_),
    .Q(\vgadonut.donut.donuthit.ryin[15] ));
 sg13g2_dfrbp_1 _14398_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net109),
    .D(net2013),
    .Q_N(_07018_),
    .Q(\vgadonut.donut.rx6[2] ));
 sg13g2_dfrbp_1 _14399_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net108),
    .D(_00391_),
    .Q_N(_07017_),
    .Q(\vgadonut.donut.rx6[3] ));
 sg13g2_dfrbp_1 _14400_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net107),
    .D(net2061),
    .Q_N(_07016_),
    .Q(\vgadonut.donut.rx6[4] ));
 sg13g2_dfrbp_1 _14401_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net106),
    .D(_00393_),
    .Q_N(_07015_),
    .Q(\vgadonut.donut.rx6[5] ));
 sg13g2_dfrbp_1 _14402_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net105),
    .D(_00394_),
    .Q_N(_07014_),
    .Q(\vgadonut.donut.donuthit.rxin[0] ));
 sg13g2_dfrbp_1 _14403_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net104),
    .D(_00395_),
    .Q_N(_07013_),
    .Q(\vgadonut.donut.donuthit.rxin[1] ));
 sg13g2_dfrbp_1 _14404_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net103),
    .D(_00396_),
    .Q_N(_07012_),
    .Q(\vgadonut.donut.donuthit.rxin[2] ));
 sg13g2_dfrbp_1 _14405_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net102),
    .D(_00397_),
    .Q_N(_07011_),
    .Q(\vgadonut.donut.donuthit.rxin[3] ));
 sg13g2_dfrbp_1 _14406_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net101),
    .D(_00398_),
    .Q_N(_07010_),
    .Q(\vgadonut.donut.donuthit.rxin[4] ));
 sg13g2_dfrbp_1 _14407_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net100),
    .D(_00399_),
    .Q_N(_07009_),
    .Q(\vgadonut.donut.donuthit.rxin[5] ));
 sg13g2_dfrbp_1 _14408_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net99),
    .D(_00400_),
    .Q_N(_07008_),
    .Q(\vgadonut.donut.donuthit.rxin[6] ));
 sg13g2_dfrbp_1 _14409_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net98),
    .D(_00401_),
    .Q_N(_07007_),
    .Q(\vgadonut.donut.donuthit.rxin[7] ));
 sg13g2_dfrbp_1 _14410_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net97),
    .D(_00402_),
    .Q_N(_07006_),
    .Q(\vgadonut.donut.donuthit.rxin[8] ));
 sg13g2_dfrbp_1 _14411_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net96),
    .D(_00403_),
    .Q_N(_07005_),
    .Q(\vgadonut.donut.donuthit.rxin[9] ));
 sg13g2_dfrbp_1 _14412_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net95),
    .D(_00404_),
    .Q_N(_07004_),
    .Q(\vgadonut.donut.donuthit.rxin[10] ));
 sg13g2_dfrbp_1 _14413_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net94),
    .D(_00405_),
    .Q_N(_07003_),
    .Q(\vgadonut.donut.donuthit.rxin[11] ));
 sg13g2_dfrbp_1 _14414_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net93),
    .D(_00406_),
    .Q_N(_07002_),
    .Q(\vgadonut.donut.donuthit.rxin[12] ));
 sg13g2_dfrbp_1 _14415_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net92),
    .D(_00407_),
    .Q_N(_07001_),
    .Q(\vgadonut.donut.donuthit.rxin[13] ));
 sg13g2_dfrbp_1 _14416_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net91),
    .D(_00408_),
    .Q_N(_07000_),
    .Q(\vgadonut.donut.donuthit.rxin[14] ));
 sg13g2_dfrbp_1 _14417_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net90),
    .D(_00409_),
    .Q_N(_00160_),
    .Q(\vgadonut.donut.donuthit.rxin[15] ));
 sg13g2_dfrbp_1 _14418_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1980),
    .D(_00410_),
    .Q_N(_06999_),
    .Q(\vgadonut.donut.sB[0] ));
 sg13g2_dfrbp_1 _14419_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1980),
    .D(net2169),
    .Q_N(_06998_),
    .Q(\vgadonut.donut.sB[1] ));
 sg13g2_dfrbp_1 _14420_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1979),
    .D(_00412_),
    .Q_N(_00138_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[0] ));
 sg13g2_dfrbp_1 _14421_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1978),
    .D(net2149),
    .Q_N(_00137_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[1] ));
 sg13g2_dfrbp_1 _14422_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1978),
    .D(net2289),
    .Q_N(_00136_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[2] ));
 sg13g2_dfrbp_1 _14423_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1980),
    .D(_00415_),
    .Q_N(_00135_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[3] ));
 sg13g2_dfrbp_1 _14424_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1978),
    .D(_00416_),
    .Q_N(_00134_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[4] ));
 sg13g2_dfrbp_1 _14425_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1980),
    .D(net2303),
    .Q_N(_00133_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[5] ));
 sg13g2_dfrbp_1 _14426_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1983),
    .D(_00418_),
    .Q_N(_00132_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[6] ));
 sg13g2_dfrbp_1 _14427_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1983),
    .D(_00419_),
    .Q_N(_00131_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[7] ));
 sg13g2_dfrbp_1 _14428_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1980),
    .D(_00420_),
    .Q_N(_00130_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[8] ));
 sg13g2_dfrbp_1 _14429_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1982),
    .D(net2255),
    .Q_N(_00129_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[9] ));
 sg13g2_dfrbp_1 _14430_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1982),
    .D(_00422_),
    .Q_N(_00128_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[10] ));
 sg13g2_dfrbp_1 _14431_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1982),
    .D(net2222),
    .Q_N(_00127_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[11] ));
 sg13g2_dfrbp_1 _14432_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1982),
    .D(_00424_),
    .Q_N(_00126_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[12] ));
 sg13g2_dfrbp_1 _14433_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1978),
    .D(_00425_),
    .Q_N(_00176_),
    .Q(\vgadonut.donut.donuthit.cordicxy.x2in[13] ));
 sg13g2_dfrbp_1 _14434_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1978),
    .D(_00426_),
    .Q_N(_06997_),
    .Q(\vgadonut.donut.cB[0] ));
 sg13g2_dfrbp_1 _14435_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1979),
    .D(_00427_),
    .Q_N(_06996_),
    .Q(\vgadonut.donut.cB[1] ));
 sg13g2_dfrbp_1 _14436_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1980),
    .D(_00428_),
    .Q_N(_06995_),
    .Q(\vgadonut.donut.cB[2] ));
 sg13g2_dfrbp_1 _14437_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1980),
    .D(_00429_),
    .Q_N(_06994_),
    .Q(\vgadonut.donut.cB[3] ));
 sg13g2_dfrbp_1 _14438_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1980),
    .D(_00430_),
    .Q_N(_00115_),
    .Q(\vgadonut.donut.cB[4] ));
 sg13g2_dfrbp_1 _14439_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1981),
    .D(_00431_),
    .Q_N(_00116_),
    .Q(\vgadonut.donut.cB[5] ));
 sg13g2_dfrbp_1 _14440_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1981),
    .D(_00432_),
    .Q_N(_00117_),
    .Q(\vgadonut.donut.cB[6] ));
 sg13g2_dfrbp_1 _14441_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1982),
    .D(_00433_),
    .Q_N(_00118_),
    .Q(\vgadonut.donut.cB[7] ));
 sg13g2_dfrbp_1 _14442_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1981),
    .D(_00434_),
    .Q_N(_00119_),
    .Q(\vgadonut.donut.cB[8] ));
 sg13g2_dfrbp_1 _14443_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1981),
    .D(_00435_),
    .Q_N(_00120_),
    .Q(\vgadonut.donut.cB[9] ));
 sg13g2_dfrbp_1 _14444_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1981),
    .D(_00436_),
    .Q_N(_00121_),
    .Q(\vgadonut.donut.cB[10] ));
 sg13g2_dfrbp_1 _14445_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1981),
    .D(_00437_),
    .Q_N(_00122_),
    .Q(\vgadonut.donut.cB[11] ));
 sg13g2_dfrbp_1 _14446_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1981),
    .D(_00438_),
    .Q_N(_00123_),
    .Q(\vgadonut.donut.cB[12] ));
 sg13g2_dfrbp_1 _14447_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1981),
    .D(_00439_),
    .Q_N(_00124_),
    .Q(\vgadonut.donut.cB[13] ));
 sg13g2_dfrbp_1 _14448_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1982),
    .D(_00440_),
    .Q_N(\vgadonut.donut.cB[14] ),
    .Q(_00202_));
 sg13g2_dfrbp_1 _14449_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1982),
    .D(_00441_),
    .Q_N(_00125_),
    .Q(\vgadonut.donut.cB[15] ));
 sg13g2_dfrbp_1 _14450_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net87),
    .D(_00442_),
    .Q_N(_06993_),
    .Q(\vgadonut.donut.donut_visible ));
 sg13g2_dfrbp_1 _14451_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1970),
    .D(net1462),
    .Q_N(\vgadonut.donut.sA[0] ),
    .Q(_00203_));
 sg13g2_dfrbp_1 _14452_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1970),
    .D(net1467),
    .Q_N(\vgadonut.donut.sA[1] ),
    .Q(_00204_));
 sg13g2_dfrbp_1 _14453_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1970),
    .D(net1460),
    .Q_N(\vgadonut.donut.sA[2] ),
    .Q(_00205_));
 sg13g2_dfrbp_1 _14454_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1960),
    .D(_00446_),
    .Q_N(\vgadonut.donut.sA[3] ),
    .Q(_00206_));
 sg13g2_dfrbp_1 _14455_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1969),
    .D(_00447_),
    .Q_N(\vgadonut.donut.sA[4] ),
    .Q(_00207_));
 sg13g2_dfrbp_1 _14456_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1969),
    .D(_00448_),
    .Q_N(\vgadonut.donut.sA[5] ),
    .Q(_00208_));
 sg13g2_dfrbp_1 _14457_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1967),
    .D(_00449_),
    .Q_N(_06992_),
    .Q(\vgadonut.donut.sA[6] ));
 sg13g2_dfrbp_1 _14458_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1967),
    .D(_00450_),
    .Q_N(_06991_),
    .Q(\vgadonut.donut.sA[7] ));
 sg13g2_dfrbp_1 _14459_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1967),
    .D(_00451_),
    .Q_N(\vgadonut.donut.sA[8] ),
    .Q(_00209_));
 sg13g2_dfrbp_1 _14460_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1967),
    .D(_00452_),
    .Q_N(_06990_),
    .Q(\vgadonut.donut.sA[9] ));
 sg13g2_dfrbp_1 _14461_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1968),
    .D(_00453_),
    .Q_N(\vgadonut.donut.sA[10] ),
    .Q(_00210_));
 sg13g2_dfrbp_1 _14462_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1967),
    .D(_00454_),
    .Q_N(\vgadonut.donut.sA[11] ),
    .Q(_00211_));
 sg13g2_dfrbp_1 _14463_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1971),
    .D(_00455_),
    .Q_N(_06989_),
    .Q(\vgadonut.donut.sA[12] ));
 sg13g2_dfrbp_1 _14464_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1967),
    .D(_00456_),
    .Q_N(\vgadonut.donut.sA[13] ),
    .Q(_00212_));
 sg13g2_dfrbp_1 _14465_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1972),
    .D(net2312),
    .Q_N(_00141_),
    .Q(\vgadonut.donut.sA[14] ));
 sg13g2_dfrbp_1 _14466_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1968),
    .D(_00458_),
    .Q_N(_06988_),
    .Q(\vgadonut.donut.sA[15] ));
 sg13g2_dfrbp_1 _14467_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1958),
    .D(net1484),
    .Q_N(\vgadonut.donut.cA[0] ),
    .Q(_00213_));
 sg13g2_dfrbp_1 _14468_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1958),
    .D(_00460_),
    .Q_N(\vgadonut.donut.cA[1] ),
    .Q(_00214_));
 sg13g2_dfrbp_1 _14469_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1958),
    .D(_00461_),
    .Q_N(\vgadonut.donut.cA[2] ),
    .Q(_00215_));
 sg13g2_dfrbp_1 _14470_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1958),
    .D(_00462_),
    .Q_N(\vgadonut.donut.cA[3] ),
    .Q(_00216_));
 sg13g2_dfrbp_1 _14471_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1958),
    .D(_00463_),
    .Q_N(\vgadonut.donut.cA[4] ),
    .Q(_00217_));
 sg13g2_dfrbp_1 _14472_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1960),
    .D(_00464_),
    .Q_N(\vgadonut.donut.cA[5] ),
    .Q(_00218_));
 sg13g2_dfrbp_1 _14473_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1959),
    .D(_00465_),
    .Q_N(_06987_),
    .Q(\vgadonut.donut.cA[6] ));
 sg13g2_dfrbp_1 _14474_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1969),
    .D(_00466_),
    .Q_N(_06986_),
    .Q(\vgadonut.donut.cA[7] ));
 sg13g2_dfrbp_1 _14475_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1969),
    .D(_00467_),
    .Q_N(\vgadonut.donut.cA[8] ),
    .Q(_00219_));
 sg13g2_dfrbp_1 _14476_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1970),
    .D(_00468_),
    .Q_N(_06985_),
    .Q(\vgadonut.donut.cA[9] ));
 sg13g2_dfrbp_1 _14477_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1970),
    .D(_00469_),
    .Q_N(\vgadonut.donut.cA[10] ),
    .Q(_00220_));
 sg13g2_dfrbp_1 _14478_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1970),
    .D(_00470_),
    .Q_N(\vgadonut.donut.cA[11] ),
    .Q(_00221_));
 sg13g2_dfrbp_1 _14479_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1968),
    .D(_00471_),
    .Q_N(_06984_),
    .Q(\vgadonut.donut.cA[12] ));
 sg13g2_dfrbp_1 _14480_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1967),
    .D(_00472_),
    .Q_N(\vgadonut.donut.cA[13] ),
    .Q(_00222_));
 sg13g2_dfrbp_1 _14481_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1967),
    .D(_00473_),
    .Q_N(_06983_),
    .Q(\vgadonut.donut.cA[14] ));
 sg13g2_dfrbp_1 _14482_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1968),
    .D(_00474_),
    .Q_N(_06982_),
    .Q(\vgadonut.donut.cA[15] ));
 sg13g2_dfrbp_1 _14483_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net161),
    .D(_00475_),
    .Q_N(_00170_),
    .Q(_00031_));
 sg13g2_dfrbp_1 _14484_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net163),
    .D(_00476_),
    .Q_N(_07150_),
    .Q(\vgadonut.donut.donuthit.hit ));
 sg13g2_dfrbp_1 _14485_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net164),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[8] ),
    .Q_N(_07151_),
    .Q(\vgadonut.donut.donuthit.light[8] ));
 sg13g2_dfrbp_1 _14486_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net165),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[9] ),
    .Q_N(_07152_),
    .Q(\vgadonut.donut.donuthit.light[9] ));
 sg13g2_dfrbp_1 _14487_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net166),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[10] ),
    .Q_N(_07153_),
    .Q(\vgadonut.donut.donuthit.light[10] ));
 sg13g2_dfrbp_1 _14488_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net167),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[11] ),
    .Q_N(_07154_),
    .Q(\vgadonut.donut.donuthit.light[11] ));
 sg13g2_dfrbp_1 _14489_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net179),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[12] ),
    .Q_N(_07155_),
    .Q(\vgadonut.donut.donuthit.light[12] ));
 sg13g2_dfrbp_1 _14490_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net160),
    .D(\vgadonut.donut.donuthit.cordicxz.x2out[13] ),
    .Q_N(_00045_),
    .Q(\vgadonut.donut.donuthit.light[13] ));
 sg13g2_dfrbp_1 _14491_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net159),
    .D(net2016),
    .Q_N(_06981_),
    .Q(\vgadonut.donut.rz6[0] ));
 sg13g2_dfrbp_1 _14492_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net158),
    .D(net2000),
    .Q_N(_06980_),
    .Q(\vgadonut.donut.rz6[1] ));
 sg13g2_dfrbp_1 _14493_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net157),
    .D(_00479_),
    .Q_N(_06979_),
    .Q(\vgadonut.donut.rz6[2] ));
 sg13g2_dfrbp_1 _14494_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net156),
    .D(_00480_),
    .Q_N(_06978_),
    .Q(\vgadonut.donut.rz6[3] ));
 sg13g2_dfrbp_1 _14495_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net155),
    .D(_00481_),
    .Q_N(_06977_),
    .Q(\vgadonut.donut.rz6[4] ));
 sg13g2_dfrbp_1 _14496_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net154),
    .D(_00482_),
    .Q_N(_06976_),
    .Q(\vgadonut.donut.rz6[5] ));
 sg13g2_dfrbp_1 _14497_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net153),
    .D(_00483_),
    .Q_N(_06975_),
    .Q(\vgadonut.donut.donuthit.rzin[0] ));
 sg13g2_dfrbp_1 _14498_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net152),
    .D(_00484_),
    .Q_N(_06974_),
    .Q(\vgadonut.donut.donuthit.rzin[1] ));
 sg13g2_dfrbp_1 _14499_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net151),
    .D(_00485_),
    .Q_N(_06973_),
    .Q(\vgadonut.donut.donuthit.rzin[2] ));
 sg13g2_dfrbp_1 _14500_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net150),
    .D(_00486_),
    .Q_N(_06972_),
    .Q(\vgadonut.donut.donuthit.rzin[3] ));
 sg13g2_dfrbp_1 _14501_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net149),
    .D(_00487_),
    .Q_N(_06971_),
    .Q(\vgadonut.donut.donuthit.rzin[4] ));
 sg13g2_dfrbp_1 _14502_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net148),
    .D(_00488_),
    .Q_N(_06970_),
    .Q(\vgadonut.donut.donuthit.rzin[5] ));
 sg13g2_dfrbp_1 _14503_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net147),
    .D(_00489_),
    .Q_N(_06969_),
    .Q(\vgadonut.donut.donuthit.rzin[6] ));
 sg13g2_dfrbp_1 _14504_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net146),
    .D(_00490_),
    .Q_N(_06968_),
    .Q(\vgadonut.donut.donuthit.rzin[7] ));
 sg13g2_dfrbp_1 _14505_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net145),
    .D(_00491_),
    .Q_N(_06967_),
    .Q(\vgadonut.donut.donuthit.rzin[8] ));
 sg13g2_dfrbp_1 _14506_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net144),
    .D(_00492_),
    .Q_N(_06966_),
    .Q(\vgadonut.donut.donuthit.rzin[9] ));
 sg13g2_dfrbp_1 _14507_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net143),
    .D(_00493_),
    .Q_N(_06965_),
    .Q(\vgadonut.donut.donuthit.rzin[10] ));
 sg13g2_dfrbp_1 _14508_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net142),
    .D(_00494_),
    .Q_N(_06964_),
    .Q(\vgadonut.donut.donuthit.rzin[11] ));
 sg13g2_dfrbp_1 _14509_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net141),
    .D(_00495_),
    .Q_N(_06963_),
    .Q(\vgadonut.donut.donuthit.rzin[12] ));
 sg13g2_dfrbp_1 _14510_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net140),
    .D(_00496_),
    .Q_N(_06962_),
    .Q(\vgadonut.donut.donuthit.rzin[13] ));
 sg13g2_dfrbp_1 _14511_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net139),
    .D(_00497_),
    .Q_N(_06961_),
    .Q(\vgadonut.donut.donuthit.rzin[14] ));
 sg13g2_dfrbp_1 _14512_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net180),
    .D(_00498_),
    .Q_N(_00169_),
    .Q(\vgadonut.donut.donuthit.rzin[15] ));
 sg13g2_dfrbp_1 _14513_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net181),
    .D(_00078_),
    .Q_N(_00154_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[0] ));
 sg13g2_dfrbp_1 _14514_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net182),
    .D(_00085_),
    .Q_N(_00153_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[1] ));
 sg13g2_dfrbp_1 _14515_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net183),
    .D(_00086_),
    .Q_N(_00152_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[2] ));
 sg13g2_dfrbp_1 _14516_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net184),
    .D(_00087_),
    .Q_N(_00151_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[3] ));
 sg13g2_dfrbp_1 _14517_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net185),
    .D(_00088_),
    .Q_N(_00150_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[4] ));
 sg13g2_dfrbp_1 _14518_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net186),
    .D(_00089_),
    .Q_N(_00149_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[5] ));
 sg13g2_dfrbp_1 _14519_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net187),
    .D(_00090_),
    .Q_N(_00148_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[6] ));
 sg13g2_dfrbp_1 _14520_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net188),
    .D(_00091_),
    .Q_N(_00147_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[7] ));
 sg13g2_dfrbp_1 _14521_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net189),
    .D(_00092_),
    .Q_N(_00146_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[8] ));
 sg13g2_dfrbp_1 _14522_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net190),
    .D(_00093_),
    .Q_N(_00145_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[9] ));
 sg13g2_dfrbp_1 _14523_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net191),
    .D(_00079_),
    .Q_N(_00144_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[10] ));
 sg13g2_dfrbp_1 _14524_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net192),
    .D(_00080_),
    .Q_N(_00143_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[11] ));
 sg13g2_dfrbp_1 _14525_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net193),
    .D(_00081_),
    .Q_N(_00155_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[12] ));
 sg13g2_dfrbp_1 _14526_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net194),
    .D(_00082_),
    .Q_N(_00157_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[13] ));
 sg13g2_dfrbp_1 _14527_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net195),
    .D(_00083_),
    .Q_N(_00158_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[14] ));
 sg13g2_dfrbp_1 _14528_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net196),
    .D(_00084_),
    .Q_N(_00156_),
    .Q(\vgadonut.donut.donuthit.cordicxz.xin[15] ));
 sg13g2_dfrbp_1 _14529_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net197),
    .D(net2339),
    .Q_N(_07156_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[0] ));
 sg13g2_dfrbp_1 _14530_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net198),
    .D(_00069_),
    .Q_N(_07157_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[1] ));
 sg13g2_dfrbp_1 _14531_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net199),
    .D(_00070_),
    .Q_N(_07158_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[2] ));
 sg13g2_dfrbp_1 _14532_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net200),
    .D(_00071_),
    .Q_N(_07159_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[3] ));
 sg13g2_dfrbp_1 _14533_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net201),
    .D(_00072_),
    .Q_N(_07160_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[4] ));
 sg13g2_dfrbp_1 _14534_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net202),
    .D(_00073_),
    .Q_N(_07161_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[5] ));
 sg13g2_dfrbp_1 _14535_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net203),
    .D(_00074_),
    .Q_N(_07162_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[6] ));
 sg13g2_dfrbp_1 _14536_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net204),
    .D(_00075_),
    .Q_N(_07163_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[7] ));
 sg13g2_dfrbp_1 _14537_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net205),
    .D(_00076_),
    .Q_N(_07164_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[8] ));
 sg13g2_dfrbp_1 _14538_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net206),
    .D(_00077_),
    .Q_N(_07165_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[9] ));
 sg13g2_dfrbp_1 _14539_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net207),
    .D(_00063_),
    .Q_N(_07166_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[10] ));
 sg13g2_dfrbp_1 _14540_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net208),
    .D(_00064_),
    .Q_N(_00164_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[11] ));
 sg13g2_dfrbp_1 _14541_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net209),
    .D(_00065_),
    .Q_N(_00166_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[12] ));
 sg13g2_dfrbp_1 _14542_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net210),
    .D(_00066_),
    .Q_N(_00167_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[13] ));
 sg13g2_dfrbp_1 _14543_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net211),
    .D(_00067_),
    .Q_N(_00168_),
    .Q(\vgadonut.donut.donuthit.cordicxy.yin[14] ));
 sg13g2_dfrbp_1 _14544_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net212),
    .D(_00068_),
    .Q_N(_00142_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xinvert ));
 sg13g2_dfrbp_1 _14545_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net213),
    .D(_00046_),
    .Q_N(_07167_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[0] ));
 sg13g2_dfrbp_1 _14546_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net214),
    .D(_00053_),
    .Q_N(_07168_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[1] ));
 sg13g2_dfrbp_1 _14547_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net215),
    .D(_00054_),
    .Q_N(_07169_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[2] ));
 sg13g2_dfrbp_1 _14548_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net216),
    .D(_00055_),
    .Q_N(_07170_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[3] ));
 sg13g2_dfrbp_1 _14549_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net217),
    .D(_00056_),
    .Q_N(_07171_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[4] ));
 sg13g2_dfrbp_1 _14550_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net218),
    .D(_00057_),
    .Q_N(_07172_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[5] ));
 sg13g2_dfrbp_1 _14551_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net219),
    .D(_00058_),
    .Q_N(_07173_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[6] ));
 sg13g2_dfrbp_1 _14552_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net220),
    .D(_00059_),
    .Q_N(_07174_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[7] ));
 sg13g2_dfrbp_1 _14553_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net221),
    .D(_00060_),
    .Q_N(_07175_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[8] ));
 sg13g2_dfrbp_1 _14554_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net222),
    .D(_00061_),
    .Q_N(_07176_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[9] ));
 sg13g2_dfrbp_1 _14555_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net223),
    .D(_00047_),
    .Q_N(_07177_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[10] ));
 sg13g2_dfrbp_1 _14556_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net224),
    .D(_00048_),
    .Q_N(_00159_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[11] ));
 sg13g2_dfrbp_1 _14557_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net225),
    .D(_00049_),
    .Q_N(_00161_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[12] ));
 sg13g2_dfrbp_1 _14558_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net226),
    .D(_00050_),
    .Q_N(_00162_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[13] ));
 sg13g2_dfrbp_1 _14559_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net257),
    .D(_00051_),
    .Q_N(_00163_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[14] ));
 sg13g2_dfrbp_1 _14560_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net138),
    .D(_00052_),
    .Q_N(_06960_),
    .Q(\vgadonut.donut.donuthit.cordicxy.xin[15] ));
 sg13g2_dfrbp_1 _14561_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net137),
    .D(net2157),
    .Q_N(_06959_),
    .Q(\vgadonut.donut.donuthit.rx[5] ));
 sg13g2_dfrbp_1 _14562_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net136),
    .D(net2105),
    .Q_N(_06958_),
    .Q(\vgadonut.donut.donuthit.rx[6] ));
 sg13g2_dfrbp_1 _14563_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net135),
    .D(net2111),
    .Q_N(_06957_),
    .Q(\vgadonut.donut.donuthit.rx[7] ));
 sg13g2_dfrbp_1 _14564_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net134),
    .D(net2072),
    .Q_N(_06956_),
    .Q(\vgadonut.donut.donuthit.rx[8] ));
 sg13g2_dfrbp_1 _14565_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net133),
    .D(net2093),
    .Q_N(_06955_),
    .Q(\vgadonut.donut.donuthit.rx[9] ));
 sg13g2_dfrbp_1 _14566_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net132),
    .D(net2123),
    .Q_N(_06954_),
    .Q(\vgadonut.donut.donuthit.rx[10] ));
 sg13g2_dfrbp_1 _14567_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net89),
    .D(net2121),
    .Q_N(_06953_),
    .Q(\vgadonut.donut.donuthit.rx[11] ));
 sg13g2_dfrbp_1 _14568_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net88),
    .D(net2199),
    .Q_N(_06952_),
    .Q(\vgadonut.donut.donuthit.rx[12] ));
 sg13g2_dfrbp_1 _14569_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net86),
    .D(net2193),
    .Q_N(_06951_),
    .Q(\vgadonut.donut.donuthit.rx[13] ));
 sg13g2_dfrbp_1 _14570_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net85),
    .D(net2204),
    .Q_N(_06950_),
    .Q(\vgadonut.donut.donuthit.rx[14] ));
 sg13g2_dfrbp_1 _14571_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net84),
    .D(net2145),
    .Q_N(_06949_),
    .Q(\vgadonut.donut.donuthit.rx[15] ));
 sg13g2_dfrbp_1 _14572_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net83),
    .D(net2163),
    .Q_N(_06948_),
    .Q(\vgadonut.donut.donuthit.ry[5] ));
 sg13g2_dfrbp_1 _14573_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net82),
    .D(net2042),
    .Q_N(_06947_),
    .Q(\vgadonut.donut.donuthit.ry[6] ));
 sg13g2_dfrbp_1 _14574_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net81),
    .D(net2135),
    .Q_N(_06946_),
    .Q(\vgadonut.donut.donuthit.ry[7] ));
 sg13g2_dfrbp_1 _14575_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net80),
    .D(net2052),
    .Q_N(_06945_),
    .Q(\vgadonut.donut.donuthit.ry[8] ));
 sg13g2_dfrbp_1 _14576_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net79),
    .D(net2088),
    .Q_N(_06944_),
    .Q(\vgadonut.donut.donuthit.ry[9] ));
 sg13g2_dfrbp_1 _14577_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net78),
    .D(net2050),
    .Q_N(_06943_),
    .Q(\vgadonut.donut.donuthit.ry[10] ));
 sg13g2_dfrbp_1 _14578_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net77),
    .D(net2057),
    .Q_N(_06942_),
    .Q(\vgadonut.donut.donuthit.ry[11] ));
 sg13g2_dfrbp_1 _14579_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net76),
    .D(net2021),
    .Q_N(_06941_),
    .Q(\vgadonut.donut.donuthit.ry[12] ));
 sg13g2_dfrbp_1 _14580_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net75),
    .D(net2036),
    .Q_N(_06940_),
    .Q(\vgadonut.donut.donuthit.ry[13] ));
 sg13g2_dfrbp_1 _14581_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net74),
    .D(net2129),
    .Q_N(_06939_),
    .Q(\vgadonut.donut.donuthit.ry[14] ));
 sg13g2_dfrbp_1 _14582_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net73),
    .D(net2117),
    .Q_N(_06938_),
    .Q(\vgadonut.donut.donuthit.ry[15] ));
 sg13g2_dfrbp_1 _14583_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net72),
    .D(net2101),
    .Q_N(_06937_),
    .Q(\vgadonut.donut.donuthit.rz[5] ));
 sg13g2_dfrbp_1 _14584_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net71),
    .D(_00522_),
    .Q_N(_06936_),
    .Q(\vgadonut.donut.donuthit.rz[6] ));
 sg13g2_dfrbp_1 _14585_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net70),
    .D(net2115),
    .Q_N(_06935_),
    .Q(\vgadonut.donut.donuthit.rz[7] ));
 sg13g2_dfrbp_1 _14586_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net69),
    .D(net2068),
    .Q_N(_06934_),
    .Q(\vgadonut.donut.donuthit.rz[8] ));
 sg13g2_dfrbp_1 _14587_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net68),
    .D(net2047),
    .Q_N(_06933_),
    .Q(\vgadonut.donut.donuthit.rz[9] ));
 sg13g2_dfrbp_1 _14588_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net67),
    .D(net2055),
    .Q_N(_06932_),
    .Q(\vgadonut.donut.donuthit.rz[10] ));
 sg13g2_dfrbp_1 _14589_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net66),
    .D(net2132),
    .Q_N(_06931_),
    .Q(\vgadonut.donut.donuthit.rz[11] ));
 sg13g2_dfrbp_1 _14590_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net65),
    .D(net2024),
    .Q_N(_06930_),
    .Q(\vgadonut.donut.donuthit.rz[12] ));
 sg13g2_dfrbp_1 _14591_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net64),
    .D(net2139),
    .Q_N(_06929_),
    .Q(\vgadonut.donut.donuthit.rz[13] ));
 sg13g2_dfrbp_1 _14592_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net63),
    .D(net2075),
    .Q_N(_06928_),
    .Q(\vgadonut.donut.donuthit.rz[14] ));
 sg13g2_dfrbp_1 _14593_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net62),
    .D(net2030),
    .Q_N(_06927_),
    .Q(\vgadonut.donut.donuthit.rz[15] ));
 sg13g2_dfrbp_1 _14594_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net61),
    .D(_00532_),
    .Q_N(_06926_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _14595_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net258),
    .D(_00533_),
    .Q_N(_07178_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _14596_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1974),
    .D(_00014_),
    .Q_N(_07179_),
    .Q(\vgadonut.donut.h_count[0] ));
 sg13g2_dfrbp_1 _14597_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1974),
    .D(net2003),
    .Q_N(_07180_),
    .Q(\vgadonut.donut.h_count[1] ));
 sg13g2_dfrbp_1 _14598_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1974),
    .D(_00017_),
    .Q_N(_00177_),
    .Q(\vgadonut.donut.h_count[2] ));
 sg13g2_dfrbp_1 _14599_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1974),
    .D(_00018_),
    .Q_N(_00178_),
    .Q(\vgadonut.donut.h_count[3] ));
 sg13g2_dfrbp_1 _14600_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1971),
    .D(_00019_),
    .Q_N(_07181_),
    .Q(\vgadonut.donut.h_count[4] ));
 sg13g2_dfrbp_1 _14601_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1971),
    .D(_00020_),
    .Q_N(_07182_),
    .Q(\vgadonut.donut.h_count[5] ));
 sg13g2_dfrbp_1 _14602_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1971),
    .D(_00021_),
    .Q_N(_07183_),
    .Q(\vgadonut.donut.h_count[6] ));
 sg13g2_dfrbp_1 _14603_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1971),
    .D(_00022_),
    .Q_N(_07184_),
    .Q(\vgadonut.donut.h_count[7] ));
 sg13g2_dfrbp_1 _14604_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1971),
    .D(_00023_),
    .Q_N(_07185_),
    .Q(\vgadonut.donut.h_count[8] ));
 sg13g2_dfrbp_1 _14605_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1971),
    .D(net2063),
    .Q_N(_07186_),
    .Q(\vgadonut.donut.h_count[9] ));
 sg13g2_dfrbp_1 _14606_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1972),
    .D(net1446),
    .Q_N(_00179_),
    .Q(\vgadonut.donut.h_count[10] ));
 sg13g2_dfrbp_1 _14607_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net60),
    .D(_00534_),
    .Q_N(_06925_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _14608_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net59),
    .D(_00535_),
    .Q_N(_06924_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _14609_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net58),
    .D(_00536_),
    .Q_N(_06923_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _14610_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net263),
    .D(_00537_),
    .Q_N(_07187_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _14611_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net168),
    .D(net2219),
    .Q_N(_07188_),
    .Q(\vgadonut.vsync ));
 sg13g2_dfrbp_1 _14612_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net57),
    .D(net2078),
    .Q_N(_06922_),
    .Q(hsync));
 sg13g2_dfrbp_1 _14613_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net55),
    .D(net1448),
    .Q_N(_00181_),
    .Q(\vgadonut.donut.frame ));
 sg13g2_dfrbp_1 _14614_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net234),
    .D(net2034),
    .Q_N(_06921_),
    .Q(\vgadonut.frame[1] ));
 sg13g2_dfrbp_1 _14615_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net231),
    .D(net2083),
    .Q_N(_06920_),
    .Q(\vgadonut.frame[2] ));
 sg13g2_dfrbp_1 _14616_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net227),
    .D(_00541_),
    .Q_N(_06919_),
    .Q(\vgadonut.frame[3] ));
 sg13g2_dfrbp_1 _14617_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net172),
    .D(_00542_),
    .Q_N(_06918_),
    .Q(\vgadonut.frame[4] ));
 sg13g2_dfrbp_1 _14618_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net171),
    .D(_00543_),
    .Q_N(_06917_),
    .Q(\vgadonut.frame[5] ));
 sg13g2_dfrbp_1 _14619_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net170),
    .D(net2090),
    .Q_N(_06916_),
    .Q(\vgadonut.frame[6] ));
 sg13g2_dfrbp_1 _14620_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net169),
    .D(net2045),
    .Q_N(_06915_),
    .Q(\vgadonut.frame[7] ));
 sg13g2_tiehi _14255__18 (.L_HI(net18));
 sg13g2_tiehi _14217__19 (.L_HI(net19));
 sg13g2_tiehi _14218__20 (.L_HI(net20));
 sg13g2_tiehi _14219__21 (.L_HI(net21));
 sg13g2_tiehi _14220__22 (.L_HI(net22));
 sg13g2_tiehi _14221__23 (.L_HI(net23));
 sg13g2_tiehi _14222__24 (.L_HI(net24));
 sg13g2_tiehi _14223__25 (.L_HI(net25));
 sg13g2_tiehi _14224__26 (.L_HI(net26));
 sg13g2_tiehi _14225__27 (.L_HI(net27));
 sg13g2_tiehi _14226__28 (.L_HI(net28));
 sg13g2_tiehi _14227__29 (.L_HI(net29));
 sg13g2_tiehi _14228__30 (.L_HI(net30));
 sg13g2_tiehi _14229__31 (.L_HI(net31));
 sg13g2_tiehi _14230__32 (.L_HI(net32));
 sg13g2_tiehi _14254__33 (.L_HI(net33));
 sg13g2_tiehi _14253__34 (.L_HI(net34));
 sg13g2_tiehi _14252__35 (.L_HI(net35));
 sg13g2_tiehi _14251__36 (.L_HI(net36));
 sg13g2_tiehi _14250__37 (.L_HI(net37));
 sg13g2_tiehi _14249__38 (.L_HI(net38));
 sg13g2_tiehi _14248__39 (.L_HI(net39));
 sg13g2_tiehi _14247__40 (.L_HI(net40));
 sg13g2_tiehi _14246__41 (.L_HI(net41));
 sg13g2_tiehi _14245__42 (.L_HI(net42));
 sg13g2_tiehi _14244__43 (.L_HI(net43));
 sg13g2_tiehi _14243__44 (.L_HI(net44));
 sg13g2_tiehi _14242__45 (.L_HI(net45));
 sg13g2_tiehi _14241__46 (.L_HI(net46));
 sg13g2_tiehi _14240__47 (.L_HI(net47));
 sg13g2_tiehi _14239__48 (.L_HI(net48));
 sg13g2_tiehi _14238__49 (.L_HI(net49));
 sg13g2_tiehi _14237__50 (.L_HI(net50));
 sg13g2_tiehi _14236__51 (.L_HI(net51));
 sg13g2_tiehi _14235__52 (.L_HI(net52));
 sg13g2_tiehi _14234__53 (.L_HI(net53));
 sg13g2_tiehi _14233__54 (.L_HI(net54));
 sg13g2_tiehi _14613__55 (.L_HI(net55));
 sg13g2_tiehi _14232__56 (.L_HI(net56));
 sg13g2_tiehi _14612__57 (.L_HI(net57));
 sg13g2_tiehi _14609__58 (.L_HI(net58));
 sg13g2_tiehi _14608__59 (.L_HI(net59));
 sg13g2_tiehi _14607__60 (.L_HI(net60));
 sg13g2_tiehi _14594__61 (.L_HI(net61));
 sg13g2_tiehi _14593__62 (.L_HI(net62));
 sg13g2_tiehi _14592__63 (.L_HI(net63));
 sg13g2_tiehi _14591__64 (.L_HI(net64));
 sg13g2_tiehi _14590__65 (.L_HI(net65));
 sg13g2_tiehi _14589__66 (.L_HI(net66));
 sg13g2_tiehi _14588__67 (.L_HI(net67));
 sg13g2_tiehi _14587__68 (.L_HI(net68));
 sg13g2_tiehi _14586__69 (.L_HI(net69));
 sg13g2_tiehi _14585__70 (.L_HI(net70));
 sg13g2_tiehi _14584__71 (.L_HI(net71));
 sg13g2_tiehi _14583__72 (.L_HI(net72));
 sg13g2_tiehi _14582__73 (.L_HI(net73));
 sg13g2_tiehi _14581__74 (.L_HI(net74));
 sg13g2_tiehi _14580__75 (.L_HI(net75));
 sg13g2_tiehi _14579__76 (.L_HI(net76));
 sg13g2_tiehi _14578__77 (.L_HI(net77));
 sg13g2_tiehi _14577__78 (.L_HI(net78));
 sg13g2_tiehi _14576__79 (.L_HI(net79));
 sg13g2_tiehi _14575__80 (.L_HI(net80));
 sg13g2_tiehi _14574__81 (.L_HI(net81));
 sg13g2_tiehi _14573__82 (.L_HI(net82));
 sg13g2_tiehi _14572__83 (.L_HI(net83));
 sg13g2_tiehi _14571__84 (.L_HI(net84));
 sg13g2_tiehi _14570__85 (.L_HI(net85));
 sg13g2_tiehi _14569__86 (.L_HI(net86));
 sg13g2_tiehi _14450__87 (.L_HI(net87));
 sg13g2_tiehi _14568__88 (.L_HI(net88));
 sg13g2_tiehi _14567__89 (.L_HI(net89));
 sg13g2_tiehi _14417__90 (.L_HI(net90));
 sg13g2_tiehi _14416__91 (.L_HI(net91));
 sg13g2_tiehi _14415__92 (.L_HI(net92));
 sg13g2_tiehi _14414__93 (.L_HI(net93));
 sg13g2_tiehi _14413__94 (.L_HI(net94));
 sg13g2_tiehi _14412__95 (.L_HI(net95));
 sg13g2_tiehi _14411__96 (.L_HI(net96));
 sg13g2_tiehi _14410__97 (.L_HI(net97));
 sg13g2_tiehi _14409__98 (.L_HI(net98));
 sg13g2_tiehi _14408__99 (.L_HI(net99));
 sg13g2_tiehi _14407__100 (.L_HI(net100));
 sg13g2_tiehi _14406__101 (.L_HI(net101));
 sg13g2_tiehi _14405__102 (.L_HI(net102));
 sg13g2_tiehi _14404__103 (.L_HI(net103));
 sg13g2_tiehi _14403__104 (.L_HI(net104));
 sg13g2_tiehi _14402__105 (.L_HI(net105));
 sg13g2_tiehi _14401__106 (.L_HI(net106));
 sg13g2_tiehi _14400__107 (.L_HI(net107));
 sg13g2_tiehi _14399__108 (.L_HI(net108));
 sg13g2_tiehi _14398__109 (.L_HI(net109));
 sg13g2_tiehi _14397__110 (.L_HI(net110));
 sg13g2_tiehi _14396__111 (.L_HI(net111));
 sg13g2_tiehi _14395__112 (.L_HI(net112));
 sg13g2_tiehi _14394__113 (.L_HI(net113));
 sg13g2_tiehi _14393__114 (.L_HI(net114));
 sg13g2_tiehi _14392__115 (.L_HI(net115));
 sg13g2_tiehi _14391__116 (.L_HI(net116));
 sg13g2_tiehi _14390__117 (.L_HI(net117));
 sg13g2_tiehi _14389__118 (.L_HI(net118));
 sg13g2_tiehi _14388__119 (.L_HI(net119));
 sg13g2_tiehi _14387__120 (.L_HI(net120));
 sg13g2_tiehi _14386__121 (.L_HI(net121));
 sg13g2_tiehi _14385__122 (.L_HI(net122));
 sg13g2_tiehi _14384__123 (.L_HI(net123));
 sg13g2_tiehi _14383__124 (.L_HI(net124));
 sg13g2_tiehi _14382__125 (.L_HI(net125));
 sg13g2_tiehi _14381__126 (.L_HI(net126));
 sg13g2_tiehi _14380__127 (.L_HI(net127));
 sg13g2_tiehi _14379__128 (.L_HI(net128));
 sg13g2_tiehi _14378__129 (.L_HI(net129));
 sg13g2_tiehi _14377__130 (.L_HI(net130));
 sg13g2_tiehi _14376__131 (.L_HI(net131));
 sg13g2_tiehi _14566__132 (.L_HI(net132));
 sg13g2_tiehi _14565__133 (.L_HI(net133));
 sg13g2_tiehi _14564__134 (.L_HI(net134));
 sg13g2_tiehi _14563__135 (.L_HI(net135));
 sg13g2_tiehi _14562__136 (.L_HI(net136));
 sg13g2_tiehi _14561__137 (.L_HI(net137));
 sg13g2_tiehi _14560__138 (.L_HI(net138));
 sg13g2_tiehi _14511__139 (.L_HI(net139));
 sg13g2_tiehi _14510__140 (.L_HI(net140));
 sg13g2_tiehi _14509__141 (.L_HI(net141));
 sg13g2_tiehi _14508__142 (.L_HI(net142));
 sg13g2_tiehi _14507__143 (.L_HI(net143));
 sg13g2_tiehi _14506__144 (.L_HI(net144));
 sg13g2_tiehi _14505__145 (.L_HI(net145));
 sg13g2_tiehi _14504__146 (.L_HI(net146));
 sg13g2_tiehi _14503__147 (.L_HI(net147));
 sg13g2_tiehi _14502__148 (.L_HI(net148));
 sg13g2_tiehi _14501__149 (.L_HI(net149));
 sg13g2_tiehi _14500__150 (.L_HI(net150));
 sg13g2_tiehi _14499__151 (.L_HI(net151));
 sg13g2_tiehi _14498__152 (.L_HI(net152));
 sg13g2_tiehi _14497__153 (.L_HI(net153));
 sg13g2_tiehi _14496__154 (.L_HI(net154));
 sg13g2_tiehi _14495__155 (.L_HI(net155));
 sg13g2_tiehi _14494__156 (.L_HI(net156));
 sg13g2_tiehi _14493__157 (.L_HI(net157));
 sg13g2_tiehi _14492__158 (.L_HI(net158));
 sg13g2_tiehi _14491__159 (.L_HI(net159));
 sg13g2_tiehi _14490__160 (.L_HI(net160));
 sg13g2_tiehi _14483__161 (.L_HI(net161));
 sg13g2_tiehi _14231__162 (.L_HI(net162));
 sg13g2_tiehi _14484__163 (.L_HI(net163));
 sg13g2_tiehi _14485__164 (.L_HI(net164));
 sg13g2_tiehi _14486__165 (.L_HI(net165));
 sg13g2_tiehi _14487__166 (.L_HI(net166));
 sg13g2_tiehi _14488__167 (.L_HI(net167));
 sg13g2_tiehi _14611__168 (.L_HI(net168));
 sg13g2_tiehi _14620__169 (.L_HI(net169));
 sg13g2_tiehi _14619__170 (.L_HI(net170));
 sg13g2_tiehi _14618__171 (.L_HI(net171));
 sg13g2_tiehi _14617__172 (.L_HI(net172));
 sg13g2_tiehi _14301__173 (.L_HI(net173));
 sg13g2_tiehi _14300__174 (.L_HI(net174));
 sg13g2_tiehi _14299__175 (.L_HI(net175));
 sg13g2_tiehi _14298__176 (.L_HI(net176));
 sg13g2_tiehi _14297__177 (.L_HI(net177));
 sg13g2_tiehi _14296__178 (.L_HI(net178));
 sg13g2_tiehi _14489__179 (.L_HI(net179));
 sg13g2_tiehi _14512__180 (.L_HI(net180));
 sg13g2_tiehi _14513__181 (.L_HI(net181));
 sg13g2_tiehi _14514__182 (.L_HI(net182));
 sg13g2_tiehi _14515__183 (.L_HI(net183));
 sg13g2_tiehi _14516__184 (.L_HI(net184));
 sg13g2_tiehi _14517__185 (.L_HI(net185));
 sg13g2_tiehi _14518__186 (.L_HI(net186));
 sg13g2_tiehi _14519__187 (.L_HI(net187));
 sg13g2_tiehi _14520__188 (.L_HI(net188));
 sg13g2_tiehi _14521__189 (.L_HI(net189));
 sg13g2_tiehi _14522__190 (.L_HI(net190));
 sg13g2_tiehi _14523__191 (.L_HI(net191));
 sg13g2_tiehi _14524__192 (.L_HI(net192));
 sg13g2_tiehi _14525__193 (.L_HI(net193));
 sg13g2_tiehi _14526__194 (.L_HI(net194));
 sg13g2_tiehi _14527__195 (.L_HI(net195));
 sg13g2_tiehi _14528__196 (.L_HI(net196));
 sg13g2_tiehi _14529__197 (.L_HI(net197));
 sg13g2_tiehi _14530__198 (.L_HI(net198));
 sg13g2_tiehi _14531__199 (.L_HI(net199));
 sg13g2_tiehi _14532__200 (.L_HI(net200));
 sg13g2_tiehi _14533__201 (.L_HI(net201));
 sg13g2_tiehi _14534__202 (.L_HI(net202));
 sg13g2_tiehi _14535__203 (.L_HI(net203));
 sg13g2_tiehi _14536__204 (.L_HI(net204));
 sg13g2_tiehi _14537__205 (.L_HI(net205));
 sg13g2_tiehi _14538__206 (.L_HI(net206));
 sg13g2_tiehi _14539__207 (.L_HI(net207));
 sg13g2_tiehi _14540__208 (.L_HI(net208));
 sg13g2_tiehi _14541__209 (.L_HI(net209));
 sg13g2_tiehi _14542__210 (.L_HI(net210));
 sg13g2_tiehi _14543__211 (.L_HI(net211));
 sg13g2_tiehi _14544__212 (.L_HI(net212));
 sg13g2_tiehi _14545__213 (.L_HI(net213));
 sg13g2_tiehi _14546__214 (.L_HI(net214));
 sg13g2_tiehi _14547__215 (.L_HI(net215));
 sg13g2_tiehi _14548__216 (.L_HI(net216));
 sg13g2_tiehi _14549__217 (.L_HI(net217));
 sg13g2_tiehi _14550__218 (.L_HI(net218));
 sg13g2_tiehi _14551__219 (.L_HI(net219));
 sg13g2_tiehi _14552__220 (.L_HI(net220));
 sg13g2_tiehi _14553__221 (.L_HI(net221));
 sg13g2_tiehi _14554__222 (.L_HI(net222));
 sg13g2_tiehi _14555__223 (.L_HI(net223));
 sg13g2_tiehi _14556__224 (.L_HI(net224));
 sg13g2_tiehi _14557__225 (.L_HI(net225));
 sg13g2_tiehi _14558__226 (.L_HI(net226));
 sg13g2_tiehi _14616__227 (.L_HI(net227));
 sg13g2_tiehi _14295__228 (.L_HI(net228));
 sg13g2_tiehi _14294__229 (.L_HI(net229));
 sg13g2_tiehi _14293__230 (.L_HI(net230));
 sg13g2_tiehi _14615__231 (.L_HI(net231));
 sg13g2_tiehi _14292__232 (.L_HI(net232));
 sg13g2_tiehi _14291__233 (.L_HI(net233));
 sg13g2_tiehi _14614__234 (.L_HI(net234));
 sg13g2_tiehi _14290__235 (.L_HI(net235));
 sg13g2_tiehi _14289__236 (.L_HI(net236));
 sg13g2_tiehi _14288__237 (.L_HI(net237));
 sg13g2_tiehi _14287__238 (.L_HI(net238));
 sg13g2_tiehi _14286__239 (.L_HI(net239));
 sg13g2_tiehi _14285__240 (.L_HI(net240));
 sg13g2_tiehi _14284__241 (.L_HI(net241));
 sg13g2_tiehi _14283__242 (.L_HI(net242));
 sg13g2_tiehi _14282__243 (.L_HI(net243));
 sg13g2_tiehi _14281__244 (.L_HI(net244));
 sg13g2_tiehi _14280__245 (.L_HI(net245));
 sg13g2_tiehi _14279__246 (.L_HI(net246));
 sg13g2_tiehi _14278__247 (.L_HI(net247));
 sg13g2_tiehi _14277__248 (.L_HI(net248));
 sg13g2_tiehi _14276__249 (.L_HI(net249));
 sg13g2_tiehi _14275__250 (.L_HI(net250));
 sg13g2_tiehi _14274__251 (.L_HI(net251));
 sg13g2_tiehi _14273__252 (.L_HI(net252));
 sg13g2_tiehi _14272__253 (.L_HI(net253));
 sg13g2_tiehi _14271__254 (.L_HI(net254));
 sg13g2_tiehi _14270__255 (.L_HI(net255));
 sg13g2_tiehi _14269__256 (.L_HI(net256));
 sg13g2_tiehi _14559__257 (.L_HI(net257));
 sg13g2_tiehi _14595__258 (.L_HI(net258));
 sg13g2_tiehi _14268__259 (.L_HI(net259));
 sg13g2_tiehi _14267__260 (.L_HI(net260));
 sg13g2_tiehi _14266__261 (.L_HI(net261));
 sg13g2_tiehi _14265__262 (.L_HI(net262));
 sg13g2_tiehi _14610__263 (.L_HI(net263));
 sg13g2_tiehi _14264__264 (.L_HI(net264));
 sg13g2_tiehi _14263__265 (.L_HI(net265));
 sg13g2_tiehi _14262__266 (.L_HI(net266));
 sg13g2_tiehi _14261__267 (.L_HI(net267));
 sg13g2_tiehi _14260__268 (.L_HI(net268));
 sg13g2_tiehi _14259__269 (.L_HI(net269));
 sg13g2_tiehi _14258__270 (.L_HI(net270));
 sg13g2_tiehi _14257__271 (.L_HI(net271));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_a1k0n_vgadonut_2 (.L_LO(net2));
 sg13g2_tielo tt_um_a1k0n_vgadonut_3 (.L_LO(net3));
 sg13g2_tielo tt_um_a1k0n_vgadonut_4 (.L_LO(net4));
 sg13g2_tielo tt_um_a1k0n_vgadonut_5 (.L_LO(net5));
 sg13g2_tielo tt_um_a1k0n_vgadonut_6 (.L_LO(net6));
 sg13g2_tielo tt_um_a1k0n_vgadonut_7 (.L_LO(net7));
 sg13g2_tielo tt_um_a1k0n_vgadonut_8 (.L_LO(net8));
 sg13g2_tielo tt_um_a1k0n_vgadonut_9 (.L_LO(net9));
 sg13g2_tielo tt_um_a1k0n_vgadonut_10 (.L_LO(net10));
 sg13g2_tielo tt_um_a1k0n_vgadonut_11 (.L_LO(net11));
 sg13g2_tielo tt_um_a1k0n_vgadonut_12 (.L_LO(net12));
 sg13g2_tielo tt_um_a1k0n_vgadonut_13 (.L_LO(net13));
 sg13g2_tielo tt_um_a1k0n_vgadonut_14 (.L_LO(net14));
 sg13g2_tielo tt_um_a1k0n_vgadonut_15 (.L_LO(net15));
 sg13g2_tielo tt_um_a1k0n_vgadonut_16 (.L_LO(net16));
 sg13g2_tiehi _14256__17 (.L_HI(net17));
 sg13g2_buf_2 _14892_ (.A(\vgadonut.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _14893_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout1492 (.A(_02860_),
    .X(net1492));
 sg13g2_buf_8 fanout1493 (.A(_02660_),
    .X(net1493));
 sg13g2_buf_8 fanout1494 (.A(_02320_),
    .X(net1494));
 sg13g2_buf_4 fanout1495 (.X(net1495),
    .A(_01896_));
 sg13g2_buf_2 fanout1496 (.A(_01884_),
    .X(net1496));
 sg13g2_buf_4 fanout1497 (.X(net1497),
    .A(_01877_));
 sg13g2_buf_4 fanout1498 (.X(net1498),
    .A(_01873_));
 sg13g2_buf_2 fanout1499 (.A(net1501),
    .X(net1499));
 sg13g2_buf_1 fanout1500 (.A(net1501),
    .X(net1500));
 sg13g2_buf_2 fanout1501 (.A(_01869_),
    .X(net1501));
 sg13g2_buf_2 fanout1502 (.A(net1503),
    .X(net1502));
 sg13g2_buf_4 fanout1503 (.X(net1503),
    .A(_01862_));
 sg13g2_buf_2 fanout1504 (.A(net1506),
    .X(net1504));
 sg13g2_buf_1 fanout1505 (.A(net1506),
    .X(net1505));
 sg13g2_buf_2 fanout1506 (.A(_01859_),
    .X(net1506));
 sg13g2_buf_4 fanout1507 (.X(net1507),
    .A(net1508));
 sg13g2_buf_8 fanout1508 (.A(_01853_),
    .X(net1508));
 sg13g2_buf_2 fanout1509 (.A(_01868_),
    .X(net1509));
 sg13g2_buf_2 fanout1510 (.A(net1512),
    .X(net1510));
 sg13g2_buf_2 fanout1511 (.A(net1512),
    .X(net1511));
 sg13g2_buf_4 fanout1512 (.X(net1512),
    .A(_01840_));
 sg13g2_buf_2 fanout1513 (.A(_01839_),
    .X(net1513));
 sg13g2_buf_1 fanout1514 (.A(_01839_),
    .X(net1514));
 sg13g2_buf_2 fanout1515 (.A(net1523),
    .X(net1515));
 sg13g2_buf_1 fanout1516 (.A(net1523),
    .X(net1516));
 sg13g2_buf_2 fanout1517 (.A(net1518),
    .X(net1517));
 sg13g2_buf_2 fanout1518 (.A(net1523),
    .X(net1518));
 sg13g2_buf_2 fanout1519 (.A(net1520),
    .X(net1519));
 sg13g2_buf_1 fanout1520 (.A(net1522),
    .X(net1520));
 sg13g2_buf_2 fanout1521 (.A(net1522),
    .X(net1521));
 sg13g2_buf_8 fanout1522 (.A(net1523),
    .X(net1522));
 sg13g2_buf_2 fanout1523 (.A(_01826_),
    .X(net1523));
 sg13g2_buf_2 fanout1524 (.A(_01825_),
    .X(net1524));
 sg13g2_buf_2 fanout1525 (.A(_01825_),
    .X(net1525));
 sg13g2_buf_2 fanout1526 (.A(net1529),
    .X(net1526));
 sg13g2_buf_2 fanout1527 (.A(net1529),
    .X(net1527));
 sg13g2_buf_2 fanout1528 (.A(net1529),
    .X(net1528));
 sg13g2_buf_2 fanout1529 (.A(_01820_),
    .X(net1529));
 sg13g2_buf_2 fanout1530 (.A(net1531),
    .X(net1530));
 sg13g2_buf_2 fanout1531 (.A(_01819_),
    .X(net1531));
 sg13g2_buf_4 fanout1532 (.X(net1532),
    .A(net1533));
 sg13g2_buf_1 fanout1533 (.A(net1534),
    .X(net1533));
 sg13g2_buf_2 fanout1534 (.A(net1537),
    .X(net1534));
 sg13g2_buf_2 fanout1535 (.A(net1536),
    .X(net1535));
 sg13g2_buf_2 fanout1536 (.A(net1537),
    .X(net1536));
 sg13g2_buf_4 fanout1537 (.X(net1537),
    .A(_01796_));
 sg13g2_buf_4 fanout1538 (.X(net1538),
    .A(net1539));
 sg13g2_buf_2 fanout1539 (.A(_01796_),
    .X(net1539));
 sg13g2_buf_2 fanout1540 (.A(net1541),
    .X(net1540));
 sg13g2_buf_2 fanout1541 (.A(_01793_),
    .X(net1541));
 sg13g2_buf_2 fanout1542 (.A(_01792_),
    .X(net1542));
 sg13g2_buf_2 fanout1543 (.A(net1544),
    .X(net1543));
 sg13g2_buf_2 fanout1544 (.A(_01791_),
    .X(net1544));
 sg13g2_buf_4 fanout1545 (.X(net1545),
    .A(_01790_));
 sg13g2_buf_2 fanout1546 (.A(_04988_),
    .X(net1546));
 sg13g2_buf_2 fanout1547 (.A(_04988_),
    .X(net1547));
 sg13g2_buf_4 fanout1548 (.X(net1548),
    .A(net1549));
 sg13g2_buf_2 fanout1549 (.A(_01530_),
    .X(net1549));
 sg13g2_buf_4 fanout1550 (.X(net1550),
    .A(_01530_));
 sg13g2_buf_2 fanout1551 (.A(net1552),
    .X(net1551));
 sg13g2_buf_2 fanout1552 (.A(net1569),
    .X(net1552));
 sg13g2_buf_4 fanout1553 (.X(net1553),
    .A(net1556));
 sg13g2_buf_4 fanout1554 (.X(net1554),
    .A(net1556));
 sg13g2_buf_1 fanout1555 (.A(net1556),
    .X(net1555));
 sg13g2_buf_2 fanout1556 (.A(net1569),
    .X(net1556));
 sg13g2_buf_4 fanout1557 (.X(net1557),
    .A(net1559));
 sg13g2_buf_1 fanout1558 (.A(net1559),
    .X(net1558));
 sg13g2_buf_2 fanout1559 (.A(net1563),
    .X(net1559));
 sg13g2_buf_2 fanout1560 (.A(net1563),
    .X(net1560));
 sg13g2_buf_2 fanout1561 (.A(net1563),
    .X(net1561));
 sg13g2_buf_2 fanout1562 (.A(net1563),
    .X(net1562));
 sg13g2_buf_2 fanout1563 (.A(net1569),
    .X(net1563));
 sg13g2_buf_4 fanout1564 (.X(net1564),
    .A(net1569));
 sg13g2_buf_2 fanout1565 (.A(net1567),
    .X(net1565));
 sg13g2_buf_2 fanout1566 (.A(net1567),
    .X(net1566));
 sg13g2_buf_2 fanout1567 (.A(net1568),
    .X(net1567));
 sg13g2_buf_2 fanout1568 (.A(net1569),
    .X(net1568));
 sg13g2_buf_4 fanout1569 (.X(net1569),
    .A(_04585_));
 sg13g2_buf_4 fanout1570 (.X(net1570),
    .A(_04584_));
 sg13g2_buf_4 fanout1571 (.X(net1571),
    .A(_04584_));
 sg13g2_buf_2 fanout1572 (.A(net1573),
    .X(net1572));
 sg13g2_buf_2 fanout1573 (.A(net1574),
    .X(net1573));
 sg13g2_buf_2 fanout1574 (.A(net1575),
    .X(net1574));
 sg13g2_buf_2 fanout1575 (.A(net1580),
    .X(net1575));
 sg13g2_buf_4 fanout1576 (.X(net1576),
    .A(net1577));
 sg13g2_buf_4 fanout1577 (.X(net1577),
    .A(net1579));
 sg13g2_buf_2 fanout1578 (.A(net1579),
    .X(net1578));
 sg13g2_buf_8 fanout1579 (.A(net1580),
    .X(net1579));
 sg13g2_buf_2 fanout1580 (.A(_01379_),
    .X(net1580));
 sg13g2_buf_2 fanout1581 (.A(net1582),
    .X(net1581));
 sg13g2_buf_2 fanout1582 (.A(net1583),
    .X(net1582));
 sg13g2_buf_2 fanout1583 (.A(net1584),
    .X(net1583));
 sg13g2_buf_2 fanout1584 (.A(_01378_),
    .X(net1584));
 sg13g2_buf_2 fanout1585 (.A(net1587),
    .X(net1585));
 sg13g2_buf_1 fanout1586 (.A(net1587),
    .X(net1586));
 sg13g2_buf_1 fanout1587 (.A(net1588),
    .X(net1587));
 sg13g2_buf_2 fanout1588 (.A(net1590),
    .X(net1588));
 sg13g2_buf_2 fanout1589 (.A(net1590),
    .X(net1589));
 sg13g2_buf_2 fanout1590 (.A(_01378_),
    .X(net1590));
 sg13g2_buf_4 fanout1591 (.X(net1591),
    .A(net1593));
 sg13g2_buf_2 fanout1592 (.A(net1593),
    .X(net1592));
 sg13g2_buf_4 fanout1593 (.X(net1593),
    .A(_01377_));
 sg13g2_buf_4 fanout1594 (.X(net1594),
    .A(net1596));
 sg13g2_buf_2 fanout1595 (.A(net1596),
    .X(net1595));
 sg13g2_buf_8 fanout1596 (.A(_01377_),
    .X(net1596));
 sg13g2_buf_4 fanout1597 (.X(net1597),
    .A(_04781_));
 sg13g2_buf_2 fanout1598 (.A(net1599),
    .X(net1598));
 sg13g2_buf_2 fanout1599 (.A(_04926_),
    .X(net1599));
 sg13g2_buf_2 fanout1600 (.A(_04523_),
    .X(net1600));
 sg13g2_buf_1 fanout1601 (.A(_04523_),
    .X(net1601));
 sg13g2_buf_2 fanout1602 (.A(_06179_),
    .X(net1602));
 sg13g2_buf_2 fanout1603 (.A(_06179_),
    .X(net1603));
 sg13g2_buf_2 fanout1604 (.A(net1607),
    .X(net1604));
 sg13g2_buf_4 fanout1605 (.X(net1605),
    .A(net1606));
 sg13g2_buf_2 fanout1606 (.A(net1607),
    .X(net1606));
 sg13g2_buf_2 fanout1607 (.A(_04712_),
    .X(net1607));
 sg13g2_buf_4 fanout1608 (.X(net1608),
    .A(net1609));
 sg13g2_buf_4 fanout1609 (.X(net1609),
    .A(net1612));
 sg13g2_buf_8 fanout1610 (.A(net1611),
    .X(net1610));
 sg13g2_buf_4 fanout1611 (.X(net1611),
    .A(net1612));
 sg13g2_buf_4 fanout1612 (.X(net1612),
    .A(_01106_));
 sg13g2_buf_2 fanout1613 (.A(net1614),
    .X(net1613));
 sg13g2_buf_4 fanout1614 (.X(net1614),
    .A(_05508_));
 sg13g2_buf_2 fanout1615 (.A(_00672_),
    .X(net1615));
 sg13g2_buf_4 fanout1616 (.X(net1616),
    .A(net1618));
 sg13g2_buf_2 fanout1617 (.A(net1618),
    .X(net1617));
 sg13g2_buf_2 fanout1618 (.A(_00921_),
    .X(net1618));
 sg13g2_buf_4 fanout1619 (.X(net1619),
    .A(_05418_));
 sg13g2_buf_4 fanout1620 (.X(net1620),
    .A(net1621));
 sg13g2_buf_2 fanout1621 (.A(net1622),
    .X(net1621));
 sg13g2_buf_2 fanout1622 (.A(net1628),
    .X(net1622));
 sg13g2_buf_4 fanout1623 (.X(net1623),
    .A(net1626));
 sg13g2_buf_4 fanout1624 (.X(net1624),
    .A(net1625));
 sg13g2_buf_2 fanout1625 (.A(net1626),
    .X(net1625));
 sg13g2_buf_2 fanout1626 (.A(net1627),
    .X(net1626));
 sg13g2_buf_2 fanout1627 (.A(net1628),
    .X(net1627));
 sg13g2_buf_2 fanout1628 (.A(_00898_),
    .X(net1628));
 sg13g2_buf_2 fanout1629 (.A(net1631),
    .X(net1629));
 sg13g2_buf_1 fanout1630 (.A(net1631),
    .X(net1630));
 sg13g2_buf_1 fanout1631 (.A(_00293_),
    .X(net1631));
 sg13g2_buf_2 fanout1632 (.A(net1633),
    .X(net1632));
 sg13g2_buf_1 fanout1633 (.A(net1634),
    .X(net1633));
 sg13g2_buf_2 fanout1634 (.A(_00291_),
    .X(net1634));
 sg13g2_buf_2 fanout1635 (.A(net1636),
    .X(net1635));
 sg13g2_buf_2 fanout1636 (.A(_00290_),
    .X(net1636));
 sg13g2_buf_2 fanout1637 (.A(net1638),
    .X(net1637));
 sg13g2_buf_1 fanout1638 (.A(net1639),
    .X(net1638));
 sg13g2_buf_1 fanout1639 (.A(_00292_),
    .X(net1639));
 sg13g2_buf_4 fanout1640 (.X(net1640),
    .A(_06705_));
 sg13g2_buf_2 fanout1641 (.A(_06705_),
    .X(net1641));
 sg13g2_buf_2 fanout1642 (.A(_00681_),
    .X(net1642));
 sg13g2_buf_2 fanout1643 (.A(net1645),
    .X(net1643));
 sg13g2_buf_2 fanout1644 (.A(net1645),
    .X(net1644));
 sg13g2_buf_1 fanout1645 (.A(_00674_),
    .X(net1645));
 sg13g2_buf_4 fanout1646 (.X(net1646),
    .A(_00666_));
 sg13g2_buf_4 fanout1647 (.X(net1647),
    .A(_00288_));
 sg13g2_buf_2 fanout1648 (.A(net1649),
    .X(net1648));
 sg13g2_buf_2 fanout1649 (.A(net1650),
    .X(net1649));
 sg13g2_buf_1 fanout1650 (.A(net1652),
    .X(net1650));
 sg13g2_buf_2 fanout1651 (.A(net1652),
    .X(net1651));
 sg13g2_buf_2 fanout1652 (.A(net1653),
    .X(net1652));
 sg13g2_buf_4 fanout1653 (.X(net1653),
    .A(net1669));
 sg13g2_buf_2 fanout1654 (.A(net1655),
    .X(net1654));
 sg13g2_buf_2 fanout1655 (.A(net1656),
    .X(net1655));
 sg13g2_buf_2 fanout1656 (.A(net1669),
    .X(net1656));
 sg13g2_buf_2 fanout1657 (.A(net1669),
    .X(net1657));
 sg13g2_buf_2 fanout1658 (.A(net1659),
    .X(net1658));
 sg13g2_buf_2 fanout1659 (.A(net1661),
    .X(net1659));
 sg13g2_buf_2 fanout1660 (.A(net1661),
    .X(net1660));
 sg13g2_buf_2 fanout1661 (.A(net1668),
    .X(net1661));
 sg13g2_buf_2 fanout1662 (.A(net1663),
    .X(net1662));
 sg13g2_buf_2 fanout1663 (.A(net1667),
    .X(net1663));
 sg13g2_buf_2 fanout1664 (.A(net1665),
    .X(net1664));
 sg13g2_buf_1 fanout1665 (.A(net1666),
    .X(net1665));
 sg13g2_buf_1 fanout1666 (.A(net1667),
    .X(net1666));
 sg13g2_buf_2 fanout1667 (.A(net1668),
    .X(net1667));
 sg13g2_buf_4 fanout1668 (.X(net1668),
    .A(net1669));
 sg13g2_buf_4 fanout1669 (.X(net1669),
    .A(_03935_));
 sg13g2_buf_8 fanout1670 (.A(_03934_),
    .X(net1670));
 sg13g2_buf_2 fanout1671 (.A(net1672),
    .X(net1671));
 sg13g2_buf_2 fanout1672 (.A(_00664_),
    .X(net1672));
 sg13g2_buf_4 fanout1673 (.X(net1673),
    .A(_00663_));
 sg13g2_buf_2 fanout1674 (.A(net1675),
    .X(net1674));
 sg13g2_buf_4 fanout1675 (.X(net1675),
    .A(_00663_));
 sg13g2_buf_4 fanout1676 (.X(net1676),
    .A(net1677));
 sg13g2_buf_4 fanout1677 (.X(net1677),
    .A(net1680));
 sg13g2_buf_2 fanout1678 (.A(net1679),
    .X(net1678));
 sg13g2_buf_4 fanout1679 (.X(net1679),
    .A(net1680));
 sg13g2_buf_2 fanout1680 (.A(_00663_),
    .X(net1680));
 sg13g2_buf_2 fanout1681 (.A(net1682),
    .X(net1681));
 sg13g2_buf_2 fanout1682 (.A(net1685),
    .X(net1682));
 sg13g2_buf_2 fanout1683 (.A(net1685),
    .X(net1683));
 sg13g2_buf_2 fanout1684 (.A(net1685),
    .X(net1684));
 sg13g2_buf_4 fanout1685 (.X(net1685),
    .A(net1700));
 sg13g2_buf_2 fanout1686 (.A(net1687),
    .X(net1686));
 sg13g2_buf_2 fanout1687 (.A(net1688),
    .X(net1687));
 sg13g2_buf_4 fanout1688 (.X(net1688),
    .A(net1689));
 sg13g2_buf_4 fanout1689 (.X(net1689),
    .A(net1700));
 sg13g2_buf_2 fanout1690 (.A(net1691),
    .X(net1690));
 sg13g2_buf_2 fanout1691 (.A(net1692),
    .X(net1691));
 sg13g2_buf_2 fanout1692 (.A(net1693),
    .X(net1692));
 sg13g2_buf_2 fanout1693 (.A(net1699),
    .X(net1693));
 sg13g2_buf_2 fanout1694 (.A(net1698),
    .X(net1694));
 sg13g2_buf_1 fanout1695 (.A(net1698),
    .X(net1695));
 sg13g2_buf_2 fanout1696 (.A(net1697),
    .X(net1696));
 sg13g2_buf_4 fanout1697 (.X(net1697),
    .A(net1698));
 sg13g2_buf_2 fanout1698 (.A(net1699),
    .X(net1698));
 sg13g2_buf_8 fanout1699 (.A(net1700),
    .X(net1699));
 sg13g2_buf_4 fanout1700 (.X(net1700),
    .A(_00662_));
 sg13g2_buf_4 fanout1701 (.X(net1701),
    .A(_05251_));
 sg13g2_buf_4 fanout1702 (.X(net1702),
    .A(net1703));
 sg13g2_buf_4 fanout1703 (.X(net1703),
    .A(net1705));
 sg13g2_buf_4 fanout1704 (.X(net1704),
    .A(net1705));
 sg13g2_buf_2 fanout1705 (.A(_04046_),
    .X(net1705));
 sg13g2_buf_4 fanout1706 (.X(net1706),
    .A(net1708));
 sg13g2_buf_1 fanout1707 (.A(net1708),
    .X(net1707));
 sg13g2_buf_4 fanout1708 (.X(net1708),
    .A(net1709));
 sg13g2_buf_4 fanout1709 (.X(net1709),
    .A(_04045_));
 sg13g2_buf_2 fanout1710 (.A(net1711),
    .X(net1710));
 sg13g2_buf_2 fanout1711 (.A(net1712),
    .X(net1711));
 sg13g2_buf_2 fanout1712 (.A(net1713),
    .X(net1712));
 sg13g2_buf_4 fanout1713 (.X(net1713),
    .A(_04044_));
 sg13g2_buf_4 fanout1714 (.X(net1714),
    .A(net1716));
 sg13g2_buf_2 fanout1715 (.A(net1716),
    .X(net1715));
 sg13g2_buf_4 fanout1716 (.X(net1716),
    .A(_04044_));
 sg13g2_buf_2 fanout1717 (.A(net1718),
    .X(net1717));
 sg13g2_buf_4 fanout1718 (.X(net1718),
    .A(net1730));
 sg13g2_buf_2 fanout1719 (.A(net1723),
    .X(net1719));
 sg13g2_buf_2 fanout1720 (.A(net1723),
    .X(net1720));
 sg13g2_buf_4 fanout1721 (.X(net1721),
    .A(net1723));
 sg13g2_buf_1 fanout1722 (.A(net1723),
    .X(net1722));
 sg13g2_buf_2 fanout1723 (.A(net1730),
    .X(net1723));
 sg13g2_buf_2 fanout1724 (.A(net1725),
    .X(net1724));
 sg13g2_buf_2 fanout1725 (.A(net1726),
    .X(net1725));
 sg13g2_buf_2 fanout1726 (.A(net1727),
    .X(net1726));
 sg13g2_buf_2 fanout1727 (.A(net1730),
    .X(net1727));
 sg13g2_buf_4 fanout1728 (.X(net1728),
    .A(net1730));
 sg13g2_buf_2 fanout1729 (.A(net1730),
    .X(net1729));
 sg13g2_buf_4 fanout1730 (.X(net1730),
    .A(_03925_));
 sg13g2_buf_2 fanout1731 (.A(net1733),
    .X(net1731));
 sg13g2_buf_2 fanout1732 (.A(net1733),
    .X(net1732));
 sg13g2_buf_2 fanout1733 (.A(_03925_),
    .X(net1733));
 sg13g2_buf_2 fanout1734 (.A(net1736),
    .X(net1734));
 sg13g2_buf_2 fanout1735 (.A(net1736),
    .X(net1735));
 sg13g2_buf_2 fanout1736 (.A(net1737),
    .X(net1736));
 sg13g2_buf_2 fanout1737 (.A(_03925_),
    .X(net1737));
 sg13g2_buf_2 fanout1738 (.A(net1739),
    .X(net1738));
 sg13g2_buf_1 fanout1739 (.A(net1740),
    .X(net1739));
 sg13g2_buf_2 fanout1740 (.A(net1741),
    .X(net1740));
 sg13g2_buf_2 fanout1741 (.A(_02949_),
    .X(net1741));
 sg13g2_buf_4 fanout1742 (.X(net1742),
    .A(net1743));
 sg13g2_buf_4 fanout1743 (.X(net1743),
    .A(net1747));
 sg13g2_buf_4 fanout1744 (.X(net1744),
    .A(net1747));
 sg13g2_buf_4 fanout1745 (.X(net1745),
    .A(net1746));
 sg13g2_buf_4 fanout1746 (.X(net1746),
    .A(net1747));
 sg13g2_buf_4 fanout1747 (.X(net1747),
    .A(_03932_));
 sg13g2_buf_8 fanout1748 (.A(net1749),
    .X(net1748));
 sg13g2_buf_8 fanout1749 (.A(_03931_),
    .X(net1749));
 sg13g2_buf_4 fanout1750 (.X(net1750),
    .A(net1752));
 sg13g2_buf_1 fanout1751 (.A(net1752),
    .X(net1751));
 sg13g2_buf_8 fanout1752 (.A(_03929_),
    .X(net1752));
 sg13g2_buf_4 fanout1753 (.X(net1753),
    .A(net1756));
 sg13g2_buf_2 fanout1754 (.A(net1755),
    .X(net1754));
 sg13g2_buf_4 fanout1755 (.X(net1755),
    .A(net1756));
 sg13g2_buf_4 fanout1756 (.X(net1756),
    .A(_03929_));
 sg13g2_buf_8 fanout1757 (.A(net1759),
    .X(net1757));
 sg13g2_buf_2 fanout1758 (.A(net1759),
    .X(net1758));
 sg13g2_buf_8 fanout1759 (.A(_03928_),
    .X(net1759));
 sg13g2_buf_8 fanout1760 (.A(_03927_),
    .X(net1760));
 sg13g2_buf_4 fanout1761 (.X(net1761),
    .A(net1764));
 sg13g2_buf_2 fanout1762 (.A(net1764),
    .X(net1762));
 sg13g2_buf_4 fanout1763 (.X(net1763),
    .A(net1764));
 sg13g2_buf_8 fanout1764 (.A(_03924_),
    .X(net1764));
 sg13g2_buf_2 fanout1765 (.A(net1766),
    .X(net1765));
 sg13g2_buf_2 fanout1766 (.A(net1769),
    .X(net1766));
 sg13g2_buf_2 fanout1767 (.A(net1768),
    .X(net1767));
 sg13g2_buf_1 fanout1768 (.A(net1769),
    .X(net1768));
 sg13g2_buf_2 fanout1769 (.A(net1773),
    .X(net1769));
 sg13g2_buf_4 fanout1770 (.X(net1770),
    .A(net1773));
 sg13g2_buf_4 fanout1771 (.X(net1771),
    .A(net1772));
 sg13g2_buf_2 fanout1772 (.A(net1773),
    .X(net1772));
 sg13g2_buf_4 fanout1773 (.X(net1773),
    .A(_03923_));
 sg13g2_buf_4 fanout1774 (.X(net1774),
    .A(net1775));
 sg13g2_buf_4 fanout1775 (.X(net1775),
    .A(net1776));
 sg13g2_buf_4 fanout1776 (.X(net1776),
    .A(net1777));
 sg13g2_buf_8 fanout1777 (.A(_03922_),
    .X(net1777));
 sg13g2_buf_2 fanout1778 (.A(net1780),
    .X(net1778));
 sg13g2_buf_1 fanout1779 (.A(net1780),
    .X(net1779));
 sg13g2_buf_2 fanout1780 (.A(net1786),
    .X(net1780));
 sg13g2_buf_2 fanout1781 (.A(net1786),
    .X(net1781));
 sg13g2_buf_2 fanout1782 (.A(net1783),
    .X(net1782));
 sg13g2_buf_2 fanout1783 (.A(net1784),
    .X(net1783));
 sg13g2_buf_2 fanout1784 (.A(net1786),
    .X(net1784));
 sg13g2_buf_2 fanout1785 (.A(net1786),
    .X(net1785));
 sg13g2_buf_2 fanout1786 (.A(_00788_),
    .X(net1786));
 sg13g2_buf_2 fanout1787 (.A(net1789),
    .X(net1787));
 sg13g2_buf_1 fanout1788 (.A(net1789),
    .X(net1788));
 sg13g2_buf_2 fanout1789 (.A(net1790),
    .X(net1789));
 sg13g2_buf_2 fanout1790 (.A(net1796),
    .X(net1790));
 sg13g2_buf_2 fanout1791 (.A(net1795),
    .X(net1791));
 sg13g2_buf_2 fanout1792 (.A(net1795),
    .X(net1792));
 sg13g2_buf_2 fanout1793 (.A(net1794),
    .X(net1793));
 sg13g2_buf_2 fanout1794 (.A(net1795),
    .X(net1794));
 sg13g2_buf_2 fanout1795 (.A(net1796),
    .X(net1795));
 sg13g2_buf_2 fanout1796 (.A(_00787_),
    .X(net1796));
 sg13g2_buf_4 fanout1797 (.X(net1797),
    .A(_00599_));
 sg13g2_buf_2 fanout1798 (.A(_00599_),
    .X(net1798));
 sg13g2_buf_4 fanout1799 (.X(net1799),
    .A(\vgadonut.donut.frame ));
 sg13g2_buf_2 fanout1800 (.A(\vgadonut.donut.h_count[4] ),
    .X(net1800));
 sg13g2_buf_4 fanout1801 (.X(net1801),
    .A(\vgadonut.donut.h_count[2] ));
 sg13g2_buf_4 fanout1802 (.X(net1802),
    .A(\vgadonut.donut.h_count[1] ));
 sg13g2_buf_2 fanout1803 (.A(net2322),
    .X(net1803));
 sg13g2_buf_4 fanout1804 (.X(net1804),
    .A(net1805));
 sg13g2_buf_4 fanout1805 (.X(net1805),
    .A(\vgadonut.donut.donuthit.cordicxy.xinvert ));
 sg13g2_buf_4 fanout1806 (.X(net1806),
    .A(net1807));
 sg13g2_buf_4 fanout1807 (.X(net1807),
    .A(net1808));
 sg13g2_buf_4 fanout1808 (.X(net1808),
    .A(\vgadonut.donut.donuthit.cordicxy.xinvert ));
 sg13g2_buf_4 fanout1809 (.X(net1809),
    .A(net1812));
 sg13g2_buf_2 fanout1810 (.A(net1811),
    .X(net1810));
 sg13g2_buf_2 fanout1811 (.A(net1812),
    .X(net1811));
 sg13g2_buf_2 fanout1812 (.A(net1813),
    .X(net1812));
 sg13g2_buf_8 fanout1813 (.A(net2212),
    .X(net1813));
 sg13g2_buf_4 fanout1814 (.X(net1814),
    .A(\vgadonut.donut.cA[14] ));
 sg13g2_buf_4 fanout1815 (.X(net1815),
    .A(\vgadonut.donut.cA[13] ));
 sg13g2_buf_4 fanout1816 (.X(net1816),
    .A(\vgadonut.donut.cA[13] ));
 sg13g2_buf_4 fanout1817 (.X(net1817),
    .A(\vgadonut.donut.cA[12] ));
 sg13g2_buf_2 fanout1818 (.A(\vgadonut.donut.cA[12] ),
    .X(net1818));
 sg13g2_buf_4 fanout1819 (.X(net1819),
    .A(\vgadonut.donut.cA[11] ));
 sg13g2_buf_2 fanout1820 (.A(\vgadonut.donut.cA[11] ),
    .X(net1820));
 sg13g2_buf_8 fanout1821 (.A(\vgadonut.donut.cA[10] ),
    .X(net1821));
 sg13g2_buf_4 fanout1822 (.X(net1822),
    .A(\vgadonut.donut.cA[9] ));
 sg13g2_buf_4 fanout1823 (.X(net1823),
    .A(\vgadonut.donut.cA[8] ));
 sg13g2_buf_4 fanout1824 (.X(net1824),
    .A(net2278));
 sg13g2_buf_4 fanout1825 (.X(net1825),
    .A(\vgadonut.donut.cA[2] ));
 sg13g2_buf_4 fanout1826 (.X(net1826),
    .A(net1830));
 sg13g2_buf_2 fanout1827 (.A(net1830),
    .X(net1827));
 sg13g2_buf_2 fanout1828 (.A(net1829),
    .X(net1828));
 sg13g2_buf_2 fanout1829 (.A(net1830),
    .X(net1829));
 sg13g2_buf_4 fanout1830 (.X(net1830),
    .A(\vgadonut.donut.sA[15] ));
 sg13g2_buf_4 fanout1831 (.X(net1831),
    .A(\vgadonut.donut.sA[14] ));
 sg13g2_buf_4 fanout1832 (.X(net1832),
    .A(net1833));
 sg13g2_buf_2 fanout1833 (.A(\vgadonut.donut.sA[13] ),
    .X(net1833));
 sg13g2_buf_4 fanout1834 (.X(net1834),
    .A(net1836));
 sg13g2_buf_2 fanout1835 (.A(net1836),
    .X(net1835));
 sg13g2_buf_2 fanout1836 (.A(net2350),
    .X(net1836));
 sg13g2_buf_4 fanout1837 (.X(net1837),
    .A(net1839));
 sg13g2_buf_2 fanout1838 (.A(net1839),
    .X(net1838));
 sg13g2_buf_2 fanout1839 (.A(\vgadonut.donut.sA[11] ),
    .X(net1839));
 sg13g2_buf_4 fanout1840 (.X(net1840),
    .A(net1841));
 sg13g2_buf_2 fanout1841 (.A(\vgadonut.donut.sA[10] ),
    .X(net1841));
 sg13g2_buf_4 fanout1842 (.X(net1842),
    .A(\vgadonut.donut.sA[9] ));
 sg13g2_buf_2 fanout1843 (.A(net2230),
    .X(net1843));
 sg13g2_buf_4 fanout1844 (.X(net1844),
    .A(\vgadonut.donut.sA[8] ));
 sg13g2_buf_2 fanout1845 (.A(\vgadonut.donut.sA[8] ),
    .X(net1845));
 sg13g2_buf_4 fanout1846 (.X(net1846),
    .A(net2251));
 sg13g2_buf_2 fanout1847 (.A(\vgadonut.donut.sA[7] ),
    .X(net1847));
 sg13g2_buf_4 fanout1848 (.X(net1848),
    .A(net1849));
 sg13g2_buf_4 fanout1849 (.X(net1849),
    .A(\vgadonut.donut.sA[6] ));
 sg13g2_buf_4 fanout1850 (.X(net1850),
    .A(\vgadonut.donut.sA[5] ));
 sg13g2_buf_2 fanout1851 (.A(\vgadonut.donut.sA[5] ),
    .X(net1851));
 sg13g2_buf_4 fanout1852 (.X(net1852),
    .A(\vgadonut.donut.sA[4] ));
 sg13g2_buf_4 fanout1853 (.X(net1853),
    .A(\vgadonut.donut.sA[3] ));
 sg13g2_buf_4 fanout1854 (.X(net1854),
    .A(\vgadonut.donut.sA[2] ));
 sg13g2_buf_2 fanout1855 (.A(net1856),
    .X(net1855));
 sg13g2_buf_4 fanout1856 (.X(net1856),
    .A(net1857));
 sg13g2_buf_2 fanout1857 (.A(net2059),
    .X(net1857));
 sg13g2_buf_2 fanout1858 (.A(_00125_),
    .X(net1858));
 sg13g2_buf_4 fanout1859 (.X(net1859),
    .A(net1860));
 sg13g2_buf_2 fanout1860 (.A(net1861),
    .X(net1860));
 sg13g2_buf_2 fanout1861 (.A(net2200),
    .X(net1861));
 sg13g2_buf_2 fanout1862 (.A(\vgadonut.donut.cB[14] ),
    .X(net1862));
 sg13g2_buf_4 fanout1863 (.X(net1863),
    .A(net2285));
 sg13g2_buf_4 fanout1864 (.X(net1864),
    .A(net2220));
 sg13g2_buf_1 fanout1865 (.A(\vgadonut.donut.cB[2] ),
    .X(net1865));
 sg13g2_buf_4 fanout1866 (.X(net1866),
    .A(net2294));
 sg13g2_buf_4 fanout1867 (.X(net1867),
    .A(net2313));
 sg13g2_buf_2 fanout1868 (.A(net1869),
    .X(net1868));
 sg13g2_buf_2 fanout1869 (.A(net1870),
    .X(net1869));
 sg13g2_buf_2 fanout1870 (.A(net2240),
    .X(net1870));
 sg13g2_buf_4 fanout1871 (.X(net1871),
    .A(net2266));
 sg13g2_buf_1 fanout1872 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[12] ),
    .X(net1872));
 sg13g2_buf_4 fanout1873 (.X(net1873),
    .A(net2221));
 sg13g2_buf_1 fanout1874 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[11] ),
    .X(net1874));
 sg13g2_buf_4 fanout1875 (.X(net1875),
    .A(net1876));
 sg13g2_buf_2 fanout1876 (.A(net2228),
    .X(net1876));
 sg13g2_buf_4 fanout1877 (.X(net1877),
    .A(net2254));
 sg13g2_buf_1 fanout1878 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[9] ),
    .X(net1878));
 sg13g2_buf_4 fanout1879 (.X(net1879),
    .A(\vgadonut.donut.donuthit.cordicxy.x2in[8] ));
 sg13g2_buf_4 fanout1880 (.X(net1880),
    .A(net2267));
 sg13g2_buf_1 fanout1881 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[7] ),
    .X(net1881));
 sg13g2_buf_4 fanout1882 (.X(net1882),
    .A(net2341));
 sg13g2_buf_4 fanout1883 (.X(net1883),
    .A(net2331));
 sg13g2_buf_4 fanout1884 (.X(net1884),
    .A(net2288));
 sg13g2_buf_2 fanout1885 (.A(net1886),
    .X(net1885));
 sg13g2_buf_2 fanout1886 (.A(net2272),
    .X(net1886));
 sg13g2_buf_4 fanout1887 (.X(net1887),
    .A(net2340));
 sg13g2_buf_4 fanout1888 (.X(net1888),
    .A(net2348));
 sg13g2_buf_4 fanout1889 (.X(net1889),
    .A(net2304));
 sg13g2_buf_2 fanout1890 (.A(\vgadonut.donut.sAsB[2] ),
    .X(net1890));
 sg13g2_buf_4 fanout1891 (.X(net1891),
    .A(net2317));
 sg13g2_buf_2 fanout1892 (.A(net2270),
    .X(net1892));
 sg13g2_buf_2 fanout1893 (.A(\vgadonut.donut.sAsB[0] ),
    .X(net1893));
 sg13g2_buf_4 fanout1894 (.X(net1894),
    .A(net1896));
 sg13g2_buf_4 fanout1895 (.X(net1895),
    .A(net1896));
 sg13g2_buf_2 fanout1896 (.A(\vgadonut.donut.cAsB[15] ),
    .X(net1896));
 sg13g2_buf_4 fanout1897 (.X(net1897),
    .A(net2306));
 sg13g2_buf_4 fanout1898 (.X(net1898),
    .A(net1899));
 sg13g2_buf_2 fanout1899 (.A(net2213),
    .X(net1899));
 sg13g2_buf_4 fanout1900 (.X(net1900),
    .A(net2334));
 sg13g2_buf_4 fanout1901 (.X(net1901),
    .A(net2298));
 sg13g2_buf_4 fanout1902 (.X(net1902),
    .A(\vgadonut.donut.cAsB[10] ));
 sg13g2_buf_2 fanout1903 (.A(\vgadonut.donut.cAsB[9] ),
    .X(net1903));
 sg13g2_buf_2 fanout1904 (.A(\vgadonut.donut.cAsB[8] ),
    .X(net1904));
 sg13g2_buf_4 fanout1905 (.X(net1905),
    .A(net2231));
 sg13g2_buf_2 fanout1906 (.A(net2284),
    .X(net1906));
 sg13g2_buf_2 fanout1907 (.A(\vgadonut.donut.cAsB[5] ),
    .X(net1907));
 sg13g2_buf_4 fanout1908 (.X(net1908),
    .A(net2281));
 sg13g2_buf_4 fanout1909 (.X(net1909),
    .A(\vgadonut.donut.cAsB[3] ));
 sg13g2_buf_2 fanout1910 (.A(\vgadonut.donut.cAsB[2] ),
    .X(net1910));
 sg13g2_buf_4 fanout1911 (.X(net1911),
    .A(net2269));
 sg13g2_buf_2 fanout1912 (.A(\vgadonut.donut.cAsB[0] ),
    .X(net1912));
 sg13g2_buf_2 fanout1913 (.A(net2305),
    .X(net1913));
 sg13g2_buf_2 fanout1914 (.A(net2218),
    .X(net1914));
 sg13g2_buf_2 fanout1915 (.A(net1478),
    .X(net1915));
 sg13g2_buf_2 fanout1916 (.A(net1917),
    .X(net1916));
 sg13g2_buf_2 fanout1917 (.A(net1918),
    .X(net1917));
 sg13g2_buf_4 fanout1918 (.X(net1918),
    .A(net2279));
 sg13g2_buf_4 fanout1919 (.X(net1919),
    .A(net2318));
 sg13g2_buf_2 fanout1920 (.A(net1921),
    .X(net1920));
 sg13g2_buf_4 fanout1921 (.X(net1921),
    .A(\vgadonut.donut.sAcB[13] ));
 sg13g2_buf_4 fanout1922 (.X(net1922),
    .A(net2349));
 sg13g2_buf_1 fanout1923 (.A(\vgadonut.donut.sAcB[12] ),
    .X(net1923));
 sg13g2_buf_2 fanout1924 (.A(net1925),
    .X(net1924));
 sg13g2_buf_4 fanout1925 (.X(net1925),
    .A(\vgadonut.donut.sAcB[11] ));
 sg13g2_buf_4 fanout1926 (.X(net1926),
    .A(net1927));
 sg13g2_buf_2 fanout1927 (.A(\vgadonut.donut.sAcB[10] ),
    .X(net1927));
 sg13g2_buf_4 fanout1928 (.X(net1928),
    .A(net2333));
 sg13g2_buf_4 fanout1929 (.X(net1929),
    .A(\vgadonut.donut.sAcB[8] ));
 sg13g2_buf_4 fanout1930 (.X(net1930),
    .A(net2330));
 sg13g2_buf_4 fanout1931 (.X(net1931),
    .A(net2324));
 sg13g2_buf_4 fanout1932 (.X(net1932),
    .A(\vgadonut.donut.sAcB[5] ));
 sg13g2_buf_2 fanout1933 (.A(\vgadonut.donut.sAcB[5] ),
    .X(net1933));
 sg13g2_buf_4 fanout1934 (.X(net1934),
    .A(\vgadonut.donut.sAcB[4] ));
 sg13g2_buf_4 fanout1935 (.X(net1935),
    .A(net2347));
 sg13g2_buf_4 fanout1936 (.X(net1936),
    .A(net1937));
 sg13g2_buf_2 fanout1937 (.A(net2256),
    .X(net1937));
 sg13g2_buf_4 fanout1938 (.X(net1938),
    .A(net1939));
 sg13g2_buf_4 fanout1939 (.X(net1939),
    .A(\vgadonut.donut.cAcB[13] ));
 sg13g2_buf_4 fanout1940 (.X(net1940),
    .A(net1941));
 sg13g2_buf_2 fanout1941 (.A(net2226),
    .X(net1941));
 sg13g2_buf_4 fanout1942 (.X(net1942),
    .A(net1943));
 sg13g2_buf_4 fanout1943 (.X(net1943),
    .A(\vgadonut.donut.cAcB[11] ));
 sg13g2_buf_4 fanout1944 (.X(net1944),
    .A(net1945));
 sg13g2_buf_2 fanout1945 (.A(\vgadonut.donut.cAcB[10] ),
    .X(net1945));
 sg13g2_buf_4 fanout1946 (.X(net1946),
    .A(net1947));
 sg13g2_buf_4 fanout1947 (.X(net1947),
    .A(net2217));
 sg13g2_buf_4 fanout1948 (.X(net1948),
    .A(\vgadonut.donut.cAcB[8] ));
 sg13g2_buf_4 fanout1949 (.X(net1949),
    .A(net1950));
 sg13g2_buf_2 fanout1950 (.A(net2225),
    .X(net1950));
 sg13g2_buf_4 fanout1951 (.X(net1951),
    .A(net1952));
 sg13g2_buf_2 fanout1952 (.A(net2229),
    .X(net1952));
 sg13g2_buf_4 fanout1953 (.X(net1953),
    .A(net1954));
 sg13g2_buf_2 fanout1954 (.A(\vgadonut.donut.cAcB[5] ),
    .X(net1954));
 sg13g2_buf_2 fanout1955 (.A(net1956),
    .X(net1955));
 sg13g2_buf_4 fanout1956 (.X(net1956),
    .A(\vgadonut.donut.cAcB[4] ));
 sg13g2_buf_4 fanout1957 (.X(net1957),
    .A(\vgadonut.donut.cAcB[3] ));
 sg13g2_buf_4 fanout1958 (.X(net1958),
    .A(net1960));
 sg13g2_buf_4 fanout1959 (.X(net1959),
    .A(net1960));
 sg13g2_buf_4 fanout1960 (.X(net1960),
    .A(net1966));
 sg13g2_buf_4 fanout1961 (.X(net1961),
    .A(net1966));
 sg13g2_buf_4 fanout1962 (.X(net1962),
    .A(net1966));
 sg13g2_buf_4 fanout1963 (.X(net1963),
    .A(net1965));
 sg13g2_buf_4 fanout1964 (.X(net1964),
    .A(net1965));
 sg13g2_buf_2 fanout1965 (.A(net1966),
    .X(net1965));
 sg13g2_buf_4 fanout1966 (.X(net1966),
    .A(rst_n));
 sg13g2_buf_4 fanout1967 (.X(net1967),
    .A(net1968));
 sg13g2_buf_4 fanout1968 (.X(net1968),
    .A(net1969));
 sg13g2_buf_4 fanout1969 (.X(net1969),
    .A(net1970));
 sg13g2_buf_4 fanout1970 (.X(net1970),
    .A(net1976));
 sg13g2_buf_4 fanout1971 (.X(net1971),
    .A(net1972));
 sg13g2_buf_4 fanout1972 (.X(net1972),
    .A(net1975));
 sg13g2_buf_2 fanout1973 (.A(net1975),
    .X(net1973));
 sg13g2_buf_4 fanout1974 (.X(net1974),
    .A(net1975));
 sg13g2_buf_2 fanout1975 (.A(net1976),
    .X(net1975));
 sg13g2_buf_4 fanout1976 (.X(net1976),
    .A(rst_n));
 sg13g2_buf_4 fanout1977 (.X(net1977),
    .A(net1978));
 sg13g2_buf_4 fanout1978 (.X(net1978),
    .A(net1979));
 sg13g2_buf_4 fanout1979 (.X(net1979),
    .A(net1984));
 sg13g2_buf_4 fanout1980 (.X(net1980),
    .A(net1983));
 sg13g2_buf_4 fanout1981 (.X(net1981),
    .A(net1982));
 sg13g2_buf_4 fanout1982 (.X(net1982),
    .A(net1983));
 sg13g2_buf_2 fanout1983 (.A(net1984),
    .X(net1983));
 sg13g2_buf_4 fanout1984 (.X(net1984),
    .A(rst_n));
 sg13g2_tielo tt_um_a1k0n_vgadonut_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_4_8_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_9_0_clk));
 sg13g2_buf_1 clkload10 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload12 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_13_0_clk));
 sg13g2_buf_2 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_70_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_71_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_7_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_64_clk));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_67_clk));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_68_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_10_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_63_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_14_clk));
 sg13g2_inv_2 clkload30 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload31 (.A(clknet_leaf_17_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_19_clk));
 sg13g2_inv_1 clkload33 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload34 (.A(clknet_leaf_22_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_23_clk));
 sg13g2_inv_4 clkload36 (.A(clknet_leaf_12_clk));
 sg13g2_inv_2 clkload37 (.A(clknet_leaf_13_clk));
 sg13g2_inv_2 clkload38 (.A(clknet_leaf_18_clk));
 sg13g2_inv_4 clkload39 (.A(clknet_leaf_25_clk));
 sg13g2_inv_8 clkload40 (.A(clknet_leaf_24_clk));
 sg13g2_inv_1 clkload41 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload42 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload43 (.A(clknet_leaf_57_clk));
 sg13g2_inv_4 clkload44 (.A(clknet_leaf_66_clk));
 sg13g2_inv_2 clkload45 (.A(clknet_leaf_58_clk));
 sg13g2_inv_4 clkload46 (.A(clknet_leaf_59_clk));
 sg13g2_inv_1 clkload47 (.A(clknet_leaf_61_clk));
 sg13g2_inv_1 clkload48 (.A(clknet_leaf_51_clk));
 sg13g2_inv_1 clkload49 (.A(clknet_leaf_52_clk));
 sg13g2_inv_4 clkload50 (.A(clknet_leaf_53_clk));
 sg13g2_inv_1 clkload51 (.A(clknet_leaf_54_clk));
 sg13g2_inv_1 clkload52 (.A(clknet_leaf_47_clk));
 sg13g2_inv_1 clkload53 (.A(clknet_leaf_50_clk));
 sg13g2_inv_4 clkload54 (.A(clknet_leaf_60_clk));
 sg13g2_inv_1 clkload55 (.A(clknet_leaf_11_clk));
 sg13g2_inv_8 clkload56 (.A(clknet_leaf_30_clk));
 sg13g2_inv_4 clkload57 (.A(clknet_leaf_32_clk));
 sg13g2_inv_4 clkload58 (.A(clknet_leaf_33_clk));
 sg13g2_inv_2 clkload59 (.A(clknet_leaf_34_clk));
 sg13g2_inv_4 clkload60 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload61 (.A(clknet_leaf_40_clk));
 sg13g2_inv_4 clkload62 (.A(clknet_leaf_45_clk));
 sg13g2_inv_2 clkload63 (.A(clknet_leaf_46_clk));
 sg13g2_inv_4 clkload64 (.A(clknet_leaf_36_clk));
 sg13g2_inv_4 clkload65 (.A(clknet_leaf_38_clk));
 sg13g2_buf_1 rebuffer1 (.A(_01222_),
    .X(net272));
 sg13g2_buf_1 rebuffer2 (.A(_01317_),
    .X(net273));
 sg13g2_dlygate4sd1_1 rebuffer3 (.A(_00810_),
    .X(net274));
 sg13g2_dlygate4sd1_1 rebuffer4 (.A(_00810_),
    .X(net275));
 sg13g2_buf_1 rebuffer5 (.A(_00804_),
    .X(net276));
 sg13g2_dlygate4sd1_1 rebuffer6 (.A(_00804_),
    .X(net277));
 sg13g2_dlygate4sd1_1 rebuffer7 (.A(net281),
    .X(net278));
 sg13g2_dlygate4sd1_1 rebuffer8 (.A(_01031_),
    .X(net279));
 sg13g2_dlygate4sd1_1 rebuffer9 (.A(_00872_),
    .X(net280));
 sg13g2_dlygate4sd3_1 rebuffer10 (.A(net282),
    .X(net281));
 sg13g2_buf_1 rebuffer11 (.A(_00868_),
    .X(net282));
 sg13g2_dlygate4sd1_1 rebuffer12 (.A(_00897_),
    .X(net283));
 sg13g2_buf_1 rebuffer13 (.A(net283),
    .X(net284));
 sg13g2_dlygate4sd1_1 rebuffer14 (.A(_00865_),
    .X(net285));
 sg13g2_dlygate4sd1_1 rebuffer15 (.A(_00817_),
    .X(net286));
 sg13g2_dlygate4sd1_1 rebuffer16 (.A(_01007_),
    .X(net287));
 sg13g2_dlygate4sd1_1 rebuffer17 (.A(_01010_),
    .X(net288));
 sg13g2_dlygate4sd1_1 rebuffer18 (.A(net288),
    .X(net289));
 sg13g2_dlygate4sd1_1 rebuffer19 (.A(_00876_),
    .X(net290));
 sg13g2_dlygate4sd1_1 rebuffer20 (.A(\vgadonut.donut.donuthit.cordicxy.yin[1] ),
    .X(net291));
 sg13g2_dlygate4sd1_1 rebuffer21 (.A(\vgadonut.donut.donuthit.cordicxy.yin[1] ),
    .X(net292));
 sg13g2_buf_1 rebuffer22 (.A(\vgadonut.donut.donuthit.cordicxy.yin[1] ),
    .X(net293));
 sg13g2_dlygate4sd1_1 rebuffer23 (.A(\vgadonut.donut.donuthit.cordicxy.yin[5] ),
    .X(net294));
 sg13g2_buf_1 rebuffer24 (.A(\vgadonut.donut.donuthit.cordicxy.yin[5] ),
    .X(net295));
 sg13g2_dlygate4sd1_1 rebuffer25 (.A(\vgadonut.donut.donuthit.cordicxy.yin[2] ),
    .X(net296));
 sg13g2_dlygate4sd1_1 rebuffer26 (.A(\vgadonut.donut.donuthit.cordicxy.yin[2] ),
    .X(net297));
 sg13g2_buf_1 rebuffer27 (.A(\vgadonut.donut.donuthit.cordicxy.yin[2] ),
    .X(net298));
 sg13g2_buf_8 rebuffer28 (.A(_01478_),
    .X(net299));
 sg13g2_buf_8 rebuffer29 (.A(net1363),
    .X(net300));
 sg13g2_buf_8 rebuffer1092 (.A(net1364),
    .X(net1363));
 sg13g2_buf_2 rebuffer1093 (.A(net1365),
    .X(net1364));
 sg13g2_buf_2 rebuffer1094 (.A(net1366),
    .X(net1365));
 sg13g2_dlygate4sd1_1 rebuffer1095 (.A(net1367),
    .X(net1366));
 sg13g2_dlygate4sd1_1 rebuffer1096 (.A(net1368),
    .X(net1367));
 sg13g2_dlygate4sd1_1 rebuffer1097 (.A(net1369),
    .X(net1368));
 sg13g2_dlygate4sd1_1 rebuffer1098 (.A(net1370),
    .X(net1369));
 sg13g2_dlygate4sd1_1 rebuffer1099 (.A(net1371),
    .X(net1370));
 sg13g2_dlygate4sd1_1 rebuffer1100 (.A(net1372),
    .X(net1371));
 sg13g2_dlygate4sd1_1 rebuffer1101 (.A(net1373),
    .X(net1372));
 sg13g2_dlygate4sd1_1 rebuffer1102 (.A(net1374),
    .X(net1373));
 sg13g2_dlygate4sd1_1 rebuffer1103 (.A(net1375),
    .X(net1374));
 sg13g2_dlygate4sd1_1 rebuffer1104 (.A(net1376),
    .X(net1375));
 sg13g2_dlygate4sd1_1 rebuffer1105 (.A(net1377),
    .X(net1376));
 sg13g2_dlygate4sd1_1 rebuffer1106 (.A(net1378),
    .X(net1377));
 sg13g2_dlygate4sd1_1 rebuffer1107 (.A(net1379),
    .X(net1378));
 sg13g2_dlygate4sd1_1 rebuffer1108 (.A(net1380),
    .X(net1379));
 sg13g2_dlygate4sd1_1 rebuffer1109 (.A(net1381),
    .X(net1380));
 sg13g2_dlygate4sd1_1 rebuffer1110 (.A(net1382),
    .X(net1381));
 sg13g2_dlygate4sd1_1 rebuffer1111 (.A(net1383),
    .X(net1382));
 sg13g2_dlygate4sd1_1 rebuffer1112 (.A(net1384),
    .X(net1383));
 sg13g2_dlygate4sd1_1 rebuffer1113 (.A(net1385),
    .X(net1384));
 sg13g2_dlygate4sd1_1 rebuffer1114 (.A(net1386),
    .X(net1385));
 sg13g2_dlygate4sd1_1 rebuffer1115 (.A(net1387),
    .X(net1386));
 sg13g2_dlygate4sd1_1 rebuffer1116 (.A(net1388),
    .X(net1387));
 sg13g2_dlygate4sd1_1 rebuffer1117 (.A(net1389),
    .X(net1388));
 sg13g2_dlygate4sd1_1 rebuffer1118 (.A(net1390),
    .X(net1389));
 sg13g2_dlygate4sd1_1 rebuffer1119 (.A(net1391),
    .X(net1390));
 sg13g2_dlygate4sd1_1 rebuffer1120 (.A(net1392),
    .X(net1391));
 sg13g2_dlygate4sd1_1 rebuffer1121 (.A(net1393),
    .X(net1392));
 sg13g2_dlygate4sd1_1 rebuffer1122 (.A(net1394),
    .X(net1393));
 sg13g2_dlygate4sd1_1 rebuffer1123 (.A(net1395),
    .X(net1394));
 sg13g2_dlygate4sd1_1 rebuffer1124 (.A(net1396),
    .X(net1395));
 sg13g2_dlygate4sd1_1 rebuffer1125 (.A(net1397),
    .X(net1396));
 sg13g2_dlygate4sd1_1 rebuffer1126 (.A(net1398),
    .X(net1397));
 sg13g2_dlygate4sd1_1 rebuffer1127 (.A(net1399),
    .X(net1398));
 sg13g2_dlygate4sd1_1 rebuffer1128 (.A(net1400),
    .X(net1399));
 sg13g2_dlygate4sd1_1 rebuffer1129 (.A(net1401),
    .X(net1400));
 sg13g2_dlygate4sd1_1 rebuffer1130 (.A(net1402),
    .X(net1401));
 sg13g2_dlygate4sd1_1 rebuffer1131 (.A(net1403),
    .X(net1402));
 sg13g2_dlygate4sd1_1 rebuffer1132 (.A(net1404),
    .X(net1403));
 sg13g2_dlygate4sd1_1 rebuffer1133 (.A(net1405),
    .X(net1404));
 sg13g2_dlygate4sd1_1 rebuffer1134 (.A(net1406),
    .X(net1405));
 sg13g2_dlygate4sd1_1 rebuffer1135 (.A(net1407),
    .X(net1406));
 sg13g2_dlygate4sd1_1 rebuffer1136 (.A(net1408),
    .X(net1407));
 sg13g2_dlygate4sd1_1 rebuffer1137 (.A(net1409),
    .X(net1408));
 sg13g2_dlygate4sd1_1 rebuffer1138 (.A(net1410),
    .X(net1409));
 sg13g2_dlygate4sd1_1 rebuffer1139 (.A(net1411),
    .X(net1410));
 sg13g2_dlygate4sd1_1 rebuffer1140 (.A(net1412),
    .X(net1411));
 sg13g2_dlygate4sd1_1 rebuffer1141 (.A(net1413),
    .X(net1412));
 sg13g2_dlygate4sd1_1 rebuffer1142 (.A(net1414),
    .X(net1413));
 sg13g2_dlygate4sd1_1 rebuffer1143 (.A(net1415),
    .X(net1414));
 sg13g2_dlygate4sd1_1 rebuffer1144 (.A(net1416),
    .X(net1415));
 sg13g2_dlygate4sd1_1 rebuffer1145 (.A(net1417),
    .X(net1416));
 sg13g2_dlygate4sd1_1 rebuffer1146 (.A(net1418),
    .X(net1417));
 sg13g2_dlygate4sd1_1 rebuffer1147 (.A(net1419),
    .X(net1418));
 sg13g2_dlygate4sd1_1 rebuffer1148 (.A(net1420),
    .X(net1419));
 sg13g2_dlygate4sd1_1 rebuffer1149 (.A(net1421),
    .X(net1420));
 sg13g2_dlygate4sd1_1 rebuffer1150 (.A(net1422),
    .X(net1421));
 sg13g2_dlygate4sd1_1 rebuffer1151 (.A(net1423),
    .X(net1422));
 sg13g2_dlygate4sd1_1 rebuffer1152 (.A(net1424),
    .X(net1423));
 sg13g2_dlygate4sd1_1 rebuffer1153 (.A(net1425),
    .X(net1424));
 sg13g2_dlygate4sd1_1 rebuffer1154 (.A(net1426),
    .X(net1425));
 sg13g2_dlygate4sd1_1 rebuffer1155 (.A(net1427),
    .X(net1426));
 sg13g2_dlygate4sd1_1 rebuffer1156 (.A(net1428),
    .X(net1427));
 sg13g2_dlygate4sd1_1 rebuffer1157 (.A(net1429),
    .X(net1428));
 sg13g2_dlygate4sd1_1 rebuffer1158 (.A(net1430),
    .X(net1429));
 sg13g2_dlygate4sd1_1 rebuffer1159 (.A(net1431),
    .X(net1430));
 sg13g2_dlygate4sd1_1 rebuffer1160 (.A(net1432),
    .X(net1431));
 sg13g2_dlygate4sd1_1 rebuffer1161 (.A(net1433),
    .X(net1432));
 sg13g2_dlygate4sd1_1 rebuffer1162 (.A(net1434),
    .X(net1433));
 sg13g2_dlygate4sd1_1 rebuffer1163 (.A(net1435),
    .X(net1434));
 sg13g2_dlygate4sd1_1 rebuffer1164 (.A(net1436),
    .X(net1435));
 sg13g2_dlygate4sd1_1 rebuffer1165 (.A(net1437),
    .X(net1436));
 sg13g2_dlygate4sd1_1 rebuffer1166 (.A(net1438),
    .X(net1437));
 sg13g2_dlygate4sd1_1 rebuffer1167 (.A(net1439),
    .X(net1438));
 sg13g2_dlygate4sd1_1 rebuffer1168 (.A(net1440),
    .X(net1439));
 sg13g2_dlygate4sd1_1 rebuffer1169 (.A(net1441),
    .X(net1440));
 sg13g2_dlygate4sd1_1 rebuffer1170 (.A(net1442),
    .X(net1441));
 sg13g2_buf_2 rebuffer1171 (.A(net1443),
    .X(net1442));
 sg13g2_buf_2 rebuffer1172 (.A(\vgadonut.donut.donuthit.cordicxy.yin[1] ),
    .X(net1443));
 sg13g2_dlygate4sd1_1 rebuffer1173 (.A(_01317_),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold1174 (.A(_00179_),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold1175 (.A(_00015_),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold1176 (.A(_00181_),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold1177 (.A(_00538_),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold1178 (.A(_00189_),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold1179 (.A(_00194_),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold1180 (.A(_00202_),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold1181 (.A(_00199_),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold1182 (.A(_00193_),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold1183 (.A(_00198_),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold1184 (.A(_00183_),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold1185 (.A(_00182_),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold1186 (.A(_00196_),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold1187 (.A(_00191_),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold1188 (.A(_00205_),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold1189 (.A(_00445_),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold1190 (.A(_00203_),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold1191 (.A(_00443_),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold1192 (.A(_00218_),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold1193 (.A(_00222_),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold1194 (.A(_00220_),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold1195 (.A(_00204_),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold1196 (.A(_00444_),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold1197 (.A(_00190_),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold1198 (.A(_00188_),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold1199 (.A(_00210_),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold1200 (.A(_00209_),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold1201 (.A(_00197_),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold1202 (.A(_00221_),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold1203 (.A(_00184_),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold1204 (.A(_00192_),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold1205 (.A(_00310_),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold1206 (.A(_00187_),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\vgadonut.bayer_j[0] ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold1208 (.A(_00185_),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold1209 (.A(_00195_),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold1210 (.A(_00217_),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold1211 (.A(_00207_),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold1212 (.A(_00213_),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold1213 (.A(_00459_),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold1214 (.A(_00215_),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold1215 (.A(_00216_),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold1216 (.A(_00219_),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold1217 (.A(_00214_),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold1218 (.A(_00186_),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold1219 (.A(_00212_),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold1220 (.A(_00211_),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold1221 (.A(_00208_),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\vgadonut.donut.cAsB[0] ),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\vgadonut.donut.rx6[0] ),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold1224 (.A(_03936_),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\vgadonut.donut.sAsB[2] ),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold1226 (.A(_00206_),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold1227 (.A(_00177_),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\vgadonut.donut.cAsB[8] ),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\vgadonut.donut.ycA[0] ),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold1230 (.A(_04432_),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\vgadonut.donut.cAsB[9] ),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\vgadonut.donut.rz6[2] ),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\vgadonut.donut.cAsB[5] ),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\vgadonut.donut.ry6[4] ),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\vgadonut.donut.rz6[1] ),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold1236 (.A(_00478_),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\vgadonut.donut.ry6[3] ),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\vgadonut.donut.h_count[1] ),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold1239 (.A(_00016_),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\vgadonut.donut.donuthit.hit ),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\vgadonut.donut.ry6[0] ),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\vgadonut.donut.cAsB[3] ),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\vgadonut.donut.donuthit.light[8] ),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold1244 (.A(_00288_),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\vgadonut.donut.ry6[1] ),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold1246 (.A(_00369_),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\vgadonut.donut.rx6[3] ),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\vgadonut.donut.rx6[2] ),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold1249 (.A(_00390_),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\vgadonut.donut.donuthit.rz[6] ),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\vgadonut.donut.rz6[0] ),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold1252 (.A(_00477_),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\vgadonut.donut.donuthit.t[0] ),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\vgadonut.donut.ysA[0] ),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold1255 (.A(_04441_),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\vgadonut.donut.donuthit.ryin[12] ),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold1257 (.A(_00517_),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\vgadonut.donut.sAsB[3] ),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\vgadonut.donut.donuthit.rz[12] ),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold1260 (.A(_00528_),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold1261 (.A(_00178_),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\vgadonut.donut.v_count[7] ),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold1263 (.A(_00333_),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\vgadonut.donut.cAsB[2] ),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\vgadonut.donut.donuthit.rz[15] ),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold1266 (.A(_00531_),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\vgadonut.donut.ycA[3] ),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\vgadonut.donut.ycA[21] ),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\vgadonut.frame[1] ),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold1270 (.A(_00539_),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\vgadonut.donut.donuthit.ry[13] ),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold1272 (.A(_00518_),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\vgadonut.donut.rz6[3] ),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\vgadonut.donut.ysA[1] ),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\vgadonut.donut.cA[9] ),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\vgadonut.donut.donuthit.ryin[2] ),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\vgadonut.donut.donuthit.ryin[6] ),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold1278 (.A(_00511_),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\vgadonut.donut.donuthit.rxin[0] ),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\vgadonut.frame[7] ),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold1281 (.A(_00545_),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\vgadonut.donut.donuthit.rz[9] ),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold1283 (.A(_00525_),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\vgadonut.donut.donuthit.ryin[3] ),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\vgadonut.donut.donuthit.ry[10] ),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold1286 (.A(_00515_),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\vgadonut.donut.donuthit.ry[8] ),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold1288 (.A(_00513_),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\vgadonut.donut.ysA[2] ),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\vgadonut.donut.donuthit.rz[10] ),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold1291 (.A(_00526_),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\vgadonut.donut.donuthit.ry[11] ),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold1293 (.A(_00516_),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\vgadonut.donut.donuthit.rxin[4] ),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\vgadonut.donut.donut_visible ),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\vgadonut.donut.rx6[4] ),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold1297 (.A(_00392_),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\vgadonut.donut.h_count[9] ),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold1299 (.A(_00024_),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\vgadonut.donut.ry6[2] ),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\vgadonut.donut.donuthit.ryin[1] ),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\vgadonut.donut.donuthit.rzin[1] ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\vgadonut.donut.donuthit.rz[8] ),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold1304 (.A(_00524_),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\vgadonut.donut.v_count[8] ),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold1306 (.A(_00334_),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\vgadonut.donut.donuthit.rx[8] ),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold1308 (.A(_00502_),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\vgadonut.donut.rx6[1] ),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\vgadonut.donut.donuthit.rz[14] ),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold1311 (.A(_00530_),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\vgadonut.donut.h_count[7] ),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold1313 (.A(_02986_),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold1314 (.A(_00025_),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\vgadonut.donut.donuthit.ryin[4] ),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\vgadonut.donut.donuthit.ryin[0] ),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold1317 (.A(_00374_),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\vgadonut.frame[2] ),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold1319 (.A(_00540_),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\vgadonut.donut.donuthit.rxin[1] ),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\vgadonut.donut.donuthit.rzin[2] ),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\vgadonut.donut.donuthit.rzin[0] ),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\vgadonut.donut.donuthit.ry[9] ),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold1324 (.A(_00514_),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\vgadonut.frame[6] ),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold1326 (.A(_00544_),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\vgadonut.donut.ycA[1] ),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\vgadonut.donut.donuthit.rx[9] ),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold1329 (.A(_00503_),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold1330 (.A(_00154_),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\vgadonut.donut.donuthit.rxin[2] ),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\vgadonut.donut.ycA[20] ),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\vgadonut.donut.ysA[4] ),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\vgadonut.donut.rx6[5] ),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\vgadonut.donut.donuthit.rxin[3] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\vgadonut.donut.donuthit.rz[5] ),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold1337 (.A(_00521_),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\vgadonut.frame[5] ),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold1339 (.A(_06843_),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\vgadonut.donut.donuthit.rxin[6] ),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold1341 (.A(_00500_),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\vgadonut.donut.rz6[4] ),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\vgadonut.donut.rz6[5] ),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\vgadonut.donut.h_count[4] ),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\vgadonut.donut.ry6[5] ),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\vgadonut.donut.donuthit.rx[7] ),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold1347 (.A(_00501_),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\vgadonut.donut.v_count[6] ),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold1349 (.A(_00332_),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\vgadonut.donut.donuthit.rz[7] ),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold1351 (.A(_00523_),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\vgadonut.donut.donuthit.ry[15] ),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold1353 (.A(_00520_),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\vgadonut.donut.donuthit.rzin[4] ),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold1355 (.A(_00200_),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\vgadonut.donut.donuthit.rx[11] ),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold1357 (.A(_00505_),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\vgadonut.donut.donuthit.rx[10] ),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold1359 (.A(_00504_),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\vgadonut.donut.sA[15] ),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold1361 (.A(_04235_),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\vgadonut.frame[3] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold1363 (.A(_00201_),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\vgadonut.donut.donuthit.ry[14] ),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold1365 (.A(_00519_),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\vgadonut.donut.donuthit.rzin[3] ),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\vgadonut.donut.donuthit.rz[11] ),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold1368 (.A(_00527_),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\vgadonut.donut.ycA[14] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\vgadonut.donut.donuthit.ry[7] ),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold1371 (.A(_00512_),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\vgadonut.donut.ycA[2] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\vgadonut.donut.ycA[7] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\vgadonut.donut.donuthit.rz[13] ),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold1375 (.A(_00529_),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\vgadonut.donut.ysA[19] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\vgadonut.donut.sB[0] ),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\vgadonut.donut.h_count[6] ),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold1379 (.A(_02961_),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\vgadonut.donut.donuthit.rx[15] ),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold1381 (.A(_00509_),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold1382 (.A(_00180_),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold1383 (.A(_00331_),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[1] ),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold1385 (.A(_00413_),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\vgadonut.donut.ycA[15] ),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\vgadonut.donut.donuthit.rzin[14] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\vgadonut.donut.ysA[14] ),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\vgadonut.donut.sAsB[10] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\vgadonut.donut.donuthit.light[11] ),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold1391 (.A(_00674_),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\vgadonut.donut.donuthit.rx[5] ),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold1393 (.A(_00499_),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\vgadonut.donut.ycA[16] ),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\vgadonut.donut.h_count[6] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\vgadonut.frame[4] ),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\vgadonut.donut.h_count[8] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\vgadonut.donut.donuthit.ry[5] ),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold1399 (.A(_00510_),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\vgadonut.donut.donuthit.rzin[11] ),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\vgadonut.donut.ysA[15] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\vgadonut.donut.v_count[9] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\vgadonut.donut.ysA[6] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\vgadonut.donut.sB[1] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold1405 (.A(_00411_),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\vgadonut.donut.ysA[20] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\vgadonut.donut.donuthit.rzin[9] ),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\vgadonut.donut.ysA[7] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\vgadonut.donut.donuthit.rzin[12] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\vgadonut.donut.ysA[8] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\vgadonut.donut.ycA[19] ),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\vgadonut.donut.cB[11] ),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\vgadonut.donut.ysA[3] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\vgadonut.donut.ysA[11] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\vgadonut.donut.donuthit.rzin[10] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[3] ),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\vgadonut.donut.h_count[5] ),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold1418 (.A(_00160_),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold1419 (.A(_02200_),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\vgadonut.donut.ycA[4] ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold1421 (.A(_00261_),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\vgadonut.donut.donuthit.cordicxy.xin[15] ),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\vgadonut.donut.donuthit.ryin[9] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\vgadonut.donut.ysA[9] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\vgadonut.donut.donuthit.rzin[13] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\vgadonut.bayer_j[1] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\vgadonut.donut.ycA[6] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\vgadonut.donut.donuthit.rxin[13] ),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold1429 (.A(_00507_),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\vgadonut.donut.cA[2] ),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold1431 (.A(_00265_),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\vgadonut.donut.sAsB[13] ),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold1433 (.A(_00162_),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\vgadonut.donut.donuthit.rx[12] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold1435 (.A(_00506_),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\vgadonut.donut.cB[15] ),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\vgadonut.donut.ysA[16] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold1438 (.A(_00161_),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\vgadonut.donut.donuthit.rx[14] ),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold1440 (.A(_00508_),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\vgadonut.donut.cB[9] ),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\vgadonut.donut.donuthit.rxin[10] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\vgadonut.donut.donuthit.t[4] ),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold1444 (.A(_00231_),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\vgadonut.donut.donuthit.ryin[13] ),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\vgadonut.donut.ysA[5] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold1447 (.A(_00244_),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\vgadonut.donut.cA[15] ),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\vgadonut.donut.cAsB[13] ),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\vgadonut.donut.donuthit.rxin[11] ),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\vgadonut.donut.donuthit.ryin[15] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\vgadonut.donut.ysA[17] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\vgadonut.donut.cAcB[9] ),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\vgadonut.donut.v_count[2] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold1455 (.A(_00026_),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\vgadonut.donut.cB[2] ),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[11] ),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold1458 (.A(_00423_),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\vgadonut.donut.ycA[17] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\vgadonut.donut.cB[10] ),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\vgadonut.donut.cAcB[7] ),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\vgadonut.donut.cAcB[12] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\vgadonut.donut.donuthit.ryin[14] ),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[10] ),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\vgadonut.donut.cAcB[6] ),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\vgadonut.donut.sA[9] ),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\vgadonut.donut.cAsB[7] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\vgadonut.donut.donuthit.rzin[7] ),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\vgadonut.donut.cB[7] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\vgadonut.donut.donuthit.ryin[11] ),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\vgadonut.donut.v_count[4] ),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold1472 (.A(_00330_),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\vgadonut.donut.sAsB[7] ),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\vgadonut.donut.ycA[5] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\vgadonut.donut.ysA[13] ),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[13] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\vgadonut.donut.sAsB[14] ),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\vgadonut.donut.cB[8] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[8] ),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\vgadonut.donut.donuthit.rxin[8] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\vgadonut.donut.donuthit.rzin[8] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\vgadonut.donut.sAsB[8] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\vgadonut.donut.ycA[9] ),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\vgadonut.donut.cB[12] ),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\vgadonut.donut.donuthit.t[2] ),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold1486 (.A(_00229_),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\vgadonut.donut.sA[7] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\vgadonut.donut.donuthit.t[1] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold1489 (.A(_00168_),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[9] ),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold1491 (.A(_00421_),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\vgadonut.donut.cAcB[14] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\vgadonut.donut.donuthit.t[8] ),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold1494 (.A(_00234_),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\vgadonut.donut.cB[4] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\vgadonut.donut.ysA[18] ),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\vgadonut.donut.cB[6] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\vgadonut.donut.ycA[18] ),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\vgadonut.donut.sAsB[4] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\vgadonut.donut.donuthit.rzin[5] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[0] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[12] ),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[7] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\vgadonut.donut.cB[13] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\vgadonut.donut.cAsB[1] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\vgadonut.donut.sAsB[0] ),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\vgadonut.donut.donuthit.rxin[9] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\vgadonut.donut.sAsB[15] ),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\vgadonut.donut.donuthit.rxin[14] ),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\vgadonut.donut.donuthit.ryin[10] ),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\vgadonut.donut.donuthit.cordicxy.xin[0] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\vgadonut.donut.sAsB[9] ),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\vgadonut.donut.ycA[11] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\vgadonut.donut.cA[7] ),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\vgadonut.donut.sAcB[15] ),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\vgadonut.donut.ysA[12] ),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\vgadonut.donut.cAsB[4] ),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\vgadonut.donut.donuthit.ryin[7] ),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\vgadonut.donut.ysA[10] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\vgadonut.donut.cAsB[6] ),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\vgadonut.donut.cB[3] ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold1522 (.A(_00156_),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\vgadonut.donut.ycA[10] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[2] ),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold1525 (.A(_00414_),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\vgadonut.donut.donuthit.cordicxz.xin[0] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold1527 (.A(_02644_),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold1528 (.A(_02646_),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\vgadonut.donut.cB[5] ),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\vgadonut.donut.cB[1] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\vgadonut.donut.donuthit.t[6] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold1532 (.A(_03969_),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\vgadonut.donut.donuthit.rxin[15] ),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\vgadonut.donut.cAsB[11] ),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\vgadonut.donut.donuthit.rxin[7] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\vgadonut.donut.donuthit.t[10] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold1537 (.A(_00236_),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[5] ),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold1539 (.A(_00417_),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\vgadonut.donut.sAsB[5] ),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\vgadonut.donut.v_count[3] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\vgadonut.donut.cAsB[14] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold1543 (.A(_00167_),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\vgadonut.donut.donuthit.rxin[12] ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\vgadonut.donut.ycA[12] ),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\vgadonut.donut.donuthit.rzin[6] ),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold1547 (.A(_00141_),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold1548 (.A(_00457_),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\vgadonut.donut.cB[0] ),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\vgadonut.donut.donuthit.t[7] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\vgadonut.donut.donuthit.t[13] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold1552 (.A(_04032_),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\vgadonut.donut.sAsB[1] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\vgadonut.donut.sAcB[14] ),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\vgadonut.donut.donuthit.rzin[15] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\vgadonut.donut.sAsB[6] ),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold1557 (.A(_00142_),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\vgadonut.donut.h_count[0] ),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\vgadonut.donut.donuthit.t[15] ),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\vgadonut.donut.sAcB[6] ),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold1561 (.A(_00169_),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold1562 (.A(_00110_),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\vgadonut.donut.donuthit.ryin[8] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\vgadonut.donut.donuthit.t[11] ),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold1565 (.A(_00166_),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\vgadonut.donut.sAcB[7] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[4] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\vgadonut.donut.donuthit.rxin[5] ),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\vgadonut.donut.sAcB[9] ),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\vgadonut.donut.cAsB[12] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold1571 (.A(_00045_),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold1572 (.A(_00681_),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\vgadonut.donut.ycA[13] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\vgadonut.donut.donuthit.ryin[5] ),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold1575 (.A(_00062_),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\vgadonut.donut.sAsB[12] ),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\vgadonut.donut.donuthit.cordicxy.x2in[6] ),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold1578 (.A(_00043_),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold1579 (.A(_06832_),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold1580 (.A(_00032_),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold1581 (.A(_00114_),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\vgadonut.donut.donuthit.t[14] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\vgadonut.donut.cAcB[15] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\vgadonut.donut.sAsB[11] ),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\vgadonut.donut.sAcB[12] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\vgadonut.donut.sA[12] ),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\vgadonut.donut.v_count[8] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold1588 (.A(_00163_),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold1589 (.A(_00159_),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold1590 (.A(_00143_),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\vgadonut.donut.donuthit.t[15] ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\vgadonut.donut.donuthit.rzin[12] ),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold1593 (.A(_00166_),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\vgadonut.donut.donuthit.t[14] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold1595 (.A(_00164_),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\vgadonut.donut.ysA[2] ),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold1597 (.A(_00161_),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold1598 (.A(_00163_),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold1599 (.A(\vgadonut.donut.ysA[2] ),
    .X(net2363));
 sg13g2_antennanp ANTENNA_1 (.A(net1764));
 sg13g2_antennanp ANTENNA_2 (.A(net1764));
 sg13g2_antennanp ANTENNA_3 (.A(net1764));
 sg13g2_antennanp ANTENNA_4 (.A(net1764));
 sg13g2_antennanp ANTENNA_5 (.A(net1764));
 sg13g2_antennanp ANTENNA_6 (.A(net1764));
 sg13g2_antennanp ANTENNA_7 (.A(net1764));
 sg13g2_antennanp ANTENNA_8 (.A(net1764));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_fill_1 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_114 ();
 sg13g2_decap_4 FILLER_0_147 ();
 sg13g2_fill_1 FILLER_0_151 ();
 sg13g2_fill_2 FILLER_0_157 ();
 sg13g2_fill_2 FILLER_0_195 ();
 sg13g2_fill_1 FILLER_0_197 ();
 sg13g2_fill_2 FILLER_0_205 ();
 sg13g2_fill_2 FILLER_0_252 ();
 sg13g2_fill_1 FILLER_0_279 ();
 sg13g2_decap_4 FILLER_0_286 ();
 sg13g2_fill_2 FILLER_0_305 ();
 sg13g2_decap_4 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_fill_1 FILLER_0_438 ();
 sg13g2_fill_2 FILLER_0_465 ();
 sg13g2_decap_4 FILLER_0_493 ();
 sg13g2_decap_8 FILLER_0_534 ();
 sg13g2_fill_2 FILLER_0_541 ();
 sg13g2_decap_8 FILLER_0_556 ();
 sg13g2_decap_8 FILLER_0_563 ();
 sg13g2_fill_2 FILLER_0_575 ();
 sg13g2_fill_1 FILLER_0_602 ();
 sg13g2_fill_2 FILLER_0_607 ();
 sg13g2_fill_1 FILLER_0_609 ();
 sg13g2_decap_4 FILLER_0_615 ();
 sg13g2_fill_2 FILLER_0_623 ();
 sg13g2_fill_2 FILLER_0_638 ();
 sg13g2_decap_8 FILLER_0_653 ();
 sg13g2_decap_4 FILLER_0_660 ();
 sg13g2_fill_1 FILLER_0_721 ();
 sg13g2_fill_2 FILLER_0_748 ();
 sg13g2_fill_1 FILLER_0_750 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_fill_2 FILLER_1_28 ();
 sg13g2_fill_2 FILLER_1_39 ();
 sg13g2_fill_1 FILLER_1_74 ();
 sg13g2_decap_4 FILLER_1_120 ();
 sg13g2_fill_2 FILLER_1_134 ();
 sg13g2_fill_1 FILLER_1_163 ();
 sg13g2_fill_2 FILLER_1_178 ();
 sg13g2_fill_1 FILLER_1_273 ();
 sg13g2_fill_2 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_4 FILLER_1_366 ();
 sg13g2_fill_1 FILLER_1_370 ();
 sg13g2_decap_4 FILLER_1_380 ();
 sg13g2_fill_2 FILLER_1_410 ();
 sg13g2_fill_2 FILLER_1_426 ();
 sg13g2_fill_1 FILLER_1_428 ();
 sg13g2_fill_2 FILLER_1_520 ();
 sg13g2_fill_1 FILLER_1_522 ();
 sg13g2_fill_1 FILLER_1_535 ();
 sg13g2_fill_1 FILLER_1_608 ();
 sg13g2_fill_2 FILLER_1_635 ();
 sg13g2_fill_1 FILLER_1_637 ();
 sg13g2_fill_2 FILLER_1_671 ();
 sg13g2_decap_4 FILLER_1_698 ();
 sg13g2_decap_8 FILLER_1_746 ();
 sg13g2_fill_2 FILLER_1_753 ();
 sg13g2_decap_4 FILLER_1_761 ();
 sg13g2_decap_8 FILLER_1_788 ();
 sg13g2_decap_8 FILLER_1_795 ();
 sg13g2_decap_8 FILLER_1_802 ();
 sg13g2_decap_8 FILLER_1_809 ();
 sg13g2_decap_8 FILLER_1_816 ();
 sg13g2_decap_8 FILLER_1_823 ();
 sg13g2_decap_8 FILLER_1_830 ();
 sg13g2_decap_8 FILLER_1_837 ();
 sg13g2_decap_8 FILLER_1_844 ();
 sg13g2_decap_8 FILLER_1_851 ();
 sg13g2_decap_4 FILLER_1_858 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_4 FILLER_2_14 ();
 sg13g2_fill_1 FILLER_2_18 ();
 sg13g2_fill_2 FILLER_2_54 ();
 sg13g2_fill_1 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_fill_2 FILLER_2_84 ();
 sg13g2_fill_2 FILLER_2_112 ();
 sg13g2_fill_2 FILLER_2_124 ();
 sg13g2_fill_1 FILLER_2_153 ();
 sg13g2_fill_2 FILLER_2_166 ();
 sg13g2_fill_2 FILLER_2_177 ();
 sg13g2_fill_1 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_fill_2 FILLER_2_203 ();
 sg13g2_fill_1 FILLER_2_205 ();
 sg13g2_decap_4 FILLER_2_237 ();
 sg13g2_fill_1 FILLER_2_259 ();
 sg13g2_decap_4 FILLER_2_265 ();
 sg13g2_fill_1 FILLER_2_315 ();
 sg13g2_decap_4 FILLER_2_329 ();
 sg13g2_fill_1 FILLER_2_333 ();
 sg13g2_decap_4 FILLER_2_384 ();
 sg13g2_fill_1 FILLER_2_388 ();
 sg13g2_fill_2 FILLER_2_496 ();
 sg13g2_fill_1 FILLER_2_514 ();
 sg13g2_decap_4 FILLER_2_543 ();
 sg13g2_fill_2 FILLER_2_547 ();
 sg13g2_decap_4 FILLER_2_559 ();
 sg13g2_fill_1 FILLER_2_563 ();
 sg13g2_fill_2 FILLER_2_576 ();
 sg13g2_decap_4 FILLER_2_616 ();
 sg13g2_fill_2 FILLER_2_625 ();
 sg13g2_fill_2 FILLER_2_639 ();
 sg13g2_fill_2 FILLER_2_648 ();
 sg13g2_fill_1 FILLER_2_650 ();
 sg13g2_decap_4 FILLER_2_660 ();
 sg13g2_fill_1 FILLER_2_664 ();
 sg13g2_decap_4 FILLER_2_695 ();
 sg13g2_fill_1 FILLER_2_699 ();
 sg13g2_fill_2 FILLER_2_724 ();
 sg13g2_fill_1 FILLER_2_726 ();
 sg13g2_decap_8 FILLER_2_785 ();
 sg13g2_decap_8 FILLER_2_792 ();
 sg13g2_decap_8 FILLER_2_799 ();
 sg13g2_decap_8 FILLER_2_806 ();
 sg13g2_decap_8 FILLER_2_813 ();
 sg13g2_decap_8 FILLER_2_820 ();
 sg13g2_decap_8 FILLER_2_827 ();
 sg13g2_decap_8 FILLER_2_834 ();
 sg13g2_decap_8 FILLER_2_841 ();
 sg13g2_decap_8 FILLER_2_848 ();
 sg13g2_decap_8 FILLER_2_855 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_4 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_25 ();
 sg13g2_fill_1 FILLER_3_44 ();
 sg13g2_decap_4 FILLER_3_61 ();
 sg13g2_fill_2 FILLER_3_77 ();
 sg13g2_fill_1 FILLER_3_79 ();
 sg13g2_decap_4 FILLER_3_88 ();
 sg13g2_fill_1 FILLER_3_92 ();
 sg13g2_decap_4 FILLER_3_117 ();
 sg13g2_fill_2 FILLER_3_121 ();
 sg13g2_fill_2 FILLER_3_135 ();
 sg13g2_fill_2 FILLER_3_149 ();
 sg13g2_fill_1 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_fill_2 FILLER_3_203 ();
 sg13g2_fill_1 FILLER_3_205 ();
 sg13g2_fill_1 FILLER_3_226 ();
 sg13g2_fill_1 FILLER_3_238 ();
 sg13g2_fill_1 FILLER_3_249 ();
 sg13g2_fill_1 FILLER_3_277 ();
 sg13g2_fill_2 FILLER_3_294 ();
 sg13g2_fill_1 FILLER_3_296 ();
 sg13g2_fill_2 FILLER_3_333 ();
 sg13g2_fill_1 FILLER_3_335 ();
 sg13g2_decap_8 FILLER_3_339 ();
 sg13g2_decap_8 FILLER_3_346 ();
 sg13g2_decap_4 FILLER_3_364 ();
 sg13g2_fill_1 FILLER_3_368 ();
 sg13g2_fill_1 FILLER_3_373 ();
 sg13g2_decap_4 FILLER_3_381 ();
 sg13g2_fill_2 FILLER_3_411 ();
 sg13g2_fill_2 FILLER_3_442 ();
 sg13g2_fill_2 FILLER_3_449 ();
 sg13g2_fill_2 FILLER_3_463 ();
 sg13g2_fill_2 FILLER_3_470 ();
 sg13g2_fill_2 FILLER_3_480 ();
 sg13g2_fill_2 FILLER_3_580 ();
 sg13g2_decap_4 FILLER_3_608 ();
 sg13g2_decap_8 FILLER_3_632 ();
 sg13g2_decap_4 FILLER_3_639 ();
 sg13g2_fill_1 FILLER_3_643 ();
 sg13g2_fill_2 FILLER_3_649 ();
 sg13g2_fill_2 FILLER_3_674 ();
 sg13g2_fill_1 FILLER_3_711 ();
 sg13g2_fill_2 FILLER_3_736 ();
 sg13g2_fill_1 FILLER_3_738 ();
 sg13g2_decap_4 FILLER_3_753 ();
 sg13g2_fill_1 FILLER_3_757 ();
 sg13g2_decap_4 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_799 ();
 sg13g2_decap_8 FILLER_3_806 ();
 sg13g2_decap_8 FILLER_3_813 ();
 sg13g2_decap_8 FILLER_3_820 ();
 sg13g2_decap_8 FILLER_3_827 ();
 sg13g2_decap_8 FILLER_3_834 ();
 sg13g2_decap_8 FILLER_3_841 ();
 sg13g2_decap_8 FILLER_3_848 ();
 sg13g2_decap_8 FILLER_3_855 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_4 FILLER_4_14 ();
 sg13g2_fill_2 FILLER_4_18 ();
 sg13g2_fill_1 FILLER_4_52 ();
 sg13g2_fill_1 FILLER_4_60 ();
 sg13g2_decap_4 FILLER_4_69 ();
 sg13g2_fill_1 FILLER_4_76 ();
 sg13g2_fill_2 FILLER_4_90 ();
 sg13g2_decap_4 FILLER_4_119 ();
 sg13g2_fill_2 FILLER_4_123 ();
 sg13g2_fill_2 FILLER_4_166 ();
 sg13g2_fill_1 FILLER_4_168 ();
 sg13g2_fill_2 FILLER_4_192 ();
 sg13g2_fill_2 FILLER_4_219 ();
 sg13g2_fill_1 FILLER_4_221 ();
 sg13g2_fill_2 FILLER_4_270 ();
 sg13g2_fill_2 FILLER_4_293 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_4 FILLER_4_310 ();
 sg13g2_fill_1 FILLER_4_314 ();
 sg13g2_fill_2 FILLER_4_325 ();
 sg13g2_fill_1 FILLER_4_327 ();
 sg13g2_fill_2 FILLER_4_355 ();
 sg13g2_fill_2 FILLER_4_382 ();
 sg13g2_fill_1 FILLER_4_384 ();
 sg13g2_fill_2 FILLER_4_393 ();
 sg13g2_fill_1 FILLER_4_395 ();
 sg13g2_fill_2 FILLER_4_409 ();
 sg13g2_fill_1 FILLER_4_411 ();
 sg13g2_decap_8 FILLER_4_487 ();
 sg13g2_decap_4 FILLER_4_576 ();
 sg13g2_fill_1 FILLER_4_606 ();
 sg13g2_fill_1 FILLER_4_632 ();
 sg13g2_decap_4 FILLER_4_661 ();
 sg13g2_fill_2 FILLER_4_665 ();
 sg13g2_fill_2 FILLER_4_672 ();
 sg13g2_fill_1 FILLER_4_674 ();
 sg13g2_decap_8 FILLER_4_691 ();
 sg13g2_decap_4 FILLER_4_718 ();
 sg13g2_fill_1 FILLER_4_722 ();
 sg13g2_decap_4 FILLER_4_755 ();
 sg13g2_fill_2 FILLER_4_759 ();
 sg13g2_fill_2 FILLER_4_776 ();
 sg13g2_fill_1 FILLER_4_778 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_fill_1 FILLER_5_26 ();
 sg13g2_fill_1 FILLER_5_44 ();
 sg13g2_decap_8 FILLER_5_65 ();
 sg13g2_decap_4 FILLER_5_72 ();
 sg13g2_fill_1 FILLER_5_76 ();
 sg13g2_fill_1 FILLER_5_91 ();
 sg13g2_fill_2 FILLER_5_100 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_fill_1 FILLER_5_123 ();
 sg13g2_fill_1 FILLER_5_137 ();
 sg13g2_fill_2 FILLER_5_148 ();
 sg13g2_fill_1 FILLER_5_171 ();
 sg13g2_decap_4 FILLER_5_176 ();
 sg13g2_fill_1 FILLER_5_204 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_fill_1 FILLER_5_217 ();
 sg13g2_decap_4 FILLER_5_223 ();
 sg13g2_fill_2 FILLER_5_237 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_decap_4 FILLER_5_249 ();
 sg13g2_fill_2 FILLER_5_253 ();
 sg13g2_fill_2 FILLER_5_260 ();
 sg13g2_fill_1 FILLER_5_262 ();
 sg13g2_fill_1 FILLER_5_271 ();
 sg13g2_decap_4 FILLER_5_285 ();
 sg13g2_fill_1 FILLER_5_289 ();
 sg13g2_decap_4 FILLER_5_297 ();
 sg13g2_fill_1 FILLER_5_301 ();
 sg13g2_decap_4 FILLER_5_310 ();
 sg13g2_fill_2 FILLER_5_336 ();
 sg13g2_fill_1 FILLER_5_338 ();
 sg13g2_fill_1 FILLER_5_368 ();
 sg13g2_fill_2 FILLER_5_390 ();
 sg13g2_fill_1 FILLER_5_392 ();
 sg13g2_fill_1 FILLER_5_428 ();
 sg13g2_fill_2 FILLER_5_453 ();
 sg13g2_fill_1 FILLER_5_455 ();
 sg13g2_fill_1 FILLER_5_530 ();
 sg13g2_fill_1 FILLER_5_588 ();
 sg13g2_decap_4 FILLER_5_592 ();
 sg13g2_fill_1 FILLER_5_616 ();
 sg13g2_fill_2 FILLER_5_656 ();
 sg13g2_fill_1 FILLER_5_658 ();
 sg13g2_fill_2 FILLER_5_683 ();
 sg13g2_fill_1 FILLER_5_685 ();
 sg13g2_fill_2 FILLER_5_703 ();
 sg13g2_decap_4 FILLER_5_726 ();
 sg13g2_fill_1 FILLER_5_730 ();
 sg13g2_decap_4 FILLER_5_735 ();
 sg13g2_fill_1 FILLER_5_739 ();
 sg13g2_fill_2 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_766 ();
 sg13g2_fill_2 FILLER_5_773 ();
 sg13g2_fill_1 FILLER_5_775 ();
 sg13g2_fill_2 FILLER_5_788 ();
 sg13g2_decap_4 FILLER_5_794 ();
 sg13g2_fill_2 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_14 ();
 sg13g2_fill_2 FILLER_6_25 ();
 sg13g2_fill_1 FILLER_6_58 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_fill_2 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_85 ();
 sg13g2_fill_1 FILLER_6_115 ();
 sg13g2_decap_4 FILLER_6_123 ();
 sg13g2_fill_2 FILLER_6_127 ();
 sg13g2_fill_1 FILLER_6_134 ();
 sg13g2_fill_1 FILLER_6_155 ();
 sg13g2_fill_2 FILLER_6_164 ();
 sg13g2_fill_1 FILLER_6_166 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_4 FILLER_6_189 ();
 sg13g2_fill_2 FILLER_6_197 ();
 sg13g2_fill_1 FILLER_6_199 ();
 sg13g2_fill_2 FILLER_6_222 ();
 sg13g2_fill_1 FILLER_6_246 ();
 sg13g2_decap_4 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_289 ();
 sg13g2_fill_2 FILLER_6_316 ();
 sg13g2_fill_2 FILLER_6_342 ();
 sg13g2_fill_1 FILLER_6_354 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_fill_2 FILLER_6_367 ();
 sg13g2_fill_1 FILLER_6_399 ();
 sg13g2_fill_1 FILLER_6_417 ();
 sg13g2_fill_1 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_436 ();
 sg13g2_fill_2 FILLER_6_441 ();
 sg13g2_fill_1 FILLER_6_457 ();
 sg13g2_fill_1 FILLER_6_484 ();
 sg13g2_fill_1 FILLER_6_496 ();
 sg13g2_decap_4 FILLER_6_501 ();
 sg13g2_fill_2 FILLER_6_531 ();
 sg13g2_fill_2 FILLER_6_538 ();
 sg13g2_fill_1 FILLER_6_540 ();
 sg13g2_fill_2 FILLER_6_546 ();
 sg13g2_fill_1 FILLER_6_548 ();
 sg13g2_fill_1 FILLER_6_589 ();
 sg13g2_decap_4 FILLER_6_630 ();
 sg13g2_fill_1 FILLER_6_634 ();
 sg13g2_fill_1 FILLER_6_681 ();
 sg13g2_fill_2 FILLER_6_698 ();
 sg13g2_fill_1 FILLER_6_700 ();
 sg13g2_fill_1 FILLER_6_729 ();
 sg13g2_decap_4 FILLER_6_751 ();
 sg13g2_fill_1 FILLER_6_797 ();
 sg13g2_decap_8 FILLER_6_814 ();
 sg13g2_decap_8 FILLER_6_821 ();
 sg13g2_decap_8 FILLER_6_828 ();
 sg13g2_decap_8 FILLER_6_835 ();
 sg13g2_decap_8 FILLER_6_842 ();
 sg13g2_decap_8 FILLER_6_849 ();
 sg13g2_decap_4 FILLER_6_856 ();
 sg13g2_fill_2 FILLER_6_860 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_76 ();
 sg13g2_fill_1 FILLER_7_78 ();
 sg13g2_fill_1 FILLER_7_106 ();
 sg13g2_decap_4 FILLER_7_118 ();
 sg13g2_fill_1 FILLER_7_138 ();
 sg13g2_fill_2 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_fill_1 FILLER_7_160 ();
 sg13g2_decap_4 FILLER_7_166 ();
 sg13g2_fill_2 FILLER_7_183 ();
 sg13g2_fill_2 FILLER_7_198 ();
 sg13g2_fill_1 FILLER_7_200 ();
 sg13g2_fill_2 FILLER_7_214 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_decap_4 FILLER_7_222 ();
 sg13g2_fill_1 FILLER_7_226 ();
 sg13g2_fill_2 FILLER_7_232 ();
 sg13g2_decap_4 FILLER_7_242 ();
 sg13g2_fill_2 FILLER_7_251 ();
 sg13g2_fill_2 FILLER_7_261 ();
 sg13g2_fill_1 FILLER_7_263 ();
 sg13g2_fill_1 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_fill_2 FILLER_7_336 ();
 sg13g2_fill_2 FILLER_7_362 ();
 sg13g2_fill_2 FILLER_7_383 ();
 sg13g2_fill_1 FILLER_7_385 ();
 sg13g2_fill_1 FILLER_7_412 ();
 sg13g2_fill_2 FILLER_7_447 ();
 sg13g2_fill_1 FILLER_7_453 ();
 sg13g2_fill_1 FILLER_7_507 ();
 sg13g2_fill_1 FILLER_7_529 ();
 sg13g2_fill_1 FILLER_7_550 ();
 sg13g2_fill_2 FILLER_7_559 ();
 sg13g2_fill_1 FILLER_7_561 ();
 sg13g2_fill_2 FILLER_7_604 ();
 sg13g2_fill_1 FILLER_7_606 ();
 sg13g2_decap_4 FILLER_7_622 ();
 sg13g2_decap_8 FILLER_7_692 ();
 sg13g2_decap_4 FILLER_7_699 ();
 sg13g2_fill_1 FILLER_7_703 ();
 sg13g2_fill_1 FILLER_7_713 ();
 sg13g2_fill_1 FILLER_7_718 ();
 sg13g2_fill_2 FILLER_7_744 ();
 sg13g2_fill_1 FILLER_7_746 ();
 sg13g2_decap_8 FILLER_7_752 ();
 sg13g2_fill_2 FILLER_7_763 ();
 sg13g2_decap_4 FILLER_7_772 ();
 sg13g2_decap_8 FILLER_7_786 ();
 sg13g2_fill_2 FILLER_7_793 ();
 sg13g2_fill_1 FILLER_7_795 ();
 sg13g2_decap_8 FILLER_7_817 ();
 sg13g2_decap_8 FILLER_7_824 ();
 sg13g2_decap_8 FILLER_7_831 ();
 sg13g2_decap_8 FILLER_7_838 ();
 sg13g2_decap_8 FILLER_7_845 ();
 sg13g2_decap_8 FILLER_7_852 ();
 sg13g2_fill_2 FILLER_7_859 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_40 ();
 sg13g2_fill_2 FILLER_8_106 ();
 sg13g2_fill_1 FILLER_8_108 ();
 sg13g2_decap_8 FILLER_8_118 ();
 sg13g2_decap_4 FILLER_8_125 ();
 sg13g2_fill_2 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_135 ();
 sg13g2_fill_2 FILLER_8_149 ();
 sg13g2_decap_4 FILLER_8_164 ();
 sg13g2_fill_2 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_fill_2 FILLER_8_225 ();
 sg13g2_fill_1 FILLER_8_227 ();
 sg13g2_fill_1 FILLER_8_268 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_4 FILLER_8_300 ();
 sg13g2_fill_2 FILLER_8_340 ();
 sg13g2_fill_1 FILLER_8_342 ();
 sg13g2_fill_1 FILLER_8_364 ();
 sg13g2_fill_2 FILLER_8_375 ();
 sg13g2_fill_2 FILLER_8_391 ();
 sg13g2_fill_2 FILLER_8_401 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_fill_2 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_451 ();
 sg13g2_fill_2 FILLER_8_465 ();
 sg13g2_fill_1 FILLER_8_480 ();
 sg13g2_decap_8 FILLER_8_493 ();
 sg13g2_decap_8 FILLER_8_500 ();
 sg13g2_decap_4 FILLER_8_507 ();
 sg13g2_decap_4 FILLER_8_535 ();
 sg13g2_fill_2 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_fill_2 FILLER_8_620 ();
 sg13g2_fill_2 FILLER_8_647 ();
 sg13g2_fill_1 FILLER_8_649 ();
 sg13g2_fill_2 FILLER_8_654 ();
 sg13g2_fill_1 FILLER_8_656 ();
 sg13g2_fill_1 FILLER_8_699 ();
 sg13g2_fill_2 FILLER_8_720 ();
 sg13g2_fill_1 FILLER_8_722 ();
 sg13g2_fill_1 FILLER_8_751 ();
 sg13g2_fill_2 FILLER_8_797 ();
 sg13g2_fill_2 FILLER_8_809 ();
 sg13g2_fill_2 FILLER_8_824 ();
 sg13g2_decap_8 FILLER_8_830 ();
 sg13g2_decap_8 FILLER_8_837 ();
 sg13g2_decap_8 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_851 ();
 sg13g2_decap_4 FILLER_8_858 ();
 sg13g2_fill_1 FILLER_9_26 ();
 sg13g2_fill_2 FILLER_9_74 ();
 sg13g2_fill_1 FILLER_9_76 ();
 sg13g2_fill_2 FILLER_9_119 ();
 sg13g2_fill_1 FILLER_9_132 ();
 sg13g2_fill_2 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_143 ();
 sg13g2_fill_1 FILLER_9_157 ();
 sg13g2_fill_2 FILLER_9_166 ();
 sg13g2_fill_1 FILLER_9_168 ();
 sg13g2_fill_2 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_decap_8 FILLER_9_244 ();
 sg13g2_decap_4 FILLER_9_251 ();
 sg13g2_decap_8 FILLER_9_281 ();
 sg13g2_fill_1 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_fill_2 FILLER_9_322 ();
 sg13g2_fill_1 FILLER_9_324 ();
 sg13g2_fill_2 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_fill_2 FILLER_9_347 ();
 sg13g2_fill_2 FILLER_9_365 ();
 sg13g2_fill_2 FILLER_9_385 ();
 sg13g2_fill_2 FILLER_9_403 ();
 sg13g2_fill_1 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_9_419 ();
 sg13g2_fill_2 FILLER_9_426 ();
 sg13g2_fill_1 FILLER_9_428 ();
 sg13g2_fill_1 FILLER_9_470 ();
 sg13g2_fill_2 FILLER_9_514 ();
 sg13g2_fill_1 FILLER_9_567 ();
 sg13g2_fill_1 FILLER_9_584 ();
 sg13g2_fill_2 FILLER_9_589 ();
 sg13g2_fill_2 FILLER_9_616 ();
 sg13g2_fill_2 FILLER_9_654 ();
 sg13g2_fill_1 FILLER_9_656 ();
 sg13g2_fill_2 FILLER_9_692 ();
 sg13g2_decap_8 FILLER_9_725 ();
 sg13g2_fill_2 FILLER_9_737 ();
 sg13g2_decap_8 FILLER_9_752 ();
 sg13g2_fill_1 FILLER_9_759 ();
 sg13g2_decap_4 FILLER_9_764 ();
 sg13g2_fill_1 FILLER_9_778 ();
 sg13g2_fill_2 FILLER_9_796 ();
 sg13g2_fill_1 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_845 ();
 sg13g2_decap_8 FILLER_9_852 ();
 sg13g2_fill_2 FILLER_9_859 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_fill_1 FILLER_10_86 ();
 sg13g2_fill_2 FILLER_10_99 ();
 sg13g2_fill_2 FILLER_10_135 ();
 sg13g2_fill_1 FILLER_10_142 ();
 sg13g2_fill_2 FILLER_10_163 ();
 sg13g2_fill_2 FILLER_10_195 ();
 sg13g2_fill_1 FILLER_10_197 ();
 sg13g2_fill_1 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_243 ();
 sg13g2_fill_2 FILLER_10_250 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_281 ();
 sg13g2_fill_2 FILLER_10_309 ();
 sg13g2_fill_1 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_419 ();
 sg13g2_fill_2 FILLER_10_450 ();
 sg13g2_fill_2 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_534 ();
 sg13g2_fill_2 FILLER_10_541 ();
 sg13g2_fill_1 FILLER_10_543 ();
 sg13g2_fill_2 FILLER_10_548 ();
 sg13g2_fill_1 FILLER_10_550 ();
 sg13g2_fill_1 FILLER_10_590 ();
 sg13g2_fill_2 FILLER_10_604 ();
 sg13g2_fill_1 FILLER_10_606 ();
 sg13g2_fill_2 FILLER_10_628 ();
 sg13g2_fill_1 FILLER_10_630 ();
 sg13g2_fill_1 FILLER_10_641 ();
 sg13g2_fill_2 FILLER_10_669 ();
 sg13g2_decap_4 FILLER_10_705 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_fill_2 FILLER_10_766 ();
 sg13g2_fill_2 FILLER_10_792 ();
 sg13g2_fill_1 FILLER_10_794 ();
 sg13g2_fill_1 FILLER_10_808 ();
 sg13g2_fill_1 FILLER_10_821 ();
 sg13g2_fill_1 FILLER_10_830 ();
 sg13g2_fill_2 FILLER_10_841 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_4 FILLER_10_858 ();
 sg13g2_fill_1 FILLER_11_44 ();
 sg13g2_fill_2 FILLER_11_80 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_fill_1 FILLER_11_87 ();
 sg13g2_fill_2 FILLER_11_93 ();
 sg13g2_decap_8 FILLER_11_114 ();
 sg13g2_decap_4 FILLER_11_121 ();
 sg13g2_fill_2 FILLER_11_125 ();
 sg13g2_decap_4 FILLER_11_144 ();
 sg13g2_fill_2 FILLER_11_205 ();
 sg13g2_fill_2 FILLER_11_219 ();
 sg13g2_fill_1 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_231 ();
 sg13g2_fill_1 FILLER_11_233 ();
 sg13g2_fill_1 FILLER_11_249 ();
 sg13g2_fill_1 FILLER_11_283 ();
 sg13g2_decap_8 FILLER_11_288 ();
 sg13g2_decap_8 FILLER_11_295 ();
 sg13g2_fill_2 FILLER_11_314 ();
 sg13g2_fill_1 FILLER_11_323 ();
 sg13g2_decap_8 FILLER_11_337 ();
 sg13g2_decap_4 FILLER_11_344 ();
 sg13g2_decap_4 FILLER_11_352 ();
 sg13g2_fill_1 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_430 ();
 sg13g2_fill_2 FILLER_11_437 ();
 sg13g2_fill_1 FILLER_11_443 ();
 sg13g2_decap_4 FILLER_11_449 ();
 sg13g2_decap_4 FILLER_11_475 ();
 sg13g2_decap_4 FILLER_11_510 ();
 sg13g2_decap_4 FILLER_11_539 ();
 sg13g2_decap_4 FILLER_11_598 ();
 sg13g2_fill_1 FILLER_11_602 ();
 sg13g2_fill_2 FILLER_11_629 ();
 sg13g2_fill_2 FILLER_11_634 ();
 sg13g2_decap_8 FILLER_11_701 ();
 sg13g2_fill_1 FILLER_11_708 ();
 sg13g2_fill_2 FILLER_11_715 ();
 sg13g2_decap_4 FILLER_11_726 ();
 sg13g2_fill_1 FILLER_11_730 ();
 sg13g2_decap_4 FILLER_11_777 ();
 sg13g2_fill_1 FILLER_11_790 ();
 sg13g2_decap_8 FILLER_11_799 ();
 sg13g2_decap_8 FILLER_11_806 ();
 sg13g2_fill_2 FILLER_11_813 ();
 sg13g2_fill_1 FILLER_11_815 ();
 sg13g2_fill_1 FILLER_11_828 ();
 sg13g2_fill_1 FILLER_11_834 ();
 sg13g2_fill_2 FILLER_11_843 ();
 sg13g2_decap_8 FILLER_11_853 ();
 sg13g2_fill_2 FILLER_11_860 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_11 ();
 sg13g2_fill_1 FILLER_12_25 ();
 sg13g2_fill_1 FILLER_12_57 ();
 sg13g2_fill_2 FILLER_12_93 ();
 sg13g2_fill_1 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_106 ();
 sg13g2_decap_4 FILLER_12_119 ();
 sg13g2_fill_2 FILLER_12_123 ();
 sg13g2_fill_1 FILLER_12_160 ();
 sg13g2_fill_2 FILLER_12_210 ();
 sg13g2_fill_1 FILLER_12_242 ();
 sg13g2_decap_4 FILLER_12_297 ();
 sg13g2_decap_4 FILLER_12_327 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_decap_4 FILLER_12_352 ();
 sg13g2_fill_2 FILLER_12_380 ();
 sg13g2_fill_1 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_409 ();
 sg13g2_fill_1 FILLER_12_421 ();
 sg13g2_decap_4 FILLER_12_470 ();
 sg13g2_fill_2 FILLER_12_490 ();
 sg13g2_fill_1 FILLER_12_492 ();
 sg13g2_fill_2 FILLER_12_498 ();
 sg13g2_fill_2 FILLER_12_505 ();
 sg13g2_fill_2 FILLER_12_522 ();
 sg13g2_fill_2 FILLER_12_550 ();
 sg13g2_fill_1 FILLER_12_560 ();
 sg13g2_fill_2 FILLER_12_570 ();
 sg13g2_fill_2 FILLER_12_586 ();
 sg13g2_fill_1 FILLER_12_588 ();
 sg13g2_decap_4 FILLER_12_602 ();
 sg13g2_fill_2 FILLER_12_606 ();
 sg13g2_fill_1 FILLER_12_639 ();
 sg13g2_fill_1 FILLER_12_662 ();
 sg13g2_fill_2 FILLER_12_666 ();
 sg13g2_fill_1 FILLER_12_668 ();
 sg13g2_fill_2 FILLER_12_678 ();
 sg13g2_fill_1 FILLER_12_680 ();
 sg13g2_fill_1 FILLER_12_741 ();
 sg13g2_fill_2 FILLER_12_750 ();
 sg13g2_fill_1 FILLER_12_752 ();
 sg13g2_fill_2 FILLER_12_758 ();
 sg13g2_fill_1 FILLER_12_760 ();
 sg13g2_fill_2 FILLER_12_813 ();
 sg13g2_decap_4 FILLER_12_835 ();
 sg13g2_fill_1 FILLER_12_846 ();
 sg13g2_fill_1 FILLER_12_851 ();
 sg13g2_decap_4 FILLER_12_858 ();
 sg13g2_fill_2 FILLER_13_43 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_decap_4 FILLER_13_76 ();
 sg13g2_fill_2 FILLER_13_80 ();
 sg13g2_fill_1 FILLER_13_99 ();
 sg13g2_fill_2 FILLER_13_148 ();
 sg13g2_fill_1 FILLER_13_150 ();
 sg13g2_fill_1 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_229 ();
 sg13g2_fill_2 FILLER_13_248 ();
 sg13g2_fill_1 FILLER_13_250 ();
 sg13g2_fill_2 FILLER_13_264 ();
 sg13g2_fill_2 FILLER_13_292 ();
 sg13g2_fill_2 FILLER_13_321 ();
 sg13g2_fill_1 FILLER_13_323 ();
 sg13g2_fill_2 FILLER_13_391 ();
 sg13g2_fill_1 FILLER_13_393 ();
 sg13g2_decap_4 FILLER_13_444 ();
 sg13g2_decap_4 FILLER_13_456 ();
 sg13g2_fill_2 FILLER_13_465 ();
 sg13g2_fill_1 FILLER_13_467 ();
 sg13g2_fill_2 FILLER_13_490 ();
 sg13g2_fill_1 FILLER_13_492 ();
 sg13g2_decap_8 FILLER_13_527 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_4 FILLER_13_546 ();
 sg13g2_fill_2 FILLER_13_558 ();
 sg13g2_fill_1 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_592 ();
 sg13g2_fill_1 FILLER_13_599 ();
 sg13g2_fill_1 FILLER_13_628 ();
 sg13g2_fill_1 FILLER_13_647 ();
 sg13g2_fill_2 FILLER_13_660 ();
 sg13g2_fill_1 FILLER_13_662 ();
 sg13g2_fill_2 FILLER_13_680 ();
 sg13g2_fill_1 FILLER_13_682 ();
 sg13g2_fill_2 FILLER_13_718 ();
 sg13g2_fill_2 FILLER_13_738 ();
 sg13g2_fill_2 FILLER_13_758 ();
 sg13g2_decap_4 FILLER_13_783 ();
 sg13g2_fill_2 FILLER_13_787 ();
 sg13g2_fill_2 FILLER_13_794 ();
 sg13g2_decap_4 FILLER_13_809 ();
 sg13g2_fill_1 FILLER_13_813 ();
 sg13g2_fill_1 FILLER_13_835 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_33 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_fill_2 FILLER_14_111 ();
 sg13g2_fill_1 FILLER_14_113 ();
 sg13g2_fill_2 FILLER_14_118 ();
 sg13g2_fill_2 FILLER_14_128 ();
 sg13g2_decap_4 FILLER_14_155 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_209 ();
 sg13g2_fill_2 FILLER_14_223 ();
 sg13g2_fill_1 FILLER_14_225 ();
 sg13g2_fill_2 FILLER_14_240 ();
 sg13g2_fill_1 FILLER_14_242 ();
 sg13g2_fill_2 FILLER_14_264 ();
 sg13g2_fill_1 FILLER_14_266 ();
 sg13g2_decap_4 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_fill_2 FILLER_14_331 ();
 sg13g2_fill_1 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_fill_1 FILLER_14_364 ();
 sg13g2_fill_2 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_410 ();
 sg13g2_decap_8 FILLER_14_417 ();
 sg13g2_decap_8 FILLER_14_424 ();
 sg13g2_fill_2 FILLER_14_431 ();
 sg13g2_fill_2 FILLER_14_465 ();
 sg13g2_fill_1 FILLER_14_467 ();
 sg13g2_fill_1 FILLER_14_506 ();
 sg13g2_fill_1 FILLER_14_523 ();
 sg13g2_fill_1 FILLER_14_565 ();
 sg13g2_fill_2 FILLER_14_578 ();
 sg13g2_fill_1 FILLER_14_606 ();
 sg13g2_fill_2 FILLER_14_620 ();
 sg13g2_fill_2 FILLER_14_656 ();
 sg13g2_fill_2 FILLER_14_692 ();
 sg13g2_decap_8 FILLER_14_737 ();
 sg13g2_fill_2 FILLER_14_744 ();
 sg13g2_decap_4 FILLER_14_754 ();
 sg13g2_fill_1 FILLER_14_767 ();
 sg13g2_fill_1 FILLER_14_773 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_4 FILLER_14_805 ();
 sg13g2_fill_2 FILLER_14_809 ();
 sg13g2_fill_1 FILLER_14_821 ();
 sg13g2_fill_2 FILLER_15_55 ();
 sg13g2_fill_1 FILLER_15_57 ();
 sg13g2_fill_1 FILLER_15_79 ();
 sg13g2_decap_8 FILLER_15_143 ();
 sg13g2_decap_4 FILLER_15_150 ();
 sg13g2_fill_2 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_179 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_2 FILLER_15_248 ();
 sg13g2_fill_1 FILLER_15_250 ();
 sg13g2_fill_1 FILLER_15_263 ();
 sg13g2_fill_2 FILLER_15_269 ();
 sg13g2_fill_2 FILLER_15_296 ();
 sg13g2_fill_1 FILLER_15_298 ();
 sg13g2_fill_1 FILLER_15_312 ();
 sg13g2_fill_2 FILLER_15_346 ();
 sg13g2_fill_2 FILLER_15_359 ();
 sg13g2_fill_1 FILLER_15_361 ();
 sg13g2_decap_4 FILLER_15_390 ();
 sg13g2_decap_4 FILLER_15_422 ();
 sg13g2_fill_2 FILLER_15_426 ();
 sg13g2_fill_2 FILLER_15_452 ();
 sg13g2_fill_2 FILLER_15_508 ();
 sg13g2_fill_1 FILLER_15_515 ();
 sg13g2_fill_1 FILLER_15_521 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_fill_2 FILLER_15_599 ();
 sg13g2_fill_1 FILLER_15_601 ();
 sg13g2_fill_2 FILLER_15_611 ();
 sg13g2_fill_1 FILLER_15_635 ();
 sg13g2_fill_2 FILLER_15_692 ();
 sg13g2_fill_1 FILLER_15_694 ();
 sg13g2_fill_1 FILLER_15_759 ();
 sg13g2_fill_2 FILLER_15_775 ();
 sg13g2_fill_1 FILLER_15_777 ();
 sg13g2_fill_1 FILLER_15_812 ();
 sg13g2_fill_2 FILLER_15_825 ();
 sg13g2_fill_1 FILLER_15_827 ();
 sg13g2_fill_2 FILLER_15_860 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_1 FILLER_16_25 ();
 sg13g2_fill_2 FILLER_16_34 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_62 ();
 sg13g2_fill_1 FILLER_16_96 ();
 sg13g2_decap_4 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_198 ();
 sg13g2_fill_1 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_decap_4 FILLER_16_225 ();
 sg13g2_fill_1 FILLER_16_229 ();
 sg13g2_decap_4 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_243 ();
 sg13g2_fill_2 FILLER_16_262 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_fill_1 FILLER_16_281 ();
 sg13g2_fill_1 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_297 ();
 sg13g2_decap_4 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_332 ();
 sg13g2_fill_2 FILLER_16_351 ();
 sg13g2_fill_1 FILLER_16_381 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_2 FILLER_16_418 ();
 sg13g2_fill_1 FILLER_16_420 ();
 sg13g2_fill_1 FILLER_16_464 ();
 sg13g2_fill_1 FILLER_16_491 ();
 sg13g2_fill_2 FILLER_16_504 ();
 sg13g2_fill_2 FILLER_16_585 ();
 sg13g2_fill_1 FILLER_16_587 ();
 sg13g2_fill_2 FILLER_16_627 ();
 sg13g2_fill_1 FILLER_16_634 ();
 sg13g2_fill_2 FILLER_16_648 ();
 sg13g2_fill_1 FILLER_16_661 ();
 sg13g2_decap_4 FILLER_16_692 ();
 sg13g2_fill_2 FILLER_16_704 ();
 sg13g2_fill_2 FILLER_16_710 ();
 sg13g2_fill_2 FILLER_16_730 ();
 sg13g2_fill_1 FILLER_16_743 ();
 sg13g2_decap_8 FILLER_16_761 ();
 sg13g2_decap_4 FILLER_16_768 ();
 sg13g2_fill_1 FILLER_16_772 ();
 sg13g2_fill_1 FILLER_16_812 ();
 sg13g2_fill_2 FILLER_16_834 ();
 sg13g2_fill_2 FILLER_17_26 ();
 sg13g2_fill_2 FILLER_17_55 ();
 sg13g2_fill_1 FILLER_17_57 ();
 sg13g2_fill_2 FILLER_17_68 ();
 sg13g2_fill_1 FILLER_17_74 ();
 sg13g2_fill_2 FILLER_17_132 ();
 sg13g2_fill_1 FILLER_17_139 ();
 sg13g2_fill_2 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_155 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_fill_2 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_fill_2 FILLER_17_334 ();
 sg13g2_fill_1 FILLER_17_336 ();
 sg13g2_fill_2 FILLER_17_359 ();
 sg13g2_decap_4 FILLER_17_373 ();
 sg13g2_decap_4 FILLER_17_385 ();
 sg13g2_fill_2 FILLER_17_398 ();
 sg13g2_fill_1 FILLER_17_400 ();
 sg13g2_fill_1 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_411 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_4 FILLER_17_427 ();
 sg13g2_fill_2 FILLER_17_431 ();
 sg13g2_fill_1 FILLER_17_454 ();
 sg13g2_fill_2 FILLER_17_464 ();
 sg13g2_fill_1 FILLER_17_466 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_fill_2 FILLER_17_492 ();
 sg13g2_fill_1 FILLER_17_494 ();
 sg13g2_decap_4 FILLER_17_540 ();
 sg13g2_fill_2 FILLER_17_548 ();
 sg13g2_fill_2 FILLER_17_555 ();
 sg13g2_decap_4 FILLER_17_562 ();
 sg13g2_fill_2 FILLER_17_579 ();
 sg13g2_fill_1 FILLER_17_581 ();
 sg13g2_fill_1 FILLER_17_594 ();
 sg13g2_decap_4 FILLER_17_600 ();
 sg13g2_fill_2 FILLER_17_604 ();
 sg13g2_fill_2 FILLER_17_626 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_fill_2 FILLER_17_663 ();
 sg13g2_fill_2 FILLER_17_692 ();
 sg13g2_decap_4 FILLER_17_699 ();
 sg13g2_fill_1 FILLER_17_703 ();
 sg13g2_fill_1 FILLER_17_720 ();
 sg13g2_fill_1 FILLER_17_733 ();
 sg13g2_fill_2 FILLER_17_772 ();
 sg13g2_fill_1 FILLER_17_774 ();
 sg13g2_decap_4 FILLER_17_806 ();
 sg13g2_fill_2 FILLER_17_813 ();
 sg13g2_fill_1 FILLER_17_852 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_24 ();
 sg13g2_fill_1 FILLER_18_44 ();
 sg13g2_fill_2 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_155 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_fill_2 FILLER_18_199 ();
 sg13g2_fill_1 FILLER_18_201 ();
 sg13g2_fill_1 FILLER_18_212 ();
 sg13g2_fill_1 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_291 ();
 sg13g2_fill_2 FILLER_18_300 ();
 sg13g2_fill_2 FILLER_18_318 ();
 sg13g2_fill_1 FILLER_18_320 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_fill_2 FILLER_18_386 ();
 sg13g2_fill_2 FILLER_18_420 ();
 sg13g2_fill_1 FILLER_18_422 ();
 sg13g2_fill_2 FILLER_18_454 ();
 sg13g2_fill_1 FILLER_18_456 ();
 sg13g2_decap_4 FILLER_18_518 ();
 sg13g2_fill_2 FILLER_18_530 ();
 sg13g2_decap_8 FILLER_18_568 ();
 sg13g2_decap_4 FILLER_18_595 ();
 sg13g2_fill_1 FILLER_18_611 ();
 sg13g2_fill_1 FILLER_18_634 ();
 sg13g2_fill_2 FILLER_18_678 ();
 sg13g2_fill_2 FILLER_18_705 ();
 sg13g2_fill_1 FILLER_18_707 ();
 sg13g2_fill_1 FILLER_18_718 ();
 sg13g2_fill_2 FILLER_18_739 ();
 sg13g2_fill_2 FILLER_18_782 ();
 sg13g2_fill_1 FILLER_18_835 ();
 sg13g2_fill_2 FILLER_19_26 ();
 sg13g2_fill_2 FILLER_19_42 ();
 sg13g2_fill_2 FILLER_19_96 ();
 sg13g2_fill_1 FILLER_19_125 ();
 sg13g2_fill_1 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_206 ();
 sg13g2_decap_4 FILLER_19_215 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_decap_4 FILLER_19_256 ();
 sg13g2_fill_2 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_277 ();
 sg13g2_fill_2 FILLER_19_302 ();
 sg13g2_fill_2 FILLER_19_312 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_decap_4 FILLER_19_323 ();
 sg13g2_fill_1 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_fill_1 FILLER_19_340 ();
 sg13g2_fill_2 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_4 FILLER_19_390 ();
 sg13g2_fill_2 FILLER_19_402 ();
 sg13g2_fill_2 FILLER_19_416 ();
 sg13g2_decap_4 FILLER_19_426 ();
 sg13g2_fill_1 FILLER_19_430 ();
 sg13g2_decap_8 FILLER_19_439 ();
 sg13g2_decap_4 FILLER_19_446 ();
 sg13g2_fill_1 FILLER_19_450 ();
 sg13g2_decap_4 FILLER_19_461 ();
 sg13g2_decap_8 FILLER_19_474 ();
 sg13g2_decap_4 FILLER_19_484 ();
 sg13g2_fill_2 FILLER_19_488 ();
 sg13g2_fill_2 FILLER_19_498 ();
 sg13g2_fill_1 FILLER_19_512 ();
 sg13g2_decap_4 FILLER_19_551 ();
 sg13g2_fill_2 FILLER_19_555 ();
 sg13g2_fill_2 FILLER_19_563 ();
 sg13g2_fill_2 FILLER_19_568 ();
 sg13g2_fill_1 FILLER_19_570 ();
 sg13g2_fill_1 FILLER_19_580 ();
 sg13g2_fill_1 FILLER_19_586 ();
 sg13g2_fill_2 FILLER_19_612 ();
 sg13g2_fill_1 FILLER_19_614 ();
 sg13g2_fill_2 FILLER_19_628 ();
 sg13g2_fill_2 FILLER_19_673 ();
 sg13g2_decap_4 FILLER_19_684 ();
 sg13g2_fill_1 FILLER_19_733 ();
 sg13g2_fill_1 FILLER_19_755 ();
 sg13g2_fill_1 FILLER_19_760 ();
 sg13g2_fill_2 FILLER_19_773 ();
 sg13g2_fill_2 FILLER_19_794 ();
 sg13g2_fill_1 FILLER_19_829 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_9 ();
 sg13g2_fill_1 FILLER_20_27 ();
 sg13g2_fill_2 FILLER_20_44 ();
 sg13g2_fill_2 FILLER_20_65 ();
 sg13g2_fill_1 FILLER_20_67 ();
 sg13g2_fill_2 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_74 ();
 sg13g2_fill_2 FILLER_20_78 ();
 sg13g2_fill_2 FILLER_20_102 ();
 sg13g2_fill_2 FILLER_20_118 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_139 ();
 sg13g2_fill_2 FILLER_20_145 ();
 sg13g2_fill_1 FILLER_20_166 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_239 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_fill_1 FILLER_20_322 ();
 sg13g2_fill_1 FILLER_20_339 ();
 sg13g2_fill_2 FILLER_20_350 ();
 sg13g2_decap_4 FILLER_20_361 ();
 sg13g2_fill_2 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_370 ();
 sg13g2_fill_2 FILLER_20_393 ();
 sg13g2_fill_1 FILLER_20_395 ();
 sg13g2_fill_1 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_fill_2 FILLER_20_441 ();
 sg13g2_fill_2 FILLER_20_498 ();
 sg13g2_fill_1 FILLER_20_500 ();
 sg13g2_fill_2 FILLER_20_515 ();
 sg13g2_decap_4 FILLER_20_540 ();
 sg13g2_fill_2 FILLER_20_553 ();
 sg13g2_fill_1 FILLER_20_563 ();
 sg13g2_fill_2 FILLER_20_572 ();
 sg13g2_fill_1 FILLER_20_574 ();
 sg13g2_fill_1 FILLER_20_591 ();
 sg13g2_decap_4 FILLER_20_595 ();
 sg13g2_fill_2 FILLER_20_599 ();
 sg13g2_fill_2 FILLER_20_710 ();
 sg13g2_fill_1 FILLER_20_721 ();
 sg13g2_fill_2 FILLER_20_749 ();
 sg13g2_fill_1 FILLER_20_751 ();
 sg13g2_fill_1 FILLER_20_762 ();
 sg13g2_decap_8 FILLER_20_772 ();
 sg13g2_fill_2 FILLER_20_784 ();
 sg13g2_fill_1 FILLER_20_808 ();
 sg13g2_fill_1 FILLER_20_835 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_fill_2 FILLER_21_52 ();
 sg13g2_fill_1 FILLER_21_54 ();
 sg13g2_fill_1 FILLER_21_114 ();
 sg13g2_fill_2 FILLER_21_157 ();
 sg13g2_fill_2 FILLER_21_172 ();
 sg13g2_decap_4 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_224 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_decap_4 FILLER_21_253 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_decap_8 FILLER_21_269 ();
 sg13g2_decap_4 FILLER_21_276 ();
 sg13g2_decap_4 FILLER_21_306 ();
 sg13g2_fill_1 FILLER_21_341 ();
 sg13g2_fill_2 FILLER_21_346 ();
 sg13g2_fill_1 FILLER_21_348 ();
 sg13g2_fill_2 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_4 FILLER_21_394 ();
 sg13g2_fill_2 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_21_412 ();
 sg13g2_fill_2 FILLER_21_419 ();
 sg13g2_decap_4 FILLER_21_441 ();
 sg13g2_fill_1 FILLER_21_453 ();
 sg13g2_decap_8 FILLER_21_464 ();
 sg13g2_fill_2 FILLER_21_474 ();
 sg13g2_fill_1 FILLER_21_476 ();
 sg13g2_decap_4 FILLER_21_528 ();
 sg13g2_fill_1 FILLER_21_545 ();
 sg13g2_fill_2 FILLER_21_559 ();
 sg13g2_fill_1 FILLER_21_561 ();
 sg13g2_fill_1 FILLER_21_569 ();
 sg13g2_fill_2 FILLER_21_582 ();
 sg13g2_fill_2 FILLER_21_602 ();
 sg13g2_fill_1 FILLER_21_604 ();
 sg13g2_fill_2 FILLER_21_630 ();
 sg13g2_fill_1 FILLER_21_632 ();
 sg13g2_fill_2 FILLER_21_651 ();
 sg13g2_fill_1 FILLER_21_674 ();
 sg13g2_fill_2 FILLER_21_705 ();
 sg13g2_fill_1 FILLER_21_707 ();
 sg13g2_fill_2 FILLER_21_738 ();
 sg13g2_fill_2 FILLER_21_772 ();
 sg13g2_fill_2 FILLER_21_796 ();
 sg13g2_fill_1 FILLER_21_810 ();
 sg13g2_fill_1 FILLER_21_851 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_fill_2 FILLER_22_61 ();
 sg13g2_fill_2 FILLER_22_75 ();
 sg13g2_decap_8 FILLER_22_87 ();
 sg13g2_decap_4 FILLER_22_94 ();
 sg13g2_fill_2 FILLER_22_98 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_decap_4 FILLER_22_180 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_195 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_203 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_232 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_257 ();
 sg13g2_fill_2 FILLER_22_263 ();
 sg13g2_fill_1 FILLER_22_265 ();
 sg13g2_fill_1 FILLER_22_276 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_fill_2 FILLER_22_327 ();
 sg13g2_fill_1 FILLER_22_337 ();
 sg13g2_decap_4 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_367 ();
 sg13g2_fill_2 FILLER_22_418 ();
 sg13g2_decap_4 FILLER_22_425 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_fill_2 FILLER_22_464 ();
 sg13g2_fill_2 FILLER_22_476 ();
 sg13g2_fill_1 FILLER_22_526 ();
 sg13g2_decap_4 FILLER_22_540 ();
 sg13g2_fill_2 FILLER_22_544 ();
 sg13g2_fill_2 FILLER_22_563 ();
 sg13g2_fill_1 FILLER_22_565 ();
 sg13g2_fill_1 FILLER_22_581 ();
 sg13g2_fill_2 FILLER_22_597 ();
 sg13g2_fill_2 FILLER_22_630 ();
 sg13g2_fill_2 FILLER_22_648 ();
 sg13g2_fill_1 FILLER_22_692 ();
 sg13g2_fill_2 FILLER_22_728 ();
 sg13g2_fill_1 FILLER_22_810 ();
 sg13g2_fill_2 FILLER_22_834 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_20 ();
 sg13g2_fill_1 FILLER_23_22 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_30 ();
 sg13g2_fill_1 FILLER_23_57 ();
 sg13g2_fill_1 FILLER_23_62 ();
 sg13g2_decap_8 FILLER_23_92 ();
 sg13g2_decap_8 FILLER_23_99 ();
 sg13g2_decap_4 FILLER_23_106 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_decap_4 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_decap_4 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_decap_4 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_269 ();
 sg13g2_fill_2 FILLER_23_278 ();
 sg13g2_fill_2 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_318 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_4 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_fill_2 FILLER_23_397 ();
 sg13g2_fill_1 FILLER_23_399 ();
 sg13g2_decap_4 FILLER_23_410 ();
 sg13g2_fill_1 FILLER_23_414 ();
 sg13g2_fill_1 FILLER_23_444 ();
 sg13g2_fill_2 FILLER_23_466 ();
 sg13g2_fill_1 FILLER_23_468 ();
 sg13g2_fill_2 FILLER_23_495 ();
 sg13g2_fill_1 FILLER_23_497 ();
 sg13g2_fill_2 FILLER_23_502 ();
 sg13g2_fill_1 FILLER_23_509 ();
 sg13g2_fill_2 FILLER_23_526 ();
 sg13g2_decap_8 FILLER_23_533 ();
 sg13g2_fill_2 FILLER_23_540 ();
 sg13g2_fill_1 FILLER_23_542 ();
 sg13g2_fill_1 FILLER_23_548 ();
 sg13g2_fill_2 FILLER_23_595 ();
 sg13g2_fill_1 FILLER_23_597 ();
 sg13g2_fill_2 FILLER_23_621 ();
 sg13g2_fill_1 FILLER_23_623 ();
 sg13g2_fill_2 FILLER_23_633 ();
 sg13g2_fill_1 FILLER_23_635 ();
 sg13g2_fill_2 FILLER_23_715 ();
 sg13g2_fill_1 FILLER_23_722 ();
 sg13g2_fill_1 FILLER_23_794 ();
 sg13g2_fill_2 FILLER_23_799 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_2 FILLER_24_23 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_121 ();
 sg13g2_fill_1 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_196 ();
 sg13g2_fill_2 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_204 ();
 sg13g2_decap_4 FILLER_24_219 ();
 sg13g2_decap_8 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_234 ();
 sg13g2_fill_2 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_248 ();
 sg13g2_fill_2 FILLER_24_262 ();
 sg13g2_fill_2 FILLER_24_272 ();
 sg13g2_fill_2 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_fill_2 FILLER_24_339 ();
 sg13g2_fill_2 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_24_379 ();
 sg13g2_fill_1 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_fill_1 FILLER_24_423 ();
 sg13g2_fill_2 FILLER_24_429 ();
 sg13g2_decap_4 FILLER_24_434 ();
 sg13g2_fill_1 FILLER_24_438 ();
 sg13g2_fill_1 FILLER_24_444 ();
 sg13g2_fill_2 FILLER_24_450 ();
 sg13g2_fill_1 FILLER_24_452 ();
 sg13g2_fill_1 FILLER_24_458 ();
 sg13g2_fill_2 FILLER_24_464 ();
 sg13g2_fill_1 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_472 ();
 sg13g2_fill_1 FILLER_24_479 ();
 sg13g2_fill_2 FILLER_24_484 ();
 sg13g2_fill_1 FILLER_24_489 ();
 sg13g2_decap_4 FILLER_24_499 ();
 sg13g2_fill_1 FILLER_24_503 ();
 sg13g2_fill_1 FILLER_24_526 ();
 sg13g2_decap_8 FILLER_24_566 ();
 sg13g2_fill_2 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_594 ();
 sg13g2_fill_2 FILLER_24_601 ();
 sg13g2_fill_1 FILLER_24_603 ();
 sg13g2_fill_2 FILLER_24_627 ();
 sg13g2_fill_1 FILLER_24_629 ();
 sg13g2_fill_2 FILLER_24_650 ();
 sg13g2_fill_2 FILLER_24_660 ();
 sg13g2_fill_1 FILLER_24_669 ();
 sg13g2_fill_2 FILLER_24_687 ();
 sg13g2_fill_1 FILLER_24_689 ();
 sg13g2_fill_2 FILLER_24_704 ();
 sg13g2_fill_1 FILLER_24_706 ();
 sg13g2_fill_1 FILLER_24_794 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_9 ();
 sg13g2_fill_2 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_50 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_79 ();
 sg13g2_fill_1 FILLER_25_81 ();
 sg13g2_fill_2 FILLER_25_92 ();
 sg13g2_fill_1 FILLER_25_120 ();
 sg13g2_fill_2 FILLER_25_164 ();
 sg13g2_fill_1 FILLER_25_166 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_fill_2 FILLER_25_285 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_fill_1 FILLER_25_371 ();
 sg13g2_fill_1 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_399 ();
 sg13g2_fill_1 FILLER_25_412 ();
 sg13g2_decap_4 FILLER_25_437 ();
 sg13g2_fill_1 FILLER_25_441 ();
 sg13g2_fill_2 FILLER_25_450 ();
 sg13g2_fill_1 FILLER_25_460 ();
 sg13g2_fill_2 FILLER_25_477 ();
 sg13g2_fill_1 FILLER_25_499 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_fill_1 FILLER_25_532 ();
 sg13g2_fill_1 FILLER_25_540 ();
 sg13g2_decap_4 FILLER_25_554 ();
 sg13g2_fill_2 FILLER_25_558 ();
 sg13g2_decap_8 FILLER_25_576 ();
 sg13g2_fill_2 FILLER_25_609 ();
 sg13g2_fill_1 FILLER_25_632 ();
 sg13g2_fill_2 FILLER_25_761 ();
 sg13g2_fill_2 FILLER_25_776 ();
 sg13g2_fill_2 FILLER_25_783 ();
 sg13g2_fill_1 FILLER_25_789 ();
 sg13g2_fill_1 FILLER_25_795 ();
 sg13g2_fill_2 FILLER_25_800 ();
 sg13g2_fill_1 FILLER_25_852 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_fill_1 FILLER_26_62 ();
 sg13g2_fill_1 FILLER_26_76 ();
 sg13g2_decap_4 FILLER_26_117 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_decap_4 FILLER_26_199 ();
 sg13g2_fill_2 FILLER_26_208 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_318 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_fill_2 FILLER_26_354 ();
 sg13g2_fill_1 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_fill_2 FILLER_26_397 ();
 sg13g2_fill_1 FILLER_26_420 ();
 sg13g2_decap_4 FILLER_26_433 ();
 sg13g2_decap_8 FILLER_26_459 ();
 sg13g2_decap_4 FILLER_26_466 ();
 sg13g2_fill_2 FILLER_26_470 ();
 sg13g2_decap_8 FILLER_26_499 ();
 sg13g2_fill_1 FILLER_26_506 ();
 sg13g2_decap_8 FILLER_26_517 ();
 sg13g2_decap_8 FILLER_26_524 ();
 sg13g2_decap_4 FILLER_26_531 ();
 sg13g2_fill_2 FILLER_26_553 ();
 sg13g2_fill_1 FILLER_26_566 ();
 sg13g2_fill_2 FILLER_26_583 ();
 sg13g2_fill_2 FILLER_26_592 ();
 sg13g2_fill_1 FILLER_26_652 ();
 sg13g2_fill_2 FILLER_26_657 ();
 sg13g2_fill_1 FILLER_26_677 ();
 sg13g2_fill_2 FILLER_26_687 ();
 sg13g2_fill_1 FILLER_26_701 ();
 sg13g2_fill_2 FILLER_26_721 ();
 sg13g2_fill_1 FILLER_26_749 ();
 sg13g2_fill_2 FILLER_26_834 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_51 ();
 sg13g2_fill_2 FILLER_27_67 ();
 sg13g2_fill_2 FILLER_27_85 ();
 sg13g2_decap_4 FILLER_27_102 ();
 sg13g2_fill_1 FILLER_27_106 ();
 sg13g2_fill_2 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_decap_4 FILLER_27_141 ();
 sg13g2_fill_2 FILLER_27_145 ();
 sg13g2_fill_2 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_fill_2 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_164 ();
 sg13g2_decap_4 FILLER_27_171 ();
 sg13g2_fill_2 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_decap_4 FILLER_27_217 ();
 sg13g2_fill_2 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_fill_1 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_decap_4 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_fill_2 FILLER_27_354 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_fill_1 FILLER_27_401 ();
 sg13g2_decap_4 FILLER_27_428 ();
 sg13g2_fill_1 FILLER_27_432 ();
 sg13g2_fill_2 FILLER_27_438 ();
 sg13g2_fill_1 FILLER_27_440 ();
 sg13g2_fill_2 FILLER_27_484 ();
 sg13g2_fill_2 FILLER_27_500 ();
 sg13g2_fill_1 FILLER_27_502 ();
 sg13g2_fill_2 FILLER_27_508 ();
 sg13g2_fill_1 FILLER_27_510 ();
 sg13g2_fill_2 FILLER_27_532 ();
 sg13g2_fill_2 FILLER_27_549 ();
 sg13g2_fill_1 FILLER_27_559 ();
 sg13g2_fill_2 FILLER_27_575 ();
 sg13g2_fill_1 FILLER_27_612 ();
 sg13g2_fill_2 FILLER_27_631 ();
 sg13g2_fill_1 FILLER_27_670 ();
 sg13g2_fill_2 FILLER_27_696 ();
 sg13g2_fill_2 FILLER_27_748 ();
 sg13g2_decap_8 FILLER_27_779 ();
 sg13g2_decap_4 FILLER_27_786 ();
 sg13g2_fill_1 FILLER_27_790 ();
 sg13g2_decap_4 FILLER_27_795 ();
 sg13g2_fill_2 FILLER_27_804 ();
 sg13g2_fill_2 FILLER_27_826 ();
 sg13g2_fill_2 FILLER_28_26 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_108 ();
 sg13g2_decap_4 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_183 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_decap_4 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_fill_2 FILLER_28_237 ();
 sg13g2_fill_1 FILLER_28_239 ();
 sg13g2_decap_4 FILLER_28_267 ();
 sg13g2_decap_8 FILLER_28_320 ();
 sg13g2_fill_2 FILLER_28_327 ();
 sg13g2_fill_1 FILLER_28_329 ();
 sg13g2_fill_2 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_4 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_361 ();
 sg13g2_fill_2 FILLER_28_372 ();
 sg13g2_fill_1 FILLER_28_379 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_4 FILLER_28_442 ();
 sg13g2_fill_1 FILLER_28_446 ();
 sg13g2_decap_8 FILLER_28_456 ();
 sg13g2_fill_2 FILLER_28_463 ();
 sg13g2_fill_1 FILLER_28_465 ();
 sg13g2_decap_4 FILLER_28_483 ();
 sg13g2_decap_4 FILLER_28_497 ();
 sg13g2_fill_1 FILLER_28_501 ();
 sg13g2_fill_1 FILLER_28_516 ();
 sg13g2_fill_1 FILLER_28_528 ();
 sg13g2_fill_1 FILLER_28_538 ();
 sg13g2_fill_1 FILLER_28_583 ();
 sg13g2_fill_1 FILLER_28_588 ();
 sg13g2_fill_2 FILLER_28_597 ();
 sg13g2_fill_2 FILLER_28_634 ();
 sg13g2_fill_2 FILLER_28_651 ();
 sg13g2_fill_1 FILLER_28_653 ();
 sg13g2_fill_1 FILLER_28_658 ();
 sg13g2_fill_2 FILLER_28_679 ();
 sg13g2_fill_2 FILLER_28_719 ();
 sg13g2_fill_2 FILLER_28_752 ();
 sg13g2_fill_2 FILLER_28_768 ();
 sg13g2_decap_4 FILLER_28_783 ();
 sg13g2_fill_1 FILLER_28_787 ();
 sg13g2_fill_1 FILLER_28_811 ();
 sg13g2_fill_2 FILLER_28_848 ();
 sg13g2_fill_2 FILLER_28_859 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_85 ();
 sg13g2_decap_4 FILLER_29_137 ();
 sg13g2_fill_2 FILLER_29_186 ();
 sg13g2_fill_2 FILLER_29_207 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_232 ();
 sg13g2_decap_4 FILLER_29_301 ();
 sg13g2_fill_2 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_4 FILLER_29_376 ();
 sg13g2_fill_1 FILLER_29_380 ();
 sg13g2_decap_4 FILLER_29_412 ();
 sg13g2_fill_2 FILLER_29_425 ();
 sg13g2_fill_2 FILLER_29_440 ();
 sg13g2_decap_8 FILLER_29_463 ();
 sg13g2_fill_2 FILLER_29_483 ();
 sg13g2_fill_1 FILLER_29_485 ();
 sg13g2_fill_1 FILLER_29_563 ();
 sg13g2_fill_1 FILLER_29_572 ();
 sg13g2_fill_2 FILLER_29_599 ();
 sg13g2_fill_2 FILLER_29_685 ();
 sg13g2_fill_1 FILLER_29_742 ();
 sg13g2_fill_2 FILLER_29_769 ();
 sg13g2_fill_2 FILLER_29_791 ();
 sg13g2_fill_1 FILLER_29_793 ();
 sg13g2_fill_2 FILLER_29_798 ();
 sg13g2_fill_1 FILLER_29_828 ();
 sg13g2_fill_1 FILLER_29_850 ();
 sg13g2_fill_2 FILLER_29_859 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_7 ();
 sg13g2_fill_2 FILLER_30_32 ();
 sg13g2_fill_1 FILLER_30_34 ();
 sg13g2_fill_2 FILLER_30_118 ();
 sg13g2_fill_2 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_131 ();
 sg13g2_fill_1 FILLER_30_145 ();
 sg13g2_fill_1 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_219 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_fill_2 FILLER_30_282 ();
 sg13g2_fill_2 FILLER_30_302 ();
 sg13g2_fill_2 FILLER_30_330 ();
 sg13g2_decap_4 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_364 ();
 sg13g2_fill_1 FILLER_30_366 ();
 sg13g2_decap_4 FILLER_30_395 ();
 sg13g2_fill_2 FILLER_30_459 ();
 sg13g2_fill_1 FILLER_30_461 ();
 sg13g2_fill_1 FILLER_30_487 ();
 sg13g2_fill_2 FILLER_30_496 ();
 sg13g2_fill_1 FILLER_30_498 ();
 sg13g2_fill_2 FILLER_30_532 ();
 sg13g2_fill_2 FILLER_30_542 ();
 sg13g2_fill_2 FILLER_30_573 ();
 sg13g2_fill_2 FILLER_30_579 ();
 sg13g2_fill_1 FILLER_30_585 ();
 sg13g2_fill_1 FILLER_30_647 ();
 sg13g2_fill_1 FILLER_30_653 ();
 sg13g2_fill_1 FILLER_30_690 ();
 sg13g2_fill_1 FILLER_30_721 ();
 sg13g2_fill_1 FILLER_30_731 ();
 sg13g2_fill_1 FILLER_30_758 ();
 sg13g2_fill_1 FILLER_30_767 ();
 sg13g2_fill_1 FILLER_30_798 ();
 sg13g2_fill_2 FILLER_31_90 ();
 sg13g2_fill_1 FILLER_31_92 ();
 sg13g2_fill_2 FILLER_31_106 ();
 sg13g2_fill_2 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_131 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_244 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_fill_2 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_282 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_decap_8 FILLER_31_382 ();
 sg13g2_fill_1 FILLER_31_389 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_31_419 ();
 sg13g2_fill_1 FILLER_31_421 ();
 sg13g2_decap_4 FILLER_31_443 ();
 sg13g2_fill_1 FILLER_31_447 ();
 sg13g2_fill_1 FILLER_31_456 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_fill_1 FILLER_31_469 ();
 sg13g2_fill_2 FILLER_31_476 ();
 sg13g2_fill_2 FILLER_31_491 ();
 sg13g2_fill_1 FILLER_31_510 ();
 sg13g2_fill_1 FILLER_31_516 ();
 sg13g2_fill_1 FILLER_31_545 ();
 sg13g2_fill_1 FILLER_31_561 ();
 sg13g2_fill_2 FILLER_31_659 ();
 sg13g2_fill_1 FILLER_31_661 ();
 sg13g2_fill_1 FILLER_31_675 ();
 sg13g2_fill_1 FILLER_31_696 ();
 sg13g2_fill_1 FILLER_31_770 ();
 sg13g2_fill_1 FILLER_31_784 ();
 sg13g2_fill_1 FILLER_31_819 ();
 sg13g2_fill_1 FILLER_31_828 ();
 sg13g2_fill_1 FILLER_31_834 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_18 ();
 sg13g2_fill_2 FILLER_32_43 ();
 sg13g2_fill_1 FILLER_32_45 ();
 sg13g2_fill_2 FILLER_32_76 ();
 sg13g2_fill_1 FILLER_32_88 ();
 sg13g2_decap_4 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_101 ();
 sg13g2_fill_2 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_136 ();
 sg13g2_decap_8 FILLER_32_153 ();
 sg13g2_decap_4 FILLER_32_160 ();
 sg13g2_fill_1 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_fill_2 FILLER_32_208 ();
 sg13g2_decap_8 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_230 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_decap_4 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_310 ();
 sg13g2_fill_2 FILLER_32_341 ();
 sg13g2_decap_4 FILLER_32_363 ();
 sg13g2_fill_2 FILLER_32_384 ();
 sg13g2_fill_1 FILLER_32_386 ();
 sg13g2_fill_1 FILLER_32_413 ();
 sg13g2_fill_2 FILLER_32_440 ();
 sg13g2_fill_1 FILLER_32_442 ();
 sg13g2_decap_4 FILLER_32_455 ();
 sg13g2_decap_4 FILLER_32_466 ();
 sg13g2_fill_2 FILLER_32_470 ();
 sg13g2_fill_1 FILLER_32_487 ();
 sg13g2_fill_2 FILLER_32_511 ();
 sg13g2_fill_2 FILLER_32_590 ();
 sg13g2_fill_2 FILLER_32_602 ();
 sg13g2_fill_1 FILLER_32_633 ();
 sg13g2_fill_2 FILLER_32_721 ();
 sg13g2_fill_1 FILLER_32_723 ();
 sg13g2_fill_2 FILLER_32_765 ();
 sg13g2_fill_1 FILLER_32_807 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_27 ();
 sg13g2_fill_2 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_61 ();
 sg13g2_decap_4 FILLER_33_69 ();
 sg13g2_decap_4 FILLER_33_94 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_107 ();
 sg13g2_fill_1 FILLER_33_109 ();
 sg13g2_fill_2 FILLER_33_115 ();
 sg13g2_fill_1 FILLER_33_117 ();
 sg13g2_decap_8 FILLER_33_131 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_fill_2 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_204 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_fill_1 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_267 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_fill_2 FILLER_33_340 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_fill_2 FILLER_33_369 ();
 sg13g2_fill_2 FILLER_33_380 ();
 sg13g2_fill_2 FILLER_33_410 ();
 sg13g2_fill_2 FILLER_33_421 ();
 sg13g2_fill_1 FILLER_33_423 ();
 sg13g2_fill_1 FILLER_33_436 ();
 sg13g2_fill_1 FILLER_33_447 ();
 sg13g2_fill_2 FILLER_33_528 ();
 sg13g2_fill_2 FILLER_33_544 ();
 sg13g2_fill_1 FILLER_33_598 ();
 sg13g2_fill_2 FILLER_33_616 ();
 sg13g2_fill_1 FILLER_33_664 ();
 sg13g2_fill_1 FILLER_33_740 ();
 sg13g2_fill_2 FILLER_33_787 ();
 sg13g2_decap_4 FILLER_34_43 ();
 sg13g2_fill_1 FILLER_34_62 ();
 sg13g2_fill_1 FILLER_34_89 ();
 sg13g2_decap_4 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_115 ();
 sg13g2_fill_2 FILLER_34_129 ();
 sg13g2_fill_1 FILLER_34_135 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_4 FILLER_34_168 ();
 sg13g2_fill_2 FILLER_34_180 ();
 sg13g2_fill_1 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_189 ();
 sg13g2_decap_4 FILLER_34_204 ();
 sg13g2_decap_4 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_220 ();
 sg13g2_fill_2 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_314 ();
 sg13g2_fill_1 FILLER_34_320 ();
 sg13g2_decap_4 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_431 ();
 sg13g2_fill_2 FILLER_34_451 ();
 sg13g2_fill_1 FILLER_34_453 ();
 sg13g2_decap_8 FILLER_34_462 ();
 sg13g2_decap_4 FILLER_34_469 ();
 sg13g2_fill_1 FILLER_34_473 ();
 sg13g2_fill_2 FILLER_34_491 ();
 sg13g2_fill_1 FILLER_34_503 ();
 sg13g2_fill_1 FILLER_34_561 ();
 sg13g2_fill_2 FILLER_34_571 ();
 sg13g2_fill_2 FILLER_34_582 ();
 sg13g2_fill_1 FILLER_34_584 ();
 sg13g2_fill_2 FILLER_34_594 ();
 sg13g2_fill_1 FILLER_34_601 ();
 sg13g2_fill_1 FILLER_34_768 ();
 sg13g2_fill_2 FILLER_34_774 ();
 sg13g2_fill_1 FILLER_34_776 ();
 sg13g2_fill_1 FILLER_34_810 ();
 sg13g2_fill_1 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_34 ();
 sg13g2_fill_2 FILLER_35_41 ();
 sg13g2_fill_1 FILLER_35_43 ();
 sg13g2_fill_1 FILLER_35_58 ();
 sg13g2_decap_8 FILLER_35_76 ();
 sg13g2_decap_4 FILLER_35_95 ();
 sg13g2_fill_2 FILLER_35_121 ();
 sg13g2_decap_4 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_220 ();
 sg13g2_decap_8 FILLER_35_227 ();
 sg13g2_fill_2 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_276 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_fill_2 FILLER_35_302 ();
 sg13g2_fill_1 FILLER_35_304 ();
 sg13g2_decap_4 FILLER_35_337 ();
 sg13g2_fill_1 FILLER_35_341 ();
 sg13g2_decap_4 FILLER_35_368 ();
 sg13g2_fill_1 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_fill_2 FILLER_35_409 ();
 sg13g2_fill_1 FILLER_35_439 ();
 sg13g2_decap_4 FILLER_35_445 ();
 sg13g2_fill_2 FILLER_35_449 ();
 sg13g2_decap_4 FILLER_35_468 ();
 sg13g2_fill_1 FILLER_35_472 ();
 sg13g2_fill_2 FILLER_35_502 ();
 sg13g2_fill_1 FILLER_35_544 ();
 sg13g2_fill_1 FILLER_35_564 ();
 sg13g2_fill_2 FILLER_35_752 ();
 sg13g2_fill_2 FILLER_35_786 ();
 sg13g2_fill_1 FILLER_35_788 ();
 sg13g2_fill_2 FILLER_35_813 ();
 sg13g2_fill_1 FILLER_35_857 ();
 sg13g2_fill_2 FILLER_36_26 ();
 sg13g2_decap_4 FILLER_36_71 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_fill_2 FILLER_36_118 ();
 sg13g2_fill_1 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_fill_2 FILLER_36_150 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_fill_2 FILLER_36_169 ();
 sg13g2_decap_4 FILLER_36_216 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_decap_4 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_fill_2 FILLER_36_368 ();
 sg13g2_fill_1 FILLER_36_370 ();
 sg13g2_fill_1 FILLER_36_384 ();
 sg13g2_fill_2 FILLER_36_398 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_fill_1 FILLER_36_430 ();
 sg13g2_fill_2 FILLER_36_451 ();
 sg13g2_fill_1 FILLER_36_453 ();
 sg13g2_fill_1 FILLER_36_462 ();
 sg13g2_fill_1 FILLER_36_471 ();
 sg13g2_fill_1 FILLER_36_482 ();
 sg13g2_fill_1 FILLER_36_488 ();
 sg13g2_fill_1 FILLER_36_497 ();
 sg13g2_fill_2 FILLER_36_517 ();
 sg13g2_fill_2 FILLER_36_528 ();
 sg13g2_fill_2 FILLER_36_546 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_fill_1 FILLER_36_585 ();
 sg13g2_fill_2 FILLER_36_726 ();
 sg13g2_fill_1 FILLER_36_787 ();
 sg13g2_fill_1 FILLER_36_829 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_86 ();
 sg13g2_fill_2 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_107 ();
 sg13g2_fill_2 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_139 ();
 sg13g2_decap_4 FILLER_37_145 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_fill_2 FILLER_37_176 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_decap_4 FILLER_37_213 ();
 sg13g2_fill_1 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_308 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_decap_8 FILLER_37_388 ();
 sg13g2_fill_2 FILLER_37_395 ();
 sg13g2_fill_1 FILLER_37_405 ();
 sg13g2_fill_2 FILLER_37_422 ();
 sg13g2_fill_2 FILLER_37_444 ();
 sg13g2_fill_1 FILLER_37_446 ();
 sg13g2_fill_2 FILLER_37_460 ();
 sg13g2_fill_1 FILLER_37_462 ();
 sg13g2_fill_1 FILLER_37_471 ();
 sg13g2_decap_4 FILLER_37_488 ();
 sg13g2_fill_2 FILLER_37_492 ();
 sg13g2_fill_2 FILLER_37_553 ();
 sg13g2_fill_1 FILLER_37_555 ();
 sg13g2_fill_2 FILLER_37_564 ();
 sg13g2_fill_1 FILLER_37_566 ();
 sg13g2_fill_2 FILLER_37_576 ();
 sg13g2_fill_1 FILLER_37_790 ();
 sg13g2_fill_2 FILLER_37_826 ();
 sg13g2_fill_1 FILLER_37_828 ();
 sg13g2_fill_2 FILLER_37_834 ();
 sg13g2_decap_4 FILLER_38_26 ();
 sg13g2_fill_1 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_115 ();
 sg13g2_fill_2 FILLER_38_149 ();
 sg13g2_fill_1 FILLER_38_160 ();
 sg13g2_fill_2 FILLER_38_175 ();
 sg13g2_fill_2 FILLER_38_204 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_288 ();
 sg13g2_fill_2 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_fill_2 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_329 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_fill_2 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_371 ();
 sg13g2_fill_2 FILLER_38_396 ();
 sg13g2_decap_8 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_450 ();
 sg13g2_decap_8 FILLER_38_467 ();
 sg13g2_decap_8 FILLER_38_486 ();
 sg13g2_decap_4 FILLER_38_493 ();
 sg13g2_fill_1 FILLER_38_497 ();
 sg13g2_decap_4 FILLER_38_506 ();
 sg13g2_fill_2 FILLER_38_534 ();
 sg13g2_fill_1 FILLER_38_536 ();
 sg13g2_fill_1 FILLER_38_541 ();
 sg13g2_fill_2 FILLER_38_552 ();
 sg13g2_decap_4 FILLER_38_567 ();
 sg13g2_fill_2 FILLER_38_673 ();
 sg13g2_fill_2 FILLER_38_841 ();
 sg13g2_fill_1 FILLER_38_843 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_21 ();
 sg13g2_decap_4 FILLER_39_54 ();
 sg13g2_fill_1 FILLER_39_58 ();
 sg13g2_fill_2 FILLER_39_74 ();
 sg13g2_fill_1 FILLER_39_85 ();
 sg13g2_decap_4 FILLER_39_178 ();
 sg13g2_fill_2 FILLER_39_214 ();
 sg13g2_decap_4 FILLER_39_246 ();
 sg13g2_fill_2 FILLER_39_250 ();
 sg13g2_fill_1 FILLER_39_270 ();
 sg13g2_fill_1 FILLER_39_290 ();
 sg13g2_decap_8 FILLER_39_317 ();
 sg13g2_fill_1 FILLER_39_324 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_fill_1 FILLER_39_350 ();
 sg13g2_decap_4 FILLER_39_364 ();
 sg13g2_fill_2 FILLER_39_373 ();
 sg13g2_fill_1 FILLER_39_375 ();
 sg13g2_decap_4 FILLER_39_409 ();
 sg13g2_decap_4 FILLER_39_443 ();
 sg13g2_fill_2 FILLER_39_492 ();
 sg13g2_decap_8 FILLER_39_518 ();
 sg13g2_fill_1 FILLER_39_525 ();
 sg13g2_fill_2 FILLER_39_539 ();
 sg13g2_decap_8 FILLER_39_557 ();
 sg13g2_fill_1 FILLER_39_564 ();
 sg13g2_fill_1 FILLER_39_586 ();
 sg13g2_fill_1 FILLER_39_597 ();
 sg13g2_fill_2 FILLER_39_650 ();
 sg13g2_fill_1 FILLER_39_652 ();
 sg13g2_fill_2 FILLER_39_795 ();
 sg13g2_fill_2 FILLER_39_810 ();
 sg13g2_fill_1 FILLER_39_822 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_fill_2 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_37 ();
 sg13g2_fill_1 FILLER_40_80 ();
 sg13g2_decap_4 FILLER_40_149 ();
 sg13g2_fill_2 FILLER_40_166 ();
 sg13g2_fill_1 FILLER_40_168 ();
 sg13g2_fill_2 FILLER_40_185 ();
 sg13g2_fill_2 FILLER_40_203 ();
 sg13g2_fill_1 FILLER_40_205 ();
 sg13g2_fill_2 FILLER_40_232 ();
 sg13g2_fill_1 FILLER_40_234 ();
 sg13g2_fill_2 FILLER_40_243 ();
 sg13g2_fill_1 FILLER_40_245 ();
 sg13g2_fill_2 FILLER_40_251 ();
 sg13g2_decap_4 FILLER_40_257 ();
 sg13g2_fill_1 FILLER_40_261 ();
 sg13g2_fill_2 FILLER_40_285 ();
 sg13g2_fill_1 FILLER_40_287 ();
 sg13g2_fill_2 FILLER_40_310 ();
 sg13g2_decap_4 FILLER_40_365 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_fill_2 FILLER_40_399 ();
 sg13g2_fill_1 FILLER_40_401 ();
 sg13g2_decap_4 FILLER_40_407 ();
 sg13g2_decap_4 FILLER_40_434 ();
 sg13g2_fill_1 FILLER_40_438 ();
 sg13g2_fill_1 FILLER_40_452 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_fill_1 FILLER_40_476 ();
 sg13g2_fill_2 FILLER_40_482 ();
 sg13g2_fill_1 FILLER_40_484 ();
 sg13g2_decap_8 FILLER_40_523 ();
 sg13g2_fill_1 FILLER_40_530 ();
 sg13g2_decap_8 FILLER_40_554 ();
 sg13g2_decap_4 FILLER_40_578 ();
 sg13g2_fill_2 FILLER_40_582 ();
 sg13g2_fill_2 FILLER_40_713 ();
 sg13g2_fill_1 FILLER_40_754 ();
 sg13g2_fill_1 FILLER_40_795 ();
 sg13g2_fill_2 FILLER_40_836 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_4 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_15 ();
 sg13g2_fill_2 FILLER_41_19 ();
 sg13g2_fill_2 FILLER_41_35 ();
 sg13g2_fill_1 FILLER_41_37 ();
 sg13g2_decap_8 FILLER_41_43 ();
 sg13g2_fill_2 FILLER_41_50 ();
 sg13g2_fill_1 FILLER_41_73 ();
 sg13g2_fill_1 FILLER_41_82 ();
 sg13g2_fill_2 FILLER_41_90 ();
 sg13g2_fill_1 FILLER_41_92 ();
 sg13g2_decap_4 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_105 ();
 sg13g2_decap_4 FILLER_41_111 ();
 sg13g2_fill_1 FILLER_41_115 ();
 sg13g2_fill_2 FILLER_41_133 ();
 sg13g2_fill_1 FILLER_41_135 ();
 sg13g2_decap_4 FILLER_41_155 ();
 sg13g2_decap_8 FILLER_41_188 ();
 sg13g2_decap_8 FILLER_41_195 ();
 sg13g2_decap_8 FILLER_41_202 ();
 sg13g2_decap_4 FILLER_41_209 ();
 sg13g2_fill_1 FILLER_41_213 ();
 sg13g2_fill_2 FILLER_41_242 ();
 sg13g2_fill_1 FILLER_41_244 ();
 sg13g2_fill_2 FILLER_41_253 ();
 sg13g2_fill_1 FILLER_41_255 ();
 sg13g2_fill_1 FILLER_41_259 ();
 sg13g2_fill_1 FILLER_41_264 ();
 sg13g2_fill_2 FILLER_41_273 ();
 sg13g2_fill_1 FILLER_41_306 ();
 sg13g2_fill_2 FILLER_41_315 ();
 sg13g2_fill_1 FILLER_41_317 ();
 sg13g2_fill_1 FILLER_41_331 ();
 sg13g2_fill_2 FILLER_41_337 ();
 sg13g2_fill_1 FILLER_41_339 ();
 sg13g2_fill_1 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_367 ();
 sg13g2_fill_2 FILLER_41_382 ();
 sg13g2_fill_1 FILLER_41_384 ();
 sg13g2_fill_2 FILLER_41_411 ();
 sg13g2_fill_1 FILLER_41_413 ();
 sg13g2_decap_4 FILLER_41_435 ();
 sg13g2_fill_2 FILLER_41_439 ();
 sg13g2_fill_2 FILLER_41_453 ();
 sg13g2_decap_8 FILLER_41_463 ();
 sg13g2_fill_2 FILLER_41_470 ();
 sg13g2_fill_1 FILLER_41_472 ();
 sg13g2_decap_8 FILLER_41_530 ();
 sg13g2_decap_4 FILLER_41_537 ();
 sg13g2_fill_1 FILLER_41_541 ();
 sg13g2_fill_2 FILLER_41_558 ();
 sg13g2_fill_2 FILLER_41_586 ();
 sg13g2_fill_2 FILLER_41_605 ();
 sg13g2_fill_1 FILLER_41_607 ();
 sg13g2_fill_1 FILLER_41_629 ();
 sg13g2_fill_1 FILLER_41_726 ();
 sg13g2_fill_2 FILLER_41_743 ();
 sg13g2_fill_1 FILLER_41_745 ();
 sg13g2_fill_1 FILLER_41_759 ();
 sg13g2_fill_2 FILLER_41_769 ();
 sg13g2_fill_2 FILLER_41_788 ();
 sg13g2_fill_2 FILLER_41_795 ();
 sg13g2_fill_1 FILLER_41_813 ();
 sg13g2_fill_2 FILLER_41_833 ();
 sg13g2_fill_2 FILLER_41_842 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_7 ();
 sg13g2_decap_4 FILLER_42_15 ();
 sg13g2_fill_2 FILLER_42_19 ();
 sg13g2_decap_8 FILLER_42_51 ();
 sg13g2_fill_1 FILLER_42_58 ();
 sg13g2_fill_1 FILLER_42_67 ();
 sg13g2_fill_1 FILLER_42_77 ();
 sg13g2_fill_1 FILLER_42_83 ();
 sg13g2_fill_1 FILLER_42_89 ();
 sg13g2_fill_2 FILLER_42_94 ();
 sg13g2_fill_1 FILLER_42_96 ();
 sg13g2_fill_2 FILLER_42_137 ();
 sg13g2_decap_8 FILLER_42_155 ();
 sg13g2_fill_1 FILLER_42_162 ();
 sg13g2_fill_2 FILLER_42_187 ();
 sg13g2_fill_2 FILLER_42_203 ();
 sg13g2_fill_1 FILLER_42_205 ();
 sg13g2_fill_2 FILLER_42_223 ();
 sg13g2_fill_2 FILLER_42_247 ();
 sg13g2_fill_1 FILLER_42_330 ();
 sg13g2_fill_1 FILLER_42_353 ();
 sg13g2_decap_4 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_415 ();
 sg13g2_decap_8 FILLER_42_486 ();
 sg13g2_decap_4 FILLER_42_493 ();
 sg13g2_fill_1 FILLER_42_497 ();
 sg13g2_decap_4 FILLER_42_506 ();
 sg13g2_fill_2 FILLER_42_510 ();
 sg13g2_decap_4 FILLER_42_536 ();
 sg13g2_fill_2 FILLER_42_540 ();
 sg13g2_decap_8 FILLER_42_554 ();
 sg13g2_decap_8 FILLER_42_561 ();
 sg13g2_decap_4 FILLER_42_568 ();
 sg13g2_fill_1 FILLER_42_576 ();
 sg13g2_decap_8 FILLER_42_582 ();
 sg13g2_fill_2 FILLER_42_589 ();
 sg13g2_fill_2 FILLER_42_607 ();
 sg13g2_fill_1 FILLER_42_626 ();
 sg13g2_fill_1 FILLER_42_681 ();
 sg13g2_fill_1 FILLER_42_822 ();
 sg13g2_fill_2 FILLER_42_845 ();
 sg13g2_fill_2 FILLER_42_860 ();
 sg13g2_decap_4 FILLER_43_26 ();
 sg13g2_fill_2 FILLER_43_74 ();
 sg13g2_decap_4 FILLER_43_94 ();
 sg13g2_fill_1 FILLER_43_98 ();
 sg13g2_fill_2 FILLER_43_111 ();
 sg13g2_fill_1 FILLER_43_113 ();
 sg13g2_decap_8 FILLER_43_124 ();
 sg13g2_fill_2 FILLER_43_151 ();
 sg13g2_fill_2 FILLER_43_177 ();
 sg13g2_fill_1 FILLER_43_179 ();
 sg13g2_decap_8 FILLER_43_185 ();
 sg13g2_fill_2 FILLER_43_192 ();
 sg13g2_fill_2 FILLER_43_202 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_4 FILLER_43_224 ();
 sg13g2_fill_2 FILLER_43_228 ();
 sg13g2_fill_2 FILLER_43_235 ();
 sg13g2_fill_1 FILLER_43_253 ();
 sg13g2_fill_2 FILLER_43_259 ();
 sg13g2_fill_1 FILLER_43_261 ();
 sg13g2_fill_2 FILLER_43_288 ();
 sg13g2_decap_8 FILLER_43_298 ();
 sg13g2_fill_1 FILLER_43_305 ();
 sg13g2_fill_1 FILLER_43_311 ();
 sg13g2_fill_2 FILLER_43_321 ();
 sg13g2_fill_2 FILLER_43_358 ();
 sg13g2_fill_1 FILLER_43_360 ();
 sg13g2_decap_8 FILLER_43_373 ();
 sg13g2_decap_4 FILLER_43_380 ();
 sg13g2_fill_1 FILLER_43_384 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_4 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_419 ();
 sg13g2_decap_4 FILLER_43_434 ();
 sg13g2_fill_2 FILLER_43_438 ();
 sg13g2_decap_8 FILLER_43_453 ();
 sg13g2_decap_8 FILLER_43_460 ();
 sg13g2_fill_2 FILLER_43_467 ();
 sg13g2_decap_8 FILLER_43_482 ();
 sg13g2_fill_1 FILLER_43_489 ();
 sg13g2_decap_4 FILLER_43_506 ();
 sg13g2_fill_2 FILLER_43_510 ();
 sg13g2_fill_1 FILLER_43_520 ();
 sg13g2_fill_1 FILLER_43_675 ();
 sg13g2_fill_1 FILLER_43_766 ();
 sg13g2_decap_4 FILLER_43_836 ();
 sg13g2_fill_2 FILLER_43_840 ();
 sg13g2_decap_4 FILLER_43_858 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_4 FILLER_44_7 ();
 sg13g2_decap_4 FILLER_44_15 ();
 sg13g2_decap_4 FILLER_44_40 ();
 sg13g2_fill_2 FILLER_44_70 ();
 sg13g2_fill_2 FILLER_44_76 ();
 sg13g2_decap_4 FILLER_44_85 ();
 sg13g2_fill_1 FILLER_44_89 ();
 sg13g2_fill_2 FILLER_44_106 ();
 sg13g2_fill_2 FILLER_44_139 ();
 sg13g2_decap_4 FILLER_44_170 ();
 sg13g2_decap_4 FILLER_44_204 ();
 sg13g2_fill_1 FILLER_44_220 ();
 sg13g2_fill_2 FILLER_44_237 ();
 sg13g2_fill_1 FILLER_44_239 ();
 sg13g2_fill_1 FILLER_44_253 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_8 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_306 ();
 sg13g2_fill_2 FILLER_44_313 ();
 sg13g2_decap_8 FILLER_44_354 ();
 sg13g2_decap_4 FILLER_44_361 ();
 sg13g2_fill_1 FILLER_44_400 ();
 sg13g2_fill_1 FILLER_44_436 ();
 sg13g2_fill_2 FILLER_44_444 ();
 sg13g2_fill_1 FILLER_44_446 ();
 sg13g2_decap_4 FILLER_44_462 ();
 sg13g2_fill_1 FILLER_44_466 ();
 sg13g2_decap_8 FILLER_44_487 ();
 sg13g2_decap_4 FILLER_44_510 ();
 sg13g2_fill_1 FILLER_44_514 ();
 sg13g2_fill_2 FILLER_44_523 ();
 sg13g2_fill_1 FILLER_44_525 ();
 sg13g2_fill_2 FILLER_44_546 ();
 sg13g2_decap_4 FILLER_44_560 ();
 sg13g2_fill_2 FILLER_44_564 ();
 sg13g2_decap_4 FILLER_44_574 ();
 sg13g2_fill_1 FILLER_44_578 ();
 sg13g2_decap_8 FILLER_44_587 ();
 sg13g2_decap_4 FILLER_44_594 ();
 sg13g2_decap_4 FILLER_44_606 ();
 sg13g2_fill_1 FILLER_44_610 ();
 sg13g2_fill_1 FILLER_44_629 ();
 sg13g2_fill_2 FILLER_44_746 ();
 sg13g2_fill_1 FILLER_44_748 ();
 sg13g2_fill_1 FILLER_44_765 ();
 sg13g2_fill_1 FILLER_44_776 ();
 sg13g2_fill_1 FILLER_44_790 ();
 sg13g2_decap_4 FILLER_44_826 ();
 sg13g2_fill_1 FILLER_44_834 ();
 sg13g2_fill_2 FILLER_44_860 ();
 sg13g2_fill_1 FILLER_45_34 ();
 sg13g2_decap_4 FILLER_45_43 ();
 sg13g2_fill_1 FILLER_45_54 ();
 sg13g2_fill_2 FILLER_45_92 ();
 sg13g2_fill_1 FILLER_45_94 ();
 sg13g2_fill_2 FILLER_45_118 ();
 sg13g2_fill_1 FILLER_45_143 ();
 sg13g2_decap_8 FILLER_45_148 ();
 sg13g2_fill_2 FILLER_45_176 ();
 sg13g2_fill_1 FILLER_45_178 ();
 sg13g2_decap_4 FILLER_45_219 ();
 sg13g2_fill_2 FILLER_45_223 ();
 sg13g2_fill_2 FILLER_45_234 ();
 sg13g2_fill_1 FILLER_45_236 ();
 sg13g2_fill_2 FILLER_45_249 ();
 sg13g2_fill_1 FILLER_45_251 ();
 sg13g2_fill_1 FILLER_45_265 ();
 sg13g2_decap_8 FILLER_45_270 ();
 sg13g2_decap_8 FILLER_45_277 ();
 sg13g2_decap_8 FILLER_45_290 ();
 sg13g2_decap_4 FILLER_45_297 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_fill_2 FILLER_45_326 ();
 sg13g2_decap_4 FILLER_45_337 ();
 sg13g2_fill_2 FILLER_45_388 ();
 sg13g2_fill_1 FILLER_45_390 ();
 sg13g2_fill_2 FILLER_45_403 ();
 sg13g2_fill_2 FILLER_45_437 ();
 sg13g2_fill_2 FILLER_45_452 ();
 sg13g2_fill_1 FILLER_45_459 ();
 sg13g2_fill_2 FILLER_45_481 ();
 sg13g2_fill_1 FILLER_45_483 ();
 sg13g2_fill_2 FILLER_45_513 ();
 sg13g2_fill_2 FILLER_45_523 ();
 sg13g2_decap_4 FILLER_45_537 ();
 sg13g2_fill_2 FILLER_45_541 ();
 sg13g2_decap_8 FILLER_45_555 ();
 sg13g2_fill_1 FILLER_45_562 ();
 sg13g2_decap_8 FILLER_45_587 ();
 sg13g2_decap_8 FILLER_45_594 ();
 sg13g2_fill_1 FILLER_45_619 ();
 sg13g2_fill_1 FILLER_45_664 ();
 sg13g2_fill_1 FILLER_45_677 ();
 sg13g2_fill_2 FILLER_45_684 ();
 sg13g2_fill_1 FILLER_45_686 ();
 sg13g2_fill_1 FILLER_45_740 ();
 sg13g2_decap_4 FILLER_45_821 ();
 sg13g2_fill_2 FILLER_45_841 ();
 sg13g2_fill_1 FILLER_45_857 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_41 ();
 sg13g2_decap_4 FILLER_46_65 ();
 sg13g2_fill_1 FILLER_46_69 ();
 sg13g2_decap_4 FILLER_46_98 ();
 sg13g2_fill_1 FILLER_46_102 ();
 sg13g2_fill_2 FILLER_46_129 ();
 sg13g2_fill_1 FILLER_46_131 ();
 sg13g2_fill_2 FILLER_46_167 ();
 sg13g2_fill_1 FILLER_46_169 ();
 sg13g2_fill_2 FILLER_46_183 ();
 sg13g2_fill_1 FILLER_46_193 ();
 sg13g2_fill_1 FILLER_46_210 ();
 sg13g2_fill_2 FILLER_46_227 ();
 sg13g2_decap_4 FILLER_46_250 ();
 sg13g2_fill_2 FILLER_46_254 ();
 sg13g2_fill_1 FILLER_46_277 ();
 sg13g2_decap_8 FILLER_46_348 ();
 sg13g2_fill_1 FILLER_46_414 ();
 sg13g2_decap_4 FILLER_46_444 ();
 sg13g2_fill_1 FILLER_46_448 ();
 sg13g2_fill_2 FILLER_46_457 ();
 sg13g2_fill_1 FILLER_46_459 ();
 sg13g2_fill_2 FILLER_46_480 ();
 sg13g2_fill_1 FILLER_46_482 ();
 sg13g2_fill_1 FILLER_46_495 ();
 sg13g2_fill_2 FILLER_46_508 ();
 sg13g2_fill_1 FILLER_46_510 ();
 sg13g2_fill_2 FILLER_46_529 ();
 sg13g2_fill_2 FILLER_46_593 ();
 sg13g2_fill_1 FILLER_46_595 ();
 sg13g2_fill_2 FILLER_46_623 ();
 sg13g2_fill_1 FILLER_46_685 ();
 sg13g2_fill_2 FILLER_46_736 ();
 sg13g2_fill_1 FILLER_46_747 ();
 sg13g2_fill_2 FILLER_46_761 ();
 sg13g2_fill_1 FILLER_46_771 ();
 sg13g2_fill_2 FILLER_46_817 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_decap_4 FILLER_47_60 ();
 sg13g2_decap_4 FILLER_47_79 ();
 sg13g2_decap_8 FILLER_47_88 ();
 sg13g2_fill_1 FILLER_47_95 ();
 sg13g2_fill_1 FILLER_47_125 ();
 sg13g2_decap_8 FILLER_47_135 ();
 sg13g2_fill_2 FILLER_47_150 ();
 sg13g2_fill_1 FILLER_47_152 ();
 sg13g2_fill_2 FILLER_47_178 ();
 sg13g2_fill_1 FILLER_47_180 ();
 sg13g2_decap_8 FILLER_47_197 ();
 sg13g2_fill_2 FILLER_47_204 ();
 sg13g2_fill_2 FILLER_47_227 ();
 sg13g2_fill_1 FILLER_47_229 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_4 FILLER_47_245 ();
 sg13g2_fill_2 FILLER_47_266 ();
 sg13g2_fill_1 FILLER_47_268 ();
 sg13g2_fill_2 FILLER_47_302 ();
 sg13g2_fill_1 FILLER_47_304 ();
 sg13g2_fill_2 FILLER_47_313 ();
 sg13g2_fill_1 FILLER_47_315 ();
 sg13g2_fill_1 FILLER_47_324 ();
 sg13g2_fill_2 FILLER_47_338 ();
 sg13g2_fill_2 FILLER_47_366 ();
 sg13g2_fill_1 FILLER_47_381 ();
 sg13g2_fill_1 FILLER_47_414 ();
 sg13g2_fill_1 FILLER_47_459 ();
 sg13g2_fill_2 FILLER_47_494 ();
 sg13g2_fill_1 FILLER_47_496 ();
 sg13g2_fill_2 FILLER_47_541 ();
 sg13g2_fill_1 FILLER_47_543 ();
 sg13g2_decap_4 FILLER_47_552 ();
 sg13g2_fill_2 FILLER_47_564 ();
 sg13g2_fill_1 FILLER_47_566 ();
 sg13g2_decap_4 FILLER_47_571 ();
 sg13g2_decap_4 FILLER_47_586 ();
 sg13g2_fill_1 FILLER_47_590 ();
 sg13g2_fill_1 FILLER_47_596 ();
 sg13g2_decap_4 FILLER_47_601 ();
 sg13g2_fill_1 FILLER_47_630 ();
 sg13g2_fill_2 FILLER_47_656 ();
 sg13g2_fill_1 FILLER_47_677 ();
 sg13g2_fill_2 FILLER_47_700 ();
 sg13g2_fill_2 FILLER_47_738 ();
 sg13g2_fill_1 FILLER_47_761 ();
 sg13g2_fill_2 FILLER_47_767 ();
 sg13g2_fill_1 FILLER_47_791 ();
 sg13g2_fill_2 FILLER_47_815 ();
 sg13g2_fill_2 FILLER_47_843 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_22 ();
 sg13g2_fill_2 FILLER_48_38 ();
 sg13g2_fill_2 FILLER_48_45 ();
 sg13g2_decap_8 FILLER_48_80 ();
 sg13g2_decap_8 FILLER_48_108 ();
 sg13g2_fill_1 FILLER_48_115 ();
 sg13g2_decap_4 FILLER_48_142 ();
 sg13g2_fill_2 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_153 ();
 sg13g2_fill_2 FILLER_48_160 ();
 sg13g2_fill_2 FILLER_48_183 ();
 sg13g2_fill_1 FILLER_48_185 ();
 sg13g2_fill_2 FILLER_48_199 ();
 sg13g2_fill_1 FILLER_48_201 ();
 sg13g2_fill_2 FILLER_48_210 ();
 sg13g2_fill_1 FILLER_48_212 ();
 sg13g2_decap_8 FILLER_48_254 ();
 sg13g2_fill_1 FILLER_48_273 ();
 sg13g2_fill_2 FILLER_48_279 ();
 sg13g2_decap_4 FILLER_48_311 ();
 sg13g2_decap_8 FILLER_48_330 ();
 sg13g2_decap_4 FILLER_48_337 ();
 sg13g2_fill_1 FILLER_48_360 ();
 sg13g2_decap_4 FILLER_48_385 ();
 sg13g2_fill_2 FILLER_48_394 ();
 sg13g2_fill_1 FILLER_48_396 ();
 sg13g2_fill_1 FILLER_48_435 ();
 sg13g2_decap_4 FILLER_48_459 ();
 sg13g2_fill_2 FILLER_48_463 ();
 sg13g2_decap_4 FILLER_48_475 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_fill_1 FILLER_48_490 ();
 sg13g2_fill_1 FILLER_48_535 ();
 sg13g2_decap_4 FILLER_48_548 ();
 sg13g2_fill_1 FILLER_48_552 ();
 sg13g2_fill_1 FILLER_48_569 ();
 sg13g2_fill_2 FILLER_48_646 ();
 sg13g2_fill_2 FILLER_48_653 ();
 sg13g2_fill_1 FILLER_48_708 ();
 sg13g2_fill_1 FILLER_48_733 ();
 sg13g2_fill_2 FILLER_48_759 ();
 sg13g2_fill_1 FILLER_48_761 ();
 sg13g2_fill_1 FILLER_48_772 ();
 sg13g2_fill_1 FILLER_48_790 ();
 sg13g2_fill_1 FILLER_48_812 ();
 sg13g2_decap_4 FILLER_48_817 ();
 sg13g2_fill_1 FILLER_48_821 ();
 sg13g2_fill_1 FILLER_48_843 ();
 sg13g2_fill_2 FILLER_49_89 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_106 ();
 sg13g2_fill_1 FILLER_49_137 ();
 sg13g2_fill_2 FILLER_49_164 ();
 sg13g2_fill_2 FILLER_49_182 ();
 sg13g2_fill_1 FILLER_49_184 ();
 sg13g2_fill_2 FILLER_49_215 ();
 sg13g2_fill_2 FILLER_49_232 ();
 sg13g2_fill_1 FILLER_49_234 ();
 sg13g2_fill_2 FILLER_49_244 ();
 sg13g2_fill_2 FILLER_49_258 ();
 sg13g2_fill_1 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_278 ();
 sg13g2_fill_2 FILLER_49_285 ();
 sg13g2_fill_2 FILLER_49_301 ();
 sg13g2_fill_2 FILLER_49_311 ();
 sg13g2_decap_4 FILLER_49_342 ();
 sg13g2_fill_1 FILLER_49_346 ();
 sg13g2_fill_2 FILLER_49_382 ();
 sg13g2_decap_4 FILLER_49_393 ();
 sg13g2_fill_1 FILLER_49_401 ();
 sg13g2_fill_2 FILLER_49_435 ();
 sg13g2_fill_1 FILLER_49_445 ();
 sg13g2_fill_2 FILLER_49_459 ();
 sg13g2_fill_1 FILLER_49_461 ();
 sg13g2_decap_4 FILLER_49_512 ();
 sg13g2_fill_2 FILLER_49_529 ();
 sg13g2_fill_1 FILLER_49_531 ();
 sg13g2_fill_2 FILLER_49_556 ();
 sg13g2_fill_1 FILLER_49_558 ();
 sg13g2_fill_2 FILLER_49_573 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_4 FILLER_49_595 ();
 sg13g2_decap_4 FILLER_49_611 ();
 sg13g2_fill_2 FILLER_49_615 ();
 sg13g2_decap_8 FILLER_49_622 ();
 sg13g2_fill_1 FILLER_49_629 ();
 sg13g2_decap_4 FILLER_49_635 ();
 sg13g2_fill_2 FILLER_49_639 ();
 sg13g2_fill_1 FILLER_49_650 ();
 sg13g2_fill_2 FILLER_49_690 ();
 sg13g2_fill_2 FILLER_49_702 ();
 sg13g2_fill_2 FILLER_49_726 ();
 sg13g2_fill_2 FILLER_49_748 ();
 sg13g2_fill_1 FILLER_49_750 ();
 sg13g2_decap_4 FILLER_49_786 ();
 sg13g2_fill_1 FILLER_49_790 ();
 sg13g2_fill_2 FILLER_49_800 ();
 sg13g2_fill_1 FILLER_49_802 ();
 sg13g2_fill_1 FILLER_49_812 ();
 sg13g2_fill_1 FILLER_49_835 ();
 sg13g2_fill_2 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_31 ();
 sg13g2_fill_1 FILLER_50_62 ();
 sg13g2_decap_8 FILLER_50_109 ();
 sg13g2_fill_1 FILLER_50_116 ();
 sg13g2_decap_4 FILLER_50_171 ();
 sg13g2_fill_2 FILLER_50_180 ();
 sg13g2_fill_1 FILLER_50_182 ();
 sg13g2_fill_1 FILLER_50_187 ();
 sg13g2_decap_4 FILLER_50_193 ();
 sg13g2_fill_1 FILLER_50_205 ();
 sg13g2_decap_8 FILLER_50_211 ();
 sg13g2_fill_2 FILLER_50_218 ();
 sg13g2_fill_1 FILLER_50_254 ();
 sg13g2_decap_8 FILLER_50_307 ();
 sg13g2_fill_2 FILLER_50_314 ();
 sg13g2_fill_1 FILLER_50_316 ();
 sg13g2_fill_1 FILLER_50_345 ();
 sg13g2_fill_1 FILLER_50_374 ();
 sg13g2_fill_2 FILLER_50_412 ();
 sg13g2_fill_1 FILLER_50_423 ();
 sg13g2_fill_1 FILLER_50_432 ();
 sg13g2_fill_1 FILLER_50_437 ();
 sg13g2_fill_2 FILLER_50_450 ();
 sg13g2_fill_1 FILLER_50_463 ();
 sg13g2_fill_2 FILLER_50_481 ();
 sg13g2_fill_1 FILLER_50_499 ();
 sg13g2_fill_2 FILLER_50_516 ();
 sg13g2_fill_1 FILLER_50_518 ();
 sg13g2_decap_8 FILLER_50_543 ();
 sg13g2_fill_2 FILLER_50_550 ();
 sg13g2_decap_4 FILLER_50_596 ();
 sg13g2_fill_1 FILLER_50_600 ();
 sg13g2_decap_8 FILLER_50_620 ();
 sg13g2_decap_4 FILLER_50_627 ();
 sg13g2_decap_4 FILLER_50_646 ();
 sg13g2_fill_1 FILLER_50_650 ();
 sg13g2_fill_2 FILLER_50_671 ();
 sg13g2_fill_1 FILLER_50_700 ();
 sg13g2_decap_4 FILLER_50_728 ();
 sg13g2_fill_2 FILLER_50_732 ();
 sg13g2_decap_4 FILLER_50_779 ();
 sg13g2_decap_4 FILLER_50_791 ();
 sg13g2_fill_2 FILLER_50_795 ();
 sg13g2_fill_2 FILLER_50_810 ();
 sg13g2_fill_1 FILLER_50_812 ();
 sg13g2_fill_1 FILLER_50_821 ();
 sg13g2_fill_2 FILLER_50_840 ();
 sg13g2_fill_1 FILLER_50_842 ();
 sg13g2_fill_2 FILLER_50_859 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_53 ();
 sg13g2_fill_1 FILLER_51_90 ();
 sg13g2_fill_1 FILLER_51_130 ();
 sg13g2_fill_2 FILLER_51_141 ();
 sg13g2_fill_1 FILLER_51_148 ();
 sg13g2_fill_1 FILLER_51_191 ();
 sg13g2_fill_1 FILLER_51_216 ();
 sg13g2_decap_8 FILLER_51_221 ();
 sg13g2_fill_2 FILLER_51_228 ();
 sg13g2_fill_1 FILLER_51_235 ();
 sg13g2_fill_2 FILLER_51_259 ();
 sg13g2_fill_1 FILLER_51_261 ();
 sg13g2_decap_8 FILLER_51_280 ();
 sg13g2_decap_4 FILLER_51_287 ();
 sg13g2_fill_2 FILLER_51_291 ();
 sg13g2_decap_8 FILLER_51_314 ();
 sg13g2_fill_2 FILLER_51_321 ();
 sg13g2_fill_1 FILLER_51_323 ();
 sg13g2_fill_1 FILLER_51_342 ();
 sg13g2_fill_1 FILLER_51_368 ();
 sg13g2_fill_2 FILLER_51_387 ();
 sg13g2_fill_1 FILLER_51_398 ();
 sg13g2_decap_4 FILLER_51_407 ();
 sg13g2_fill_1 FILLER_51_411 ();
 sg13g2_fill_2 FILLER_51_416 ();
 sg13g2_fill_2 FILLER_51_439 ();
 sg13g2_fill_2 FILLER_51_488 ();
 sg13g2_fill_1 FILLER_51_506 ();
 sg13g2_fill_1 FILLER_51_520 ();
 sg13g2_fill_1 FILLER_51_548 ();
 sg13g2_decap_4 FILLER_51_562 ();
 sg13g2_fill_1 FILLER_51_566 ();
 sg13g2_decap_8 FILLER_51_575 ();
 sg13g2_fill_2 FILLER_51_624 ();
 sg13g2_fill_2 FILLER_51_668 ();
 sg13g2_fill_1 FILLER_51_670 ();
 sg13g2_fill_1 FILLER_51_676 ();
 sg13g2_fill_1 FILLER_51_717 ();
 sg13g2_fill_2 FILLER_51_723 ();
 sg13g2_fill_1 FILLER_51_738 ();
 sg13g2_fill_2 FILLER_51_749 ();
 sg13g2_fill_1 FILLER_51_782 ();
 sg13g2_fill_2 FILLER_51_788 ();
 sg13g2_decap_8 FILLER_51_806 ();
 sg13g2_fill_2 FILLER_51_833 ();
 sg13g2_decap_4 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_4 ();
 sg13g2_decap_8 FILLER_52_32 ();
 sg13g2_decap_4 FILLER_52_39 ();
 sg13g2_fill_1 FILLER_52_43 ();
 sg13g2_fill_2 FILLER_52_61 ();
 sg13g2_fill_1 FILLER_52_63 ();
 sg13g2_fill_1 FILLER_52_91 ();
 sg13g2_fill_2 FILLER_52_106 ();
 sg13g2_decap_8 FILLER_52_113 ();
 sg13g2_fill_1 FILLER_52_120 ();
 sg13g2_fill_2 FILLER_52_155 ();
 sg13g2_fill_1 FILLER_52_162 ();
 sg13g2_decap_8 FILLER_52_198 ();
 sg13g2_fill_2 FILLER_52_205 ();
 sg13g2_decap_4 FILLER_52_235 ();
 sg13g2_fill_2 FILLER_52_244 ();
 sg13g2_fill_1 FILLER_52_246 ();
 sg13g2_fill_1 FILLER_52_256 ();
 sg13g2_fill_2 FILLER_52_273 ();
 sg13g2_fill_2 FILLER_52_285 ();
 sg13g2_fill_1 FILLER_52_287 ();
 sg13g2_fill_2 FILLER_52_300 ();
 sg13g2_decap_8 FILLER_52_306 ();
 sg13g2_fill_2 FILLER_52_313 ();
 sg13g2_fill_1 FILLER_52_323 ();
 sg13g2_fill_2 FILLER_52_334 ();
 sg13g2_fill_1 FILLER_52_336 ();
 sg13g2_fill_1 FILLER_52_374 ();
 sg13g2_fill_2 FILLER_52_399 ();
 sg13g2_fill_1 FILLER_52_401 ();
 sg13g2_decap_8 FILLER_52_438 ();
 sg13g2_fill_2 FILLER_52_488 ();
 sg13g2_fill_1 FILLER_52_490 ();
 sg13g2_fill_1 FILLER_52_499 ();
 sg13g2_fill_1 FILLER_52_521 ();
 sg13g2_fill_2 FILLER_52_544 ();
 sg13g2_fill_2 FILLER_52_558 ();
 sg13g2_decap_8 FILLER_52_578 ();
 sg13g2_decap_4 FILLER_52_593 ();
 sg13g2_fill_1 FILLER_52_597 ();
 sg13g2_decap_4 FILLER_52_618 ();
 sg13g2_fill_1 FILLER_52_622 ();
 sg13g2_fill_2 FILLER_52_646 ();
 sg13g2_fill_1 FILLER_52_648 ();
 sg13g2_fill_2 FILLER_52_653 ();
 sg13g2_decap_8 FILLER_52_689 ();
 sg13g2_fill_2 FILLER_52_696 ();
 sg13g2_fill_1 FILLER_52_698 ();
 sg13g2_fill_2 FILLER_52_709 ();
 sg13g2_fill_1 FILLER_52_711 ();
 sg13g2_decap_4 FILLER_52_775 ();
 sg13g2_decap_8 FILLER_52_808 ();
 sg13g2_fill_1 FILLER_52_815 ();
 sg13g2_decap_8 FILLER_52_832 ();
 sg13g2_fill_2 FILLER_52_859 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_48 ();
 sg13g2_fill_1 FILLER_53_50 ();
 sg13g2_decap_4 FILLER_53_69 ();
 sg13g2_fill_2 FILLER_53_73 ();
 sg13g2_fill_2 FILLER_53_80 ();
 sg13g2_fill_2 FILLER_53_106 ();
 sg13g2_fill_1 FILLER_53_108 ();
 sg13g2_fill_1 FILLER_53_114 ();
 sg13g2_fill_1 FILLER_53_127 ();
 sg13g2_decap_4 FILLER_53_131 ();
 sg13g2_fill_2 FILLER_53_140 ();
 sg13g2_fill_2 FILLER_53_147 ();
 sg13g2_fill_1 FILLER_53_169 ();
 sg13g2_fill_2 FILLER_53_218 ();
 sg13g2_fill_1 FILLER_53_220 ();
 sg13g2_fill_1 FILLER_53_246 ();
 sg13g2_fill_1 FILLER_53_251 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_fill_1 FILLER_53_299 ();
 sg13g2_fill_2 FILLER_53_312 ();
 sg13g2_fill_1 FILLER_53_314 ();
 sg13g2_decap_4 FILLER_53_328 ();
 sg13g2_fill_1 FILLER_53_345 ();
 sg13g2_decap_4 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_53_358 ();
 sg13g2_decap_8 FILLER_53_363 ();
 sg13g2_decap_4 FILLER_53_370 ();
 sg13g2_fill_1 FILLER_53_374 ();
 sg13g2_fill_1 FILLER_53_385 ();
 sg13g2_fill_2 FILLER_53_390 ();
 sg13g2_fill_1 FILLER_53_392 ();
 sg13g2_decap_4 FILLER_53_405 ();
 sg13g2_decap_4 FILLER_53_413 ();
 sg13g2_fill_2 FILLER_53_417 ();
 sg13g2_fill_2 FILLER_53_423 ();
 sg13g2_fill_1 FILLER_53_425 ();
 sg13g2_fill_1 FILLER_53_513 ();
 sg13g2_fill_2 FILLER_53_530 ();
 sg13g2_fill_1 FILLER_53_532 ();
 sg13g2_fill_2 FILLER_53_559 ();
 sg13g2_fill_1 FILLER_53_561 ();
 sg13g2_decap_8 FILLER_53_570 ();
 sg13g2_decap_4 FILLER_53_577 ();
 sg13g2_fill_2 FILLER_53_597 ();
 sg13g2_fill_1 FILLER_53_599 ();
 sg13g2_fill_2 FILLER_53_615 ();
 sg13g2_fill_1 FILLER_53_617 ();
 sg13g2_fill_2 FILLER_53_622 ();
 sg13g2_fill_2 FILLER_53_632 ();
 sg13g2_fill_1 FILLER_53_634 ();
 sg13g2_decap_8 FILLER_53_688 ();
 sg13g2_decap_4 FILLER_53_695 ();
 sg13g2_fill_1 FILLER_53_699 ();
 sg13g2_fill_1 FILLER_53_721 ();
 sg13g2_decap_4 FILLER_53_731 ();
 sg13g2_fill_1 FILLER_53_735 ();
 sg13g2_fill_1 FILLER_53_757 ();
 sg13g2_decap_8 FILLER_53_778 ();
 sg13g2_decap_4 FILLER_53_785 ();
 sg13g2_fill_1 FILLER_53_789 ();
 sg13g2_decap_8 FILLER_53_805 ();
 sg13g2_fill_2 FILLER_53_836 ();
 sg13g2_decap_4 FILLER_53_854 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_2 ();
 sg13g2_fill_2 FILLER_54_17 ();
 sg13g2_fill_1 FILLER_54_19 ();
 sg13g2_fill_1 FILLER_54_41 ();
 sg13g2_fill_2 FILLER_54_50 ();
 sg13g2_decap_4 FILLER_54_101 ();
 sg13g2_fill_2 FILLER_54_125 ();
 sg13g2_decap_8 FILLER_54_142 ();
 sg13g2_fill_1 FILLER_54_167 ();
 sg13g2_fill_2 FILLER_54_172 ();
 sg13g2_fill_1 FILLER_54_179 ();
 sg13g2_fill_1 FILLER_54_185 ();
 sg13g2_decap_4 FILLER_54_216 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_fill_2 FILLER_54_241 ();
 sg13g2_fill_2 FILLER_54_252 ();
 sg13g2_fill_1 FILLER_54_254 ();
 sg13g2_fill_2 FILLER_54_315 ();
 sg13g2_fill_1 FILLER_54_317 ();
 sg13g2_fill_1 FILLER_54_344 ();
 sg13g2_fill_2 FILLER_54_409 ();
 sg13g2_fill_1 FILLER_54_411 ();
 sg13g2_decap_4 FILLER_54_420 ();
 sg13g2_decap_8 FILLER_54_436 ();
 sg13g2_fill_2 FILLER_54_443 ();
 sg13g2_fill_1 FILLER_54_445 ();
 sg13g2_fill_1 FILLER_54_449 ();
 sg13g2_fill_1 FILLER_54_463 ();
 sg13g2_fill_1 FILLER_54_507 ();
 sg13g2_fill_2 FILLER_54_557 ();
 sg13g2_decap_4 FILLER_54_583 ();
 sg13g2_fill_2 FILLER_54_601 ();
 sg13g2_fill_1 FILLER_54_603 ();
 sg13g2_fill_2 FILLER_54_644 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_2 FILLER_54_655 ();
 sg13g2_fill_2 FILLER_54_669 ();
 sg13g2_fill_1 FILLER_54_671 ();
 sg13g2_fill_2 FILLER_54_683 ();
 sg13g2_fill_1 FILLER_54_685 ();
 sg13g2_decap_8 FILLER_54_701 ();
 sg13g2_fill_1 FILLER_54_708 ();
 sg13g2_decap_8 FILLER_54_820 ();
 sg13g2_decap_4 FILLER_54_827 ();
 sg13g2_fill_1 FILLER_54_831 ();
 sg13g2_fill_1 FILLER_54_861 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_4 ();
 sg13g2_fill_1 FILLER_55_83 ();
 sg13g2_fill_2 FILLER_55_115 ();
 sg13g2_fill_1 FILLER_55_122 ();
 sg13g2_fill_1 FILLER_55_128 ();
 sg13g2_fill_2 FILLER_55_168 ();
 sg13g2_decap_4 FILLER_55_183 ();
 sg13g2_fill_1 FILLER_55_190 ();
 sg13g2_fill_2 FILLER_55_207 ();
 sg13g2_fill_2 FILLER_55_217 ();
 sg13g2_fill_2 FILLER_55_264 ();
 sg13g2_fill_2 FILLER_55_306 ();
 sg13g2_decap_4 FILLER_55_312 ();
 sg13g2_fill_1 FILLER_55_316 ();
 sg13g2_decap_8 FILLER_55_338 ();
 sg13g2_decap_4 FILLER_55_345 ();
 sg13g2_fill_2 FILLER_55_377 ();
 sg13g2_fill_1 FILLER_55_379 ();
 sg13g2_decap_4 FILLER_55_394 ();
 sg13g2_fill_2 FILLER_55_398 ();
 sg13g2_decap_8 FILLER_55_439 ();
 sg13g2_decap_4 FILLER_55_446 ();
 sg13g2_fill_2 FILLER_55_464 ();
 sg13g2_fill_2 FILLER_55_480 ();
 sg13g2_fill_1 FILLER_55_482 ();
 sg13g2_fill_2 FILLER_55_554 ();
 sg13g2_fill_2 FILLER_55_608 ();
 sg13g2_fill_2 FILLER_55_667 ();
 sg13g2_fill_2 FILLER_55_678 ();
 sg13g2_decap_8 FILLER_55_699 ();
 sg13g2_fill_2 FILLER_55_706 ();
 sg13g2_decap_4 FILLER_55_733 ();
 sg13g2_fill_2 FILLER_55_745 ();
 sg13g2_fill_1 FILLER_55_747 ();
 sg13g2_fill_2 FILLER_55_760 ();
 sg13g2_fill_1 FILLER_55_762 ();
 sg13g2_fill_2 FILLER_55_788 ();
 sg13g2_fill_2 FILLER_55_811 ();
 sg13g2_fill_1 FILLER_55_813 ();
 sg13g2_decap_4 FILLER_55_830 ();
 sg13g2_decap_4 FILLER_55_858 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_37 ();
 sg13g2_fill_1 FILLER_56_105 ();
 sg13g2_decap_4 FILLER_56_149 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_185 ();
 sg13g2_fill_2 FILLER_56_222 ();
 sg13g2_fill_2 FILLER_56_232 ();
 sg13g2_decap_4 FILLER_56_251 ();
 sg13g2_fill_2 FILLER_56_255 ();
 sg13g2_fill_2 FILLER_56_297 ();
 sg13g2_fill_1 FILLER_56_299 ();
 sg13g2_fill_1 FILLER_56_309 ();
 sg13g2_decap_8 FILLER_56_318 ();
 sg13g2_decap_8 FILLER_56_325 ();
 sg13g2_decap_8 FILLER_56_340 ();
 sg13g2_fill_2 FILLER_56_347 ();
 sg13g2_fill_2 FILLER_56_354 ();
 sg13g2_fill_2 FILLER_56_369 ();
 sg13g2_fill_1 FILLER_56_371 ();
 sg13g2_fill_2 FILLER_56_421 ();
 sg13g2_fill_1 FILLER_56_423 ();
 sg13g2_fill_2 FILLER_56_451 ();
 sg13g2_fill_1 FILLER_56_453 ();
 sg13g2_fill_1 FILLER_56_466 ();
 sg13g2_fill_2 FILLER_56_475 ();
 sg13g2_fill_1 FILLER_56_477 ();
 sg13g2_fill_1 FILLER_56_483 ();
 sg13g2_fill_2 FILLER_56_493 ();
 sg13g2_fill_1 FILLER_56_504 ();
 sg13g2_fill_2 FILLER_56_510 ();
 sg13g2_fill_2 FILLER_56_521 ();
 sg13g2_fill_1 FILLER_56_523 ();
 sg13g2_fill_1 FILLER_56_588 ();
 sg13g2_fill_1 FILLER_56_603 ();
 sg13g2_decap_8 FILLER_56_624 ();
 sg13g2_decap_4 FILLER_56_631 ();
 sg13g2_fill_2 FILLER_56_650 ();
 sg13g2_decap_8 FILLER_56_668 ();
 sg13g2_fill_2 FILLER_56_675 ();
 sg13g2_fill_1 FILLER_56_677 ();
 sg13g2_fill_2 FILLER_56_706 ();
 sg13g2_fill_1 FILLER_56_708 ();
 sg13g2_fill_1 FILLER_56_714 ();
 sg13g2_decap_4 FILLER_56_725 ();
 sg13g2_fill_1 FILLER_56_729 ();
 sg13g2_decap_8 FILLER_56_741 ();
 sg13g2_fill_1 FILLER_56_748 ();
 sg13g2_fill_1 FILLER_56_759 ();
 sg13g2_fill_2 FILLER_56_776 ();
 sg13g2_fill_2 FILLER_56_786 ();
 sg13g2_fill_1 FILLER_56_813 ();
 sg13g2_fill_1 FILLER_56_861 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_2 FILLER_57_21 ();
 sg13g2_fill_2 FILLER_57_33 ();
 sg13g2_fill_2 FILLER_57_40 ();
 sg13g2_fill_1 FILLER_57_42 ();
 sg13g2_fill_2 FILLER_57_48 ();
 sg13g2_fill_1 FILLER_57_50 ();
 sg13g2_fill_2 FILLER_57_91 ();
 sg13g2_fill_1 FILLER_57_93 ();
 sg13g2_fill_1 FILLER_57_110 ();
 sg13g2_fill_1 FILLER_57_119 ();
 sg13g2_fill_2 FILLER_57_148 ();
 sg13g2_fill_1 FILLER_57_150 ();
 sg13g2_fill_1 FILLER_57_169 ();
 sg13g2_fill_2 FILLER_57_182 ();
 sg13g2_fill_2 FILLER_57_193 ();
 sg13g2_fill_1 FILLER_57_195 ();
 sg13g2_decap_4 FILLER_57_200 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_4 FILLER_57_224 ();
 sg13g2_fill_2 FILLER_57_228 ();
 sg13g2_decap_8 FILLER_57_252 ();
 sg13g2_decap_4 FILLER_57_259 ();
 sg13g2_fill_2 FILLER_57_263 ();
 sg13g2_decap_8 FILLER_57_274 ();
 sg13g2_decap_4 FILLER_57_318 ();
 sg13g2_fill_2 FILLER_57_322 ();
 sg13g2_fill_1 FILLER_57_371 ();
 sg13g2_fill_2 FILLER_57_404 ();
 sg13g2_fill_1 FILLER_57_410 ();
 sg13g2_fill_2 FILLER_57_434 ();
 sg13g2_fill_1 FILLER_57_436 ();
 sg13g2_fill_2 FILLER_57_485 ();
 sg13g2_fill_1 FILLER_57_487 ();
 sg13g2_fill_2 FILLER_57_553 ();
 sg13g2_fill_1 FILLER_57_562 ();
 sg13g2_fill_1 FILLER_57_573 ();
 sg13g2_decap_8 FILLER_57_589 ();
 sg13g2_decap_8 FILLER_57_596 ();
 sg13g2_fill_2 FILLER_57_608 ();
 sg13g2_fill_1 FILLER_57_610 ();
 sg13g2_fill_1 FILLER_57_616 ();
 sg13g2_fill_1 FILLER_57_627 ();
 sg13g2_fill_1 FILLER_57_640 ();
 sg13g2_fill_1 FILLER_57_655 ();
 sg13g2_decap_8 FILLER_57_676 ();
 sg13g2_fill_2 FILLER_57_683 ();
 sg13g2_decap_4 FILLER_57_717 ();
 sg13g2_decap_8 FILLER_57_742 ();
 sg13g2_fill_2 FILLER_57_749 ();
 sg13g2_fill_1 FILLER_57_755 ();
 sg13g2_fill_2 FILLER_57_769 ();
 sg13g2_fill_2 FILLER_57_776 ();
 sg13g2_fill_2 FILLER_57_789 ();
 sg13g2_decap_8 FILLER_57_800 ();
 sg13g2_fill_1 FILLER_57_807 ();
 sg13g2_fill_2 FILLER_57_837 ();
 sg13g2_fill_1 FILLER_57_839 ();
 sg13g2_fill_1 FILLER_57_845 ();
 sg13g2_fill_2 FILLER_57_860 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_30 ();
 sg13g2_fill_1 FILLER_58_75 ();
 sg13g2_fill_2 FILLER_58_114 ();
 sg13g2_fill_2 FILLER_58_126 ();
 sg13g2_fill_2 FILLER_58_136 ();
 sg13g2_fill_1 FILLER_58_138 ();
 sg13g2_decap_4 FILLER_58_153 ();
 sg13g2_fill_1 FILLER_58_157 ();
 sg13g2_decap_4 FILLER_58_179 ();
 sg13g2_fill_2 FILLER_58_183 ();
 sg13g2_decap_8 FILLER_58_211 ();
 sg13g2_fill_1 FILLER_58_230 ();
 sg13g2_decap_8 FILLER_58_255 ();
 sg13g2_fill_1 FILLER_58_262 ();
 sg13g2_fill_1 FILLER_58_276 ();
 sg13g2_fill_2 FILLER_58_294 ();
 sg13g2_fill_1 FILLER_58_296 ();
 sg13g2_fill_1 FILLER_58_305 ();
 sg13g2_decap_4 FILLER_58_328 ();
 sg13g2_decap_8 FILLER_58_340 ();
 sg13g2_fill_2 FILLER_58_347 ();
 sg13g2_fill_2 FILLER_58_363 ();
 sg13g2_decap_4 FILLER_58_373 ();
 sg13g2_fill_2 FILLER_58_385 ();
 sg13g2_fill_1 FILLER_58_421 ();
 sg13g2_fill_2 FILLER_58_456 ();
 sg13g2_fill_2 FILLER_58_469 ();
 sg13g2_fill_1 FILLER_58_471 ();
 sg13g2_fill_1 FILLER_58_502 ();
 sg13g2_fill_2 FILLER_58_522 ();
 sg13g2_fill_2 FILLER_58_533 ();
 sg13g2_fill_2 FILLER_58_583 ();
 sg13g2_fill_2 FILLER_58_615 ();
 sg13g2_fill_2 FILLER_58_641 ();
 sg13g2_fill_2 FILLER_58_656 ();
 sg13g2_fill_1 FILLER_58_658 ();
 sg13g2_fill_2 FILLER_58_690 ();
 sg13g2_decap_4 FILLER_58_708 ();
 sg13g2_fill_1 FILLER_58_712 ();
 sg13g2_fill_1 FILLER_58_726 ();
 sg13g2_decap_4 FILLER_58_738 ();
 sg13g2_fill_1 FILLER_58_753 ();
 sg13g2_fill_2 FILLER_58_762 ();
 sg13g2_fill_2 FILLER_58_768 ();
 sg13g2_decap_4 FILLER_58_783 ();
 sg13g2_fill_2 FILLER_58_787 ();
 sg13g2_decap_4 FILLER_58_797 ();
 sg13g2_fill_2 FILLER_58_801 ();
 sg13g2_fill_2 FILLER_58_835 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_fill_1 FILLER_59_26 ();
 sg13g2_fill_2 FILLER_59_32 ();
 sg13g2_fill_1 FILLER_59_34 ();
 sg13g2_fill_2 FILLER_59_45 ();
 sg13g2_fill_1 FILLER_59_69 ();
 sg13g2_fill_2 FILLER_59_117 ();
 sg13g2_fill_1 FILLER_59_119 ();
 sg13g2_fill_2 FILLER_59_128 ();
 sg13g2_fill_2 FILLER_59_147 ();
 sg13g2_fill_1 FILLER_59_149 ();
 sg13g2_fill_2 FILLER_59_178 ();
 sg13g2_fill_2 FILLER_59_206 ();
 sg13g2_fill_1 FILLER_59_208 ();
 sg13g2_fill_2 FILLER_59_237 ();
 sg13g2_decap_4 FILLER_59_252 ();
 sg13g2_fill_1 FILLER_59_256 ();
 sg13g2_decap_8 FILLER_59_262 ();
 sg13g2_decap_4 FILLER_59_269 ();
 sg13g2_fill_2 FILLER_59_273 ();
 sg13g2_fill_1 FILLER_59_304 ();
 sg13g2_fill_2 FILLER_59_315 ();
 sg13g2_decap_8 FILLER_59_322 ();
 sg13g2_fill_2 FILLER_59_329 ();
 sg13g2_fill_1 FILLER_59_331 ();
 sg13g2_decap_4 FILLER_59_392 ();
 sg13g2_fill_2 FILLER_59_396 ();
 sg13g2_decap_4 FILLER_59_402 ();
 sg13g2_fill_1 FILLER_59_415 ();
 sg13g2_fill_1 FILLER_59_433 ();
 sg13g2_fill_1 FILLER_59_439 ();
 sg13g2_fill_2 FILLER_59_443 ();
 sg13g2_fill_1 FILLER_59_445 ();
 sg13g2_fill_2 FILLER_59_458 ();
 sg13g2_fill_2 FILLER_59_475 ();
 sg13g2_fill_1 FILLER_59_482 ();
 sg13g2_fill_2 FILLER_59_502 ();
 sg13g2_fill_1 FILLER_59_504 ();
 sg13g2_fill_1 FILLER_59_574 ();
 sg13g2_fill_1 FILLER_59_585 ();
 sg13g2_decap_4 FILLER_59_591 ();
 sg13g2_fill_2 FILLER_59_595 ();
 sg13g2_fill_1 FILLER_59_602 ();
 sg13g2_fill_2 FILLER_59_660 ();
 sg13g2_decap_8 FILLER_59_703 ();
 sg13g2_fill_2 FILLER_59_710 ();
 sg13g2_fill_1 FILLER_59_712 ();
 sg13g2_fill_2 FILLER_59_737 ();
 sg13g2_decap_8 FILLER_59_763 ();
 sg13g2_fill_1 FILLER_59_778 ();
 sg13g2_fill_2 FILLER_59_800 ();
 sg13g2_fill_1 FILLER_59_802 ();
 sg13g2_decap_4 FILLER_59_830 ();
 sg13g2_fill_2 FILLER_59_834 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_2 ();
 sg13g2_fill_2 FILLER_60_52 ();
 sg13g2_fill_1 FILLER_60_54 ();
 sg13g2_fill_2 FILLER_60_98 ();
 sg13g2_decap_4 FILLER_60_148 ();
 sg13g2_fill_1 FILLER_60_152 ();
 sg13g2_fill_2 FILLER_60_181 ();
 sg13g2_fill_1 FILLER_60_183 ();
 sg13g2_decap_4 FILLER_60_201 ();
 sg13g2_fill_1 FILLER_60_205 ();
 sg13g2_decap_8 FILLER_60_246 ();
 sg13g2_decap_4 FILLER_60_253 ();
 sg13g2_fill_1 FILLER_60_257 ();
 sg13g2_fill_2 FILLER_60_269 ();
 sg13g2_fill_2 FILLER_60_279 ();
 sg13g2_fill_1 FILLER_60_281 ();
 sg13g2_decap_4 FILLER_60_299 ();
 sg13g2_fill_1 FILLER_60_303 ();
 sg13g2_decap_4 FILLER_60_316 ();
 sg13g2_fill_2 FILLER_60_320 ();
 sg13g2_decap_4 FILLER_60_348 ();
 sg13g2_fill_1 FILLER_60_352 ();
 sg13g2_fill_2 FILLER_60_358 ();
 sg13g2_fill_1 FILLER_60_360 ();
 sg13g2_decap_8 FILLER_60_378 ();
 sg13g2_decap_8 FILLER_60_385 ();
 sg13g2_fill_2 FILLER_60_392 ();
 sg13g2_fill_2 FILLER_60_402 ();
 sg13g2_fill_2 FILLER_60_412 ();
 sg13g2_fill_1 FILLER_60_414 ();
 sg13g2_fill_1 FILLER_60_532 ();
 sg13g2_decap_4 FILLER_60_553 ();
 sg13g2_fill_2 FILLER_60_578 ();
 sg13g2_fill_1 FILLER_60_580 ();
 sg13g2_decap_4 FILLER_60_605 ();
 sg13g2_fill_2 FILLER_60_631 ();
 sg13g2_fill_1 FILLER_60_633 ();
 sg13g2_decap_8 FILLER_60_663 ();
 sg13g2_fill_1 FILLER_60_691 ();
 sg13g2_decap_4 FILLER_60_704 ();
 sg13g2_fill_1 FILLER_60_708 ();
 sg13g2_decap_4 FILLER_60_740 ();
 sg13g2_decap_4 FILLER_60_770 ();
 sg13g2_fill_2 FILLER_60_827 ();
 sg13g2_fill_2 FILLER_60_860 ();
 sg13g2_fill_2 FILLER_61_73 ();
 sg13g2_fill_2 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_fill_2 FILLER_61_127 ();
 sg13g2_decap_4 FILLER_61_141 ();
 sg13g2_fill_2 FILLER_61_145 ();
 sg13g2_decap_4 FILLER_61_151 ();
 sg13g2_fill_2 FILLER_61_155 ();
 sg13g2_fill_2 FILLER_61_162 ();
 sg13g2_fill_1 FILLER_61_173 ();
 sg13g2_decap_4 FILLER_61_200 ();
 sg13g2_fill_1 FILLER_61_204 ();
 sg13g2_fill_2 FILLER_61_218 ();
 sg13g2_fill_1 FILLER_61_220 ();
 sg13g2_decap_8 FILLER_61_245 ();
 sg13g2_decap_4 FILLER_61_252 ();
 sg13g2_fill_1 FILLER_61_256 ();
 sg13g2_decap_8 FILLER_61_291 ();
 sg13g2_fill_2 FILLER_61_298 ();
 sg13g2_decap_4 FILLER_61_313 ();
 sg13g2_fill_1 FILLER_61_317 ();
 sg13g2_fill_2 FILLER_61_322 ();
 sg13g2_fill_1 FILLER_61_324 ();
 sg13g2_fill_1 FILLER_61_332 ();
 sg13g2_fill_1 FILLER_61_345 ();
 sg13g2_decap_8 FILLER_61_354 ();
 sg13g2_decap_4 FILLER_61_361 ();
 sg13g2_fill_2 FILLER_61_365 ();
 sg13g2_fill_2 FILLER_61_391 ();
 sg13g2_decap_8 FILLER_61_425 ();
 sg13g2_fill_1 FILLER_61_432 ();
 sg13g2_fill_2 FILLER_61_437 ();
 sg13g2_fill_2 FILLER_61_443 ();
 sg13g2_fill_2 FILLER_61_471 ();
 sg13g2_fill_1 FILLER_61_473 ();
 sg13g2_fill_1 FILLER_61_479 ();
 sg13g2_fill_2 FILLER_61_489 ();
 sg13g2_fill_2 FILLER_61_495 ();
 sg13g2_fill_1 FILLER_61_497 ();
 sg13g2_fill_2 FILLER_61_502 ();
 sg13g2_fill_1 FILLER_61_504 ();
 sg13g2_fill_1 FILLER_61_517 ();
 sg13g2_fill_2 FILLER_61_541 ();
 sg13g2_fill_1 FILLER_61_556 ();
 sg13g2_decap_4 FILLER_61_572 ();
 sg13g2_fill_1 FILLER_61_576 ();
 sg13g2_fill_2 FILLER_61_605 ();
 sg13g2_fill_1 FILLER_61_607 ();
 sg13g2_fill_1 FILLER_61_613 ();
 sg13g2_fill_1 FILLER_61_627 ();
 sg13g2_decap_8 FILLER_61_649 ();
 sg13g2_fill_2 FILLER_61_656 ();
 sg13g2_fill_1 FILLER_61_658 ();
 sg13g2_fill_1 FILLER_61_667 ();
 sg13g2_decap_4 FILLER_61_676 ();
 sg13g2_fill_2 FILLER_61_680 ();
 sg13g2_fill_1 FILLER_61_686 ();
 sg13g2_fill_1 FILLER_61_738 ();
 sg13g2_fill_1 FILLER_61_753 ();
 sg13g2_fill_2 FILLER_61_770 ();
 sg13g2_decap_4 FILLER_61_790 ();
 sg13g2_decap_8 FILLER_61_823 ();
 sg13g2_decap_4 FILLER_61_830 ();
 sg13g2_fill_2 FILLER_61_834 ();
 sg13g2_decap_4 FILLER_61_857 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_1 FILLER_62_71 ();
 sg13g2_fill_1 FILLER_62_117 ();
 sg13g2_fill_2 FILLER_62_123 ();
 sg13g2_decap_4 FILLER_62_183 ();
 sg13g2_fill_1 FILLER_62_187 ();
 sg13g2_fill_2 FILLER_62_219 ();
 sg13g2_decap_8 FILLER_62_238 ();
 sg13g2_fill_2 FILLER_62_245 ();
 sg13g2_fill_1 FILLER_62_273 ();
 sg13g2_fill_2 FILLER_62_286 ();
 sg13g2_decap_4 FILLER_62_301 ();
 sg13g2_fill_2 FILLER_62_323 ();
 sg13g2_fill_2 FILLER_62_338 ();
 sg13g2_fill_1 FILLER_62_340 ();
 sg13g2_decap_4 FILLER_62_371 ();
 sg13g2_fill_1 FILLER_62_375 ();
 sg13g2_decap_4 FILLER_62_380 ();
 sg13g2_fill_2 FILLER_62_401 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_62_414 ();
 sg13g2_fill_1 FILLER_62_421 ();
 sg13g2_fill_1 FILLER_62_443 ();
 sg13g2_fill_1 FILLER_62_475 ();
 sg13g2_decap_8 FILLER_62_541 ();
 sg13g2_decap_4 FILLER_62_548 ();
 sg13g2_decap_8 FILLER_62_560 ();
 sg13g2_fill_2 FILLER_62_567 ();
 sg13g2_fill_1 FILLER_62_569 ();
 sg13g2_decap_8 FILLER_62_574 ();
 sg13g2_decap_4 FILLER_62_581 ();
 sg13g2_fill_1 FILLER_62_616 ();
 sg13g2_decap_8 FILLER_62_643 ();
 sg13g2_decap_4 FILLER_62_662 ();
 sg13g2_decap_4 FILLER_62_683 ();
 sg13g2_decap_4 FILLER_62_719 ();
 sg13g2_fill_2 FILLER_62_735 ();
 sg13g2_decap_4 FILLER_62_765 ();
 sg13g2_fill_1 FILLER_62_769 ();
 sg13g2_fill_2 FILLER_62_791 ();
 sg13g2_decap_4 FILLER_62_806 ();
 sg13g2_decap_4 FILLER_62_826 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_2 ();
 sg13g2_fill_2 FILLER_63_38 ();
 sg13g2_fill_1 FILLER_63_81 ();
 sg13g2_fill_1 FILLER_63_146 ();
 sg13g2_fill_1 FILLER_63_156 ();
 sg13g2_fill_1 FILLER_63_170 ();
 sg13g2_decap_4 FILLER_63_205 ();
 sg13g2_fill_1 FILLER_63_209 ();
 sg13g2_decap_4 FILLER_63_240 ();
 sg13g2_fill_1 FILLER_63_244 ();
 sg13g2_fill_1 FILLER_63_266 ();
 sg13g2_fill_2 FILLER_63_282 ();
 sg13g2_fill_2 FILLER_63_323 ();
 sg13g2_fill_1 FILLER_63_325 ();
 sg13g2_fill_1 FILLER_63_331 ();
 sg13g2_fill_2 FILLER_63_348 ();
 sg13g2_fill_1 FILLER_63_350 ();
 sg13g2_decap_4 FILLER_63_382 ();
 sg13g2_fill_1 FILLER_63_413 ();
 sg13g2_fill_2 FILLER_63_426 ();
 sg13g2_decap_4 FILLER_63_433 ();
 sg13g2_decap_4 FILLER_63_447 ();
 sg13g2_fill_1 FILLER_63_451 ();
 sg13g2_decap_8 FILLER_63_467 ();
 sg13g2_decap_8 FILLER_63_474 ();
 sg13g2_fill_1 FILLER_63_486 ();
 sg13g2_fill_1 FILLER_63_525 ();
 sg13g2_fill_2 FILLER_63_539 ();
 sg13g2_fill_1 FILLER_63_541 ();
 sg13g2_fill_1 FILLER_63_594 ();
 sg13g2_fill_2 FILLER_63_615 ();
 sg13g2_fill_1 FILLER_63_617 ();
 sg13g2_decap_4 FILLER_63_632 ();
 sg13g2_fill_1 FILLER_63_654 ();
 sg13g2_decap_8 FILLER_63_684 ();
 sg13g2_fill_2 FILLER_63_691 ();
 sg13g2_fill_1 FILLER_63_693 ();
 sg13g2_fill_1 FILLER_63_712 ();
 sg13g2_fill_1 FILLER_63_718 ();
 sg13g2_fill_2 FILLER_63_727 ();
 sg13g2_decap_4 FILLER_63_734 ();
 sg13g2_decap_4 FILLER_63_741 ();
 sg13g2_fill_1 FILLER_63_745 ();
 sg13g2_decap_4 FILLER_63_763 ();
 sg13g2_fill_1 FILLER_63_767 ();
 sg13g2_decap_4 FILLER_63_771 ();
 sg13g2_fill_1 FILLER_63_779 ();
 sg13g2_decap_8 FILLER_63_784 ();
 sg13g2_decap_8 FILLER_63_791 ();
 sg13g2_fill_1 FILLER_63_798 ();
 sg13g2_fill_2 FILLER_63_833 ();
 sg13g2_fill_2 FILLER_63_848 ();
 sg13g2_decap_8 FILLER_63_854 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_fill_2 FILLER_64_38 ();
 sg13g2_fill_2 FILLER_64_94 ();
 sg13g2_fill_2 FILLER_64_115 ();
 sg13g2_fill_2 FILLER_64_177 ();
 sg13g2_fill_1 FILLER_64_179 ();
 sg13g2_decap_8 FILLER_64_206 ();
 sg13g2_fill_2 FILLER_64_213 ();
 sg13g2_fill_1 FILLER_64_215 ();
 sg13g2_fill_1 FILLER_64_219 ();
 sg13g2_fill_2 FILLER_64_248 ();
 sg13g2_decap_4 FILLER_64_268 ();
 sg13g2_fill_2 FILLER_64_301 ();
 sg13g2_fill_1 FILLER_64_303 ();
 sg13g2_fill_2 FILLER_64_314 ();
 sg13g2_fill_1 FILLER_64_316 ();
 sg13g2_decap_8 FILLER_64_333 ();
 sg13g2_fill_1 FILLER_64_353 ();
 sg13g2_fill_2 FILLER_64_366 ();
 sg13g2_fill_1 FILLER_64_368 ();
 sg13g2_decap_4 FILLER_64_385 ();
 sg13g2_fill_2 FILLER_64_389 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_2 FILLER_64_422 ();
 sg13g2_fill_2 FILLER_64_439 ();
 sg13g2_fill_2 FILLER_64_458 ();
 sg13g2_decap_4 FILLER_64_465 ();
 sg13g2_fill_1 FILLER_64_499 ();
 sg13g2_fill_2 FILLER_64_503 ();
 sg13g2_fill_1 FILLER_64_505 ();
 sg13g2_fill_2 FILLER_64_514 ();
 sg13g2_fill_1 FILLER_64_516 ();
 sg13g2_decap_8 FILLER_64_546 ();
 sg13g2_decap_8 FILLER_64_553 ();
 sg13g2_fill_1 FILLER_64_578 ();
 sg13g2_fill_2 FILLER_64_583 ();
 sg13g2_fill_2 FILLER_64_595 ();
 sg13g2_fill_2 FILLER_64_610 ();
 sg13g2_fill_1 FILLER_64_625 ();
 sg13g2_fill_1 FILLER_64_666 ();
 sg13g2_decap_8 FILLER_64_675 ();
 sg13g2_fill_2 FILLER_64_682 ();
 sg13g2_fill_2 FILLER_64_717 ();
 sg13g2_decap_8 FILLER_64_765 ();
 sg13g2_fill_1 FILLER_64_772 ();
 sg13g2_fill_2 FILLER_64_794 ();
 sg13g2_decap_4 FILLER_64_814 ();
 sg13g2_fill_1 FILLER_64_818 ();
 sg13g2_decap_4 FILLER_64_835 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_fill_1 FILLER_65_59 ();
 sg13g2_fill_1 FILLER_65_68 ();
 sg13g2_fill_1 FILLER_65_135 ();
 sg13g2_fill_1 FILLER_65_141 ();
 sg13g2_fill_2 FILLER_65_151 ();
 sg13g2_fill_2 FILLER_65_179 ();
 sg13g2_fill_1 FILLER_65_181 ();
 sg13g2_decap_8 FILLER_65_203 ();
 sg13g2_fill_2 FILLER_65_210 ();
 sg13g2_fill_1 FILLER_65_212 ();
 sg13g2_fill_1 FILLER_65_243 ();
 sg13g2_decap_4 FILLER_65_265 ();
 sg13g2_fill_2 FILLER_65_285 ();
 sg13g2_decap_4 FILLER_65_297 ();
 sg13g2_fill_2 FILLER_65_337 ();
 sg13g2_fill_1 FILLER_65_339 ();
 sg13g2_fill_1 FILLER_65_352 ();
 sg13g2_decap_8 FILLER_65_363 ();
 sg13g2_fill_2 FILLER_65_370 ();
 sg13g2_fill_1 FILLER_65_372 ();
 sg13g2_decap_4 FILLER_65_377 ();
 sg13g2_fill_1 FILLER_65_381 ();
 sg13g2_fill_2 FILLER_65_390 ();
 sg13g2_fill_1 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_401 ();
 sg13g2_fill_2 FILLER_65_408 ();
 sg13g2_decap_4 FILLER_65_418 ();
 sg13g2_decap_4 FILLER_65_426 ();
 sg13g2_fill_2 FILLER_65_440 ();
 sg13g2_decap_4 FILLER_65_458 ();
 sg13g2_fill_1 FILLER_65_462 ();
 sg13g2_decap_4 FILLER_65_471 ();
 sg13g2_fill_1 FILLER_65_475 ();
 sg13g2_decap_8 FILLER_65_491 ();
 sg13g2_decap_4 FILLER_65_524 ();
 sg13g2_fill_1 FILLER_65_532 ();
 sg13g2_fill_1 FILLER_65_565 ();
 sg13g2_fill_1 FILLER_65_595 ();
 sg13g2_decap_4 FILLER_65_617 ();
 sg13g2_fill_2 FILLER_65_621 ();
 sg13g2_decap_8 FILLER_65_635 ();
 sg13g2_fill_2 FILLER_65_642 ();
 sg13g2_decap_8 FILLER_65_654 ();
 sg13g2_decap_4 FILLER_65_661 ();
 sg13g2_decap_8 FILLER_65_683 ();
 sg13g2_fill_1 FILLER_65_690 ();
 sg13g2_fill_1 FILLER_65_712 ();
 sg13g2_fill_1 FILLER_65_718 ();
 sg13g2_decap_4 FILLER_65_740 ();
 sg13g2_fill_1 FILLER_65_744 ();
 sg13g2_fill_1 FILLER_65_755 ();
 sg13g2_fill_1 FILLER_65_762 ();
 sg13g2_fill_2 FILLER_65_769 ();
 sg13g2_fill_1 FILLER_65_797 ();
 sg13g2_decap_8 FILLER_65_811 ();
 sg13g2_fill_1 FILLER_65_818 ();
 sg13g2_fill_1 FILLER_66_62 ();
 sg13g2_fill_1 FILLER_66_87 ();
 sg13g2_fill_2 FILLER_66_166 ();
 sg13g2_fill_1 FILLER_66_168 ();
 sg13g2_fill_1 FILLER_66_191 ();
 sg13g2_fill_2 FILLER_66_275 ();
 sg13g2_fill_1 FILLER_66_277 ();
 sg13g2_decap_8 FILLER_66_298 ();
 sg13g2_decap_8 FILLER_66_305 ();
 sg13g2_fill_1 FILLER_66_326 ();
 sg13g2_fill_2 FILLER_66_352 ();
 sg13g2_fill_1 FILLER_66_354 ();
 sg13g2_decap_4 FILLER_66_365 ();
 sg13g2_fill_1 FILLER_66_369 ();
 sg13g2_fill_2 FILLER_66_375 ();
 sg13g2_fill_1 FILLER_66_409 ();
 sg13g2_decap_4 FILLER_66_428 ();
 sg13g2_fill_2 FILLER_66_437 ();
 sg13g2_fill_2 FILLER_66_444 ();
 sg13g2_decap_4 FILLER_66_456 ();
 sg13g2_fill_1 FILLER_66_460 ();
 sg13g2_decap_8 FILLER_66_503 ();
 sg13g2_decap_8 FILLER_66_510 ();
 sg13g2_decap_4 FILLER_66_517 ();
 sg13g2_fill_1 FILLER_66_521 ();
 sg13g2_decap_4 FILLER_66_563 ();
 sg13g2_fill_2 FILLER_66_567 ();
 sg13g2_fill_2 FILLER_66_577 ();
 sg13g2_fill_1 FILLER_66_579 ();
 sg13g2_fill_2 FILLER_66_590 ();
 sg13g2_decap_8 FILLER_66_602 ();
 sg13g2_decap_8 FILLER_66_609 ();
 sg13g2_decap_4 FILLER_66_616 ();
 sg13g2_fill_1 FILLER_66_620 ();
 sg13g2_fill_2 FILLER_66_639 ();
 sg13g2_fill_2 FILLER_66_649 ();
 sg13g2_fill_1 FILLER_66_651 ();
 sg13g2_decap_4 FILLER_66_690 ();
 sg13g2_fill_1 FILLER_66_694 ();
 sg13g2_fill_2 FILLER_66_707 ();
 sg13g2_fill_1 FILLER_66_709 ();
 sg13g2_fill_2 FILLER_66_722 ();
 sg13g2_decap_8 FILLER_66_769 ();
 sg13g2_decap_8 FILLER_66_776 ();
 sg13g2_fill_1 FILLER_66_783 ();
 sg13g2_fill_1 FILLER_66_797 ();
 sg13g2_decap_4 FILLER_66_834 ();
 sg13g2_fill_2 FILLER_66_846 ();
 sg13g2_fill_1 FILLER_66_861 ();
 sg13g2_fill_1 FILLER_67_44 ();
 sg13g2_fill_1 FILLER_67_50 ();
 sg13g2_decap_8 FILLER_67_137 ();
 sg13g2_fill_1 FILLER_67_192 ();
 sg13g2_fill_1 FILLER_67_205 ();
 sg13g2_fill_2 FILLER_67_249 ();
 sg13g2_decap_8 FILLER_67_271 ();
 sg13g2_fill_1 FILLER_67_278 ();
 sg13g2_fill_1 FILLER_67_289 ();
 sg13g2_decap_8 FILLER_67_295 ();
 sg13g2_decap_8 FILLER_67_302 ();
 sg13g2_fill_2 FILLER_67_309 ();
 sg13g2_fill_1 FILLER_67_311 ();
 sg13g2_decap_4 FILLER_67_320 ();
 sg13g2_fill_1 FILLER_67_324 ();
 sg13g2_fill_2 FILLER_67_373 ();
 sg13g2_fill_1 FILLER_67_375 ();
 sg13g2_decap_4 FILLER_67_389 ();
 sg13g2_fill_1 FILLER_67_413 ();
 sg13g2_decap_4 FILLER_67_422 ();
 sg13g2_fill_2 FILLER_67_434 ();
 sg13g2_fill_1 FILLER_67_436 ();
 sg13g2_decap_8 FILLER_67_463 ();
 sg13g2_fill_2 FILLER_67_470 ();
 sg13g2_fill_1 FILLER_67_491 ();
 sg13g2_decap_8 FILLER_67_507 ();
 sg13g2_fill_2 FILLER_67_514 ();
 sg13g2_fill_1 FILLER_67_521 ();
 sg13g2_fill_1 FILLER_67_546 ();
 sg13g2_fill_1 FILLER_67_579 ();
 sg13g2_decap_8 FILLER_67_590 ();
 sg13g2_fill_2 FILLER_67_597 ();
 sg13g2_fill_2 FILLER_67_617 ();
 sg13g2_fill_1 FILLER_67_670 ();
 sg13g2_decap_8 FILLER_67_680 ();
 sg13g2_fill_1 FILLER_67_687 ();
 sg13g2_fill_2 FILLER_67_729 ();
 sg13g2_decap_4 FILLER_67_744 ();
 sg13g2_fill_1 FILLER_67_762 ();
 sg13g2_fill_1 FILLER_67_771 ();
 sg13g2_decap_4 FILLER_67_793 ();
 sg13g2_fill_1 FILLER_67_797 ();
 sg13g2_decap_4 FILLER_67_802 ();
 sg13g2_decap_4 FILLER_67_826 ();
 sg13g2_fill_1 FILLER_67_830 ();
 sg13g2_fill_2 FILLER_67_843 ();
 sg13g2_fill_2 FILLER_67_860 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_22 ();
 sg13g2_fill_2 FILLER_68_32 ();
 sg13g2_fill_1 FILLER_68_39 ();
 sg13g2_fill_1 FILLER_68_63 ();
 sg13g2_fill_2 FILLER_68_68 ();
 sg13g2_fill_1 FILLER_68_137 ();
 sg13g2_fill_2 FILLER_68_181 ();
 sg13g2_fill_1 FILLER_68_183 ();
 sg13g2_decap_4 FILLER_68_220 ();
 sg13g2_fill_2 FILLER_68_224 ();
 sg13g2_fill_2 FILLER_68_241 ();
 sg13g2_fill_1 FILLER_68_243 ();
 sg13g2_decap_8 FILLER_68_275 ();
 sg13g2_decap_8 FILLER_68_282 ();
 sg13g2_fill_2 FILLER_68_289 ();
 sg13g2_fill_2 FILLER_68_333 ();
 sg13g2_fill_1 FILLER_68_343 ();
 sg13g2_decap_8 FILLER_68_359 ();
 sg13g2_fill_2 FILLER_68_366 ();
 sg13g2_fill_1 FILLER_68_368 ();
 sg13g2_fill_1 FILLER_68_385 ();
 sg13g2_decap_8 FILLER_68_394 ();
 sg13g2_fill_2 FILLER_68_405 ();
 sg13g2_fill_1 FILLER_68_407 ();
 sg13g2_fill_2 FILLER_68_416 ();
 sg13g2_fill_1 FILLER_68_418 ();
 sg13g2_fill_1 FILLER_68_432 ();
 sg13g2_decap_4 FILLER_68_441 ();
 sg13g2_fill_2 FILLER_68_458 ();
 sg13g2_fill_1 FILLER_68_460 ();
 sg13g2_fill_1 FILLER_68_502 ();
 sg13g2_fill_1 FILLER_68_538 ();
 sg13g2_decap_4 FILLER_68_555 ();
 sg13g2_fill_2 FILLER_68_567 ();
 sg13g2_fill_2 FILLER_68_594 ();
 sg13g2_fill_1 FILLER_68_596 ();
 sg13g2_decap_8 FILLER_68_647 ();
 sg13g2_decap_8 FILLER_68_684 ();
 sg13g2_decap_4 FILLER_68_691 ();
 sg13g2_fill_1 FILLER_68_695 ();
 sg13g2_decap_4 FILLER_68_707 ();
 sg13g2_fill_1 FILLER_68_711 ();
 sg13g2_decap_8 FILLER_68_721 ();
 sg13g2_fill_1 FILLER_68_728 ();
 sg13g2_fill_2 FILLER_68_753 ();
 sg13g2_fill_2 FILLER_68_780 ();
 sg13g2_decap_8 FILLER_68_786 ();
 sg13g2_fill_1 FILLER_68_793 ();
 sg13g2_fill_2 FILLER_68_802 ();
 sg13g2_fill_1 FILLER_68_804 ();
 sg13g2_decap_8 FILLER_68_821 ();
 sg13g2_fill_1 FILLER_68_828 ();
 sg13g2_fill_1 FILLER_68_841 ();
 sg13g2_fill_1 FILLER_68_847 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_fill_1 FILLER_69_35 ();
 sg13g2_fill_2 FILLER_69_64 ();
 sg13g2_fill_2 FILLER_69_80 ();
 sg13g2_decap_4 FILLER_69_130 ();
 sg13g2_fill_1 FILLER_69_134 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_decap_8 FILLER_69_215 ();
 sg13g2_decap_8 FILLER_69_222 ();
 sg13g2_decap_8 FILLER_69_229 ();
 sg13g2_fill_2 FILLER_69_236 ();
 sg13g2_fill_2 FILLER_69_246 ();
 sg13g2_fill_1 FILLER_69_267 ();
 sg13g2_decap_8 FILLER_69_276 ();
 sg13g2_fill_2 FILLER_69_283 ();
 sg13g2_fill_1 FILLER_69_285 ();
 sg13g2_decap_4 FILLER_69_302 ();
 sg13g2_fill_2 FILLER_69_306 ();
 sg13g2_fill_1 FILLER_69_333 ();
 sg13g2_decap_4 FILLER_69_347 ();
 sg13g2_fill_1 FILLER_69_351 ();
 sg13g2_fill_2 FILLER_69_371 ();
 sg13g2_fill_1 FILLER_69_373 ();
 sg13g2_fill_2 FILLER_69_379 ();
 sg13g2_fill_1 FILLER_69_381 ();
 sg13g2_fill_1 FILLER_69_390 ();
 sg13g2_fill_2 FILLER_69_404 ();
 sg13g2_fill_1 FILLER_69_406 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_fill_1 FILLER_69_435 ();
 sg13g2_decap_8 FILLER_69_462 ();
 sg13g2_fill_2 FILLER_69_469 ();
 sg13g2_fill_1 FILLER_69_471 ();
 sg13g2_fill_2 FILLER_69_481 ();
 sg13g2_fill_2 FILLER_69_491 ();
 sg13g2_fill_1 FILLER_69_493 ();
 sg13g2_decap_4 FILLER_69_544 ();
 sg13g2_fill_1 FILLER_69_548 ();
 sg13g2_fill_2 FILLER_69_561 ();
 sg13g2_fill_1 FILLER_69_563 ();
 sg13g2_fill_2 FILLER_69_579 ();
 sg13g2_fill_1 FILLER_69_581 ();
 sg13g2_decap_8 FILLER_69_585 ();
 sg13g2_decap_8 FILLER_69_592 ();
 sg13g2_fill_1 FILLER_69_599 ();
 sg13g2_decap_8 FILLER_69_611 ();
 sg13g2_decap_4 FILLER_69_618 ();
 sg13g2_fill_1 FILLER_69_622 ();
 sg13g2_fill_2 FILLER_69_628 ();
 sg13g2_fill_1 FILLER_69_630 ();
 sg13g2_decap_8 FILLER_69_656 ();
 sg13g2_fill_2 FILLER_69_663 ();
 sg13g2_decap_8 FILLER_69_694 ();
 sg13g2_fill_2 FILLER_69_701 ();
 sg13g2_decap_4 FILLER_69_728 ();
 sg13g2_fill_2 FILLER_69_732 ();
 sg13g2_fill_2 FILLER_69_762 ();
 sg13g2_fill_1 FILLER_69_764 ();
 sg13g2_fill_2 FILLER_69_794 ();
 sg13g2_decap_4 FILLER_69_804 ();
 sg13g2_decap_4 FILLER_69_831 ();
 sg13g2_fill_1 FILLER_69_835 ();
 sg13g2_fill_2 FILLER_69_860 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_2 ();
 sg13g2_fill_1 FILLER_70_56 ();
 sg13g2_fill_2 FILLER_70_67 ();
 sg13g2_fill_1 FILLER_70_109 ();
 sg13g2_fill_2 FILLER_70_127 ();
 sg13g2_decap_4 FILLER_70_145 ();
 sg13g2_fill_2 FILLER_70_149 ();
 sg13g2_fill_2 FILLER_70_155 ();
 sg13g2_fill_1 FILLER_70_157 ();
 sg13g2_fill_2 FILLER_70_170 ();
 sg13g2_fill_1 FILLER_70_207 ();
 sg13g2_decap_8 FILLER_70_234 ();
 sg13g2_fill_2 FILLER_70_241 ();
 sg13g2_fill_1 FILLER_70_243 ();
 sg13g2_fill_2 FILLER_70_287 ();
 sg13g2_fill_2 FILLER_70_329 ();
 sg13g2_fill_2 FILLER_70_339 ();
 sg13g2_fill_1 FILLER_70_369 ();
 sg13g2_fill_1 FILLER_70_378 ();
 sg13g2_fill_2 FILLER_70_383 ();
 sg13g2_fill_2 FILLER_70_402 ();
 sg13g2_fill_1 FILLER_70_404 ();
 sg13g2_decap_8 FILLER_70_413 ();
 sg13g2_fill_2 FILLER_70_425 ();
 sg13g2_decap_4 FILLER_70_439 ();
 sg13g2_fill_1 FILLER_70_443 ();
 sg13g2_decap_4 FILLER_70_456 ();
 sg13g2_fill_2 FILLER_70_460 ();
 sg13g2_decap_4 FILLER_70_482 ();
 sg13g2_fill_2 FILLER_70_486 ();
 sg13g2_fill_1 FILLER_70_496 ();
 sg13g2_fill_2 FILLER_70_504 ();
 sg13g2_decap_8 FILLER_70_513 ();
 sg13g2_fill_2 FILLER_70_520 ();
 sg13g2_fill_1 FILLER_70_522 ();
 sg13g2_fill_1 FILLER_70_540 ();
 sg13g2_decap_4 FILLER_70_559 ();
 sg13g2_fill_1 FILLER_70_563 ();
 sg13g2_decap_4 FILLER_70_569 ();
 sg13g2_decap_8 FILLER_70_617 ();
 sg13g2_fill_2 FILLER_70_624 ();
 sg13g2_fill_1 FILLER_70_626 ();
 sg13g2_fill_1 FILLER_70_649 ();
 sg13g2_fill_2 FILLER_70_658 ();
 sg13g2_fill_1 FILLER_70_660 ();
 sg13g2_fill_2 FILLER_70_678 ();
 sg13g2_fill_1 FILLER_70_680 ();
 sg13g2_decap_8 FILLER_70_693 ();
 sg13g2_fill_2 FILLER_70_700 ();
 sg13g2_decap_8 FILLER_70_735 ();
 sg13g2_decap_4 FILLER_70_752 ();
 sg13g2_fill_2 FILLER_70_756 ();
 sg13g2_decap_4 FILLER_70_784 ();
 sg13g2_fill_2 FILLER_70_788 ();
 sg13g2_decap_4 FILLER_70_798 ();
 sg13g2_fill_1 FILLER_70_802 ();
 sg13g2_decap_4 FILLER_70_838 ();
 sg13g2_fill_1 FILLER_70_842 ();
 sg13g2_fill_2 FILLER_70_860 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_28 ();
 sg13g2_fill_1 FILLER_71_71 ();
 sg13g2_fill_1 FILLER_71_77 ();
 sg13g2_fill_2 FILLER_71_139 ();
 sg13g2_decap_8 FILLER_71_145 ();
 sg13g2_fill_2 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_251 ();
 sg13g2_fill_2 FILLER_71_283 ();
 sg13g2_decap_4 FILLER_71_321 ();
 sg13g2_decap_4 FILLER_71_341 ();
 sg13g2_fill_2 FILLER_71_345 ();
 sg13g2_decap_4 FILLER_71_354 ();
 sg13g2_fill_2 FILLER_71_358 ();
 sg13g2_decap_8 FILLER_71_372 ();
 sg13g2_fill_1 FILLER_71_379 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_fill_1 FILLER_71_409 ();
 sg13g2_decap_4 FILLER_71_435 ();
 sg13g2_fill_2 FILLER_71_439 ();
 sg13g2_fill_2 FILLER_71_467 ();
 sg13g2_fill_1 FILLER_71_469 ();
 sg13g2_decap_4 FILLER_71_482 ();
 sg13g2_fill_2 FILLER_71_486 ();
 sg13g2_fill_1 FILLER_71_501 ();
 sg13g2_fill_1 FILLER_71_510 ();
 sg13g2_fill_2 FILLER_71_516 ();
 sg13g2_decap_4 FILLER_71_530 ();
 sg13g2_fill_1 FILLER_71_534 ();
 sg13g2_decap_8 FILLER_71_640 ();
 sg13g2_fill_1 FILLER_71_672 ();
 sg13g2_decap_8 FILLER_71_699 ();
 sg13g2_decap_4 FILLER_71_706 ();
 sg13g2_fill_2 FILLER_71_710 ();
 sg13g2_fill_1 FILLER_71_742 ();
 sg13g2_fill_2 FILLER_71_774 ();
 sg13g2_fill_1 FILLER_71_776 ();
 sg13g2_fill_2 FILLER_71_785 ();
 sg13g2_fill_1 FILLER_71_816 ();
 sg13g2_fill_1 FILLER_71_835 ();
 sg13g2_fill_1 FILLER_72_48 ();
 sg13g2_fill_2 FILLER_72_89 ();
 sg13g2_fill_1 FILLER_72_95 ();
 sg13g2_fill_1 FILLER_72_109 ();
 sg13g2_fill_2 FILLER_72_125 ();
 sg13g2_fill_1 FILLER_72_127 ();
 sg13g2_fill_1 FILLER_72_158 ();
 sg13g2_fill_2 FILLER_72_178 ();
 sg13g2_fill_2 FILLER_72_212 ();
 sg13g2_decap_8 FILLER_72_244 ();
 sg13g2_fill_2 FILLER_72_251 ();
 sg13g2_decap_4 FILLER_72_279 ();
 sg13g2_fill_1 FILLER_72_326 ();
 sg13g2_fill_2 FILLER_72_340 ();
 sg13g2_fill_2 FILLER_72_366 ();
 sg13g2_fill_1 FILLER_72_368 ();
 sg13g2_fill_1 FILLER_72_382 ();
 sg13g2_fill_2 FILLER_72_387 ();
 sg13g2_decap_8 FILLER_72_405 ();
 sg13g2_decap_4 FILLER_72_412 ();
 sg13g2_fill_2 FILLER_72_416 ();
 sg13g2_decap_8 FILLER_72_427 ();
 sg13g2_decap_8 FILLER_72_434 ();
 sg13g2_decap_4 FILLER_72_441 ();
 sg13g2_fill_1 FILLER_72_503 ();
 sg13g2_decap_8 FILLER_72_529 ();
 sg13g2_fill_1 FILLER_72_536 ();
 sg13g2_decap_8 FILLER_72_546 ();
 sg13g2_decap_4 FILLER_72_553 ();
 sg13g2_fill_2 FILLER_72_557 ();
 sg13g2_fill_2 FILLER_72_567 ();
 sg13g2_fill_1 FILLER_72_569 ();
 sg13g2_fill_2 FILLER_72_585 ();
 sg13g2_fill_1 FILLER_72_603 ();
 sg13g2_fill_1 FILLER_72_622 ();
 sg13g2_fill_1 FILLER_72_631 ();
 sg13g2_fill_2 FILLER_72_649 ();
 sg13g2_fill_1 FILLER_72_651 ();
 sg13g2_decap_4 FILLER_72_657 ();
 sg13g2_fill_2 FILLER_72_689 ();
 sg13g2_fill_1 FILLER_72_691 ();
 sg13g2_decap_8 FILLER_72_725 ();
 sg13g2_fill_2 FILLER_72_732 ();
 sg13g2_decap_8 FILLER_72_743 ();
 sg13g2_fill_1 FILLER_72_766 ();
 sg13g2_fill_2 FILLER_72_787 ();
 sg13g2_fill_1 FILLER_72_789 ();
 sg13g2_decap_8 FILLER_72_798 ();
 sg13g2_fill_2 FILLER_72_805 ();
 sg13g2_fill_2 FILLER_72_812 ();
 sg13g2_fill_1 FILLER_72_814 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_48 ();
 sg13g2_fill_2 FILLER_73_75 ();
 sg13g2_fill_2 FILLER_73_103 ();
 sg13g2_fill_1 FILLER_73_122 ();
 sg13g2_fill_1 FILLER_73_127 ();
 sg13g2_fill_2 FILLER_73_141 ();
 sg13g2_decap_8 FILLER_73_149 ();
 sg13g2_decap_4 FILLER_73_156 ();
 sg13g2_fill_1 FILLER_73_195 ();
 sg13g2_fill_2 FILLER_73_218 ();
 sg13g2_fill_1 FILLER_73_220 ();
 sg13g2_fill_2 FILLER_73_230 ();
 sg13g2_fill_1 FILLER_73_270 ();
 sg13g2_decap_8 FILLER_73_297 ();
 sg13g2_decap_8 FILLER_73_304 ();
 sg13g2_decap_8 FILLER_73_311 ();
 sg13g2_decap_4 FILLER_73_351 ();
 sg13g2_fill_1 FILLER_73_355 ();
 sg13g2_fill_2 FILLER_73_361 ();
 sg13g2_fill_1 FILLER_73_363 ();
 sg13g2_decap_4 FILLER_73_373 ();
 sg13g2_fill_1 FILLER_73_377 ();
 sg13g2_fill_2 FILLER_73_410 ();
 sg13g2_fill_1 FILLER_73_438 ();
 sg13g2_fill_1 FILLER_73_470 ();
 sg13g2_fill_2 FILLER_73_485 ();
 sg13g2_decap_4 FILLER_73_524 ();
 sg13g2_fill_2 FILLER_73_528 ();
 sg13g2_fill_2 FILLER_73_550 ();
 sg13g2_fill_1 FILLER_73_552 ();
 sg13g2_decap_8 FILLER_73_568 ();
 sg13g2_decap_8 FILLER_73_575 ();
 sg13g2_decap_8 FILLER_73_582 ();
 sg13g2_decap_8 FILLER_73_589 ();
 sg13g2_decap_4 FILLER_73_596 ();
 sg13g2_fill_1 FILLER_73_608 ();
 sg13g2_decap_8 FILLER_73_617 ();
 sg13g2_decap_8 FILLER_73_624 ();
 sg13g2_decap_4 FILLER_73_666 ();
 sg13g2_fill_2 FILLER_73_683 ();
 sg13g2_decap_8 FILLER_73_729 ();
 sg13g2_fill_2 FILLER_73_736 ();
 sg13g2_fill_1 FILLER_73_738 ();
 sg13g2_decap_4 FILLER_73_747 ();
 sg13g2_fill_2 FILLER_73_788 ();
 sg13g2_fill_2 FILLER_73_816 ();
 sg13g2_fill_2 FILLER_74_79 ();
 sg13g2_fill_1 FILLER_74_85 ();
 sg13g2_fill_1 FILLER_74_99 ();
 sg13g2_decap_4 FILLER_74_161 ();
 sg13g2_fill_2 FILLER_74_165 ();
 sg13g2_fill_2 FILLER_74_177 ();
 sg13g2_fill_1 FILLER_74_179 ();
 sg13g2_fill_2 FILLER_74_188 ();
 sg13g2_fill_1 FILLER_74_190 ();
 sg13g2_fill_2 FILLER_74_213 ();
 sg13g2_fill_1 FILLER_74_215 ();
 sg13g2_fill_2 FILLER_74_221 ();
 sg13g2_fill_1 FILLER_74_223 ();
 sg13g2_decap_8 FILLER_74_228 ();
 sg13g2_fill_2 FILLER_74_235 ();
 sg13g2_fill_2 FILLER_74_241 ();
 sg13g2_decap_4 FILLER_74_247 ();
 sg13g2_fill_2 FILLER_74_263 ();
 sg13g2_decap_8 FILLER_74_270 ();
 sg13g2_decap_4 FILLER_74_277 ();
 sg13g2_decap_4 FILLER_74_285 ();
 sg13g2_fill_2 FILLER_74_289 ();
 sg13g2_decap_4 FILLER_74_305 ();
 sg13g2_fill_2 FILLER_74_309 ();
 sg13g2_decap_8 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_322 ();
 sg13g2_fill_2 FILLER_74_329 ();
 sg13g2_fill_2 FILLER_74_383 ();
 sg13g2_fill_1 FILLER_74_394 ();
 sg13g2_fill_1 FILLER_74_400 ();
 sg13g2_decap_4 FILLER_74_427 ();
 sg13g2_fill_1 FILLER_74_431 ();
 sg13g2_decap_8 FILLER_74_493 ();
 sg13g2_decap_4 FILLER_74_500 ();
 sg13g2_decap_4 FILLER_74_520 ();
 sg13g2_fill_1 FILLER_74_524 ();
 sg13g2_fill_1 FILLER_74_538 ();
 sg13g2_decap_4 FILLER_74_566 ();
 sg13g2_decap_8 FILLER_74_599 ();
 sg13g2_decap_8 FILLER_74_616 ();
 sg13g2_fill_2 FILLER_74_623 ();
 sg13g2_fill_1 FILLER_74_625 ();
 sg13g2_fill_2 FILLER_74_634 ();
 sg13g2_fill_2 FILLER_74_640 ();
 sg13g2_fill_1 FILLER_74_642 ();
 sg13g2_fill_2 FILLER_74_676 ();
 sg13g2_fill_1 FILLER_74_708 ();
 sg13g2_fill_2 FILLER_74_736 ();
 sg13g2_fill_1 FILLER_74_764 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_2 ();
 sg13g2_fill_2 FILLER_75_72 ();
 sg13g2_fill_2 FILLER_75_79 ();
 sg13g2_fill_1 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_115 ();
 sg13g2_decap_8 FILLER_75_121 ();
 sg13g2_fill_2 FILLER_75_128 ();
 sg13g2_decap_8 FILLER_75_134 ();
 sg13g2_decap_4 FILLER_75_141 ();
 sg13g2_fill_1 FILLER_75_145 ();
 sg13g2_fill_1 FILLER_75_150 ();
 sg13g2_fill_2 FILLER_75_177 ();
 sg13g2_fill_1 FILLER_75_187 ();
 sg13g2_fill_1 FILLER_75_196 ();
 sg13g2_fill_2 FILLER_75_223 ();
 sg13g2_fill_1 FILLER_75_233 ();
 sg13g2_fill_1 FILLER_75_249 ();
 sg13g2_fill_1 FILLER_75_309 ();
 sg13g2_decap_4 FILLER_75_324 ();
 sg13g2_fill_1 FILLER_75_328 ();
 sg13g2_decap_8 FILLER_75_333 ();
 sg13g2_decap_8 FILLER_75_340 ();
 sg13g2_decap_8 FILLER_75_351 ();
 sg13g2_decap_4 FILLER_75_358 ();
 sg13g2_fill_1 FILLER_75_362 ();
 sg13g2_decap_4 FILLER_75_398 ();
 sg13g2_fill_2 FILLER_75_402 ();
 sg13g2_fill_2 FILLER_75_410 ();
 sg13g2_fill_2 FILLER_75_416 ();
 sg13g2_decap_8 FILLER_75_422 ();
 sg13g2_decap_4 FILLER_75_429 ();
 sg13g2_fill_1 FILLER_75_438 ();
 sg13g2_decap_4 FILLER_75_448 ();
 sg13g2_fill_2 FILLER_75_452 ();
 sg13g2_fill_2 FILLER_75_466 ();
 sg13g2_decap_8 FILLER_75_508 ();
 sg13g2_fill_1 FILLER_75_515 ();
 sg13g2_fill_2 FILLER_75_526 ();
 sg13g2_fill_2 FILLER_75_543 ();
 sg13g2_fill_1 FILLER_75_545 ();
 sg13g2_decap_8 FILLER_75_565 ();
 sg13g2_fill_2 FILLER_75_580 ();
 sg13g2_fill_1 FILLER_75_582 ();
 sg13g2_fill_2 FILLER_75_609 ();
 sg13g2_fill_2 FILLER_75_627 ();
 sg13g2_fill_1 FILLER_75_629 ();
 sg13g2_fill_2 FILLER_75_634 ();
 sg13g2_fill_1 FILLER_75_644 ();
 sg13g2_fill_2 FILLER_75_649 ();
 sg13g2_decap_8 FILLER_75_668 ();
 sg13g2_decap_4 FILLER_75_675 ();
 sg13g2_fill_1 FILLER_75_679 ();
 sg13g2_fill_2 FILLER_75_687 ();
 sg13g2_decap_4 FILLER_75_694 ();
 sg13g2_fill_2 FILLER_75_703 ();
 sg13g2_decap_8 FILLER_75_724 ();
 sg13g2_decap_8 FILLER_75_731 ();
 sg13g2_fill_1 FILLER_75_770 ();
 sg13g2_fill_2 FILLER_75_789 ();
 sg13g2_fill_1 FILLER_75_821 ();
 sg13g2_fill_2 FILLER_75_826 ();
 sg13g2_fill_1 FILLER_75_828 ();
 sg13g2_fill_1 FILLER_76_31 ();
 sg13g2_fill_2 FILLER_76_59 ();
 sg13g2_fill_2 FILLER_76_65 ();
 sg13g2_fill_1 FILLER_76_67 ();
 sg13g2_fill_1 FILLER_76_82 ();
 sg13g2_fill_2 FILLER_76_97 ();
 sg13g2_decap_8 FILLER_76_153 ();
 sg13g2_fill_2 FILLER_76_186 ();
 sg13g2_fill_1 FILLER_76_188 ();
 sg13g2_decap_4 FILLER_76_202 ();
 sg13g2_fill_2 FILLER_76_206 ();
 sg13g2_fill_2 FILLER_76_212 ();
 sg13g2_fill_1 FILLER_76_214 ();
 sg13g2_decap_8 FILLER_76_219 ();
 sg13g2_decap_4 FILLER_76_226 ();
 sg13g2_decap_8 FILLER_76_249 ();
 sg13g2_fill_1 FILLER_76_278 ();
 sg13g2_fill_2 FILLER_76_284 ();
 sg13g2_fill_1 FILLER_76_295 ();
 sg13g2_fill_2 FILLER_76_305 ();
 sg13g2_fill_2 FILLER_76_327 ();
 sg13g2_fill_1 FILLER_76_329 ();
 sg13g2_fill_2 FILLER_76_335 ();
 sg13g2_fill_1 FILLER_76_337 ();
 sg13g2_decap_4 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_444 ();
 sg13g2_decap_8 FILLER_76_451 ();
 sg13g2_decap_8 FILLER_76_485 ();
 sg13g2_fill_1 FILLER_76_492 ();
 sg13g2_decap_8 FILLER_76_497 ();
 sg13g2_fill_2 FILLER_76_531 ();
 sg13g2_fill_1 FILLER_76_533 ();
 sg13g2_fill_1 FILLER_76_547 ();
 sg13g2_decap_4 FILLER_76_570 ();
 sg13g2_fill_2 FILLER_76_574 ();
 sg13g2_decap_8 FILLER_76_595 ();
 sg13g2_fill_2 FILLER_76_602 ();
 sg13g2_decap_4 FILLER_76_617 ();
 sg13g2_fill_2 FILLER_76_621 ();
 sg13g2_fill_2 FILLER_76_635 ();
 sg13g2_fill_1 FILLER_76_657 ();
 sg13g2_decap_4 FILLER_76_711 ();
 sg13g2_fill_1 FILLER_76_731 ();
 sg13g2_fill_1 FILLER_76_814 ();
 sg13g2_fill_2 FILLER_76_833 ();
 sg13g2_fill_1 FILLER_76_835 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_15 ();
 sg13g2_fill_1 FILLER_77_17 ();
 sg13g2_fill_1 FILLER_77_51 ();
 sg13g2_fill_1 FILLER_77_72 ();
 sg13g2_fill_1 FILLER_77_94 ();
 sg13g2_fill_1 FILLER_77_108 ();
 sg13g2_fill_2 FILLER_77_141 ();
 sg13g2_fill_1 FILLER_77_143 ();
 sg13g2_fill_2 FILLER_77_204 ();
 sg13g2_fill_1 FILLER_77_206 ();
 sg13g2_fill_2 FILLER_77_227 ();
 sg13g2_fill_1 FILLER_77_229 ();
 sg13g2_fill_1 FILLER_77_266 ();
 sg13g2_fill_2 FILLER_77_305 ();
 sg13g2_fill_2 FILLER_77_345 ();
 sg13g2_decap_4 FILLER_77_448 ();
 sg13g2_fill_1 FILLER_77_452 ();
 sg13g2_decap_8 FILLER_77_488 ();
 sg13g2_fill_2 FILLER_77_495 ();
 sg13g2_fill_1 FILLER_77_497 ();
 sg13g2_fill_2 FILLER_77_502 ();
 sg13g2_fill_1 FILLER_77_512 ();
 sg13g2_fill_1 FILLER_77_541 ();
 sg13g2_fill_1 FILLER_77_551 ();
 sg13g2_fill_2 FILLER_77_571 ();
 sg13g2_fill_1 FILLER_77_589 ();
 sg13g2_decap_8 FILLER_77_615 ();
 sg13g2_decap_8 FILLER_77_663 ();
 sg13g2_decap_4 FILLER_77_670 ();
 sg13g2_fill_1 FILLER_77_674 ();
 sg13g2_decap_4 FILLER_77_681 ();
 sg13g2_fill_2 FILLER_77_689 ();
 sg13g2_fill_1 FILLER_77_703 ();
 sg13g2_fill_2 FILLER_77_743 ();
 sg13g2_fill_2 FILLER_77_819 ();
 sg13g2_fill_1 FILLER_77_837 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_fill_2 FILLER_78_14 ();
 sg13g2_fill_1 FILLER_78_42 ();
 sg13g2_fill_2 FILLER_78_74 ();
 sg13g2_fill_1 FILLER_78_81 ();
 sg13g2_fill_2 FILLER_78_97 ();
 sg13g2_fill_2 FILLER_78_163 ();
 sg13g2_decap_4 FILLER_78_201 ();
 sg13g2_fill_2 FILLER_78_205 ();
 sg13g2_fill_1 FILLER_78_225 ();
 sg13g2_fill_2 FILLER_78_231 ();
 sg13g2_fill_1 FILLER_78_241 ();
 sg13g2_decap_4 FILLER_78_247 ();
 sg13g2_fill_2 FILLER_78_251 ();
 sg13g2_fill_2 FILLER_78_262 ();
 sg13g2_fill_1 FILLER_78_264 ();
 sg13g2_fill_2 FILLER_78_277 ();
 sg13g2_fill_1 FILLER_78_279 ();
 sg13g2_fill_2 FILLER_78_288 ();
 sg13g2_decap_8 FILLER_78_295 ();
 sg13g2_fill_2 FILLER_78_317 ();
 sg13g2_fill_1 FILLER_78_337 ();
 sg13g2_fill_1 FILLER_78_344 ();
 sg13g2_decap_4 FILLER_78_351 ();
 sg13g2_fill_1 FILLER_78_355 ();
 sg13g2_fill_1 FILLER_78_360 ();
 sg13g2_fill_1 FILLER_78_407 ();
 sg13g2_fill_2 FILLER_78_421 ();
 sg13g2_fill_2 FILLER_78_445 ();
 sg13g2_fill_2 FILLER_78_464 ();
 sg13g2_fill_1 FILLER_78_466 ();
 sg13g2_fill_2 FILLER_78_475 ();
 sg13g2_decap_4 FILLER_78_522 ();
 sg13g2_fill_1 FILLER_78_534 ();
 sg13g2_fill_1 FILLER_78_550 ();
 sg13g2_fill_2 FILLER_78_569 ();
 sg13g2_decap_8 FILLER_78_576 ();
 sg13g2_fill_1 FILLER_78_595 ();
 sg13g2_fill_2 FILLER_78_622 ();
 sg13g2_fill_1 FILLER_78_624 ();
 sg13g2_fill_2 FILLER_78_632 ();
 sg13g2_fill_2 FILLER_78_642 ();
 sg13g2_fill_1 FILLER_78_647 ();
 sg13g2_fill_1 FILLER_78_655 ();
 sg13g2_decap_4 FILLER_78_664 ();
 sg13g2_fill_2 FILLER_78_693 ();
 sg13g2_fill_1 FILLER_78_695 ();
 sg13g2_decap_8 FILLER_78_709 ();
 sg13g2_fill_2 FILLER_78_716 ();
 sg13g2_fill_1 FILLER_78_718 ();
 sg13g2_fill_2 FILLER_78_725 ();
 sg13g2_fill_1 FILLER_78_753 ();
 sg13g2_fill_1 FILLER_78_818 ();
 sg13g2_fill_2 FILLER_78_834 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_4 FILLER_79_21 ();
 sg13g2_fill_1 FILLER_79_61 ();
 sg13g2_fill_2 FILLER_79_88 ();
 sg13g2_fill_1 FILLER_79_189 ();
 sg13g2_fill_1 FILLER_79_223 ();
 sg13g2_fill_2 FILLER_79_247 ();
 sg13g2_fill_2 FILLER_79_259 ();
 sg13g2_fill_2 FILLER_79_284 ();
 sg13g2_fill_2 FILLER_79_322 ();
 sg13g2_fill_1 FILLER_79_324 ();
 sg13g2_fill_2 FILLER_79_339 ();
 sg13g2_fill_2 FILLER_79_349 ();
 sg13g2_fill_2 FILLER_79_377 ();
 sg13g2_fill_1 FILLER_79_379 ();
 sg13g2_fill_2 FILLER_79_500 ();
 sg13g2_fill_1 FILLER_79_502 ();
 sg13g2_fill_2 FILLER_79_532 ();
 sg13g2_fill_1 FILLER_79_534 ();
 sg13g2_fill_1 FILLER_79_550 ();
 sg13g2_fill_2 FILLER_79_609 ();
 sg13g2_fill_1 FILLER_79_611 ();
 sg13g2_fill_2 FILLER_79_628 ();
 sg13g2_fill_1 FILLER_79_630 ();
 sg13g2_fill_1 FILLER_79_768 ();
 sg13g2_fill_2 FILLER_79_777 ();
 sg13g2_fill_2 FILLER_79_803 ();
 sg13g2_decap_4 FILLER_79_857 ();
 sg13g2_fill_1 FILLER_79_861 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_51 ();
 sg13g2_fill_1 FILLER_80_64 ();
 sg13g2_fill_2 FILLER_80_133 ();
 sg13g2_fill_1 FILLER_80_135 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_fill_2 FILLER_80_233 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_decap_4 FILLER_80_249 ();
 sg13g2_fill_1 FILLER_80_253 ();
 sg13g2_fill_2 FILLER_80_270 ();
 sg13g2_decap_4 FILLER_80_277 ();
 sg13g2_fill_1 FILLER_80_281 ();
 sg13g2_fill_1 FILLER_80_286 ();
 sg13g2_decap_8 FILLER_80_297 ();
 sg13g2_fill_1 FILLER_80_304 ();
 sg13g2_decap_4 FILLER_80_323 ();
 sg13g2_fill_1 FILLER_80_327 ();
 sg13g2_decap_4 FILLER_80_344 ();
 sg13g2_decap_8 FILLER_80_352 ();
 sg13g2_fill_2 FILLER_80_359 ();
 sg13g2_fill_1 FILLER_80_361 ();
 sg13g2_decap_8 FILLER_80_366 ();
 sg13g2_fill_1 FILLER_80_373 ();
 sg13g2_fill_1 FILLER_80_388 ();
 sg13g2_fill_1 FILLER_80_398 ();
 sg13g2_fill_2 FILLER_80_408 ();
 sg13g2_fill_2 FILLER_80_431 ();
 sg13g2_fill_1 FILLER_80_433 ();
 sg13g2_fill_1 FILLER_80_447 ();
 sg13g2_fill_1 FILLER_80_504 ();
 sg13g2_fill_2 FILLER_80_513 ();
 sg13g2_decap_8 FILLER_80_524 ();
 sg13g2_decap_8 FILLER_80_531 ();
 sg13g2_fill_2 FILLER_80_538 ();
 sg13g2_fill_1 FILLER_80_540 ();
 sg13g2_fill_2 FILLER_80_546 ();
 sg13g2_decap_8 FILLER_80_558 ();
 sg13g2_decap_4 FILLER_80_565 ();
 sg13g2_fill_1 FILLER_80_569 ();
 sg13g2_decap_4 FILLER_80_578 ();
 sg13g2_fill_2 FILLER_80_582 ();
 sg13g2_decap_8 FILLER_80_601 ();
 sg13g2_decap_4 FILLER_80_613 ();
 sg13g2_decap_4 FILLER_80_630 ();
 sg13g2_decap_8 FILLER_80_638 ();
 sg13g2_decap_8 FILLER_80_645 ();
 sg13g2_decap_4 FILLER_80_652 ();
 sg13g2_fill_2 FILLER_80_656 ();
 sg13g2_decap_8 FILLER_80_663 ();
 sg13g2_fill_2 FILLER_80_670 ();
 sg13g2_fill_1 FILLER_80_672 ();
 sg13g2_decap_4 FILLER_80_690 ();
 sg13g2_fill_1 FILLER_80_738 ();
 sg13g2_fill_2 FILLER_80_773 ();
 sg13g2_decap_4 FILLER_80_814 ();
 sg13g2_decap_8 FILLER_80_853 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule

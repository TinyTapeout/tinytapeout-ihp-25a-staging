module tt_um_anas_7193 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \PWM_Generator._pwm_cnt_T_1[0] ;
 wire \PWM_Generator.fprev[0] ;
 wire \PWM_Generator.fprev[1] ;
 wire \PWM_Generator.fprev[2] ;
 wire \PWM_Generator.fprev[3] ;
 wire \PWM_Generator.fprev[4] ;
 wire \PWM_Generator.fprev[5] ;
 wire \PWM_Generator.pwm_cnt[0] ;
 wire \PWM_Generator.pwm_cnt[10] ;
 wire \PWM_Generator.pwm_cnt[11] ;
 wire \PWM_Generator.pwm_cnt[12] ;
 wire \PWM_Generator.pwm_cnt[13] ;
 wire \PWM_Generator.pwm_cnt[14] ;
 wire \PWM_Generator.pwm_cnt[15] ;
 wire \PWM_Generator.pwm_cnt[16] ;
 wire \PWM_Generator.pwm_cnt[17] ;
 wire \PWM_Generator.pwm_cnt[18] ;
 wire \PWM_Generator.pwm_cnt[19] ;
 wire \PWM_Generator.pwm_cnt[1] ;
 wire \PWM_Generator.pwm_cnt[20] ;
 wire \PWM_Generator.pwm_cnt[21] ;
 wire \PWM_Generator.pwm_cnt[22] ;
 wire \PWM_Generator.pwm_cnt[23] ;
 wire \PWM_Generator.pwm_cnt[24] ;
 wire \PWM_Generator.pwm_cnt[25] ;
 wire \PWM_Generator.pwm_cnt[26] ;
 wire \PWM_Generator.pwm_cnt[27] ;
 wire \PWM_Generator.pwm_cnt[28] ;
 wire \PWM_Generator.pwm_cnt[29] ;
 wire \PWM_Generator.pwm_cnt[2] ;
 wire \PWM_Generator.pwm_cnt[30] ;
 wire \PWM_Generator.pwm_cnt[31] ;
 wire \PWM_Generator.pwm_cnt[32] ;
 wire \PWM_Generator.pwm_cnt[33] ;
 wire \PWM_Generator.pwm_cnt[34] ;
 wire \PWM_Generator.pwm_cnt[35] ;
 wire \PWM_Generator.pwm_cnt[3] ;
 wire \PWM_Generator.pwm_cnt[4] ;
 wire \PWM_Generator.pwm_cnt[5] ;
 wire \PWM_Generator.pwm_cnt[6] ;
 wire \PWM_Generator.pwm_cnt[7] ;
 wire \PWM_Generator.pwm_cnt[8] ;
 wire \PWM_Generator.pwm_cnt[9] ;
 wire \PWM_Generator.pwm_out ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire clknet_0_clk;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;

 sg13g2_inv_1 _0599_ (.Y(_0063_),
    .A(net171));
 sg13g2_inv_1 _0600_ (.Y(_0064_),
    .A(net173));
 sg13g2_inv_1 _0601_ (.Y(_0065_),
    .A(net174));
 sg13g2_inv_2 _0602_ (.Y(_0066_),
    .A(net166));
 sg13g2_inv_1 _0603_ (.Y(_0067_),
    .A(_0000_));
 sg13g2_inv_1 _0604_ (.Y(_0068_),
    .A(\PWM_Generator.pwm_cnt[29] ));
 sg13g2_inv_1 _0605_ (.Y(_0069_),
    .A(\PWM_Generator.pwm_cnt[22] ));
 sg13g2_inv_1 _0606_ (.Y(_0070_),
    .A(\PWM_Generator.pwm_cnt[20] ));
 sg13g2_inv_1 _0607_ (.Y(_0071_),
    .A(\PWM_Generator.pwm_cnt[18] ));
 sg13g2_inv_2 _0608_ (.Y(_0072_),
    .A(\PWM_Generator.pwm_cnt[16] ));
 sg13g2_inv_1 _0609_ (.Y(_0073_),
    .A(_0007_));
 sg13g2_inv_2 _0610_ (.Y(_0074_),
    .A(\PWM_Generator.pwm_cnt[8] ));
 sg13g2_inv_1 _0611_ (.Y(_0075_),
    .A(net105));
 sg13g2_inv_1 _0612_ (.Y(_0076_),
    .A(\PWM_Generator.pwm_cnt[6] ));
 sg13g2_inv_1 _0613_ (.Y(_0077_),
    .A(net96));
 sg13g2_inv_1 _0614_ (.Y(_0078_),
    .A(net156));
 sg13g2_inv_1 _0615_ (.Y(_0079_),
    .A(net159));
 sg13g2_inv_1 _0616_ (.Y(_0080_),
    .A(net1));
 sg13g2_and2_1 _0617_ (.A(net8),
    .B(net12),
    .X(_0081_));
 sg13g2_mux2_1 _0618_ (.A0(net11),
    .A1(net10),
    .S(net8),
    .X(_0082_));
 sg13g2_mux2_1 _0619_ (.A0(_0081_),
    .A1(_0082_),
    .S(net9),
    .X(_0083_));
 sg13g2_nor2b_2 _0620_ (.A(net161),
    .B_N(_0083_),
    .Y(_0084_));
 sg13g2_nand3_1 _0621_ (.B(net158),
    .C(_0084_),
    .A(net148),
    .Y(_0085_));
 sg13g2_xor2_1 _0622_ (.B(_0085_),
    .A(\PWM_Generator.pwm_cnt[11] ),
    .X(_0086_));
 sg13g2_nand2b_1 _0623_ (.Y(_0087_),
    .B(net10),
    .A_N(net8));
 sg13g2_or2_1 _0624_ (.X(_0088_),
    .B(_0087_),
    .A(net163));
 sg13g2_nor3_1 _0625_ (.A(net163),
    .B(net162),
    .C(_0087_),
    .Y(_0089_));
 sg13g2_mux2_1 _0626_ (.A0(net12),
    .A1(net11),
    .S(net8),
    .X(_0090_));
 sg13g2_nand3_1 _0627_ (.B(net162),
    .C(_0090_),
    .A(net163),
    .Y(_0091_));
 sg13g2_nand2_1 _0628_ (.Y(_0092_),
    .A(net146),
    .B(_0091_));
 sg13g2_o21ai_1 _0629_ (.B1(_0092_),
    .Y(_0093_),
    .A1(net146),
    .A2(_0089_));
 sg13g2_or2_1 _0630_ (.X(_0094_),
    .B(_0093_),
    .A(net148));
 sg13g2_or2_1 _0631_ (.X(_0095_),
    .B(_0094_),
    .A(\PWM_Generator.pwm_cnt[24] ));
 sg13g2_nor2_1 _0632_ (.A(net163),
    .B(_0090_),
    .Y(_0096_));
 sg13g2_a21oi_2 _0633_ (.B1(_0096_),
    .Y(_0097_),
    .A2(_0087_),
    .A1(net163));
 sg13g2_nand3_1 _0634_ (.B(net158),
    .C(_0097_),
    .A(net161),
    .Y(_0098_));
 sg13g2_nand4_1 _0635_ (.B(net161),
    .C(net159),
    .A(net157),
    .Y(_0099_),
    .D(_0097_));
 sg13g2_and2_2 _0636_ (.A(net161),
    .B(_0083_),
    .X(_0100_));
 sg13g2_nand3_1 _0637_ (.B(net146),
    .C(_0100_),
    .A(net148),
    .Y(_0101_));
 sg13g2_xnor2_1 _0638_ (.Y(_0102_),
    .A(\PWM_Generator.pwm_cnt[7] ),
    .B(_0101_));
 sg13g2_nor2_1 _0639_ (.A(net156),
    .B(_0093_),
    .Y(_0103_));
 sg13g2_nand3_1 _0640_ (.B(net147),
    .C(_0100_),
    .A(net154),
    .Y(_0104_));
 sg13g2_nor2_1 _0641_ (.A(\PWM_Generator.pwm_cnt[23] ),
    .B(_0104_),
    .Y(_0105_));
 sg13g2_nand2_1 _0642_ (.Y(_0106_),
    .A(net158),
    .B(_0100_));
 sg13g2_nand3_1 _0643_ (.B(net158),
    .C(_0100_),
    .A(net154),
    .Y(_0107_));
 sg13g2_nor2b_1 _0644_ (.A(net161),
    .B_N(_0097_),
    .Y(_0108_));
 sg13g2_nand3_1 _0645_ (.B(net158),
    .C(_0108_),
    .A(net149),
    .Y(_0109_));
 sg13g2_nand2b_2 _0646_ (.Y(_0110_),
    .B(_0082_),
    .A_N(net163));
 sg13g2_or4_1 _0647_ (.A(net157),
    .B(net162),
    .C(net159),
    .D(_0110_),
    .X(_0111_));
 sg13g2_nand2_1 _0648_ (.Y(_0112_),
    .A(net9),
    .B(_0081_));
 sg13g2_mux2_2 _0649_ (.A0(_0112_),
    .A1(_0110_),
    .S(net162),
    .X(_0113_));
 sg13g2_nor3_1 _0650_ (.A(net148),
    .B(net158),
    .C(_0113_),
    .Y(_0114_));
 sg13g2_a21oi_1 _0651_ (.A1(net163),
    .A2(_0090_),
    .Y(_0115_),
    .B1(net162));
 sg13g2_a21oi_2 _0652_ (.B1(_0115_),
    .Y(_0116_),
    .A2(_0088_),
    .A1(net162));
 sg13g2_and3_1 _0653_ (.X(_0117_),
    .A(net149),
    .B(net147),
    .C(_0116_));
 sg13g2_xnor2_1 _0654_ (.Y(_0118_),
    .A(\PWM_Generator.pwm_cnt[4] ),
    .B(_0117_));
 sg13g2_nand3_1 _0655_ (.B(net147),
    .C(_0084_),
    .A(net157),
    .Y(_0119_));
 sg13g2_xor2_1 _0656_ (.B(_0119_),
    .A(\PWM_Generator.pwm_cnt[19] ),
    .X(_0120_));
 sg13g2_nand3_1 _0657_ (.B(net158),
    .C(_0116_),
    .A(net148),
    .Y(_0121_));
 sg13g2_nor2_1 _0658_ (.A(net146),
    .B(_0091_),
    .Y(_0122_));
 sg13g2_nand2_1 _0659_ (.Y(_0123_),
    .A(net154),
    .B(_0122_));
 sg13g2_and2_1 _0660_ (.A(net147),
    .B(_0108_),
    .X(_0124_));
 sg13g2_nor2_1 _0661_ (.A(\PWM_Generator.pwm_cnt[18] ),
    .B(\PWM_Generator.pwm_cnt[2] ),
    .Y(_0125_));
 sg13g2_a21oi_1 _0662_ (.A1(\PWM_Generator.pwm_cnt[18] ),
    .A2(net149),
    .Y(_0126_),
    .B1(_0125_));
 sg13g2_and2_1 _0663_ (.A(net146),
    .B(_0089_),
    .X(_0127_));
 sg13g2_and2_1 _0664_ (.A(net149),
    .B(_0127_),
    .X(_0128_));
 sg13g2_nor2_1 _0665_ (.A(\PWM_Generator._pwm_cnt_T_1[0] ),
    .B(_0128_),
    .Y(_0129_));
 sg13g2_and4_1 _0666_ (.A(net163),
    .B(net8),
    .C(net162),
    .D(net12),
    .X(_0130_));
 sg13g2_and2_1 _0667_ (.A(net160),
    .B(_0130_),
    .X(_0131_));
 sg13g2_nand3_1 _0668_ (.B(net159),
    .C(_0130_),
    .A(net157),
    .Y(_0132_));
 sg13g2_or2_1 _0669_ (.X(_0133_),
    .B(\PWM_Generator.pwm_cnt[34] ),
    .A(\PWM_Generator.pwm_cnt[35] ));
 sg13g2_nand3_1 _0670_ (.B(net146),
    .C(_0084_),
    .A(net148),
    .Y(_0134_));
 sg13g2_xnor2_1 _0671_ (.Y(_0135_),
    .A(\PWM_Generator.pwm_cnt[3] ),
    .B(_0134_));
 sg13g2_nand3_1 _0672_ (.B(net160),
    .C(_0108_),
    .A(net157),
    .Y(_0136_));
 sg13g2_xor2_1 _0673_ (.B(_0136_),
    .A(\PWM_Generator.pwm_cnt[26] ),
    .X(_0137_));
 sg13g2_nor4_1 _0674_ (.A(net149),
    .B(net161),
    .C(net159),
    .D(_0110_),
    .Y(_0138_));
 sg13g2_a21oi_1 _0675_ (.A1(net149),
    .A2(_0131_),
    .Y(_0139_),
    .B1(_0138_));
 sg13g2_nor3_1 _0676_ (.A(net156),
    .B(net159),
    .C(_0113_),
    .Y(_0140_));
 sg13g2_nand3_1 _0677_ (.B(net158),
    .C(_0084_),
    .A(net155),
    .Y(_0141_));
 sg13g2_nor2_1 _0678_ (.A(\PWM_Generator.pwm_cnt[27] ),
    .B(_0141_),
    .Y(_0142_));
 sg13g2_nor2_1 _0679_ (.A(net147),
    .B(_0113_),
    .Y(_0143_));
 sg13g2_a21oi_1 _0680_ (.A1(net155),
    .A2(_0143_),
    .Y(_0144_),
    .B1(_0068_));
 sg13g2_nand3_1 _0681_ (.B(net147),
    .C(_0116_),
    .A(net154),
    .Y(_0145_));
 sg13g2_nand2_1 _0682_ (.Y(_0146_),
    .A(\PWM_Generator.pwm_cnt[20] ),
    .B(_0145_));
 sg13g2_mux2_1 _0683_ (.A0(_0122_),
    .A1(_0127_),
    .S(net154),
    .X(_0147_));
 sg13g2_nand4_1 _0684_ (.B(net161),
    .C(net146),
    .A(net154),
    .Y(_0148_),
    .D(_0097_));
 sg13g2_nor2_1 _0685_ (.A(\PWM_Generator.pwm_cnt[22] ),
    .B(_0148_),
    .Y(_0149_));
 sg13g2_o21ai_1 _0686_ (.B1(\PWM_Generator.pwm_cnt[8] ),
    .Y(_0150_),
    .A1(net155),
    .A2(_0093_));
 sg13g2_nor3_1 _0687_ (.A(\PWM_Generator.pwm_cnt[14] ),
    .B(net154),
    .C(_0098_),
    .Y(_0151_));
 sg13g2_nand3_1 _0688_ (.B(net160),
    .C(_0116_),
    .A(net157),
    .Y(_0152_));
 sg13g2_o21ai_1 _0689_ (.B1(net159),
    .Y(_0153_),
    .A1(net162),
    .A2(_0110_));
 sg13g2_o21ai_1 _0690_ (.B1(_0153_),
    .Y(_0154_),
    .A1(net159),
    .A2(_0130_));
 sg13g2_nand2b_1 _0691_ (.Y(_0155_),
    .B(net148),
    .A_N(_0154_));
 sg13g2_nor3_1 _0692_ (.A(\PWM_Generator.pwm_cnt[15] ),
    .B(net155),
    .C(_0106_),
    .Y(_0156_));
 sg13g2_and4_1 _0693_ (.A(net148),
    .B(net161),
    .C(net146),
    .D(_0097_),
    .X(_0157_));
 sg13g2_o21ai_1 _0694_ (.B1(\PWM_Generator.pwm_cnt[15] ),
    .Y(_0158_),
    .A1(net155),
    .A2(_0106_));
 sg13g2_nor3_1 _0695_ (.A(net155),
    .B(net147),
    .C(_0113_),
    .Y(_0159_));
 sg13g2_nor2b_1 _0696_ (.A(_0159_),
    .B_N(\PWM_Generator.pwm_cnt[13] ),
    .Y(_0160_));
 sg13g2_nor2b_1 _0697_ (.A(\PWM_Generator.pwm_cnt[13] ),
    .B_N(_0159_),
    .Y(_0161_));
 sg13g2_nor2_1 _0698_ (.A(net149),
    .B(_0154_),
    .Y(_0162_));
 sg13g2_nor2_1 _0699_ (.A(\PWM_Generator.pwm_cnt[20] ),
    .B(_0145_),
    .Y(_0163_));
 sg13g2_nor2_1 _0700_ (.A(\PWM_Generator.pwm_cnt[9] ),
    .B(_0155_),
    .Y(_0164_));
 sg13g2_nand3_1 _0701_ (.B(net155),
    .C(_0143_),
    .A(_0068_),
    .Y(_0165_));
 sg13g2_xor2_1 _0702_ (.B(_0107_),
    .A(\PWM_Generator.pwm_cnt[31] ),
    .X(_0166_));
 sg13g2_xor2_1 _0703_ (.B(_0140_),
    .A(\PWM_Generator.pwm_cnt[5] ),
    .X(_0167_));
 sg13g2_xnor2_1 _0704_ (.Y(_0168_),
    .A(\PWM_Generator.pwm_cnt[6] ),
    .B(_0157_));
 sg13g2_a21oi_1 _0705_ (.A1(\PWM_Generator.pwm_cnt[2] ),
    .A2(net157),
    .Y(_0169_),
    .B1(_0129_));
 sg13g2_xnor2_1 _0706_ (.Y(_0170_),
    .A(\PWM_Generator.pwm_cnt[21] ),
    .B(_0114_));
 sg13g2_o21ai_1 _0707_ (.B1(_0146_),
    .Y(_0171_),
    .A1(\PWM_Generator.pwm_cnt[17] ),
    .A2(_0139_));
 sg13g2_a22oi_1 _0708_ (.Y(_0172_),
    .B1(_0147_),
    .B2(_0072_),
    .A2(_0104_),
    .A1(\PWM_Generator.pwm_cnt[23] ));
 sg13g2_o21ai_1 _0709_ (.B1(_0172_),
    .Y(_0173_),
    .A1(_0072_),
    .A2(_0147_));
 sg13g2_nor4_1 _0710_ (.A(_0144_),
    .B(_0151_),
    .C(_0171_),
    .D(_0173_),
    .Y(_0174_));
 sg13g2_a21oi_1 _0711_ (.A1(\PWM_Generator.pwm_cnt[12] ),
    .A2(_0121_),
    .Y(_0175_),
    .B1(_0160_));
 sg13g2_a21oi_1 _0712_ (.A1(\PWM_Generator.pwm_cnt[22] ),
    .A2(_0148_),
    .Y(_0176_),
    .B1(_0142_));
 sg13g2_nor2_1 _0713_ (.A(\PWM_Generator.pwm_cnt[12] ),
    .B(_0121_),
    .Y(_0177_));
 sg13g2_xnor2_1 _0714_ (.Y(_0178_),
    .A(\PWM_Generator.pwm_cnt[33] ),
    .B(_0132_));
 sg13g2_a22oi_1 _0715_ (.Y(_0179_),
    .B1(_0141_),
    .B2(\PWM_Generator.pwm_cnt[27] ),
    .A2(_0103_),
    .A1(_0074_));
 sg13g2_xor2_1 _0716_ (.B(_0123_),
    .A(\PWM_Generator.pwm_cnt[32] ),
    .X(_0180_));
 sg13g2_nor2_1 _0717_ (.A(_0105_),
    .B(_0163_),
    .Y(_0181_));
 sg13g2_nand4_1 _0718_ (.B(_0179_),
    .C(_0180_),
    .A(_0158_),
    .Y(_0182_),
    .D(_0181_));
 sg13g2_nor3_1 _0719_ (.A(_0161_),
    .B(_0177_),
    .C(_0182_),
    .Y(_0183_));
 sg13g2_a21oi_1 _0720_ (.A1(\PWM_Generator.pwm_cnt[9] ),
    .A2(_0155_),
    .Y(_0184_),
    .B1(_0156_));
 sg13g2_nand4_1 _0721_ (.B(_0165_),
    .C(_0176_),
    .A(_0150_),
    .Y(_0185_),
    .D(_0184_));
 sg13g2_nor3_1 _0722_ (.A(_0149_),
    .B(_0164_),
    .C(_0185_),
    .Y(_0186_));
 sg13g2_a221oi_1 _0723_ (.B2(\PWM_Generator.pwm_cnt[17] ),
    .C1(_0167_),
    .B1(_0139_),
    .A1(\PWM_Generator.pwm_cnt[24] ),
    .Y(_0187_),
    .A2(_0094_));
 sg13g2_and4_1 _0724_ (.A(_0166_),
    .B(_0174_),
    .C(_0175_),
    .D(_0187_),
    .X(_0188_));
 sg13g2_xnor2_1 _0725_ (.Y(_0189_),
    .A(\PWM_Generator.pwm_cnt[25] ),
    .B(_0162_));
 sg13g2_mux2_1 _0726_ (.A0(_0125_),
    .A1(_0126_),
    .S(_0124_),
    .X(_0190_));
 sg13g2_a21oi_1 _0727_ (.A1(\PWM_Generator._pwm_cnt_T_1[0] ),
    .A2(_0128_),
    .Y(_0191_),
    .B1(_0133_));
 sg13g2_nand4_1 _0728_ (.B(_0189_),
    .C(_0190_),
    .A(_0169_),
    .Y(_0192_),
    .D(_0191_));
 sg13g2_o21ai_1 _0729_ (.B1(\PWM_Generator.pwm_cnt[14] ),
    .Y(_0193_),
    .A1(net154),
    .A2(_0098_));
 sg13g2_xnor2_1 _0730_ (.Y(_0194_),
    .A(\PWM_Generator.pwm_cnt[30] ),
    .B(_0099_));
 sg13g2_a21oi_1 _0731_ (.A1(\PWM_Generator.pwm_cnt[1] ),
    .A2(_0111_),
    .Y(_0195_),
    .B1(_0178_));
 sg13g2_o21ai_1 _0732_ (.B1(_0195_),
    .Y(_0196_),
    .A1(\PWM_Generator.pwm_cnt[1] ),
    .A2(_0111_));
 sg13g2_nor4_1 _0733_ (.A(_0102_),
    .B(_0135_),
    .C(_0194_),
    .D(_0196_),
    .Y(_0197_));
 sg13g2_nand4_1 _0734_ (.B(_0095_),
    .C(_0193_),
    .A(_0086_),
    .Y(_0198_),
    .D(_0197_));
 sg13g2_xor2_1 _0735_ (.B(_0109_),
    .A(\PWM_Generator.pwm_cnt[10] ),
    .X(_0199_));
 sg13g2_xor2_1 _0736_ (.B(_0152_),
    .A(\PWM_Generator.pwm_cnt[28] ),
    .X(_0200_));
 sg13g2_nand4_1 _0737_ (.B(_0170_),
    .C(_0199_),
    .A(_0120_),
    .Y(_0201_),
    .D(_0200_));
 sg13g2_nand3_1 _0738_ (.B(_0137_),
    .C(_0168_),
    .A(_0118_),
    .Y(_0202_));
 sg13g2_nor4_1 _0739_ (.A(_0192_),
    .B(_0198_),
    .C(_0201_),
    .D(_0202_),
    .Y(_0203_));
 sg13g2_nand4_1 _0740_ (.B(_0186_),
    .C(_0188_),
    .A(_0183_),
    .Y(_0204_),
    .D(_0203_));
 sg13g2_nand2_1 _0741_ (.Y(_0205_),
    .A(net1),
    .B(net142));
 sg13g2_nor2_1 _0742_ (.A(_0077_),
    .B(net138),
    .Y(_0014_));
 sg13g2_xnor2_1 _0743_ (.Y(_0206_),
    .A(\PWM_Generator.pwm_cnt[1] ),
    .B(net112));
 sg13g2_nor2_1 _0744_ (.A(net138),
    .B(net113),
    .Y(_0015_));
 sg13g2_and3_1 _0745_ (.X(_0207_),
    .A(net123),
    .B(\PWM_Generator.pwm_cnt[1] ),
    .C(net112));
 sg13g2_a21oi_1 _0746_ (.A1(\PWM_Generator.pwm_cnt[1] ),
    .A2(net112),
    .Y(_0208_),
    .B1(net123));
 sg13g2_nor3_1 _0747_ (.A(net137),
    .B(_0207_),
    .C(net124),
    .Y(_0016_));
 sg13g2_and4_2 _0748_ (.A(net108),
    .B(\PWM_Generator.pwm_cnt[2] ),
    .C(\PWM_Generator.pwm_cnt[1] ),
    .D(net112),
    .X(_0209_));
 sg13g2_nor2_1 _0749_ (.A(net108),
    .B(_0207_),
    .Y(_0210_));
 sg13g2_nor3_1 _0750_ (.A(net137),
    .B(_0209_),
    .C(net109),
    .Y(_0017_));
 sg13g2_and2_1 _0751_ (.A(net130),
    .B(_0209_),
    .X(_0211_));
 sg13g2_nor2_1 _0752_ (.A(net130),
    .B(_0209_),
    .Y(_0212_));
 sg13g2_nor3_1 _0753_ (.A(net137),
    .B(_0211_),
    .C(_0212_),
    .Y(_0018_));
 sg13g2_xnor2_1 _0754_ (.Y(_0213_),
    .A(net126),
    .B(_0211_));
 sg13g2_nor2_1 _0755_ (.A(net137),
    .B(net127),
    .Y(_0019_));
 sg13g2_nand4_1 _0756_ (.B(\PWM_Generator.pwm_cnt[5] ),
    .C(\PWM_Generator.pwm_cnt[4] ),
    .A(\PWM_Generator.pwm_cnt[6] ),
    .Y(_0214_),
    .D(_0209_));
 sg13g2_inv_1 _0757_ (.Y(_0215_),
    .A(_0214_));
 sg13g2_a21oi_1 _0758_ (.A1(\PWM_Generator.pwm_cnt[5] ),
    .A2(_0211_),
    .Y(_0216_),
    .B1(net103));
 sg13g2_nor3_1 _0759_ (.A(net135),
    .B(_0215_),
    .C(net104),
    .Y(_0020_));
 sg13g2_nor2_1 _0760_ (.A(net105),
    .B(_0215_),
    .Y(_0217_));
 sg13g2_nor2_1 _0761_ (.A(_0075_),
    .B(_0214_),
    .Y(_0218_));
 sg13g2_nor3_1 _0762_ (.A(net135),
    .B(_0217_),
    .C(_0218_),
    .Y(_0021_));
 sg13g2_nor3_2 _0763_ (.A(_0074_),
    .B(_0075_),
    .C(_0214_),
    .Y(_0219_));
 sg13g2_nor2_1 _0764_ (.A(net116),
    .B(_0218_),
    .Y(_0220_));
 sg13g2_nor3_1 _0765_ (.A(net138),
    .B(_0219_),
    .C(_0220_),
    .Y(_0022_));
 sg13g2_xnor2_1 _0766_ (.Y(_0221_),
    .A(net114),
    .B(_0219_));
 sg13g2_nor2_1 _0767_ (.A(net135),
    .B(_0221_),
    .Y(_0023_));
 sg13g2_nand2_1 _0768_ (.Y(_0222_),
    .A(\PWM_Generator.pwm_cnt[10] ),
    .B(net114));
 sg13g2_nor4_2 _0769_ (.A(_0074_),
    .B(_0075_),
    .C(_0214_),
    .Y(_0223_),
    .D(_0222_));
 sg13g2_a21oi_1 _0770_ (.A1(net114),
    .A2(_0219_),
    .Y(_0224_),
    .B1(\PWM_Generator.pwm_cnt[10] ));
 sg13g2_nor3_1 _0771_ (.A(net135),
    .B(_0223_),
    .C(net115),
    .Y(_0024_));
 sg13g2_and2_1 _0772_ (.A(net110),
    .B(_0223_),
    .X(_0225_));
 sg13g2_nor2_1 _0773_ (.A(net110),
    .B(_0223_),
    .Y(_0226_));
 sg13g2_nor3_1 _0774_ (.A(net135),
    .B(_0225_),
    .C(net111),
    .Y(_0025_));
 sg13g2_xnor2_1 _0775_ (.Y(_0227_),
    .A(net178),
    .B(_0225_));
 sg13g2_nor2_1 _0776_ (.A(net133),
    .B(_0227_),
    .Y(_0026_));
 sg13g2_and4_1 _0777_ (.A(net83),
    .B(\PWM_Generator.pwm_cnt[12] ),
    .C(net110),
    .D(_0223_),
    .X(_0228_));
 sg13g2_a21oi_1 _0778_ (.A1(\PWM_Generator.pwm_cnt[12] ),
    .A2(_0225_),
    .Y(_0229_),
    .B1(net83));
 sg13g2_nor3_1 _0779_ (.A(net133),
    .B(_0228_),
    .C(net84),
    .Y(_0027_));
 sg13g2_and2_1 _0780_ (.A(net132),
    .B(_0228_),
    .X(_0230_));
 sg13g2_nor2_1 _0781_ (.A(net132),
    .B(_0228_),
    .Y(_0231_));
 sg13g2_nor3_1 _0782_ (.A(net133),
    .B(_0230_),
    .C(_0231_),
    .Y(_0028_));
 sg13g2_and2_1 _0783_ (.A(net106),
    .B(_0230_),
    .X(_0232_));
 sg13g2_nor2_1 _0784_ (.A(net106),
    .B(_0230_),
    .Y(_0233_));
 sg13g2_nor3_1 _0785_ (.A(net133),
    .B(_0232_),
    .C(net107),
    .Y(_0029_));
 sg13g2_xnor2_1 _0786_ (.Y(_0234_),
    .A(net119),
    .B(_0232_));
 sg13g2_nor2_1 _0787_ (.A(net133),
    .B(_0234_),
    .Y(_0030_));
 sg13g2_a21oi_1 _0788_ (.A1(net119),
    .A2(_0232_),
    .Y(_0235_),
    .B1(net120));
 sg13g2_and2_1 _0789_ (.A(\PWM_Generator.pwm_cnt[17] ),
    .B(\PWM_Generator.pwm_cnt[16] ),
    .X(_0236_));
 sg13g2_and4_2 _0790_ (.A(net106),
    .B(\PWM_Generator.pwm_cnt[14] ),
    .C(_0228_),
    .D(_0236_),
    .X(_0237_));
 sg13g2_nor3_1 _0791_ (.A(net133),
    .B(_0235_),
    .C(_0237_),
    .Y(_0031_));
 sg13g2_nor2_1 _0792_ (.A(net184),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_and2_1 _0793_ (.A(net184),
    .B(_0237_),
    .X(_0239_));
 sg13g2_nor3_1 _0794_ (.A(net137),
    .B(_0238_),
    .C(_0239_),
    .Y(_0032_));
 sg13g2_nor2_1 _0795_ (.A(net125),
    .B(_0239_),
    .Y(_0240_));
 sg13g2_and2_1 _0796_ (.A(net125),
    .B(_0239_),
    .X(_0241_));
 sg13g2_nor3_1 _0797_ (.A(net137),
    .B(_0240_),
    .C(_0241_),
    .Y(_0033_));
 sg13g2_nor2_1 _0798_ (.A(net175),
    .B(_0241_),
    .Y(_0242_));
 sg13g2_and4_1 _0799_ (.A(\PWM_Generator.pwm_cnt[20] ),
    .B(\PWM_Generator.pwm_cnt[19] ),
    .C(\PWM_Generator.pwm_cnt[18] ),
    .D(_0237_),
    .X(_0243_));
 sg13g2_nor3_1 _0800_ (.A(net136),
    .B(_0242_),
    .C(_0243_),
    .Y(_0034_));
 sg13g2_nor2_1 _0801_ (.A(net128),
    .B(_0243_),
    .Y(_0244_));
 sg13g2_and2_1 _0802_ (.A(net128),
    .B(_0243_),
    .X(_0245_));
 sg13g2_nor3_1 _0803_ (.A(net136),
    .B(net129),
    .C(_0245_),
    .Y(_0035_));
 sg13g2_nor2_1 _0804_ (.A(net186),
    .B(_0245_),
    .Y(_0246_));
 sg13g2_and2_1 _0805_ (.A(net186),
    .B(_0245_),
    .X(_0247_));
 sg13g2_nor3_1 _0806_ (.A(net136),
    .B(_0246_),
    .C(_0247_),
    .Y(_0036_));
 sg13g2_nor2_1 _0807_ (.A(net117),
    .B(_0247_),
    .Y(_0248_));
 sg13g2_and4_2 _0808_ (.A(net117),
    .B(\PWM_Generator.pwm_cnt[22] ),
    .C(\PWM_Generator.pwm_cnt[21] ),
    .D(_0243_),
    .X(_0249_));
 sg13g2_nor3_1 _0809_ (.A(net137),
    .B(net118),
    .C(_0249_),
    .Y(_0037_));
 sg13g2_nor2_1 _0810_ (.A(net182),
    .B(_0249_),
    .Y(_0250_));
 sg13g2_and2_1 _0811_ (.A(net182),
    .B(_0249_),
    .X(_0251_));
 sg13g2_nor3_1 _0812_ (.A(net136),
    .B(net183),
    .C(_0251_),
    .Y(_0038_));
 sg13g2_nor2_1 _0813_ (.A(net121),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_and2_1 _0814_ (.A(\PWM_Generator.pwm_cnt[25] ),
    .B(\PWM_Generator.pwm_cnt[24] ),
    .X(_0253_));
 sg13g2_and2_1 _0815_ (.A(_0249_),
    .B(_0253_),
    .X(_0254_));
 sg13g2_nor3_1 _0816_ (.A(net133),
    .B(net122),
    .C(_0254_),
    .Y(_0039_));
 sg13g2_xnor2_1 _0817_ (.Y(_0255_),
    .A(net188),
    .B(_0254_));
 sg13g2_nor2_1 _0818_ (.A(net134),
    .B(_0255_),
    .Y(_0040_));
 sg13g2_a21oi_1 _0819_ (.A1(\PWM_Generator.pwm_cnt[26] ),
    .A2(_0254_),
    .Y(_0256_),
    .B1(net101));
 sg13g2_and4_2 _0820_ (.A(net101),
    .B(\PWM_Generator.pwm_cnt[26] ),
    .C(_0249_),
    .D(_0253_),
    .X(_0257_));
 sg13g2_nor3_1 _0821_ (.A(net134),
    .B(net102),
    .C(_0257_),
    .Y(_0041_));
 sg13g2_xnor2_1 _0822_ (.Y(_0258_),
    .A(net179),
    .B(_0257_));
 sg13g2_nor2_1 _0823_ (.A(net133),
    .B(_0258_),
    .Y(_0042_));
 sg13g2_a21oi_1 _0824_ (.A1(\PWM_Generator.pwm_cnt[28] ),
    .A2(_0257_),
    .Y(_0259_),
    .B1(net78));
 sg13g2_and2_1 _0825_ (.A(\PWM_Generator.pwm_cnt[29] ),
    .B(\PWM_Generator.pwm_cnt[28] ),
    .X(_0260_));
 sg13g2_and2_1 _0826_ (.A(_0257_),
    .B(_0260_),
    .X(_0261_));
 sg13g2_nor3_1 _0827_ (.A(net134),
    .B(net79),
    .C(_0261_),
    .Y(_0043_));
 sg13g2_xnor2_1 _0828_ (.Y(_0262_),
    .A(net189),
    .B(_0261_));
 sg13g2_nor2_1 _0829_ (.A(net134),
    .B(_0262_),
    .Y(_0044_));
 sg13g2_a21oi_1 _0830_ (.A1(\PWM_Generator.pwm_cnt[30] ),
    .A2(_0261_),
    .Y(_0263_),
    .B1(net90));
 sg13g2_and4_1 _0831_ (.A(net90),
    .B(\PWM_Generator.pwm_cnt[30] ),
    .C(_0257_),
    .D(_0260_),
    .X(_0264_));
 sg13g2_nor3_1 _0832_ (.A(net134),
    .B(net91),
    .C(_0264_),
    .Y(_0045_));
 sg13g2_nor2_1 _0833_ (.A(net190),
    .B(_0264_),
    .Y(_0265_));
 sg13g2_and2_1 _0834_ (.A(\PWM_Generator.pwm_cnt[32] ),
    .B(_0264_),
    .X(_0266_));
 sg13g2_nor3_1 _0835_ (.A(net136),
    .B(_0265_),
    .C(_0266_),
    .Y(_0046_));
 sg13g2_nor2_1 _0836_ (.A(net187),
    .B(_0266_),
    .Y(_0267_));
 sg13g2_a21oi_1 _0837_ (.A1(net187),
    .A2(_0266_),
    .Y(_0268_),
    .B1(net136));
 sg13g2_nor2b_1 _0838_ (.A(_0267_),
    .B_N(_0268_),
    .Y(_0047_));
 sg13g2_a21oi_1 _0839_ (.A1(\PWM_Generator.pwm_cnt[33] ),
    .A2(_0266_),
    .Y(_0269_),
    .B1(net81));
 sg13g2_and4_1 _0840_ (.A(net81),
    .B(\PWM_Generator.pwm_cnt[33] ),
    .C(\PWM_Generator.pwm_cnt[32] ),
    .D(_0264_),
    .X(_0270_));
 sg13g2_nor3_1 _0841_ (.A(net136),
    .B(net82),
    .C(_0270_),
    .Y(_0048_));
 sg13g2_nor2_1 _0842_ (.A(net87),
    .B(_0270_),
    .Y(_0271_));
 sg13g2_a21oi_1 _0843_ (.A1(net87),
    .A2(_0270_),
    .Y(_0272_),
    .B1(net136));
 sg13g2_nor2b_1 _0844_ (.A(_0271_),
    .B_N(_0272_),
    .Y(_0049_));
 sg13g2_and2_1 _0845_ (.A(net7),
    .B(net2),
    .X(_0273_));
 sg13g2_and4_1 _0846_ (.A(net4),
    .B(net7),
    .C(net2),
    .D(net3),
    .X(_0274_));
 sg13g2_and2_1 _0847_ (.A(net171),
    .B(_0274_),
    .X(_0275_));
 sg13g2_nand2_1 _0848_ (.Y(_0276_),
    .A(net168),
    .B(_0275_));
 sg13g2_or2_1 _0849_ (.X(_0277_),
    .B(_0276_),
    .A(\PWM_Generator.pwm_cnt[33] ));
 sg13g2_mux2_1 _0850_ (.A0(net7),
    .A1(net6),
    .S(net2),
    .X(_0278_));
 sg13g2_and4_1 _0851_ (.A(net170),
    .B(net172),
    .C(net174),
    .D(_0278_),
    .X(_0279_));
 sg13g2_nand2_1 _0852_ (.Y(_0280_),
    .A(net168),
    .B(_0279_));
 sg13g2_o21ai_1 _0853_ (.B1(_0277_),
    .Y(_0281_),
    .A1(\PWM_Generator.pwm_cnt[32] ),
    .A2(_0280_));
 sg13g2_nand2_1 _0854_ (.Y(_0282_),
    .A(\PWM_Generator.pwm_cnt[32] ),
    .B(_0280_));
 sg13g2_a21oi_1 _0855_ (.A1(\PWM_Generator.pwm_cnt[33] ),
    .A2(_0276_),
    .Y(_0283_),
    .B1(_0133_));
 sg13g2_nand3b_1 _0856_ (.B(_0282_),
    .C(_0283_),
    .Y(_0284_),
    .A_N(_0281_));
 sg13g2_mux2_2 _0857_ (.A0(net6),
    .A1(net5),
    .S(net2),
    .X(_0285_));
 sg13g2_and2_1 _0858_ (.A(_0065_),
    .B(_0285_),
    .X(_0286_));
 sg13g2_a21oi_2 _0859_ (.B1(net152),
    .Y(_0287_),
    .A2(_0285_),
    .A1(_0065_));
 sg13g2_a21oi_2 _0860_ (.B1(net172),
    .Y(_0288_),
    .A2(_0273_),
    .A1(net174));
 sg13g2_nor3_2 _0861_ (.A(net153),
    .B(_0287_),
    .C(_0288_),
    .Y(_0289_));
 sg13g2_nand3_1 _0862_ (.B(_0001_),
    .C(_0289_),
    .A(net164),
    .Y(_0290_));
 sg13g2_inv_1 _0863_ (.Y(_0291_),
    .A(_0290_));
 sg13g2_nor2b_1 _0864_ (.A(net2),
    .B_N(net5),
    .Y(_0292_));
 sg13g2_nand2b_1 _0865_ (.Y(_0293_),
    .B(net5),
    .A_N(net2));
 sg13g2_o21ai_1 _0866_ (.B1(net172),
    .Y(_0294_),
    .A1(net174),
    .A2(_0293_));
 sg13g2_a21o_1 _0867_ (.A2(_0278_),
    .A1(net174),
    .B1(net172),
    .X(_0295_));
 sg13g2_nand3_1 _0868_ (.B(_0294_),
    .C(_0295_),
    .A(net170),
    .Y(_0296_));
 sg13g2_nor2_1 _0869_ (.A(net150),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_a21o_1 _0870_ (.A2(net2),
    .A1(net7),
    .B1(net3),
    .X(_0298_));
 sg13g2_mux2_1 _0871_ (.A0(_0273_),
    .A1(_0285_),
    .S(net3),
    .X(_0299_));
 sg13g2_o21ai_1 _0872_ (.B1(_0298_),
    .Y(_0300_),
    .A1(_0065_),
    .A2(_0285_));
 sg13g2_nor2_1 _0873_ (.A(net173),
    .B(_0300_),
    .Y(_0301_));
 sg13g2_nand3_1 _0874_ (.B(net164),
    .C(_0301_),
    .A(net169),
    .Y(_0302_));
 sg13g2_nand2b_1 _0875_ (.Y(_0303_),
    .B(_0302_),
    .A_N(_0002_));
 sg13g2_nand4_1 _0876_ (.B(net173),
    .C(net166),
    .A(net169),
    .Y(_0304_),
    .D(_0299_));
 sg13g2_inv_1 _0877_ (.Y(_0305_),
    .A(_0304_));
 sg13g2_mux2_2 _0878_ (.A0(_0278_),
    .A1(_0292_),
    .S(net174),
    .X(_0306_));
 sg13g2_nand3_1 _0879_ (.B(net173),
    .C(_0306_),
    .A(net169),
    .Y(_0307_));
 sg13g2_or2_1 _0880_ (.X(_0308_),
    .B(_0307_),
    .A(net150));
 sg13g2_nor2_1 _0881_ (.A(\PWM_Generator.pwm_cnt[30] ),
    .B(_0308_),
    .Y(_0309_));
 sg13g2_a21oi_1 _0882_ (.A1(_0000_),
    .A2(_0305_),
    .Y(_0310_),
    .B1(_0309_));
 sg13g2_nand2_1 _0883_ (.Y(_0311_),
    .A(\PWM_Generator.pwm_cnt[30] ),
    .B(_0308_));
 sg13g2_nand2_1 _0884_ (.Y(_0312_),
    .A(_0067_),
    .B(_0304_));
 sg13g2_a21oi_1 _0885_ (.A1(net164),
    .A2(_0289_),
    .Y(_0313_),
    .B1(_0001_));
 sg13g2_xor2_1 _0886_ (.B(_0297_),
    .A(\PWM_Generator.pwm_cnt[28] ),
    .X(_0314_));
 sg13g2_nor3_1 _0887_ (.A(_0291_),
    .B(_0313_),
    .C(_0314_),
    .Y(_0315_));
 sg13g2_nand4_1 _0888_ (.B(_0311_),
    .C(_0312_),
    .A(_0310_),
    .Y(_0316_),
    .D(_0315_));
 sg13g2_nor2b_1 _0889_ (.A(_0316_),
    .B_N(_0303_),
    .Y(_0317_));
 sg13g2_nand4_1 _0890_ (.B(net164),
    .C(_0002_),
    .A(net169),
    .Y(_0318_),
    .D(_0301_));
 sg13g2_nand3_1 _0891_ (.B(net152),
    .C(_0306_),
    .A(net169),
    .Y(_0319_));
 sg13g2_or2_1 _0892_ (.X(_0320_),
    .B(_0319_),
    .A(net150));
 sg13g2_o21ai_1 _0893_ (.B1(_0318_),
    .Y(_0321_),
    .A1(\PWM_Generator.pwm_cnt[26] ),
    .A2(_0320_));
 sg13g2_nand2_1 _0894_ (.Y(_0322_),
    .A(net152),
    .B(_0286_));
 sg13g2_nor2_1 _0895_ (.A(net170),
    .B(_0274_),
    .Y(_0323_));
 sg13g2_a21oi_2 _0896_ (.B1(_0323_),
    .Y(_0324_),
    .A2(_0322_),
    .A1(net170));
 sg13g2_and2_1 _0897_ (.A(net164),
    .B(_0324_),
    .X(_0325_));
 sg13g2_a21oi_1 _0898_ (.A1(net164),
    .A2(_0324_),
    .Y(_0326_),
    .B1(_0003_));
 sg13g2_a21oi_1 _0899_ (.A1(\PWM_Generator.pwm_cnt[26] ),
    .A2(_0320_),
    .Y(_0327_),
    .B1(_0326_));
 sg13g2_nand4_1 _0900_ (.B(net172),
    .C(net174),
    .A(net153),
    .Y(_0328_),
    .D(_0278_));
 sg13g2_nand4_1 _0901_ (.B(net152),
    .C(_0065_),
    .A(net170),
    .Y(_0329_),
    .D(_0292_));
 sg13g2_and2_1 _0902_ (.A(_0328_),
    .B(_0329_),
    .X(_0330_));
 sg13g2_or2_1 _0903_ (.X(_0331_),
    .B(_0330_),
    .A(net150));
 sg13g2_nor2_1 _0904_ (.A(\PWM_Generator.pwm_cnt[24] ),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_a21oi_1 _0905_ (.A1(_0003_),
    .A2(_0325_),
    .Y(_0333_),
    .B1(_0332_));
 sg13g2_nand2_1 _0906_ (.Y(_0334_),
    .A(\PWM_Generator.pwm_cnt[24] ),
    .B(_0331_));
 sg13g2_and4_1 _0907_ (.A(net153),
    .B(net173),
    .C(net166),
    .D(_0306_),
    .X(_0335_));
 sg13g2_nor4_1 _0908_ (.A(net169),
    .B(net152),
    .C(net151),
    .D(_0300_),
    .Y(_0336_));
 sg13g2_a22oi_1 _0909_ (.Y(_0337_),
    .B1(_0336_),
    .B2(_0004_),
    .A2(_0335_),
    .A1(_0069_));
 sg13g2_nand2b_1 _0910_ (.Y(_0338_),
    .B(\PWM_Generator.pwm_cnt[22] ),
    .A_N(_0335_));
 sg13g2_or2_1 _0911_ (.X(_0339_),
    .B(_0336_),
    .A(_0004_));
 sg13g2_and3_1 _0912_ (.X(_0340_),
    .A(_0337_),
    .B(_0338_),
    .C(_0339_));
 sg13g2_nor3_2 _0913_ (.A(net170),
    .B(_0287_),
    .C(_0288_),
    .Y(_0341_));
 sg13g2_and2_1 _0914_ (.A(net166),
    .B(_0341_),
    .X(_0342_));
 sg13g2_nand3_1 _0915_ (.B(_0294_),
    .C(_0295_),
    .A(_0063_),
    .Y(_0343_));
 sg13g2_nor2_1 _0916_ (.A(net150),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_a22oi_1 _0917_ (.Y(_0345_),
    .B1(_0344_),
    .B2(_0070_),
    .A2(_0342_),
    .A1(_0005_));
 sg13g2_or2_1 _0918_ (.X(_0346_),
    .B(_0342_),
    .A(_0005_));
 sg13g2_o21ai_1 _0919_ (.B1(\PWM_Generator.pwm_cnt[20] ),
    .Y(_0347_),
    .A1(net150),
    .A2(_0343_));
 sg13g2_nand4_1 _0920_ (.B(_0345_),
    .C(_0346_),
    .A(_0340_),
    .Y(_0348_),
    .D(_0347_));
 sg13g2_nor4_2 _0921_ (.A(net169),
    .B(net173),
    .C(net150),
    .Y(_0349_),
    .D(_0300_));
 sg13g2_or2_1 _0922_ (.X(_0350_),
    .B(_0349_),
    .A(_0006_));
 sg13g2_and4_1 _0923_ (.A(net153),
    .B(net152),
    .C(net166),
    .D(_0306_),
    .X(_0351_));
 sg13g2_a22oi_1 _0924_ (.Y(_0352_),
    .B1(_0351_),
    .B2(_0071_),
    .A2(_0349_),
    .A1(_0006_));
 sg13g2_inv_1 _0925_ (.Y(_0353_),
    .A(_0352_));
 sg13g2_nand2_1 _0926_ (.Y(_0354_),
    .A(_0350_),
    .B(_0353_));
 sg13g2_nand2b_1 _0927_ (.Y(_0355_),
    .B(\PWM_Generator.pwm_cnt[18] ),
    .A_N(_0351_));
 sg13g2_nand3_1 _0928_ (.B(_0352_),
    .C(_0355_),
    .A(_0350_),
    .Y(_0356_));
 sg13g2_nor4_2 _0929_ (.A(net170),
    .B(net172),
    .C(net174),
    .Y(_0357_),
    .D(_0293_));
 sg13g2_mux2_1 _0930_ (.A0(_0279_),
    .A1(_0357_),
    .S(net168),
    .X(_0358_));
 sg13g2_nand2_1 _0931_ (.Y(_0359_),
    .A(_0072_),
    .B(_0358_));
 sg13g2_nand3_1 _0932_ (.B(net152),
    .C(_0286_),
    .A(net153),
    .Y(_0360_));
 sg13g2_nor2_1 _0933_ (.A(net168),
    .B(_0275_),
    .Y(_0361_));
 sg13g2_a21o_1 _0934_ (.A2(_0360_),
    .A1(net167),
    .B1(_0361_),
    .X(_0362_));
 sg13g2_o21ai_1 _0935_ (.B1(_0359_),
    .Y(_0363_),
    .A1(\PWM_Generator.pwm_cnt[17] ),
    .A2(_0362_));
 sg13g2_nand2_1 _0936_ (.Y(_0364_),
    .A(\PWM_Generator.pwm_cnt[17] ),
    .B(_0362_));
 sg13g2_nand3b_1 _0937_ (.B(_0363_),
    .C(_0364_),
    .Y(_0365_),
    .A_N(_0356_));
 sg13g2_a21oi_1 _0938_ (.A1(_0354_),
    .A2(_0365_),
    .Y(_0366_),
    .B1(_0348_));
 sg13g2_nor2b_1 _0939_ (.A(_0345_),
    .B_N(_0346_),
    .Y(_0367_));
 sg13g2_and2_1 _0940_ (.A(_0340_),
    .B(_0367_),
    .X(_0368_));
 sg13g2_nor2b_1 _0941_ (.A(_0337_),
    .B_N(_0339_),
    .Y(_0369_));
 sg13g2_nor3_1 _0942_ (.A(_0366_),
    .B(_0368_),
    .C(_0369_),
    .Y(_0370_));
 sg13g2_nor4_1 _0943_ (.A(net150),
    .B(\PWM_Generator.pwm_cnt[28] ),
    .C(_0296_),
    .D(_0313_),
    .Y(_0371_));
 sg13g2_o21ai_1 _0944_ (.B1(_0311_),
    .Y(_0372_),
    .A1(_0291_),
    .A2(_0371_));
 sg13g2_a22oi_1 _0945_ (.Y(_0373_),
    .B1(_0310_),
    .B2(_0372_),
    .A2(_0304_),
    .A1(_0067_));
 sg13g2_nand4_1 _0946_ (.B(net173),
    .C(net151),
    .A(net169),
    .Y(_0374_),
    .D(_0299_));
 sg13g2_nor2_1 _0947_ (.A(_0073_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_nor3_1 _0948_ (.A(net164),
    .B(\PWM_Generator.pwm_cnt[14] ),
    .C(_0307_),
    .Y(_0376_));
 sg13g2_nor2_1 _0949_ (.A(_0375_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_o21ai_1 _0950_ (.B1(\PWM_Generator.pwm_cnt[14] ),
    .Y(_0378_),
    .A1(net165),
    .A2(_0307_));
 sg13g2_nand2_1 _0951_ (.Y(_0379_),
    .A(_0073_),
    .B(_0374_));
 sg13g2_nand3_1 _0952_ (.B(_0378_),
    .C(_0379_),
    .A(_0377_),
    .Y(_0380_));
 sg13g2_nor4_2 _0953_ (.A(net153),
    .B(net167),
    .C(_0287_),
    .Y(_0381_),
    .D(_0288_));
 sg13g2_nand2_1 _0954_ (.Y(_0382_),
    .A(_0008_),
    .B(_0381_));
 sg13g2_or3_1 _0955_ (.A(net165),
    .B(\PWM_Generator.pwm_cnt[12] ),
    .C(_0296_),
    .X(_0383_));
 sg13g2_nand2_1 _0956_ (.Y(_0384_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_or2_1 _0957_ (.X(_0385_),
    .B(_0381_),
    .A(_0008_));
 sg13g2_o21ai_1 _0958_ (.B1(\PWM_Generator.pwm_cnt[12] ),
    .Y(_0386_),
    .A1(net165),
    .A2(_0296_));
 sg13g2_nor4_2 _0959_ (.A(net153),
    .B(net173),
    .C(net166),
    .Y(_0387_),
    .D(_0300_));
 sg13g2_or2_1 _0960_ (.X(_0388_),
    .B(_0387_),
    .A(_0009_));
 sg13g2_nand3_1 _0961_ (.B(_0386_),
    .C(_0388_),
    .A(_0385_),
    .Y(_0389_));
 sg13g2_o21ai_1 _0962_ (.B1(\PWM_Generator.pwm_cnt[10] ),
    .Y(_0390_),
    .A1(net165),
    .A2(_0319_));
 sg13g2_a21oi_1 _0963_ (.A1(_0066_),
    .A2(_0324_),
    .Y(_0391_),
    .B1(_0010_));
 sg13g2_nand3b_1 _0964_ (.B(_0074_),
    .C(_0066_),
    .Y(_0392_),
    .A_N(_0330_));
 sg13g2_nor3_1 _0965_ (.A(net164),
    .B(\PWM_Generator.pwm_cnt[10] ),
    .C(_0319_),
    .Y(_0393_));
 sg13g2_a21oi_1 _0966_ (.A1(_0009_),
    .A2(_0387_),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_nand3_1 _0967_ (.B(_0010_),
    .C(_0324_),
    .A(net151),
    .Y(_0395_));
 sg13g2_o21ai_1 _0968_ (.B1(\PWM_Generator.pwm_cnt[8] ),
    .Y(_0396_),
    .A1(net167),
    .A2(_0330_));
 sg13g2_and4_1 _0969_ (.A(_0382_),
    .B(_0383_),
    .C(_0385_),
    .D(_0386_),
    .X(_0397_));
 sg13g2_nand4_1 _0970_ (.B(_0378_),
    .C(_0379_),
    .A(_0377_),
    .Y(_0398_),
    .D(_0397_));
 sg13g2_nand3_1 _0971_ (.B(_0390_),
    .C(_0394_),
    .A(_0388_),
    .Y(_0399_));
 sg13g2_and2_1 _0972_ (.A(_0392_),
    .B(_0396_),
    .X(_0400_));
 sg13g2_nand3b_1 _0973_ (.B(_0395_),
    .C(_0400_),
    .Y(_0401_),
    .A_N(_0391_));
 sg13g2_nor3_2 _0974_ (.A(_0398_),
    .B(_0399_),
    .C(_0401_),
    .Y(_0402_));
 sg13g2_nor4_2 _0975_ (.A(net171),
    .B(net172),
    .C(net168),
    .Y(_0403_),
    .D(_0300_));
 sg13g2_nand2_1 _0976_ (.Y(_0404_),
    .A(_0013_),
    .B(_0403_));
 sg13g2_nand4_1 _0977_ (.B(_0064_),
    .C(net151),
    .A(_0063_),
    .Y(_0405_),
    .D(_0306_));
 sg13g2_o21ai_1 _0978_ (.B1(_0404_),
    .Y(_0406_),
    .A1(\PWM_Generator.pwm_cnt[2] ),
    .A2(_0405_));
 sg13g2_nand2_1 _0979_ (.Y(_0407_),
    .A(\PWM_Generator.pwm_cnt[2] ),
    .B(_0405_));
 sg13g2_nor3_1 _0980_ (.A(net167),
    .B(\PWM_Generator.pwm_cnt[1] ),
    .C(_0360_),
    .Y(_0408_));
 sg13g2_o21ai_1 _0981_ (.B1(\PWM_Generator.pwm_cnt[1] ),
    .Y(_0409_),
    .A1(net167),
    .A2(_0360_));
 sg13g2_nand2_1 _0982_ (.Y(_0410_),
    .A(_0066_),
    .B(_0357_));
 sg13g2_nand2_1 _0983_ (.Y(_0411_),
    .A(\PWM_Generator.pwm_cnt[0] ),
    .B(_0410_));
 sg13g2_a21o_1 _0984_ (.A2(_0411_),
    .A1(_0409_),
    .B1(_0408_),
    .X(_0412_));
 sg13g2_a21oi_1 _0985_ (.A1(_0407_),
    .A2(_0412_),
    .Y(_0413_),
    .B1(_0406_));
 sg13g2_nor4_2 _0986_ (.A(net170),
    .B(net152),
    .C(net167),
    .Y(_0414_),
    .D(_0300_));
 sg13g2_and4_1 _0987_ (.A(net153),
    .B(net172),
    .C(net151),
    .D(_0306_),
    .X(_0415_));
 sg13g2_a22oi_1 _0988_ (.Y(_0416_),
    .B1(_0415_),
    .B2(_0076_),
    .A2(_0414_),
    .A1(_0011_));
 sg13g2_nand2b_1 _0989_ (.Y(_0417_),
    .B(\PWM_Generator.pwm_cnt[6] ),
    .A_N(_0415_));
 sg13g2_or2_1 _0990_ (.X(_0418_),
    .B(_0414_),
    .A(_0011_));
 sg13g2_and3_1 _0991_ (.X(_0419_),
    .A(_0416_),
    .B(_0417_),
    .C(_0418_));
 sg13g2_or3_1 _0992_ (.A(net167),
    .B(\PWM_Generator.pwm_cnt[4] ),
    .C(_0343_),
    .X(_0420_));
 sg13g2_nand3_1 _0993_ (.B(_0012_),
    .C(_0341_),
    .A(net151),
    .Y(_0421_));
 sg13g2_a21oi_1 _0994_ (.A1(net151),
    .A2(_0341_),
    .Y(_0422_),
    .B1(_0012_));
 sg13g2_o21ai_1 _0995_ (.B1(\PWM_Generator.pwm_cnt[4] ),
    .Y(_0423_),
    .A1(net167),
    .A2(_0343_));
 sg13g2_nor2b_1 _0996_ (.A(_0422_),
    .B_N(_0423_),
    .Y(_0424_));
 sg13g2_nand4_1 _0997_ (.B(_0420_),
    .C(_0421_),
    .A(_0419_),
    .Y(_0425_),
    .D(_0424_));
 sg13g2_nor2_1 _0998_ (.A(_0013_),
    .B(_0403_),
    .Y(_0426_));
 sg13g2_or2_1 _0999_ (.X(_0427_),
    .B(_0403_),
    .A(_0013_));
 sg13g2_nor3_1 _1000_ (.A(_0413_),
    .B(_0425_),
    .C(_0426_),
    .Y(_0428_));
 sg13g2_o21ai_1 _1001_ (.B1(_0421_),
    .Y(_0429_),
    .A1(_0420_),
    .A2(_0422_));
 sg13g2_nand2b_1 _1002_ (.Y(_0430_),
    .B(_0418_),
    .A_N(_0416_));
 sg13g2_nand2_1 _1003_ (.Y(_0431_),
    .A(_0419_),
    .B(_0429_));
 sg13g2_nand2_1 _1004_ (.Y(_0432_),
    .A(_0430_),
    .B(_0431_));
 sg13g2_o21ai_1 _1005_ (.B1(_0402_),
    .Y(_0433_),
    .A1(_0428_),
    .A2(_0432_));
 sg13g2_o21ai_1 _1006_ (.B1(_0395_),
    .Y(_0434_),
    .A1(_0391_),
    .A2(_0392_));
 sg13g2_a221oi_1 _1007_ (.B2(_0434_),
    .C1(_0393_),
    .B1(_0390_),
    .A1(_0009_),
    .Y(_0435_),
    .A2(_0387_));
 sg13g2_or4_1 _1008_ (.A(_0380_),
    .B(_0384_),
    .C(_0389_),
    .D(_0435_),
    .X(_0436_));
 sg13g2_o21ai_1 _1009_ (.B1(_0379_),
    .Y(_0437_),
    .A1(_0375_),
    .A2(_0376_));
 sg13g2_nand3b_1 _1010_ (.B(_0384_),
    .C(_0385_),
    .Y(_0438_),
    .A_N(_0380_));
 sg13g2_nand4_1 _1011_ (.B(_0436_),
    .C(_0437_),
    .A(_0433_),
    .Y(_0439_),
    .D(_0438_));
 sg13g2_nand4_1 _1012_ (.B(_0327_),
    .C(_0333_),
    .A(_0303_),
    .Y(_0440_),
    .D(_0334_));
 sg13g2_or3_1 _1013_ (.A(_0316_),
    .B(_0321_),
    .C(_0440_),
    .X(_0441_));
 sg13g2_o21ai_1 _1014_ (.B1(_0364_),
    .Y(_0442_),
    .A1(_0072_),
    .A2(_0358_));
 sg13g2_or2_1 _1015_ (.X(_0443_),
    .B(_0442_),
    .A(_0363_));
 sg13g2_nand2b_1 _1016_ (.Y(_0444_),
    .B(_0327_),
    .A_N(_0333_));
 sg13g2_nand2b_1 _1017_ (.Y(_0445_),
    .B(_0444_),
    .A_N(_0321_));
 sg13g2_nor2_1 _1018_ (.A(_0370_),
    .B(_0441_),
    .Y(_0446_));
 sg13g2_a21oi_1 _1019_ (.A1(_0317_),
    .A2(_0445_),
    .Y(_0447_),
    .B1(_0373_));
 sg13g2_nor4_2 _1020_ (.A(_0348_),
    .B(_0356_),
    .C(_0441_),
    .Y(_0448_),
    .D(_0443_));
 sg13g2_a21oi_1 _1021_ (.A1(_0439_),
    .A2(_0448_),
    .Y(_0449_),
    .B1(_0446_));
 sg13g2_a21o_1 _1022_ (.A2(_0449_),
    .A1(_0447_),
    .B1(_0284_),
    .X(_0450_));
 sg13g2_xnor2_1 _1023_ (.Y(_0451_),
    .A(_0077_),
    .B(_0410_));
 sg13g2_nor2_1 _1024_ (.A(_0408_),
    .B(_0451_),
    .Y(_0452_));
 sg13g2_nand4_1 _1025_ (.B(_0409_),
    .C(_0427_),
    .A(_0407_),
    .Y(_0453_),
    .D(_0452_));
 sg13g2_nor4_1 _1026_ (.A(_0284_),
    .B(_0406_),
    .C(_0425_),
    .D(_0453_),
    .Y(_0454_));
 sg13g2_and2_1 _1027_ (.A(_0402_),
    .B(_0454_),
    .X(_0455_));
 sg13g2_a22oi_1 _1028_ (.Y(_0456_),
    .B1(_0448_),
    .B2(_0455_),
    .A2(_0283_),
    .A1(_0281_));
 sg13g2_a21oi_1 _1029_ (.A1(_0450_),
    .A2(_0456_),
    .Y(_0050_),
    .B1(net145));
 sg13g2_and4_1 _1030_ (.A(uo_out[6]),
    .B(uo_out[5]),
    .C(uo_out[3]),
    .D(uo_out[1]),
    .X(_0457_));
 sg13g2_nand3b_1 _1031_ (.B(uo_out[2]),
    .C(_0457_),
    .Y(_0458_),
    .A_N(uo_out[4]));
 sg13g2_xnor2_1 _1032_ (.Y(_0459_),
    .A(\PWM_Generator.fprev[0] ),
    .B(uo_out[1]));
 sg13g2_nand3_1 _1033_ (.B(net143),
    .C(_0459_),
    .A(net1),
    .Y(_0460_));
 sg13g2_nor2_1 _1034_ (.A(net142),
    .B(_0460_),
    .Y(_0461_));
 sg13g2_nor2_1 _1035_ (.A(net181),
    .B(net135),
    .Y(_0462_));
 sg13g2_nor2_1 _1036_ (.A(_0461_),
    .B(_0462_),
    .Y(_0051_));
 sg13g2_nor2b_1 _1037_ (.A(net177),
    .B_N(_0204_),
    .Y(_0463_));
 sg13g2_nand2_1 _1038_ (.Y(_0464_),
    .A(\PWM_Generator.fprev[1] ),
    .B(uo_out[2]));
 sg13g2_xor2_1 _1039_ (.B(uo_out[2]),
    .A(\PWM_Generator.fprev[1] ),
    .X(_0465_));
 sg13g2_a21o_1 _1040_ (.A2(uo_out[1]),
    .A1(\PWM_Generator.fprev[0] ),
    .B1(_0465_),
    .X(_0466_));
 sg13g2_nand3_1 _1041_ (.B(uo_out[1]),
    .C(_0465_),
    .A(\PWM_Generator.fprev[0] ),
    .Y(_0467_));
 sg13g2_nand3_1 _1042_ (.B(_0466_),
    .C(_0467_),
    .A(_0458_),
    .Y(_0468_));
 sg13g2_nor2b_1 _1043_ (.A(net142),
    .B_N(_0468_),
    .Y(_0469_));
 sg13g2_nor3_1 _1044_ (.A(net145),
    .B(_0463_),
    .C(_0469_),
    .Y(_0052_));
 sg13g2_nor2b_1 _1045_ (.A(net176),
    .B_N(net141),
    .Y(_0470_));
 sg13g2_nand2_1 _1046_ (.Y(_0471_),
    .A(\PWM_Generator.fprev[2] ),
    .B(uo_out[3]));
 sg13g2_xnor2_1 _1047_ (.Y(_0472_),
    .A(\PWM_Generator.fprev[2] ),
    .B(uo_out[3]));
 sg13g2_nand3_1 _1048_ (.B(_0467_),
    .C(_0472_),
    .A(_0464_),
    .Y(_0473_));
 sg13g2_a21o_1 _1049_ (.A2(_0467_),
    .A1(_0464_),
    .B1(_0472_),
    .X(_0474_));
 sg13g2_nand3_1 _1050_ (.B(_0473_),
    .C(_0474_),
    .A(net143),
    .Y(_0475_));
 sg13g2_nor2b_1 _1051_ (.A(net141),
    .B_N(_0475_),
    .Y(_0476_));
 sg13g2_nor3_1 _1052_ (.A(net144),
    .B(_0470_),
    .C(_0476_),
    .Y(_0053_));
 sg13g2_nor2b_1 _1053_ (.A(net185),
    .B_N(net139),
    .Y(_0477_));
 sg13g2_nand2_1 _1054_ (.Y(_0478_),
    .A(\PWM_Generator.fprev[3] ),
    .B(uo_out[4]));
 sg13g2_xnor2_1 _1055_ (.Y(_0479_),
    .A(net94),
    .B(uo_out[4]));
 sg13g2_and2_1 _1056_ (.A(_0471_),
    .B(_0474_),
    .X(_0480_));
 sg13g2_or2_1 _1057_ (.X(_0481_),
    .B(_0480_),
    .A(_0479_));
 sg13g2_nand2_1 _1058_ (.Y(_0482_),
    .A(net143),
    .B(_0481_));
 sg13g2_a21oi_1 _1059_ (.A1(_0479_),
    .A2(_0480_),
    .Y(_0483_),
    .B1(_0482_));
 sg13g2_nor2_1 _1060_ (.A(net139),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_nor3_1 _1061_ (.A(net144),
    .B(_0477_),
    .C(_0484_),
    .Y(_0054_));
 sg13g2_nand2_1 _1062_ (.Y(_0485_),
    .A(_0478_),
    .B(_0481_));
 sg13g2_xnor2_1 _1063_ (.Y(_0486_),
    .A(\PWM_Generator.fprev[4] ),
    .B(uo_out[5]));
 sg13g2_inv_1 _1064_ (.Y(_0487_),
    .A(_0486_));
 sg13g2_a21oi_1 _1065_ (.A1(_0478_),
    .A2(_0481_),
    .Y(_0488_),
    .B1(_0486_));
 sg13g2_o21ai_1 _1066_ (.B1(net143),
    .Y(_0489_),
    .A1(_0485_),
    .A2(_0487_));
 sg13g2_nor2_1 _1067_ (.A(_0488_),
    .B(_0489_),
    .Y(_0490_));
 sg13g2_nor2b_1 _1068_ (.A(net180),
    .B_N(net140),
    .Y(_0491_));
 sg13g2_nor2_1 _1069_ (.A(net140),
    .B(_0490_),
    .Y(_0492_));
 sg13g2_nor3_1 _1070_ (.A(net144),
    .B(_0491_),
    .C(_0492_),
    .Y(_0055_));
 sg13g2_nor2b_1 _1071_ (.A(net131),
    .B_N(net139),
    .Y(_0493_));
 sg13g2_a21oi_1 _1072_ (.A1(net92),
    .A2(uo_out[5]),
    .Y(_0494_),
    .B1(_0488_));
 sg13g2_xnor2_1 _1073_ (.Y(_0495_),
    .A(net85),
    .B(uo_out[6]));
 sg13g2_o21ai_1 _1074_ (.B1(net143),
    .Y(_0496_),
    .A1(_0494_),
    .A2(_0495_));
 sg13g2_a21oi_1 _1075_ (.A1(_0494_),
    .A2(_0495_),
    .Y(_0497_),
    .B1(_0496_));
 sg13g2_nor2_1 _1076_ (.A(net139),
    .B(_0497_),
    .Y(_0498_));
 sg13g2_nor3_1 _1077_ (.A(net144),
    .B(_0493_),
    .C(_0498_),
    .Y(_0056_));
 sg13g2_nand2_1 _1078_ (.Y(_0499_),
    .A(net99),
    .B(net142));
 sg13g2_nand2_1 _1079_ (.Y(_0500_),
    .A(uo_out[1]),
    .B(_0458_));
 sg13g2_or2_1 _1080_ (.X(_0501_),
    .B(_0500_),
    .A(net142));
 sg13g2_a21oi_1 _1081_ (.A1(_0499_),
    .A2(_0501_),
    .Y(_0057_),
    .B1(net145));
 sg13g2_nand2_1 _1082_ (.Y(_0502_),
    .A(net88),
    .B(net142));
 sg13g2_nand2_1 _1083_ (.Y(_0503_),
    .A(uo_out[2]),
    .B(_0458_));
 sg13g2_or2_1 _1084_ (.X(_0504_),
    .B(_0503_),
    .A(net142));
 sg13g2_a21oi_1 _1085_ (.A1(_0502_),
    .A2(_0504_),
    .Y(_0058_),
    .B1(net145));
 sg13g2_nand2_1 _1086_ (.Y(_0505_),
    .A(net97),
    .B(net141));
 sg13g2_nand2_1 _1087_ (.Y(_0506_),
    .A(uo_out[3]),
    .B(net143));
 sg13g2_or2_1 _1088_ (.X(_0507_),
    .B(_0506_),
    .A(net141));
 sg13g2_a21oi_1 _1089_ (.A1(_0505_),
    .A2(_0507_),
    .Y(_0059_),
    .B1(net144));
 sg13g2_nor2b_1 _1090_ (.A(net94),
    .B_N(net139),
    .Y(_0508_));
 sg13g2_nor2_1 _1091_ (.A(uo_out[4]),
    .B(net139),
    .Y(_0509_));
 sg13g2_nor3_1 _1092_ (.A(net144),
    .B(_0508_),
    .C(_0509_),
    .Y(_0060_));
 sg13g2_nand2_1 _1093_ (.Y(_0510_),
    .A(net92),
    .B(net139));
 sg13g2_nand2_1 _1094_ (.Y(_0511_),
    .A(uo_out[5]),
    .B(net143));
 sg13g2_or2_1 _1095_ (.X(_0512_),
    .B(_0511_),
    .A(net139));
 sg13g2_a21oi_1 _1096_ (.A1(_0510_),
    .A2(_0512_),
    .Y(_0061_),
    .B1(net144));
 sg13g2_nand2_1 _1097_ (.Y(_0513_),
    .A(net85),
    .B(net140));
 sg13g2_nand2_1 _1098_ (.Y(_0514_),
    .A(uo_out[6]),
    .B(net143));
 sg13g2_or2_1 _1099_ (.X(_0515_),
    .B(_0514_),
    .A(net140));
 sg13g2_a21oi_1 _1100_ (.A1(_0513_),
    .A2(_0515_),
    .Y(_0062_),
    .B1(net144));
 sg13g2_dfrbp_1 _1101_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net71),
    .D(_0014_),
    .Q_N(\PWM_Generator._pwm_cnt_T_1[0] ),
    .Q(\PWM_Generator.pwm_cnt[0] ));
 sg13g2_dfrbp_1 _1102_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net67),
    .D(_0015_),
    .Q_N(_0549_),
    .Q(\PWM_Generator.pwm_cnt[1] ));
 sg13g2_dfrbp_1 _1103_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net66),
    .D(_0016_),
    .Q_N(_0548_),
    .Q(\PWM_Generator.pwm_cnt[2] ));
 sg13g2_dfrbp_1 _1104_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net65),
    .D(_0017_),
    .Q_N(_0013_),
    .Q(\PWM_Generator.pwm_cnt[3] ));
 sg13g2_dfrbp_1 _1105_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net64),
    .D(_0018_),
    .Q_N(_0547_),
    .Q(\PWM_Generator.pwm_cnt[4] ));
 sg13g2_dfrbp_1 _1106_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net63),
    .D(_0019_),
    .Q_N(_0012_),
    .Q(\PWM_Generator.pwm_cnt[5] ));
 sg13g2_dfrbp_1 _1107_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net62),
    .D(_0020_),
    .Q_N(_0546_),
    .Q(\PWM_Generator.pwm_cnt[6] ));
 sg13g2_dfrbp_1 _1108_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net61),
    .D(_0021_),
    .Q_N(_0011_),
    .Q(\PWM_Generator.pwm_cnt[7] ));
 sg13g2_dfrbp_1 _1109_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net60),
    .D(_0022_),
    .Q_N(_0545_),
    .Q(\PWM_Generator.pwm_cnt[8] ));
 sg13g2_dfrbp_1 _1110_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net59),
    .D(_0023_),
    .Q_N(_0010_),
    .Q(\PWM_Generator.pwm_cnt[9] ));
 sg13g2_dfrbp_1 _1111_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net58),
    .D(_0024_),
    .Q_N(_0544_),
    .Q(\PWM_Generator.pwm_cnt[10] ));
 sg13g2_dfrbp_1 _1112_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net57),
    .D(_0025_),
    .Q_N(_0009_),
    .Q(\PWM_Generator.pwm_cnt[11] ));
 sg13g2_dfrbp_1 _1113_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net56),
    .D(_0026_),
    .Q_N(_0543_),
    .Q(\PWM_Generator.pwm_cnt[12] ));
 sg13g2_dfrbp_1 _1114_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net55),
    .D(_0027_),
    .Q_N(_0008_),
    .Q(\PWM_Generator.pwm_cnt[13] ));
 sg13g2_dfrbp_1 _1115_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net54),
    .D(_0028_),
    .Q_N(_0542_),
    .Q(\PWM_Generator.pwm_cnt[14] ));
 sg13g2_dfrbp_1 _1116_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net53),
    .D(_0029_),
    .Q_N(_0007_),
    .Q(\PWM_Generator.pwm_cnt[15] ));
 sg13g2_dfrbp_1 _1117_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net52),
    .D(_0030_),
    .Q_N(_0541_),
    .Q(\PWM_Generator.pwm_cnt[16] ));
 sg13g2_dfrbp_1 _1118_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net51),
    .D(_0031_),
    .Q_N(_0540_),
    .Q(\PWM_Generator.pwm_cnt[17] ));
 sg13g2_dfrbp_1 _1119_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net50),
    .D(_0032_),
    .Q_N(_0539_),
    .Q(\PWM_Generator.pwm_cnt[18] ));
 sg13g2_dfrbp_1 _1120_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net49),
    .D(_0033_),
    .Q_N(_0006_),
    .Q(\PWM_Generator.pwm_cnt[19] ));
 sg13g2_dfrbp_1 _1121_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net48),
    .D(_0034_),
    .Q_N(_0538_),
    .Q(\PWM_Generator.pwm_cnt[20] ));
 sg13g2_dfrbp_1 _1122_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net47),
    .D(_0035_),
    .Q_N(_0005_),
    .Q(\PWM_Generator.pwm_cnt[21] ));
 sg13g2_dfrbp_1 _1123_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net46),
    .D(_0036_),
    .Q_N(_0537_),
    .Q(\PWM_Generator.pwm_cnt[22] ));
 sg13g2_dfrbp_1 _1124_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net45),
    .D(_0037_),
    .Q_N(_0004_),
    .Q(\PWM_Generator.pwm_cnt[23] ));
 sg13g2_dfrbp_1 _1125_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net44),
    .D(_0038_),
    .Q_N(_0536_),
    .Q(\PWM_Generator.pwm_cnt[24] ));
 sg13g2_dfrbp_1 _1126_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net43),
    .D(_0039_),
    .Q_N(_0003_),
    .Q(\PWM_Generator.pwm_cnt[25] ));
 sg13g2_dfrbp_1 _1127_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net42),
    .D(_0040_),
    .Q_N(_0535_),
    .Q(\PWM_Generator.pwm_cnt[26] ));
 sg13g2_dfrbp_1 _1128_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net41),
    .D(_0041_),
    .Q_N(_0002_),
    .Q(\PWM_Generator.pwm_cnt[27] ));
 sg13g2_dfrbp_1 _1129_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net40),
    .D(_0042_),
    .Q_N(_0534_),
    .Q(\PWM_Generator.pwm_cnt[28] ));
 sg13g2_dfrbp_1 _1130_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net39),
    .D(net80),
    .Q_N(_0001_),
    .Q(\PWM_Generator.pwm_cnt[29] ));
 sg13g2_dfrbp_1 _1131_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net38),
    .D(_0044_),
    .Q_N(_0533_),
    .Q(\PWM_Generator.pwm_cnt[30] ));
 sg13g2_dfrbp_1 _1132_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net37),
    .D(_0045_),
    .Q_N(_0000_),
    .Q(\PWM_Generator.pwm_cnt[31] ));
 sg13g2_dfrbp_1 _1133_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net36),
    .D(_0046_),
    .Q_N(_0532_),
    .Q(\PWM_Generator.pwm_cnt[32] ));
 sg13g2_dfrbp_1 _1134_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net35),
    .D(_0047_),
    .Q_N(_0531_),
    .Q(\PWM_Generator.pwm_cnt[33] ));
 sg13g2_dfrbp_1 _1135_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net34),
    .D(_0048_),
    .Q_N(_0530_),
    .Q(\PWM_Generator.pwm_cnt[34] ));
 sg13g2_dfrbp_1 _1136_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net33),
    .D(_0049_),
    .Q_N(_0529_),
    .Q(\PWM_Generator.pwm_cnt[35] ));
 sg13g2_dfrbp_1 _1137_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net32),
    .D(_0050_),
    .Q_N(_0528_),
    .Q(\PWM_Generator.pwm_out ));
 sg13g2_dfrbp_1 _1138_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net31),
    .D(_0051_),
    .Q_N(_0527_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1139_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net29),
    .D(_0052_),
    .Q_N(_0526_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1140_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net76),
    .D(_0053_),
    .Q_N(_0525_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1141_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net74),
    .D(_0054_),
    .Q_N(_0524_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1142_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net72),
    .D(_0055_),
    .Q_N(_0523_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1143_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net70),
    .D(_0056_),
    .Q_N(_0522_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1144_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net68),
    .D(net100),
    .Q_N(_0521_),
    .Q(\PWM_Generator.fprev[0] ));
 sg13g2_dfrbp_1 _1145_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net77),
    .D(net89),
    .Q_N(_0520_),
    .Q(\PWM_Generator.fprev[1] ));
 sg13g2_dfrbp_1 _1146_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net73),
    .D(net98),
    .Q_N(_0519_),
    .Q(\PWM_Generator.fprev[2] ));
 sg13g2_dfrbp_1 _1147_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net69),
    .D(net95),
    .Q_N(_0518_),
    .Q(\PWM_Generator.fprev[3] ));
 sg13g2_dfrbp_1 _1148_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net75),
    .D(net93),
    .Q_N(_0517_),
    .Q(\PWM_Generator.fprev[4] ));
 sg13g2_dfrbp_1 _1149_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net30),
    .D(net86),
    .Q_N(_0516_),
    .Q(\PWM_Generator.fprev[5] ));
 sg13g2_tiehi _1149__30 (.L_HI(net30));
 sg13g2_tiehi _1138__31 (.L_HI(net31));
 sg13g2_tiehi _1137__32 (.L_HI(net32));
 sg13g2_tiehi _1136__33 (.L_HI(net33));
 sg13g2_tiehi _1135__34 (.L_HI(net34));
 sg13g2_tiehi _1134__35 (.L_HI(net35));
 sg13g2_tiehi _1133__36 (.L_HI(net36));
 sg13g2_tiehi _1132__37 (.L_HI(net37));
 sg13g2_tiehi _1131__38 (.L_HI(net38));
 sg13g2_tiehi _1130__39 (.L_HI(net39));
 sg13g2_tiehi _1129__40 (.L_HI(net40));
 sg13g2_tiehi _1128__41 (.L_HI(net41));
 sg13g2_tiehi _1127__42 (.L_HI(net42));
 sg13g2_tiehi _1126__43 (.L_HI(net43));
 sg13g2_tiehi _1125__44 (.L_HI(net44));
 sg13g2_tiehi _1124__45 (.L_HI(net45));
 sg13g2_tiehi _1123__46 (.L_HI(net46));
 sg13g2_tiehi _1122__47 (.L_HI(net47));
 sg13g2_tiehi _1121__48 (.L_HI(net48));
 sg13g2_tiehi _1120__49 (.L_HI(net49));
 sg13g2_tiehi _1119__50 (.L_HI(net50));
 sg13g2_tiehi _1118__51 (.L_HI(net51));
 sg13g2_tiehi _1117__52 (.L_HI(net52));
 sg13g2_tiehi _1116__53 (.L_HI(net53));
 sg13g2_tiehi _1115__54 (.L_HI(net54));
 sg13g2_tiehi _1114__55 (.L_HI(net55));
 sg13g2_tiehi _1113__56 (.L_HI(net56));
 sg13g2_tiehi _1112__57 (.L_HI(net57));
 sg13g2_tiehi _1111__58 (.L_HI(net58));
 sg13g2_tiehi _1110__59 (.L_HI(net59));
 sg13g2_tiehi _1109__60 (.L_HI(net60));
 sg13g2_tiehi _1108__61 (.L_HI(net61));
 sg13g2_tiehi _1107__62 (.L_HI(net62));
 sg13g2_tiehi _1106__63 (.L_HI(net63));
 sg13g2_tiehi _1105__64 (.L_HI(net64));
 sg13g2_tiehi _1104__65 (.L_HI(net65));
 sg13g2_tiehi _1103__66 (.L_HI(net66));
 sg13g2_tiehi _1102__67 (.L_HI(net67));
 sg13g2_tiehi _1144__68 (.L_HI(net68));
 sg13g2_tiehi _1147__69 (.L_HI(net69));
 sg13g2_tiehi _1143__70 (.L_HI(net70));
 sg13g2_tiehi _1101__71 (.L_HI(net71));
 sg13g2_tiehi _1142__72 (.L_HI(net72));
 sg13g2_tiehi _1146__73 (.L_HI(net73));
 sg13g2_tiehi _1141__74 (.L_HI(net74));
 sg13g2_tiehi _1148__75 (.L_HI(net75));
 sg13g2_tiehi _1140__76 (.L_HI(net76));
 sg13g2_tiehi _1145__77 (.L_HI(net77));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_anas_7193_14 (.L_LO(net14));
 sg13g2_tielo tt_um_anas_7193_15 (.L_LO(net15));
 sg13g2_tielo tt_um_anas_7193_16 (.L_LO(net16));
 sg13g2_tielo tt_um_anas_7193_17 (.L_LO(net17));
 sg13g2_tielo tt_um_anas_7193_18 (.L_LO(net18));
 sg13g2_tielo tt_um_anas_7193_19 (.L_LO(net19));
 sg13g2_tielo tt_um_anas_7193_20 (.L_LO(net20));
 sg13g2_tielo tt_um_anas_7193_21 (.L_LO(net21));
 sg13g2_tielo tt_um_anas_7193_22 (.L_LO(net22));
 sg13g2_tielo tt_um_anas_7193_23 (.L_LO(net23));
 sg13g2_tielo tt_um_anas_7193_24 (.L_LO(net24));
 sg13g2_tielo tt_um_anas_7193_25 (.L_LO(net25));
 sg13g2_tielo tt_um_anas_7193_26 (.L_LO(net26));
 sg13g2_tielo tt_um_anas_7193_27 (.L_LO(net27));
 sg13g2_tielo tt_um_anas_7193_28 (.L_LO(net28));
 sg13g2_tiehi _1139__29 (.L_HI(net29));
 sg13g2_buf_1 _1215_ (.A(\PWM_Generator.pwm_out ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1216_ (.A(ena),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout133 (.A(net135),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net138));
 sg13g2_buf_2 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net138));
 sg13g2_buf_2 fanout138 (.A(_0205_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net141),
    .X(net139));
 sg13g2_buf_1 fanout140 (.A(net141),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_0204_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_0458_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(net145),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_0080_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(net147),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_0079_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(net149),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_0078_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(net151),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_0066_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_0064_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_0063_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(net155),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(net156),
    .X(net155));
 sg13g2_buf_1 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(uio_in[4]),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(net160),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(uio_in[3]),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(uio_in[2]),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(uio_in[2]),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(net9),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(net166),
    .X(net164));
 sg13g2_buf_1 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(ui_in[4]),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(ui_in[4]),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(ui_in[4]),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(net171),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(ui_in[3]),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(net4),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(net4),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(net3),
    .X(net174));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[5]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[6]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[7]),
    .X(net12));
 sg13g2_tielo tt_um_anas_7193_13 (.L_LO(net13));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\PWM_Generator.pwm_cnt[29] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0259_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0043_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold4 (.A(\PWM_Generator.pwm_cnt[34] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0269_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold6 (.A(\PWM_Generator.pwm_cnt[13] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0229_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold8 (.A(\PWM_Generator.fprev[5] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0062_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold10 (.A(\PWM_Generator.pwm_cnt[35] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold11 (.A(\PWM_Generator.fprev[1] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0058_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold13 (.A(\PWM_Generator.pwm_cnt[31] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0263_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold15 (.A(\PWM_Generator.fprev[4] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0061_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold17 (.A(\PWM_Generator.fprev[3] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0060_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold19 (.A(\PWM_Generator._pwm_cnt_T_1[0] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold20 (.A(\PWM_Generator.fprev[2] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0059_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold22 (.A(\PWM_Generator.fprev[0] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0057_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold24 (.A(\PWM_Generator.pwm_cnt[27] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0256_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold26 (.A(\PWM_Generator.pwm_cnt[6] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0216_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold28 (.A(\PWM_Generator.pwm_cnt[7] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold29 (.A(\PWM_Generator.pwm_cnt[15] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0233_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold31 (.A(\PWM_Generator.pwm_cnt[3] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0210_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold33 (.A(\PWM_Generator.pwm_cnt[11] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0226_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold35 (.A(\PWM_Generator.pwm_cnt[0] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0206_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold37 (.A(\PWM_Generator.pwm_cnt[9] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0224_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold39 (.A(\PWM_Generator.pwm_cnt[8] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold40 (.A(\PWM_Generator.pwm_cnt[23] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0248_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold42 (.A(\PWM_Generator.pwm_cnt[16] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold43 (.A(\PWM_Generator.pwm_cnt[17] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold44 (.A(\PWM_Generator.pwm_cnt[25] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0252_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold46 (.A(\PWM_Generator.pwm_cnt[2] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0208_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold48 (.A(\PWM_Generator.pwm_cnt[19] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold49 (.A(\PWM_Generator.pwm_cnt[5] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0213_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold51 (.A(\PWM_Generator.pwm_cnt[21] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0244_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold53 (.A(\PWM_Generator.pwm_cnt[4] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold54 (.A(uo_out[6]),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold55 (.A(\PWM_Generator.pwm_cnt[14] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold56 (.A(\PWM_Generator.pwm_cnt[20] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold57 (.A(uo_out[3]),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold58 (.A(uo_out[2]),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold59 (.A(\PWM_Generator.pwm_cnt[12] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold60 (.A(\PWM_Generator.pwm_cnt[28] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold61 (.A(uo_out[5]),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold62 (.A(uo_out[1]),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold63 (.A(\PWM_Generator.pwm_cnt[24] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0250_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold65 (.A(\PWM_Generator.pwm_cnt[18] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold66 (.A(uo_out[4]),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold67 (.A(\PWM_Generator.pwm_cnt[22] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold68 (.A(\PWM_Generator.pwm_cnt[33] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold69 (.A(\PWM_Generator.pwm_cnt[26] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold70 (.A(\PWM_Generator.pwm_cnt[30] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold71 (.A(\PWM_Generator.pwm_cnt[32] ),
    .X(net190));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_4 FILLER_18_294 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_decap_4 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_307 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_fill_2 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_fill_2 FILLER_20_203 ();
 sg13g2_fill_1 FILLER_20_213 ();
 sg13g2_decap_8 FILLER_20_227 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_fill_1 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_241 ();
 sg13g2_fill_1 FILLER_20_309 ();
 sg13g2_fill_2 FILLER_20_319 ();
 sg13g2_fill_1 FILLER_20_321 ();
 sg13g2_fill_1 FILLER_20_335 ();
 sg13g2_fill_2 FILLER_20_341 ();
 sg13g2_fill_1 FILLER_20_343 ();
 sg13g2_fill_1 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_fill_2 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_198 ();
 sg13g2_fill_2 FILLER_21_250 ();
 sg13g2_fill_1 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_266 ();
 sg13g2_fill_1 FILLER_21_342 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_159 ();
 sg13g2_decap_4 FILLER_22_170 ();
 sg13g2_fill_1 FILLER_22_200 ();
 sg13g2_decap_4 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_fill_2 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_276 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_decap_4 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_4 FILLER_23_119 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_fill_2 FILLER_23_220 ();
 sg13g2_fill_1 FILLER_23_222 ();
 sg13g2_fill_1 FILLER_23_242 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_decap_4 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_146 ();
 sg13g2_decap_4 FILLER_24_166 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_decap_8 FILLER_24_184 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_fill_2 FILLER_24_269 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_310 ();
 sg13g2_decap_4 FILLER_24_316 ();
 sg13g2_fill_1 FILLER_24_328 ();
 sg13g2_fill_1 FILLER_24_348 ();
 sg13g2_decap_4 FILLER_24_358 ();
 sg13g2_decap_4 FILLER_24_388 ();
 sg13g2_fill_2 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_137 ();
 sg13g2_decap_4 FILLER_25_190 ();
 sg13g2_fill_1 FILLER_25_194 ();
 sg13g2_decap_8 FILLER_25_212 ();
 sg13g2_decap_4 FILLER_25_219 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_fill_2 FILLER_25_285 ();
 sg13g2_decap_4 FILLER_25_307 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_333 ();
 sg13g2_fill_2 FILLER_25_368 ();
 sg13g2_fill_2 FILLER_25_392 ();
 sg13g2_fill_1 FILLER_25_394 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_196 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_fill_2 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_decap_4 FILLER_26_285 ();
 sg13g2_fill_1 FILLER_26_294 ();
 sg13g2_decap_4 FILLER_26_299 ();
 sg13g2_decap_8 FILLER_26_318 ();
 sg13g2_fill_2 FILLER_26_325 ();
 sg13g2_fill_1 FILLER_26_327 ();
 sg13g2_decap_8 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_4 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_129 ();
 sg13g2_fill_1 FILLER_27_176 ();
 sg13g2_fill_2 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_fill_1 FILLER_27_211 ();
 sg13g2_fill_2 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_241 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_fill_2 FILLER_27_254 ();
 sg13g2_decap_8 FILLER_27_261 ();
 sg13g2_decap_4 FILLER_27_268 ();
 sg13g2_fill_1 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_286 ();
 sg13g2_decap_4 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_314 ();
 sg13g2_fill_2 FILLER_27_321 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_decap_8 FILLER_27_369 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_decap_4 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_146 ();
 sg13g2_decap_4 FILLER_28_155 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_216 ();
 sg13g2_decap_8 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_233 ();
 sg13g2_fill_2 FILLER_28_248 ();
 sg13g2_fill_1 FILLER_28_250 ();
 sg13g2_fill_1 FILLER_28_263 ();
 sg13g2_decap_4 FILLER_28_289 ();
 sg13g2_fill_2 FILLER_28_293 ();
 sg13g2_fill_2 FILLER_28_317 ();
 sg13g2_decap_8 FILLER_28_347 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_4 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_46 ();
 sg13g2_decap_8 FILLER_29_52 ();
 sg13g2_decap_8 FILLER_29_59 ();
 sg13g2_decap_8 FILLER_29_66 ();
 sg13g2_decap_8 FILLER_29_73 ();
 sg13g2_decap_8 FILLER_29_80 ();
 sg13g2_decap_8 FILLER_29_87 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_decap_8 FILLER_29_101 ();
 sg13g2_fill_1 FILLER_29_108 ();
 sg13g2_decap_8 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_fill_2 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_188 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_fill_2 FILLER_29_202 ();
 sg13g2_fill_1 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_263 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_fill_2 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_decap_4 FILLER_29_320 ();
 sg13g2_fill_2 FILLER_29_324 ();
 sg13g2_decap_4 FILLER_29_345 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_356 ();
 sg13g2_fill_1 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_59 ();
 sg13g2_decap_8 FILLER_30_66 ();
 sg13g2_decap_8 FILLER_30_73 ();
 sg13g2_decap_8 FILLER_30_80 ();
 sg13g2_fill_2 FILLER_30_87 ();
 sg13g2_fill_1 FILLER_30_119 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_204 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_fill_1 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_decap_8 FILLER_30_299 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_352 ();
 sg13g2_decap_4 FILLER_30_359 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_fill_1 FILLER_30_395 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_32 ();
 sg13g2_fill_2 FILLER_31_47 ();
 sg13g2_fill_1 FILLER_31_49 ();
 sg13g2_fill_2 FILLER_31_85 ();
 sg13g2_fill_2 FILLER_31_96 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_117 ();
 sg13g2_decap_8 FILLER_31_163 ();
 sg13g2_fill_2 FILLER_31_170 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_decap_4 FILLER_31_196 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_decap_8 FILLER_31_242 ();
 sg13g2_fill_2 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_251 ();
 sg13g2_decap_4 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_fill_2 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_319 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_decap_4 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_331 ();
 sg13g2_decap_8 FILLER_31_359 ();
 sg13g2_fill_1 FILLER_31_366 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_48 ();
 sg13g2_fill_1 FILLER_32_68 ();
 sg13g2_fill_2 FILLER_32_118 ();
 sg13g2_decap_4 FILLER_32_124 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_decap_8 FILLER_32_134 ();
 sg13g2_decap_4 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_fill_2 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_decap_8 FILLER_32_192 ();
 sg13g2_decap_4 FILLER_32_199 ();
 sg13g2_fill_2 FILLER_32_203 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_fill_2 FILLER_32_227 ();
 sg13g2_fill_1 FILLER_32_229 ();
 sg13g2_fill_2 FILLER_32_243 ();
 sg13g2_decap_4 FILLER_32_270 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_fill_1 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_fill_1 FILLER_32_384 ();
 sg13g2_fill_1 FILLER_32_393 ();
 sg13g2_fill_2 FILLER_32_398 ();
 sg13g2_fill_1 FILLER_33_31 ();
 sg13g2_fill_2 FILLER_33_50 ();
 sg13g2_fill_2 FILLER_33_78 ();
 sg13g2_fill_2 FILLER_33_87 ();
 sg13g2_decap_4 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_110 ();
 sg13g2_fill_1 FILLER_33_145 ();
 sg13g2_decap_4 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_decap_4 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_190 ();
 sg13g2_decap_4 FILLER_33_207 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_248 ();
 sg13g2_decap_8 FILLER_33_263 ();
 sg13g2_decap_4 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_fill_2 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_303 ();
 sg13g2_fill_2 FILLER_33_313 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_334 ();
 sg13g2_fill_2 FILLER_33_352 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_fill_2 FILLER_33_361 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_33_383 ();
 sg13g2_fill_1 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_33 ();
 sg13g2_decap_8 FILLER_34_52 ();
 sg13g2_fill_2 FILLER_34_67 ();
 sg13g2_fill_1 FILLER_34_69 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_decap_4 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_decap_4 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_210 ();
 sg13g2_decap_4 FILLER_34_226 ();
 sg13g2_fill_1 FILLER_34_238 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_267 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_decap_4 FILLER_34_342 ();
 sg13g2_fill_2 FILLER_34_346 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_368 ();
 sg13g2_fill_1 FILLER_34_376 ();
 sg13g2_fill_1 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_11 ();
 sg13g2_fill_2 FILLER_35_16 ();
 sg13g2_fill_1 FILLER_35_18 ();
 sg13g2_fill_1 FILLER_35_49 ();
 sg13g2_fill_1 FILLER_35_71 ();
 sg13g2_fill_1 FILLER_35_87 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_decap_4 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_127 ();
 sg13g2_decap_8 FILLER_35_142 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_decap_4 FILLER_35_199 ();
 sg13g2_fill_2 FILLER_35_245 ();
 sg13g2_decap_4 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_269 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_325 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_decap_8 FILLER_35_346 ();
 sg13g2_decap_4 FILLER_35_353 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_39 ();
 sg13g2_fill_2 FILLER_36_81 ();
 sg13g2_fill_1 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_135 ();
 sg13g2_fill_1 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_153 ();
 sg13g2_decap_8 FILLER_36_160 ();
 sg13g2_decap_8 FILLER_36_167 ();
 sg13g2_decap_4 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_178 ();
 sg13g2_fill_1 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_193 ();
 sg13g2_decap_4 FILLER_36_200 ();
 sg13g2_decap_4 FILLER_36_212 ();
 sg13g2_fill_2 FILLER_36_216 ();
 sg13g2_decap_8 FILLER_36_232 ();
 sg13g2_decap_4 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_243 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_321 ();
 sg13g2_fill_2 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_389 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_27 ();
 sg13g2_fill_2 FILLER_37_43 ();
 sg13g2_fill_1 FILLER_37_45 ();
 sg13g2_fill_1 FILLER_37_55 ();
 sg13g2_fill_1 FILLER_37_89 ();
 sg13g2_fill_2 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_174 ();
 sg13g2_fill_2 FILLER_37_179 ();
 sg13g2_decap_4 FILLER_37_217 ();
 sg13g2_fill_2 FILLER_37_221 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_fill_1 FILLER_37_269 ();
 sg13g2_fill_1 FILLER_37_291 ();
 sg13g2_fill_1 FILLER_37_332 ();
 sg13g2_fill_2 FILLER_37_342 ();
 sg13g2_fill_2 FILLER_37_360 ();
 sg13g2_fill_1 FILLER_37_362 ();
 sg13g2_fill_2 FILLER_37_397 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_101 ();
 sg13g2_fill_2 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_156 ();
 sg13g2_fill_1 FILLER_38_158 ();
 sg13g2_fill_1 FILLER_38_167 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_195 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_fill_1 FILLER_38_214 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_338 ();
 sg13g2_fill_1 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net17;
 assign uio_oe[5] = net18;
 assign uio_oe[6] = net19;
 assign uio_oe[7] = net20;
 assign uio_out[0] = net21;
 assign uio_out[1] = net22;
 assign uio_out[2] = net23;
 assign uio_out[3] = net24;
 assign uio_out[4] = net25;
 assign uio_out[5] = net26;
 assign uio_out[6] = net27;
 assign uio_out[7] = net28;
endmodule

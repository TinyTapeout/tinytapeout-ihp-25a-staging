module tt_um_wrapper (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire \dc4.clkcnt[0] ;
 wire \dc4.clkcnt[10] ;
 wire \dc4.clkcnt[11] ;
 wire \dc4.clkcnt[12] ;
 wire \dc4.clkcnt[13] ;
 wire \dc4.clkcnt[14] ;
 wire \dc4.clkcnt[1] ;
 wire \dc4.clkcnt[2] ;
 wire \dc4.clkcnt[3] ;
 wire \dc4.clkcnt[4] ;
 wire \dc4.clkcnt[5] ;
 wire \dc4.clkcnt[6] ;
 wire \dc4.clkcnt[7] ;
 wire \dc4.clkcnt[8] ;
 wire \dc4.clkcnt[9] ;
 wire \dc4.dot ;
 wire \dc4.ho[0] ;
 wire \dc4.ho[1] ;
 wire \dc4.ho[2] ;
 wire \dc4.ho[3] ;
 wire \dc4.ht[0] ;
 wire \dc4.ht[1] ;
 wire \dc4.ht[2] ;
 wire \dc4.ht[3] ;
 wire \dc4.mo[0] ;
 wire \dc4.mo[1] ;
 wire \dc4.mo[2] ;
 wire \dc4.mo[3] ;
 wire \dc4.mt[0] ;
 wire \dc4.mt[1] ;
 wire \dc4.mt[2] ;
 wire \dc4.mt[3] ;
 wire \dc4.pb_sreg[0][0] ;
 wire \dc4.pb_sreg[0][1] ;
 wire \dc4.pb_sreg[0][2] ;
 wire \dc4.pb_sreg[0][3] ;
 wire \dc4.pb_sreg[1][0] ;
 wire \dc4.pb_sreg[1][1] ;
 wire \dc4.pb_sreg[1][2] ;
 wire \dc4.pb_sreg[1][3] ;
 wire \dc4.sel[0] ;
 wire \dc4.sel[1] ;
 wire \dc4.sel[2] ;
 wire \dc4.so[0] ;
 wire \dc4.so[1] ;
 wire \dc4.so[2] ;
 wire \dc4.so[3] ;
 wire \dc4.st[0] ;
 wire \dc4.st[1] ;
 wire \dc4.st[2] ;
 wire \dc4.st[3] ;
 wire net4;
 wire clknet_0_clk;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;

 sg13g2_inv_1 _236_ (.Y(_046_),
    .A(net45));
 sg13g2_inv_2 _237_ (.Y(_047_),
    .A(net48));
 sg13g2_inv_1 _238_ (.Y(_048_),
    .A(\dc4.ho[2] ));
 sg13g2_inv_1 _239_ (.Y(_049_),
    .A(\dc4.ht[1] ));
 sg13g2_inv_1 _240_ (.Y(_050_),
    .A(net78));
 sg13g2_inv_1 _241_ (.Y(_051_),
    .A(net29));
 sg13g2_inv_1 _242_ (.Y(_052_),
    .A(net17));
 sg13g2_inv_1 _243_ (.Y(_053_),
    .A(net108));
 sg13g2_inv_1 _244_ (.Y(_054_),
    .A(net67));
 sg13g2_inv_1 _245_ (.Y(_055_),
    .A(net10));
 sg13g2_nor2b_1 _246_ (.A(net46),
    .B_N(net48),
    .Y(_056_));
 sg13g2_nand2b_1 _247_ (.Y(_057_),
    .B(net48),
    .A_N(net46));
 sg13g2_nor2_1 _248_ (.A(net44),
    .B(_057_),
    .Y(_058_));
 sg13g2_nor2b_1 _249_ (.A(\dc4.sel[2] ),
    .B_N(net46),
    .Y(_059_));
 sg13g2_nor2_1 _250_ (.A(net45),
    .B(\dc4.sel[0] ),
    .Y(_060_));
 sg13g2_and2_1 _251_ (.A(_047_),
    .B(_059_),
    .X(_061_));
 sg13g2_nor3_2 _252_ (.A(net45),
    .B(net46),
    .C(net48),
    .Y(_062_));
 sg13g2_nor2_1 _253_ (.A(net45),
    .B(_057_),
    .Y(_063_));
 sg13g2_a22oi_1 _254_ (.Y(_064_),
    .B1(_063_),
    .B2(\dc4.st[3] ),
    .A2(_062_),
    .A1(\dc4.so[3] ));
 sg13g2_and2_1 _255_ (.A(net48),
    .B(_059_),
    .X(_065_));
 sg13g2_nand3b_1 _256_ (.B(net47),
    .C(\dc4.sel[0] ),
    .Y(_066_),
    .A_N(net45));
 sg13g2_nor3_2 _257_ (.A(net46),
    .B(net48),
    .C(net44),
    .Y(_067_));
 sg13g2_a22oi_1 _258_ (.Y(_068_),
    .B1(_065_),
    .B2(\dc4.mt[3] ),
    .A2(_058_),
    .A1(\dc4.ht[3] ));
 sg13g2_a22oi_1 _259_ (.Y(_069_),
    .B1(_067_),
    .B2(\dc4.ho[3] ),
    .A2(_061_),
    .A1(\dc4.mo[3] ));
 sg13g2_and3_1 _260_ (.X(_070_),
    .A(_064_),
    .B(_068_),
    .C(_069_));
 sg13g2_nand2_1 _261_ (.Y(_071_),
    .A(net47),
    .B(_000_));
 sg13g2_a21oi_1 _262_ (.A1(net45),
    .A2(net44),
    .Y(_072_),
    .B1(net46));
 sg13g2_nor2b_1 _263_ (.A(_072_),
    .B_N(_071_),
    .Y(_073_));
 sg13g2_nand2b_1 _264_ (.Y(_074_),
    .B(_071_),
    .A_N(_072_));
 sg13g2_a22oi_1 _265_ (.Y(_075_),
    .B1(_063_),
    .B2(\dc4.st[1] ),
    .A2(_062_),
    .A1(\dc4.so[1] ));
 sg13g2_nor3_1 _266_ (.A(net44),
    .B(_049_),
    .C(_057_),
    .Y(_076_));
 sg13g2_nor2_1 _267_ (.A(_050_),
    .B(_066_),
    .Y(_077_));
 sg13g2_and2_1 _268_ (.A(\dc4.ho[1] ),
    .B(_067_),
    .X(_078_));
 sg13g2_and3_1 _269_ (.X(_079_),
    .A(net47),
    .B(\dc4.mo[1] ),
    .C(_060_));
 sg13g2_nor4_1 _270_ (.A(_076_),
    .B(_077_),
    .C(_078_),
    .D(_079_),
    .Y(_080_));
 sg13g2_a21o_2 _271_ (.A2(_080_),
    .A1(_075_),
    .B1(_073_),
    .X(_081_));
 sg13g2_nand2_1 _272_ (.Y(_082_),
    .A(\dc4.ho[2] ),
    .B(_067_));
 sg13g2_nand2_1 _273_ (.Y(_083_),
    .A(\dc4.so[2] ),
    .B(_062_));
 sg13g2_or3_1 _274_ (.A(net44),
    .B(_001_),
    .C(_057_),
    .X(_084_));
 sg13g2_nand3_1 _275_ (.B(\dc4.st[2] ),
    .C(_056_),
    .A(_046_),
    .Y(_085_));
 sg13g2_nand3_1 _276_ (.B(\dc4.mo[2] ),
    .C(_060_),
    .A(net47),
    .Y(_086_));
 sg13g2_o21ai_1 _277_ (.B1(_082_),
    .Y(_087_),
    .A1(_051_),
    .A2(_066_));
 sg13g2_nand4_1 _278_ (.B(_084_),
    .C(_085_),
    .A(_083_),
    .Y(_088_),
    .D(_086_));
 sg13g2_or2_1 _279_ (.X(_089_),
    .B(_088_),
    .A(_087_));
 sg13g2_inv_1 _280_ (.Y(_090_),
    .A(_089_));
 sg13g2_o21ai_1 _281_ (.B1(_074_),
    .Y(_091_),
    .A1(_087_),
    .A2(_088_));
 sg13g2_nand2_1 _282_ (.Y(_092_),
    .A(_081_),
    .B(_091_));
 sg13g2_a21oi_2 _283_ (.B1(_070_),
    .Y(_093_),
    .A2(_091_),
    .A1(_081_));
 sg13g2_nand2b_1 _284_ (.Y(_094_),
    .B(_074_),
    .A_N(_070_));
 sg13g2_nand2_1 _285_ (.Y(_095_),
    .A(\dc4.ho[0] ),
    .B(_067_));
 sg13g2_nand3_1 _286_ (.B(\dc4.mt[0] ),
    .C(_059_),
    .A(\dc4.sel[0] ),
    .Y(_096_));
 sg13g2_nand2_1 _287_ (.Y(_097_),
    .A(\dc4.so[0] ),
    .B(_062_));
 sg13g2_nand3_1 _288_ (.B(\dc4.st[0] ),
    .C(_056_),
    .A(_046_),
    .Y(_098_));
 sg13g2_a22oi_1 _289_ (.Y(_099_),
    .B1(_061_),
    .B2(\dc4.mo[0] ),
    .A2(_058_),
    .A1(_055_));
 sg13g2_and4_1 _290_ (.A(_095_),
    .B(_096_),
    .C(_097_),
    .D(_098_),
    .X(_100_));
 sg13g2_and2_1 _291_ (.A(_099_),
    .B(_100_),
    .X(_101_));
 sg13g2_a21oi_1 _292_ (.A1(_099_),
    .A2(_100_),
    .Y(_102_),
    .B1(_073_));
 sg13g2_or2_1 _293_ (.X(_103_),
    .B(_101_),
    .A(_081_));
 sg13g2_o21ai_1 _294_ (.B1(_092_),
    .Y(_104_),
    .A1(_090_),
    .A2(_103_));
 sg13g2_a21o_1 _295_ (.A2(_104_),
    .A1(_094_),
    .B1(_093_),
    .X(uo_out[0]));
 sg13g2_nand2_1 _296_ (.Y(_105_),
    .A(_089_),
    .B(_103_));
 sg13g2_o21ai_1 _297_ (.B1(_081_),
    .Y(_106_),
    .A1(_073_),
    .A2(_101_));
 sg13g2_inv_1 _298_ (.Y(_107_),
    .A(_106_));
 sg13g2_and2_1 _299_ (.A(_094_),
    .B(_106_),
    .X(_108_));
 sg13g2_a21o_1 _300_ (.A2(_108_),
    .A1(_105_),
    .B1(_093_),
    .X(uo_out[1]));
 sg13g2_nor2b_1 _301_ (.A(_081_),
    .B_N(_101_),
    .Y(_109_));
 sg13g2_a22oi_1 _302_ (.Y(uo_out[2]),
    .B1(_109_),
    .B2(_070_),
    .A2(_107_),
    .A1(_091_));
 sg13g2_mux2_1 _303_ (.A0(_101_),
    .A1(_102_),
    .S(_081_),
    .X(_110_));
 sg13g2_nand3_1 _304_ (.B(_091_),
    .C(_102_),
    .A(_081_),
    .Y(_111_));
 sg13g2_o21ai_1 _305_ (.B1(_111_),
    .Y(_112_),
    .A1(_091_),
    .A2(_110_));
 sg13g2_a21o_1 _306_ (.A2(_112_),
    .A1(_094_),
    .B1(_093_),
    .X(uo_out[3]));
 sg13g2_a21o_1 _307_ (.A2(_109_),
    .A1(_090_),
    .B1(_093_),
    .X(uo_out[4]));
 sg13g2_nand2b_1 _308_ (.Y(_113_),
    .B(_110_),
    .A_N(_091_));
 sg13g2_nand2b_1 _309_ (.Y(uo_out[5]),
    .B(_113_),
    .A_N(_093_));
 sg13g2_o21ai_1 _310_ (.B1(_111_),
    .Y(_114_),
    .A1(_091_),
    .A2(_106_));
 sg13g2_a21o_1 _311_ (.A2(_114_),
    .A1(_094_),
    .B1(_093_),
    .X(uo_out[6]));
 sg13g2_nand2_1 _312_ (.Y(uio_out[0]),
    .A(_000_),
    .B(_062_));
 sg13g2_nand2_1 _313_ (.Y(uio_out[1]),
    .A(_000_),
    .B(_063_));
 sg13g2_nand2b_1 _314_ (.Y(uio_out[2]),
    .B(_047_),
    .A_N(_071_));
 sg13g2_nand3_1 _315_ (.B(net48),
    .C(net44),
    .A(net46),
    .Y(uio_out[3]));
 sg13g2_nand2_2 _316_ (.Y(uio_out[4]),
    .A(net45),
    .B(_067_));
 sg13g2_nand2_2 _317_ (.Y(uio_out[5]),
    .A(net45),
    .B(_058_));
 sg13g2_nand2b_1 _318_ (.Y(_115_),
    .B(\dc4.clkcnt[14] ),
    .A_N(_067_));
 sg13g2_o21ai_1 _319_ (.B1(_115_),
    .Y(\dc4.dot ),
    .A1(\dc4.clkcnt[14] ),
    .A2(_061_));
 sg13g2_nand3_1 _320_ (.B(net40),
    .C(net100),
    .A(\dc4.clkcnt[0] ),
    .Y(_116_));
 sg13g2_and4_1 _321_ (.A(\dc4.clkcnt[0] ),
    .B(\dc4.clkcnt[1] ),
    .C(net19),
    .D(\dc4.clkcnt[2] ),
    .X(_117_));
 sg13g2_and2_1 _322_ (.A(net32),
    .B(_117_),
    .X(_118_));
 sg13g2_and2_2 _323_ (.A(net69),
    .B(_118_),
    .X(_119_));
 sg13g2_nand2_2 _324_ (.Y(_120_),
    .A(net69),
    .B(_118_));
 sg13g2_nand4_1 _325_ (.B(net32),
    .C(net15),
    .A(\dc4.clkcnt[5] ),
    .Y(_121_),
    .D(_117_));
 sg13g2_nor3_1 _326_ (.A(_052_),
    .B(_053_),
    .C(_121_),
    .Y(_122_));
 sg13g2_nor4_2 _327_ (.A(_052_),
    .B(_053_),
    .C(_054_),
    .Y(_123_),
    .D(_121_));
 sg13g2_and3_2 _328_ (.X(_124_),
    .A(net12),
    .B(net34),
    .C(_123_));
 sg13g2_a21oi_1 _329_ (.A1(\dc4.clkcnt[12] ),
    .A2(_124_),
    .Y(_125_),
    .B1(net23));
 sg13g2_and3_1 _330_ (.X(_126_),
    .A(net23),
    .B(net58),
    .C(_124_));
 sg13g2_nor2_1 _331_ (.A(net24),
    .B(_126_),
    .Y(_006_));
 sg13g2_and3_1 _332_ (.X(_127_),
    .A(net23),
    .B(\dc4.clkcnt[12] ),
    .C(\dc4.clkcnt[14] ));
 sg13g2_nand2_1 _333_ (.Y(_128_),
    .A(_124_),
    .B(_127_));
 sg13g2_o21ai_1 _334_ (.B1(_128_),
    .Y(_129_),
    .A1(net95),
    .A2(_126_));
 sg13g2_inv_1 _335_ (.Y(_007_),
    .A(_129_));
 sg13g2_xor2_1 _336_ (.B(net40),
    .A(\dc4.clkcnt[0] ),
    .X(_008_));
 sg13g2_a21o_1 _337_ (.A2(net40),
    .A1(\dc4.clkcnt[0] ),
    .B1(net100),
    .X(_130_));
 sg13g2_and2_1 _338_ (.A(_116_),
    .B(net101),
    .X(_009_));
 sg13g2_xnor2_1 _339_ (.Y(_010_),
    .A(net19),
    .B(_116_));
 sg13g2_xor2_1 _340_ (.B(_117_),
    .A(net32),
    .X(_011_));
 sg13g2_xor2_1 _341_ (.B(_118_),
    .A(net69),
    .X(_012_));
 sg13g2_xnor2_1 _342_ (.Y(_013_),
    .A(net15),
    .B(_120_));
 sg13g2_xnor2_1 _343_ (.Y(_014_),
    .A(net17),
    .B(_121_));
 sg13g2_o21ai_1 _344_ (.B1(_053_),
    .Y(_131_),
    .A1(_052_),
    .A2(_121_));
 sg13g2_nor2b_1 _345_ (.A(_122_),
    .B_N(net109),
    .Y(_015_));
 sg13g2_xnor2_1 _346_ (.Y(_016_),
    .A(_054_),
    .B(_122_));
 sg13g2_xor2_1 _347_ (.B(_123_),
    .A(net34),
    .X(_003_));
 sg13g2_a21oi_1 _348_ (.A1(\dc4.clkcnt[10] ),
    .A2(_123_),
    .Y(_132_),
    .B1(net12));
 sg13g2_nor2_1 _349_ (.A(_124_),
    .B(net13),
    .Y(_004_));
 sg13g2_xor2_1 _350_ (.B(_124_),
    .A(net58),
    .X(_005_));
 sg13g2_nand3_1 _351_ (.B(_124_),
    .C(_127_),
    .A(\dc4.so[0] ),
    .Y(_133_));
 sg13g2_nand2_1 _352_ (.Y(_134_),
    .A(net70),
    .B(net59));
 sg13g2_nor3_2 _353_ (.A(net99),
    .B(net81),
    .C(_134_),
    .Y(_135_));
 sg13g2_xor2_1 _354_ (.B(_128_),
    .A(net99),
    .X(_136_));
 sg13g2_nor2_1 _355_ (.A(_135_),
    .B(_136_),
    .Y(_017_));
 sg13g2_nor2b_1 _356_ (.A(net70),
    .B_N(_133_),
    .Y(_137_));
 sg13g2_and4_1 _357_ (.A(net70),
    .B(\dc4.so[0] ),
    .C(_124_),
    .D(_127_),
    .X(_138_));
 sg13g2_nor3_1 _358_ (.A(_135_),
    .B(net71),
    .C(_138_),
    .Y(_018_));
 sg13g2_xor2_1 _359_ (.B(_138_),
    .A(net81),
    .X(_019_));
 sg13g2_a21oi_1 _360_ (.A1(\dc4.so[2] ),
    .A2(_138_),
    .Y(_139_),
    .B1(net59));
 sg13g2_and3_1 _361_ (.X(_140_),
    .A(\dc4.so[2] ),
    .B(net59),
    .C(_138_));
 sg13g2_nor3_1 _362_ (.A(_135_),
    .B(net60),
    .C(_140_),
    .Y(_020_));
 sg13g2_nand2_1 _363_ (.Y(_141_),
    .A(net75),
    .B(net42));
 sg13g2_nor3_2 _364_ (.A(net88),
    .B(net65),
    .C(_141_),
    .Y(_142_));
 sg13g2_nor2b_1 _365_ (.A(net105),
    .B_N(net8),
    .Y(_143_));
 sg13g2_nor2_1 _366_ (.A(_142_),
    .B(_143_),
    .Y(_144_));
 sg13g2_nor3_1 _367_ (.A(\dc4.mo[0] ),
    .B(_142_),
    .C(_143_),
    .Y(_145_));
 sg13g2_nand2_1 _368_ (.Y(_146_),
    .A(net92),
    .B(net83));
 sg13g2_nor3_2 _369_ (.A(\dc4.mo[0] ),
    .B(net62),
    .C(_146_),
    .Y(_147_));
 sg13g2_nor2b_2 _370_ (.A(_144_),
    .B_N(\dc4.mo[0] ),
    .Y(_148_));
 sg13g2_nor3_1 _371_ (.A(net106),
    .B(_147_),
    .C(_148_),
    .Y(_021_));
 sg13g2_xnor2_1 _372_ (.Y(_149_),
    .A(net92),
    .B(_148_));
 sg13g2_nor2_1 _373_ (.A(_147_),
    .B(net93),
    .Y(_022_));
 sg13g2_a21oi_1 _374_ (.A1(\dc4.mo[1] ),
    .A2(_148_),
    .Y(_150_),
    .B1(net62));
 sg13g2_nand3_1 _375_ (.B(net62),
    .C(_148_),
    .A(\dc4.mo[1] ),
    .Y(_151_));
 sg13g2_nor2b_1 _376_ (.A(net63),
    .B_N(_151_),
    .Y(_023_));
 sg13g2_xor2_1 _377_ (.B(_151_),
    .A(net83),
    .X(_152_));
 sg13g2_nor2_1 _378_ (.A(_147_),
    .B(net84),
    .Y(_024_));
 sg13g2_nand2_1 _379_ (.Y(_153_),
    .A(\dc4.ho[1] ),
    .B(\dc4.ho[3] ));
 sg13g2_nor3_2 _380_ (.A(\dc4.ho[0] ),
    .B(\dc4.ho[2] ),
    .C(_153_),
    .Y(_154_));
 sg13g2_nor4_1 _381_ (.A(_049_),
    .B(\dc4.ht[0] ),
    .C(\dc4.ht[3] ),
    .D(\dc4.ht[2] ),
    .Y(_155_));
 sg13g2_nor4_1 _382_ (.A(\dc4.ho[1] ),
    .B(\dc4.ho[0] ),
    .C(_048_),
    .D(\dc4.ho[3] ),
    .Y(_156_));
 sg13g2_and2_1 _383_ (.A(_155_),
    .B(_156_),
    .X(_157_));
 sg13g2_or2_1 _384_ (.X(_158_),
    .B(_157_),
    .A(_154_));
 sg13g2_nor4_2 _385_ (.A(_050_),
    .B(net86),
    .C(net73),
    .Y(_159_),
    .D(_051_));
 sg13g2_nand2b_1 _386_ (.Y(_160_),
    .B(\dc4.pb_sreg[1][2] ),
    .A_N(\dc4.pb_sreg[1][3] ));
 sg13g2_nand2b_2 _387_ (.Y(_161_),
    .B(_160_),
    .A_N(_159_));
 sg13g2_nor2_1 _388_ (.A(_158_),
    .B(_161_),
    .Y(_162_));
 sg13g2_nor2b_1 _389_ (.A(_158_),
    .B_N(_161_),
    .Y(_163_));
 sg13g2_mux2_1 _390_ (.A0(_163_),
    .A1(_162_),
    .S(net111),
    .X(_025_));
 sg13g2_xor2_1 _391_ (.B(\dc4.ho[0] ),
    .A(net97),
    .X(_164_));
 sg13g2_a22oi_1 _392_ (.Y(_165_),
    .B1(_163_),
    .B2(_164_),
    .A2(_162_),
    .A1(net97));
 sg13g2_inv_1 _393_ (.Y(_026_),
    .A(net98));
 sg13g2_nand3_1 _394_ (.B(\dc4.ho[0] ),
    .C(_161_),
    .A(net97),
    .Y(_166_));
 sg13g2_nand4_1 _395_ (.B(\dc4.ho[0] ),
    .C(\dc4.ho[2] ),
    .A(\dc4.ho[1] ),
    .Y(_167_),
    .D(_161_));
 sg13g2_xor2_1 _396_ (.B(_166_),
    .A(net103),
    .X(_168_));
 sg13g2_nor2_1 _397_ (.A(_158_),
    .B(net104),
    .Y(_027_));
 sg13g2_xor2_1 _398_ (.B(_167_),
    .A(net90),
    .X(_169_));
 sg13g2_nor2_1 _399_ (.A(_158_),
    .B(net91),
    .Y(_028_));
 sg13g2_nor2_1 _400_ (.A(\dc4.ht[0] ),
    .B(_154_),
    .Y(_170_));
 sg13g2_a21oi_1 _401_ (.A1(_055_),
    .A2(_154_),
    .Y(_029_),
    .B1(_170_));
 sg13g2_a21oi_1 _402_ (.A1(\dc4.ht[0] ),
    .A2(_154_),
    .Y(_171_),
    .B1(net26));
 sg13g2_nand3_1 _403_ (.B(\dc4.ht[0] ),
    .C(_154_),
    .A(net26),
    .Y(_172_));
 sg13g2_nand2b_1 _404_ (.Y(_173_),
    .B(_172_),
    .A_N(_157_));
 sg13g2_nor2_1 _405_ (.A(net27),
    .B(_173_),
    .Y(_030_));
 sg13g2_xnor2_1 _406_ (.Y(_031_),
    .A(net21),
    .B(_172_));
 sg13g2_nor2_1 _407_ (.A(_001_),
    .B(_172_),
    .Y(_174_));
 sg13g2_xor2_1 _408_ (.B(_174_),
    .A(net38),
    .X(_032_));
 sg13g2_xnor2_1 _409_ (.Y(_033_),
    .A(_047_),
    .B(_119_));
 sg13g2_o21ai_1 _410_ (.B1(net46),
    .Y(_175_),
    .A1(_047_),
    .A2(_120_));
 sg13g2_nand3_1 _411_ (.B(_056_),
    .C(_119_),
    .A(net44),
    .Y(_176_));
 sg13g2_nand2_1 _412_ (.Y(_034_),
    .A(_175_),
    .B(_176_));
 sg13g2_o21ai_1 _413_ (.B1(uio_out[3]),
    .Y(_177_),
    .A1(net48),
    .A2(net44));
 sg13g2_nor2_1 _414_ (.A(_120_),
    .B(_177_),
    .Y(_178_));
 sg13g2_a21oi_1 _415_ (.A1(_046_),
    .A2(_120_),
    .Y(_035_),
    .B1(_178_));
 sg13g2_nor2_1 _416_ (.A(net88),
    .B(_135_),
    .Y(_179_));
 sg13g2_and2_1 _417_ (.A(net88),
    .B(_135_),
    .X(_180_));
 sg13g2_nor3_1 _418_ (.A(_142_),
    .B(net89),
    .C(_180_),
    .Y(_036_));
 sg13g2_xnor2_1 _419_ (.Y(_181_),
    .A(net75),
    .B(_180_));
 sg13g2_nor2_1 _420_ (.A(_142_),
    .B(net76),
    .Y(_037_));
 sg13g2_a21oi_1 _421_ (.A1(\dc4.st[1] ),
    .A2(_180_),
    .Y(_182_),
    .B1(net42));
 sg13g2_nor2b_1 _422_ (.A(_141_),
    .B_N(_180_),
    .Y(_183_));
 sg13g2_nor3_1 _423_ (.A(_142_),
    .B(net43),
    .C(_183_),
    .Y(_038_));
 sg13g2_xor2_1 _424_ (.B(_183_),
    .A(net65),
    .X(_039_));
 sg13g2_mux2_1 _425_ (.A0(net8),
    .A1(net36),
    .S(_119_),
    .X(_040_));
 sg13g2_mux2_1 _426_ (.A0(net9),
    .A1(net37),
    .S(_119_),
    .X(_041_));
 sg13g2_nor2_1 _427_ (.A(net86),
    .B(_147_),
    .Y(_184_));
 sg13g2_and2_1 _428_ (.A(net86),
    .B(_147_),
    .X(_185_));
 sg13g2_nor3_1 _429_ (.A(_159_),
    .B(net87),
    .C(_185_),
    .Y(_042_));
 sg13g2_xnor2_1 _430_ (.Y(_186_),
    .A(net78),
    .B(_185_));
 sg13g2_nor2_1 _431_ (.A(_159_),
    .B(net79),
    .Y(_043_));
 sg13g2_a21oi_1 _432_ (.A1(\dc4.mt[1] ),
    .A2(_185_),
    .Y(_187_),
    .B1(net29));
 sg13g2_and3_1 _433_ (.X(_188_),
    .A(\dc4.mt[1] ),
    .B(net29),
    .C(_185_));
 sg13g2_nor3_1 _434_ (.A(_159_),
    .B(net30),
    .C(_188_),
    .Y(_044_));
 sg13g2_xor2_1 _435_ (.B(_188_),
    .A(net73),
    .X(_045_));
 sg13g2_dfrbp_1 _436_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net54),
    .D(net2),
    .Q_N(_217_),
    .Q(\dc4.pb_sreg[1][0] ));
 sg13g2_dfrbp_1 _437_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net54),
    .D(net7),
    .Q_N(_218_),
    .Q(\dc4.pb_sreg[1][1] ));
 sg13g2_dfrbp_1 _438_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net56),
    .D(net9),
    .Q_N(_219_),
    .Q(\dc4.pb_sreg[1][3] ));
 sg13g2_dfrbp_1 _439_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net54),
    .D(net1),
    .Q_N(_220_),
    .Q(\dc4.pb_sreg[0][0] ));
 sg13g2_dfrbp_1 _440_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net54),
    .D(net6),
    .Q_N(_221_),
    .Q(\dc4.pb_sreg[0][1] ));
 sg13g2_dfrbp_1 _441_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net54),
    .D(net8),
    .Q_N(_216_),
    .Q(\dc4.pb_sreg[0][3] ));
 sg13g2_dfrbp_1 _442_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net49),
    .D(_017_),
    .Q_N(_215_),
    .Q(\dc4.so[0] ));
 sg13g2_dfrbp_1 _443_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net49),
    .D(net72),
    .Q_N(_214_),
    .Q(\dc4.so[1] ));
 sg13g2_dfrbp_1 _444_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net49),
    .D(net82),
    .Q_N(_213_),
    .Q(\dc4.so[2] ));
 sg13g2_dfrbp_1 _445_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net51),
    .D(net61),
    .Q_N(_212_),
    .Q(\dc4.so[3] ));
 sg13g2_dfrbp_1 _446_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net53),
    .D(net107),
    .Q_N(_211_),
    .Q(\dc4.mo[0] ));
 sg13g2_dfrbp_1 _447_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net52),
    .D(net94),
    .Q_N(_210_),
    .Q(\dc4.mo[1] ));
 sg13g2_dfrbp_1 _448_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net52),
    .D(net64),
    .Q_N(_209_),
    .Q(\dc4.mo[2] ));
 sg13g2_dfrbp_1 _449_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net53),
    .D(net85),
    .Q_N(_208_),
    .Q(\dc4.mo[3] ));
 sg13g2_dfrbp_1 _450_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net52),
    .D(_025_),
    .Q_N(_207_),
    .Q(\dc4.ho[0] ));
 sg13g2_dfrbp_1 _451_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net51),
    .D(_026_),
    .Q_N(_206_),
    .Q(\dc4.ho[1] ));
 sg13g2_dfrbp_1 _452_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net52),
    .D(_027_),
    .Q_N(_205_),
    .Q(\dc4.ho[2] ));
 sg13g2_dfrbp_1 _453_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net52),
    .D(_028_),
    .Q_N(_204_),
    .Q(\dc4.ho[3] ));
 sg13g2_dfrbp_1 _454_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net51),
    .D(net11),
    .Q_N(_002_),
    .Q(\dc4.ht[0] ));
 sg13g2_dfrbp_1 _455_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net51),
    .D(net28),
    .Q_N(_203_),
    .Q(\dc4.ht[1] ));
 sg13g2_dfrbp_1 _456_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net51),
    .D(net22),
    .Q_N(_001_),
    .Q(\dc4.ht[2] ));
 sg13g2_dfrbp_1 _457_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net51),
    .D(net39),
    .Q_N(_202_),
    .Q(\dc4.ht[3] ));
 sg13g2_dfrbp_1 _458_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net50),
    .D(_033_),
    .Q_N(_201_),
    .Q(\dc4.sel[0] ));
 sg13g2_dfrbp_1 _459_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net49),
    .D(_034_),
    .Q_N(_200_),
    .Q(\dc4.sel[1] ));
 sg13g2_dfrbp_1 _460_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net50),
    .D(_035_),
    .Q_N(_000_),
    .Q(\dc4.sel[2] ));
 sg13g2_dfrbp_1 _461_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net50),
    .D(_036_),
    .Q_N(_199_),
    .Q(\dc4.st[0] ));
 sg13g2_dfrbp_1 _462_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net50),
    .D(net77),
    .Q_N(_198_),
    .Q(\dc4.st[1] ));
 sg13g2_dfrbp_1 _463_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net50),
    .D(net57),
    .Q_N(_197_),
    .Q(\dc4.st[2] ));
 sg13g2_dfrbp_1 _464_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net50),
    .D(net66),
    .Q_N(_196_),
    .Q(\dc4.st[3] ));
 sg13g2_dfrbp_1 _465_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net54),
    .D(_040_),
    .Q_N(_195_),
    .Q(\dc4.pb_sreg[0][2] ));
 sg13g2_dfrbp_1 _466_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net54),
    .D(_041_),
    .Q_N(_194_),
    .Q(\dc4.pb_sreg[1][2] ));
 sg13g2_dfrbp_1 _467_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net53),
    .D(_042_),
    .Q_N(_193_),
    .Q(\dc4.mt[0] ));
 sg13g2_dfrbp_1 _468_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net53),
    .D(net80),
    .Q_N(_192_),
    .Q(\dc4.mt[1] ));
 sg13g2_dfrbp_1 _469_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net52),
    .D(net31),
    .Q_N(_191_),
    .Q(\dc4.mt[2] ));
 sg13g2_dfrbp_1 _470_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net53),
    .D(net74),
    .Q_N(_222_),
    .Q(\dc4.mt[3] ));
 sg13g2_dfrbp_1 _471_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net55),
    .D(net5),
    .Q_N(_189_),
    .Q(\dc4.clkcnt[0] ));
 sg13g2_dfrbp_1 _472_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net55),
    .D(net41),
    .Q_N(_223_),
    .Q(\dc4.clkcnt[1] ));
 sg13g2_dfrbp_1 _473_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net55),
    .D(net102),
    .Q_N(_224_),
    .Q(\dc4.clkcnt[2] ));
 sg13g2_dfrbp_1 _474_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net55),
    .D(net20),
    .Q_N(_225_),
    .Q(\dc4.clkcnt[3] ));
 sg13g2_dfrbp_1 _475_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net55),
    .D(net33),
    .Q_N(_226_),
    .Q(\dc4.clkcnt[4] ));
 sg13g2_dfrbp_1 _476_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net54),
    .D(_012_),
    .Q_N(_227_),
    .Q(\dc4.clkcnt[5] ));
 sg13g2_dfrbp_1 _477_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net55),
    .D(net16),
    .Q_N(_228_),
    .Q(\dc4.clkcnt[6] ));
 sg13g2_dfrbp_1 _478_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net52),
    .D(net18),
    .Q_N(_229_),
    .Q(\dc4.clkcnt[7] ));
 sg13g2_dfrbp_1 _479_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net55),
    .D(net110),
    .Q_N(_230_),
    .Q(\dc4.clkcnt[8] ));
 sg13g2_dfrbp_1 _480_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net52),
    .D(net68),
    .Q_N(_231_),
    .Q(\dc4.clkcnt[9] ));
 sg13g2_dfrbp_1 _481_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net49),
    .D(net35),
    .Q_N(_232_),
    .Q(\dc4.clkcnt[10] ));
 sg13g2_dfrbp_1 _482_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net49),
    .D(net14),
    .Q_N(_233_),
    .Q(\dc4.clkcnt[11] ));
 sg13g2_dfrbp_1 _483_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net49),
    .D(_005_),
    .Q_N(_234_),
    .Q(\dc4.clkcnt[12] ));
 sg13g2_dfrbp_1 _484_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net49),
    .D(net25),
    .Q_N(_235_),
    .Q(\dc4.clkcnt[13] ));
 sg13g2_dfrbp_1 _485_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net50),
    .D(_007_),
    .Q_N(_190_),
    .Q(\dc4.clkcnt[14] ));
 sg13g2_tielo tt_um_wrapper_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _488_ (.A(ena),
    .X(uio_oe[0]));
 sg13g2_buf_1 _489_ (.A(ena),
    .X(uio_oe[1]));
 sg13g2_buf_1 _490_ (.A(ena),
    .X(uio_oe[2]));
 sg13g2_buf_1 _491_ (.A(ena),
    .X(uio_oe[3]));
 sg13g2_buf_1 _492_ (.A(ena),
    .X(uio_oe[4]));
 sg13g2_buf_1 _493_ (.A(ena),
    .X(uio_oe[5]));
 sg13g2_buf_1 _494_ (.A(ena),
    .X(uio_oe[6]));
 sg13g2_buf_1 _495_ (.A(ena),
    .X(uio_oe[7]));
 sg13g2_buf_1 _496_ (.A(\dc4.dot ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout44 (.A(net112),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(net96),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_1 fanout47 (.A(\dc4.sel[1] ),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(\dc4.sel[0] ),
    .X(net48));
 sg13g2_buf_4 fanout49 (.X(net49),
    .A(net50));
 sg13g2_buf_4 fanout50 (.X(net50),
    .A(net51));
 sg13g2_buf_4 fanout51 (.X(net51),
    .A(rst_n));
 sg13g2_buf_4 fanout52 (.X(net52),
    .A(net56));
 sg13g2_buf_4 fanout53 (.X(net53),
    .A(net56));
 sg13g2_buf_4 fanout54 (.X(net54),
    .A(net55));
 sg13g2_buf_4 fanout55 (.X(net55),
    .A(net56));
 sg13g2_buf_2 fanout56 (.A(rst_n),
    .X(net56));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_wrapper_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_189_),
    .X(net5));
 sg13g2_dlygate4sd3_1 hold2 (.A(\dc4.pb_sreg[0][0] ),
    .X(net6));
 sg13g2_dlygate4sd3_1 hold3 (.A(\dc4.pb_sreg[1][0] ),
    .X(net7));
 sg13g2_dlygate4sd3_1 hold4 (.A(\dc4.pb_sreg[0][2] ),
    .X(net8));
 sg13g2_dlygate4sd3_1 hold5 (.A(\dc4.pb_sreg[1][2] ),
    .X(net9));
 sg13g2_dlygate4sd3_1 hold6 (.A(_002_),
    .X(net10));
 sg13g2_dlygate4sd3_1 hold7 (.A(_029_),
    .X(net11));
 sg13g2_dlygate4sd3_1 hold8 (.A(\dc4.clkcnt[11] ),
    .X(net12));
 sg13g2_dlygate4sd3_1 hold9 (.A(_132_),
    .X(net13));
 sg13g2_dlygate4sd3_1 hold10 (.A(_004_),
    .X(net14));
 sg13g2_dlygate4sd3_1 hold11 (.A(\dc4.clkcnt[6] ),
    .X(net15));
 sg13g2_dlygate4sd3_1 hold12 (.A(_013_),
    .X(net16));
 sg13g2_dlygate4sd3_1 hold13 (.A(\dc4.clkcnt[7] ),
    .X(net17));
 sg13g2_dlygate4sd3_1 hold14 (.A(_014_),
    .X(net18));
 sg13g2_dlygate4sd3_1 hold15 (.A(\dc4.clkcnt[3] ),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold16 (.A(_010_),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold17 (.A(\dc4.ht[2] ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold18 (.A(_031_),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold19 (.A(\dc4.clkcnt[13] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold20 (.A(_125_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold21 (.A(_006_),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold22 (.A(\dc4.ht[1] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold23 (.A(_171_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold24 (.A(_030_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold25 (.A(\dc4.mt[2] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold26 (.A(_187_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold27 (.A(_044_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold28 (.A(\dc4.clkcnt[4] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold29 (.A(_011_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold30 (.A(\dc4.clkcnt[10] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold31 (.A(_003_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold32 (.A(\dc4.pb_sreg[0][1] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold33 (.A(\dc4.pb_sreg[1][1] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold34 (.A(\dc4.ht[3] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold35 (.A(_032_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold36 (.A(\dc4.clkcnt[1] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold37 (.A(_008_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold38 (.A(\dc4.st[2] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold39 (.A(_182_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold40 (.A(_038_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold41 (.A(\dc4.clkcnt[12] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold42 (.A(\dc4.so[3] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold43 (.A(_139_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold44 (.A(_020_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold45 (.A(\dc4.mo[2] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold46 (.A(_150_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold47 (.A(_023_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold48 (.A(\dc4.st[3] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold49 (.A(_039_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold50 (.A(\dc4.clkcnt[9] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold51 (.A(_016_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold52 (.A(\dc4.clkcnt[5] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold53 (.A(\dc4.so[1] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold54 (.A(_137_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold55 (.A(_018_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold56 (.A(\dc4.mt[3] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold57 (.A(_045_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold58 (.A(\dc4.st[1] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold59 (.A(_181_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold60 (.A(_037_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold61 (.A(\dc4.mt[1] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold62 (.A(_186_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold63 (.A(_043_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold64 (.A(\dc4.so[2] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold65 (.A(_019_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold66 (.A(\dc4.mo[3] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold67 (.A(_152_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold68 (.A(_024_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold69 (.A(\dc4.mt[0] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold70 (.A(_184_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold71 (.A(\dc4.st[0] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold72 (.A(_179_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold73 (.A(\dc4.ho[3] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold74 (.A(_169_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold75 (.A(\dc4.mo[1] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold76 (.A(_149_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold77 (.A(_022_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold78 (.A(\dc4.clkcnt[14] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold79 (.A(\dc4.sel[2] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold80 (.A(\dc4.ho[1] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold81 (.A(_165_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold82 (.A(\dc4.so[0] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold83 (.A(\dc4.clkcnt[2] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold84 (.A(_130_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold85 (.A(_009_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold86 (.A(\dc4.ho[2] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold87 (.A(_168_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold88 (.A(\dc4.pb_sreg[0][3] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold89 (.A(_145_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold90 (.A(_021_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold91 (.A(\dc4.clkcnt[8] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold92 (.A(_131_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold93 (.A(_015_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold94 (.A(\dc4.ho[0] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold95 (.A(_000_),
    .X(net112));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_210 ();
 sg13g2_decap_4 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_fill_1 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_320 ();
 sg13g2_decap_8 FILLER_24_327 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_4 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_123 ();
 sg13g2_decap_4 FILLER_25_138 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_decap_4 FILLER_25_151 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_decap_8 FILLER_25_166 ();
 sg13g2_decap_8 FILLER_25_173 ();
 sg13g2_decap_8 FILLER_25_180 ();
 sg13g2_decap_8 FILLER_25_187 ();
 sg13g2_fill_2 FILLER_25_194 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_decap_4 FILLER_25_268 ();
 sg13g2_fill_2 FILLER_25_272 ();
 sg13g2_fill_2 FILLER_25_309 ();
 sg13g2_decap_8 FILLER_25_320 ();
 sg13g2_fill_2 FILLER_25_327 ();
 sg13g2_fill_2 FILLER_25_332 ();
 sg13g2_decap_4 FILLER_25_348 ();
 sg13g2_fill_1 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_93 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_289 ();
 sg13g2_fill_2 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_4 FILLER_27_163 ();
 sg13g2_fill_1 FILLER_27_167 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_fill_2 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_fill_1 FILLER_27_339 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_4 FILLER_28_84 ();
 sg13g2_fill_1 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_fill_1 FILLER_28_176 ();
 sg13g2_fill_1 FILLER_28_181 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_4 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_154 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_297 ();
 sg13g2_fill_2 FILLER_29_335 ();
 sg13g2_fill_1 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_165 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_267 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_decap_4 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_4 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_decap_4 FILLER_31_164 ();
 sg13g2_decap_4 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_fill_2 FILLER_31_223 ();
 sg13g2_fill_2 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_323 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_160 ();
 sg13g2_fill_2 FILLER_32_166 ();
 sg13g2_decap_4 FILLER_32_182 ();
 sg13g2_fill_1 FILLER_32_207 ();
 sg13g2_fill_2 FILLER_32_276 ();
 sg13g2_fill_1 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_4 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_102 ();
 sg13g2_fill_2 FILLER_33_135 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_152 ();
 sg13g2_fill_2 FILLER_33_166 ();
 sg13g2_fill_1 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_198 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_2 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_358 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_4 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_172 ();
 sg13g2_decap_8 FILLER_34_181 ();
 sg13g2_decap_8 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_228 ();
 sg13g2_fill_2 FILLER_34_243 ();
 sg13g2_fill_2 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_decap_8 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_138 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_decap_4 FILLER_35_212 ();
 sg13g2_fill_2 FILLER_35_216 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_fill_2 FILLER_35_256 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_114 ();
 sg13g2_decap_4 FILLER_36_163 ();
 sg13g2_decap_8 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_193 ();
 sg13g2_fill_1 FILLER_36_195 ();
 sg13g2_fill_1 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_221 ();
 sg13g2_decap_8 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_121 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_fill_2 FILLER_37_218 ();
 sg13g2_fill_1 FILLER_37_306 ();
 sg13g2_decap_4 FILLER_37_334 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_4 FILLER_38_105 ();
 sg13g2_fill_2 FILLER_38_109 ();
 sg13g2_fill_2 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_145 ();
 sg13g2_decap_8 FILLER_38_176 ();
 sg13g2_decap_8 FILLER_38_183 ();
 sg13g2_decap_4 FILLER_38_190 ();
 sg13g2_fill_2 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_214 ();
 sg13g2_fill_2 FILLER_38_221 ();
 sg13g2_fill_1 FILLER_38_223 ();
 sg13g2_decap_4 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_4 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_out[6] = net3;
 assign uio_out[7] = net4;
endmodule

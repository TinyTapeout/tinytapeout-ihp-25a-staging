module tt_um_Rapoport (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire \perceptron1.out ;
 wire \perceptron1.we1[0] ;
 wire \perceptron1.we1[10] ;
 wire \perceptron1.we1[11] ;
 wire \perceptron1.we1[12] ;
 wire \perceptron1.we1[13] ;
 wire \perceptron1.we1[14] ;
 wire \perceptron1.we1[15] ;
 wire \perceptron1.we1[1] ;
 wire \perceptron1.we1[2] ;
 wire \perceptron1.we1[3] ;
 wire \perceptron1.we1[4] ;
 wire \perceptron1.we1[5] ;
 wire \perceptron1.we1[6] ;
 wire \perceptron1.we1[7] ;
 wire \perceptron1.we1[8] ;
 wire \perceptron1.we1[9] ;
 wire \perceptron1.we2[0] ;
 wire \perceptron1.we2[10] ;
 wire \perceptron1.we2[11] ;
 wire \perceptron1.we2[12] ;
 wire \perceptron1.we2[13] ;
 wire \perceptron1.we2[14] ;
 wire \perceptron1.we2[15] ;
 wire \perceptron1.we2[1] ;
 wire \perceptron1.we2[2] ;
 wire \perceptron1.we2[3] ;
 wire \perceptron1.we2[4] ;
 wire \perceptron1.we2[5] ;
 wire \perceptron1.we2[6] ;
 wire \perceptron1.we2[7] ;
 wire \perceptron1.we2[8] ;
 wire \perceptron1.we2[9] ;
 wire \perceptron1.we3[0] ;
 wire \perceptron1.we3[10] ;
 wire \perceptron1.we3[11] ;
 wire \perceptron1.we3[12] ;
 wire \perceptron1.we3[13] ;
 wire \perceptron1.we3[14] ;
 wire \perceptron1.we3[15] ;
 wire \perceptron1.we3[1] ;
 wire \perceptron1.we3[2] ;
 wire \perceptron1.we3[3] ;
 wire \perceptron1.we3[4] ;
 wire \perceptron1.we3[5] ;
 wire \perceptron1.we3[6] ;
 wire \perceptron1.we3[7] ;
 wire \perceptron1.we3[8] ;
 wire \perceptron1.we3[9] ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;

 sg13g2_inv_1 _1298_ (.Y(_0335_),
    .A(net40));
 sg13g2_inv_1 _1299_ (.Y(_0342_),
    .A(net298));
 sg13g2_inv_1 _1300_ (.Y(_0353_),
    .A(net286));
 sg13g2_inv_1 _1301_ (.Y(_0362_),
    .A(net279));
 sg13g2_inv_1 _1302_ (.Y(_0371_),
    .A(net281));
 sg13g2_inv_1 _1303_ (.Y(_0379_),
    .A(net59));
 sg13g2_inv_1 _1304_ (.Y(_0387_),
    .A(_0001_));
 sg13g2_and4_1 _1305_ (.A(net323),
    .B(net327),
    .C(\perceptron1.we1[2] ),
    .D(net274),
    .X(_0396_));
 sg13g2_nand2_1 _1306_ (.Y(_0402_),
    .A(net331),
    .B(\perceptron1.we1[4] ));
 sg13g2_a22oi_1 _1307_ (.Y(_0403_),
    .B1(net274),
    .B2(net327),
    .A2(\perceptron1.we1[2] ),
    .A1(net323));
 sg13g2_nor3_1 _1308_ (.A(_0396_),
    .B(_0402_),
    .C(_0403_),
    .Y(_0404_));
 sg13g2_or2_1 _1309_ (.X(_0405_),
    .B(_0404_),
    .A(_0396_));
 sg13g2_nand2_1 _1310_ (.Y(_0406_),
    .A(net331),
    .B(\perceptron1.we1[5] ));
 sg13g2_nand2_1 _1311_ (.Y(_0407_),
    .A(net323),
    .B(\perceptron1.we1[4] ));
 sg13g2_and4_1 _1312_ (.A(net323),
    .B(net327),
    .C(net274),
    .D(\perceptron1.we1[4] ),
    .X(_0408_));
 sg13g2_a22oi_1 _1313_ (.Y(_0409_),
    .B1(\perceptron1.we1[4] ),
    .B2(net327),
    .A2(net274),
    .A1(net323));
 sg13g2_nor3_1 _1314_ (.A(_0406_),
    .B(_0408_),
    .C(_0409_),
    .Y(_0410_));
 sg13g2_o21ai_1 _1315_ (.B1(_0406_),
    .Y(_0411_),
    .A1(_0408_),
    .A2(_0409_));
 sg13g2_nor2b_1 _1316_ (.A(_0410_),
    .B_N(_0411_),
    .Y(_0412_));
 sg13g2_nand2_1 _1317_ (.Y(_0413_),
    .A(_0405_),
    .B(_0412_));
 sg13g2_xnor2_1 _1318_ (.Y(_0414_),
    .A(_0405_),
    .B(_0412_));
 sg13g2_nand2_1 _1319_ (.Y(_0415_),
    .A(net303),
    .B(net280));
 sg13g2_and4_1 _1320_ (.A(net335),
    .B(net305),
    .C(\perceptron1.we1[6] ),
    .D(net279),
    .X(_0416_));
 sg13g2_a22oi_1 _1321_ (.Y(_0417_),
    .B1(net279),
    .B2(net305),
    .A2(\perceptron1.we1[6] ),
    .A1(net335));
 sg13g2_nor3_1 _1322_ (.A(_0415_),
    .B(_0416_),
    .C(_0417_),
    .Y(_0418_));
 sg13g2_o21ai_1 _1323_ (.B1(_0415_),
    .Y(_0419_),
    .A1(_0416_),
    .A2(_0417_));
 sg13g2_nand2b_1 _1324_ (.Y(_0420_),
    .B(_0419_),
    .A_N(_0418_));
 sg13g2_o21ai_1 _1325_ (.B1(_0413_),
    .Y(_0421_),
    .A1(_0414_),
    .A2(_0420_));
 sg13g2_nand2_1 _1326_ (.Y(_0422_),
    .A(net300),
    .B(\perceptron1.we3[6] ));
 sg13g2_and4_1 _1327_ (.A(net335),
    .B(net305),
    .C(\perceptron1.we1[7] ),
    .D(\perceptron1.we3[7] ),
    .X(_0423_));
 sg13g2_a22oi_1 _1328_ (.Y(_0424_),
    .B1(\perceptron1.we3[7] ),
    .B2(net304),
    .A2(\perceptron1.we1[7] ),
    .A1(net335));
 sg13g2_nor3_1 _1329_ (.A(_0422_),
    .B(_0423_),
    .C(_0424_),
    .Y(_0425_));
 sg13g2_o21ai_1 _1330_ (.B1(_0422_),
    .Y(_0426_),
    .A1(_0423_),
    .A2(_0424_));
 sg13g2_nand2b_1 _1331_ (.Y(_0427_),
    .B(_0426_),
    .A_N(_0425_));
 sg13g2_or2_1 _1332_ (.X(_0428_),
    .B(_0410_),
    .A(_0408_));
 sg13g2_nand2_1 _1333_ (.Y(_0429_),
    .A(net332),
    .B(\perceptron1.we1[6] ));
 sg13g2_nand2_1 _1334_ (.Y(_0430_),
    .A(net327),
    .B(net273));
 sg13g2_or2_1 _1335_ (.X(_0431_),
    .B(_0430_),
    .A(_0407_));
 sg13g2_and2_1 _1336_ (.A(_0407_),
    .B(_0430_),
    .X(_0432_));
 sg13g2_xor2_1 _1337_ (.B(_0430_),
    .A(_0407_),
    .X(_0433_));
 sg13g2_xnor2_1 _1338_ (.Y(_0434_),
    .A(_0429_),
    .B(_0433_));
 sg13g2_nand2_1 _1339_ (.Y(_0435_),
    .A(_0428_),
    .B(_0434_));
 sg13g2_xnor2_1 _1340_ (.Y(_0436_),
    .A(_0428_),
    .B(_0434_));
 sg13g2_xor2_1 _1341_ (.B(_0436_),
    .A(_0427_),
    .X(_0437_));
 sg13g2_nand2_1 _1342_ (.Y(_0438_),
    .A(_0421_),
    .B(_0437_));
 sg13g2_nand2_1 _1343_ (.Y(_0439_),
    .A(net294),
    .B(net281));
 sg13g2_and4_1 _1344_ (.A(net283),
    .B(net299),
    .C(net296),
    .D(\perceptron1.we3[4] ),
    .X(_0440_));
 sg13g2_nand2_1 _1345_ (.Y(_0441_),
    .A(\perceptron1.we3[2] ),
    .B(net293));
 sg13g2_a22oi_1 _1346_ (.Y(_0442_),
    .B1(\perceptron1.we3[4] ),
    .B2(net298),
    .A2(net296),
    .A1(net283));
 sg13g2_nor3_1 _1347_ (.A(_0440_),
    .B(_0441_),
    .C(_0442_),
    .Y(_0443_));
 sg13g2_or2_1 _1348_ (.X(_0444_),
    .B(_0443_),
    .A(_0440_));
 sg13g2_or2_1 _1349_ (.X(_0445_),
    .B(_0418_),
    .A(_0416_));
 sg13g2_nand2_1 _1350_ (.Y(_0446_),
    .A(net283),
    .B(net293));
 sg13g2_nand2_1 _1351_ (.Y(_0447_),
    .A(net294),
    .B(\perceptron1.we3[5] ));
 sg13g2_nand2_1 _1352_ (.Y(_0448_),
    .A(net297),
    .B(\perceptron1.we3[5] ));
 sg13g2_or2_1 _1353_ (.X(_0449_),
    .B(_0448_),
    .A(_0439_));
 sg13g2_xnor2_1 _1354_ (.Y(_0450_),
    .A(_0439_),
    .B(_0448_));
 sg13g2_xor2_1 _1355_ (.B(_0450_),
    .A(_0446_),
    .X(_0451_));
 sg13g2_xnor2_1 _1356_ (.Y(_0452_),
    .A(_0445_),
    .B(_0451_));
 sg13g2_nor2b_1 _1357_ (.A(_0452_),
    .B_N(_0444_),
    .Y(_0453_));
 sg13g2_xor2_1 _1358_ (.B(_0452_),
    .A(_0444_),
    .X(_0454_));
 sg13g2_xnor2_1 _1359_ (.Y(_0455_),
    .A(_0421_),
    .B(_0437_));
 sg13g2_o21ai_1 _1360_ (.B1(_0438_),
    .Y(_0456_),
    .A1(_0454_),
    .A2(_0455_));
 sg13g2_o21ai_1 _1361_ (.B1(_0435_),
    .Y(_0457_),
    .A1(_0427_),
    .A2(_0436_));
 sg13g2_o21ai_1 _1362_ (.B1(_0431_),
    .Y(_0458_),
    .A1(_0429_),
    .A2(_0432_));
 sg13g2_nand2_1 _1363_ (.Y(_0459_),
    .A(net330),
    .B(\perceptron1.we1[7] ));
 sg13g2_nand2_1 _1364_ (.Y(_0460_),
    .A(net322),
    .B(\perceptron1.we1[6] ));
 sg13g2_and4_1 _1365_ (.A(net322),
    .B(net325),
    .C(net273),
    .D(\perceptron1.we1[6] ),
    .X(_0461_));
 sg13g2_a22oi_1 _1366_ (.Y(_0462_),
    .B1(\perceptron1.we1[6] ),
    .B2(net326),
    .A2(net273),
    .A1(net321));
 sg13g2_nor3_1 _1367_ (.A(_0459_),
    .B(_0461_),
    .C(_0462_),
    .Y(_0463_));
 sg13g2_o21ai_1 _1368_ (.B1(_0459_),
    .Y(_0464_),
    .A1(_0461_),
    .A2(_0462_));
 sg13g2_nor2b_1 _1369_ (.A(_0463_),
    .B_N(_0464_),
    .Y(_0465_));
 sg13g2_nand2_1 _1370_ (.Y(_0466_),
    .A(_0458_),
    .B(_0465_));
 sg13g2_xnor2_1 _1371_ (.Y(_0467_),
    .A(_0458_),
    .B(_0465_));
 sg13g2_nand2_1 _1372_ (.Y(_0468_),
    .A(net300),
    .B(net278));
 sg13g2_and4_1 _1373_ (.A(net335),
    .B(net305),
    .C(net277),
    .D(\perceptron1.we1[8] ),
    .X(_0469_));
 sg13g2_a22oi_1 _1374_ (.Y(_0470_),
    .B1(\perceptron1.we1[8] ),
    .B2(net335),
    .A2(net277),
    .A1(net305));
 sg13g2_nor3_1 _1375_ (.A(_0468_),
    .B(_0469_),
    .C(_0470_),
    .Y(_0471_));
 sg13g2_o21ai_1 _1376_ (.B1(_0468_),
    .Y(_0472_),
    .A1(_0469_),
    .A2(_0470_));
 sg13g2_nand2b_1 _1377_ (.Y(_0473_),
    .B(_0472_),
    .A_N(_0471_));
 sg13g2_xor2_1 _1378_ (.B(_0473_),
    .A(_0467_),
    .X(_0474_));
 sg13g2_nand2_1 _1379_ (.Y(_0475_),
    .A(_0457_),
    .B(_0474_));
 sg13g2_xnor2_1 _1380_ (.Y(_0476_),
    .A(_0457_),
    .B(_0474_));
 sg13g2_o21ai_1 _1381_ (.B1(_0449_),
    .Y(_0477_),
    .A1(_0446_),
    .A2(_0450_));
 sg13g2_or2_1 _1382_ (.X(_0478_),
    .B(_0425_),
    .A(_0423_));
 sg13g2_nand2_1 _1383_ (.Y(_0479_),
    .A(net281),
    .B(net292));
 sg13g2_nand2_1 _1384_ (.Y(_0480_),
    .A(net294),
    .B(net279));
 sg13g2_nand2_1 _1385_ (.Y(_0481_),
    .A(net297),
    .B(net279));
 sg13g2_or2_1 _1386_ (.X(_0482_),
    .B(_0480_),
    .A(_0448_));
 sg13g2_xnor2_1 _1387_ (.Y(_0483_),
    .A(_0447_),
    .B(_0481_));
 sg13g2_xor2_1 _1388_ (.B(_0483_),
    .A(_0479_),
    .X(_0484_));
 sg13g2_xnor2_1 _1389_ (.Y(_0485_),
    .A(_0478_),
    .B(_0484_));
 sg13g2_nor2b_1 _1390_ (.A(_0485_),
    .B_N(_0477_),
    .Y(_0486_));
 sg13g2_xor2_1 _1391_ (.B(_0485_),
    .A(_0477_),
    .X(_0487_));
 sg13g2_xor2_1 _1392_ (.B(_0487_),
    .A(_0476_),
    .X(_0488_));
 sg13g2_nand2_1 _1393_ (.Y(_0489_),
    .A(_0456_),
    .B(_0488_));
 sg13g2_xnor2_1 _1394_ (.Y(_0490_),
    .A(_0456_),
    .B(_0488_));
 sg13g2_nand2_1 _1395_ (.Y(_0491_),
    .A(\perceptron1.we3[1] ),
    .B(net288));
 sg13g2_nand2_1 _1396_ (.Y(_0492_),
    .A(\perceptron1.we3[1] ),
    .B(net290));
 sg13g2_nand2_1 _1397_ (.Y(_0493_),
    .A(\perceptron1.we3[0] ),
    .B(net287));
 sg13g2_nand2_1 _1398_ (.Y(_0494_),
    .A(net318),
    .B(\perceptron1.we2[6] ));
 sg13g2_xor2_1 _1399_ (.B(_0493_),
    .A(_0492_),
    .X(_0495_));
 sg13g2_nand2b_1 _1400_ (.Y(_0496_),
    .B(_0495_),
    .A_N(_0494_));
 sg13g2_o21ai_1 _1401_ (.B1(_0496_),
    .Y(_0497_),
    .A1(_0492_),
    .A2(_0493_));
 sg13g2_nand2_1 _1402_ (.Y(_0498_),
    .A(net319),
    .B(\perceptron1.we2[7] ));
 sg13g2_nand2_1 _1403_ (.Y(_0499_),
    .A(\perceptron1.we3[2] ),
    .B(net287));
 sg13g2_nand2_1 _1404_ (.Y(_0500_),
    .A(net284),
    .B(net290));
 sg13g2_xor2_1 _1405_ (.B(_0500_),
    .A(_0491_),
    .X(_0501_));
 sg13g2_nand2b_1 _1406_ (.Y(_0502_),
    .B(_0501_),
    .A_N(_0498_));
 sg13g2_xnor2_1 _1407_ (.Y(_0503_),
    .A(_0498_),
    .B(_0501_));
 sg13g2_nand2_1 _1408_ (.Y(_0504_),
    .A(_0497_),
    .B(_0503_));
 sg13g2_nand2_1 _1409_ (.Y(_0505_),
    .A(net311),
    .B(\perceptron1.we2[4] ));
 sg13g2_nand2_1 _1410_ (.Y(_0506_),
    .A(net312),
    .B(\perceptron1.we2[6] ));
 sg13g2_nand2_1 _1411_ (.Y(_0507_),
    .A(net313),
    .B(\perceptron1.we2[5] ));
 sg13g2_nand2_1 _1412_ (.Y(_0508_),
    .A(net315),
    .B(\perceptron1.we2[6] ));
 sg13g2_xor2_1 _1413_ (.B(_0508_),
    .A(_0507_),
    .X(_0509_));
 sg13g2_nand2b_1 _1414_ (.Y(_0510_),
    .B(_0509_),
    .A_N(_0505_));
 sg13g2_xnor2_1 _1415_ (.Y(_0511_),
    .A(_0505_),
    .B(_0509_));
 sg13g2_inv_1 _1416_ (.Y(_0512_),
    .A(_0511_));
 sg13g2_xnor2_1 _1417_ (.Y(_0513_),
    .A(_0497_),
    .B(_0503_));
 sg13g2_o21ai_1 _1418_ (.B1(_0504_),
    .Y(_0514_),
    .A1(_0512_),
    .A2(_0513_));
 sg13g2_a21o_1 _1419_ (.A2(_0451_),
    .A1(_0445_),
    .B1(_0453_),
    .X(_0515_));
 sg13g2_o21ai_1 _1420_ (.B1(_0502_),
    .Y(_0516_),
    .A1(_0491_),
    .A2(_0500_));
 sg13g2_nand2_1 _1421_ (.Y(_0517_),
    .A(net320),
    .B(\perceptron1.we2[8] ));
 sg13g2_nand2_1 _1422_ (.Y(_0518_),
    .A(net283),
    .B(net288));
 sg13g2_nand2_1 _1423_ (.Y(_0519_),
    .A(net282),
    .B(net290));
 sg13g2_xor2_1 _1424_ (.B(_0519_),
    .A(_0499_),
    .X(_0520_));
 sg13g2_nand2b_1 _1425_ (.Y(_0521_),
    .B(_0520_),
    .A_N(_0517_));
 sg13g2_xnor2_1 _1426_ (.Y(_0522_),
    .A(_0517_),
    .B(_0520_));
 sg13g2_xnor2_1 _1427_ (.Y(_0523_),
    .A(_0516_),
    .B(_0522_));
 sg13g2_nand2_1 _1428_ (.Y(_0524_),
    .A(net310),
    .B(\perceptron1.we2[5] ));
 sg13g2_nand2_1 _1429_ (.Y(_0525_),
    .A(net312),
    .B(\perceptron1.we2[7] ));
 sg13g2_nand2_1 _1430_ (.Y(_0526_),
    .A(net315),
    .B(\perceptron1.we2[7] ));
 sg13g2_xor2_1 _1431_ (.B(_0526_),
    .A(_0506_),
    .X(_0527_));
 sg13g2_nand2b_1 _1432_ (.Y(_0528_),
    .B(_0527_),
    .A_N(_0524_));
 sg13g2_xnor2_1 _1433_ (.Y(_0529_),
    .A(_0524_),
    .B(_0527_));
 sg13g2_nor2b_1 _1434_ (.A(_0523_),
    .B_N(_0529_),
    .Y(_0530_));
 sg13g2_xnor2_1 _1435_ (.Y(_0531_),
    .A(_0523_),
    .B(_0529_));
 sg13g2_xnor2_1 _1436_ (.Y(_0532_),
    .A(_0515_),
    .B(_0531_));
 sg13g2_nor2b_1 _1437_ (.A(_0532_),
    .B_N(_0514_),
    .Y(_0533_));
 sg13g2_xor2_1 _1438_ (.B(_0532_),
    .A(_0514_),
    .X(_0534_));
 sg13g2_o21ai_1 _1439_ (.B1(_0489_),
    .Y(_0535_),
    .A1(_0490_),
    .A2(_0534_));
 sg13g2_o21ai_1 _1440_ (.B1(_0475_),
    .Y(_0536_),
    .A1(_0476_),
    .A2(_0487_));
 sg13g2_o21ai_1 _1441_ (.B1(_0466_),
    .Y(_0537_),
    .A1(_0467_),
    .A2(_0473_));
 sg13g2_or2_1 _1442_ (.X(_0538_),
    .B(_0463_),
    .A(_0461_));
 sg13g2_nand2_1 _1443_ (.Y(_0539_),
    .A(net330),
    .B(\perceptron1.we1[8] ));
 sg13g2_nand2_1 _1444_ (.Y(_0540_),
    .A(net326),
    .B(\perceptron1.we1[7] ));
 sg13g2_or2_1 _1445_ (.X(_0541_),
    .B(_0540_),
    .A(_0460_));
 sg13g2_and2_1 _1446_ (.A(_0460_),
    .B(_0540_),
    .X(_0542_));
 sg13g2_xor2_1 _1447_ (.B(_0540_),
    .A(_0460_),
    .X(_0543_));
 sg13g2_xnor2_1 _1448_ (.Y(_0544_),
    .A(_0539_),
    .B(_0543_));
 sg13g2_nand2_1 _1449_ (.Y(_0545_),
    .A(_0538_),
    .B(_0544_));
 sg13g2_xnor2_1 _1450_ (.Y(_0546_),
    .A(_0538_),
    .B(_0544_));
 sg13g2_nand2_1 _1451_ (.Y(_0547_),
    .A(net300),
    .B(net277));
 sg13g2_and4_1 _1452_ (.A(net334),
    .B(net304),
    .C(\perceptron1.we1[9] ),
    .D(\perceptron1.we3[9] ),
    .X(_0548_));
 sg13g2_a22oi_1 _1453_ (.Y(_0549_),
    .B1(\perceptron1.we3[9] ),
    .B2(net304),
    .A2(\perceptron1.we1[9] ),
    .A1(net334));
 sg13g2_nor3_1 _1454_ (.A(_0547_),
    .B(_0548_),
    .C(_0549_),
    .Y(_0550_));
 sg13g2_o21ai_1 _1455_ (.B1(_0547_),
    .Y(_0551_),
    .A1(_0548_),
    .A2(_0549_));
 sg13g2_nand2b_1 _1456_ (.Y(_0552_),
    .B(_0551_),
    .A_N(_0550_));
 sg13g2_xor2_1 _1457_ (.B(_0552_),
    .A(_0546_),
    .X(_0553_));
 sg13g2_nand2_1 _1458_ (.Y(_0554_),
    .A(_0537_),
    .B(_0553_));
 sg13g2_xnor2_1 _1459_ (.Y(_0555_),
    .A(_0537_),
    .B(_0553_));
 sg13g2_o21ai_1 _1460_ (.B1(_0482_),
    .Y(_0556_),
    .A1(_0479_),
    .A2(_0483_));
 sg13g2_or2_1 _1461_ (.X(_0557_),
    .B(_0471_),
    .A(_0469_));
 sg13g2_nand2_1 _1462_ (.Y(_0558_),
    .A(net280),
    .B(net292));
 sg13g2_nand2_1 _1463_ (.Y(_0559_),
    .A(net294),
    .B(net278));
 sg13g2_nand2_1 _1464_ (.Y(_0560_),
    .A(net297),
    .B(net278));
 sg13g2_or2_1 _1465_ (.X(_0561_),
    .B(_0559_),
    .A(_0481_));
 sg13g2_xnor2_1 _1466_ (.Y(_0562_),
    .A(_0480_),
    .B(_0560_));
 sg13g2_xor2_1 _1467_ (.B(_0562_),
    .A(_0558_),
    .X(_0563_));
 sg13g2_xnor2_1 _1468_ (.Y(_0564_),
    .A(_0557_),
    .B(_0563_));
 sg13g2_nor2b_1 _1469_ (.A(_0564_),
    .B_N(_0556_),
    .Y(_0565_));
 sg13g2_xor2_1 _1470_ (.B(_0564_),
    .A(_0556_),
    .X(_0566_));
 sg13g2_xor2_1 _1471_ (.B(_0566_),
    .A(_0555_),
    .X(_0567_));
 sg13g2_nand2_1 _1472_ (.Y(_0568_),
    .A(_0536_),
    .B(_0567_));
 sg13g2_xnor2_1 _1473_ (.Y(_0569_),
    .A(_0536_),
    .B(_0567_));
 sg13g2_a21o_1 _1474_ (.A2(_0522_),
    .A1(_0516_),
    .B1(_0530_),
    .X(_0570_));
 sg13g2_a21o_1 _1475_ (.A2(_0484_),
    .A1(_0478_),
    .B1(_0486_),
    .X(_0571_));
 sg13g2_o21ai_1 _1476_ (.B1(_0521_),
    .Y(_0572_),
    .A1(_0499_),
    .A2(_0519_));
 sg13g2_nand2_1 _1477_ (.Y(_0573_),
    .A(net320),
    .B(\perceptron1.we2[9] ));
 sg13g2_nand2_1 _1478_ (.Y(_0574_),
    .A(net281),
    .B(net287));
 sg13g2_nand2_1 _1479_ (.Y(_0575_),
    .A(net281),
    .B(net289));
 sg13g2_xor2_1 _1480_ (.B(_0575_),
    .A(_0518_),
    .X(_0576_));
 sg13g2_nand2b_1 _1481_ (.Y(_0577_),
    .B(_0576_),
    .A_N(_0573_));
 sg13g2_xnor2_1 _1482_ (.Y(_0578_),
    .A(_0573_),
    .B(_0576_));
 sg13g2_xnor2_1 _1483_ (.Y(_0579_),
    .A(_0572_),
    .B(_0578_));
 sg13g2_nand2_1 _1484_ (.Y(_0580_),
    .A(net310),
    .B(\perceptron1.we2[6] ));
 sg13g2_nand2_1 _1485_ (.Y(_0581_),
    .A(net314),
    .B(\perceptron1.we2[8] ));
 sg13g2_nand2_1 _1486_ (.Y(_0582_),
    .A(net317),
    .B(\perceptron1.we2[8] ));
 sg13g2_xor2_1 _1487_ (.B(_0582_),
    .A(_0525_),
    .X(_0583_));
 sg13g2_nand2b_1 _1488_ (.Y(_0584_),
    .B(_0583_),
    .A_N(_0580_));
 sg13g2_xnor2_1 _1489_ (.Y(_0585_),
    .A(_0580_),
    .B(_0583_));
 sg13g2_nor2b_1 _1490_ (.A(_0579_),
    .B_N(_0585_),
    .Y(_0586_));
 sg13g2_xnor2_1 _1491_ (.Y(_0587_),
    .A(_0579_),
    .B(_0585_));
 sg13g2_xnor2_1 _1492_ (.Y(_0588_),
    .A(_0571_),
    .B(_0587_));
 sg13g2_nor2b_1 _1493_ (.A(_0588_),
    .B_N(_0570_),
    .Y(_0589_));
 sg13g2_xor2_1 _1494_ (.B(_0588_),
    .A(_0570_),
    .X(_0590_));
 sg13g2_xor2_1 _1495_ (.B(_0590_),
    .A(_0569_),
    .X(_0591_));
 sg13g2_a21o_1 _1496_ (.A2(_0531_),
    .A1(_0515_),
    .B1(_0533_),
    .X(_0592_));
 sg13g2_xnor2_1 _1497_ (.Y(_0593_),
    .A(_0535_),
    .B(_0591_));
 sg13g2_nor2b_1 _1498_ (.A(_0593_),
    .B_N(_0592_),
    .Y(_0594_));
 sg13g2_a21o_1 _1499_ (.A2(_0591_),
    .A1(_0535_),
    .B1(_0594_),
    .X(_0595_));
 sg13g2_a21o_1 _1500_ (.A2(_0587_),
    .A1(_0571_),
    .B1(_0589_),
    .X(_0596_));
 sg13g2_o21ai_1 _1501_ (.B1(_0568_),
    .Y(_0597_),
    .A1(_0569_),
    .A2(_0590_));
 sg13g2_o21ai_1 _1502_ (.B1(_0554_),
    .Y(_0598_),
    .A1(_0555_),
    .A2(_0566_));
 sg13g2_o21ai_1 _1503_ (.B1(_0545_),
    .Y(_0599_),
    .A1(_0546_),
    .A2(_0552_));
 sg13g2_o21ai_1 _1504_ (.B1(_0541_),
    .Y(_0600_),
    .A1(_0539_),
    .A2(_0542_));
 sg13g2_nand2_1 _1505_ (.Y(_0601_),
    .A(net330),
    .B(\perceptron1.we1[9] ));
 sg13g2_nand2_1 _1506_ (.Y(_0602_),
    .A(net321),
    .B(\perceptron1.we1[8] ));
 sg13g2_and4_1 _1507_ (.A(net322),
    .B(net326),
    .C(\perceptron1.we1[7] ),
    .D(\perceptron1.we1[8] ),
    .X(_0603_));
 sg13g2_a22oi_1 _1508_ (.Y(_0604_),
    .B1(\perceptron1.we1[8] ),
    .B2(net326),
    .A2(\perceptron1.we1[7] ),
    .A1(net322));
 sg13g2_nor3_1 _1509_ (.A(_0601_),
    .B(_0603_),
    .C(_0604_),
    .Y(_0605_));
 sg13g2_o21ai_1 _1510_ (.B1(_0601_),
    .Y(_0606_),
    .A1(_0603_),
    .A2(_0604_));
 sg13g2_nor2b_1 _1511_ (.A(_0605_),
    .B_N(_0606_),
    .Y(_0607_));
 sg13g2_nand2_1 _1512_ (.Y(_0608_),
    .A(_0600_),
    .B(_0607_));
 sg13g2_xnor2_1 _1513_ (.Y(_0609_),
    .A(_0600_),
    .B(_0607_));
 sg13g2_nand2_1 _1514_ (.Y(_0610_),
    .A(net300),
    .B(net276));
 sg13g2_and4_1 _1515_ (.A(net333),
    .B(net304),
    .C(\perceptron1.we1[10] ),
    .D(net275),
    .X(_0611_));
 sg13g2_a22oi_1 _1516_ (.Y(_0612_),
    .B1(net275),
    .B2(net304),
    .A2(\perceptron1.we1[10] ),
    .A1(net333));
 sg13g2_nor3_1 _1517_ (.A(_0610_),
    .B(_0611_),
    .C(_0612_),
    .Y(_0613_));
 sg13g2_o21ai_1 _1518_ (.B1(_0610_),
    .Y(_0614_),
    .A1(_0611_),
    .A2(_0612_));
 sg13g2_nand2b_1 _1519_ (.Y(_0615_),
    .B(_0614_),
    .A_N(_0613_));
 sg13g2_xor2_1 _1520_ (.B(_0615_),
    .A(_0609_),
    .X(_0616_));
 sg13g2_nand2_1 _1521_ (.Y(_0617_),
    .A(_0599_),
    .B(_0616_));
 sg13g2_xnor2_1 _1522_ (.Y(_0618_),
    .A(_0599_),
    .B(_0616_));
 sg13g2_o21ai_1 _1523_ (.B1(_0561_),
    .Y(_0619_),
    .A1(_0558_),
    .A2(_0562_));
 sg13g2_or2_1 _1524_ (.X(_0620_),
    .B(_0550_),
    .A(_0548_));
 sg13g2_nand2_1 _1525_ (.Y(_0621_),
    .A(net279),
    .B(net292));
 sg13g2_nand2_1 _1526_ (.Y(_0622_),
    .A(net294),
    .B(net277));
 sg13g2_nand2_1 _1527_ (.Y(_0623_),
    .A(net297),
    .B(net277));
 sg13g2_or2_1 _1528_ (.X(_0624_),
    .B(_0622_),
    .A(_0560_));
 sg13g2_xnor2_1 _1529_ (.Y(_0625_),
    .A(_0559_),
    .B(_0623_));
 sg13g2_xor2_1 _1530_ (.B(_0625_),
    .A(_0621_),
    .X(_0626_));
 sg13g2_xnor2_1 _1531_ (.Y(_0627_),
    .A(_0620_),
    .B(_0626_));
 sg13g2_nor2b_1 _1532_ (.A(_0627_),
    .B_N(_0619_),
    .Y(_0628_));
 sg13g2_xor2_1 _1533_ (.B(_0627_),
    .A(_0619_),
    .X(_0629_));
 sg13g2_xor2_1 _1534_ (.B(_0629_),
    .A(_0618_),
    .X(_0630_));
 sg13g2_nand2_1 _1535_ (.Y(_0631_),
    .A(_0598_),
    .B(_0630_));
 sg13g2_xnor2_1 _1536_ (.Y(_0632_),
    .A(_0598_),
    .B(_0630_));
 sg13g2_a21o_1 _1537_ (.A2(_0578_),
    .A1(_0572_),
    .B1(_0586_),
    .X(_0633_));
 sg13g2_a21o_1 _1538_ (.A2(_0563_),
    .A1(_0557_),
    .B1(_0565_),
    .X(_0634_));
 sg13g2_o21ai_1 _1539_ (.B1(_0577_),
    .Y(_0635_),
    .A1(_0518_),
    .A2(_0575_));
 sg13g2_nand2_1 _1540_ (.Y(_0636_),
    .A(net320),
    .B(\perceptron1.we2[10] ));
 sg13g2_nand2_1 _1541_ (.Y(_0637_),
    .A(net280),
    .B(net287));
 sg13g2_nand2_1 _1542_ (.Y(_0638_),
    .A(net280),
    .B(net289));
 sg13g2_xor2_1 _1543_ (.B(_0638_),
    .A(_0574_),
    .X(_0639_));
 sg13g2_nand2b_1 _1544_ (.Y(_0640_),
    .B(_0639_),
    .A_N(_0636_));
 sg13g2_xnor2_1 _1545_ (.Y(_0641_),
    .A(_0636_),
    .B(_0639_));
 sg13g2_xnor2_1 _1546_ (.Y(_0642_),
    .A(_0635_),
    .B(_0641_));
 sg13g2_nand2_1 _1547_ (.Y(_0643_),
    .A(net311),
    .B(\perceptron1.we2[7] ));
 sg13g2_nand2_1 _1548_ (.Y(_0644_),
    .A(net314),
    .B(\perceptron1.we2[9] ));
 sg13g2_nand2_1 _1549_ (.Y(_0645_),
    .A(net317),
    .B(\perceptron1.we2[9] ));
 sg13g2_xor2_1 _1550_ (.B(_0645_),
    .A(_0581_),
    .X(_0646_));
 sg13g2_nand2b_1 _1551_ (.Y(_0647_),
    .B(_0646_),
    .A_N(_0643_));
 sg13g2_xnor2_1 _1552_ (.Y(_0648_),
    .A(_0643_),
    .B(_0646_));
 sg13g2_nor2b_1 _1553_ (.A(_0642_),
    .B_N(_0648_),
    .Y(_0649_));
 sg13g2_xnor2_1 _1554_ (.Y(_0650_),
    .A(_0642_),
    .B(_0648_));
 sg13g2_xnor2_1 _1555_ (.Y(_0651_),
    .A(_0634_),
    .B(_0650_));
 sg13g2_nor2b_1 _1556_ (.A(_0651_),
    .B_N(_0633_),
    .Y(_0652_));
 sg13g2_xor2_1 _1557_ (.B(_0651_),
    .A(_0633_),
    .X(_0653_));
 sg13g2_xor2_1 _1558_ (.B(_0653_),
    .A(_0632_),
    .X(_0654_));
 sg13g2_nand2_1 _1559_ (.Y(_0655_),
    .A(_0597_),
    .B(_0654_));
 sg13g2_xnor2_1 _1560_ (.Y(_0656_),
    .A(_0597_),
    .B(_0654_));
 sg13g2_nand2b_1 _1561_ (.Y(_0657_),
    .B(_0596_),
    .A_N(_0656_));
 sg13g2_xor2_1 _1562_ (.B(_0656_),
    .A(_0596_),
    .X(_0658_));
 sg13g2_nand2b_1 _1563_ (.Y(_0659_),
    .B(_0595_),
    .A_N(_0658_));
 sg13g2_o21ai_1 _1564_ (.B1(_0584_),
    .Y(_0660_),
    .A1(_0525_),
    .A2(_0582_));
 sg13g2_inv_1 _1565_ (.Y(_0661_),
    .A(_0660_));
 sg13g2_xor2_1 _1566_ (.B(_0658_),
    .A(_0595_),
    .X(_0662_));
 sg13g2_o21ai_1 _1567_ (.B1(_0659_),
    .Y(_0663_),
    .A1(_0661_),
    .A2(_0662_));
 sg13g2_o21ai_1 _1568_ (.B1(_0647_),
    .Y(_0664_),
    .A1(_0581_),
    .A2(_0645_));
 sg13g2_nand2_1 _1569_ (.Y(_0665_),
    .A(_0655_),
    .B(_0657_));
 sg13g2_a21o_1 _1570_ (.A2(_0650_),
    .A1(_0634_),
    .B1(_0652_),
    .X(_0666_));
 sg13g2_o21ai_1 _1571_ (.B1(_0631_),
    .Y(_0667_),
    .A1(_0632_),
    .A2(_0653_));
 sg13g2_o21ai_1 _1572_ (.B1(_0617_),
    .Y(_0668_),
    .A1(_0618_),
    .A2(_0629_));
 sg13g2_o21ai_1 _1573_ (.B1(_0608_),
    .Y(_0669_),
    .A1(_0609_),
    .A2(_0615_));
 sg13g2_or2_1 _1574_ (.X(_0670_),
    .B(_0605_),
    .A(_0603_));
 sg13g2_nand2_1 _1575_ (.Y(_0671_),
    .A(net330),
    .B(\perceptron1.we1[10] ));
 sg13g2_nand2_1 _1576_ (.Y(_0672_),
    .A(net325),
    .B(\perceptron1.we1[9] ));
 sg13g2_or2_1 _1577_ (.X(_0673_),
    .B(_0672_),
    .A(_0602_));
 sg13g2_and2_1 _1578_ (.A(_0602_),
    .B(_0672_),
    .X(_0674_));
 sg13g2_xor2_1 _1579_ (.B(_0672_),
    .A(_0602_),
    .X(_0675_));
 sg13g2_xnor2_1 _1580_ (.Y(_0676_),
    .A(_0671_),
    .B(_0675_));
 sg13g2_nand2_1 _1581_ (.Y(_0677_),
    .A(_0670_),
    .B(_0676_));
 sg13g2_xnor2_1 _1582_ (.Y(_0678_),
    .A(_0670_),
    .B(_0676_));
 sg13g2_nand2_1 _1583_ (.Y(_0679_),
    .A(net303),
    .B(net275));
 sg13g2_and4_1 _1584_ (.A(net334),
    .B(net304),
    .C(net272),
    .D(\perceptron1.we3[11] ),
    .X(_0680_));
 sg13g2_a22oi_1 _1585_ (.Y(_0681_),
    .B1(\perceptron1.we3[11] ),
    .B2(net304),
    .A2(net272),
    .A1(net334));
 sg13g2_nor3_1 _1586_ (.A(_0679_),
    .B(_0680_),
    .C(_0681_),
    .Y(_0682_));
 sg13g2_o21ai_1 _1587_ (.B1(_0679_),
    .Y(_0683_),
    .A1(_0680_),
    .A2(_0681_));
 sg13g2_nand2b_1 _1588_ (.Y(_0684_),
    .B(_0683_),
    .A_N(_0682_));
 sg13g2_xor2_1 _1589_ (.B(_0684_),
    .A(_0678_),
    .X(_0685_));
 sg13g2_nand2_1 _1590_ (.Y(_0686_),
    .A(_0669_),
    .B(_0685_));
 sg13g2_xnor2_1 _1591_ (.Y(_0687_),
    .A(_0669_),
    .B(_0685_));
 sg13g2_o21ai_1 _1592_ (.B1(_0624_),
    .Y(_0688_),
    .A1(_0621_),
    .A2(_0625_));
 sg13g2_or2_1 _1593_ (.X(_0689_),
    .B(_0613_),
    .A(_0611_));
 sg13g2_nand2_1 _1594_ (.Y(_0690_),
    .A(net278),
    .B(net292));
 sg13g2_nand2_1 _1595_ (.Y(_0691_),
    .A(net1),
    .B(net276));
 sg13g2_nand2_1 _1596_ (.Y(_0692_),
    .A(net299),
    .B(net276));
 sg13g2_or2_1 _1597_ (.X(_0693_),
    .B(_0691_),
    .A(_0623_));
 sg13g2_xnor2_1 _1598_ (.Y(_0694_),
    .A(_0622_),
    .B(_0692_));
 sg13g2_xor2_1 _1599_ (.B(_0694_),
    .A(_0690_),
    .X(_0695_));
 sg13g2_xnor2_1 _1600_ (.Y(_0696_),
    .A(_0689_),
    .B(_0695_));
 sg13g2_nor2b_1 _1601_ (.A(_0696_),
    .B_N(_0688_),
    .Y(_0697_));
 sg13g2_xor2_1 _1602_ (.B(_0696_),
    .A(_0688_),
    .X(_0698_));
 sg13g2_xor2_1 _1603_ (.B(_0698_),
    .A(_0687_),
    .X(_0699_));
 sg13g2_nand2_1 _1604_ (.Y(_0700_),
    .A(_0668_),
    .B(_0699_));
 sg13g2_xnor2_1 _1605_ (.Y(_0701_),
    .A(_0668_),
    .B(_0699_));
 sg13g2_a21o_1 _1606_ (.A2(_0641_),
    .A1(_0635_),
    .B1(_0649_),
    .X(_0702_));
 sg13g2_a21o_1 _1607_ (.A2(_0626_),
    .A1(_0620_),
    .B1(_0628_),
    .X(_0703_));
 sg13g2_o21ai_1 _1608_ (.B1(_0640_),
    .Y(_0704_),
    .A1(_0574_),
    .A2(_0638_));
 sg13g2_nand2_1 _1609_ (.Y(_0705_),
    .A(net320),
    .B(\perceptron1.we2[11] ));
 sg13g2_nand2_1 _1610_ (.Y(_0706_),
    .A(\perceptron1.we3[6] ),
    .B(net287));
 sg13g2_nand2_1 _1611_ (.Y(_0707_),
    .A(net279),
    .B(net289));
 sg13g2_xor2_1 _1612_ (.B(_0707_),
    .A(_0637_),
    .X(_0708_));
 sg13g2_nand2b_1 _1613_ (.Y(_0709_),
    .B(_0708_),
    .A_N(_0705_));
 sg13g2_xnor2_1 _1614_ (.Y(_0710_),
    .A(_0705_),
    .B(_0708_));
 sg13g2_xnor2_1 _1615_ (.Y(_0711_),
    .A(_0704_),
    .B(_0710_));
 sg13g2_nand2_1 _1616_ (.Y(_0712_),
    .A(net311),
    .B(\perceptron1.we2[8] ));
 sg13g2_nand2_2 _1617_ (.Y(_0713_),
    .A(net317),
    .B(\perceptron1.we2[10] ));
 sg13g2_xor2_1 _1618_ (.B(_0713_),
    .A(_0644_),
    .X(_0714_));
 sg13g2_nand2b_1 _1619_ (.Y(_0715_),
    .B(_0714_),
    .A_N(_0712_));
 sg13g2_xnor2_1 _1620_ (.Y(_0716_),
    .A(_0712_),
    .B(_0714_));
 sg13g2_nor2b_1 _1621_ (.A(_0711_),
    .B_N(_0716_),
    .Y(_0717_));
 sg13g2_xnor2_1 _1622_ (.Y(_0718_),
    .A(_0711_),
    .B(_0716_));
 sg13g2_xnor2_1 _1623_ (.Y(_0719_),
    .A(_0703_),
    .B(_0718_));
 sg13g2_nor2b_1 _1624_ (.A(_0719_),
    .B_N(_0702_),
    .Y(_0720_));
 sg13g2_xor2_1 _1625_ (.B(_0719_),
    .A(_0702_),
    .X(_0721_));
 sg13g2_xor2_1 _1626_ (.B(_0721_),
    .A(_0701_),
    .X(_0722_));
 sg13g2_xnor2_1 _1627_ (.Y(_0723_),
    .A(_0667_),
    .B(_0722_));
 sg13g2_nor2b_1 _1628_ (.A(_0723_),
    .B_N(_0666_),
    .Y(_0724_));
 sg13g2_xor2_1 _1629_ (.B(_0723_),
    .A(_0666_),
    .X(_0725_));
 sg13g2_a21oi_1 _1630_ (.A1(_0655_),
    .A2(_0657_),
    .Y(_0726_),
    .B1(_0725_));
 sg13g2_xor2_1 _1631_ (.B(_0725_),
    .A(_0665_),
    .X(_0727_));
 sg13g2_nor2b_1 _1632_ (.A(_0727_),
    .B_N(_0664_),
    .Y(_0728_));
 sg13g2_xor2_1 _1633_ (.B(_0727_),
    .A(_0664_),
    .X(_0729_));
 sg13g2_nand2b_1 _1634_ (.Y(_0730_),
    .B(_0663_),
    .A_N(_0729_));
 sg13g2_xnor2_1 _1635_ (.Y(_0731_),
    .A(_0663_),
    .B(_0729_));
 sg13g2_nand2_2 _1636_ (.Y(_0732_),
    .A(net328),
    .B(\perceptron1.we1[1] ));
 sg13g2_and4_1 _1637_ (.A(net324),
    .B(net328),
    .C(\perceptron1.we1[1] ),
    .D(\perceptron1.we1[2] ),
    .X(_0733_));
 sg13g2_nand2_1 _1638_ (.Y(_0734_),
    .A(net332),
    .B(\perceptron1.we1[3] ));
 sg13g2_a22oi_1 _1639_ (.Y(_0735_),
    .B1(\perceptron1.we1[2] ),
    .B2(net328),
    .A2(\perceptron1.we1[1] ),
    .A1(net323));
 sg13g2_nor3_1 _1640_ (.A(_0733_),
    .B(_0734_),
    .C(_0735_),
    .Y(_0736_));
 sg13g2_or2_1 _1641_ (.X(_0737_),
    .B(_0736_),
    .A(_0733_));
 sg13g2_o21ai_1 _1642_ (.B1(_0402_),
    .Y(_0738_),
    .A1(_0396_),
    .A2(_0403_));
 sg13g2_nor2b_1 _1643_ (.A(_0404_),
    .B_N(_0738_),
    .Y(_0739_));
 sg13g2_nand2_1 _1644_ (.Y(_0740_),
    .A(_0737_),
    .B(_0739_));
 sg13g2_xnor2_1 _1645_ (.Y(_0741_),
    .A(_0737_),
    .B(_0739_));
 sg13g2_nand2_1 _1646_ (.Y(_0742_),
    .A(net302),
    .B(net281));
 sg13g2_and4_1 _1647_ (.A(net336),
    .B(net309),
    .C(net273),
    .D(net280),
    .X(_0743_));
 sg13g2_a22oi_1 _1648_ (.Y(_0744_),
    .B1(net280),
    .B2(net309),
    .A2(net273),
    .A1(net336));
 sg13g2_nor3_1 _1649_ (.A(_0742_),
    .B(_0743_),
    .C(_0744_),
    .Y(_0745_));
 sg13g2_o21ai_1 _1650_ (.B1(_0742_),
    .Y(_0746_),
    .A1(_0743_),
    .A2(_0744_));
 sg13g2_nand2b_1 _1651_ (.Y(_0747_),
    .B(_0746_),
    .A_N(_0745_));
 sg13g2_o21ai_1 _1652_ (.B1(_0740_),
    .Y(_0748_),
    .A1(_0741_),
    .A2(_0747_));
 sg13g2_xor2_1 _1653_ (.B(_0420_),
    .A(_0414_),
    .X(_0749_));
 sg13g2_nand2_1 _1654_ (.Y(_0750_),
    .A(_0748_),
    .B(_0749_));
 sg13g2_xnor2_1 _1655_ (.Y(_0751_),
    .A(_0748_),
    .B(_0749_));
 sg13g2_and4_1 _1656_ (.A(net282),
    .B(net284),
    .C(net299),
    .D(net296),
    .X(_0752_));
 sg13g2_nand2_1 _1657_ (.Y(_0753_),
    .A(\perceptron1.we3[1] ),
    .B(net293));
 sg13g2_a22oi_1 _1658_ (.Y(_0754_),
    .B1(net296),
    .B2(\perceptron1.we3[2] ),
    .A2(net299),
    .A1(net283));
 sg13g2_nor3_1 _1659_ (.A(_0752_),
    .B(_0753_),
    .C(_0754_),
    .Y(_0755_));
 sg13g2_or2_1 _1660_ (.X(_0756_),
    .B(_0755_),
    .A(_0752_));
 sg13g2_or2_1 _1661_ (.X(_0757_),
    .B(_0745_),
    .A(_0743_));
 sg13g2_o21ai_1 _1662_ (.B1(_0441_),
    .Y(_0758_),
    .A1(_0440_),
    .A2(_0442_));
 sg13g2_nor2b_1 _1663_ (.A(_0443_),
    .B_N(_0758_),
    .Y(_0759_));
 sg13g2_xnor2_1 _1664_ (.Y(_0760_),
    .A(_0757_),
    .B(_0759_));
 sg13g2_nor2b_1 _1665_ (.A(_0760_),
    .B_N(_0756_),
    .Y(_0761_));
 sg13g2_xor2_1 _1666_ (.B(_0760_),
    .A(_0756_),
    .X(_0762_));
 sg13g2_o21ai_1 _1667_ (.B1(_0750_),
    .Y(_0763_),
    .A1(_0751_),
    .A2(_0762_));
 sg13g2_xor2_1 _1668_ (.B(_0455_),
    .A(_0454_),
    .X(_0764_));
 sg13g2_nand2_1 _1669_ (.Y(_0765_),
    .A(_0763_),
    .B(_0764_));
 sg13g2_and4_1 _1670_ (.A(net286),
    .B(net318),
    .C(net290),
    .D(\perceptron1.we2[5] ),
    .X(_0766_));
 sg13g2_xnor2_1 _1671_ (.Y(_0767_),
    .A(_0494_),
    .B(_0495_));
 sg13g2_and2_1 _1672_ (.A(_0766_),
    .B(_0767_),
    .X(_0768_));
 sg13g2_xor2_1 _1673_ (.B(_0767_),
    .A(_0766_),
    .X(_0769_));
 sg13g2_nand2_1 _1674_ (.Y(_0770_),
    .A(\perceptron1.we2[3] ),
    .B(net310));
 sg13g2_nand2_1 _1675_ (.Y(_0771_),
    .A(net315),
    .B(\perceptron1.we2[4] ));
 sg13g2_nor2_1 _1676_ (.A(_0507_),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_a22oi_1 _1677_ (.Y(_0773_),
    .B1(\perceptron1.we2[4] ),
    .B2(net312),
    .A2(\perceptron1.we2[5] ),
    .A1(net315));
 sg13g2_nor3_1 _1678_ (.A(_0770_),
    .B(_0772_),
    .C(_0773_),
    .Y(_0774_));
 sg13g2_o21ai_1 _1679_ (.B1(_0770_),
    .Y(_0775_),
    .A1(_0772_),
    .A2(_0773_));
 sg13g2_nor2b_1 _1680_ (.A(_0774_),
    .B_N(_0775_),
    .Y(_0776_));
 sg13g2_a21o_1 _1681_ (.A2(_0776_),
    .A1(_0769_),
    .B1(_0768_),
    .X(_0777_));
 sg13g2_a21o_1 _1682_ (.A2(_0759_),
    .A1(_0757_),
    .B1(_0761_),
    .X(_0778_));
 sg13g2_inv_1 _1683_ (.Y(_0779_),
    .A(_0778_));
 sg13g2_xnor2_1 _1684_ (.Y(_0780_),
    .A(_0512_),
    .B(_0513_));
 sg13g2_xor2_1 _1685_ (.B(_0780_),
    .A(_0778_),
    .X(_0781_));
 sg13g2_nand2b_1 _1686_ (.Y(_0782_),
    .B(_0777_),
    .A_N(_0781_));
 sg13g2_xor2_1 _1687_ (.B(_0781_),
    .A(_0777_),
    .X(_0783_));
 sg13g2_xnor2_1 _1688_ (.Y(_0784_),
    .A(_0763_),
    .B(_0764_));
 sg13g2_o21ai_1 _1689_ (.B1(_0765_),
    .Y(_0785_),
    .A1(_0783_),
    .A2(_0784_));
 sg13g2_xor2_1 _1690_ (.B(_0534_),
    .A(_0490_),
    .X(_0786_));
 sg13g2_o21ai_1 _1691_ (.B1(_0782_),
    .Y(_0787_),
    .A1(_0779_),
    .A2(_0780_));
 sg13g2_xnor2_1 _1692_ (.Y(_0788_),
    .A(_0785_),
    .B(_0786_));
 sg13g2_nor2b_1 _1693_ (.A(_0788_),
    .B_N(_0787_),
    .Y(_0789_));
 sg13g2_a21o_1 _1694_ (.A2(_0786_),
    .A1(_0785_),
    .B1(_0789_),
    .X(_0790_));
 sg13g2_xor2_1 _1695_ (.B(_0593_),
    .A(_0592_),
    .X(_0791_));
 sg13g2_nand2b_1 _1696_ (.Y(_0792_),
    .B(_0790_),
    .A_N(_0791_));
 sg13g2_o21ai_1 _1697_ (.B1(_0528_),
    .Y(_0793_),
    .A1(_0506_),
    .A2(_0526_));
 sg13g2_xor2_1 _1698_ (.B(_0791_),
    .A(_0790_),
    .X(_0794_));
 sg13g2_nand2b_1 _1699_ (.Y(_0795_),
    .B(_0793_),
    .A_N(_0794_));
 sg13g2_xnor2_1 _1700_ (.Y(_0796_),
    .A(_0661_),
    .B(_0662_));
 sg13g2_a21oi_1 _1701_ (.A1(_0792_),
    .A2(_0795_),
    .Y(_0797_),
    .B1(_0796_));
 sg13g2_a21o_1 _1702_ (.A2(_0795_),
    .A1(_0792_),
    .B1(_0796_),
    .X(_0798_));
 sg13g2_nand3_1 _1703_ (.B(_0795_),
    .C(_0796_),
    .A(_0792_),
    .Y(_0799_));
 sg13g2_and3_1 _1704_ (.X(_0800_),
    .A(_0731_),
    .B(_0798_),
    .C(_0799_));
 sg13g2_nand2_1 _1705_ (.Y(_0801_),
    .A(net323),
    .B(\perceptron1.we1[0] ));
 sg13g2_or2_1 _1706_ (.X(_0802_),
    .B(_0801_),
    .A(_0732_));
 sg13g2_nand2_1 _1707_ (.Y(_0803_),
    .A(net331),
    .B(\perceptron1.we1[2] ));
 sg13g2_and2_1 _1708_ (.A(_0732_),
    .B(_0801_),
    .X(_0804_));
 sg13g2_xor2_1 _1709_ (.B(_0801_),
    .A(_0732_),
    .X(_0805_));
 sg13g2_o21ai_1 _1710_ (.B1(_0802_),
    .Y(_0806_),
    .A1(_0803_),
    .A2(_0804_));
 sg13g2_o21ai_1 _1711_ (.B1(_0734_),
    .Y(_0807_),
    .A1(_0733_),
    .A2(_0735_));
 sg13g2_nor2b_1 _1712_ (.A(_0736_),
    .B_N(_0807_),
    .Y(_0808_));
 sg13g2_nand2_1 _1713_ (.Y(_0809_),
    .A(_0806_),
    .B(_0808_));
 sg13g2_xnor2_1 _1714_ (.Y(_0810_),
    .A(_0806_),
    .B(_0808_));
 sg13g2_nand2_1 _1715_ (.Y(_0811_),
    .A(net282),
    .B(net302));
 sg13g2_and4_1 _1716_ (.A(net336),
    .B(net309),
    .C(\perceptron1.we1[4] ),
    .D(net281),
    .X(_0812_));
 sg13g2_a22oi_1 _1717_ (.Y(_0813_),
    .B1(net281),
    .B2(net309),
    .A2(\perceptron1.we1[4] ),
    .A1(net336));
 sg13g2_nor3_1 _1718_ (.A(_0811_),
    .B(_0812_),
    .C(_0813_),
    .Y(_0814_));
 sg13g2_o21ai_1 _1719_ (.B1(_0811_),
    .Y(_0815_),
    .A1(_0812_),
    .A2(_0813_));
 sg13g2_nand2b_1 _1720_ (.Y(_0816_),
    .B(_0815_),
    .A_N(_0814_));
 sg13g2_o21ai_1 _1721_ (.B1(_0809_),
    .Y(_0817_),
    .A1(_0810_),
    .A2(_0816_));
 sg13g2_xor2_1 _1722_ (.B(_0747_),
    .A(_0741_),
    .X(_0818_));
 sg13g2_nand2_1 _1723_ (.Y(_0819_),
    .A(_0817_),
    .B(_0818_));
 sg13g2_xnor2_1 _1724_ (.Y(_0820_),
    .A(_0817_),
    .B(_0818_));
 sg13g2_and4_1 _1725_ (.A(net284),
    .B(net285),
    .C(net298),
    .D(net296),
    .X(_0821_));
 sg13g2_nand2_1 _1726_ (.Y(_0822_),
    .A(net286),
    .B(net293));
 sg13g2_a22oi_1 _1727_ (.Y(_0823_),
    .B1(net295),
    .B2(net285),
    .A2(net298),
    .A1(net284));
 sg13g2_nor3_1 _1728_ (.A(_0821_),
    .B(_0822_),
    .C(_0823_),
    .Y(_0824_));
 sg13g2_or2_1 _1729_ (.X(_0825_),
    .B(_0824_),
    .A(_0821_));
 sg13g2_or2_1 _1730_ (.X(_0826_),
    .B(_0814_),
    .A(_0812_));
 sg13g2_o21ai_1 _1731_ (.B1(_0753_),
    .Y(_0827_),
    .A1(_0752_),
    .A2(_0754_));
 sg13g2_nor2b_1 _1732_ (.A(_0755_),
    .B_N(_0827_),
    .Y(_0828_));
 sg13g2_xnor2_1 _1733_ (.Y(_0829_),
    .A(_0826_),
    .B(_0828_));
 sg13g2_nor2b_1 _1734_ (.A(_0829_),
    .B_N(_0825_),
    .Y(_0830_));
 sg13g2_xor2_1 _1735_ (.B(_0829_),
    .A(_0825_),
    .X(_0831_));
 sg13g2_o21ai_1 _1736_ (.B1(_0819_),
    .Y(_0832_),
    .A1(_0820_),
    .A2(_0831_));
 sg13g2_xor2_1 _1737_ (.B(_0762_),
    .A(_0751_),
    .X(_0833_));
 sg13g2_nand2_1 _1738_ (.Y(_0834_),
    .A(_0832_),
    .B(_0833_));
 sg13g2_xnor2_1 _1739_ (.Y(_0835_),
    .A(_0832_),
    .B(_0833_));
 sg13g2_a22oi_1 _1740_ (.Y(_0836_),
    .B1(\perceptron1.we2[5] ),
    .B2(net319),
    .A2(net289),
    .A1(net286));
 sg13g2_nor2_1 _1741_ (.A(_0766_),
    .B(_0836_),
    .Y(_0837_));
 sg13g2_nand2_1 _1742_ (.Y(_0838_),
    .A(\perceptron1.we2[2] ),
    .B(net310));
 sg13g2_nand2_1 _1743_ (.Y(_0839_),
    .A(\perceptron1.we2[3] ),
    .B(net313));
 sg13g2_or2_1 _1744_ (.X(_0840_),
    .B(_0839_),
    .A(_0771_));
 sg13g2_xor2_1 _1745_ (.B(_0839_),
    .A(_0771_),
    .X(_0841_));
 sg13g2_nand2b_1 _1746_ (.Y(_0842_),
    .B(_0841_),
    .A_N(_0838_));
 sg13g2_xnor2_1 _1747_ (.Y(_0843_),
    .A(_0838_),
    .B(_0841_));
 sg13g2_nand2_1 _1748_ (.Y(_0844_),
    .A(_0837_),
    .B(_0843_));
 sg13g2_a21o_1 _1749_ (.A2(_0828_),
    .A1(_0826_),
    .B1(_0830_),
    .X(_0845_));
 sg13g2_xnor2_1 _1750_ (.Y(_0846_),
    .A(_0769_),
    .B(_0776_));
 sg13g2_nand2b_1 _1751_ (.Y(_0847_),
    .B(_0845_),
    .A_N(_0846_));
 sg13g2_xor2_1 _1752_ (.B(_0846_),
    .A(_0845_),
    .X(_0848_));
 sg13g2_xnor2_1 _1753_ (.Y(_0849_),
    .A(_0844_),
    .B(_0848_));
 sg13g2_o21ai_1 _1754_ (.B1(_0834_),
    .Y(_0850_),
    .A1(_0835_),
    .A2(_0849_));
 sg13g2_xor2_1 _1755_ (.B(_0784_),
    .A(_0783_),
    .X(_0851_));
 sg13g2_o21ai_1 _1756_ (.B1(_0847_),
    .Y(_0852_),
    .A1(_0844_),
    .A2(_0848_));
 sg13g2_xnor2_1 _1757_ (.Y(_0853_),
    .A(_0850_),
    .B(_0851_));
 sg13g2_nor2b_1 _1758_ (.A(_0853_),
    .B_N(_0852_),
    .Y(_0854_));
 sg13g2_a21o_1 _1759_ (.A2(_0851_),
    .A1(_0850_),
    .B1(_0854_),
    .X(_0855_));
 sg13g2_xor2_1 _1760_ (.B(_0788_),
    .A(_0787_),
    .X(_0856_));
 sg13g2_nand2b_1 _1761_ (.Y(_0857_),
    .B(_0855_),
    .A_N(_0856_));
 sg13g2_o21ai_1 _1762_ (.B1(_0510_),
    .Y(_0858_),
    .A1(_0507_),
    .A2(_0508_));
 sg13g2_inv_1 _1763_ (.Y(_0859_),
    .A(_0858_));
 sg13g2_xor2_1 _1764_ (.B(_0856_),
    .A(_0855_),
    .X(_0860_));
 sg13g2_o21ai_1 _1765_ (.B1(_0857_),
    .Y(_0861_),
    .A1(_0859_),
    .A2(_0860_));
 sg13g2_xor2_1 _1766_ (.B(_0794_),
    .A(_0793_),
    .X(_0862_));
 sg13g2_nor2b_1 _1767_ (.A(_0862_),
    .B_N(_0861_),
    .Y(_0863_));
 sg13g2_nand2_2 _1768_ (.Y(_0864_),
    .A(\perceptron1.we1[0] ),
    .B(net332));
 sg13g2_nor2_1 _1769_ (.A(_0732_),
    .B(_0864_),
    .Y(_0865_));
 sg13g2_xnor2_1 _1770_ (.Y(_0866_),
    .A(_0803_),
    .B(_0805_));
 sg13g2_nand2_1 _1771_ (.Y(_0867_),
    .A(_0865_),
    .B(_0866_));
 sg13g2_nand2_1 _1772_ (.Y(_0868_),
    .A(net301),
    .B(net284));
 sg13g2_and4_1 _1773_ (.A(net336),
    .B(net274),
    .C(net282),
    .D(net307),
    .X(_0869_));
 sg13g2_a22oi_1 _1774_ (.Y(_0870_),
    .B1(net282),
    .B2(net307),
    .A2(net274),
    .A1(net336));
 sg13g2_nor3_1 _1775_ (.A(_0868_),
    .B(_0869_),
    .C(_0870_),
    .Y(_0871_));
 sg13g2_o21ai_1 _1776_ (.B1(_0868_),
    .Y(_0872_),
    .A1(_0869_),
    .A2(_0870_));
 sg13g2_nand2b_1 _1777_ (.Y(_0873_),
    .B(_0872_),
    .A_N(_0871_));
 sg13g2_xnor2_1 _1778_ (.Y(_0874_),
    .A(_0865_),
    .B(_0866_));
 sg13g2_o21ai_1 _1779_ (.B1(_0867_),
    .Y(_0875_),
    .A1(_0873_),
    .A2(_0874_));
 sg13g2_xor2_1 _1780_ (.B(_0816_),
    .A(_0810_),
    .X(_0876_));
 sg13g2_nand2_1 _1781_ (.Y(_0877_),
    .A(_0875_),
    .B(_0876_));
 sg13g2_xnor2_1 _1782_ (.Y(_0878_),
    .A(_0875_),
    .B(_0876_));
 sg13g2_nor2_2 _1783_ (.A(_0342_),
    .B(_0353_),
    .Y(_0879_));
 sg13g2_nand3_1 _1784_ (.B(net295),
    .C(_0879_),
    .A(net285),
    .Y(_0880_));
 sg13g2_inv_1 _1785_ (.Y(_0881_),
    .A(_0880_));
 sg13g2_or2_1 _1786_ (.X(_0882_),
    .B(_0871_),
    .A(_0869_));
 sg13g2_o21ai_1 _1787_ (.B1(_0822_),
    .Y(_0883_),
    .A1(_0821_),
    .A2(_0823_));
 sg13g2_nor2b_1 _1788_ (.A(_0824_),
    .B_N(_0883_),
    .Y(_0884_));
 sg13g2_nand2_1 _1789_ (.Y(_0885_),
    .A(_0882_),
    .B(_0884_));
 sg13g2_xnor2_1 _1790_ (.Y(_0886_),
    .A(_0882_),
    .B(_0884_));
 sg13g2_xnor2_1 _1791_ (.Y(_0887_),
    .A(_0880_),
    .B(_0886_));
 sg13g2_o21ai_1 _1792_ (.B1(_0877_),
    .Y(_0888_),
    .A1(_0878_),
    .A2(_0887_));
 sg13g2_xor2_1 _1793_ (.B(_0831_),
    .A(_0820_),
    .X(_0889_));
 sg13g2_nand2_1 _1794_ (.Y(_0890_),
    .A(_0888_),
    .B(_0889_));
 sg13g2_xnor2_1 _1795_ (.Y(_0891_),
    .A(_0888_),
    .B(_0889_));
 sg13g2_nand2_1 _1796_ (.Y(_0892_),
    .A(net318),
    .B(\perceptron1.we2[4] ));
 sg13g2_and2_1 _1797_ (.A(\perceptron1.we2[1] ),
    .B(net310),
    .X(_0893_));
 sg13g2_nand2_1 _1798_ (.Y(_0894_),
    .A(\perceptron1.we2[2] ),
    .B(net316));
 sg13g2_or2_1 _1799_ (.X(_0895_),
    .B(_0894_),
    .A(_0839_));
 sg13g2_inv_1 _1800_ (.Y(_0896_),
    .A(_0895_));
 sg13g2_a22oi_1 _1801_ (.Y(_0897_),
    .B1(net313),
    .B2(\perceptron1.we2[2] ),
    .A2(net316),
    .A1(\perceptron1.we2[3] ));
 sg13g2_nor2_1 _1802_ (.A(_0896_),
    .B(_0897_),
    .Y(_0898_));
 sg13g2_xor2_1 _1803_ (.B(_0898_),
    .A(_0893_),
    .X(_0899_));
 sg13g2_nand2b_1 _1804_ (.Y(_0900_),
    .B(_0899_),
    .A_N(_0892_));
 sg13g2_xnor2_1 _1805_ (.Y(_0901_),
    .A(_0837_),
    .B(_0843_));
 sg13g2_o21ai_1 _1806_ (.B1(_0885_),
    .Y(_0902_),
    .A1(_0880_),
    .A2(_0886_));
 sg13g2_nand2b_1 _1807_ (.Y(_0903_),
    .B(_0902_),
    .A_N(_0901_));
 sg13g2_xor2_1 _1808_ (.B(_0902_),
    .A(_0901_),
    .X(_0904_));
 sg13g2_xnor2_1 _1809_ (.Y(_0905_),
    .A(_0900_),
    .B(_0904_));
 sg13g2_o21ai_1 _1810_ (.B1(_0890_),
    .Y(_0906_),
    .A1(_0891_),
    .A2(_0905_));
 sg13g2_xor2_1 _1811_ (.B(_0849_),
    .A(_0835_),
    .X(_0907_));
 sg13g2_nand2_1 _1812_ (.Y(_0908_),
    .A(_0906_),
    .B(_0907_));
 sg13g2_o21ai_1 _1813_ (.B1(_0903_),
    .Y(_0909_),
    .A1(_0900_),
    .A2(_0904_));
 sg13g2_inv_1 _1814_ (.Y(_0910_),
    .A(_0909_));
 sg13g2_xnor2_1 _1815_ (.Y(_0911_),
    .A(_0906_),
    .B(_0907_));
 sg13g2_o21ai_1 _1816_ (.B1(_0908_),
    .Y(_0912_),
    .A1(_0910_),
    .A2(_0911_));
 sg13g2_xor2_1 _1817_ (.B(_0853_),
    .A(_0852_),
    .X(_0913_));
 sg13g2_nor2b_1 _1818_ (.A(_0913_),
    .B_N(_0912_),
    .Y(_0914_));
 sg13g2_or2_1 _1819_ (.X(_0915_),
    .B(_0774_),
    .A(_0772_));
 sg13g2_xor2_1 _1820_ (.B(_0913_),
    .A(_0912_),
    .X(_0916_));
 sg13g2_nor2b_1 _1821_ (.A(_0916_),
    .B_N(_0915_),
    .Y(_0917_));
 sg13g2_xnor2_1 _1822_ (.Y(_0918_),
    .A(_0858_),
    .B(_0860_));
 sg13g2_o21ai_1 _1823_ (.B1(_0918_),
    .Y(_0919_),
    .A1(_0914_),
    .A2(_0917_));
 sg13g2_xor2_1 _1824_ (.B(_0862_),
    .A(_0861_),
    .X(_0920_));
 sg13g2_inv_1 _1825_ (.Y(_0921_),
    .A(_0920_));
 sg13g2_nor2_1 _1826_ (.A(_0919_),
    .B(_0920_),
    .Y(_0922_));
 sg13g2_nor2_1 _1827_ (.A(_0863_),
    .B(_0922_),
    .Y(_0923_));
 sg13g2_o21ai_1 _1828_ (.B1(_0800_),
    .Y(_0924_),
    .A1(_0863_),
    .A2(_0922_));
 sg13g2_nand2_1 _1829_ (.Y(_0925_),
    .A(_0731_),
    .B(_0797_));
 sg13g2_nand3_1 _1830_ (.B(_0924_),
    .C(_0925_),
    .A(_0730_),
    .Y(_0926_));
 sg13g2_a22oi_1 _1831_ (.Y(_0927_),
    .B1(\perceptron1.we1[1] ),
    .B2(net331),
    .A2(net328),
    .A1(\perceptron1.we1[0] ));
 sg13g2_nor2_1 _1832_ (.A(_0865_),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_and2_1 _1833_ (.A(net302),
    .B(net285),
    .X(_0929_));
 sg13g2_nand2_1 _1834_ (.Y(_0930_),
    .A(net308),
    .B(net284));
 sg13g2_nand2_1 _1835_ (.Y(_0931_),
    .A(\perceptron1.we1[2] ),
    .B(net337));
 sg13g2_nor2_1 _1836_ (.A(_0930_),
    .B(_0931_),
    .Y(_0932_));
 sg13g2_xor2_1 _1837_ (.B(_0931_),
    .A(_0930_),
    .X(_0933_));
 sg13g2_xor2_1 _1838_ (.B(_0933_),
    .A(_0929_),
    .X(_0934_));
 sg13g2_nand2_1 _1839_ (.Y(_0935_),
    .A(_0928_),
    .B(_0934_));
 sg13g2_xnor2_1 _1840_ (.Y(_0936_),
    .A(_0873_),
    .B(_0874_));
 sg13g2_or2_1 _1841_ (.X(_0937_),
    .B(_0936_),
    .A(_0935_));
 sg13g2_a22oi_1 _1842_ (.Y(_0938_),
    .B1(net286),
    .B2(net295),
    .A2(net298),
    .A1(net285));
 sg13g2_nor2_1 _1843_ (.A(_0881_),
    .B(_0938_),
    .Y(_0939_));
 sg13g2_a21oi_1 _1844_ (.A1(_0929_),
    .A2(_0933_),
    .Y(_0940_),
    .B1(_0932_));
 sg13g2_nand2b_1 _1845_ (.Y(_0941_),
    .B(_0939_),
    .A_N(_0940_));
 sg13g2_xor2_1 _1846_ (.B(_0940_),
    .A(_0939_),
    .X(_0942_));
 sg13g2_and2_1 _1847_ (.A(_0935_),
    .B(_0936_),
    .X(_0943_));
 sg13g2_xor2_1 _1848_ (.B(_0936_),
    .A(_0935_),
    .X(_0944_));
 sg13g2_o21ai_1 _1849_ (.B1(_0937_),
    .Y(_0945_),
    .A1(_0942_),
    .A2(_0943_));
 sg13g2_xor2_1 _1850_ (.B(_0887_),
    .A(_0878_),
    .X(_0946_));
 sg13g2_nand2_1 _1851_ (.Y(_0947_),
    .A(_0945_),
    .B(_0946_));
 sg13g2_xnor2_1 _1852_ (.Y(_0948_),
    .A(_0945_),
    .B(_0946_));
 sg13g2_nand2_1 _1853_ (.Y(_0949_),
    .A(net310),
    .B(\perceptron1.we2[0] ));
 sg13g2_nand2_2 _1854_ (.Y(_0950_),
    .A(net313),
    .B(\perceptron1.we2[1] ));
 sg13g2_xor2_1 _1855_ (.B(_0950_),
    .A(_0894_),
    .X(_0951_));
 sg13g2_nand2b_1 _1856_ (.Y(_0952_),
    .B(_0951_),
    .A_N(_0949_));
 sg13g2_xnor2_1 _1857_ (.Y(_0953_),
    .A(_0949_),
    .B(_0951_));
 sg13g2_nand3_1 _1858_ (.B(net318),
    .C(_0953_),
    .A(\perceptron1.we2[3] ),
    .Y(_0954_));
 sg13g2_inv_1 _1859_ (.Y(_0955_),
    .A(_0954_));
 sg13g2_xnor2_1 _1860_ (.Y(_0956_),
    .A(_0892_),
    .B(_0899_));
 sg13g2_nor2b_1 _1861_ (.A(_0941_),
    .B_N(_0956_),
    .Y(_0957_));
 sg13g2_xnor2_1 _1862_ (.Y(_0958_),
    .A(_0941_),
    .B(_0956_));
 sg13g2_xnor2_1 _1863_ (.Y(_0959_),
    .A(_0954_),
    .B(_0958_));
 sg13g2_inv_1 _1864_ (.Y(_0960_),
    .A(_0959_));
 sg13g2_o21ai_1 _1865_ (.B1(_0947_),
    .Y(_0961_),
    .A1(_0948_),
    .A2(_0960_));
 sg13g2_xor2_1 _1866_ (.B(_0905_),
    .A(_0891_),
    .X(_0962_));
 sg13g2_nand2_1 _1867_ (.Y(_0963_),
    .A(_0961_),
    .B(_0962_));
 sg13g2_a21oi_1 _1868_ (.A1(_0955_),
    .A2(_0958_),
    .Y(_0964_),
    .B1(_0957_));
 sg13g2_xnor2_1 _1869_ (.Y(_0965_),
    .A(_0961_),
    .B(_0962_));
 sg13g2_o21ai_1 _1870_ (.B1(_0963_),
    .Y(_0966_),
    .A1(_0964_),
    .A2(_0965_));
 sg13g2_xnor2_1 _1871_ (.Y(_0967_),
    .A(_0910_),
    .B(_0911_));
 sg13g2_nand2b_1 _1872_ (.Y(_0968_),
    .B(_0966_),
    .A_N(_0967_));
 sg13g2_and2_1 _1873_ (.A(_0840_),
    .B(_0842_),
    .X(_0969_));
 sg13g2_xor2_1 _1874_ (.B(_0967_),
    .A(_0966_),
    .X(_0970_));
 sg13g2_o21ai_1 _1875_ (.B1(_0968_),
    .Y(_0971_),
    .A1(_0969_),
    .A2(_0970_));
 sg13g2_xor2_1 _1876_ (.B(_0916_),
    .A(_0915_),
    .X(_0972_));
 sg13g2_nor2b_1 _1877_ (.A(_0972_),
    .B_N(_0971_),
    .Y(_0973_));
 sg13g2_nand2_1 _1878_ (.Y(_0974_),
    .A(net301),
    .B(net286));
 sg13g2_nand2_1 _1879_ (.Y(_0975_),
    .A(net308),
    .B(net285));
 sg13g2_nand2_1 _1880_ (.Y(_0976_),
    .A(\perceptron1.we1[1] ),
    .B(net337));
 sg13g2_nor2_1 _1881_ (.A(_0975_),
    .B(_0976_),
    .Y(_0977_));
 sg13g2_xor2_1 _1882_ (.B(_0976_),
    .A(_0975_),
    .X(_0978_));
 sg13g2_nor2b_1 _1883_ (.A(_0974_),
    .B_N(_0978_),
    .Y(_0979_));
 sg13g2_xnor2_1 _1884_ (.Y(_0980_),
    .A(_0974_),
    .B(_0978_));
 sg13g2_nand2b_1 _1885_ (.Y(_0981_),
    .B(_0980_),
    .A_N(_0864_));
 sg13g2_xnor2_1 _1886_ (.Y(_0982_),
    .A(_0928_),
    .B(_0934_));
 sg13g2_nor2_1 _1887_ (.A(_0981_),
    .B(_0982_),
    .Y(_0983_));
 sg13g2_nor2_1 _1888_ (.A(_0977_),
    .B(_0979_),
    .Y(_0984_));
 sg13g2_o21ai_1 _1889_ (.B1(_0879_),
    .Y(_0985_),
    .A1(_0977_),
    .A2(_0979_));
 sg13g2_xnor2_1 _1890_ (.Y(_0986_),
    .A(_0879_),
    .B(_0984_));
 sg13g2_xor2_1 _1891_ (.B(_0982_),
    .A(_0981_),
    .X(_0987_));
 sg13g2_a21oi_1 _1892_ (.A1(_0986_),
    .A2(_0987_),
    .Y(_0988_),
    .B1(_0983_));
 sg13g2_xnor2_1 _1893_ (.Y(_0989_),
    .A(_0942_),
    .B(_0944_));
 sg13g2_nor2b_1 _1894_ (.A(_0988_),
    .B_N(_0989_),
    .Y(_0990_));
 sg13g2_nand2_1 _1895_ (.Y(_0991_),
    .A(net318),
    .B(\perceptron1.we2[2] ));
 sg13g2_a22oi_1 _1896_ (.Y(_0992_),
    .B1(\perceptron1.we2[0] ),
    .B2(net312),
    .A2(\perceptron1.we2[1] ),
    .A1(net316));
 sg13g2_nand2_2 _1897_ (.Y(_0993_),
    .A(net316),
    .B(\perceptron1.we2[0] ));
 sg13g2_nor2_2 _1898_ (.A(_0950_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_or2_1 _1899_ (.X(_0995_),
    .B(_0993_),
    .A(_0950_));
 sg13g2_nor3_2 _1900_ (.A(_0991_),
    .B(_0992_),
    .C(_0994_),
    .Y(_0996_));
 sg13g2_a21o_1 _1901_ (.A2(net318),
    .A1(\perceptron1.we2[3] ),
    .B1(_0953_),
    .X(_0997_));
 sg13g2_nand2_1 _1902_ (.Y(_0998_),
    .A(_0954_),
    .B(_0997_));
 sg13g2_nor2_1 _1903_ (.A(_0985_),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_xor2_1 _1904_ (.B(_0998_),
    .A(_0985_),
    .X(_1000_));
 sg13g2_xnor2_1 _1905_ (.Y(_1001_),
    .A(_0996_),
    .B(_1000_));
 sg13g2_inv_1 _1906_ (.Y(_1002_),
    .A(_1001_));
 sg13g2_xnor2_1 _1907_ (.Y(_1003_),
    .A(_0988_),
    .B(_0989_));
 sg13g2_a21oi_1 _1908_ (.A1(_1002_),
    .A2(_1003_),
    .Y(_1004_),
    .B1(_0990_));
 sg13g2_xnor2_1 _1909_ (.Y(_1005_),
    .A(_0948_),
    .B(_0959_));
 sg13g2_nand2b_1 _1910_ (.Y(_1006_),
    .B(_1005_),
    .A_N(_1004_));
 sg13g2_a21oi_1 _1911_ (.A1(_0996_),
    .A2(_1000_),
    .Y(_1007_),
    .B1(_0999_));
 sg13g2_xnor2_1 _1912_ (.Y(_1008_),
    .A(_1004_),
    .B(_1005_));
 sg13g2_nand2b_1 _1913_ (.Y(_1009_),
    .B(_1008_),
    .A_N(_1007_));
 sg13g2_nand2_1 _1914_ (.Y(_1010_),
    .A(_1006_),
    .B(_1009_));
 sg13g2_xor2_1 _1915_ (.B(_0965_),
    .A(_0964_),
    .X(_1011_));
 sg13g2_nand2_1 _1916_ (.Y(_1012_),
    .A(_1010_),
    .B(_1011_));
 sg13g2_a21oi_1 _1917_ (.A1(_0893_),
    .A2(_0898_),
    .Y(_1013_),
    .B1(_0896_));
 sg13g2_xnor2_1 _1918_ (.Y(_1014_),
    .A(_1010_),
    .B(_1011_));
 sg13g2_o21ai_1 _1919_ (.B1(_1012_),
    .Y(_1015_),
    .A1(_1013_),
    .A2(_1014_));
 sg13g2_xor2_1 _1920_ (.B(_0970_),
    .A(_0969_),
    .X(_1016_));
 sg13g2_nand2_1 _1921_ (.Y(_1017_),
    .A(_1015_),
    .B(_1016_));
 sg13g2_nand4_1 _1922_ (.B(net337),
    .C(net308),
    .A(\perceptron1.we1[0] ),
    .Y(_1018_),
    .D(net286));
 sg13g2_xnor2_1 _1923_ (.Y(_1019_),
    .A(_0864_),
    .B(_0980_));
 sg13g2_nand2b_1 _1924_ (.Y(_1020_),
    .B(_1019_),
    .A_N(_1018_));
 sg13g2_xnor2_1 _1925_ (.Y(_1021_),
    .A(_0986_),
    .B(_0987_));
 sg13g2_nor2_1 _1926_ (.A(_1020_),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_nand2_1 _1927_ (.Y(_1023_),
    .A(net318),
    .B(\perceptron1.we2[1] ));
 sg13g2_or2_1 _1928_ (.X(_1024_),
    .B(_1023_),
    .A(_0993_));
 sg13g2_o21ai_1 _1929_ (.B1(_0991_),
    .Y(_1025_),
    .A1(_0992_),
    .A2(_0994_));
 sg13g2_nor2b_1 _1930_ (.A(_0996_),
    .B_N(_1025_),
    .Y(_1026_));
 sg13g2_nor2b_1 _1931_ (.A(_1024_),
    .B_N(_1026_),
    .Y(_1027_));
 sg13g2_xnor2_1 _1932_ (.Y(_1028_),
    .A(_1024_),
    .B(_1026_));
 sg13g2_xnor2_1 _1933_ (.Y(_1029_),
    .A(_1020_),
    .B(_1021_));
 sg13g2_inv_1 _1934_ (.Y(_1030_),
    .A(_1029_));
 sg13g2_a21oi_1 _1935_ (.A1(_1028_),
    .A2(_1030_),
    .Y(_1031_),
    .B1(_1022_));
 sg13g2_xnor2_1 _1936_ (.Y(_1032_),
    .A(_1001_),
    .B(_1003_));
 sg13g2_nor2b_1 _1937_ (.A(_1031_),
    .B_N(_1032_),
    .Y(_1033_));
 sg13g2_xnor2_1 _1938_ (.Y(_1034_),
    .A(_1031_),
    .B(_1032_));
 sg13g2_a21oi_1 _1939_ (.A1(_1027_),
    .A2(_1034_),
    .Y(_1035_),
    .B1(_1033_));
 sg13g2_xnor2_1 _1940_ (.Y(_1036_),
    .A(_1007_),
    .B(_1008_));
 sg13g2_nor2b_1 _1941_ (.A(_1035_),
    .B_N(_1036_),
    .Y(_1037_));
 sg13g2_o21ai_1 _1942_ (.B1(_0952_),
    .Y(_1038_),
    .A1(_0894_),
    .A2(_0950_));
 sg13g2_xnor2_1 _1943_ (.Y(_1039_),
    .A(_1035_),
    .B(_1036_));
 sg13g2_a21o_1 _1944_ (.A2(_1039_),
    .A1(_1038_),
    .B1(_1037_),
    .X(_1040_));
 sg13g2_xnor2_1 _1945_ (.Y(_1041_),
    .A(_1013_),
    .B(_1014_));
 sg13g2_nand2b_1 _1946_ (.Y(_1042_),
    .B(_1041_),
    .A_N(_1040_));
 sg13g2_xor2_1 _1947_ (.B(_1039_),
    .A(_1038_),
    .X(_1043_));
 sg13g2_xor2_1 _1948_ (.B(_1023_),
    .A(_0993_),
    .X(_1044_));
 sg13g2_xnor2_1 _1949_ (.Y(_1045_),
    .A(_1018_),
    .B(_1019_));
 sg13g2_nand2_1 _1950_ (.Y(_1046_),
    .A(_1044_),
    .B(_1045_));
 sg13g2_xor2_1 _1951_ (.B(_1029_),
    .A(_1028_),
    .X(_1047_));
 sg13g2_nor2_1 _1952_ (.A(_1046_),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_xor2_1 _1953_ (.B(_1034_),
    .A(_1027_),
    .X(_1049_));
 sg13g2_nand2_1 _1954_ (.Y(_1050_),
    .A(_1048_),
    .B(_1049_));
 sg13g2_xnor2_1 _1955_ (.Y(_1051_),
    .A(_1048_),
    .B(_1049_));
 sg13g2_o21ai_1 _1956_ (.B1(_1050_),
    .Y(_1052_),
    .A1(_0995_),
    .A2(_1051_));
 sg13g2_nand2_1 _1957_ (.Y(_1053_),
    .A(_1043_),
    .B(_1052_));
 sg13g2_xor2_1 _1958_ (.B(_1052_),
    .A(_1043_),
    .X(_1054_));
 sg13g2_xnor2_1 _1959_ (.Y(_1055_),
    .A(_0994_),
    .B(_1051_));
 sg13g2_nor2_1 _1960_ (.A(_1044_),
    .B(_1045_),
    .Y(_1056_));
 sg13g2_a22oi_1 _1961_ (.Y(_1057_),
    .B1(net308),
    .B2(net286),
    .A2(net337),
    .A1(\perceptron1.we1[0] ));
 sg13g2_inv_1 _1962_ (.Y(_1058_),
    .A(_1057_));
 sg13g2_nand2_1 _1963_ (.Y(_1059_),
    .A(_1018_),
    .B(_1058_));
 sg13g2_nand3_1 _1964_ (.B(\perceptron1.we2[0] ),
    .C(_1046_),
    .A(net318),
    .Y(_1060_));
 sg13g2_nor4_2 _1965_ (.A(_1047_),
    .B(_1056_),
    .C(_1059_),
    .Y(_1061_),
    .D(_1060_));
 sg13g2_nand3_1 _1966_ (.B(_1055_),
    .C(_1061_),
    .A(_1054_),
    .Y(_1062_));
 sg13g2_nand2b_1 _1967_ (.Y(_1063_),
    .B(_1040_),
    .A_N(_1041_));
 sg13g2_nand3_1 _1968_ (.B(_1062_),
    .C(_1063_),
    .A(_1053_),
    .Y(_1064_));
 sg13g2_xor2_1 _1969_ (.B(_1016_),
    .A(_1015_),
    .X(_1065_));
 sg13g2_nand3_1 _1970_ (.B(_1064_),
    .C(_1065_),
    .A(_1042_),
    .Y(_1066_));
 sg13g2_xor2_1 _1971_ (.B(_0972_),
    .A(_0971_),
    .X(_1067_));
 sg13g2_a21oi_1 _1972_ (.A1(_1017_),
    .A2(_1066_),
    .Y(_1068_),
    .B1(_1067_));
 sg13g2_or2_1 _1973_ (.X(_1069_),
    .B(_1068_),
    .A(_0973_));
 sg13g2_nor2_1 _1974_ (.A(_0926_),
    .B(_1069_),
    .Y(_1070_));
 sg13g2_o21ai_1 _1975_ (.B1(_0686_),
    .Y(_1071_),
    .A1(_0687_),
    .A2(_0698_));
 sg13g2_o21ai_1 _1976_ (.B1(_0677_),
    .Y(_1072_),
    .A1(_0678_),
    .A2(_0684_));
 sg13g2_o21ai_1 _1977_ (.B1(_0673_),
    .Y(_1073_),
    .A1(_0671_),
    .A2(_0674_));
 sg13g2_nand2_1 _1978_ (.Y(_1074_),
    .A(net330),
    .B(net272));
 sg13g2_nand2_1 _1979_ (.Y(_1075_),
    .A(net321),
    .B(\perceptron1.we1[10] ));
 sg13g2_and4_1 _1980_ (.A(net321),
    .B(net325),
    .C(\perceptron1.we1[10] ),
    .D(\perceptron1.we1[9] ),
    .X(_1076_));
 sg13g2_a22oi_1 _1981_ (.Y(_1077_),
    .B1(\perceptron1.we1[9] ),
    .B2(net321),
    .A2(\perceptron1.we1[10] ),
    .A1(net325));
 sg13g2_nor3_1 _1982_ (.A(_1074_),
    .B(_1076_),
    .C(_1077_),
    .Y(_1078_));
 sg13g2_o21ai_1 _1983_ (.B1(_1074_),
    .Y(_1079_),
    .A1(_1076_),
    .A2(_1077_));
 sg13g2_nor2b_1 _1984_ (.A(_1078_),
    .B_N(_1079_),
    .Y(_1080_));
 sg13g2_nand2_1 _1985_ (.Y(_1081_),
    .A(_1073_),
    .B(_1080_));
 sg13g2_xnor2_1 _1986_ (.Y(_1082_),
    .A(_1073_),
    .B(_1080_));
 sg13g2_nand2_1 _1987_ (.Y(_1083_),
    .A(net300),
    .B(\perceptron1.we3[11] ));
 sg13g2_and4_1 _1988_ (.A(net333),
    .B(net306),
    .C(\perceptron1.we1[12] ),
    .D(\perceptron1.we3[12] ),
    .X(_1084_));
 sg13g2_a22oi_1 _1989_ (.Y(_1085_),
    .B1(\perceptron1.we3[12] ),
    .B2(net304),
    .A2(\perceptron1.we1[12] ),
    .A1(net334));
 sg13g2_nor3_1 _1990_ (.A(_1083_),
    .B(_1084_),
    .C(_1085_),
    .Y(_1086_));
 sg13g2_o21ai_1 _1991_ (.B1(_1083_),
    .Y(_1087_),
    .A1(_1084_),
    .A2(_1085_));
 sg13g2_nand2b_1 _1992_ (.Y(_1088_),
    .B(_1087_),
    .A_N(_1086_));
 sg13g2_xor2_1 _1993_ (.B(_1088_),
    .A(_1082_),
    .X(_1089_));
 sg13g2_nand2_1 _1994_ (.Y(_1090_),
    .A(_1072_),
    .B(_1089_));
 sg13g2_xnor2_1 _1995_ (.Y(_1091_),
    .A(_1072_),
    .B(_1089_));
 sg13g2_o21ai_1 _1996_ (.B1(_0693_),
    .Y(_1092_),
    .A1(_0690_),
    .A2(_0694_));
 sg13g2_or2_1 _1997_ (.X(_1093_),
    .B(_0682_),
    .A(_0680_));
 sg13g2_nand2_1 _1998_ (.Y(_1094_),
    .A(net292),
    .B(\perceptron1.we3[8] ));
 sg13g2_nand2_1 _1999_ (.Y(_1095_),
    .A(net294),
    .B(net275));
 sg13g2_nand2_1 _2000_ (.Y(_1096_),
    .A(net297),
    .B(net275));
 sg13g2_or2_1 _2001_ (.X(_1097_),
    .B(_1095_),
    .A(_0692_));
 sg13g2_xnor2_1 _2002_ (.Y(_1098_),
    .A(_0691_),
    .B(_1096_));
 sg13g2_xor2_1 _2003_ (.B(_1098_),
    .A(_1094_),
    .X(_1099_));
 sg13g2_xnor2_1 _2004_ (.Y(_1100_),
    .A(_1093_),
    .B(_1099_));
 sg13g2_nor2b_1 _2005_ (.A(_1100_),
    .B_N(_1092_),
    .Y(_1101_));
 sg13g2_xor2_1 _2006_ (.B(_1100_),
    .A(_1092_),
    .X(_1102_));
 sg13g2_xor2_1 _2007_ (.B(_1102_),
    .A(_1091_),
    .X(_1103_));
 sg13g2_nand2_1 _2008_ (.Y(_1104_),
    .A(_1071_),
    .B(_1103_));
 sg13g2_xnor2_1 _2009_ (.Y(_1105_),
    .A(_1071_),
    .B(_1103_));
 sg13g2_a21o_1 _2010_ (.A2(_0710_),
    .A1(_0704_),
    .B1(_0717_),
    .X(_1106_));
 sg13g2_a21o_1 _2011_ (.A2(_0695_),
    .A1(_0689_),
    .B1(_0697_),
    .X(_1107_));
 sg13g2_o21ai_1 _2012_ (.B1(_0709_),
    .Y(_1108_),
    .A1(_0637_),
    .A2(_0707_));
 sg13g2_nand2_1 _2013_ (.Y(_1109_),
    .A(net320),
    .B(\perceptron1.we2[12] ));
 sg13g2_nand2_1 _2014_ (.Y(_1110_),
    .A(net278),
    .B(net287));
 sg13g2_nand2_1 _2015_ (.Y(_1111_),
    .A(net278),
    .B(net289));
 sg13g2_xor2_1 _2016_ (.B(_1111_),
    .A(_0706_),
    .X(_1112_));
 sg13g2_nand2b_1 _2017_ (.Y(_1113_),
    .B(_1112_),
    .A_N(_1109_));
 sg13g2_xnor2_1 _2018_ (.Y(_1114_),
    .A(_1109_),
    .B(_1112_));
 sg13g2_xnor2_1 _2019_ (.Y(_1115_),
    .A(_1108_),
    .B(_1114_));
 sg13g2_nand2_1 _2020_ (.Y(_1116_),
    .A(net311),
    .B(\perceptron1.we2[9] ));
 sg13g2_nand2_2 _2021_ (.Y(_1117_),
    .A(net314),
    .B(\perceptron1.we2[11] ));
 sg13g2_nor2_1 _2022_ (.A(_0713_),
    .B(_1117_),
    .Y(_1118_));
 sg13g2_or2_1 _2023_ (.X(_1119_),
    .B(_1117_),
    .A(_0713_));
 sg13g2_a22oi_1 _2024_ (.Y(_1120_),
    .B1(\perceptron1.we2[10] ),
    .B2(net314),
    .A2(\perceptron1.we2[11] ),
    .A1(net317));
 sg13g2_nor2_1 _2025_ (.A(_1118_),
    .B(_1120_),
    .Y(_1121_));
 sg13g2_xnor2_1 _2026_ (.Y(_1122_),
    .A(_1116_),
    .B(_1121_));
 sg13g2_nor2b_1 _2027_ (.A(_1115_),
    .B_N(_1122_),
    .Y(_1123_));
 sg13g2_xnor2_1 _2028_ (.Y(_1124_),
    .A(_1115_),
    .B(_1122_));
 sg13g2_xnor2_1 _2029_ (.Y(_1125_),
    .A(_1107_),
    .B(_1124_));
 sg13g2_nor2b_1 _2030_ (.A(_1125_),
    .B_N(_1106_),
    .Y(_1126_));
 sg13g2_xor2_1 _2031_ (.B(_1125_),
    .A(_1106_),
    .X(_1127_));
 sg13g2_o21ai_1 _2032_ (.B1(_1104_),
    .Y(_1128_),
    .A1(_1105_),
    .A2(_1127_));
 sg13g2_o21ai_1 _2033_ (.B1(_1090_),
    .Y(_1129_),
    .A1(_1091_),
    .A2(_1102_));
 sg13g2_o21ai_1 _2034_ (.B1(_1081_),
    .Y(_1130_),
    .A1(_1082_),
    .A2(_1088_));
 sg13g2_or2_1 _2035_ (.X(_1131_),
    .B(_1078_),
    .A(_1076_));
 sg13g2_nand2_1 _2036_ (.Y(_1132_),
    .A(net330),
    .B(\perceptron1.we1[12] ));
 sg13g2_nand2_1 _2037_ (.Y(_1133_),
    .A(net325),
    .B(\perceptron1.we1[11] ));
 sg13g2_or2_1 _2038_ (.X(_1134_),
    .B(_1133_),
    .A(_1075_));
 sg13g2_and2_1 _2039_ (.A(_1075_),
    .B(_1133_),
    .X(_1135_));
 sg13g2_xor2_1 _2040_ (.B(_1133_),
    .A(_1075_),
    .X(_1136_));
 sg13g2_xnor2_1 _2041_ (.Y(_1137_),
    .A(_1132_),
    .B(_1136_));
 sg13g2_nand2_1 _2042_ (.Y(_1138_),
    .A(_1131_),
    .B(_1137_));
 sg13g2_xnor2_1 _2043_ (.Y(_1139_),
    .A(_1131_),
    .B(_1137_));
 sg13g2_nand2_1 _2044_ (.Y(_1140_),
    .A(net300),
    .B(\perceptron1.we3[12] ));
 sg13g2_and4_1 _2045_ (.A(net333),
    .B(net306),
    .C(\perceptron1.we1[13] ),
    .D(\perceptron1.we3[13] ),
    .X(_1141_));
 sg13g2_a22oi_1 _2046_ (.Y(_1142_),
    .B1(\perceptron1.we3[13] ),
    .B2(net306),
    .A2(\perceptron1.we1[13] ),
    .A1(net333));
 sg13g2_nor3_1 _2047_ (.A(_1140_),
    .B(_1141_),
    .C(_1142_),
    .Y(_1143_));
 sg13g2_o21ai_1 _2048_ (.B1(_1140_),
    .Y(_1144_),
    .A1(_1141_),
    .A2(_1142_));
 sg13g2_nand2b_1 _2049_ (.Y(_1145_),
    .B(_1144_),
    .A_N(_1143_));
 sg13g2_xor2_1 _2050_ (.B(_1145_),
    .A(_1139_),
    .X(_1146_));
 sg13g2_nand2_1 _2051_ (.Y(_1147_),
    .A(_1130_),
    .B(_1146_));
 sg13g2_xnor2_1 _2052_ (.Y(_1148_),
    .A(_1130_),
    .B(_1146_));
 sg13g2_o21ai_1 _2053_ (.B1(_1097_),
    .Y(_1149_),
    .A1(_1094_),
    .A2(_1098_));
 sg13g2_or2_1 _2054_ (.X(_1150_),
    .B(_1086_),
    .A(_1084_));
 sg13g2_nand2_1 _2055_ (.Y(_1151_),
    .A(net292),
    .B(net276));
 sg13g2_nand2_1 _2056_ (.Y(_1152_),
    .A(net294),
    .B(\perceptron1.we3[11] ));
 sg13g2_nand2_1 _2057_ (.Y(_1153_),
    .A(net297),
    .B(\perceptron1.we3[11] ));
 sg13g2_or2_1 _2058_ (.X(_1154_),
    .B(_1152_),
    .A(_1096_));
 sg13g2_xnor2_1 _2059_ (.Y(_1155_),
    .A(_1095_),
    .B(_1153_));
 sg13g2_xor2_1 _2060_ (.B(_1155_),
    .A(_1151_),
    .X(_1156_));
 sg13g2_xnor2_1 _2061_ (.Y(_1157_),
    .A(_1150_),
    .B(_1156_));
 sg13g2_nor2b_1 _2062_ (.A(_1157_),
    .B_N(_1149_),
    .Y(_1158_));
 sg13g2_xor2_1 _2063_ (.B(_1157_),
    .A(_1149_),
    .X(_1159_));
 sg13g2_xor2_1 _2064_ (.B(_1159_),
    .A(_1148_),
    .X(_1160_));
 sg13g2_nand2_1 _2065_ (.Y(_1161_),
    .A(_1129_),
    .B(_1160_));
 sg13g2_xnor2_1 _2066_ (.Y(_1162_),
    .A(_1129_),
    .B(_1160_));
 sg13g2_a21o_1 _2067_ (.A2(_1114_),
    .A1(_1108_),
    .B1(_1123_),
    .X(_1163_));
 sg13g2_a21o_1 _2068_ (.A2(_1099_),
    .A1(_1093_),
    .B1(_1101_),
    .X(_1164_));
 sg13g2_o21ai_1 _2069_ (.B1(_1113_),
    .Y(_1165_),
    .A1(_0706_),
    .A2(_1111_));
 sg13g2_nand2_1 _2070_ (.Y(_1166_),
    .A(net320),
    .B(\perceptron1.we2[13] ));
 sg13g2_nand2_1 _2071_ (.Y(_1167_),
    .A(net289),
    .B(\perceptron1.we3[8] ));
 sg13g2_xor2_1 _2072_ (.B(_1167_),
    .A(_1110_),
    .X(_1168_));
 sg13g2_nand2b_1 _2073_ (.Y(_1169_),
    .B(_1168_),
    .A_N(_1166_));
 sg13g2_xnor2_1 _2074_ (.Y(_1170_),
    .A(_1166_),
    .B(_1168_));
 sg13g2_xnor2_1 _2075_ (.Y(_1171_),
    .A(_1165_),
    .B(_1170_));
 sg13g2_nand2_1 _2076_ (.Y(_1172_),
    .A(net311),
    .B(\perceptron1.we2[10] ));
 sg13g2_nand2_1 _2077_ (.Y(_1173_),
    .A(net317),
    .B(\perceptron1.we2[12] ));
 sg13g2_xor2_1 _2078_ (.B(_1173_),
    .A(_1117_),
    .X(_1174_));
 sg13g2_nand2b_1 _2079_ (.Y(_1175_),
    .B(_1174_),
    .A_N(_1172_));
 sg13g2_xnor2_1 _2080_ (.Y(_1176_),
    .A(_1172_),
    .B(_1174_));
 sg13g2_nor2b_1 _2081_ (.A(_1171_),
    .B_N(_1176_),
    .Y(_1177_));
 sg13g2_xnor2_1 _2082_ (.Y(_1178_),
    .A(_1171_),
    .B(_1176_));
 sg13g2_xnor2_1 _2083_ (.Y(_1179_),
    .A(_1164_),
    .B(_1178_));
 sg13g2_nor2b_1 _2084_ (.A(_1179_),
    .B_N(_1163_),
    .Y(_1180_));
 sg13g2_xor2_1 _2085_ (.B(_1179_),
    .A(_1163_),
    .X(_1181_));
 sg13g2_xor2_1 _2086_ (.B(_1181_),
    .A(_1162_),
    .X(_1182_));
 sg13g2_a21o_1 _2087_ (.A2(_1124_),
    .A1(_1107_),
    .B1(_1126_),
    .X(_1183_));
 sg13g2_xnor2_1 _2088_ (.Y(_1184_),
    .A(_1128_),
    .B(_1182_));
 sg13g2_nor2b_1 _2089_ (.A(_1184_),
    .B_N(_1183_),
    .Y(_1185_));
 sg13g2_a21o_1 _2090_ (.A2(_1182_),
    .A1(_1128_),
    .B1(_1185_),
    .X(_1186_));
 sg13g2_a21o_1 _2091_ (.A2(_1178_),
    .A1(_1164_),
    .B1(_1180_),
    .X(_1187_));
 sg13g2_o21ai_1 _2092_ (.B1(_1161_),
    .Y(_1188_),
    .A1(_1162_),
    .A2(_1181_));
 sg13g2_o21ai_1 _2093_ (.B1(_1147_),
    .Y(_1189_),
    .A1(_1148_),
    .A2(_1159_));
 sg13g2_o21ai_1 _2094_ (.B1(_1138_),
    .Y(_1190_),
    .A1(_1139_),
    .A2(_1145_));
 sg13g2_o21ai_1 _2095_ (.B1(_1134_),
    .Y(_1191_),
    .A1(_1132_),
    .A2(_1135_));
 sg13g2_nand2_1 _2096_ (.Y(_1192_),
    .A(net330),
    .B(\perceptron1.we1[13] ));
 sg13g2_nand2_1 _2097_ (.Y(_1193_),
    .A(net321),
    .B(\perceptron1.we1[12] ));
 sg13g2_and4_1 _2098_ (.A(net321),
    .B(net325),
    .C(\perceptron1.we1[12] ),
    .D(net272),
    .X(_1194_));
 sg13g2_a22oi_1 _2099_ (.Y(_1195_),
    .B1(net272),
    .B2(net321),
    .A2(\perceptron1.we1[12] ),
    .A1(net325));
 sg13g2_nor3_1 _2100_ (.A(_1192_),
    .B(_1194_),
    .C(_1195_),
    .Y(_1196_));
 sg13g2_o21ai_1 _2101_ (.B1(_1192_),
    .Y(_1197_),
    .A1(_1194_),
    .A2(_1195_));
 sg13g2_nor2b_1 _2102_ (.A(_1196_),
    .B_N(_1197_),
    .Y(_1198_));
 sg13g2_nand2_1 _2103_ (.Y(_1199_),
    .A(_1191_),
    .B(_1198_));
 sg13g2_xnor2_1 _2104_ (.Y(_1200_),
    .A(_1191_),
    .B(_1198_));
 sg13g2_nand2_1 _2105_ (.Y(_1201_),
    .A(net300),
    .B(\perceptron1.we3[13] ));
 sg13g2_and4_1 _2106_ (.A(net333),
    .B(net306),
    .C(\perceptron1.we1[14] ),
    .D(\perceptron1.we3[14] ),
    .X(_1202_));
 sg13g2_a22oi_1 _2107_ (.Y(_1203_),
    .B1(\perceptron1.we3[14] ),
    .B2(net306),
    .A2(\perceptron1.we1[14] ),
    .A1(net333));
 sg13g2_nor3_1 _2108_ (.A(_1201_),
    .B(_1202_),
    .C(_1203_),
    .Y(_1204_));
 sg13g2_o21ai_1 _2109_ (.B1(_1201_),
    .Y(_1205_),
    .A1(_1202_),
    .A2(_1203_));
 sg13g2_nor2b_1 _2110_ (.A(_1204_),
    .B_N(_1205_),
    .Y(_1206_));
 sg13g2_nand2b_1 _2111_ (.Y(_1207_),
    .B(_1206_),
    .A_N(_1200_));
 sg13g2_xnor2_1 _2112_ (.Y(_1208_),
    .A(_1200_),
    .B(_1206_));
 sg13g2_nand2_1 _2113_ (.Y(_1209_),
    .A(_1190_),
    .B(_1208_));
 sg13g2_xnor2_1 _2114_ (.Y(_1210_),
    .A(_1190_),
    .B(_1208_));
 sg13g2_o21ai_1 _2115_ (.B1(_1154_),
    .Y(_1211_),
    .A1(_1151_),
    .A2(_1155_));
 sg13g2_or2_1 _2116_ (.X(_1212_),
    .B(_1143_),
    .A(_1141_));
 sg13g2_nand2_1 _2117_ (.Y(_1213_),
    .A(net292),
    .B(net275));
 sg13g2_nand2_1 _2118_ (.Y(_1214_),
    .A(net294),
    .B(\perceptron1.we3[12] ));
 sg13g2_nand2_1 _2119_ (.Y(_1215_),
    .A(net297),
    .B(\perceptron1.we3[12] ));
 sg13g2_xor2_1 _2120_ (.B(_1215_),
    .A(_1152_),
    .X(_1216_));
 sg13g2_nand2b_1 _2121_ (.Y(_1217_),
    .B(_1216_),
    .A_N(_1213_));
 sg13g2_xnor2_1 _2122_ (.Y(_1218_),
    .A(_1213_),
    .B(_1216_));
 sg13g2_xnor2_1 _2123_ (.Y(_1219_),
    .A(_1212_),
    .B(_1218_));
 sg13g2_nor2b_1 _2124_ (.A(_1219_),
    .B_N(_1211_),
    .Y(_1220_));
 sg13g2_xor2_1 _2125_ (.B(_1219_),
    .A(_1211_),
    .X(_1221_));
 sg13g2_xor2_1 _2126_ (.B(_1221_),
    .A(_1210_),
    .X(_1222_));
 sg13g2_nand2_1 _2127_ (.Y(_1223_),
    .A(_1189_),
    .B(_1222_));
 sg13g2_xnor2_1 _2128_ (.Y(_1224_),
    .A(_1189_),
    .B(_1222_));
 sg13g2_a21o_1 _2129_ (.A2(_1170_),
    .A1(_1165_),
    .B1(_1177_),
    .X(_1225_));
 sg13g2_a21o_1 _2130_ (.A2(_1156_),
    .A1(_1150_),
    .B1(_1158_),
    .X(_1226_));
 sg13g2_o21ai_1 _2131_ (.B1(_1169_),
    .Y(_1227_),
    .A1(_1110_),
    .A2(_1167_));
 sg13g2_nand2_1 _2132_ (.Y(_1228_),
    .A(net320),
    .B(\perceptron1.we2[14] ));
 sg13g2_nand2_1 _2133_ (.Y(_1229_),
    .A(net287),
    .B(\perceptron1.we3[9] ));
 sg13g2_nor2_1 _2134_ (.A(_1167_),
    .B(_1229_),
    .Y(_1230_));
 sg13g2_a22oi_1 _2135_ (.Y(_1231_),
    .B1(net277),
    .B2(net287),
    .A2(net276),
    .A1(net289));
 sg13g2_nor3_1 _2136_ (.A(_1228_),
    .B(_1230_),
    .C(_1231_),
    .Y(_1232_));
 sg13g2_o21ai_1 _2137_ (.B1(_1228_),
    .Y(_1233_),
    .A1(_1230_),
    .A2(_1231_));
 sg13g2_nor2b_1 _2138_ (.A(_1232_),
    .B_N(_1233_),
    .Y(_1234_));
 sg13g2_xnor2_1 _2139_ (.Y(_1235_),
    .A(_1227_),
    .B(_1234_));
 sg13g2_nand2_1 _2140_ (.Y(_1236_),
    .A(net311),
    .B(\perceptron1.we2[11] ));
 sg13g2_nand2_1 _2141_ (.Y(_1237_),
    .A(net314),
    .B(\perceptron1.we2[13] ));
 sg13g2_nor2_1 _2142_ (.A(_1173_),
    .B(_1237_),
    .Y(_1238_));
 sg13g2_a22oi_1 _2143_ (.Y(_1239_),
    .B1(\perceptron1.we2[12] ),
    .B2(net314),
    .A2(\perceptron1.we2[13] ),
    .A1(net317));
 sg13g2_nor3_1 _2144_ (.A(_1236_),
    .B(_1238_),
    .C(_1239_),
    .Y(_1240_));
 sg13g2_o21ai_1 _2145_ (.B1(_1236_),
    .Y(_1241_),
    .A1(_1238_),
    .A2(_1239_));
 sg13g2_nand2b_1 _2146_ (.Y(_1242_),
    .B(_1241_),
    .A_N(_1240_));
 sg13g2_nor2_1 _2147_ (.A(_1235_),
    .B(_1242_),
    .Y(_1243_));
 sg13g2_xor2_1 _2148_ (.B(_1242_),
    .A(_1235_),
    .X(_1244_));
 sg13g2_xnor2_1 _2149_ (.Y(_1245_),
    .A(_1226_),
    .B(_1244_));
 sg13g2_nor2b_1 _2150_ (.A(_1245_),
    .B_N(_1225_),
    .Y(_1246_));
 sg13g2_xor2_1 _2151_ (.B(_1245_),
    .A(_1225_),
    .X(_1247_));
 sg13g2_xor2_1 _2152_ (.B(_1247_),
    .A(_1224_),
    .X(_1248_));
 sg13g2_xnor2_1 _2153_ (.Y(_1249_),
    .A(_1188_),
    .B(_1248_));
 sg13g2_nor2b_1 _2154_ (.A(_1249_),
    .B_N(_1187_),
    .Y(_1250_));
 sg13g2_xnor2_1 _2155_ (.Y(_1251_),
    .A(_1187_),
    .B(_1249_));
 sg13g2_nand2_1 _2156_ (.Y(_1252_),
    .A(_1186_),
    .B(_1251_));
 sg13g2_o21ai_1 _2157_ (.B1(_1175_),
    .Y(_1253_),
    .A1(_1117_),
    .A2(_1173_));
 sg13g2_inv_1 _2158_ (.Y(_1254_),
    .A(_1253_));
 sg13g2_xnor2_1 _2159_ (.Y(_1255_),
    .A(_1186_),
    .B(_1251_));
 sg13g2_o21ai_1 _2160_ (.B1(_1252_),
    .Y(_1256_),
    .A1(_1254_),
    .A2(_1255_));
 sg13g2_or2_1 _2161_ (.X(_1257_),
    .B(_1240_),
    .A(_1238_));
 sg13g2_a21oi_1 _2162_ (.A1(_1188_),
    .A2(_1248_),
    .Y(_1258_),
    .B1(_1250_));
 sg13g2_a21oi_1 _2163_ (.A1(_1226_),
    .A2(_1244_),
    .Y(_1259_),
    .B1(_1246_));
 sg13g2_o21ai_1 _2164_ (.B1(_1223_),
    .Y(_1260_),
    .A1(_1224_),
    .A2(_1247_));
 sg13g2_a21oi_1 _2165_ (.A1(_1227_),
    .A2(_1234_),
    .Y(_1261_),
    .B1(_1243_));
 sg13g2_o21ai_1 _2166_ (.B1(_1209_),
    .Y(_1262_),
    .A1(_1210_),
    .A2(_1221_));
 sg13g2_xnor2_1 _2167_ (.Y(_1263_),
    .A(_1261_),
    .B(_1262_));
 sg13g2_a21oi_1 _2168_ (.A1(_1212_),
    .A2(_1218_),
    .Y(_0064_),
    .B1(_1220_));
 sg13g2_nand2_1 _2169_ (.Y(_0065_),
    .A(_1199_),
    .B(_1207_));
 sg13g2_o21ai_1 _2170_ (.B1(_1217_),
    .Y(_0066_),
    .A1(_1152_),
    .A2(_1215_));
 sg13g2_xor2_1 _2171_ (.B(_0066_),
    .A(_0065_),
    .X(_0067_));
 sg13g2_nand2_1 _2172_ (.Y(_0068_),
    .A(net325),
    .B(\perceptron1.we1[13] ));
 sg13g2_xnor2_1 _2173_ (.Y(_0069_),
    .A(_1193_),
    .B(_0068_));
 sg13g2_nand2_1 _2174_ (.Y(_0070_),
    .A(net333),
    .B(\perceptron1.we1[15] ));
 sg13g2_nand2_1 _2175_ (.Y(_0071_),
    .A(net330),
    .B(\perceptron1.we1[14] ));
 sg13g2_nand2_1 _2176_ (.Y(_0072_),
    .A(net306),
    .B(\perceptron1.we3[15] ));
 sg13g2_xnor2_1 _2177_ (.Y(_0073_),
    .A(_0071_),
    .B(_0072_));
 sg13g2_xnor2_1 _2178_ (.Y(_0074_),
    .A(_0069_),
    .B(_0073_));
 sg13g2_xnor2_1 _2179_ (.Y(_0075_),
    .A(_0070_),
    .B(_0074_));
 sg13g2_nand2_1 _2180_ (.Y(_0076_),
    .A(net311),
    .B(\perceptron1.we2[12] ));
 sg13g2_nor2_1 _2181_ (.A(_1230_),
    .B(_1232_),
    .Y(_0077_));
 sg13g2_xor2_1 _2182_ (.B(_0077_),
    .A(_0076_),
    .X(_0078_));
 sg13g2_nand2_1 _2183_ (.Y(_0079_),
    .A(net320),
    .B(\perceptron1.we2[15] ));
 sg13g2_nand2_1 _2184_ (.Y(_0080_),
    .A(net289),
    .B(\perceptron1.we3[10] ));
 sg13g2_xor2_1 _2185_ (.B(_0080_),
    .A(_1229_),
    .X(_0081_));
 sg13g2_nand2_1 _2186_ (.Y(_0082_),
    .A(net317),
    .B(\perceptron1.we2[14] ));
 sg13g2_xor2_1 _2187_ (.B(_0082_),
    .A(_1237_),
    .X(_0083_));
 sg13g2_xnor2_1 _2188_ (.Y(_0084_),
    .A(_0081_),
    .B(_0083_));
 sg13g2_xnor2_1 _2189_ (.Y(_0085_),
    .A(_0079_),
    .B(_0084_));
 sg13g2_xnor2_1 _2190_ (.Y(_0086_),
    .A(_0078_),
    .B(_0085_));
 sg13g2_nand2_1 _2191_ (.Y(_0087_),
    .A(net300),
    .B(\perceptron1.we3[14] ));
 sg13g2_nor2_1 _2192_ (.A(_1194_),
    .B(_1196_),
    .Y(_0088_));
 sg13g2_xor2_1 _2193_ (.B(_0088_),
    .A(_0087_),
    .X(_0089_));
 sg13g2_or2_1 _2194_ (.X(_0090_),
    .B(_1204_),
    .A(_1202_));
 sg13g2_nand2_1 _2195_ (.Y(_0091_),
    .A(net292),
    .B(\perceptron1.we3[11] ));
 sg13g2_nand2_1 _2196_ (.Y(_0092_),
    .A(net297),
    .B(\perceptron1.we3[13] ));
 sg13g2_xor2_1 _2197_ (.B(_0092_),
    .A(_1214_),
    .X(_0093_));
 sg13g2_xnor2_1 _2198_ (.Y(_0094_),
    .A(_0091_),
    .B(_0093_));
 sg13g2_xnor2_1 _2199_ (.Y(_0095_),
    .A(_0090_),
    .B(_0094_));
 sg13g2_xnor2_1 _2200_ (.Y(_0096_),
    .A(_0064_),
    .B(_0086_));
 sg13g2_xnor2_1 _2201_ (.Y(_0097_),
    .A(_0075_),
    .B(_0089_));
 sg13g2_xnor2_1 _2202_ (.Y(_0098_),
    .A(_0095_),
    .B(_0097_));
 sg13g2_xnor2_1 _2203_ (.Y(_0099_),
    .A(_0096_),
    .B(_0098_));
 sg13g2_xnor2_1 _2204_ (.Y(_0100_),
    .A(_0067_),
    .B(_0099_));
 sg13g2_xnor2_1 _2205_ (.Y(_0101_),
    .A(_1263_),
    .B(_0100_));
 sg13g2_xnor2_1 _2206_ (.Y(_0102_),
    .A(_1260_),
    .B(_0101_));
 sg13g2_xnor2_1 _2207_ (.Y(_0103_),
    .A(_1259_),
    .B(_0102_));
 sg13g2_xnor2_1 _2208_ (.Y(_0104_),
    .A(_1258_),
    .B(_0103_));
 sg13g2_xnor2_1 _2209_ (.Y(_0105_),
    .A(_1257_),
    .B(_0104_));
 sg13g2_xnor2_1 _2210_ (.Y(_0106_),
    .A(_1256_),
    .B(_0105_));
 sg13g2_o21ai_1 _2211_ (.B1(_0700_),
    .Y(_0107_),
    .A1(_0701_),
    .A2(_0721_));
 sg13g2_xor2_1 _2212_ (.B(_1127_),
    .A(_1105_),
    .X(_0108_));
 sg13g2_a21o_1 _2213_ (.A2(_0718_),
    .A1(_0703_),
    .B1(_0720_),
    .X(_0109_));
 sg13g2_xnor2_1 _2214_ (.Y(_0110_),
    .A(_0107_),
    .B(_0108_));
 sg13g2_nor2b_1 _2215_ (.A(_0110_),
    .B_N(_0109_),
    .Y(_0111_));
 sg13g2_a21o_1 _2216_ (.A2(_0108_),
    .A1(_0107_),
    .B1(_0111_),
    .X(_0112_));
 sg13g2_xor2_1 _2217_ (.B(_1184_),
    .A(_1183_),
    .X(_0113_));
 sg13g2_nand2b_1 _2218_ (.Y(_0114_),
    .B(_0112_),
    .A_N(_0113_));
 sg13g2_o21ai_1 _2219_ (.B1(_1119_),
    .Y(_0115_),
    .A1(_1116_),
    .A2(_1120_));
 sg13g2_xor2_1 _2220_ (.B(_0113_),
    .A(_0112_),
    .X(_0116_));
 sg13g2_nand2b_1 _2221_ (.Y(_0117_),
    .B(_0115_),
    .A_N(_0116_));
 sg13g2_xnor2_1 _2222_ (.Y(_0118_),
    .A(_1254_),
    .B(_1255_));
 sg13g2_nand3_1 _2223_ (.B(_0117_),
    .C(_0118_),
    .A(_0114_),
    .Y(_0119_));
 sg13g2_a21o_1 _2224_ (.A2(_0117_),
    .A1(_0114_),
    .B1(_0118_),
    .X(_0120_));
 sg13g2_nand3_1 _2225_ (.B(_0119_),
    .C(_0120_),
    .A(_0106_),
    .Y(_0121_));
 sg13g2_a21o_1 _2226_ (.A2(_0722_),
    .A1(_0667_),
    .B1(_0724_),
    .X(_0122_));
 sg13g2_xnor2_1 _2227_ (.Y(_0123_),
    .A(_0109_),
    .B(_0110_));
 sg13g2_nand2_1 _2228_ (.Y(_0124_),
    .A(_0122_),
    .B(_0123_));
 sg13g2_o21ai_1 _2229_ (.B1(_0715_),
    .Y(_0125_),
    .A1(_0644_),
    .A2(_0713_));
 sg13g2_inv_1 _2230_ (.Y(_0126_),
    .A(_0125_));
 sg13g2_xnor2_1 _2231_ (.Y(_0127_),
    .A(_0122_),
    .B(_0123_));
 sg13g2_o21ai_1 _2232_ (.B1(_0124_),
    .Y(_0128_),
    .A1(_0126_),
    .A2(_0127_));
 sg13g2_xor2_1 _2233_ (.B(_0116_),
    .A(_0115_),
    .X(_0129_));
 sg13g2_nand2b_1 _2234_ (.Y(_0130_),
    .B(_0128_),
    .A_N(_0129_));
 sg13g2_xor2_1 _2235_ (.B(_0129_),
    .A(_0128_),
    .X(_0131_));
 sg13g2_xnor2_1 _2236_ (.Y(_0132_),
    .A(_0125_),
    .B(_0127_));
 sg13g2_o21ai_1 _2237_ (.B1(_0132_),
    .Y(_0133_),
    .A1(_0726_),
    .A2(_0728_));
 sg13g2_nor3_1 _2238_ (.A(_0726_),
    .B(_0728_),
    .C(_0132_),
    .Y(_0134_));
 sg13g2_nor3_1 _2239_ (.A(_0121_),
    .B(_0131_),
    .C(_0134_),
    .Y(_0135_));
 sg13g2_a21oi_1 _2240_ (.A1(_0133_),
    .A2(_0135_),
    .Y(_0136_),
    .B1(_1070_));
 sg13g2_and3_1 _2241_ (.X(_0137_),
    .A(_1017_),
    .B(_1066_),
    .C(_1067_));
 sg13g2_a21o_1 _2242_ (.A2(_1064_),
    .A1(_1042_),
    .B1(_1065_),
    .X(_0138_));
 sg13g2_or3_1 _2243_ (.A(_1054_),
    .B(_1055_),
    .C(_1061_),
    .X(_0139_));
 sg13g2_nand2_1 _2244_ (.Y(_0140_),
    .A(_1042_),
    .B(_1063_));
 sg13g2_xnor2_1 _2245_ (.Y(_0141_),
    .A(_1043_),
    .B(_0140_));
 sg13g2_a21oi_1 _2246_ (.A1(_1062_),
    .A2(_0139_),
    .Y(_0142_),
    .B1(_0141_));
 sg13g2_nand2_1 _2247_ (.Y(_0143_),
    .A(_1066_),
    .B(_0138_));
 sg13g2_nor4_2 _2248_ (.A(_1068_),
    .B(_0137_),
    .C(_0142_),
    .Y(_0144_),
    .D(_0143_));
 sg13g2_nor2_1 _2249_ (.A(_0131_),
    .B(_0133_),
    .Y(_0145_));
 sg13g2_o21ai_1 _2250_ (.B1(_0130_),
    .Y(_0146_),
    .A1(_0131_),
    .A2(_0133_));
 sg13g2_nor2_1 _2251_ (.A(_0106_),
    .B(_0120_),
    .Y(_0147_));
 sg13g2_o21ai_1 _2252_ (.B1(_0121_),
    .Y(_0148_),
    .A1(_0146_),
    .A2(_0147_));
 sg13g2_nand2b_1 _2253_ (.Y(_0149_),
    .B(_0148_),
    .A_N(_0144_));
 sg13g2_a21oi_1 _2254_ (.A1(_0131_),
    .A2(_0134_),
    .Y(_0150_),
    .B1(_0145_));
 sg13g2_o21ai_1 _2255_ (.B1(_0120_),
    .Y(_0151_),
    .A1(_0106_),
    .A2(_0119_));
 sg13g2_nor2_1 _2256_ (.A(_0146_),
    .B(_0151_),
    .Y(_0152_));
 sg13g2_nor2_1 _2257_ (.A(_0150_),
    .B(_0152_),
    .Y(_0153_));
 sg13g2_nor2_1 _2258_ (.A(_0926_),
    .B(_0153_),
    .Y(_0154_));
 sg13g2_or3_1 _2259_ (.A(_0914_),
    .B(_0917_),
    .C(_0918_),
    .X(_0155_));
 sg13g2_nand2b_1 _2260_ (.Y(_0156_),
    .B(_0920_),
    .A_N(_0155_));
 sg13g2_nand2b_1 _2261_ (.Y(_0157_),
    .B(_0156_),
    .A_N(_0922_));
 sg13g2_o21ai_1 _2262_ (.B1(_0925_),
    .Y(_0158_),
    .A1(_0731_),
    .A2(_0799_));
 sg13g2_nand2_1 _2263_ (.Y(_0159_),
    .A(_0923_),
    .B(_0158_));
 sg13g2_nand2_1 _2264_ (.Y(_0160_),
    .A(_0924_),
    .B(_0159_));
 sg13g2_nand3b_1 _2265_ (.B(_0157_),
    .C(_0160_),
    .Y(_0161_),
    .A_N(_0154_));
 sg13g2_nand4_1 _2266_ (.B(_0919_),
    .C(_0921_),
    .A(_0800_),
    .Y(_0162_),
    .D(_0155_));
 sg13g2_mux2_1 _2267_ (.A0(_0161_),
    .A1(_0162_),
    .S(_1069_),
    .X(_0163_));
 sg13g2_or3_1 _2268_ (.A(_0136_),
    .B(_0149_),
    .C(_0163_),
    .X(_0000_));
 sg13g2_nor2b_1 _2269_ (.A(net2),
    .B_N(\perceptron1.out ),
    .Y(_0164_));
 sg13g2_nand2b_2 _2270_ (.Y(_0165_),
    .B(\perceptron1.out ),
    .A_N(net2));
 sg13g2_nor2b_1 _2271_ (.A(\perceptron1.out ),
    .B_N(net2),
    .Y(_0166_));
 sg13g2_nor2_1 _2272_ (.A(net269),
    .B(_0166_),
    .Y(_0167_));
 sg13g2_xor2_1 _2273_ (.B(\perceptron1.out ),
    .A(net2),
    .X(_0168_));
 sg13g2_nand3_1 _2274_ (.B(net301),
    .C(net270),
    .A(net307),
    .Y(_0169_));
 sg13g2_and4_1 _2275_ (.A(net307),
    .B(net301),
    .C(net298),
    .D(net269),
    .X(_0170_));
 sg13g2_nand4_1 _2276_ (.B(net301),
    .C(net298),
    .A(net307),
    .Y(_0171_),
    .D(net269));
 sg13g2_nor3_2 _2277_ (.A(net307),
    .B(net301),
    .C(net298),
    .Y(_0172_));
 sg13g2_o21ai_1 _2278_ (.B1(net270),
    .Y(_0173_),
    .A1(net307),
    .A2(net301));
 sg13g2_nor2_1 _2279_ (.A(_0165_),
    .B(_0172_),
    .Y(_0174_));
 sg13g2_nand2b_1 _2280_ (.Y(_0175_),
    .B(net269),
    .A_N(_0172_));
 sg13g2_nor2_1 _2281_ (.A(net295),
    .B(net293),
    .Y(_0176_));
 sg13g2_xor2_1 _2282_ (.B(net293),
    .A(net295),
    .X(_0177_));
 sg13g2_a22oi_1 _2283_ (.Y(_0178_),
    .B1(_0177_),
    .B2(net269),
    .A2(_0166_),
    .A1(net293));
 sg13g2_nand3b_1 _2284_ (.B(_0171_),
    .C(_0174_),
    .Y(_0179_),
    .A_N(_0178_));
 sg13g2_o21ai_1 _2285_ (.B1(_0178_),
    .Y(_0180_),
    .A1(_0170_),
    .A2(_0175_));
 sg13g2_and2_1 _2286_ (.A(net295),
    .B(net265),
    .X(_0181_));
 sg13g2_nand3b_1 _2287_ (.B(net269),
    .C(net295),
    .Y(_0182_),
    .A_N(_0172_));
 sg13g2_mux2_1 _2288_ (.A0(_0181_),
    .A1(_0182_),
    .S(_0171_),
    .X(_0183_));
 sg13g2_a21oi_1 _2289_ (.A1(_0179_),
    .A2(_0180_),
    .Y(_0184_),
    .B1(_0183_));
 sg13g2_nand3_1 _2290_ (.B(_0180_),
    .C(_0183_),
    .A(_0179_),
    .Y(_0185_));
 sg13g2_nor2b_1 _2291_ (.A(_0184_),
    .B_N(_0185_),
    .Y(_0186_));
 sg13g2_nand2b_1 _2292_ (.Y(_0187_),
    .B(_0185_),
    .A_N(_0184_));
 sg13g2_nand2_1 _2293_ (.Y(_0188_),
    .A(net288),
    .B(net267));
 sg13g2_nor3_1 _2294_ (.A(net295),
    .B(net293),
    .C(net291),
    .Y(_0189_));
 sg13g2_a21oi_2 _2295_ (.B1(_0165_),
    .Y(_0190_),
    .A2(_0189_),
    .A1(_0172_));
 sg13g2_xnor2_1 _2296_ (.Y(_0191_),
    .A(_0188_),
    .B(_0190_));
 sg13g2_inv_1 _2297_ (.Y(_0192_),
    .A(_0191_));
 sg13g2_a21oi_1 _2298_ (.A1(_0172_),
    .A2(_0176_),
    .Y(_0193_),
    .B1(net2));
 sg13g2_or2_1 _2299_ (.X(_0194_),
    .B(_0193_),
    .A(net291));
 sg13g2_a21oi_1 _2300_ (.A1(net291),
    .A2(_0193_),
    .Y(_0195_),
    .B1(net264));
 sg13g2_and2_1 _2301_ (.A(_0194_),
    .B(_0195_),
    .X(_0196_));
 sg13g2_nand2_1 _2302_ (.Y(_0197_),
    .A(_0194_),
    .B(_0195_));
 sg13g2_a21oi_2 _2303_ (.B1(_0190_),
    .Y(_0198_),
    .A2(net269),
    .A1(net288));
 sg13g2_a21o_2 _2304_ (.A2(net269),
    .A1(net288),
    .B1(_0190_),
    .X(_0199_));
 sg13g2_o21ai_1 _2305_ (.B1(_0199_),
    .Y(_0200_),
    .A1(_0191_),
    .A2(_0196_));
 sg13g2_a21oi_2 _2306_ (.B1(_0192_),
    .Y(_0201_),
    .A2(_0199_),
    .A1(_0197_));
 sg13g2_nand3_1 _2307_ (.B(_0195_),
    .C(_0198_),
    .A(_0194_),
    .Y(_0202_));
 sg13g2_nand3b_1 _2308_ (.B(_0185_),
    .C(_0202_),
    .Y(_0203_),
    .A_N(_0184_));
 sg13g2_xnor2_1 _2309_ (.Y(_0204_),
    .A(_0197_),
    .B(_0200_));
 sg13g2_nor3_2 _2310_ (.A(_0191_),
    .B(_0196_),
    .C(_0198_),
    .Y(_0205_));
 sg13g2_a21oi_1 _2311_ (.A1(_0201_),
    .A2(_0203_),
    .Y(_0206_),
    .B1(_0205_));
 sg13g2_a21o_1 _2312_ (.A2(_0203_),
    .A1(_0201_),
    .B1(_0205_),
    .X(_0207_));
 sg13g2_xnor2_1 _2313_ (.Y(_0208_),
    .A(_0186_),
    .B(_0206_));
 sg13g2_inv_1 _2314_ (.Y(_0209_),
    .A(_0208_));
 sg13g2_xnor2_1 _2315_ (.Y(_0210_),
    .A(_0174_),
    .B(_0181_));
 sg13g2_and2_1 _2316_ (.A(_0208_),
    .B(_0210_),
    .X(_0211_));
 sg13g2_nand2_1 _2317_ (.Y(_0212_),
    .A(_0208_),
    .B(_0210_));
 sg13g2_a21oi_1 _2318_ (.A1(_0187_),
    .A2(_0205_),
    .Y(_0213_),
    .B1(_0201_));
 sg13g2_a21oi_2 _2319_ (.B1(_0213_),
    .Y(_0214_),
    .A2(_0203_),
    .A1(_0201_));
 sg13g2_a21o_1 _2320_ (.A2(_0207_),
    .A1(_0186_),
    .B1(_0204_),
    .X(_0215_));
 sg13g2_nand2_1 _2321_ (.Y(_0216_),
    .A(_0186_),
    .B(_0205_));
 sg13g2_nand2_1 _2322_ (.Y(_0217_),
    .A(_0215_),
    .B(_0216_));
 sg13g2_a22oi_1 _2323_ (.Y(_0218_),
    .B1(_0215_),
    .B2(_0216_),
    .A2(_0210_),
    .A1(_0208_));
 sg13g2_nor2_1 _2324_ (.A(_0214_),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_o21ai_1 _2325_ (.B1(_0210_),
    .Y(_0220_),
    .A1(_0214_),
    .A2(_0218_));
 sg13g2_a22oi_1 _2326_ (.Y(_0221_),
    .B1(_0220_),
    .B2(_0209_),
    .A2(_0214_),
    .A1(_0211_));
 sg13g2_or3_1 _2327_ (.A(_0210_),
    .B(_0214_),
    .C(_0217_),
    .X(_0222_));
 sg13g2_nand2_1 _2328_ (.Y(_0223_),
    .A(_0220_),
    .B(_0222_));
 sg13g2_a21o_1 _2329_ (.A2(net270),
    .A1(net307),
    .B1(net301),
    .X(_0224_));
 sg13g2_nand3_1 _2330_ (.B(_0169_),
    .C(_0224_),
    .A(net265),
    .Y(_0225_));
 sg13g2_o21ai_1 _2331_ (.B1(_0173_),
    .Y(_0226_),
    .A1(_0342_),
    .A2(net263));
 sg13g2_o21ai_1 _2332_ (.B1(_0226_),
    .Y(_0227_),
    .A1(_0342_),
    .A2(_0173_));
 sg13g2_and2_1 _2333_ (.A(_0225_),
    .B(_0227_),
    .X(_0228_));
 sg13g2_a21o_1 _2334_ (.A2(_0222_),
    .A1(_0220_),
    .B1(_0228_),
    .X(_0229_));
 sg13g2_nand3_1 _2335_ (.B(_0222_),
    .C(_0227_),
    .A(_0220_),
    .Y(_0230_));
 sg13g2_nor2b_1 _2336_ (.A(_0221_),
    .B_N(_0230_),
    .Y(_0231_));
 sg13g2_mux2_1 _2337_ (.A0(_0230_),
    .A1(_0229_),
    .S(_0221_),
    .X(_0232_));
 sg13g2_a21oi_1 _2338_ (.A1(_0212_),
    .A2(_0214_),
    .Y(_0233_),
    .B1(_0217_));
 sg13g2_nor2_1 _2339_ (.A(_0218_),
    .B(_0233_),
    .Y(_0234_));
 sg13g2_nor2_1 _2340_ (.A(_0225_),
    .B(_0227_),
    .Y(_0235_));
 sg13g2_a21oi_1 _2341_ (.A1(_0223_),
    .A2(_0235_),
    .Y(_0236_),
    .B1(_0234_));
 sg13g2_a21o_1 _2342_ (.A2(_0236_),
    .A1(_0232_),
    .B1(net61),
    .X(_0237_));
 sg13g2_nand3_1 _2343_ (.B(_0232_),
    .C(_0236_),
    .A(net61),
    .Y(_0238_));
 sg13g2_a21oi_1 _2344_ (.A1(_0237_),
    .A2(_0238_),
    .Y(_0239_),
    .B1(net263));
 sg13g2_a21oi_1 _2345_ (.A1(_0353_),
    .A2(net263),
    .Y(_0016_),
    .B1(_0239_));
 sg13g2_nor2_1 _2346_ (.A(net32),
    .B(net266),
    .Y(_0240_));
 sg13g2_nor3_1 _2347_ (.A(net285),
    .B(_0231_),
    .C(_0234_),
    .Y(_0241_));
 sg13g2_o21ai_1 _2348_ (.B1(net285),
    .Y(_0242_),
    .A1(_0231_),
    .A2(_0234_));
 sg13g2_nor2b_1 _2349_ (.A(_0241_),
    .B_N(_0242_),
    .Y(_0243_));
 sg13g2_xnor2_1 _2350_ (.Y(_0244_),
    .A(_0237_),
    .B(_0243_));
 sg13g2_a21oi_1 _2351_ (.A1(net266),
    .A2(_0244_),
    .Y(_0017_),
    .B1(_0240_));
 sg13g2_o21ai_1 _2352_ (.B1(_0242_),
    .Y(_0245_),
    .A1(_0237_),
    .A2(_0241_));
 sg13g2_nor2b_1 _2353_ (.A(_0219_),
    .B_N(net284),
    .Y(_0246_));
 sg13g2_xnor2_1 _2354_ (.Y(_0247_),
    .A(net284),
    .B(_0219_));
 sg13g2_xnor2_1 _2355_ (.Y(_0248_),
    .A(_0245_),
    .B(_0247_));
 sg13g2_mux2_1 _2356_ (.A0(net29),
    .A1(_0248_),
    .S(net265),
    .X(_0018_));
 sg13g2_nor2_1 _2357_ (.A(net34),
    .B(net267),
    .Y(_0249_));
 sg13g2_a21oi_1 _2358_ (.A1(_0245_),
    .A2(_0247_),
    .Y(_0250_),
    .B1(_0246_));
 sg13g2_nor2_1 _2359_ (.A(net282),
    .B(_0207_),
    .Y(_0251_));
 sg13g2_xnor2_1 _2360_ (.Y(_0252_),
    .A(net282),
    .B(_0206_));
 sg13g2_xnor2_1 _2361_ (.Y(_0253_),
    .A(_0250_),
    .B(_0252_));
 sg13g2_a21oi_1 _2362_ (.A1(net267),
    .A2(_0253_),
    .Y(_0019_),
    .B1(_0249_));
 sg13g2_nor2_1 _2363_ (.A(_0371_),
    .B(_0200_),
    .Y(_0254_));
 sg13g2_xnor2_1 _2364_ (.Y(_0255_),
    .A(_0371_),
    .B(_0200_));
 sg13g2_a221oi_1 _2365_ (.B2(_0247_),
    .C1(_0246_),
    .B1(_0245_),
    .A1(net282),
    .Y(_0256_),
    .A2(_0207_));
 sg13g2_o21ai_1 _2366_ (.B1(_0255_),
    .Y(_0257_),
    .A1(_0251_),
    .A2(_0256_));
 sg13g2_nor3_1 _2367_ (.A(_0251_),
    .B(_0255_),
    .C(_0256_),
    .Y(_0258_));
 sg13g2_nor2_1 _2368_ (.A(net263),
    .B(_0258_),
    .Y(_0259_));
 sg13g2_a22oi_1 _2369_ (.Y(_0020_),
    .B1(_0257_),
    .B2(_0259_),
    .A2(net263),
    .A1(_0335_));
 sg13g2_nor2_1 _2370_ (.A(_0254_),
    .B(_0258_),
    .Y(_0260_));
 sg13g2_o21ai_1 _2371_ (.B1(net280),
    .Y(_0261_),
    .A1(_0254_),
    .A2(_0258_));
 sg13g2_xnor2_1 _2372_ (.Y(_0021_),
    .A(net280),
    .B(_0260_));
 sg13g2_nor2_1 _2373_ (.A(_0362_),
    .B(_0261_),
    .Y(_0262_));
 sg13g2_xnor2_1 _2374_ (.Y(_0022_),
    .A(net279),
    .B(_0261_));
 sg13g2_nand2_1 _2375_ (.Y(_0263_),
    .A(net278),
    .B(_0199_));
 sg13g2_nand2b_1 _2376_ (.Y(_0264_),
    .B(_0198_),
    .A_N(net278));
 sg13g2_and2_1 _2377_ (.A(_0263_),
    .B(_0264_),
    .X(_0265_));
 sg13g2_xor2_1 _2378_ (.B(_0265_),
    .A(_0262_),
    .X(_0023_));
 sg13g2_nand2_1 _2379_ (.Y(_0266_),
    .A(net277),
    .B(_0199_));
 sg13g2_xnor2_1 _2380_ (.Y(_0267_),
    .A(net277),
    .B(_0198_));
 sg13g2_o21ai_1 _2381_ (.B1(_0263_),
    .Y(_0268_),
    .A1(_0362_),
    .A2(_0261_));
 sg13g2_a21oi_1 _2382_ (.A1(_0264_),
    .A2(_0268_),
    .Y(_0269_),
    .B1(_0267_));
 sg13g2_nand3_1 _2383_ (.B(_0267_),
    .C(_0268_),
    .A(_0264_),
    .Y(_0270_));
 sg13g2_nor2b_1 _2384_ (.A(_0269_),
    .B_N(_0270_),
    .Y(_0024_));
 sg13g2_nand2_1 _2385_ (.Y(_0271_),
    .A(_0266_),
    .B(_0270_));
 sg13g2_xor2_1 _2386_ (.B(_0271_),
    .A(net276),
    .X(_0025_));
 sg13g2_nand2_1 _2387_ (.Y(_0272_),
    .A(net275),
    .B(net276));
 sg13g2_a21oi_1 _2388_ (.A1(_0266_),
    .A2(_0270_),
    .Y(_0273_),
    .B1(_0272_));
 sg13g2_a21oi_1 _2389_ (.A1(net276),
    .A2(_0271_),
    .Y(_0274_),
    .B1(net275));
 sg13g2_nor2_1 _2390_ (.A(_0273_),
    .B(net70),
    .Y(_0026_));
 sg13g2_nand2_1 _2391_ (.Y(_0275_),
    .A(\perceptron1.we3[11] ),
    .B(_0199_));
 sg13g2_xnor2_1 _2392_ (.Y(_0276_),
    .A(net86),
    .B(_0198_));
 sg13g2_xor2_1 _2393_ (.B(_0276_),
    .A(_0273_),
    .X(_0027_));
 sg13g2_nor2b_1 _2394_ (.A(_0272_),
    .B_N(_0276_),
    .Y(_0277_));
 sg13g2_and4_1 _2395_ (.A(_0264_),
    .B(_0267_),
    .C(_0268_),
    .D(_0277_),
    .X(_0278_));
 sg13g2_o21ai_1 _2396_ (.B1(_0275_),
    .Y(_0279_),
    .A1(_0266_),
    .A2(_0272_));
 sg13g2_nor2_1 _2397_ (.A(_0278_),
    .B(_0279_),
    .Y(_0280_));
 sg13g2_nand2_1 _2398_ (.Y(_0281_),
    .A(\perceptron1.we3[12] ),
    .B(_0199_));
 sg13g2_xnor2_1 _2399_ (.Y(_0282_),
    .A(net82),
    .B(_0198_));
 sg13g2_o21ai_1 _2400_ (.B1(_0282_),
    .Y(_0283_),
    .A1(_0278_),
    .A2(_0279_));
 sg13g2_xnor2_1 _2401_ (.Y(_0028_),
    .A(_0280_),
    .B(_0282_));
 sg13g2_nand2_1 _2402_ (.Y(_0284_),
    .A(net50),
    .B(net263));
 sg13g2_a21oi_2 _2403_ (.B1(net43),
    .Y(_0285_),
    .A2(_0283_),
    .A1(_0281_));
 sg13g2_nand3_1 _2404_ (.B(_0281_),
    .C(_0283_),
    .A(net43),
    .Y(_0286_));
 sg13g2_nand2_1 _2405_ (.Y(_0287_),
    .A(net267),
    .B(_0286_));
 sg13g2_o21ai_1 _2406_ (.B1(_0284_),
    .Y(_0029_),
    .A1(_0285_),
    .A2(_0287_));
 sg13g2_nand2_1 _2407_ (.Y(_0288_),
    .A(\perceptron1.we3[14] ),
    .B(_0285_));
 sg13g2_xor2_1 _2408_ (.B(_0285_),
    .A(\perceptron1.we3[14] ),
    .X(_0030_));
 sg13g2_xnor2_1 _2409_ (.Y(_0031_),
    .A(net38),
    .B(_0288_));
 sg13g2_nand3_1 _2410_ (.B(net331),
    .C(net337),
    .A(net327),
    .Y(_0289_));
 sg13g2_or3_1 _2411_ (.A(net327),
    .B(net331),
    .C(net336),
    .X(_0290_));
 sg13g2_nand3_1 _2412_ (.B(_0289_),
    .C(_0290_),
    .A(net270),
    .Y(_0291_));
 sg13g2_nand2_1 _2413_ (.Y(_0292_),
    .A(net323),
    .B(net265));
 sg13g2_nand3_1 _2414_ (.B(net337),
    .C(net270),
    .A(net328),
    .Y(_0293_));
 sg13g2_nand2_1 _2415_ (.Y(_0294_),
    .A(net266),
    .B(_0293_));
 sg13g2_a221oi_1 _2416_ (.B2(net327),
    .C1(net331),
    .B1(net266),
    .A1(net336),
    .Y(_0295_),
    .A2(net270));
 sg13g2_a21o_1 _2417_ (.A2(_0294_),
    .A1(net331),
    .B1(_0295_),
    .X(_0296_));
 sg13g2_xnor2_1 _2418_ (.Y(_0297_),
    .A(_0291_),
    .B(_0292_));
 sg13g2_o21ai_1 _2419_ (.B1(_0004_),
    .Y(_0298_),
    .A1(_0296_),
    .A2(_0297_));
 sg13g2_nor3_2 _2420_ (.A(net75),
    .B(_0296_),
    .C(_0297_),
    .Y(_0299_));
 sg13g2_nand2_1 _2421_ (.Y(_0300_),
    .A(net266),
    .B(_0298_));
 sg13g2_nand2_1 _2422_ (.Y(_0301_),
    .A(net55),
    .B(net263));
 sg13g2_o21ai_1 _2423_ (.B1(_0301_),
    .Y(_0032_),
    .A1(_0299_),
    .A2(_0300_));
 sg13g2_nor2_1 _2424_ (.A(net30),
    .B(net265),
    .Y(_0302_));
 sg13g2_xor2_1 _2425_ (.B(_0299_),
    .A(\perceptron1.we1[1] ),
    .X(_0303_));
 sg13g2_a21oi_1 _2426_ (.A1(net265),
    .A2(_0303_),
    .Y(_0033_),
    .B1(_0302_));
 sg13g2_nand3_1 _2427_ (.B(\perceptron1.we1[2] ),
    .C(_0299_),
    .A(\perceptron1.we1[1] ),
    .Y(_0304_));
 sg13g2_a21o_1 _2428_ (.A2(_0299_),
    .A1(\perceptron1.we1[1] ),
    .B1(\perceptron1.we1[2] ),
    .X(_0305_));
 sg13g2_and2_1 _2429_ (.A(_0304_),
    .B(net76),
    .X(_0034_));
 sg13g2_nor2_1 _2430_ (.A(net28),
    .B(net265),
    .Y(_0306_));
 sg13g2_nor2_1 _2431_ (.A(net324),
    .B(_0290_),
    .Y(_0307_));
 sg13g2_nor2_1 _2432_ (.A(_0165_),
    .B(_0307_),
    .Y(_0308_));
 sg13g2_nand2_1 _2433_ (.Y(_0309_),
    .A(net274),
    .B(net262));
 sg13g2_xnor2_1 _2434_ (.Y(_0310_),
    .A(net274),
    .B(net262));
 sg13g2_or2_1 _2435_ (.X(_0311_),
    .B(_0310_),
    .A(_0304_));
 sg13g2_xor2_1 _2436_ (.B(_0310_),
    .A(_0304_),
    .X(_0312_));
 sg13g2_a21oi_1 _2437_ (.A1(net265),
    .A2(_0312_),
    .Y(_0035_),
    .B1(_0306_));
 sg13g2_xnor2_1 _2438_ (.Y(_0313_),
    .A(\perceptron1.we1[4] ),
    .B(net262));
 sg13g2_a21oi_1 _2439_ (.A1(_0309_),
    .A2(_0311_),
    .Y(_0314_),
    .B1(_0313_));
 sg13g2_nand3_1 _2440_ (.B(_0311_),
    .C(_0313_),
    .A(_0309_),
    .Y(_0315_));
 sg13g2_nor2b_1 _2441_ (.A(_0314_),
    .B_N(_0315_),
    .Y(_0036_));
 sg13g2_a21o_1 _2442_ (.A2(net262),
    .A1(\perceptron1.we1[4] ),
    .B1(_0314_),
    .X(_0316_));
 sg13g2_xor2_1 _2443_ (.B(_0316_),
    .A(net273),
    .X(_0037_));
 sg13g2_nand3_1 _2444_ (.B(net80),
    .C(_0316_),
    .A(net273),
    .Y(_0317_));
 sg13g2_a21o_1 _2445_ (.A2(_0316_),
    .A1(net273),
    .B1(net80),
    .X(_0318_));
 sg13g2_and2_1 _2446_ (.A(_0317_),
    .B(_0318_),
    .X(_0038_));
 sg13g2_nand2_1 _2447_ (.Y(_0319_),
    .A(\perceptron1.we1[7] ),
    .B(net262));
 sg13g2_xnor2_1 _2448_ (.Y(_0320_),
    .A(\perceptron1.we1[7] ),
    .B(net261));
 sg13g2_or2_1 _2449_ (.X(_0321_),
    .B(_0320_),
    .A(_0317_));
 sg13g2_xor2_1 _2450_ (.B(_0320_),
    .A(_0317_),
    .X(_0039_));
 sg13g2_xnor2_1 _2451_ (.Y(_0322_),
    .A(\perceptron1.we1[8] ),
    .B(net261));
 sg13g2_a21oi_1 _2452_ (.A1(_0319_),
    .A2(_0321_),
    .Y(_0323_),
    .B1(_0322_));
 sg13g2_nand3_1 _2453_ (.B(_0321_),
    .C(_0322_),
    .A(_0319_),
    .Y(_0324_));
 sg13g2_nor2b_1 _2454_ (.A(_0323_),
    .B_N(_0324_),
    .Y(_0040_));
 sg13g2_a21oi_1 _2455_ (.A1(\perceptron1.we1[8] ),
    .A2(net261),
    .Y(_0325_),
    .B1(_0323_));
 sg13g2_nor2b_1 _2456_ (.A(_0325_),
    .B_N(\perceptron1.we1[9] ),
    .Y(_0326_));
 sg13g2_xnor2_1 _2457_ (.Y(_0041_),
    .A(net67),
    .B(_0325_));
 sg13g2_nand2_1 _2458_ (.Y(_0327_),
    .A(net63),
    .B(_0326_));
 sg13g2_xor2_1 _2459_ (.B(_0326_),
    .A(net63),
    .X(_0042_));
 sg13g2_nand2_1 _2460_ (.Y(_0328_),
    .A(net272),
    .B(net261));
 sg13g2_nor2_1 _2461_ (.A(net272),
    .B(net261),
    .Y(_0329_));
 sg13g2_xor2_1 _2462_ (.B(net261),
    .A(net272),
    .X(_0330_));
 sg13g2_xnor2_1 _2463_ (.Y(_0043_),
    .A(_0327_),
    .B(_0330_));
 sg13g2_nand2_1 _2464_ (.Y(_0331_),
    .A(\perceptron1.we1[12] ),
    .B(net261));
 sg13g2_xnor2_1 _2465_ (.Y(_0332_),
    .A(net88),
    .B(net261));
 sg13g2_a21oi_1 _2466_ (.A1(_0327_),
    .A2(_0328_),
    .Y(_0333_),
    .B1(_0329_));
 sg13g2_nand2b_1 _2467_ (.Y(_0334_),
    .B(_0333_),
    .A_N(_0332_));
 sg13g2_xnor2_1 _2468_ (.Y(_0044_),
    .A(_0332_),
    .B(_0333_));
 sg13g2_nand2_1 _2469_ (.Y(_0336_),
    .A(net49),
    .B(net263));
 sg13g2_a21oi_2 _2470_ (.B1(net45),
    .Y(_0337_),
    .A2(_0334_),
    .A1(_0331_));
 sg13g2_nand3_1 _2471_ (.B(_0331_),
    .C(_0334_),
    .A(net45),
    .Y(_0338_));
 sg13g2_nand2_1 _2472_ (.Y(_0339_),
    .A(net267),
    .B(_0338_));
 sg13g2_o21ai_1 _2473_ (.B1(_0336_),
    .Y(_0045_),
    .A1(_0337_),
    .A2(_0339_));
 sg13g2_nand2_1 _2474_ (.Y(_0340_),
    .A(\perceptron1.we1[14] ),
    .B(_0337_));
 sg13g2_xor2_1 _2475_ (.B(_0337_),
    .A(\perceptron1.we1[14] ),
    .X(_0046_));
 sg13g2_xnor2_1 _2476_ (.Y(_0047_),
    .A(net36),
    .B(_0340_));
 sg13g2_nand2_1 _2477_ (.Y(_0341_),
    .A(net319),
    .B(net271));
 sg13g2_xor2_1 _2478_ (.B(_0341_),
    .A(net315),
    .X(_0343_));
 sg13g2_nor2_1 _2479_ (.A(net264),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_o21ai_1 _2480_ (.B1(net271),
    .Y(_0345_),
    .A1(net319),
    .A2(net315));
 sg13g2_a21oi_1 _2481_ (.A1(net312),
    .A2(net268),
    .Y(_0346_),
    .B1(_0345_));
 sg13g2_and3_1 _2482_ (.X(_0347_),
    .A(net312),
    .B(net268),
    .C(_0345_));
 sg13g2_nor3_1 _2483_ (.A(_0344_),
    .B(_0346_),
    .C(_0347_),
    .Y(_0348_));
 sg13g2_nand2_1 _2484_ (.Y(_0349_),
    .A(net310),
    .B(net268));
 sg13g2_a21oi_1 _2485_ (.A1(net312),
    .A2(net271),
    .Y(_0350_),
    .B1(_0346_));
 sg13g2_xnor2_1 _2486_ (.Y(_0351_),
    .A(_0349_),
    .B(_0350_));
 sg13g2_nor3_2 _2487_ (.A(_0002_),
    .B(_0348_),
    .C(_0351_),
    .Y(_0352_));
 sg13g2_o21ai_1 _2488_ (.B1(_0002_),
    .Y(_0354_),
    .A1(_0348_),
    .A2(_0351_));
 sg13g2_nand2_1 _2489_ (.Y(_0355_),
    .A(net268),
    .B(_0354_));
 sg13g2_nand2_1 _2490_ (.Y(_0356_),
    .A(net51),
    .B(net264));
 sg13g2_o21ai_1 _2491_ (.B1(_0356_),
    .Y(_0048_),
    .A1(_0352_),
    .A2(_0355_));
 sg13g2_and2_1 _2492_ (.A(_0387_),
    .B(_0352_),
    .X(_0357_));
 sg13g2_o21ai_1 _2493_ (.B1(_0168_),
    .Y(_0358_),
    .A1(_0387_),
    .A2(_0352_));
 sg13g2_nand2_1 _2494_ (.Y(_0359_),
    .A(net53),
    .B(net264));
 sg13g2_o21ai_1 _2495_ (.B1(_0359_),
    .Y(_0049_),
    .A1(_0357_),
    .A2(_0358_));
 sg13g2_and2_1 _2496_ (.A(net84),
    .B(_0357_),
    .X(_0360_));
 sg13g2_xnor2_1 _2497_ (.Y(_0361_),
    .A(\perceptron1.we2[2] ),
    .B(_0357_));
 sg13g2_mux2_1 _2498_ (.A0(net26),
    .A1(_0361_),
    .S(net268),
    .X(_0050_));
 sg13g2_nand4_1 _2499_ (.B(net315),
    .C(net312),
    .A(net319),
    .Y(_0363_),
    .D(net271));
 sg13g2_nand2_1 _2500_ (.Y(_0364_),
    .A(_0349_),
    .B(_0363_));
 sg13g2_o21ai_1 _2501_ (.B1(net271),
    .Y(_0365_),
    .A1(net315),
    .A2(net310));
 sg13g2_o21ai_1 _2502_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_0350_),
    .A2(_0364_));
 sg13g2_and2_1 _2503_ (.A(\perceptron1.we2[3] ),
    .B(net260),
    .X(_0367_));
 sg13g2_xor2_1 _2504_ (.B(net260),
    .A(\perceptron1.we2[3] ),
    .X(_0368_));
 sg13g2_xor2_1 _2505_ (.B(_0368_),
    .A(_0360_),
    .X(_0051_));
 sg13g2_nor2_1 _2506_ (.A(net35),
    .B(net268),
    .Y(_0369_));
 sg13g2_a21oi_1 _2507_ (.A1(_0360_),
    .A2(_0368_),
    .Y(_0370_),
    .B1(_0367_));
 sg13g2_xor2_1 _2508_ (.B(net260),
    .A(\perceptron1.we2[4] ),
    .X(_0372_));
 sg13g2_nor2b_1 _2509_ (.A(_0370_),
    .B_N(_0372_),
    .Y(_0373_));
 sg13g2_xnor2_1 _2510_ (.Y(_0374_),
    .A(_0370_),
    .B(_0372_));
 sg13g2_a21oi_1 _2511_ (.A1(net268),
    .A2(_0374_),
    .Y(_0052_),
    .B1(_0369_));
 sg13g2_a21oi_1 _2512_ (.A1(\perceptron1.we2[4] ),
    .A2(net260),
    .Y(_0375_),
    .B1(_0373_));
 sg13g2_nand2b_1 _2513_ (.Y(_0376_),
    .B(\perceptron1.we2[5] ),
    .A_N(_0375_));
 sg13g2_xnor2_1 _2514_ (.Y(_0053_),
    .A(net65),
    .B(_0375_));
 sg13g2_nor2_1 _2515_ (.A(_0379_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_xnor2_1 _2516_ (.Y(_0054_),
    .A(net59),
    .B(_0376_));
 sg13g2_and2_1 _2517_ (.A(net83),
    .B(net259),
    .X(_0378_));
 sg13g2_xor2_1 _2518_ (.B(net259),
    .A(net83),
    .X(_0380_));
 sg13g2_xor2_1 _2519_ (.B(_0380_),
    .A(_0377_),
    .X(_0055_));
 sg13g2_a21oi_1 _2520_ (.A1(_0377_),
    .A2(_0380_),
    .Y(_0381_),
    .B1(_0378_));
 sg13g2_nor2_1 _2521_ (.A(net77),
    .B(net259),
    .Y(_0382_));
 sg13g2_nand2_1 _2522_ (.Y(_0383_),
    .A(\perceptron1.we2[8] ),
    .B(net259));
 sg13g2_nor2b_1 _2523_ (.A(_0382_),
    .B_N(net78),
    .Y(_0384_));
 sg13g2_xnor2_1 _2524_ (.Y(_0056_),
    .A(_0381_),
    .B(_0384_));
 sg13g2_o21ai_1 _2525_ (.B1(_0383_),
    .Y(_0385_),
    .A1(_0381_),
    .A2(_0382_));
 sg13g2_xor2_1 _2526_ (.B(_0385_),
    .A(net62),
    .X(_0057_));
 sg13g2_nand3_1 _2527_ (.B(net62),
    .C(_0385_),
    .A(net71),
    .Y(_0386_));
 sg13g2_a21o_1 _2528_ (.A2(_0385_),
    .A1(net62),
    .B1(net71),
    .X(_0388_));
 sg13g2_and2_1 _2529_ (.A(_0386_),
    .B(_0388_),
    .X(_0058_));
 sg13g2_nand2_1 _2530_ (.Y(_0389_),
    .A(\perceptron1.we2[11] ),
    .B(net259));
 sg13g2_or2_1 _2531_ (.X(_0390_),
    .B(net259),
    .A(\perceptron1.we2[11] ));
 sg13g2_nand2_1 _2532_ (.Y(_0391_),
    .A(_0389_),
    .B(_0390_));
 sg13g2_xor2_1 _2533_ (.B(_0391_),
    .A(_0386_),
    .X(_0059_));
 sg13g2_nand2_1 _2534_ (.Y(_0392_),
    .A(\perceptron1.we2[12] ),
    .B(net259));
 sg13g2_xor2_1 _2535_ (.B(net259),
    .A(\perceptron1.we2[12] ),
    .X(_0393_));
 sg13g2_nand2_1 _2536_ (.Y(_0394_),
    .A(_0386_),
    .B(_0389_));
 sg13g2_nand3_1 _2537_ (.B(_0393_),
    .C(_0394_),
    .A(_0390_),
    .Y(_0395_));
 sg13g2_a21o_1 _2538_ (.A2(_0394_),
    .A1(_0390_),
    .B1(_0393_),
    .X(_0397_));
 sg13g2_and2_1 _2539_ (.A(_0395_),
    .B(_0397_),
    .X(_0060_));
 sg13g2_a21oi_2 _2540_ (.B1(_0003_),
    .Y(_0398_),
    .A2(_0395_),
    .A1(_0392_));
 sg13g2_and3_1 _2541_ (.X(_0399_),
    .A(_0003_),
    .B(_0392_),
    .C(_0395_));
 sg13g2_nor3_1 _2542_ (.A(net264),
    .B(_0398_),
    .C(_0399_),
    .Y(_0400_));
 sg13g2_a21o_1 _2543_ (.A2(net264),
    .A1(net57),
    .B1(_0400_),
    .X(_0061_));
 sg13g2_nand2_1 _2544_ (.Y(_0401_),
    .A(\perceptron1.we2[14] ),
    .B(_0398_));
 sg13g2_xor2_1 _2545_ (.B(_0398_),
    .A(net47),
    .X(_0062_));
 sg13g2_xnor2_1 _2546_ (.Y(_0063_),
    .A(net41),
    .B(_0401_));
 sg13g2_dfrbp_1 _2547_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net341),
    .D(_0016_),
    .Q_N(_0006_),
    .Q(\perceptron1.we3[0] ));
 sg13g2_dfrbp_1 _2548_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net342),
    .D(net33),
    .Q_N(\perceptron1.we3[1] ),
    .Q(_0008_));
 sg13g2_dfrbp_1 _2549_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net341),
    .D(_0018_),
    .Q_N(\perceptron1.we3[2] ),
    .Q(_0009_));
 sg13g2_dfrbp_1 _2550_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net341),
    .D(_0019_),
    .Q_N(\perceptron1.we3[3] ),
    .Q(_0010_));
 sg13g2_dfrbp_1 _2551_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net340),
    .D(_0020_),
    .Q_N(\perceptron1.we3[4] ),
    .Q(_0011_));
 sg13g2_dfrbp_1 _2552_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net340),
    .D(_0021_),
    .Q_N(_1296_),
    .Q(\perceptron1.we3[5] ));
 sg13g2_dfrbp_1 _2553_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net339),
    .D(_0022_),
    .Q_N(_1295_),
    .Q(\perceptron1.we3[6] ));
 sg13g2_dfrbp_1 _2554_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net339),
    .D(_0023_),
    .Q_N(_1294_),
    .Q(\perceptron1.we3[7] ));
 sg13g2_dfrbp_1 _2555_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net340),
    .D(_0024_),
    .Q_N(_1293_),
    .Q(\perceptron1.we3[8] ));
 sg13g2_dfrbp_1 _2556_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net342),
    .D(_0025_),
    .Q_N(_1292_),
    .Q(\perceptron1.we3[9] ));
 sg13g2_dfrbp_1 _2557_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net340),
    .D(_0026_),
    .Q_N(_1291_),
    .Q(\perceptron1.we3[10] ));
 sg13g2_dfrbp_1 _2558_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net340),
    .D(_0027_),
    .Q_N(_1290_),
    .Q(\perceptron1.we3[11] ));
 sg13g2_dfrbp_1 _2559_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net338),
    .D(_0028_),
    .Q_N(_1289_),
    .Q(\perceptron1.we3[12] ));
 sg13g2_dfrbp_1 _2560_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net338),
    .D(_0029_),
    .Q_N(_0007_),
    .Q(\perceptron1.we3[13] ));
 sg13g2_dfrbp_1 _2561_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net339),
    .D(net44),
    .Q_N(_1288_),
    .Q(\perceptron1.we3[14] ));
 sg13g2_dfrbp_1 _2562_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net339),
    .D(net39),
    .Q_N(_1287_),
    .Q(\perceptron1.we3[15] ));
 sg13g2_dfrbp_1 _2563_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net341),
    .D(net56),
    .Q_N(_0004_),
    .Q(\perceptron1.we1[0] ));
 sg13g2_dfrbp_1 _2564_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net341),
    .D(net31),
    .Q_N(\perceptron1.we1[1] ),
    .Q(_0012_));
 sg13g2_dfrbp_1 _2565_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net341),
    .D(_0034_),
    .Q_N(_1286_),
    .Q(\perceptron1.we1[2] ));
 sg13g2_dfrbp_1 _2566_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net341),
    .D(_0035_),
    .Q_N(\perceptron1.we1[3] ),
    .Q(_0013_));
 sg13g2_dfrbp_1 _2567_ (.CLK(clknet_3_2__leaf_clk),
    .RESET_B(net341),
    .D(_0036_),
    .Q_N(_1285_),
    .Q(\perceptron1.we1[4] ));
 sg13g2_dfrbp_1 _2568_ (.CLK(clknet_3_4__leaf_clk),
    .RESET_B(net340),
    .D(_0037_),
    .Q_N(_1284_),
    .Q(\perceptron1.we1[5] ));
 sg13g2_dfrbp_1 _2569_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net339),
    .D(_0038_),
    .Q_N(_1283_),
    .Q(\perceptron1.we1[6] ));
 sg13g2_dfrbp_1 _2570_ (.CLK(clknet_3_3__leaf_clk),
    .RESET_B(net340),
    .D(net81),
    .Q_N(_1282_),
    .Q(\perceptron1.we1[7] ));
 sg13g2_dfrbp_1 _2571_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net339),
    .D(_0040_),
    .Q_N(_1281_),
    .Q(\perceptron1.we1[8] ));
 sg13g2_dfrbp_1 _2572_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net338),
    .D(net68),
    .Q_N(_1280_),
    .Q(\perceptron1.we1[9] ));
 sg13g2_dfrbp_1 _2573_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net338),
    .D(net64),
    .Q_N(_1279_),
    .Q(\perceptron1.we1[10] ));
 sg13g2_dfrbp_1 _2574_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net338),
    .D(_0043_),
    .Q_N(_1278_),
    .Q(\perceptron1.we1[11] ));
 sg13g2_dfrbp_1 _2575_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net338),
    .D(_0044_),
    .Q_N(_1277_),
    .Q(\perceptron1.we1[12] ));
 sg13g2_dfrbp_1 _2576_ (.CLK(clknet_3_1__leaf_clk),
    .RESET_B(net338),
    .D(_0045_),
    .Q_N(_0005_),
    .Q(\perceptron1.we1[13] ));
 sg13g2_dfrbp_1 _2577_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net338),
    .D(net46),
    .Q_N(_1276_),
    .Q(\perceptron1.we1[14] ));
 sg13g2_dfrbp_1 _2578_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net339),
    .D(net37),
    .Q_N(_1297_),
    .Q(\perceptron1.we1[15] ));
 sg13g2_dfrbp_1 _2579_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net343),
    .D(_0000_),
    .Q_N(_1275_),
    .Q(\perceptron1.out ));
 sg13g2_dfrbp_1 _2580_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net343),
    .D(net52),
    .Q_N(_0002_),
    .Q(\perceptron1.we2[0] ));
 sg13g2_dfrbp_1 _2581_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net343),
    .D(net54),
    .Q_N(_0001_),
    .Q(\perceptron1.we2[1] ));
 sg13g2_dfrbp_1 _2582_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net343),
    .D(net27),
    .Q_N(\perceptron1.we2[2] ),
    .Q(_0014_));
 sg13g2_dfrbp_1 _2583_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net345),
    .D(net85),
    .Q_N(_1274_),
    .Q(\perceptron1.we2[3] ));
 sg13g2_dfrbp_1 _2584_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net343),
    .D(_0052_),
    .Q_N(\perceptron1.we2[4] ),
    .Q(_0015_));
 sg13g2_dfrbp_1 _2585_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net343),
    .D(net66),
    .Q_N(_1273_),
    .Q(\perceptron1.we2[5] ));
 sg13g2_dfrbp_1 _2586_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net343),
    .D(net60),
    .Q_N(_1272_),
    .Q(\perceptron1.we2[6] ));
 sg13g2_dfrbp_1 _2587_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net343),
    .D(_0055_),
    .Q_N(_1271_),
    .Q(\perceptron1.we2[7] ));
 sg13g2_dfrbp_1 _2588_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net344),
    .D(_0056_),
    .Q_N(_1270_),
    .Q(\perceptron1.we2[8] ));
 sg13g2_dfrbp_1 _2589_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net344),
    .D(_0057_),
    .Q_N(_1269_),
    .Q(\perceptron1.we2[9] ));
 sg13g2_dfrbp_1 _2590_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net344),
    .D(_0058_),
    .Q_N(_1268_),
    .Q(\perceptron1.we2[10] ));
 sg13g2_dfrbp_1 _2591_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net344),
    .D(net72),
    .Q_N(_1267_),
    .Q(\perceptron1.we2[11] ));
 sg13g2_dfrbp_1 _2592_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net344),
    .D(_0060_),
    .Q_N(_1266_),
    .Q(\perceptron1.we2[12] ));
 sg13g2_dfrbp_1 _2593_ (.CLK(clknet_3_5__leaf_clk),
    .RESET_B(net344),
    .D(net58),
    .Q_N(_0003_),
    .Q(\perceptron1.we2[13] ));
 sg13g2_dfrbp_1 _2594_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net344),
    .D(net48),
    .Q_N(_1265_),
    .Q(\perceptron1.we2[14] ));
 sg13g2_dfrbp_1 _2595_ (.CLK(clknet_3_7__leaf_clk),
    .RESET_B(net344),
    .D(net42),
    .Q_N(_1264_),
    .Q(\perceptron1.we2[15] ));
 sg13g2_tielo tt_um_Rapoport_4 (.L_LO(net4));
 sg13g2_tielo tt_um_Rapoport_5 (.L_LO(net5));
 sg13g2_tielo tt_um_Rapoport_6 (.L_LO(net6));
 sg13g2_tielo tt_um_Rapoport_7 (.L_LO(net7));
 sg13g2_tielo tt_um_Rapoport_8 (.L_LO(net8));
 sg13g2_tielo tt_um_Rapoport_9 (.L_LO(net9));
 sg13g2_tielo tt_um_Rapoport_10 (.L_LO(net10));
 sg13g2_tielo tt_um_Rapoport_11 (.L_LO(net11));
 sg13g2_tielo tt_um_Rapoport_12 (.L_LO(net12));
 sg13g2_tielo tt_um_Rapoport_13 (.L_LO(net13));
 sg13g2_tielo tt_um_Rapoport_14 (.L_LO(net14));
 sg13g2_tielo tt_um_Rapoport_15 (.L_LO(net15));
 sg13g2_tielo tt_um_Rapoport_16 (.L_LO(net16));
 sg13g2_tielo tt_um_Rapoport_17 (.L_LO(net17));
 sg13g2_tielo tt_um_Rapoport_18 (.L_LO(net18));
 sg13g2_tielo tt_um_Rapoport_19 (.L_LO(net19));
 sg13g2_tielo tt_um_Rapoport_20 (.L_LO(net20));
 sg13g2_tielo tt_um_Rapoport_21 (.L_LO(net21));
 sg13g2_tielo tt_um_Rapoport_22 (.L_LO(net22));
 sg13g2_tielo tt_um_Rapoport_23 (.L_LO(net23));
 sg13g2_tielo tt_um_Rapoport_24 (.L_LO(net24));
 sg13g2_tielo tt_um_Rapoport_25 (.L_LO(net25));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _2619_ (.A(\perceptron1.out ),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout259 (.A(_0366_),
    .X(net259));
 sg13g2_buf_1 fanout260 (.A(_0366_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(net262),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_0308_),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(net264));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_0167_));
 sg13g2_buf_2 fanout265 (.A(net266),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(net267),
    .X(net266));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(net268));
 sg13g2_buf_2 fanout268 (.A(_0168_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(net271),
    .X(net269));
 sg13g2_buf_1 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_0164_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(\perceptron1.we1[11] ),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(net74),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(\perceptron1.we1[3] ),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(net69),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(net87),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(\perceptron1.we3[8] ),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(\perceptron1.we3[7] ),
    .X(net278));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(net79));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(net73));
 sg13g2_buf_2 fanout281 (.A(\perceptron1.we3[4] ),
    .X(net281));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(\perceptron1.we3[3] ));
 sg13g2_buf_2 fanout283 (.A(\perceptron1.we3[3] ),
    .X(net283));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(\perceptron1.we3[2] ));
 sg13g2_buf_2 fanout285 (.A(\perceptron1.we3[1] ),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(\perceptron1.we3[0] ),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(uio_in[6]),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(net291),
    .X(net289));
 sg13g2_buf_1 fanout290 (.A(net291),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(uio_in[5]),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(uio_in[4]),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(uio_in[4]),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(net1),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(net1),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(net299),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(net299),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(uio_in[2]),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(net303),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(net302),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(net303),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(uio_in[1]),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(net306),
    .X(net304));
 sg13g2_buf_1 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(uio_in[0]),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(net309),
    .X(net307));
 sg13g2_buf_1 fanout308 (.A(net309),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(uio_in[0]),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(net311),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(ui_in[7]),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(net314),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net314),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(ui_in[6]),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(ui_in[5]),
    .X(net315));
 sg13g2_buf_1 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(ui_in[5]));
 sg13g2_buf_2 fanout318 (.A(net319),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(ui_in[4]),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(ui_in[4]),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(net324),
    .X(net321));
 sg13g2_buf_1 fanout322 (.A(net324),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(ui_in[3]),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(net329),
    .X(net325));
 sg13g2_buf_1 fanout326 (.A(net329),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(net329),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(net329),
    .X(net328));
 sg13g2_buf_1 fanout329 (.A(ui_in[2]),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(net332),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(net332),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(ui_in[1]),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(net335),
    .X(net333));
 sg13g2_buf_1 fanout334 (.A(net335),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(ui_in[0]),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(ui_in[0]),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(ui_in[0]),
    .X(net337));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(net339));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(net340));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(net342));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(net342));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(net345));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(net345));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(net345));
 sg13g2_buf_2 fanout345 (.A(rst_n),
    .X(net345));
 sg13g2_buf_2 input1 (.A(uio_in[3]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(uio_in[7]),
    .X(net2));
 sg13g2_tielo tt_um_Rapoport_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0014_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0050_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0013_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0009_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0012_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0033_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0008_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0017_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0010_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0015_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold11 (.A(\perceptron1.we1[15] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0047_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold13 (.A(\perceptron1.we3[15] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0031_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0011_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold16 (.A(\perceptron1.we2[15] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0063_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0007_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0030_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0005_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0046_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold22 (.A(\perceptron1.we2[14] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0062_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold24 (.A(\perceptron1.we1[13] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold25 (.A(\perceptron1.we3[13] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold26 (.A(\perceptron1.we2[0] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0048_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold28 (.A(\perceptron1.we2[1] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0049_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold30 (.A(\perceptron1.we1[0] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0032_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold32 (.A(\perceptron1.we2[13] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0061_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold34 (.A(\perceptron1.we2[6] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0054_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0006_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold37 (.A(\perceptron1.we2[9] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold38 (.A(\perceptron1.we1[10] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0042_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold40 (.A(\perceptron1.we2[5] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0053_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold42 (.A(\perceptron1.we1[9] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0041_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold44 (.A(\perceptron1.we3[10] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0274_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold46 (.A(\perceptron1.we2[10] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0059_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold48 (.A(\perceptron1.we3[5] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold49 (.A(\perceptron1.we1[5] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0004_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0305_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold52 (.A(\perceptron1.we2[8] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0383_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold54 (.A(\perceptron1.we3[6] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold55 (.A(\perceptron1.we1[6] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0039_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold57 (.A(\perceptron1.we3[12] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold58 (.A(\perceptron1.we2[7] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold59 (.A(\perceptron1.we2[2] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0051_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold61 (.A(\perceptron1.we3[11] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold62 (.A(\perceptron1.we3[9] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold63 (.A(\perceptron1.we1[12] ),
    .X(net88));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_4 FILLER_1_77 ();
 sg13g2_fill_1 FILLER_1_81 ();
 sg13g2_decap_8 FILLER_1_90 ();
 sg13g2_decap_8 FILLER_1_97 ();
 sg13g2_decap_8 FILLER_1_104 ();
 sg13g2_decap_8 FILLER_1_111 ();
 sg13g2_decap_8 FILLER_1_118 ();
 sg13g2_decap_8 FILLER_1_125 ();
 sg13g2_decap_8 FILLER_1_132 ();
 sg13g2_decap_8 FILLER_1_139 ();
 sg13g2_decap_8 FILLER_1_146 ();
 sg13g2_decap_8 FILLER_1_153 ();
 sg13g2_decap_8 FILLER_1_160 ();
 sg13g2_decap_8 FILLER_1_167 ();
 sg13g2_decap_8 FILLER_1_174 ();
 sg13g2_decap_8 FILLER_1_181 ();
 sg13g2_decap_8 FILLER_1_188 ();
 sg13g2_decap_8 FILLER_1_195 ();
 sg13g2_decap_8 FILLER_1_202 ();
 sg13g2_decap_8 FILLER_1_209 ();
 sg13g2_decap_8 FILLER_1_216 ();
 sg13g2_decap_8 FILLER_1_223 ();
 sg13g2_decap_8 FILLER_1_230 ();
 sg13g2_decap_8 FILLER_1_237 ();
 sg13g2_decap_8 FILLER_1_244 ();
 sg13g2_decap_8 FILLER_1_251 ();
 sg13g2_decap_8 FILLER_1_258 ();
 sg13g2_decap_8 FILLER_1_265 ();
 sg13g2_decap_8 FILLER_1_272 ();
 sg13g2_decap_8 FILLER_1_279 ();
 sg13g2_decap_8 FILLER_1_286 ();
 sg13g2_decap_8 FILLER_1_293 ();
 sg13g2_decap_8 FILLER_1_300 ();
 sg13g2_decap_8 FILLER_1_307 ();
 sg13g2_decap_8 FILLER_1_314 ();
 sg13g2_decap_8 FILLER_1_321 ();
 sg13g2_decap_8 FILLER_1_328 ();
 sg13g2_decap_8 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_342 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_fill_2 FILLER_2_42 ();
 sg13g2_fill_1 FILLER_2_44 ();
 sg13g2_fill_2 FILLER_2_53 ();
 sg13g2_fill_1 FILLER_2_55 ();
 sg13g2_fill_1 FILLER_2_60 ();
 sg13g2_fill_2 FILLER_2_70 ();
 sg13g2_fill_1 FILLER_2_72 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_fill_2 FILLER_2_97 ();
 sg13g2_decap_4 FILLER_2_108 ();
 sg13g2_fill_2 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_122 ();
 sg13g2_decap_8 FILLER_2_129 ();
 sg13g2_decap_8 FILLER_2_136 ();
 sg13g2_decap_8 FILLER_2_143 ();
 sg13g2_decap_8 FILLER_2_150 ();
 sg13g2_fill_2 FILLER_2_157 ();
 sg13g2_fill_1 FILLER_2_159 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_fill_2 FILLER_3_42 ();
 sg13g2_fill_2 FILLER_3_113 ();
 sg13g2_fill_1 FILLER_3_115 ();
 sg13g2_fill_2 FILLER_3_158 ();
 sg13g2_fill_1 FILLER_3_160 ();
 sg13g2_decap_8 FILLER_3_171 ();
 sg13g2_fill_2 FILLER_3_178 ();
 sg13g2_fill_1 FILLER_3_180 ();
 sg13g2_decap_8 FILLER_3_197 ();
 sg13g2_decap_8 FILLER_3_204 ();
 sg13g2_decap_4 FILLER_3_211 ();
 sg13g2_fill_1 FILLER_3_215 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_4 FILLER_4_28 ();
 sg13g2_fill_1 FILLER_4_32 ();
 sg13g2_decap_4 FILLER_4_67 ();
 sg13g2_fill_1 FILLER_4_80 ();
 sg13g2_decap_8 FILLER_4_107 ();
 sg13g2_fill_2 FILLER_4_114 ();
 sg13g2_decap_4 FILLER_4_124 ();
 sg13g2_fill_1 FILLER_4_128 ();
 sg13g2_fill_1 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_146 ();
 sg13g2_fill_2 FILLER_4_153 ();
 sg13g2_fill_1 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_198 ();
 sg13g2_decap_8 FILLER_4_205 ();
 sg13g2_fill_1 FILLER_4_212 ();
 sg13g2_decap_8 FILLER_4_229 ();
 sg13g2_decap_8 FILLER_4_236 ();
 sg13g2_decap_8 FILLER_4_243 ();
 sg13g2_decap_8 FILLER_4_250 ();
 sg13g2_decap_8 FILLER_4_257 ();
 sg13g2_decap_8 FILLER_4_264 ();
 sg13g2_decap_8 FILLER_4_271 ();
 sg13g2_decap_8 FILLER_4_278 ();
 sg13g2_decap_8 FILLER_4_285 ();
 sg13g2_decap_8 FILLER_4_292 ();
 sg13g2_decap_8 FILLER_4_299 ();
 sg13g2_decap_8 FILLER_4_306 ();
 sg13g2_decap_8 FILLER_4_313 ();
 sg13g2_decap_8 FILLER_4_320 ();
 sg13g2_decap_8 FILLER_4_327 ();
 sg13g2_decap_8 FILLER_4_334 ();
 sg13g2_decap_8 FILLER_4_341 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_decap_8 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_fill_1 FILLER_5_47 ();
 sg13g2_decap_4 FILLER_5_58 ();
 sg13g2_fill_2 FILLER_5_62 ();
 sg13g2_fill_2 FILLER_5_68 ();
 sg13g2_fill_2 FILLER_5_79 ();
 sg13g2_fill_1 FILLER_5_90 ();
 sg13g2_fill_1 FILLER_5_119 ();
 sg13g2_fill_2 FILLER_5_139 ();
 sg13g2_decap_8 FILLER_5_160 ();
 sg13g2_decap_4 FILLER_5_171 ();
 sg13g2_fill_2 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_202 ();
 sg13g2_fill_1 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_fill_2 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_16 ();
 sg13g2_fill_2 FILLER_6_39 ();
 sg13g2_fill_1 FILLER_6_115 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_137 ();
 sg13g2_fill_2 FILLER_6_172 ();
 sg13g2_fill_2 FILLER_6_190 ();
 sg13g2_fill_1 FILLER_6_192 ();
 sg13g2_decap_8 FILLER_6_202 ();
 sg13g2_fill_2 FILLER_6_209 ();
 sg13g2_decap_8 FILLER_6_223 ();
 sg13g2_fill_2 FILLER_6_230 ();
 sg13g2_fill_1 FILLER_6_232 ();
 sg13g2_decap_8 FILLER_6_267 ();
 sg13g2_decap_4 FILLER_6_274 ();
 sg13g2_fill_1 FILLER_6_278 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_4 FILLER_7_14 ();
 sg13g2_decap_4 FILLER_7_55 ();
 sg13g2_fill_2 FILLER_7_68 ();
 sg13g2_fill_1 FILLER_7_88 ();
 sg13g2_decap_4 FILLER_7_98 ();
 sg13g2_decap_4 FILLER_7_132 ();
 sg13g2_fill_2 FILLER_7_148 ();
 sg13g2_fill_2 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_166 ();
 sg13g2_decap_4 FILLER_7_173 ();
 sg13g2_fill_1 FILLER_7_177 ();
 sg13g2_decap_4 FILLER_7_182 ();
 sg13g2_fill_1 FILLER_7_194 ();
 sg13g2_fill_1 FILLER_7_200 ();
 sg13g2_fill_2 FILLER_7_214 ();
 sg13g2_decap_8 FILLER_7_248 ();
 sg13g2_fill_2 FILLER_7_255 ();
 sg13g2_decap_4 FILLER_7_265 ();
 sg13g2_fill_2 FILLER_7_269 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_4 FILLER_8_38 ();
 sg13g2_fill_1 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_fill_2 FILLER_8_105 ();
 sg13g2_fill_1 FILLER_8_107 ();
 sg13g2_fill_1 FILLER_8_116 ();
 sg13g2_decap_4 FILLER_8_141 ();
 sg13g2_fill_2 FILLER_8_153 ();
 sg13g2_fill_1 FILLER_8_155 ();
 sg13g2_decap_8 FILLER_8_174 ();
 sg13g2_decap_4 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_201 ();
 sg13g2_decap_8 FILLER_8_208 ();
 sg13g2_fill_2 FILLER_8_215 ();
 sg13g2_fill_1 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_4 FILLER_8_237 ();
 sg13g2_fill_2 FILLER_8_253 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_fill_2 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_4 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_55 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_128 ();
 sg13g2_fill_2 FILLER_9_135 ();
 sg13g2_fill_2 FILLER_9_149 ();
 sg13g2_fill_1 FILLER_9_151 ();
 sg13g2_fill_2 FILLER_9_172 ();
 sg13g2_fill_1 FILLER_9_186 ();
 sg13g2_fill_1 FILLER_9_195 ();
 sg13g2_decap_4 FILLER_9_201 ();
 sg13g2_fill_2 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_decap_4 FILLER_9_244 ();
 sg13g2_fill_1 FILLER_9_248 ();
 sg13g2_fill_1 FILLER_9_262 ();
 sg13g2_decap_4 FILLER_9_271 ();
 sg13g2_decap_4 FILLER_9_300 ();
 sg13g2_fill_1 FILLER_9_304 ();
 sg13g2_decap_8 FILLER_9_313 ();
 sg13g2_decap_8 FILLER_9_320 ();
 sg13g2_fill_1 FILLER_9_327 ();
 sg13g2_decap_4 FILLER_9_346 ();
 sg13g2_fill_2 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_11 ();
 sg13g2_fill_2 FILLER_10_57 ();
 sg13g2_fill_1 FILLER_10_59 ();
 sg13g2_fill_2 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_110 ();
 sg13g2_decap_8 FILLER_10_134 ();
 sg13g2_decap_4 FILLER_10_141 ();
 sg13g2_fill_2 FILLER_10_145 ();
 sg13g2_decap_4 FILLER_10_151 ();
 sg13g2_fill_2 FILLER_10_155 ();
 sg13g2_fill_1 FILLER_10_186 ();
 sg13g2_fill_1 FILLER_10_192 ();
 sg13g2_fill_2 FILLER_10_213 ();
 sg13g2_fill_1 FILLER_10_215 ();
 sg13g2_decap_8 FILLER_10_232 ();
 sg13g2_decap_8 FILLER_10_239 ();
 sg13g2_fill_2 FILLER_10_246 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_fill_2 FILLER_10_321 ();
 sg13g2_fill_1 FILLER_10_323 ();
 sg13g2_decap_4 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_4 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_113 ();
 sg13g2_fill_2 FILLER_11_165 ();
 sg13g2_fill_1 FILLER_11_167 ();
 sg13g2_fill_2 FILLER_11_181 ();
 sg13g2_decap_4 FILLER_11_188 ();
 sg13g2_decap_4 FILLER_11_201 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_249 ();
 sg13g2_fill_1 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_264 ();
 sg13g2_decap_4 FILLER_11_300 ();
 sg13g2_fill_2 FILLER_11_316 ();
 sg13g2_fill_1 FILLER_11_330 ();
 sg13g2_fill_2 FILLER_11_337 ();
 sg13g2_decap_4 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_4 FILLER_12_21 ();
 sg13g2_fill_2 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_63 ();
 sg13g2_fill_1 FILLER_12_65 ();
 sg13g2_decap_4 FILLER_12_94 ();
 sg13g2_fill_1 FILLER_12_124 ();
 sg13g2_fill_2 FILLER_12_163 ();
 sg13g2_fill_2 FILLER_12_170 ();
 sg13g2_fill_1 FILLER_12_172 ();
 sg13g2_fill_2 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_fill_1 FILLER_12_220 ();
 sg13g2_decap_4 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_290 ();
 sg13g2_decap_4 FILLER_12_297 ();
 sg13g2_fill_1 FILLER_12_301 ();
 sg13g2_fill_2 FILLER_12_306 ();
 sg13g2_decap_4 FILLER_12_317 ();
 sg13g2_fill_1 FILLER_12_321 ();
 sg13g2_fill_2 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_60 ();
 sg13g2_fill_1 FILLER_13_62 ();
 sg13g2_decap_4 FILLER_13_110 ();
 sg13g2_decap_8 FILLER_13_138 ();
 sg13g2_fill_2 FILLER_13_145 ();
 sg13g2_fill_2 FILLER_13_157 ();
 sg13g2_decap_8 FILLER_13_173 ();
 sg13g2_fill_2 FILLER_13_180 ();
 sg13g2_fill_1 FILLER_13_187 ();
 sg13g2_decap_4 FILLER_13_201 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_fill_2 FILLER_13_227 ();
 sg13g2_fill_1 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_fill_2 FILLER_13_250 ();
 sg13g2_fill_1 FILLER_13_252 ();
 sg13g2_decap_4 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_267 ();
 sg13g2_decap_4 FILLER_13_281 ();
 sg13g2_fill_2 FILLER_13_285 ();
 sg13g2_decap_4 FILLER_13_292 ();
 sg13g2_fill_1 FILLER_13_296 ();
 sg13g2_decap_4 FILLER_13_312 ();
 sg13g2_fill_2 FILLER_13_338 ();
 sg13g2_decap_4 FILLER_13_360 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_30 ();
 sg13g2_decap_8 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_46 ();
 sg13g2_decap_8 FILLER_14_53 ();
 sg13g2_decap_4 FILLER_14_60 ();
 sg13g2_fill_2 FILLER_14_64 ();
 sg13g2_decap_4 FILLER_14_85 ();
 sg13g2_fill_1 FILLER_14_89 ();
 sg13g2_decap_8 FILLER_14_106 ();
 sg13g2_decap_4 FILLER_14_113 ();
 sg13g2_decap_4 FILLER_14_131 ();
 sg13g2_fill_1 FILLER_14_135 ();
 sg13g2_decap_8 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_fill_1 FILLER_14_239 ();
 sg13g2_fill_1 FILLER_14_248 ();
 sg13g2_fill_2 FILLER_14_264 ();
 sg13g2_decap_4 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_317 ();
 sg13g2_decap_4 FILLER_14_322 ();
 sg13g2_decap_4 FILLER_14_339 ();
 sg13g2_fill_2 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_fill_2 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_61 ();
 sg13g2_fill_2 FILLER_15_77 ();
 sg13g2_fill_1 FILLER_15_79 ();
 sg13g2_fill_2 FILLER_15_115 ();
 sg13g2_fill_1 FILLER_15_117 ();
 sg13g2_decap_8 FILLER_15_132 ();
 sg13g2_decap_4 FILLER_15_139 ();
 sg13g2_decap_4 FILLER_15_149 ();
 sg13g2_decap_8 FILLER_15_171 ();
 sg13g2_decap_4 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_182 ();
 sg13g2_fill_1 FILLER_15_192 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_4 FILLER_15_204 ();
 sg13g2_fill_1 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_237 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_fill_2 FILLER_15_272 ();
 sg13g2_fill_1 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_fill_1 FILLER_15_301 ();
 sg13g2_fill_2 FILLER_15_321 ();
 sg13g2_fill_2 FILLER_15_342 ();
 sg13g2_fill_2 FILLER_15_362 ();
 sg13g2_fill_2 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_48 ();
 sg13g2_fill_2 FILLER_16_55 ();
 sg13g2_fill_1 FILLER_16_57 ();
 sg13g2_decap_4 FILLER_16_92 ();
 sg13g2_fill_1 FILLER_16_96 ();
 sg13g2_fill_1 FILLER_16_114 ();
 sg13g2_fill_2 FILLER_16_155 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_2 FILLER_16_168 ();
 sg13g2_fill_1 FILLER_16_170 ();
 sg13g2_fill_1 FILLER_16_184 ();
 sg13g2_fill_2 FILLER_16_198 ();
 sg13g2_fill_1 FILLER_16_200 ();
 sg13g2_fill_2 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_237 ();
 sg13g2_fill_1 FILLER_16_250 ();
 sg13g2_fill_2 FILLER_16_261 ();
 sg13g2_fill_1 FILLER_16_263 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_decap_4 FILLER_16_302 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_4 FILLER_16_345 ();
 sg13g2_fill_2 FILLER_16_374 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_2 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_30 ();
 sg13g2_fill_1 FILLER_17_65 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_93 ();
 sg13g2_decap_4 FILLER_17_102 ();
 sg13g2_fill_2 FILLER_17_106 ();
 sg13g2_fill_2 FILLER_17_116 ();
 sg13g2_fill_2 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_125 ();
 sg13g2_decap_8 FILLER_17_135 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_fill_2 FILLER_17_146 ();
 sg13g2_decap_8 FILLER_17_158 ();
 sg13g2_fill_1 FILLER_17_165 ();
 sg13g2_decap_4 FILLER_17_176 ();
 sg13g2_fill_1 FILLER_17_180 ();
 sg13g2_fill_1 FILLER_17_185 ();
 sg13g2_decap_4 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_decap_4 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_decap_8 FILLER_17_261 ();
 sg13g2_fill_2 FILLER_17_268 ();
 sg13g2_decap_4 FILLER_17_275 ();
 sg13g2_fill_2 FILLER_17_279 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_fill_1 FILLER_17_293 ();
 sg13g2_fill_2 FILLER_17_302 ();
 sg13g2_fill_1 FILLER_17_309 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_4 FILLER_17_346 ();
 sg13g2_fill_2 FILLER_17_359 ();
 sg13g2_fill_1 FILLER_17_361 ();
 sg13g2_fill_2 FILLER_17_372 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_57 ();
 sg13g2_fill_1 FILLER_18_59 ();
 sg13g2_fill_1 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_decap_4 FILLER_18_166 ();
 sg13g2_fill_2 FILLER_18_178 ();
 sg13g2_fill_1 FILLER_18_180 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_decap_4 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_235 ();
 sg13g2_fill_2 FILLER_18_276 ();
 sg13g2_decap_4 FILLER_18_286 ();
 sg13g2_fill_2 FILLER_18_327 ();
 sg13g2_fill_1 FILLER_18_329 ();
 sg13g2_fill_2 FILLER_18_335 ();
 sg13g2_fill_1 FILLER_18_337 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_fill_2 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_51 ();
 sg13g2_fill_2 FILLER_19_103 ();
 sg13g2_decap_4 FILLER_19_110 ();
 sg13g2_fill_1 FILLER_19_114 ();
 sg13g2_fill_2 FILLER_19_124 ();
 sg13g2_fill_2 FILLER_19_143 ();
 sg13g2_decap_4 FILLER_19_159 ();
 sg13g2_fill_1 FILLER_19_163 ();
 sg13g2_fill_1 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_224 ();
 sg13g2_decap_4 FILLER_19_230 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_fill_2 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_250 ();
 sg13g2_decap_4 FILLER_19_256 ();
 sg13g2_fill_1 FILLER_19_265 ();
 sg13g2_decap_4 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_316 ();
 sg13g2_decap_4 FILLER_19_323 ();
 sg13g2_fill_2 FILLER_19_331 ();
 sg13g2_fill_1 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_339 ();
 sg13g2_decap_8 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_376 ();
 sg13g2_fill_1 FILLER_19_395 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_4 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_59 ();
 sg13g2_fill_1 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_83 ();
 sg13g2_fill_2 FILLER_20_90 ();
 sg13g2_fill_1 FILLER_20_100 ();
 sg13g2_fill_2 FILLER_20_115 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_decap_4 FILLER_20_122 ();
 sg13g2_decap_4 FILLER_20_136 ();
 sg13g2_decap_4 FILLER_20_145 ();
 sg13g2_fill_1 FILLER_20_149 ();
 sg13g2_decap_4 FILLER_20_155 ();
 sg13g2_fill_1 FILLER_20_159 ();
 sg13g2_decap_4 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_decap_4 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_223 ();
 sg13g2_decap_8 FILLER_20_232 ();
 sg13g2_fill_2 FILLER_20_239 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_fill_2 FILLER_20_273 ();
 sg13g2_fill_1 FILLER_20_289 ();
 sg13g2_fill_2 FILLER_20_298 ();
 sg13g2_decap_4 FILLER_20_321 ();
 sg13g2_fill_1 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_37 ();
 sg13g2_decap_4 FILLER_21_47 ();
 sg13g2_fill_1 FILLER_21_51 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_108 ();
 sg13g2_fill_1 FILLER_21_115 ();
 sg13g2_fill_2 FILLER_21_136 ();
 sg13g2_fill_1 FILLER_21_150 ();
 sg13g2_decap_4 FILLER_21_159 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_170 ();
 sg13g2_fill_1 FILLER_21_179 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_decap_4 FILLER_21_214 ();
 sg13g2_fill_1 FILLER_21_218 ();
 sg13g2_fill_1 FILLER_21_228 ();
 sg13g2_fill_2 FILLER_21_270 ();
 sg13g2_fill_1 FILLER_21_272 ();
 sg13g2_decap_8 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_317 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_decap_4 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_decap_4 FILLER_21_360 ();
 sg13g2_decap_4 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_14 ();
 sg13g2_fill_1 FILLER_22_16 ();
 sg13g2_fill_2 FILLER_22_60 ();
 sg13g2_fill_1 FILLER_22_62 ();
 sg13g2_fill_1 FILLER_22_71 ();
 sg13g2_fill_2 FILLER_22_82 ();
 sg13g2_fill_1 FILLER_22_99 ();
 sg13g2_fill_2 FILLER_22_120 ();
 sg13g2_fill_2 FILLER_22_131 ();
 sg13g2_fill_1 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_fill_1 FILLER_22_151 ();
 sg13g2_decap_4 FILLER_22_156 ();
 sg13g2_fill_1 FILLER_22_160 ();
 sg13g2_fill_2 FILLER_22_166 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_181 ();
 sg13g2_decap_4 FILLER_22_188 ();
 sg13g2_fill_2 FILLER_22_192 ();
 sg13g2_decap_8 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_209 ();
 sg13g2_fill_2 FILLER_22_216 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_decap_4 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_4 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_4 FILLER_22_282 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_4 FILLER_22_308 ();
 sg13g2_fill_2 FILLER_22_312 ();
 sg13g2_decap_4 FILLER_22_327 ();
 sg13g2_decap_4 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_388 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_51 ();
 sg13g2_fill_1 FILLER_23_61 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_fill_1 FILLER_23_92 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_fill_1 FILLER_23_119 ();
 sg13g2_decap_4 FILLER_23_124 ();
 sg13g2_fill_2 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_fill_2 FILLER_23_158 ();
 sg13g2_fill_1 FILLER_23_160 ();
 sg13g2_fill_2 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_181 ();
 sg13g2_decap_4 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_207 ();
 sg13g2_fill_1 FILLER_23_209 ();
 sg13g2_fill_2 FILLER_23_228 ();
 sg13g2_fill_1 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_239 ();
 sg13g2_decap_4 FILLER_23_248 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_259 ();
 sg13g2_fill_1 FILLER_23_261 ();
 sg13g2_fill_2 FILLER_23_286 ();
 sg13g2_fill_2 FILLER_23_310 ();
 sg13g2_fill_1 FILLER_23_336 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_fill_1 FILLER_23_362 ();
 sg13g2_fill_1 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_61 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_4 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_fill_2 FILLER_24_128 ();
 sg13g2_decap_4 FILLER_24_141 ();
 sg13g2_fill_2 FILLER_24_145 ();
 sg13g2_fill_2 FILLER_24_157 ();
 sg13g2_fill_2 FILLER_24_164 ();
 sg13g2_decap_8 FILLER_24_171 ();
 sg13g2_decap_4 FILLER_24_178 ();
 sg13g2_fill_2 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_fill_2 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_226 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_fill_2 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_fill_2 FILLER_24_332 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_349 ();
 sg13g2_decap_4 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_fill_1 FILLER_24_378 ();
 sg13g2_decap_4 FILLER_24_395 ();
 sg13g2_fill_2 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_52 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_79 ();
 sg13g2_fill_2 FILLER_25_86 ();
 sg13g2_fill_2 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_117 ();
 sg13g2_fill_1 FILLER_25_127 ();
 sg13g2_fill_2 FILLER_25_148 ();
 sg13g2_fill_1 FILLER_25_164 ();
 sg13g2_decap_4 FILLER_25_179 ();
 sg13g2_fill_2 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_decap_8 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_262 ();
 sg13g2_fill_1 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_decap_4 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_300 ();
 sg13g2_fill_2 FILLER_25_346 ();
 sg13g2_decap_4 FILLER_25_353 ();
 sg13g2_fill_1 FILLER_25_357 ();
 sg13g2_fill_1 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_50 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_4 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_185 ();
 sg13g2_decap_8 FILLER_26_222 ();
 sg13g2_decap_4 FILLER_26_233 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_fill_2 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_293 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_23 ();
 sg13g2_fill_2 FILLER_27_34 ();
 sg13g2_fill_1 FILLER_27_36 ();
 sg13g2_decap_4 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_46 ();
 sg13g2_fill_2 FILLER_27_58 ();
 sg13g2_fill_1 FILLER_27_60 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_fill_2 FILLER_27_115 ();
 sg13g2_decap_4 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_161 ();
 sg13g2_decap_4 FILLER_27_183 ();
 sg13g2_fill_2 FILLER_27_187 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_fill_1 FILLER_27_206 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_261 ();
 sg13g2_decap_4 FILLER_27_288 ();
 sg13g2_fill_1 FILLER_27_292 ();
 sg13g2_fill_1 FILLER_27_310 ();
 sg13g2_decap_4 FILLER_27_316 ();
 sg13g2_fill_1 FILLER_27_320 ();
 sg13g2_fill_1 FILLER_27_353 ();
 sg13g2_fill_2 FILLER_27_369 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_fill_2 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_84 ();
 sg13g2_fill_2 FILLER_28_122 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_decap_8 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_fill_2 FILLER_28_211 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_233 ();
 sg13g2_fill_2 FILLER_28_240 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_286 ();
 sg13g2_decap_8 FILLER_28_293 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_4 FILLER_28_329 ();
 sg13g2_fill_1 FILLER_28_333 ();
 sg13g2_fill_1 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_decap_4 FILLER_28_360 ();
 sg13g2_fill_2 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_99 ();
 sg13g2_decap_4 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_decap_8 FILLER_29_125 ();
 sg13g2_decap_8 FILLER_29_132 ();
 sg13g2_decap_8 FILLER_29_149 ();
 sg13g2_decap_4 FILLER_29_186 ();
 sg13g2_fill_2 FILLER_29_195 ();
 sg13g2_decap_4 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_fill_1 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_fill_2 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_248 ();
 sg13g2_decap_8 FILLER_29_253 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_283 ();
 sg13g2_decap_4 FILLER_29_302 ();
 sg13g2_fill_2 FILLER_29_323 ();
 sg13g2_fill_2 FILLER_29_335 ();
 sg13g2_decap_4 FILLER_29_357 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_fill_1 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_fill_1 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_81 ();
 sg13g2_fill_2 FILLER_30_100 ();
 sg13g2_decap_4 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_153 ();
 sg13g2_decap_4 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_decap_8 FILLER_30_173 ();
 sg13g2_decap_4 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_decap_4 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_fill_2 FILLER_30_220 ();
 sg13g2_decap_4 FILLER_30_227 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_4 FILLER_30_242 ();
 sg13g2_fill_2 FILLER_30_272 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_4 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_25 ();
 sg13g2_decap_8 FILLER_31_52 ();
 sg13g2_fill_1 FILLER_31_59 ();
 sg13g2_decap_8 FILLER_31_65 ();
 sg13g2_decap_8 FILLER_31_72 ();
 sg13g2_decap_4 FILLER_31_79 ();
 sg13g2_fill_1 FILLER_31_83 ();
 sg13g2_fill_2 FILLER_31_99 ();
 sg13g2_fill_1 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_106 ();
 sg13g2_fill_2 FILLER_31_123 ();
 sg13g2_decap_4 FILLER_31_130 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_fill_1 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_173 ();
 sg13g2_fill_1 FILLER_31_186 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_220 ();
 sg13g2_fill_2 FILLER_31_229 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_263 ();
 sg13g2_decap_4 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_274 ();
 sg13g2_fill_2 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_283 ();
 sg13g2_decap_4 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_293 ();
 sg13g2_fill_2 FILLER_31_298 ();
 sg13g2_fill_1 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_358 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_fill_2 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_fill_2 FILLER_32_36 ();
 sg13g2_fill_1 FILLER_32_38 ();
 sg13g2_fill_2 FILLER_32_43 ();
 sg13g2_fill_1 FILLER_32_45 ();
 sg13g2_decap_8 FILLER_32_67 ();
 sg13g2_fill_2 FILLER_32_74 ();
 sg13g2_fill_1 FILLER_32_76 ();
 sg13g2_fill_2 FILLER_32_85 ();
 sg13g2_fill_1 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_fill_2 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_152 ();
 sg13g2_fill_1 FILLER_32_154 ();
 sg13g2_fill_2 FILLER_32_168 ();
 sg13g2_decap_4 FILLER_32_180 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_fill_2 FILLER_32_211 ();
 sg13g2_fill_2 FILLER_32_221 ();
 sg13g2_fill_1 FILLER_32_223 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_fill_2 FILLER_32_246 ();
 sg13g2_fill_1 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_339 ();
 sg13g2_fill_1 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_45 ();
 sg13g2_fill_1 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_113 ();
 sg13g2_decap_4 FILLER_33_120 ();
 sg13g2_decap_4 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_4 FILLER_33_245 ();
 sg13g2_decap_4 FILLER_33_257 ();
 sg13g2_fill_1 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_decap_4 FILLER_33_370 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_23 ();
 sg13g2_fill_1 FILLER_34_47 ();
 sg13g2_decap_8 FILLER_34_57 ();
 sg13g2_decap_8 FILLER_34_64 ();
 sg13g2_decap_4 FILLER_34_71 ();
 sg13g2_fill_2 FILLER_34_75 ();
 sg13g2_fill_1 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_106 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_fill_2 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_168 ();
 sg13g2_fill_2 FILLER_34_178 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_decap_4 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_194 ();
 sg13g2_decap_8 FILLER_34_199 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_decap_8 FILLER_34_218 ();
 sg13g2_decap_4 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_241 ();
 sg13g2_decap_4 FILLER_34_255 ();
 sg13g2_decap_4 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_fill_2 FILLER_34_346 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_4 FILLER_35_35 ();
 sg13g2_fill_2 FILLER_35_43 ();
 sg13g2_decap_8 FILLER_35_50 ();
 sg13g2_decap_8 FILLER_35_57 ();
 sg13g2_decap_8 FILLER_35_64 ();
 sg13g2_decap_8 FILLER_35_71 ();
 sg13g2_decap_4 FILLER_35_78 ();
 sg13g2_fill_2 FILLER_35_82 ();
 sg13g2_decap_8 FILLER_35_88 ();
 sg13g2_decap_8 FILLER_35_95 ();
 sg13g2_fill_1 FILLER_35_102 ();
 sg13g2_decap_8 FILLER_35_108 ();
 sg13g2_decap_4 FILLER_35_115 ();
 sg13g2_fill_1 FILLER_35_119 ();
 sg13g2_fill_1 FILLER_35_136 ();
 sg13g2_fill_2 FILLER_35_153 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_fill_1 FILLER_35_203 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_decap_4 FILLER_35_235 ();
 sg13g2_decap_8 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_262 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_291 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_4 FILLER_35_329 ();
 sg13g2_fill_2 FILLER_35_357 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_369 ();
 sg13g2_fill_1 FILLER_35_393 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_4 FILLER_36_119 ();
 sg13g2_fill_2 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_130 ();
 sg13g2_fill_2 FILLER_36_135 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_decap_8 FILLER_36_142 ();
 sg13g2_decap_8 FILLER_36_149 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_decap_4 FILLER_36_163 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_227 ();
 sg13g2_decap_8 FILLER_36_234 ();
 sg13g2_decap_4 FILLER_36_254 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_decap_4 FILLER_36_270 ();
 sg13g2_decap_4 FILLER_36_294 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_fill_1 FILLER_36_303 ();
 sg13g2_fill_2 FILLER_36_308 ();
 sg13g2_decap_4 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_353 ();
 sg13g2_fill_2 FILLER_36_374 ();
 sg13g2_fill_1 FILLER_36_376 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_fill_2 FILLER_37_224 ();
 sg13g2_fill_1 FILLER_37_226 ();
 sg13g2_decap_8 FILLER_37_239 ();
 sg13g2_decap_8 FILLER_37_246 ();
 sg13g2_fill_2 FILLER_37_253 ();
 sg13g2_fill_2 FILLER_37_271 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_fill_2 FILLER_37_308 ();
 sg13g2_fill_2 FILLER_37_318 ();
 sg13g2_decap_8 FILLER_37_330 ();
 sg13g2_fill_2 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_367 ();
 sg13g2_fill_1 FILLER_37_374 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_decap_4 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_decap_4 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_253 ();
 sg13g2_decap_8 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_267 ();
 sg13g2_decap_4 FILLER_38_274 ();
 sg13g2_fill_2 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_1 FILLER_38_317 ();
 sg13g2_decap_4 FILLER_38_331 ();
 sg13g2_decap_4 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_fill_2 FILLER_38_379 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uo_out[0] = net18;
 assign uo_out[1] = net19;
 assign uo_out[2] = net20;
 assign uo_out[3] = net21;
 assign uo_out[4] = net22;
 assign uo_out[5] = net23;
 assign uo_out[6] = net24;
 assign uo_out[7] = net25;
endmodule

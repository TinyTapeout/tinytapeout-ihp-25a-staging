module tt_um_toivoh_demo_tt10 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire \dtop.field_top.acc[0] ;
 wire \dtop.field_top.acc[10] ;
 wire \dtop.field_top.acc[11] ;
 wire \dtop.field_top.acc[12] ;
 wire \dtop.field_top.acc[13] ;
 wire \dtop.field_top.acc[14] ;
 wire \dtop.field_top.acc[15] ;
 wire \dtop.field_top.acc[16] ;
 wire \dtop.field_top.acc[1] ;
 wire \dtop.field_top.acc[2] ;
 wire \dtop.field_top.acc[3] ;
 wire \dtop.field_top.acc[4] ;
 wire \dtop.field_top.acc[5] ;
 wire \dtop.field_top.acc[6] ;
 wire \dtop.field_top.acc[7] ;
 wire \dtop.field_top.acc[8] ;
 wire \dtop.field_top.acc[9] ;
 wire \dtop.field_top.afl_alu.last_r_sum_msbs[0] ;
 wire \dtop.field_top.afl_alu.last_r_sum_msbs[1] ;
 wire \dtop.field_top.afl_alu.p ;
 wire \dtop.field_top.afl_pc[0] ;
 wire \dtop.field_top.afl_pc[1] ;
 wire \dtop.field_top.afl_pc[2] ;
 wire \dtop.field_top.afl_pc[3] ;
 wire \dtop.field_top.afl_pc[4] ;
 wire \dtop.field_top.afl_pc[5] ;
 wire \dtop.field_top.afl_pc[6] ;
 wire \dtop.field_top.afl_pc[7] ;
 wire \dtop.field_top.afl_pc[8] ;
 wire \dtop.field_top.afl_sub_pc[0] ;
 wire \dtop.field_top.afl_sub_pc[1] ;
 wire \dtop.field_top.alt_osc[1] ;
 wire \dtop.field_top.alt_osc[2] ;
 wire \dtop.field_top.alt_osc[3] ;
 wire \dtop.field_top.alt_osc[4] ;
 wire \dtop.field_top.alt_osc[5] ;
 wire \dtop.field_top.alt_osc[6] ;
 wire \dtop.field_top.alt_osc[7] ;
 wire \dtop.field_top.alt_osc[8] ;
 wire \dtop.field_top.channel[0] ;
 wire \dtop.field_top.channel[1] ;
 wire \dtop.field_top.channel[2] ;
 wire \dtop.field_top.channel[3] ;
 wire \dtop.field_top.channel_output[0] ;
 wire \dtop.field_top.channel_output[10] ;
 wire \dtop.field_top.channel_output[1] ;
 wire \dtop.field_top.channel_output[2] ;
 wire \dtop.field_top.channel_output[3] ;
 wire \dtop.field_top.channel_output[4] ;
 wire \dtop.field_top.channel_output[5] ;
 wire \dtop.field_top.channel_output[6] ;
 wire \dtop.field_top.channel_output[7] ;
 wire \dtop.field_top.channel_output[8] ;
 wire \dtop.field_top.channel_output[9] ;
 wire \dtop.field_top.comp_value0[0] ;
 wire \dtop.field_top.comp_value0[1] ;
 wire \dtop.field_top.comp_value0[2] ;
 wire \dtop.field_top.comp_value0[3] ;
 wire \dtop.field_top.comp_value0[4] ;
 wire \dtop.field_top.comp_value0[5] ;
 wire \dtop.field_top.comp_value0[6] ;
 wire \dtop.field_top.comp_value0[7] ;
 wire \dtop.field_top.comp_value0[8] ;
 wire \dtop.field_top.comp_value0_0[10] ;
 wire \dtop.field_top.comp_value0_1[0] ;
 wire \dtop.field_top.comp_value0_1[10] ;
 wire \dtop.field_top.comp_value0_1[1] ;
 wire \dtop.field_top.comp_value0_1[2] ;
 wire \dtop.field_top.comp_value0_1[3] ;
 wire \dtop.field_top.comp_value0_1[4] ;
 wire \dtop.field_top.comp_value0_1[5] ;
 wire \dtop.field_top.comp_value0_1[6] ;
 wire \dtop.field_top.comp_value0_1[7] ;
 wire \dtop.field_top.comp_value0_1[8] ;
 wire \dtop.field_top.comp_value0_1[9] ;
 wire \dtop.field_top.comp_values0[2][0] ;
 wire \dtop.field_top.comp_values0[2][10] ;
 wire \dtop.field_top.comp_values0[2][1] ;
 wire \dtop.field_top.comp_values0[2][2] ;
 wire \dtop.field_top.comp_values0[2][3] ;
 wire \dtop.field_top.comp_values0[2][4] ;
 wire \dtop.field_top.comp_values0[2][5] ;
 wire \dtop.field_top.comp_values0[2][6] ;
 wire \dtop.field_top.comp_values0[2][7] ;
 wire \dtop.field_top.comp_values0[2][8] ;
 wire \dtop.field_top.comp_values0[2][9] ;
 wire \dtop.field_top.comp_values0[3][0] ;
 wire \dtop.field_top.comp_values0[3][10] ;
 wire \dtop.field_top.comp_values0[3][1] ;
 wire \dtop.field_top.comp_values0[3][2] ;
 wire \dtop.field_top.comp_values0[3][3] ;
 wire \dtop.field_top.comp_values0[3][4] ;
 wire \dtop.field_top.comp_values0[3][5] ;
 wire \dtop.field_top.comp_values0[3][6] ;
 wire \dtop.field_top.comp_values0[3][7] ;
 wire \dtop.field_top.comp_values0[3][8] ;
 wire \dtop.field_top.comp_values0[3][9] ;
 wire \dtop.field_top.comp_values0[4][0] ;
 wire \dtop.field_top.comp_values0[4][10] ;
 wire \dtop.field_top.comp_values0[4][1] ;
 wire \dtop.field_top.comp_values0[4][2] ;
 wire \dtop.field_top.comp_values0[4][3] ;
 wire \dtop.field_top.comp_values0[4][4] ;
 wire \dtop.field_top.comp_values0[4][5] ;
 wire \dtop.field_top.comp_values0[4][6] ;
 wire \dtop.field_top.comp_values0[4][7] ;
 wire \dtop.field_top.comp_values0[4][8] ;
 wire \dtop.field_top.comp_values0[4][9] ;
 wire \dtop.field_top.controller.pattern0[0] ;
 wire \dtop.field_top.controller.pattern0[1] ;
 wire \dtop.field_top.controller.pattern0[2] ;
 wire \dtop.field_top.controller.ppos[0] ;
 wire \dtop.field_top.controller.ppos[1] ;
 wire \dtop.field_top.controller.ppos[2] ;
 wire \dtop.field_top.controller.ppos[3] ;
 wire \dtop.field_top.controller.ppos[4] ;
 wire \dtop.field_top.controller.ppos[5] ;
 wire \dtop.field_top.controller.ppos[6] ;
 wire \dtop.field_top.controller.timer[0] ;
 wire \dtop.field_top.controller.timer[1] ;
 wire \dtop.field_top.controller.timer[2] ;
 wire \dtop.field_top.fx[0] ;
 wire \dtop.field_top.fx[10] ;
 wire \dtop.field_top.fx[1] ;
 wire \dtop.field_top.fx[2] ;
 wire \dtop.field_top.fx[3] ;
 wire \dtop.field_top.fx[4] ;
 wire \dtop.field_top.fx[5] ;
 wire \dtop.field_top.fx[6] ;
 wire \dtop.field_top.fx[7] ;
 wire \dtop.field_top.fx[8] ;
 wire \dtop.field_top.fx[9] ;
 wire \dtop.field_top.fy[0] ;
 wire \dtop.field_top.fy[10] ;
 wire \dtop.field_top.fy[1] ;
 wire \dtop.field_top.fy[2] ;
 wire \dtop.field_top.fy[3] ;
 wire \dtop.field_top.fy[4] ;
 wire \dtop.field_top.fy[5] ;
 wire \dtop.field_top.fy[6] ;
 wire \dtop.field_top.fy[7] ;
 wire \dtop.field_top.fy[8] ;
 wire \dtop.field_top.fy[9] ;
 wire \dtop.field_top.hsync ;
 wire \dtop.field_top.last_wave[0] ;
 wire \dtop.field_top.last_wave[1] ;
 wire \dtop.field_top.last_wave[2] ;
 wire \dtop.field_top.last_wave[3] ;
 wire \dtop.field_top.last_wave[4] ;
 wire \dtop.field_top.last_wave[5] ;
 wire \dtop.field_top.last_wave[6] ;
 wire \dtop.field_top.last_wave[7] ;
 wire \dtop.field_top.logo_prev_pixel ;
 wire \dtop.field_top.lside ;
 wire \dtop.field_top.masked_bits[0] ;
 wire \dtop.field_top.masked_bits[1] ;
 wire \dtop.field_top.nsource.num_iter[0] ;
 wire \dtop.field_top.nsource.num_iter[1] ;
 wire \dtop.field_top.nsource.shuffle_state.in[0] ;
 wire \dtop.field_top.nsource.shuffle_state.in[1] ;
 wire \dtop.field_top.nsource.shuffle_state.in[2] ;
 wire \dtop.field_top.nsource.shuffle_state.in[3] ;
 wire \dtop.field_top.nsource.shuffle_state.in[4] ;
 wire \dtop.field_top.nsource.shuffle_state.in[5] ;
 wire \dtop.field_top.nsource.shuffle_state.in[6] ;
 wire \dtop.field_top.nsource.shuffle_state.in[7] ;
 wire \dtop.field_top.player.chan_timer[0] ;
 wire \dtop.field_top.player.chan_timer[1] ;
 wire \dtop.field_top.player.chan_timer[2] ;
 wire \dtop.field_top.player.chan_timer[3] ;
 wire \dtop.field_top.player.chan_timer[4] ;
 wire \dtop.field_top.player.chan_timer[5] ;
 wire \dtop.field_top.player.controller.pattern0[0] ;
 wire \dtop.field_top.player.controller.pattern0[1] ;
 wire \dtop.field_top.player.controller.pattern0[2] ;
 wire \dtop.field_top.player.controller.ppos[0] ;
 wire \dtop.field_top.player.controller.ppos[1] ;
 wire \dtop.field_top.player.controller.ppos[2] ;
 wire \dtop.field_top.player.controller.ppos[3] ;
 wire \dtop.field_top.player.controller.ppos[4] ;
 wire \dtop.field_top.player.controller.ppos[5] ;
 wire \dtop.field_top.player.controller.ppos[6] ;
 wire \dtop.field_top.player.controller.timer[0] ;
 wire \dtop.field_top.player.controller.timer[1] ;
 wire \dtop.field_top.player.controller.timer[2] ;
 wire \dtop.field_top.player.osc0[0] ;
 wire \dtop.field_top.player.osc0[10] ;
 wire \dtop.field_top.player.osc0[11] ;
 wire \dtop.field_top.player.osc0[12] ;
 wire \dtop.field_top.player.osc0[13] ;
 wire \dtop.field_top.player.osc0[14] ;
 wire \dtop.field_top.player.osc0[15] ;
 wire \dtop.field_top.player.osc0[16] ;
 wire \dtop.field_top.player.osc0[17] ;
 wire \dtop.field_top.player.osc0[18] ;
 wire \dtop.field_top.player.osc0[19] ;
 wire \dtop.field_top.player.osc0[1] ;
 wire \dtop.field_top.player.osc0[20] ;
 wire \dtop.field_top.player.osc0[21] ;
 wire \dtop.field_top.player.osc0[22] ;
 wire \dtop.field_top.player.osc0[2] ;
 wire \dtop.field_top.player.osc0[3] ;
 wire \dtop.field_top.player.osc0[4] ;
 wire \dtop.field_top.player.osc0[5] ;
 wire \dtop.field_top.player.osc0[6] ;
 wire \dtop.field_top.player.osc0[7] ;
 wire \dtop.field_top.player.osc0[8] ;
 wire \dtop.field_top.player.osc0[9] ;
 wire \dtop.field_top.player.out_acc[0] ;
 wire \dtop.field_top.player.out_acc[1] ;
 wire \dtop.field_top.player.out_acc[2] ;
 wire \dtop.field_top.player.out_acc[3] ;
 wire \dtop.field_top.player.out_acc[4] ;
 wire \dtop.field_top.player.out_acc[5] ;
 wire \dtop.field_top.player.out_acc[6] ;
 wire \dtop.field_top.player.out_acc[7] ;
 wire \dtop.field_top.player.out_acc[8] ;
 wire \dtop.field_top.player.out_acc[9] ;
 wire \dtop.field_top.player.out_pw[0] ;
 wire \dtop.field_top.player.out_pw[1] ;
 wire \dtop.field_top.player.out_pw[2] ;
 wire \dtop.field_top.player.out_pw[3] ;
 wire \dtop.field_top.player.out_pw[4] ;
 wire \dtop.field_top.player.out_pw[5] ;
 wire \dtop.field_top.player.out_pw[6] ;
 wire \dtop.field_top.player.out_pw[7] ;
 wire \dtop.field_top.player.out_pw[8] ;
 wire \dtop.field_top.player.out_pw[9] ;
 wire \dtop.field_top.player.out_pw_high ;
 wire \dtop.field_top.player.sched.alu.p0 ;
 wire \dtop.field_top.player.sched.alu.p1 ;
 wire \dtop.field_top.prev_wave[0] ;
 wire \dtop.field_top.prev_wave[1] ;
 wire \dtop.field_top.prev_wave[2] ;
 wire \dtop.field_top.prev_wave[3] ;
 wire \dtop.field_top.prev_wave[4] ;
 wire \dtop.field_top.prev_wave[5] ;
 wire \dtop.field_top.prev_wave[6] ;
 wire \dtop.field_top.prev_wave[7] ;
 wire \dtop.field_top.reg1[11] ;
 wire \dtop.field_top.reg1[12] ;
 wire \dtop.field_top.reg1[13] ;
 wire \dtop.field_top.reg1[14] ;
 wire \dtop.field_top.reg1[15] ;
 wire \dtop.field_top.reg1[16] ;
 wire \dtop.field_top.reg2[11] ;
 wire \dtop.field_top.reg2[12] ;
 wire \dtop.field_top.reg2[13] ;
 wire \dtop.field_top.reg2[14] ;
 wire \dtop.field_top.reg2[15] ;
 wire \dtop.field_top.reg2[16] ;
 wire \dtop.field_top.reg3[11] ;
 wire \dtop.field_top.reg3[12] ;
 wire \dtop.field_top.reg3[13] ;
 wire \dtop.field_top.reg3[14] ;
 wire \dtop.field_top.reg3[15] ;
 wire \dtop.field_top.reg3[16] ;
 wire \dtop.field_top.reg4[11] ;
 wire \dtop.field_top.reg4[12] ;
 wire \dtop.field_top.reg4[13] ;
 wire \dtop.field_top.reg4[14] ;
 wire \dtop.field_top.reg4[15] ;
 wire \dtop.field_top.reg4[16] ;
 wire \dtop.field_top.rs.scan_x.state[0] ;
 wire \dtop.field_top.rs.scan_x.state[1] ;
 wire \dtop.field_top.rs.scan_y.pos[8] ;
 wire \dtop.field_top.rs.scan_y.pos[9] ;
 wire \dtop.field_top.rs.scan_y.state[0] ;
 wire \dtop.field_top.rs.scan_y.state[1] ;
 wire \dtop.field_top.rs.vsync ;
 wire \dtop.field_top.rside ;
 wire \dtop.field_top.sflag ;
 wire \dtop.field_top.sflag2 ;
 wire \dtop.field_top.wave[0] ;
 wire \dtop.field_top.wave[1] ;
 wire \dtop.field_top.wave[2] ;
 wire \dtop.field_top.wave[3] ;
 wire \dtop.field_top.wave[4] ;
 wire \dtop.field_top.wave[5] ;
 wire \dtop.field_top.wave[6] ;
 wire \dtop.field_top.wave[7] ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_leaf_0_clk;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;

 sg13g2_inv_1 _3559_ (.Y(_2821_),
    .A(net657));
 sg13g2_inv_1 _3560_ (.Y(_2822_),
    .A(\dtop.field_top.channel_output[0] ));
 sg13g2_inv_1 _3561_ (.Y(_2823_),
    .A(\dtop.field_top.player.osc0[10] ));
 sg13g2_inv_1 _3562_ (.Y(_2824_),
    .A(\dtop.field_top.player.osc0[9] ));
 sg13g2_inv_1 _3563_ (.Y(_2825_),
    .A(net428));
 sg13g2_inv_1 _3564_ (.Y(_2826_),
    .A(net374));
 sg13g2_inv_1 _3565_ (.Y(_2827_),
    .A(net526));
 sg13g2_inv_1 _3566_ (.Y(_2828_),
    .A(net575));
 sg13g2_inv_1 _3567_ (.Y(_2829_),
    .A(net610));
 sg13g2_inv_2 _3568_ (.Y(_2830_),
    .A(net1029));
 sg13g2_inv_1 _3569_ (.Y(_2831_),
    .A(net1062));
 sg13g2_inv_2 _3570_ (.Y(_2832_),
    .A(net1066));
 sg13g2_inv_1 _3571_ (.Y(_2833_),
    .A(net1071));
 sg13g2_inv_2 _3572_ (.Y(_2834_),
    .A(net1082));
 sg13g2_inv_4 _3573_ (.A(net1088),
    .Y(_2835_));
 sg13g2_inv_4 _3574_ (.A(net1090),
    .Y(_2836_));
 sg13g2_inv_1 _3575_ (.Y(_2837_),
    .A(net1093));
 sg13g2_inv_1 _3576_ (.Y(_2838_),
    .A(\dtop.field_top.fy[10] ));
 sg13g2_inv_2 _3577_ (.Y(_2839_),
    .A(net1108));
 sg13g2_inv_1 _3578_ (.Y(_2840_),
    .A(\dtop.field_top.fy[5] ));
 sg13g2_inv_1 _3579_ (.Y(_2841_),
    .A(\dtop.field_top.fx[4] ));
 sg13g2_inv_1 _3580_ (.Y(_2842_),
    .A(net1119));
 sg13g2_inv_2 _3581_ (.Y(_2843_),
    .A(net1036));
 sg13g2_inv_1 _3582_ (.Y(_2844_),
    .A(net1041));
 sg13g2_inv_1 _3583_ (.Y(_2845_),
    .A(net1037));
 sg13g2_inv_4 _3584_ (.A(net1046),
    .Y(_2846_));
 sg13g2_inv_2 _3585_ (.Y(_2847_),
    .A(net1048));
 sg13g2_inv_1 _3586_ (.Y(_2848_),
    .A(net1044));
 sg13g2_inv_1 _3587_ (.Y(_2849_),
    .A(net1030));
 sg13g2_inv_1 _3588_ (.Y(_2850_),
    .A(net1031));
 sg13g2_inv_1 _3589_ (.Y(_2851_),
    .A(\dtop.field_top.player.controller.pattern0[2] ));
 sg13g2_inv_2 _3590_ (.Y(_2852_),
    .A(net1070));
 sg13g2_inv_2 _3591_ (.Y(_2853_),
    .A(\dtop.field_top.player.controller.ppos[5] ));
 sg13g2_inv_2 _3592_ (.Y(_2854_),
    .A(\dtop.field_top.player.controller.ppos[6] ));
 sg13g2_inv_2 _3593_ (.Y(_2855_),
    .A(\dtop.field_top.player.controller.ppos[2] ));
 sg13g2_inv_2 _3594_ (.Y(_2856_),
    .A(net1103));
 sg13g2_inv_1 _3595_ (.Y(_2857_),
    .A(net1027));
 sg13g2_inv_1 _3596_ (.Y(_2858_),
    .A(net1106));
 sg13g2_inv_1 _3597_ (.Y(_2859_),
    .A(_0115_));
 sg13g2_inv_2 _3598_ (.Y(_2860_),
    .A(net663));
 sg13g2_inv_1 _3599_ (.Y(_2861_),
    .A(\dtop.field_top.afl_sub_pc[1] ));
 sg13g2_inv_2 _3600_ (.Y(_2862_),
    .A(net1056));
 sg13g2_inv_1 _3601_ (.Y(_2863_),
    .A(net1053));
 sg13g2_inv_1 _3602_ (.Y(_2864_),
    .A(net1050));
 sg13g2_inv_1 _3603_ (.Y(_2865_),
    .A(net602));
 sg13g2_inv_1 _3604_ (.Y(_2866_),
    .A(net712));
 sg13g2_inv_1 _3605_ (.Y(_2867_),
    .A(\dtop.field_top.alt_osc[6] ));
 sg13g2_inv_1 _3606_ (.Y(_2868_),
    .A(\dtop.field_top.alt_osc[8] ));
 sg13g2_inv_2 _3607_ (.Y(_2869_),
    .A(_0017_));
 sg13g2_inv_1 _3608_ (.Y(_2870_),
    .A(_0401_));
 sg13g2_inv_1 _3609_ (.Y(_2871_),
    .A(_0020_));
 sg13g2_inv_1 _3610_ (.Y(_2872_),
    .A(net507));
 sg13g2_inv_1 _3611_ (.Y(_2873_),
    .A(\dtop.field_top.comp_values0[3][9] ));
 sg13g2_inv_1 _3612_ (.Y(_2874_),
    .A(_0027_));
 sg13g2_inv_2 _3613_ (.Y(_2875_),
    .A(net708));
 sg13g2_inv_1 _3614_ (.Y(_2876_),
    .A(_0029_));
 sg13g2_inv_4 _3615_ (.A(net673),
    .Y(_2877_));
 sg13g2_inv_2 _3616_ (.Y(_2878_),
    .A(net711));
 sg13g2_inv_1 _3617_ (.Y(_2879_),
    .A(_0035_));
 sg13g2_inv_1 _3618_ (.Y(_2880_),
    .A(_0034_));
 sg13g2_inv_2 _3619_ (.Y(_2881_),
    .A(net651));
 sg13g2_inv_1 _3620_ (.Y(_2882_),
    .A(_0043_));
 sg13g2_inv_1 _3621_ (.Y(_2883_),
    .A(_0045_));
 sg13g2_inv_1 _3622_ (.Y(_2884_),
    .A(\dtop.field_top.comp_value0_1[2] ));
 sg13g2_inv_1 _3623_ (.Y(_2885_),
    .A(net524));
 sg13g2_inv_1 _3624_ (.Y(_2886_),
    .A(\dtop.field_top.comp_values0[3][2] ));
 sg13g2_inv_1 _3625_ (.Y(_2887_),
    .A(_0049_));
 sg13g2_inv_1 _3626_ (.Y(_2888_),
    .A(net459));
 sg13g2_inv_1 _3627_ (.Y(_2889_),
    .A(net567));
 sg13g2_inv_1 _3628_ (.Y(_2890_),
    .A(net530));
 sg13g2_inv_1 _3629_ (.Y(_2891_),
    .A(\dtop.field_top.comp_values0[2][3] ));
 sg13g2_inv_1 _3630_ (.Y(_2892_),
    .A(_0050_));
 sg13g2_inv_1 _3631_ (.Y(_2893_),
    .A(\dtop.field_top.comp_value0_1[4] ));
 sg13g2_inv_1 _3632_ (.Y(_2894_),
    .A(\dtop.field_top.comp_values0[3][4] ));
 sg13g2_inv_1 _3633_ (.Y(_2895_),
    .A(net551));
 sg13g2_inv_1 _3634_ (.Y(_2896_),
    .A(_0051_));
 sg13g2_inv_1 _3635_ (.Y(_2897_),
    .A(\dtop.field_top.comp_values0[3][10] ));
 sg13g2_inv_1 _3636_ (.Y(_2898_),
    .A(net426));
 sg13g2_inv_1 _3637_ (.Y(_2899_),
    .A(net589));
 sg13g2_inv_1 _3638_ (.Y(_2900_),
    .A(net539));
 sg13g2_inv_1 _3639_ (.Y(_2901_),
    .A(\dtop.field_top.comp_values0[2][5] ));
 sg13g2_inv_1 _3640_ (.Y(_2902_),
    .A(_0057_));
 sg13g2_inv_1 _3641_ (.Y(_2903_),
    .A(net473));
 sg13g2_inv_1 _3642_ (.Y(_2904_),
    .A(\dtop.field_top.comp_values0[4][6] ));
 sg13g2_inv_1 _3643_ (.Y(_2905_),
    .A(net501));
 sg13g2_inv_1 _3644_ (.Y(_2906_),
    .A(net597));
 sg13g2_inv_1 _3645_ (.Y(_2907_),
    .A(_0058_));
 sg13g2_inv_1 _3646_ (.Y(_2908_),
    .A(net436));
 sg13g2_inv_1 _3647_ (.Y(_2909_),
    .A(net493));
 sg13g2_inv_1 _3648_ (.Y(_2910_),
    .A(_0059_));
 sg13g2_inv_1 _3649_ (.Y(_2911_),
    .A(_0060_));
 sg13g2_inv_1 _3650_ (.Y(_2912_),
    .A(\dtop.field_top.player.out_pw[5] ));
 sg13g2_inv_1 _3651_ (.Y(_2913_),
    .A(_0063_));
 sg13g2_inv_1 _3652_ (.Y(_2914_),
    .A(net333));
 sg13g2_inv_1 _3653_ (.Y(_2915_),
    .A(net375));
 sg13g2_inv_1 _3654_ (.Y(_2916_),
    .A(\dtop.field_top.wave[5] ));
 sg13g2_inv_1 _3655_ (.Y(_2917_),
    .A(net342));
 sg13g2_inv_1 _3656_ (.Y(_2918_),
    .A(\dtop.field_top.last_wave[0] ));
 sg13g2_inv_1 _3657_ (.Y(_2919_),
    .A(\dtop.field_top.last_wave[1] ));
 sg13g2_inv_1 _3658_ (.Y(_2920_),
    .A(\dtop.field_top.last_wave[4] ));
 sg13g2_inv_1 _3659_ (.Y(_2921_),
    .A(net396));
 sg13g2_inv_1 _3660_ (.Y(_2922_),
    .A(net405));
 sg13g2_inv_1 _3661_ (.Y(_2923_),
    .A(net441));
 sg13g2_inv_1 _3662_ (.Y(_2924_),
    .A(\dtop.field_top.comp_value0[1] ));
 sg13g2_inv_2 _3663_ (.Y(_2925_),
    .A(net587));
 sg13g2_inv_2 _3664_ (.Y(_2926_),
    .A(\dtop.field_top.player.controller.timer[2] ));
 sg13g2_inv_2 _3665_ (.Y(_2927_),
    .A(\dtop.field_top.player.controller.timer[1] ));
 sg13g2_inv_2 _3666_ (.Y(_2928_),
    .A(\dtop.field_top.player.controller.timer[0] ));
 sg13g2_nand2_2 _3667_ (.Y(\dtop.field_top.hsync ),
    .A(_2865_),
    .B(net692));
 sg13g2_nand2_2 _3668_ (.Y(\dtop.field_top.rs.vsync ),
    .A(net699),
    .B(net639));
 sg13g2_nand2_2 _3669_ (.Y(_2929_),
    .A(net602),
    .B(\dtop.field_top.rs.scan_x.state[0] ));
 sg13g2_nand3_1 _3670_ (.B(\dtop.field_top.rs.scan_x.state[1] ),
    .C(\dtop.field_top.rs.scan_x.state[0] ),
    .A(_0107_),
    .Y(_2930_));
 sg13g2_and2_1 _3671_ (.A(net1038),
    .B(_2930_),
    .X(_2931_));
 sg13g2_o21ai_1 _3672_ (.B1(_0009_),
    .Y(_2932_),
    .A1(net1018),
    .A2(\dtop.field_top.hsync ));
 sg13g2_nor2_1 _3673_ (.A(net1048),
    .B(_2865_),
    .Y(_2933_));
 sg13g2_nand2_1 _3674_ (.Y(_2934_),
    .A(net1016),
    .B(\dtop.field_top.rs.scan_x.state[1] ));
 sg13g2_nand3_1 _3675_ (.B(_2932_),
    .C(_2934_),
    .A(net1014),
    .Y(_2935_));
 sg13g2_o21ai_1 _3676_ (.B1(net1041),
    .Y(_2936_),
    .A1(net1016),
    .A2(\dtop.field_top.rs.scan_x.state[0] ));
 sg13g2_a21oi_1 _3677_ (.A1(\dtop.field_top.hsync ),
    .A2(_2936_),
    .Y(_2937_),
    .B1(_0009_));
 sg13g2_nand2_1 _3678_ (.Y(_2938_),
    .A(net1040),
    .B(\dtop.field_top.rs.scan_x.state[1] ));
 sg13g2_a221oi_1 _3679_ (.B2(net1047),
    .C1(net1034),
    .B1(_2938_),
    .A1(\dtop.field_top.rs.scan_x.state[1] ),
    .Y(_2939_),
    .A2(\dtop.field_top.rs.scan_x.state[0] ));
 sg13g2_nor2_1 _3680_ (.A(net1038),
    .B(_2939_),
    .Y(_2940_));
 sg13g2_nand2_1 _3681_ (.Y(_2941_),
    .A(net1058),
    .B(net686));
 sg13g2_nand2_2 _3682_ (.Y(_2942_),
    .A(net1056),
    .B(net1052));
 sg13g2_nand4_1 _3683_ (.B(\dtop.field_top.afl_sub_pc[1] ),
    .C(net1056),
    .A(net1058),
    .Y(_2943_),
    .D(net1053));
 sg13g2_nor2_2 _3684_ (.A(net648),
    .B(_2943_),
    .Y(_2944_));
 sg13g2_o21ai_1 _3685_ (.B1(_2944_),
    .Y(_2945_),
    .A1(net1037),
    .A2(_2939_));
 sg13g2_nor4_2 _3686_ (.A(_2931_),
    .B(_2935_),
    .C(_2937_),
    .Y(_2946_),
    .D(_2945_));
 sg13g2_nor2b_2 _3687_ (.A(\dtop.field_top.hsync ),
    .B_N(_2946_),
    .Y(_2947_));
 sg13g2_nand2b_2 _3688_ (.Y(_2948_),
    .B(_2946_),
    .A_N(\dtop.field_top.hsync ));
 sg13g2_nand3_1 _3689_ (.B(_0016_),
    .C(\dtop.field_top.rs.scan_y.pos[9] ),
    .A(_0015_),
    .Y(_2949_));
 sg13g2_or2_1 _3690_ (.X(_2950_),
    .B(_0011_),
    .A(\dtop.field_top.rs.scan_y.state[0] ));
 sg13g2_nand2_1 _3691_ (.Y(_2951_),
    .A(\dtop.field_top.rs.scan_y.pos[8] ),
    .B(_0014_));
 sg13g2_nor3_1 _3692_ (.A(_2949_),
    .B(_2950_),
    .C(_2951_),
    .Y(_2952_));
 sg13g2_nor2_1 _3693_ (.A(\dtop.field_top.rs.scan_y.pos[8] ),
    .B(_0016_),
    .Y(_2953_));
 sg13g2_nand2_1 _3694_ (.Y(_2954_),
    .A(_2950_),
    .B(_2953_));
 sg13g2_nor4_1 _3695_ (.A(_0014_),
    .B(_0015_),
    .C(net601),
    .D(_2954_),
    .Y(_2955_));
 sg13g2_nand2b_1 _3696_ (.Y(_2956_),
    .B(\dtop.field_top.rs.scan_y.state[1] ),
    .A_N(\dtop.field_top.rs.scan_y.state[0] ));
 sg13g2_nor2_1 _3697_ (.A(_0013_),
    .B(\dtop.field_top.alt_osc[5] ),
    .Y(_2957_));
 sg13g2_nor2_1 _3698_ (.A(_0010_),
    .B(_0012_),
    .Y(_2958_));
 sg13g2_o21ai_1 _3699_ (.B1(_2958_),
    .Y(_2959_),
    .A1(\dtop.field_top.rs.scan_y.state[1] ),
    .A2(_2957_));
 sg13g2_nand3_1 _3700_ (.B(\dtop.field_top.alt_osc[5] ),
    .C(_2950_),
    .A(_0013_),
    .Y(_2960_));
 sg13g2_a221oi_1 _3701_ (.B2(\dtop.field_top.rs.scan_y.state[1] ),
    .C1(_2959_),
    .B1(_2960_),
    .A1(_0011_),
    .Y(_2961_),
    .A2(_2956_));
 sg13g2_o21ai_1 _3702_ (.B1(_2961_),
    .Y(_2962_),
    .A1(_2952_),
    .A2(_2955_));
 sg13g2_nor2_1 _3703_ (.A(_2948_),
    .B(_2962_),
    .Y(_2963_));
 sg13g2_nand2b_1 _3704_ (.Y(_2964_),
    .B(_2963_),
    .A_N(\dtop.field_top.rs.vsync ));
 sg13g2_nor2_1 _3705_ (.A(_2937_),
    .B(_2940_),
    .Y(_2965_));
 sg13g2_nand4_1 _3706_ (.B(_2934_),
    .C(_2944_),
    .A(_2932_),
    .Y(_2966_),
    .D(_2965_));
 sg13g2_nor3_2 _3707_ (.A(net1043),
    .B(_2931_),
    .C(_2966_),
    .Y(_2967_));
 sg13g2_nand2_1 _3708_ (.Y(_2968_),
    .A(_2932_),
    .B(_2944_));
 sg13g2_nor4_1 _3709_ (.A(net1043),
    .B(_2931_),
    .C(_2933_),
    .D(_2968_),
    .Y(_2969_));
 sg13g2_and4_1 _3710_ (.A(_2865_),
    .B(\dtop.field_top.rs.scan_x.state[0] ),
    .C(_2965_),
    .D(_2969_),
    .X(_2970_));
 sg13g2_inv_2 _3711_ (.Y(_2971_),
    .A(net958));
 sg13g2_and2_1 _3712_ (.A(net1116),
    .B(_2964_),
    .X(_2972_));
 sg13g2_nand2_2 _3713_ (.Y(_2973_),
    .A(net1116),
    .B(_2964_));
 sg13g2_nand2_1 _3714_ (.Y(_2974_),
    .A(net665),
    .B(net933));
 sg13g2_o21ai_1 _3715_ (.B1(_2974_),
    .Y(_2975_),
    .A1(net1020),
    .A2(net933));
 sg13g2_inv_2 _3716_ (.Y(_0001_),
    .A(_2975_));
 sg13g2_nand2_1 _3717_ (.Y(_2976_),
    .A(\dtop.field_top.player.out_pw[7] ),
    .B(\dtop.field_top.player.out_pw[8] ));
 sg13g2_nor3_1 _3718_ (.A(\dtop.field_top.player.out_pw[6] ),
    .B(\dtop.field_top.player.out_pw[9] ),
    .C(_2976_),
    .Y(_2977_));
 sg13g2_nand2_1 _3719_ (.Y(_2978_),
    .A(\dtop.field_top.player.out_pw[3] ),
    .B(\dtop.field_top.player.out_pw[2] ));
 sg13g2_nor3_1 _3720_ (.A(\dtop.field_top.player.out_pw[5] ),
    .B(\dtop.field_top.player.out_pw[4] ),
    .C(_2978_),
    .Y(_2979_));
 sg13g2_nand4_1 _3721_ (.B(net384),
    .C(_2977_),
    .A(\dtop.field_top.player.out_pw[1] ),
    .Y(_2980_),
    .D(_2979_));
 sg13g2_inv_1 _3722_ (.Y(\dtop.field_top.player.out_pw_high ),
    .A(net385));
 sg13g2_nand2_1 _3723_ (.Y(_2981_),
    .A(net660),
    .B(net932));
 sg13g2_o21ai_1 _3724_ (.B1(_2981_),
    .Y(_2982_),
    .A1(_2834_),
    .A2(net932));
 sg13g2_nand2_1 _3725_ (.Y(_2983_),
    .A(net353),
    .B(net932));
 sg13g2_o21ai_1 _3726_ (.B1(_2983_),
    .Y(_2984_),
    .A1(_2835_),
    .A2(net932));
 sg13g2_nor2_2 _3727_ (.A(_2982_),
    .B(_2984_),
    .Y(_0163_));
 sg13g2_nor2_1 _3728_ (.A(_0001_),
    .B(_0163_),
    .Y(_2985_));
 sg13g2_nand2_1 _3729_ (.Y(_2986_),
    .A(net322),
    .B(net933));
 sg13g2_o21ai_1 _3730_ (.B1(_2986_),
    .Y(_2987_),
    .A1(_2836_),
    .A2(net932));
 sg13g2_o21ai_1 _3731_ (.B1(_2985_),
    .Y(_0285_),
    .A1(_2982_),
    .A2(_2987_));
 sg13g2_and2_1 _3732_ (.A(_2982_),
    .B(_2984_),
    .X(_2988_));
 sg13g2_inv_1 _3733_ (.Y(_0162_),
    .A(_2988_));
 sg13g2_o21ai_1 _3734_ (.B1(_2982_),
    .Y(_2989_),
    .A1(_2984_),
    .A2(_2987_));
 sg13g2_and2_1 _3735_ (.A(_0285_),
    .B(_2989_),
    .X(_0000_));
 sg13g2_a21oi_1 _3736_ (.A1(_0001_),
    .A2(_2988_),
    .Y(_0002_),
    .B1(_0163_));
 sg13g2_xnor2_1 _3737_ (.Y(_0003_),
    .A(_0001_),
    .B(_0163_));
 sg13g2_or2_1 _3738_ (.X(_2990_),
    .B(_2963_),
    .A(net699));
 sg13g2_nand2_1 _3739_ (.Y(_2991_),
    .A(net699),
    .B(_2963_));
 sg13g2_and3_1 _3740_ (.X(_0118_),
    .A(net1116),
    .B(_2990_),
    .C(_2991_));
 sg13g2_nand3_1 _3741_ (.B(net639),
    .C(_2991_),
    .A(net1116),
    .Y(_2992_));
 sg13g2_nor2b_2 _3742_ (.A(\dtop.field_top.rs.scan_y.state[1] ),
    .B_N(\dtop.field_top.rs.scan_y.state[0] ),
    .Y(_2993_));
 sg13g2_nand3_1 _3743_ (.B(net935),
    .C(_2993_),
    .A(_2947_),
    .Y(_2994_));
 sg13g2_o21ai_1 _3744_ (.B1(net640),
    .Y(_0119_),
    .A1(_2962_),
    .A2(net914));
 sg13g2_nor2_2 _3745_ (.A(net1107),
    .B(_2858_),
    .Y(_2995_));
 sg13g2_nand2_2 _3746_ (.Y(_2996_),
    .A(_2839_),
    .B(net1105));
 sg13g2_nor2_1 _3747_ (.A(\dtop.field_top.channel[1] ),
    .B(\dtop.field_top.channel[0] ),
    .Y(_2997_));
 sg13g2_nand3_1 _3748_ (.B(\dtop.field_top.channel[3] ),
    .C(_2997_),
    .A(\dtop.field_top.channel[2] ),
    .Y(_2998_));
 sg13g2_nand2_1 _3749_ (.Y(_2999_),
    .A(net1103),
    .B(net1100));
 sg13g2_nor2b_1 _3750_ (.A(net1026),
    .B_N(net1096),
    .Y(_3000_));
 sg13g2_nand3_1 _3751_ (.B(net1101),
    .C(net1098),
    .A(net1103),
    .Y(_3001_));
 sg13g2_nor3_2 _3752_ (.A(net1027),
    .B(_2998_),
    .C(_3001_),
    .Y(_3002_));
 sg13g2_inv_1 _3753_ (.Y(_3003_),
    .A(_3002_));
 sg13g2_nand2_2 _3754_ (.Y(_3004_),
    .A(_2995_),
    .B(_3002_));
 sg13g2_a21oi_2 _3755_ (.B1(net1115),
    .Y(_3005_),
    .A2(_3002_),
    .A1(_2995_));
 sg13g2_nand2_1 _3756_ (.Y(_3006_),
    .A(net1117),
    .B(_3004_));
 sg13g2_nor2_1 _3757_ (.A(_2996_),
    .B(_2999_),
    .Y(_3007_));
 sg13g2_inv_1 _3758_ (.Y(_3008_),
    .A(_3007_));
 sg13g2_nand3_1 _3759_ (.B(net1025),
    .C(_3007_),
    .A(net1095),
    .Y(_3009_));
 sg13g2_inv_2 _3760_ (.Y(_3010_),
    .A(_3009_));
 sg13g2_nand2_1 _3761_ (.Y(_3011_),
    .A(net1109),
    .B(\dtop.field_top.channel[0] ));
 sg13g2_nor2_1 _3762_ (.A(_3009_),
    .B(_3011_),
    .Y(_3012_));
 sg13g2_a21oi_1 _3763_ (.A1(net633),
    .A2(_3010_),
    .Y(_3013_),
    .B1(net1109));
 sg13g2_nor3_1 _3764_ (.A(_3006_),
    .B(_3012_),
    .C(net634),
    .Y(_0120_));
 sg13g2_xnor2_1 _3765_ (.Y(_3014_),
    .A(net635),
    .B(_3012_));
 sg13g2_nor2_1 _3766_ (.A(_3006_),
    .B(net636),
    .Y(_0121_));
 sg13g2_nand2_1 _3767_ (.Y(_0122_),
    .A(_2860_),
    .B(_3005_));
 sg13g2_nand2_2 _3768_ (.Y(_3015_),
    .A(net1108),
    .B(net1009));
 sg13g2_nand3_1 _3769_ (.B(_2996_),
    .C(_3015_),
    .A(net1117),
    .Y(_0123_));
 sg13g2_nor2_2 _3770_ (.A(_2839_),
    .B(net1009),
    .Y(_3016_));
 sg13g2_nand2_2 _3771_ (.Y(_3017_),
    .A(net1108),
    .B(net1105));
 sg13g2_nand2_1 _3772_ (.Y(_3018_),
    .A(net1103),
    .B(net1105));
 sg13g2_nor2_2 _3773_ (.A(_2856_),
    .B(_3017_),
    .Y(_3019_));
 sg13g2_nand2_1 _3774_ (.Y(_3020_),
    .A(net1104),
    .B(_3016_));
 sg13g2_nor2_1 _3775_ (.A(net1103),
    .B(_3016_),
    .Y(_3021_));
 sg13g2_o21ai_1 _3776_ (.B1(_3005_),
    .Y(_0124_),
    .A1(_3019_),
    .A2(_3021_));
 sg13g2_nor2_2 _3777_ (.A(_0115_),
    .B(_3017_),
    .Y(_3022_));
 sg13g2_xnor2_1 _3778_ (.Y(_3023_),
    .A(net1102),
    .B(_3022_));
 sg13g2_nand2_1 _3779_ (.Y(_0125_),
    .A(_3005_),
    .B(_3023_));
 sg13g2_nor2_1 _3780_ (.A(_3001_),
    .B(_3017_),
    .Y(_3024_));
 sg13g2_a21oi_1 _3781_ (.A1(net1102),
    .A2(_3019_),
    .Y(_3025_),
    .B1(net1098));
 sg13g2_o21ai_1 _3782_ (.B1(_3005_),
    .Y(_0126_),
    .A1(_3024_),
    .A2(net670));
 sg13g2_nand2b_1 _3783_ (.Y(_3026_),
    .B(net1045),
    .A_N(net1039));
 sg13g2_nand2b_2 _3784_ (.Y(_3027_),
    .B(net1055),
    .A_N(net1053));
 sg13g2_or2_2 _3785_ (.X(_3028_),
    .B(net1050),
    .A(net1047));
 sg13g2_nor2_2 _3786_ (.A(_3027_),
    .B(_3028_),
    .Y(_3029_));
 sg13g2_nor4_1 _3787_ (.A(net1040),
    .B(net1034),
    .C(_3027_),
    .D(_3028_),
    .Y(_3030_));
 sg13g2_nand4_1 _3788_ (.B(net1046),
    .C(net1014),
    .A(_2845_),
    .Y(_3031_),
    .D(_3030_));
 sg13g2_nand2b_2 _3789_ (.Y(_3032_),
    .B(net1047),
    .A_N(net1051));
 sg13g2_nor2_2 _3790_ (.A(_3027_),
    .B(_3032_),
    .Y(_3033_));
 sg13g2_nand2b_2 _3791_ (.Y(_3034_),
    .B(net1036),
    .A_N(net1040));
 sg13g2_nor3_1 _3792_ (.A(net1043),
    .B(_3026_),
    .C(_3034_),
    .Y(_3035_));
 sg13g2_nand2_2 _3793_ (.Y(_3036_),
    .A(_3033_),
    .B(net999));
 sg13g2_nand2_2 _3794_ (.Y(_3037_),
    .A(_3031_),
    .B(_3036_));
 sg13g2_nor3_2 _3795_ (.A(net1055),
    .B(net1052),
    .C(_3032_),
    .Y(_3038_));
 sg13g2_nand2b_2 _3796_ (.Y(_3039_),
    .B(net1043),
    .A_N(net1046));
 sg13g2_nor3_1 _3797_ (.A(net1037),
    .B(_3034_),
    .C(_3039_),
    .Y(_3040_));
 sg13g2_nand2b_2 _3798_ (.Y(_3041_),
    .B(net1052),
    .A_N(net1055));
 sg13g2_nor2_2 _3799_ (.A(_3032_),
    .B(_3041_),
    .Y(_3042_));
 sg13g2_nand2_1 _3800_ (.Y(_3043_),
    .A(net994),
    .B(_3042_));
 sg13g2_nand2_2 _3801_ (.Y(_3044_),
    .A(net1047),
    .B(net1051));
 sg13g2_nor3_2 _3802_ (.A(net1055),
    .B(net1052),
    .C(_3044_),
    .Y(_3045_));
 sg13g2_nand2_2 _3803_ (.Y(_3046_),
    .A(net995),
    .B(_3045_));
 sg13g2_nand2_2 _3804_ (.Y(_3047_),
    .A(net714),
    .B(net1043));
 sg13g2_nor3_1 _3805_ (.A(net1037),
    .B(_3034_),
    .C(_3047_),
    .Y(_3048_));
 sg13g2_nand2_1 _3806_ (.Y(_3049_),
    .A(_3033_),
    .B(net992));
 sg13g2_nand2_1 _3807_ (.Y(_3050_),
    .A(_3046_),
    .B(_3049_));
 sg13g2_nor2_2 _3808_ (.A(_3028_),
    .B(_3041_),
    .Y(_3051_));
 sg13g2_nand2_2 _3809_ (.Y(_3052_),
    .A(net998),
    .B(_3051_));
 sg13g2_nor2_2 _3810_ (.A(_2942_),
    .B(_3028_),
    .Y(_3053_));
 sg13g2_nand2_2 _3811_ (.Y(_3054_),
    .A(net995),
    .B(_3053_));
 sg13g2_nand2_1 _3812_ (.Y(_3055_),
    .A(net999),
    .B(_3045_));
 sg13g2_and2_1 _3813_ (.A(_3054_),
    .B(_3055_),
    .X(_3056_));
 sg13g2_nand2_1 _3814_ (.Y(_3057_),
    .A(_3054_),
    .B(_3055_));
 sg13g2_o21ai_1 _3815_ (.B1(net998),
    .Y(_3058_),
    .A1(_3038_),
    .A2(_3051_));
 sg13g2_nand2_1 _3816_ (.Y(_3059_),
    .A(_3043_),
    .B(_3058_));
 sg13g2_nor4_2 _3817_ (.A(_3037_),
    .B(_3050_),
    .C(_3057_),
    .Y(_3060_),
    .D(_3059_));
 sg13g2_nand2_1 _3818_ (.Y(_3061_),
    .A(\dtop.field_top.controller.pattern0[0] ),
    .B(net1031));
 sg13g2_nor2_2 _3819_ (.A(_0108_),
    .B(_3061_),
    .Y(_3062_));
 sg13g2_nor2_1 _3820_ (.A(_2849_),
    .B(\dtop.field_top.controller.pattern0[0] ),
    .Y(_3063_));
 sg13g2_o21ai_1 _3821_ (.B1(_3063_),
    .Y(_3064_),
    .A1(\dtop.field_top.controller.ppos[5] ),
    .A2(_2850_));
 sg13g2_nor2b_1 _3822_ (.A(_3062_),
    .B_N(_3064_),
    .Y(_3065_));
 sg13g2_nand2b_2 _3823_ (.Y(_3066_),
    .B(_3064_),
    .A_N(_3062_));
 sg13g2_nand2b_2 _3824_ (.Y(_3067_),
    .B(net1051),
    .A_N(net1047));
 sg13g2_nor2_2 _3825_ (.A(_2942_),
    .B(_3067_),
    .Y(_3068_));
 sg13g2_and2_1 _3826_ (.A(net993),
    .B(_3068_),
    .X(_3069_));
 sg13g2_nor3_2 _3827_ (.A(net1055),
    .B(net1053),
    .C(_3028_),
    .Y(_3070_));
 sg13g2_nand2_1 _3828_ (.Y(_3071_),
    .A(net996),
    .B(_3070_));
 sg13g2_o21ai_1 _3829_ (.B1(net993),
    .Y(_3072_),
    .A1(_3068_),
    .A2(_3070_));
 sg13g2_nor2_2 _3830_ (.A(_3027_),
    .B(_3044_),
    .Y(_3073_));
 sg13g2_o21ai_1 _3831_ (.B1(net992),
    .Y(_3074_),
    .A1(_3070_),
    .A2(_3073_));
 sg13g2_and3_1 _3832_ (.X(_3075_),
    .A(net969),
    .B(_3072_),
    .C(_3074_));
 sg13g2_nor2_2 _3833_ (.A(_3027_),
    .B(_3067_),
    .Y(_3076_));
 sg13g2_nand2_1 _3834_ (.Y(_3077_),
    .A(net994),
    .B(_3076_));
 sg13g2_nor2_2 _3835_ (.A(_2942_),
    .B(_3032_),
    .Y(_3078_));
 sg13g2_a22oi_1 _3836_ (.Y(_3079_),
    .B1(_3078_),
    .B2(net991),
    .A2(_3076_),
    .A1(net995));
 sg13g2_nand2b_1 _3837_ (.Y(_3080_),
    .B(net1040),
    .A_N(net1037));
 sg13g2_nor4_2 _3838_ (.A(_2843_),
    .B(net1046),
    .C(net1043),
    .Y(_3081_),
    .D(_3080_));
 sg13g2_nor2_1 _3839_ (.A(net1055),
    .B(_3067_),
    .Y(_3082_));
 sg13g2_nor3_2 _3840_ (.A(net1055),
    .B(net1052),
    .C(_3067_),
    .Y(_3083_));
 sg13g2_nand2_1 _3841_ (.Y(_3084_),
    .A(net991),
    .B(_3083_));
 sg13g2_a22oi_1 _3842_ (.Y(_3085_),
    .B1(_3083_),
    .B2(net991),
    .A2(net990),
    .A1(_3029_));
 sg13g2_nor2_2 _3843_ (.A(_3041_),
    .B(_3044_),
    .Y(_3086_));
 sg13g2_nand2_1 _3844_ (.Y(_3087_),
    .A(net993),
    .B(_3086_));
 sg13g2_o21ai_1 _3845_ (.B1(_3086_),
    .Y(_3088_),
    .A1(net998),
    .A2(net994));
 sg13g2_inv_1 _3846_ (.Y(_3089_),
    .A(_3088_));
 sg13g2_a21oi_1 _3847_ (.A1(net999),
    .A2(_3082_),
    .Y(_3090_),
    .B1(_3089_));
 sg13g2_nand4_1 _3848_ (.B(_3079_),
    .C(_3085_),
    .A(_3075_),
    .Y(_3091_),
    .D(_3090_));
 sg13g2_nor2_1 _3849_ (.A(_2942_),
    .B(_3044_),
    .Y(_3092_));
 sg13g2_nand4_1 _3850_ (.B(net1055),
    .C(net1052),
    .A(net1047),
    .Y(_3093_),
    .D(net1050));
 sg13g2_nand2_1 _3851_ (.Y(_3094_),
    .A(net991),
    .B(_3092_));
 sg13g2_nand2_2 _3852_ (.Y(_3095_),
    .A(_3033_),
    .B(net990));
 sg13g2_nand2_1 _3853_ (.Y(_3096_),
    .A(_3068_),
    .B(net990));
 sg13g2_nand3_1 _3854_ (.B(_3095_),
    .C(_3096_),
    .A(_3094_),
    .Y(_3097_));
 sg13g2_a22oi_1 _3855_ (.Y(_3098_),
    .B1(_3078_),
    .B2(net997),
    .A2(_3051_),
    .A1(net994));
 sg13g2_nand2_2 _3856_ (.Y(_3099_),
    .A(_3033_),
    .B(net993));
 sg13g2_nand2_1 _3857_ (.Y(_3100_),
    .A(_3038_),
    .B(net992));
 sg13g2_nand3_1 _3858_ (.B(_3099_),
    .C(_3100_),
    .A(_3098_),
    .Y(_3101_));
 sg13g2_a22oi_1 _3859_ (.Y(_3102_),
    .B1(_3076_),
    .B2(_3081_),
    .A2(_3051_),
    .A1(net992));
 sg13g2_nand2_1 _3860_ (.Y(_3103_),
    .A(net1000),
    .B(_3070_));
 sg13g2_nand2_1 _3861_ (.Y(_3104_),
    .A(_3102_),
    .B(_3103_));
 sg13g2_nor4_2 _3862_ (.A(_3091_),
    .B(_3097_),
    .C(_3101_),
    .Y(_3105_),
    .D(_3104_));
 sg13g2_nand2_2 _3863_ (.Y(_3106_),
    .A(net998),
    .B(_3042_));
 sg13g2_and2_2 _3864_ (.A(net966),
    .B(_3106_),
    .X(_3107_));
 sg13g2_and2_2 _3865_ (.A(_3029_),
    .B(net994),
    .X(_3108_));
 sg13g2_nand2_1 _3866_ (.Y(_3109_),
    .A(_3029_),
    .B(net994));
 sg13g2_nand3_1 _3867_ (.B(_3107_),
    .C(_3109_),
    .A(_3052_),
    .Y(_3110_));
 sg13g2_nor2_1 _3868_ (.A(_3037_),
    .B(_3110_),
    .Y(_3111_));
 sg13g2_nand2_2 _3869_ (.Y(_3112_),
    .A(net993),
    .B(_3073_));
 sg13g2_inv_1 _3870_ (.Y(_3113_),
    .A(_3112_));
 sg13g2_nor2_1 _3871_ (.A(_3069_),
    .B(_3113_),
    .Y(_3114_));
 sg13g2_nand3_1 _3872_ (.B(_3090_),
    .C(_3114_),
    .A(_3056_),
    .Y(_0402_));
 sg13g2_o21ai_1 _3873_ (.B1(net1000),
    .Y(_0403_),
    .A1(_3038_),
    .A2(_3070_));
 sg13g2_inv_1 _3874_ (.Y(_0404_),
    .A(_0403_));
 sg13g2_nand2_1 _3875_ (.Y(_0405_),
    .A(_3071_),
    .B(_3099_));
 sg13g2_nand3_1 _3876_ (.B(net995),
    .C(_3082_),
    .A(net1052),
    .Y(_0406_));
 sg13g2_nand3_1 _3877_ (.B(_0403_),
    .C(_0406_),
    .A(_3046_),
    .Y(_0407_));
 sg13g2_nor3_1 _3878_ (.A(_0402_),
    .B(_0405_),
    .C(_0407_),
    .Y(_0408_));
 sg13g2_a22oi_1 _3879_ (.Y(_0409_),
    .B1(_3111_),
    .B2(_0408_),
    .A2(_3105_),
    .A1(_3060_));
 sg13g2_o21ai_1 _3880_ (.B1(net992),
    .Y(_0410_),
    .A1(_3029_),
    .A2(_3086_));
 sg13g2_nand2_1 _3881_ (.Y(_0411_),
    .A(net998),
    .B(_3076_));
 sg13g2_nand2_1 _3882_ (.Y(_0412_),
    .A(_3045_),
    .B(net991));
 sg13g2_nor4_1 _3883_ (.A(net1037),
    .B(_3034_),
    .C(_3039_),
    .D(_3093_),
    .Y(_0413_));
 sg13g2_o21ai_1 _3884_ (.B1(_3092_),
    .Y(_0414_),
    .A1(net998),
    .A2(net994));
 sg13g2_nand4_1 _3885_ (.B(_0411_),
    .C(_0412_),
    .A(_0406_),
    .Y(_0415_),
    .D(_0414_));
 sg13g2_nor2_2 _3886_ (.A(net967),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_nand2_1 _3887_ (.Y(_0417_),
    .A(_0410_),
    .B(_0416_));
 sg13g2_nand4_1 _3888_ (.B(_2862_),
    .C(net1005),
    .A(net1016),
    .Y(_0418_),
    .D(_3081_));
 sg13g2_o21ai_1 _3889_ (.B1(net991),
    .Y(_0419_),
    .A1(_3053_),
    .A2(_3076_));
 sg13g2_nand2_1 _3890_ (.Y(_0420_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_a21oi_1 _3891_ (.A1(_3032_),
    .A2(_3067_),
    .Y(_0421_),
    .B1(_3041_));
 sg13g2_o21ai_1 _3892_ (.B1(_0421_),
    .Y(_0422_),
    .A1(net991),
    .A2(net990));
 sg13g2_o21ai_1 _3893_ (.B1(net990),
    .Y(_0423_),
    .A1(_3038_),
    .A2(_3053_));
 sg13g2_nand2_1 _3894_ (.Y(_0424_),
    .A(net997),
    .B(_3068_));
 sg13g2_nand3_1 _3895_ (.B(_0423_),
    .C(_0424_),
    .A(_0422_),
    .Y(_0425_));
 sg13g2_nand2_1 _3896_ (.Y(_0426_),
    .A(net998),
    .B(_3053_));
 sg13g2_a22oi_1 _3897_ (.Y(_0427_),
    .B1(_3083_),
    .B2(net994),
    .A2(_3073_),
    .A1(net997));
 sg13g2_nand3_1 _3898_ (.B(_0426_),
    .C(_0427_),
    .A(_3112_),
    .Y(_0428_));
 sg13g2_nor4_2 _3899_ (.A(_0417_),
    .B(_0420_),
    .C(_0425_),
    .Y(_0429_),
    .D(_0428_));
 sg13g2_o21ai_1 _3900_ (.B1(net997),
    .Y(_0430_),
    .A1(_3073_),
    .A2(_3076_));
 sg13g2_nand2_2 _3901_ (.Y(_0431_),
    .A(_0411_),
    .B(_0427_));
 sg13g2_o21ai_1 _3902_ (.B1(net998),
    .Y(_0432_),
    .A1(_3053_),
    .A2(_3092_));
 sg13g2_nand2_2 _3903_ (.Y(_0433_),
    .A(_3038_),
    .B(net993));
 sg13g2_a21oi_1 _3904_ (.A1(net993),
    .A2(_3042_),
    .Y(_0434_),
    .B1(_0413_));
 sg13g2_nand2_1 _3905_ (.Y(_0435_),
    .A(_0433_),
    .B(_0434_));
 sg13g2_nor2_1 _3906_ (.A(_0431_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_and4_1 _3907_ (.A(_3077_),
    .B(_3098_),
    .C(_0432_),
    .D(_0436_),
    .X(_0437_));
 sg13g2_nand2_1 _3908_ (.Y(_0438_),
    .A(net966),
    .B(_0406_));
 sg13g2_nand3_1 _3909_ (.B(_0406_),
    .C(_0437_),
    .A(net966),
    .Y(_0439_));
 sg13g2_nand2b_1 _3910_ (.Y(_0440_),
    .B(_0439_),
    .A_N(_0429_));
 sg13g2_nand2_1 _3911_ (.Y(_0441_),
    .A(_0409_),
    .B(_0440_));
 sg13g2_nor2b_2 _3912_ (.A(\dtop.field_top.afl_sub_pc[1] ),
    .B_N(net1059),
    .Y(_0442_));
 sg13g2_nand2_1 _3913_ (.Y(_0443_),
    .A(net1059),
    .B(_2861_));
 sg13g2_a22oi_1 _3914_ (.Y(_0444_),
    .B1(_0437_),
    .B2(_3111_),
    .A2(_0429_),
    .A1(_3060_));
 sg13g2_nand2_2 _3915_ (.Y(_0445_),
    .A(_0442_),
    .B(_0444_));
 sg13g2_nor2_2 _3916_ (.A(_0441_),
    .B(_0445_),
    .Y(_0446_));
 sg13g2_inv_1 _3917_ (.Y(_0447_),
    .A(_0446_));
 sg13g2_o21ai_1 _3918_ (.B1(_3091_),
    .Y(_0448_),
    .A1(net970),
    .A2(_0402_));
 sg13g2_nand2b_1 _3919_ (.Y(_0449_),
    .B(net686),
    .A_N(net1059));
 sg13g2_or2_1 _3920_ (.X(_0450_),
    .B(_0449_),
    .A(_0448_));
 sg13g2_nor3_2 _3921_ (.A(net1008),
    .B(_0409_),
    .C(_0440_),
    .Y(_0451_));
 sg13g2_nand3b_1 _3922_ (.B(_0448_),
    .C(_0442_),
    .Y(_0452_),
    .A_N(_0444_));
 sg13g2_nor2_2 _3923_ (.A(_0406_),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_inv_1 _3924_ (.Y(_0454_),
    .A(_0453_));
 sg13g2_a21oi_2 _3925_ (.B1(_0452_),
    .Y(_0455_),
    .A2(_0441_),
    .A1(_0406_));
 sg13g2_nor2_1 _3926_ (.A(_0446_),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_nand2b_1 _3927_ (.Y(_0457_),
    .B(_0456_),
    .A_N(_0451_));
 sg13g2_nor2b_1 _3928_ (.A(_0457_),
    .B_N(_0450_),
    .Y(_0458_));
 sg13g2_inv_4 _3929_ (.A(net879),
    .Y(_0459_));
 sg13g2_nor2_1 _3930_ (.A(_0446_),
    .B(net878),
    .Y(_0460_));
 sg13g2_nand2_2 _3931_ (.Y(_0461_),
    .A(_0447_),
    .B(_0459_));
 sg13g2_nor2b_1 _3932_ (.A(net1058),
    .B_N(_0451_),
    .Y(_0462_));
 sg13g2_nand2b_2 _3933_ (.Y(_0463_),
    .B(_0451_),
    .A_N(net1058));
 sg13g2_and2_2 _3934_ (.A(net1058),
    .B(_0451_),
    .X(_0464_));
 sg13g2_nand2_2 _3935_ (.Y(_0465_),
    .A(net1058),
    .B(_0451_));
 sg13g2_o21ai_1 _3936_ (.B1(net909),
    .Y(_0466_),
    .A1(_0443_),
    .A2(_0448_));
 sg13g2_inv_1 _3937_ (.Y(_0467_),
    .A(_0466_));
 sg13g2_and3_2 _3938_ (.X(_0468_),
    .A(_0450_),
    .B(_0456_),
    .C(_0467_));
 sg13g2_nand3_1 _3939_ (.B(_0456_),
    .C(_0467_),
    .A(_0450_),
    .Y(_0469_));
 sg13g2_nand2_1 _3940_ (.Y(_0470_),
    .A(net1058),
    .B(_0467_));
 sg13g2_nand3_1 _3941_ (.B(_0440_),
    .C(_0470_),
    .A(\dtop.field_top.afl_alu.p ),
    .Y(_0471_));
 sg13g2_nand2_1 _3942_ (.Y(_0472_),
    .A(_0469_),
    .B(_0471_));
 sg13g2_o21ai_1 _3943_ (.B1(_0451_),
    .Y(_0473_),
    .A1(net1058),
    .A2(\dtop.field_top.afl_alu.p ));
 sg13g2_inv_1 _3944_ (.Y(_0474_),
    .A(net906));
 sg13g2_nand2_1 _3945_ (.Y(_0475_),
    .A(_3046_),
    .B(_3054_));
 sg13g2_nand4_1 _3946_ (.B(_3095_),
    .C(_3096_),
    .A(_3094_),
    .Y(_0476_),
    .D(_0419_));
 sg13g2_nor4_2 _3947_ (.A(_0425_),
    .B(_0428_),
    .C(_0475_),
    .Y(_0477_),
    .D(_0476_));
 sg13g2_and4_1 _3948_ (.A(net970),
    .B(_3074_),
    .C(_3102_),
    .D(_0418_),
    .X(_0478_));
 sg13g2_and4_1 _3949_ (.A(_3043_),
    .B(_0403_),
    .C(_0477_),
    .D(_0478_),
    .X(_0479_));
 sg13g2_nand2_1 _3950_ (.Y(_0480_),
    .A(_3087_),
    .B(_3099_));
 sg13g2_nand3_1 _3951_ (.B(_3098_),
    .C(_0432_),
    .A(_3052_),
    .Y(_0481_));
 sg13g2_nand2_1 _3952_ (.Y(_0482_),
    .A(_3109_),
    .B(_0403_));
 sg13g2_nor4_2 _3953_ (.A(_0435_),
    .B(_0480_),
    .C(_0481_),
    .Y(_0483_),
    .D(_0482_));
 sg13g2_o21ai_1 _3954_ (.B1(net997),
    .Y(_0484_),
    .A1(_3042_),
    .A2(_3086_));
 sg13g2_nand2_1 _3955_ (.Y(_0485_),
    .A(_3072_),
    .B(_0484_));
 sg13g2_nand3_1 _3956_ (.B(_3077_),
    .C(_3112_),
    .A(_3046_),
    .Y(_0486_));
 sg13g2_nor4_2 _3957_ (.A(_3037_),
    .B(_0431_),
    .C(_0485_),
    .Y(_0487_),
    .D(_0486_));
 sg13g2_nor3_1 _3958_ (.A(_3108_),
    .B(_0404_),
    .C(_0481_),
    .Y(_0488_));
 sg13g2_nor2_1 _3959_ (.A(_0435_),
    .B(_0480_),
    .Y(_0489_));
 sg13g2_nand2_1 _3960_ (.Y(_0490_),
    .A(_0483_),
    .B(_0487_));
 sg13g2_a21oi_1 _3961_ (.A1(net997),
    .A2(_3086_),
    .Y(_0491_),
    .B1(_3113_));
 sg13g2_a221oi_1 _3962_ (.B2(_0487_),
    .C1(_3113_),
    .B1(_0483_),
    .A1(net997),
    .Y(_0492_),
    .A2(_3086_));
 sg13g2_nor2_1 _3963_ (.A(_3037_),
    .B(net968),
    .Y(_0493_));
 sg13g2_and4_1 _3964_ (.A(_0488_),
    .B(_0489_),
    .C(_0491_),
    .D(_0493_),
    .X(_0494_));
 sg13g2_a21oi_1 _3965_ (.A1(_0490_),
    .A2(_0494_),
    .Y(_0495_),
    .B1(_0479_));
 sg13g2_a21o_1 _3966_ (.A2(_0494_),
    .A1(_0490_),
    .B1(_0479_),
    .X(_0496_));
 sg13g2_a21oi_1 _3967_ (.A1(_3029_),
    .A2(net990),
    .Y(_0497_),
    .B1(_3101_));
 sg13g2_nand4_1 _3968_ (.B(_3036_),
    .C(_3043_),
    .A(_3031_),
    .Y(_0498_),
    .D(_0403_));
 sg13g2_nand3_1 _3969_ (.B(_3102_),
    .C(_0418_),
    .A(_3084_),
    .Y(_0499_));
 sg13g2_nor3_1 _3970_ (.A(_0415_),
    .B(_0498_),
    .C(_0499_),
    .Y(_0500_));
 sg13g2_nand3_1 _3971_ (.B(_0497_),
    .C(_0500_),
    .A(_0477_),
    .Y(_0501_));
 sg13g2_nand3_1 _3972_ (.B(_3052_),
    .C(_3055_),
    .A(_3049_),
    .Y(_0502_));
 sg13g2_nand3_1 _3973_ (.B(_3074_),
    .C(_0410_),
    .A(_3072_),
    .Y(_0503_));
 sg13g2_or2_1 _3974_ (.X(_0504_),
    .B(_0503_),
    .A(_0502_));
 sg13g2_and4_1 _3975_ (.A(_0410_),
    .B(_0416_),
    .C(_0477_),
    .D(_0497_),
    .X(_0505_));
 sg13g2_o21ai_1 _3976_ (.B1(_0505_),
    .Y(_0506_),
    .A1(_0501_),
    .A2(_0504_));
 sg13g2_nor4_1 _3977_ (.A(_3069_),
    .B(_0480_),
    .C(_0481_),
    .D(_0486_),
    .Y(_0507_));
 sg13g2_nand4_1 _3978_ (.B(_0430_),
    .C(_0490_),
    .A(net967),
    .Y(_0508_),
    .D(_0507_));
 sg13g2_nand2_1 _3979_ (.Y(_0509_),
    .A(_0506_),
    .B(_0508_));
 sg13g2_and3_2 _3980_ (.X(_0510_),
    .A(_0496_),
    .B(_0506_),
    .C(_0508_));
 sg13g2_nor3_1 _3981_ (.A(_3037_),
    .B(net969),
    .C(_0431_),
    .Y(_0511_));
 sg13g2_nor2_2 _3982_ (.A(_0416_),
    .B(_0511_),
    .Y(_0512_));
 sg13g2_nor4_1 _3983_ (.A(_0425_),
    .B(_0428_),
    .C(_0475_),
    .D(_0498_),
    .Y(_0513_));
 sg13g2_and2_1 _3984_ (.A(_3075_),
    .B(_0513_),
    .X(_0514_));
 sg13g2_o21ai_1 _3985_ (.B1(_0514_),
    .Y(_0515_),
    .A1(_0501_),
    .A2(_0504_));
 sg13g2_nand4_1 _3986_ (.B(_3072_),
    .C(_3112_),
    .A(net967),
    .Y(_0516_),
    .D(_0488_));
 sg13g2_and2_1 _3987_ (.A(_0515_),
    .B(_0516_),
    .X(_0517_));
 sg13g2_nand2_1 _3988_ (.Y(_0518_),
    .A(_3107_),
    .B(_0492_));
 sg13g2_nand2_1 _3989_ (.Y(_0519_),
    .A(net968),
    .B(_0501_));
 sg13g2_or2_1 _3990_ (.X(_0520_),
    .B(_0501_),
    .A(net967));
 sg13g2_nand2_1 _3991_ (.Y(_0521_),
    .A(_3112_),
    .B(_0484_));
 sg13g2_a21oi_1 _3992_ (.A1(_0483_),
    .A2(_0487_),
    .Y(_0522_),
    .B1(_0521_));
 sg13g2_or2_1 _3993_ (.X(_0523_),
    .B(_0522_),
    .A(net968));
 sg13g2_a22oi_1 _3994_ (.Y(_0524_),
    .B1(_0501_),
    .B2(net968),
    .A2(_0492_),
    .A1(_3107_));
 sg13g2_a21o_1 _3995_ (.A2(_0516_),
    .A1(_0515_),
    .B1(_0524_),
    .X(_0525_));
 sg13g2_a221oi_1 _3996_ (.B2(_0519_),
    .C1(_0512_),
    .B1(_0518_),
    .A1(_0515_),
    .Y(_0526_),
    .A2(_0516_));
 sg13g2_and2_1 _3997_ (.A(_0510_),
    .B(_0526_),
    .X(_0527_));
 sg13g2_a21oi_2 _3998_ (.B1(_0496_),
    .Y(_0528_),
    .A2(_0508_),
    .A1(_0506_));
 sg13g2_and2_2 _3999_ (.A(_0526_),
    .B(_0528_),
    .X(_0529_));
 sg13g2_o21ai_1 _4000_ (.B1(_0526_),
    .Y(_0530_),
    .A1(_0510_),
    .A2(_0528_));
 sg13g2_a21oi_2 _4001_ (.B1(_0495_),
    .Y(_0531_),
    .A2(_0508_),
    .A1(_0506_));
 sg13g2_a22oi_1 _4002_ (.Y(_0532_),
    .B1(_0520_),
    .B2(_0523_),
    .A2(_0516_),
    .A1(_0515_));
 sg13g2_a22oi_1 _4003_ (.Y(_0533_),
    .B1(_0531_),
    .B2(_0532_),
    .A2(_0512_),
    .A1(_0510_));
 sg13g2_nand3_1 _4004_ (.B(_0506_),
    .C(_0508_),
    .A(_0495_),
    .Y(_0534_));
 sg13g2_and3_2 _4005_ (.X(_0535_),
    .A(_0515_),
    .B(_0516_),
    .C(_0524_));
 sg13g2_nand3_1 _4006_ (.B(_0516_),
    .C(_0524_),
    .A(_0515_),
    .Y(_0536_));
 sg13g2_nand2b_2 _4007_ (.Y(_0537_),
    .B(_0535_),
    .A_N(_0534_));
 sg13g2_nand2_1 _4008_ (.Y(_0538_),
    .A(_0512_),
    .B(_0528_));
 sg13g2_nand4_1 _4009_ (.B(_0533_),
    .C(_0537_),
    .A(_0530_),
    .Y(_0539_),
    .D(_0538_));
 sg13g2_nor3_1 _4010_ (.A(_0512_),
    .B(_0525_),
    .C(_0534_),
    .Y(_0540_));
 sg13g2_and2_1 _4011_ (.A(_0510_),
    .B(_0535_),
    .X(_0541_));
 sg13g2_nor2b_1 _4012_ (.A(_0524_),
    .B_N(_0517_),
    .Y(_0542_));
 sg13g2_or2_1 _4013_ (.X(_0543_),
    .B(_0542_),
    .A(_0541_));
 sg13g2_nor4_2 _4014_ (.A(_0047_),
    .B(_0539_),
    .C(net923),
    .Y(_0544_),
    .D(_0543_));
 sg13g2_a221oi_1 _4015_ (.B2(_0523_),
    .C1(_0496_),
    .B1(_0520_),
    .A1(_0515_),
    .Y(_0545_),
    .A2(_0516_));
 sg13g2_a21oi_1 _4016_ (.A1(_0531_),
    .A2(_0535_),
    .Y(_0546_),
    .B1(_0545_));
 sg13g2_a21o_1 _4017_ (.A2(_0535_),
    .A1(_0531_),
    .B1(_0545_),
    .X(_0547_));
 sg13g2_nand2_1 _4018_ (.Y(_0548_),
    .A(_0512_),
    .B(_0531_));
 sg13g2_and3_1 _4019_ (.X(_0549_),
    .A(_0510_),
    .B(_0525_),
    .C(_0536_));
 sg13g2_nand3_1 _4020_ (.B(_0525_),
    .C(_0536_),
    .A(_0510_),
    .Y(_0550_));
 sg13g2_nand3_1 _4021_ (.B(_0548_),
    .C(_0550_),
    .A(_0546_),
    .Y(_0551_));
 sg13g2_nand2_1 _4022_ (.Y(_0552_),
    .A(_0517_),
    .B(_0528_));
 sg13g2_nand2_1 _4023_ (.Y(_0553_),
    .A(_0528_),
    .B(_0535_));
 sg13g2_nand4_1 _4024_ (.B(_0548_),
    .C(_0550_),
    .A(_0546_),
    .Y(_0554_),
    .D(_0553_));
 sg13g2_nand2_1 _4025_ (.Y(_0555_),
    .A(\dtop.field_top.reg3[11] ),
    .B(net925));
 sg13g2_nand2_1 _4026_ (.Y(_0556_),
    .A(_0537_),
    .B(_0555_));
 sg13g2_nand2_1 _4027_ (.Y(_0557_),
    .A(\dtop.field_top.reg4[11] ),
    .B(net921));
 sg13g2_nand2_1 _4028_ (.Y(_0558_),
    .A(\dtop.field_top.reg2[11] ),
    .B(net926));
 sg13g2_nand2_2 _4029_ (.Y(_0559_),
    .A(_0557_),
    .B(_0558_));
 sg13g2_nor4_2 _4030_ (.A(_0544_),
    .B(_0554_),
    .C(_0556_),
    .Y(_0560_),
    .D(_0559_));
 sg13g2_or4_2 _4031_ (.A(_0544_),
    .B(_0554_),
    .C(_0556_),
    .D(_0559_),
    .X(_0561_));
 sg13g2_nand2_1 _4032_ (.Y(_0562_),
    .A(_0046_),
    .B(net906));
 sg13g2_o21ai_1 _4033_ (.B1(_0562_),
    .Y(_0563_),
    .A1(net907),
    .A2(_0561_));
 sg13g2_o21ai_1 _4034_ (.B1(_0037_),
    .Y(_0564_),
    .A1(_2875_),
    .A2(\dtop.field_top.acc[2] ));
 sg13g2_a21oi_2 _4035_ (.B1(_2879_),
    .Y(_0565_),
    .A2(_0564_),
    .A1(_0036_));
 sg13g2_o21ai_1 _4036_ (.B1(_0033_),
    .Y(_0566_),
    .A1(_2880_),
    .A2(_0565_));
 sg13g2_a21o_1 _4037_ (.A2(_0566_),
    .A1(_0032_),
    .B1(_2874_),
    .X(_0567_));
 sg13g2_a21oi_1 _4038_ (.A1(_0031_),
    .A2(_0567_),
    .Y(_0568_),
    .B1(\dtop.field_top.afl_alu.last_r_sum_msbs[0] ));
 sg13g2_nor3_2 _4039_ (.A(\dtop.field_top.afl_alu.last_r_sum_msbs[1] ),
    .B(_0465_),
    .C(_0568_),
    .Y(_0569_));
 sg13g2_or2_1 _4040_ (.X(_0570_),
    .B(_0569_),
    .A(_0455_));
 sg13g2_a21oi_2 _4041_ (.B1(_0570_),
    .Y(_0571_),
    .A2(_0563_),
    .A1(net909));
 sg13g2_nand3_1 _4042_ (.B(_3079_),
    .C(_3088_),
    .A(net970),
    .Y(_0572_));
 sg13g2_o21ai_1 _4043_ (.B1(_0572_),
    .Y(_0573_),
    .A1(_3057_),
    .A2(_0438_));
 sg13g2_nand2_1 _4044_ (.Y(_0574_),
    .A(net999),
    .B(_3083_));
 sg13g2_nand3_1 _4045_ (.B(_0573_),
    .C(_0574_),
    .A(net907),
    .Y(_0575_));
 sg13g2_nor2_1 _4046_ (.A(_0561_),
    .B(net892),
    .Y(_0576_));
 sg13g2_a21oi_2 _4047_ (.B1(_0576_),
    .Y(_0577_),
    .A2(net892),
    .A1(_0046_));
 sg13g2_nor4_1 _4048_ (.A(_0539_),
    .B(net923),
    .C(_0543_),
    .D(_0554_),
    .Y(_0578_));
 sg13g2_inv_2 _4049_ (.Y(_0579_),
    .A(net890));
 sg13g2_a221oi_1 _4050_ (.B2(_0509_),
    .C1(_0549_),
    .B1(_0547_),
    .A1(_0510_),
    .Y(_0580_),
    .A2(_0512_));
 sg13g2_a22oi_1 _4051_ (.Y(_0581_),
    .B1(net925),
    .B2(\dtop.field_top.reg3[12] ),
    .A2(net927),
    .A1(\dtop.field_top.reg2[12] ));
 sg13g2_nand2_1 _4052_ (.Y(_0582_),
    .A(_0580_),
    .B(_0581_));
 sg13g2_a221oi_1 _4053_ (.B2(_2883_),
    .C1(_0582_),
    .B1(net890),
    .A1(\dtop.field_top.reg4[12] ),
    .Y(_0583_),
    .A2(net922));
 sg13g2_mux2_1 _4054_ (.A0(_0583_),
    .A1(_0044_),
    .S(net892),
    .X(_0584_));
 sg13g2_mux4_1 _4055_ (.S0(_0454_),
    .A0(_0583_),
    .A1(_0560_),
    .A2(_0044_),
    .A3(_0046_),
    .S1(net892),
    .X(_0585_));
 sg13g2_xnor2_1 _4056_ (.Y(_0586_),
    .A(_0469_),
    .B(_0585_));
 sg13g2_nor2b_1 _4057_ (.A(_0586_),
    .B_N(_0571_),
    .Y(_0587_));
 sg13g2_xnor2_1 _4058_ (.Y(_0588_),
    .A(_0571_),
    .B(_0586_));
 sg13g2_xnor2_1 _4059_ (.Y(_0589_),
    .A(_0472_),
    .B(_0588_));
 sg13g2_inv_1 _4060_ (.Y(_0590_),
    .A(_0589_));
 sg13g2_o21ai_1 _4061_ (.B1(_0460_),
    .Y(_0591_),
    .A1(_0463_),
    .A2(_0571_));
 sg13g2_a21oi_1 _4062_ (.A1(_0463_),
    .A2(_0589_),
    .Y(_0592_),
    .B1(_0591_));
 sg13g2_nor3_1 _4063_ (.A(\dtop.field_top.afl_alu.last_r_sum_msbs[0] ),
    .B(\dtop.field_top.afl_alu.last_r_sum_msbs[1] ),
    .C(_0465_),
    .Y(_0593_));
 sg13g2_or3_2 _4064_ (.A(\dtop.field_top.afl_alu.last_r_sum_msbs[0] ),
    .B(\dtop.field_top.afl_alu.last_r_sum_msbs[1] ),
    .C(net909),
    .X(_0594_));
 sg13g2_nor2_2 _4065_ (.A(_0455_),
    .B(_0464_),
    .Y(_0595_));
 sg13g2_nand2b_2 _4066_ (.Y(_0596_),
    .B(net909),
    .A_N(_0455_));
 sg13g2_nand2b_1 _4067_ (.Y(_0597_),
    .B(net906),
    .A_N(_0038_));
 sg13g2_a21o_1 _4068_ (.A2(_0512_),
    .A1(_0510_),
    .B1(_0551_),
    .X(_0598_));
 sg13g2_and2_1 _4069_ (.A(\dtop.field_top.reg3[15] ),
    .B(net925),
    .X(_0599_));
 sg13g2_a22oi_1 _4070_ (.Y(_0600_),
    .B1(net922),
    .B2(\dtop.field_top.reg4[15] ),
    .A2(net927),
    .A1(\dtop.field_top.reg2[15] ));
 sg13g2_o21ai_1 _4071_ (.B1(_0600_),
    .Y(_0601_),
    .A1(_0039_),
    .A2(_0579_));
 sg13g2_nor3_2 _4072_ (.A(_0598_),
    .B(_0599_),
    .C(_0601_),
    .Y(_0602_));
 sg13g2_o21ai_1 _4073_ (.B1(_0597_),
    .Y(_0603_),
    .A1(net906),
    .A2(_0602_));
 sg13g2_nor2_1 _4074_ (.A(\dtop.field_top.afl_alu.last_r_sum_msbs[0] ),
    .B(\dtop.field_top.afl_alu.last_r_sum_msbs[1] ),
    .Y(_0604_));
 sg13g2_and2_2 _4075_ (.A(_0464_),
    .B(_0604_),
    .X(_0605_));
 sg13g2_nand2_1 _4076_ (.Y(_0606_),
    .A(_0464_),
    .B(_0604_));
 sg13g2_a21o_1 _4077_ (.A2(_0603_),
    .A1(_0595_),
    .B1(net888),
    .X(_0607_));
 sg13g2_mux2_1 _4078_ (.A0(_0602_),
    .A1(_0038_),
    .S(net891),
    .X(_0608_));
 sg13g2_xnor2_1 _4079_ (.Y(_0609_),
    .A(_0468_),
    .B(_0608_));
 sg13g2_and2_1 _4080_ (.A(_0607_),
    .B(_0609_),
    .X(_0610_));
 sg13g2_nor2b_1 _4081_ (.A(_0041_),
    .B_N(net890),
    .Y(_0611_));
 sg13g2_nand2_2 _4082_ (.Y(_0612_),
    .A(\dtop.field_top.reg4[14] ),
    .B(net921));
 sg13g2_a22oi_1 _4083_ (.Y(_0613_),
    .B1(net924),
    .B2(\dtop.field_top.reg3[14] ),
    .A2(net926),
    .A1(\dtop.field_top.reg2[14] ));
 sg13g2_nand3_1 _4084_ (.B(_0612_),
    .C(_0613_),
    .A(_0537_),
    .Y(_0614_));
 sg13g2_nor3_2 _4085_ (.A(_0598_),
    .B(_0611_),
    .C(_0614_),
    .Y(_0615_));
 sg13g2_nand2b_1 _4086_ (.Y(_0616_),
    .B(net907),
    .A_N(_0040_));
 sg13g2_o21ai_1 _4087_ (.B1(_0616_),
    .Y(_0617_),
    .A1(net907),
    .A2(_0615_));
 sg13g2_nor3_2 _4088_ (.A(\dtop.field_top.acc[5] ),
    .B(\dtop.field_top.acc[4] ),
    .C(\dtop.field_top.acc[3] ),
    .Y(_0618_));
 sg13g2_nor3_1 _4089_ (.A(\dtop.field_top.acc[9] ),
    .B(\dtop.field_top.acc[8] ),
    .C(\dtop.field_top.acc[7] ),
    .Y(_0619_));
 sg13g2_nand2_1 _4090_ (.Y(_0620_),
    .A(_0618_),
    .B(_0619_));
 sg13g2_nor2_1 _4091_ (.A(\dtop.field_top.acc[6] ),
    .B(_0620_),
    .Y(_0621_));
 sg13g2_nand2_2 _4092_ (.Y(_0622_),
    .A(_0031_),
    .B(_0621_));
 sg13g2_nand2_1 _4093_ (.Y(_0623_),
    .A(net887),
    .B(_0622_));
 sg13g2_nand2_1 _4094_ (.Y(_0624_),
    .A(_0605_),
    .B(_0622_));
 sg13g2_a22oi_1 _4095_ (.Y(_0625_),
    .B1(_0622_),
    .B2(net888),
    .A2(_0617_),
    .A1(_0595_));
 sg13g2_mux2_1 _4096_ (.A0(_0615_),
    .A1(_0040_),
    .S(net891),
    .X(_0626_));
 sg13g2_and2_1 _4097_ (.A(_0454_),
    .B(_0626_),
    .X(_0627_));
 sg13g2_a21oi_1 _4098_ (.A1(_0453_),
    .A2(_0608_),
    .Y(_0628_),
    .B1(_0627_));
 sg13g2_xnor2_1 _4099_ (.Y(_0629_),
    .A(_0468_),
    .B(_0628_));
 sg13g2_or2_1 _4100_ (.X(_0630_),
    .B(_0629_),
    .A(_0625_));
 sg13g2_nand2b_1 _4101_ (.Y(_0631_),
    .B(net906),
    .A_N(_0042_));
 sg13g2_a22oi_1 _4102_ (.Y(_0632_),
    .B1(net921),
    .B2(\dtop.field_top.reg4[13] ),
    .A2(net924),
    .A1(\dtop.field_top.reg3[13] ));
 sg13g2_nand2_1 _4103_ (.Y(_0633_),
    .A(\dtop.field_top.reg2[13] ),
    .B(net927));
 sg13g2_nand3_1 _4104_ (.B(_0632_),
    .C(_0633_),
    .A(_0580_),
    .Y(_0634_));
 sg13g2_a21oi_2 _4105_ (.B1(_0634_),
    .Y(_0635_),
    .A2(net889),
    .A1(_2882_));
 sg13g2_o21ai_1 _4106_ (.B1(_0631_),
    .Y(_0636_),
    .A1(net907),
    .A2(_0635_));
 sg13g2_nand2_1 _4107_ (.Y(_0637_),
    .A(_0031_),
    .B(_0619_));
 sg13g2_a21oi_2 _4108_ (.B1(_0637_),
    .Y(_0638_),
    .A2(_0618_),
    .A1(_0034_));
 sg13g2_nor2_2 _4109_ (.A(_0594_),
    .B(_0638_),
    .Y(_0639_));
 sg13g2_a21oi_1 _4110_ (.A1(_0595_),
    .A2(_0636_),
    .Y(_0640_),
    .B1(_0639_));
 sg13g2_mux2_1 _4111_ (.A0(_0635_),
    .A1(_0042_),
    .S(net892),
    .X(_0641_));
 sg13g2_and2_1 _4112_ (.A(_0454_),
    .B(_0641_),
    .X(_0642_));
 sg13g2_a21oi_1 _4113_ (.A1(_0453_),
    .A2(_0626_),
    .Y(_0643_),
    .B1(_0642_));
 sg13g2_xnor2_1 _4114_ (.Y(_0644_),
    .A(_0468_),
    .B(_0643_));
 sg13g2_nor2_1 _4115_ (.A(_0640_),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_and2_1 _4116_ (.A(_0044_),
    .B(net907),
    .X(_0646_));
 sg13g2_a21oi_1 _4117_ (.A1(net895),
    .A2(_0583_),
    .Y(_0647_),
    .B1(_0646_));
 sg13g2_nor2_2 _4118_ (.A(\dtop.field_top.acc[1] ),
    .B(\dtop.field_top.acc[2] ),
    .Y(_0648_));
 sg13g2_nor2_1 _4119_ (.A(\dtop.field_top.acc[3] ),
    .B(_0648_),
    .Y(_0649_));
 sg13g2_a21oi_2 _4120_ (.B1(\dtop.field_top.acc[5] ),
    .Y(_0650_),
    .A2(_0649_),
    .A1(_0036_));
 sg13g2_a21oi_1 _4121_ (.A1(_0034_),
    .A2(_0650_),
    .Y(_0651_),
    .B1(\dtop.field_top.acc[7] ));
 sg13g2_a21oi_1 _4122_ (.A1(_0032_),
    .A2(_0651_),
    .Y(_0652_),
    .B1(\dtop.field_top.acc[9] ));
 sg13g2_nand2_2 _4123_ (.Y(_0653_),
    .A(_0031_),
    .B(_0652_));
 sg13g2_nand2_1 _4124_ (.Y(_0654_),
    .A(net888),
    .B(_0653_));
 sg13g2_nand2_1 _4125_ (.Y(_0655_),
    .A(_0605_),
    .B(_0653_));
 sg13g2_a22oi_1 _4126_ (.Y(_0656_),
    .B1(_0653_),
    .B2(net888),
    .A2(_0647_),
    .A1(_0595_));
 sg13g2_mux2_1 _4127_ (.A0(_0584_),
    .A1(_0641_),
    .S(_0453_),
    .X(_0657_));
 sg13g2_xnor2_1 _4128_ (.Y(_0658_),
    .A(_0469_),
    .B(_0657_));
 sg13g2_or2_1 _4129_ (.X(_0659_),
    .B(_0658_),
    .A(_0656_));
 sg13g2_a21oi_1 _4130_ (.A1(_0472_),
    .A2(_0588_),
    .Y(_0660_),
    .B1(_0587_));
 sg13g2_xnor2_1 _4131_ (.Y(_0661_),
    .A(_0656_),
    .B(_0658_));
 sg13g2_o21ai_1 _4132_ (.B1(_0659_),
    .Y(_0662_),
    .A1(_0660_),
    .A2(_0661_));
 sg13g2_nand2_1 _4133_ (.Y(_0663_),
    .A(_0640_),
    .B(_0644_));
 sg13g2_nand2b_1 _4134_ (.Y(_0664_),
    .B(_0663_),
    .A_N(_0645_));
 sg13g2_a21oi_1 _4135_ (.A1(_0662_),
    .A2(_0663_),
    .Y(_0665_),
    .B1(_0645_));
 sg13g2_xnor2_1 _4136_ (.Y(_0666_),
    .A(_0625_),
    .B(_0629_));
 sg13g2_o21ai_1 _4137_ (.B1(_0630_),
    .Y(_0667_),
    .A1(_0665_),
    .A2(_0666_));
 sg13g2_xor2_1 _4138_ (.B(_0609_),
    .A(_0607_),
    .X(_0668_));
 sg13g2_nand2b_1 _4139_ (.Y(_0669_),
    .B(_0668_),
    .A_N(_0667_));
 sg13g2_xnor2_1 _4140_ (.Y(_0670_),
    .A(_0667_),
    .B(_0668_));
 sg13g2_xor2_1 _4141_ (.B(_0668_),
    .A(_0667_),
    .X(_0671_));
 sg13g2_nor2_1 _4142_ (.A(net911),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_inv_1 _4143_ (.Y(_0673_),
    .A(_0672_));
 sg13g2_nand2_1 _4144_ (.Y(_0674_),
    .A(_0621_),
    .B(_0648_));
 sg13g2_nor4_1 _4145_ (.A(\dtop.field_top.acc[10] ),
    .B(\dtop.field_top.acc[0] ),
    .C(_0594_),
    .D(_0674_),
    .Y(_0675_));
 sg13g2_a21oi_2 _4146_ (.B1(_0675_),
    .Y(_0676_),
    .A2(_0672_),
    .A1(_0610_));
 sg13g2_inv_2 _4147_ (.Y(_0677_),
    .A(_0676_));
 sg13g2_nand2b_1 _4148_ (.Y(_0678_),
    .B(_0669_),
    .A_N(_0610_));
 sg13g2_a22oi_1 _4149_ (.Y(_0679_),
    .B1(_0592_),
    .B2(_0676_),
    .A2(_0461_),
    .A1(net655));
 sg13g2_inv_1 _4150_ (.Y(_0127_),
    .A(_0679_));
 sg13g2_xor2_1 _4151_ (.B(_0661_),
    .A(_0660_),
    .X(_0680_));
 sg13g2_nand2_1 _4152_ (.Y(_0681_),
    .A(net910),
    .B(_0656_));
 sg13g2_o21ai_1 _4153_ (.B1(_0676_),
    .Y(_0682_),
    .A1(net910),
    .A2(_0680_));
 sg13g2_nor2_1 _4154_ (.A(_0461_),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_a22oi_1 _4155_ (.Y(_0684_),
    .B1(_0681_),
    .B2(_0683_),
    .A2(_0461_),
    .A1(net553));
 sg13g2_inv_1 _4156_ (.Y(_0128_),
    .A(_0684_));
 sg13g2_xor2_1 _4157_ (.B(_0664_),
    .A(_0662_),
    .X(_0685_));
 sg13g2_nand2_1 _4158_ (.Y(_0686_),
    .A(net910),
    .B(_0640_));
 sg13g2_nand3_1 _4159_ (.B(_0676_),
    .C(_0686_),
    .A(_0460_),
    .Y(_0687_));
 sg13g2_a21oi_1 _4160_ (.A1(_0463_),
    .A2(_0685_),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_a21o_1 _4161_ (.A2(_0461_),
    .A1(net638),
    .B1(_0688_),
    .X(_0129_));
 sg13g2_xor2_1 _4162_ (.B(_0666_),
    .A(_0665_),
    .X(_0689_));
 sg13g2_nand2_1 _4163_ (.Y(_0690_),
    .A(net910),
    .B(_0625_));
 sg13g2_o21ai_1 _4164_ (.B1(_0690_),
    .Y(_0691_),
    .A1(net910),
    .A2(_0689_));
 sg13g2_nor2_1 _4165_ (.A(_0461_),
    .B(_0691_),
    .Y(_0692_));
 sg13g2_a22oi_1 _4166_ (.Y(_0693_),
    .B1(_0676_),
    .B2(_0692_),
    .A2(_0461_),
    .A1(net658));
 sg13g2_inv_1 _4167_ (.Y(_0130_),
    .A(_0693_));
 sg13g2_or2_1 _4168_ (.X(_0694_),
    .B(_0607_),
    .A(_0463_));
 sg13g2_a21oi_1 _4169_ (.A1(_0673_),
    .A2(_0694_),
    .Y(_0695_),
    .B1(_0461_));
 sg13g2_a22oi_1 _4170_ (.Y(_0131_),
    .B1(_0676_),
    .B2(_0695_),
    .A2(_0461_),
    .A1(_2881_));
 sg13g2_nand2_1 _4171_ (.Y(_0696_),
    .A(net671),
    .B(net878));
 sg13g2_and2_1 _4172_ (.A(_0531_),
    .B(_0542_),
    .X(_0697_));
 sg13g2_a22oi_1 _4173_ (.Y(_0698_),
    .B1(net905),
    .B2(\dtop.field_top.alt_osc[6] ),
    .A2(_0527_),
    .A1(\dtop.field_top.comp_values0[2][7] ));
 sg13g2_nor2_2 _4174_ (.A(_0524_),
    .B(_0552_),
    .Y(_0699_));
 sg13g2_a22oi_1 _4175_ (.Y(_0700_),
    .B1(net922),
    .B2(\dtop.field_top.comp_values0[4][7] ),
    .A2(_0529_),
    .A1(\dtop.field_top.comp_values0[3][7] ));
 sg13g2_nand2_1 _4176_ (.Y(_0701_),
    .A(_0698_),
    .B(_0700_));
 sg13g2_a221oi_1 _4177_ (.B2(\dtop.field_top.controller.timer[2] ),
    .C1(_0701_),
    .B1(_0699_),
    .A1(_2910_),
    .Y(_0702_),
    .A2(net889));
 sg13g2_nand2_1 _4178_ (.Y(_0703_),
    .A(_0033_),
    .B(net908));
 sg13g2_a21oi_1 _4179_ (.A1(net896),
    .A2(_0702_),
    .Y(_0704_),
    .B1(_0596_));
 sg13g2_nor2_2 _4180_ (.A(net911),
    .B(_0469_),
    .Y(_0705_));
 sg13g2_o21ai_1 _4181_ (.B1(net991),
    .Y(_0706_),
    .A1(_3042_),
    .A2(_3076_));
 sg13g2_o21ai_1 _4182_ (.B1(_0706_),
    .Y(_0707_),
    .A1(net1052),
    .A2(_0418_));
 sg13g2_nor2_1 _4183_ (.A(_0428_),
    .B(_0707_),
    .Y(_0708_));
 sg13g2_nand4_1 _4184_ (.B(_3077_),
    .C(_3098_),
    .A(net967),
    .Y(_0709_),
    .D(_0426_));
 sg13g2_nor2_1 _4185_ (.A(_0431_),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_a22oi_1 _4186_ (.Y(_0711_),
    .B1(_0710_),
    .B2(_0433_),
    .A2(_0708_),
    .A1(_0416_));
 sg13g2_nand2_1 _4187_ (.Y(_0712_),
    .A(net909),
    .B(_0711_));
 sg13g2_xnor2_1 _4188_ (.Y(_0713_),
    .A(_0053_),
    .B(_0712_));
 sg13g2_nor2_2 _4189_ (.A(_0054_),
    .B(_0579_),
    .Y(_0714_));
 sg13g2_o21ai_1 _4190_ (.B1(\dtop.field_top.sflag ),
    .Y(_0715_),
    .A1(_0541_),
    .A2(_0547_));
 sg13g2_nor2_1 _4191_ (.A(\dtop.field_top.sflag2 ),
    .B(_0537_),
    .Y(_0716_));
 sg13g2_a21oi_1 _4192_ (.A1(\dtop.field_top.controller.ppos[3] ),
    .A2(_0699_),
    .Y(_0717_),
    .B1(_0716_));
 sg13g2_nand2_2 _4193_ (.Y(_0718_),
    .A(\dtop.field_top.reg2[16] ),
    .B(net926));
 sg13g2_xnor2_1 _4194_ (.Y(_0719_),
    .A(\dtop.field_top.sflag ),
    .B(\dtop.field_top.sflag2 ));
 sg13g2_o21ai_1 _4195_ (.B1(_0718_),
    .Y(_0720_),
    .A1(_0553_),
    .A2(_0719_));
 sg13g2_a22oi_1 _4196_ (.Y(_0721_),
    .B1(net921),
    .B2(\dtop.field_top.reg4[16] ),
    .A2(net924),
    .A1(\dtop.field_top.reg3[16] ));
 sg13g2_nand3_1 _4197_ (.B(_0717_),
    .C(_0721_),
    .A(_0715_),
    .Y(_0722_));
 sg13g2_nor3_2 _4198_ (.A(_0714_),
    .B(_0720_),
    .C(_0722_),
    .Y(_0723_));
 sg13g2_mux2_2 _4199_ (.A0(_0723_),
    .A1(_0713_),
    .S(net894),
    .X(_0724_));
 sg13g2_inv_1 _4200_ (.Y(_0725_),
    .A(_0724_));
 sg13g2_mux2_1 _4201_ (.A0(_0713_),
    .A1(_0723_),
    .S(net896),
    .X(_0726_));
 sg13g2_inv_1 _4202_ (.Y(_0727_),
    .A(_0726_));
 sg13g2_xor2_1 _4203_ (.B(_0726_),
    .A(_0724_),
    .X(_0728_));
 sg13g2_nor2_1 _4204_ (.A(_3031_),
    .B(net966),
    .Y(_0729_));
 sg13g2_a221oi_1 _4205_ (.B2(_0446_),
    .C1(_0705_),
    .B1(_0729_),
    .A1(net911),
    .Y(_0730_),
    .A2(_0728_));
 sg13g2_inv_1 _4206_ (.Y(_0731_),
    .A(_0730_));
 sg13g2_o21ai_1 _4207_ (.B1(net910),
    .Y(_0732_),
    .A1(_0590_),
    .A2(_0671_));
 sg13g2_nand2_1 _4208_ (.Y(_0733_),
    .A(net966),
    .B(_3108_));
 sg13g2_nand2_2 _4209_ (.Y(_0734_),
    .A(_0445_),
    .B(_0705_));
 sg13g2_nand2b_2 _4210_ (.Y(_0735_),
    .B(_0734_),
    .A_N(_0733_));
 sg13g2_nand2_1 _4211_ (.Y(_0736_),
    .A(_0464_),
    .B(_0568_));
 sg13g2_a21oi_2 _4212_ (.B1(_0453_),
    .Y(_0737_),
    .A2(_0464_),
    .A1(\dtop.field_top.afl_alu.last_r_sum_msbs[1] ));
 sg13g2_and3_1 _4213_ (.X(_0738_),
    .A(_0735_),
    .B(_0736_),
    .C(_0737_));
 sg13g2_and2_1 _4214_ (.A(_0732_),
    .B(_0738_),
    .X(_0739_));
 sg13g2_nand2_1 _4215_ (.Y(_0740_),
    .A(_0732_),
    .B(_0738_));
 sg13g2_mux2_2 _4216_ (.A0(_0702_),
    .A1(_0033_),
    .S(net894),
    .X(_0741_));
 sg13g2_inv_1 _4217_ (.Y(_0742_),
    .A(_0741_));
 sg13g2_a22oi_1 _4218_ (.Y(_0743_),
    .B1(net922),
    .B2(\dtop.field_top.comp_values0[4][8] ),
    .A2(_0529_),
    .A1(\dtop.field_top.comp_values0[3][8] ));
 sg13g2_a22oi_1 _4219_ (.Y(_0744_),
    .B1(_0699_),
    .B2(\dtop.field_top.controller.ppos[0] ),
    .A2(_0527_),
    .A1(\dtop.field_top.comp_values0[2][8] ));
 sg13g2_nand2_1 _4220_ (.Y(_0745_),
    .A(_0743_),
    .B(_0744_));
 sg13g2_a221oi_1 _4221_ (.B2(\dtop.field_top.alt_osc[7] ),
    .C1(_0745_),
    .B1(_0697_),
    .A1(_2911_),
    .Y(_0746_),
    .A2(net890));
 sg13g2_nand2b_1 _4222_ (.Y(_0747_),
    .B(net893),
    .A_N(_0032_));
 sg13g2_o21ai_1 _4223_ (.B1(_0747_),
    .Y(_0748_),
    .A1(net893),
    .A2(_0746_));
 sg13g2_inv_1 _4224_ (.Y(_0749_),
    .A(_0748_));
 sg13g2_o21ai_1 _4225_ (.B1(net910),
    .Y(_0750_),
    .A1(_0671_),
    .A2(_0680_));
 sg13g2_nand2_1 _4226_ (.Y(_0751_),
    .A(_0654_),
    .B(_0750_));
 sg13g2_nand2_1 _4227_ (.Y(_0752_),
    .A(_0028_),
    .B(net890));
 sg13g2_nor2_1 _4228_ (.A(\dtop.field_top.masked_bits[0] ),
    .B(_0538_),
    .Y(_0753_));
 sg13g2_a221oi_1 _4229_ (.B2(net1060),
    .C1(_0753_),
    .B1(net905),
    .A1(\dtop.field_top.comp_values0[4][9] ),
    .Y(_0754_),
    .A2(net923));
 sg13g2_nand2_1 _4230_ (.Y(_0755_),
    .A(\dtop.field_top.comp_values0[2][9] ),
    .B(net927));
 sg13g2_a22oi_1 _4231_ (.Y(_0756_),
    .B1(_0699_),
    .B2(\dtop.field_top.controller.ppos[1] ),
    .A2(net925),
    .A1(\dtop.field_top.comp_values0[3][9] ));
 sg13g2_nand3_1 _4232_ (.B(_0755_),
    .C(_0756_),
    .A(_0754_),
    .Y(_0757_));
 sg13g2_o21ai_1 _4233_ (.B1(_0752_),
    .Y(_0758_),
    .A1(net890),
    .A2(_0757_));
 sg13g2_nand2_1 _4234_ (.Y(_0759_),
    .A(_2874_),
    .B(net893));
 sg13g2_o21ai_1 _4235_ (.B1(_0759_),
    .Y(_0760_),
    .A1(net893),
    .A2(_0758_));
 sg13g2_inv_1 _4236_ (.Y(_0761_),
    .A(_0760_));
 sg13g2_o21ai_1 _4237_ (.B1(_0552_),
    .Y(_0762_),
    .A1(_0534_),
    .A2(_0542_));
 sg13g2_nor4_1 _4238_ (.A(_0539_),
    .B(_0541_),
    .C(_0551_),
    .D(_0762_),
    .Y(_0763_));
 sg13g2_nor2_1 _4239_ (.A(\dtop.field_top.masked_bits[1] ),
    .B(_0538_),
    .Y(_0764_));
 sg13g2_a22oi_1 _4240_ (.Y(_0765_),
    .B1(net925),
    .B2(\dtop.field_top.comp_values0[3][10] ),
    .A2(net927),
    .A1(\dtop.field_top.comp_values0[2][10] ));
 sg13g2_a21oi_1 _4241_ (.A1(\dtop.field_top.controller.ppos[2] ),
    .A2(_0699_),
    .Y(_0766_),
    .B1(_0764_));
 sg13g2_a21oi_1 _4242_ (.A1(\dtop.field_top.comp_values0[4][10] ),
    .A2(net923),
    .Y(_0767_),
    .B1(_0763_));
 sg13g2_and3_1 _4243_ (.X(_0768_),
    .A(_0765_),
    .B(_0766_),
    .C(_0767_));
 sg13g2_a221oi_1 _4244_ (.B2(\dtop.field_top.rs.scan_y.pos[8] ),
    .C1(_0768_),
    .B1(net905),
    .A1(_0052_),
    .Y(_0769_),
    .A2(net889));
 sg13g2_nor2_1 _4245_ (.A(net893),
    .B(_0769_),
    .Y(_0770_));
 sg13g2_a21oi_2 _4246_ (.B1(_0770_),
    .Y(_0771_),
    .A2(net893),
    .A1(_0031_));
 sg13g2_mux4_1 _4247_ (.S0(net857),
    .A0(_0742_),
    .A1(_0748_),
    .A2(_0760_),
    .A3(_0771_),
    .S1(net854),
    .X(_0772_));
 sg13g2_nand2_1 _4248_ (.Y(_0773_),
    .A(_0670_),
    .B(_0685_));
 sg13g2_a21oi_2 _4249_ (.B1(_0463_),
    .Y(_0774_),
    .A2(_0685_),
    .A1(_0670_));
 sg13g2_nor2_1 _4250_ (.A(_0639_),
    .B(_0774_),
    .Y(_0775_));
 sg13g2_nor3_2 _4251_ (.A(_0594_),
    .B(_0639_),
    .C(_0774_),
    .Y(_0776_));
 sg13g2_a21oi_2 _4252_ (.B1(_0774_),
    .Y(_0777_),
    .A2(_0638_),
    .A1(net887));
 sg13g2_or2_2 _4253_ (.X(_0778_),
    .B(_0776_),
    .A(_0774_));
 sg13g2_nand3b_1 _4254_ (.B(_0638_),
    .C(_0605_),
    .Y(_0779_),
    .A_N(_0774_));
 sg13g2_a21oi_2 _4255_ (.B1(_0774_),
    .Y(_0780_),
    .A2(_0638_),
    .A1(_0605_));
 sg13g2_a21o_2 _4256_ (.A2(_0638_),
    .A1(_0605_),
    .B1(_0774_),
    .X(_0781_));
 sg13g2_and2_1 _4257_ (.A(_0772_),
    .B(_0777_),
    .X(_0782_));
 sg13g2_nand3_1 _4258_ (.B(_0626_),
    .C(_0641_),
    .A(_0584_),
    .Y(_0783_));
 sg13g2_nor3_1 _4259_ (.A(_0577_),
    .B(_0608_),
    .C(_0783_),
    .Y(_0784_));
 sg13g2_a21oi_2 _4260_ (.B1(_0784_),
    .Y(_0785_),
    .A2(_0724_),
    .A1(_0446_));
 sg13g2_a22oi_1 _4261_ (.Y(_0786_),
    .B1(net924),
    .B2(\dtop.field_top.comp_values0[3][0] ),
    .A2(net926),
    .A1(\dtop.field_top.comp_values0[2][0] ));
 sg13g2_o21ai_1 _4262_ (.B1(_0786_),
    .Y(_0787_),
    .A1(_0056_),
    .A2(_0579_));
 sg13g2_a21oi_2 _4263_ (.B1(_0787_),
    .Y(_0788_),
    .A2(net921),
    .A1(\dtop.field_top.comp_values0[4][0] ));
 sg13g2_nand2b_1 _4264_ (.Y(_0789_),
    .B(net893),
    .A_N(_0055_));
 sg13g2_o21ai_1 _4265_ (.B1(_0789_),
    .Y(_0790_),
    .A1(net893),
    .A2(_0788_));
 sg13g2_inv_1 _4266_ (.Y(_0791_),
    .A(_0790_));
 sg13g2_a22oi_1 _4267_ (.Y(_0792_),
    .B1(net924),
    .B2(\dtop.field_top.comp_values0[3][1] ),
    .A2(net926),
    .A1(\dtop.field_top.comp_values0[2][1] ));
 sg13g2_o21ai_1 _4268_ (.B1(_0792_),
    .Y(_0793_),
    .A1(_0030_),
    .A2(_0579_));
 sg13g2_a21oi_2 _4269_ (.B1(_0793_),
    .Y(_0794_),
    .A2(net921),
    .A1(\dtop.field_top.comp_values0[4][1] ));
 sg13g2_nand2_1 _4270_ (.Y(_0795_),
    .A(_2876_),
    .B(net891));
 sg13g2_o21ai_1 _4271_ (.B1(_0795_),
    .Y(_0796_),
    .A1(net891),
    .A2(_0794_));
 sg13g2_inv_1 _4272_ (.Y(_0797_),
    .A(_0796_));
 sg13g2_a22oi_1 _4273_ (.Y(_0798_),
    .B1(net905),
    .B2(\dtop.field_top.alt_osc[1] ),
    .A2(net926),
    .A1(\dtop.field_top.comp_values0[2][2] ));
 sg13g2_a22oi_1 _4274_ (.Y(_0799_),
    .B1(net921),
    .B2(\dtop.field_top.comp_values0[4][2] ),
    .A2(net924),
    .A1(\dtop.field_top.comp_values0[3][2] ));
 sg13g2_nand2_1 _4275_ (.Y(_0800_),
    .A(_0798_),
    .B(_0799_));
 sg13g2_a21oi_2 _4276_ (.B1(_0800_),
    .Y(_0801_),
    .A2(net889),
    .A1(_2887_));
 sg13g2_mux2_2 _4277_ (.A0(_0801_),
    .A1(_0048_),
    .S(net891),
    .X(_0802_));
 sg13g2_inv_1 _4278_ (.Y(_0803_),
    .A(_0802_));
 sg13g2_mux4_1 _4279_ (.S0(net856),
    .A0(_0785_),
    .A1(_0790_),
    .A2(_0796_),
    .A3(_0803_),
    .S1(net854),
    .X(_0804_));
 sg13g2_a21oi_1 _4280_ (.A1(_0778_),
    .A2(_0804_),
    .Y(_0805_),
    .B1(_0782_));
 sg13g2_o21ai_1 _4281_ (.B1(net910),
    .Y(_0806_),
    .A1(_0671_),
    .A2(_0689_));
 sg13g2_nand2_1 _4282_ (.Y(_0807_),
    .A(_0623_),
    .B(_0806_));
 sg13g2_xor2_1 _4283_ (.B(_0807_),
    .A(_0776_),
    .X(_0808_));
 sg13g2_nand2_1 _4284_ (.Y(_0809_),
    .A(_0624_),
    .B(_0806_));
 sg13g2_xor2_1 _4285_ (.B(_0809_),
    .A(_0779_),
    .X(_0810_));
 sg13g2_nand2_1 _4286_ (.Y(_0811_),
    .A(_0805_),
    .B(_0810_));
 sg13g2_a22oi_1 _4287_ (.Y(_0812_),
    .B1(net905),
    .B2(\dtop.field_top.alt_osc[2] ),
    .A2(net925),
    .A1(\dtop.field_top.comp_values0[3][3] ));
 sg13g2_a22oi_1 _4288_ (.Y(_0813_),
    .B1(net922),
    .B2(\dtop.field_top.comp_values0[4][3] ),
    .A2(net926),
    .A1(\dtop.field_top.comp_values0[2][3] ));
 sg13g2_nand2_1 _4289_ (.Y(_0814_),
    .A(_0812_),
    .B(_0813_));
 sg13g2_a21oi_2 _4290_ (.B1(_0814_),
    .Y(_0815_),
    .A2(net889),
    .A1(_2892_));
 sg13g2_mux2_2 _4291_ (.A0(_0815_),
    .A1(_0037_),
    .S(net891),
    .X(_0816_));
 sg13g2_inv_1 _4292_ (.Y(_0817_),
    .A(_0816_));
 sg13g2_a22oi_1 _4293_ (.Y(_0818_),
    .B1(net905),
    .B2(\dtop.field_top.alt_osc[3] ),
    .A2(net925),
    .A1(\dtop.field_top.comp_values0[3][4] ));
 sg13g2_a22oi_1 _4294_ (.Y(_0819_),
    .B1(net921),
    .B2(\dtop.field_top.comp_values0[4][4] ),
    .A2(net926),
    .A1(\dtop.field_top.comp_values0[2][4] ));
 sg13g2_nand2_1 _4295_ (.Y(_0820_),
    .A(_0818_),
    .B(_0819_));
 sg13g2_a21oi_2 _4296_ (.B1(_0820_),
    .Y(_0821_),
    .A2(net889),
    .A1(_2896_));
 sg13g2_mux2_2 _4297_ (.A0(_0821_),
    .A1(_0036_),
    .S(net892),
    .X(_0822_));
 sg13g2_inv_1 _4298_ (.Y(_0823_),
    .A(_0822_));
 sg13g2_a22oi_1 _4299_ (.Y(_0824_),
    .B1(net922),
    .B2(\dtop.field_top.comp_values0[4][5] ),
    .A2(net924),
    .A1(\dtop.field_top.comp_values0[3][5] ));
 sg13g2_a22oi_1 _4300_ (.Y(_0825_),
    .B1(_0699_),
    .B2(\dtop.field_top.controller.timer[0] ),
    .A2(net927),
    .A1(\dtop.field_top.comp_values0[2][5] ));
 sg13g2_nand2_1 _4301_ (.Y(_0826_),
    .A(_0824_),
    .B(_0825_));
 sg13g2_a221oi_1 _4302_ (.B2(\dtop.field_top.alt_osc[4] ),
    .C1(_0826_),
    .B1(net905),
    .A1(_2902_),
    .Y(_0827_),
    .A2(net889));
 sg13g2_nor2_1 _4303_ (.A(net891),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_a21oi_2 _4304_ (.B1(_0828_),
    .Y(_0829_),
    .A2(net891),
    .A1(_2879_));
 sg13g2_inv_1 _4305_ (.Y(_0830_),
    .A(_0829_));
 sg13g2_a22oi_1 _4306_ (.Y(_0831_),
    .B1(net922),
    .B2(\dtop.field_top.comp_values0[4][6] ),
    .A2(net924),
    .A1(\dtop.field_top.comp_values0[3][6] ));
 sg13g2_a22oi_1 _4307_ (.Y(_0832_),
    .B1(_0699_),
    .B2(\dtop.field_top.controller.timer[1] ),
    .A2(net927),
    .A1(\dtop.field_top.comp_values0[2][6] ));
 sg13g2_nand2_1 _4308_ (.Y(_0833_),
    .A(_0831_),
    .B(_0832_));
 sg13g2_a221oi_1 _4309_ (.B2(\dtop.field_top.alt_osc[5] ),
    .C1(_0833_),
    .B1(net905),
    .A1(_2907_),
    .Y(_0834_),
    .A2(net889));
 sg13g2_nor2_1 _4310_ (.A(net894),
    .B(_0834_),
    .Y(_0835_));
 sg13g2_a21oi_2 _4311_ (.B1(_0835_),
    .Y(_0836_),
    .A2(net894),
    .A1(_2880_));
 sg13g2_inv_1 _4312_ (.Y(_0837_),
    .A(_0836_));
 sg13g2_mux4_1 _4313_ (.S0(net857),
    .A0(_0816_),
    .A1(_0822_),
    .A2(_0829_),
    .A3(_0836_),
    .S1(net854),
    .X(_0838_));
 sg13g2_nor2_1 _4314_ (.A(_0778_),
    .B(_0838_),
    .Y(_0839_));
 sg13g2_a21oi_1 _4315_ (.A1(_0772_),
    .A2(_0778_),
    .Y(_0840_),
    .B1(_0839_));
 sg13g2_nand2_1 _4316_ (.Y(_0841_),
    .A(net852),
    .B(_0840_));
 sg13g2_a21oi_1 _4317_ (.A1(net855),
    .A2(_0778_),
    .Y(_0842_),
    .B1(net852));
 sg13g2_o21ai_1 _4318_ (.B1(_0842_),
    .Y(_0843_),
    .A1(_0739_),
    .A2(_0777_));
 sg13g2_xnor2_1 _4319_ (.Y(_0844_),
    .A(net888),
    .B(_0843_));
 sg13g2_nand3_1 _4320_ (.B(_0841_),
    .C(_0844_),
    .A(_0811_),
    .Y(_0845_));
 sg13g2_xnor2_1 _4321_ (.Y(_0846_),
    .A(net858),
    .B(_0845_));
 sg13g2_and3_1 _4322_ (.X(_0847_),
    .A(_0703_),
    .B(_0704_),
    .C(_0846_));
 sg13g2_a21o_1 _4323_ (.A2(_0834_),
    .A1(net896),
    .B1(_0596_),
    .X(_0848_));
 sg13g2_a21oi_1 _4324_ (.A1(_0034_),
    .A2(net908),
    .Y(_0849_),
    .B1(_0848_));
 sg13g2_mux4_1 _4325_ (.S0(net854),
    .A0(_0741_),
    .A1(_0761_),
    .A2(_0836_),
    .A3(_0749_),
    .S1(_0739_),
    .X(_0850_));
 sg13g2_nand2_1 _4326_ (.Y(_0851_),
    .A(_0777_),
    .B(_0850_));
 sg13g2_mux4_1 _4327_ (.S0(net856),
    .A0(_0771_),
    .A1(_0785_),
    .A2(_0790_),
    .A3(_0796_),
    .S1(net854),
    .X(_0852_));
 sg13g2_o21ai_1 _4328_ (.B1(_0851_),
    .Y(_0853_),
    .A1(_0777_),
    .A2(_0852_));
 sg13g2_mux4_1 _4329_ (.S0(net857),
    .A0(_0802_),
    .A1(_0816_),
    .A2(_0822_),
    .A3(_0829_),
    .S1(net854),
    .X(_0854_));
 sg13g2_mux2_1 _4330_ (.A0(_0850_),
    .A1(_0854_),
    .S(_0780_),
    .X(_0855_));
 sg13g2_xnor2_1 _4331_ (.Y(_0856_),
    .A(net888),
    .B(_0842_));
 sg13g2_a221oi_1 _4332_ (.B2(net852),
    .C1(_0856_),
    .B1(_0855_),
    .A1(net851),
    .Y(_0857_),
    .A2(_0853_));
 sg13g2_xnor2_1 _4333_ (.Y(_0858_),
    .A(_0730_),
    .B(_0857_));
 sg13g2_and2_1 _4334_ (.A(_0849_),
    .B(_0858_),
    .X(_0859_));
 sg13g2_inv_1 _4335_ (.Y(_0860_),
    .A(_0859_));
 sg13g2_a21oi_1 _4336_ (.A1(net895),
    .A2(_0827_),
    .Y(_0861_),
    .B1(net886));
 sg13g2_o21ai_1 _4337_ (.B1(_0861_),
    .Y(_0862_),
    .A1(_2879_),
    .A2(net895));
 sg13g2_mux4_1 _4338_ (.S0(net857),
    .A0(_0830_),
    .A1(_0837_),
    .A2(_0742_),
    .A3(_0748_),
    .S1(net854),
    .X(_0863_));
 sg13g2_mux4_1 _4339_ (.S0(net856),
    .A0(_0760_),
    .A1(_0771_),
    .A2(_0785_),
    .A3(_0790_),
    .S1(net855),
    .X(_0864_));
 sg13g2_mux2_1 _4340_ (.A0(_0863_),
    .A1(_0864_),
    .S(_0781_),
    .X(_0865_));
 sg13g2_nor2_1 _4341_ (.A(net887),
    .B(_0807_),
    .Y(_0866_));
 sg13g2_nand2_1 _4342_ (.Y(_0867_),
    .A(_0594_),
    .B(_0806_));
 sg13g2_a22oi_1 _4343_ (.Y(_0868_),
    .B1(_0750_),
    .B2(_0655_),
    .A2(_0738_),
    .A1(_0732_));
 sg13g2_and2_1 _4344_ (.A(_0781_),
    .B(_0868_),
    .X(_0869_));
 sg13g2_nor2_1 _4345_ (.A(_0605_),
    .B(_0809_),
    .Y(_0870_));
 sg13g2_o21ai_1 _4346_ (.B1(_0865_),
    .Y(_0871_),
    .A1(_0869_),
    .A2(_0870_));
 sg13g2_nand2_1 _4347_ (.Y(_0872_),
    .A(net887),
    .B(net853));
 sg13g2_nor2_1 _4348_ (.A(_0606_),
    .B(net851),
    .Y(_0873_));
 sg13g2_mux4_1 _4349_ (.S0(net856),
    .A0(_0796_),
    .A1(_0803_),
    .A2(_0817_),
    .A3(_0823_),
    .S1(net854),
    .X(_0874_));
 sg13g2_mux2_1 _4350_ (.A0(_0863_),
    .A1(_0874_),
    .S(_0780_),
    .X(_0875_));
 sg13g2_a22oi_1 _4351_ (.Y(_0876_),
    .B1(_0871_),
    .B2(_0872_),
    .A2(_0869_),
    .A1(_0606_));
 sg13g2_o21ai_1 _4352_ (.B1(_0876_),
    .Y(_0877_),
    .A1(net851),
    .A2(_0875_));
 sg13g2_xnor2_1 _4353_ (.Y(_0878_),
    .A(net858),
    .B(_0877_));
 sg13g2_nor2b_1 _4354_ (.A(_0862_),
    .B_N(_0878_),
    .Y(_0879_));
 sg13g2_a21o_1 _4355_ (.A2(_0821_),
    .A1(net895),
    .B1(net886),
    .X(_0880_));
 sg13g2_a21oi_1 _4356_ (.A1(_0036_),
    .A2(net906),
    .Y(_0881_),
    .B1(_0880_));
 sg13g2_mux4_1 _4357_ (.S0(net856),
    .A0(_0822_),
    .A1(_0829_),
    .A2(_0836_),
    .A3(_0741_),
    .S1(net855),
    .X(_0882_));
 sg13g2_nand2_1 _4358_ (.Y(_0883_),
    .A(_0777_),
    .B(_0882_));
 sg13g2_mux4_1 _4359_ (.S0(net856),
    .A0(_0748_),
    .A1(_0760_),
    .A2(_0771_),
    .A3(_0785_),
    .S1(net855),
    .X(_0884_));
 sg13g2_o21ai_1 _4360_ (.B1(_0883_),
    .Y(_0885_),
    .A1(_0777_),
    .A2(_0884_));
 sg13g2_mux4_1 _4361_ (.S0(net856),
    .A0(_0791_),
    .A1(_0797_),
    .A2(_0802_),
    .A3(_0816_),
    .S1(net855),
    .X(_0886_));
 sg13g2_mux2_1 _4362_ (.A0(_0882_),
    .A1(_0886_),
    .S(_0780_),
    .X(_0887_));
 sg13g2_or2_1 _4363_ (.X(_0888_),
    .B(_0887_),
    .A(_0872_));
 sg13g2_o21ai_1 _4364_ (.B1(_0888_),
    .Y(_0889_),
    .A1(_0867_),
    .A2(_0885_));
 sg13g2_xnor2_1 _4365_ (.Y(_0890_),
    .A(net858),
    .B(_0889_));
 sg13g2_nand2b_1 _4366_ (.Y(_0891_),
    .B(_0881_),
    .A_N(_0890_));
 sg13g2_a21o_1 _4367_ (.A2(_0815_),
    .A1(net895),
    .B1(net886),
    .X(_0892_));
 sg13g2_a21oi_1 _4368_ (.A1(_0037_),
    .A2(net906),
    .Y(_0893_),
    .B1(_0892_));
 sg13g2_nor2_1 _4369_ (.A(_0777_),
    .B(_0838_),
    .Y(_0894_));
 sg13g2_a21oi_1 _4370_ (.A1(_0780_),
    .A2(_0804_),
    .Y(_0895_),
    .B1(_0894_));
 sg13g2_nand2_1 _4371_ (.Y(_0896_),
    .A(net851),
    .B(_0840_));
 sg13g2_nand2b_1 _4372_ (.Y(_0897_),
    .B(_0777_),
    .A_N(net855));
 sg13g2_o21ai_1 _4373_ (.B1(net853),
    .Y(_0898_),
    .A1(net856),
    .A2(_0897_));
 sg13g2_xnor2_1 _4374_ (.Y(_0899_),
    .A(net887),
    .B(_0898_));
 sg13g2_a21oi_1 _4375_ (.A1(_0808_),
    .A2(_0895_),
    .Y(_0900_),
    .B1(_0899_));
 sg13g2_nand2_1 _4376_ (.Y(_0901_),
    .A(_0896_),
    .B(_0900_));
 sg13g2_xnor2_1 _4377_ (.Y(_0902_),
    .A(_0731_),
    .B(_0901_));
 sg13g2_and2_1 _4378_ (.A(_0893_),
    .B(_0902_),
    .X(_0903_));
 sg13g2_a21o_1 _4379_ (.A2(_0801_),
    .A1(net895),
    .B1(net886),
    .X(_0904_));
 sg13g2_a21oi_1 _4380_ (.A1(_0048_),
    .A2(net906),
    .Y(_0905_),
    .B1(_0904_));
 sg13g2_nor2b_1 _4381_ (.A(_0855_),
    .B_N(_0866_),
    .Y(_0906_));
 sg13g2_xnor2_1 _4382_ (.Y(_0907_),
    .A(_0594_),
    .B(_0897_));
 sg13g2_nor2b_1 _4383_ (.A(_0907_),
    .B_N(net853),
    .Y(_0908_));
 sg13g2_nor2_1 _4384_ (.A(_0778_),
    .B(_0852_),
    .Y(_0909_));
 sg13g2_and2_1 _4385_ (.A(_0781_),
    .B(_0854_),
    .X(_0910_));
 sg13g2_nor2_1 _4386_ (.A(_0909_),
    .B(_0910_),
    .Y(_0911_));
 sg13g2_o21ai_1 _4387_ (.B1(net852),
    .Y(_0912_),
    .A1(_0909_),
    .A2(_0910_));
 sg13g2_o21ai_1 _4388_ (.B1(_0912_),
    .Y(_0913_),
    .A1(_0906_),
    .A2(_0908_));
 sg13g2_xnor2_1 _4389_ (.Y(_0914_),
    .A(_0731_),
    .B(_0913_));
 sg13g2_nand2_1 _4390_ (.Y(_0915_),
    .A(_0905_),
    .B(_0914_));
 sg13g2_a21oi_1 _4391_ (.A1(net895),
    .A2(_0794_),
    .Y(_0916_),
    .B1(net886));
 sg13g2_o21ai_1 _4392_ (.B1(_0916_),
    .Y(_0917_),
    .A1(_2876_),
    .A2(net895));
 sg13g2_mux2_1 _4393_ (.A0(_0864_),
    .A1(_0874_),
    .S(_0781_),
    .X(_0918_));
 sg13g2_o21ai_1 _4394_ (.B1(_0605_),
    .Y(_0919_),
    .A1(_0781_),
    .A2(_0868_));
 sg13g2_or3_1 _4395_ (.A(_0605_),
    .B(_0781_),
    .C(_0868_),
    .X(_0920_));
 sg13g2_nand2_1 _4396_ (.Y(_0921_),
    .A(_0919_),
    .B(_0920_));
 sg13g2_a21oi_1 _4397_ (.A1(_0919_),
    .A2(_0920_),
    .Y(_0922_),
    .B1(net851));
 sg13g2_a22oi_1 _4398_ (.Y(_0923_),
    .B1(_0918_),
    .B2(_0922_),
    .A2(_0875_),
    .A1(_0866_));
 sg13g2_xnor2_1 _4399_ (.Y(_0924_),
    .A(net858),
    .B(_0923_));
 sg13g2_nor2b_1 _4400_ (.A(_0917_),
    .B_N(_0924_),
    .Y(_0925_));
 sg13g2_or3_1 _4401_ (.A(net887),
    .B(net853),
    .C(_0887_),
    .X(_0926_));
 sg13g2_nand2_1 _4402_ (.Y(_0927_),
    .A(_0778_),
    .B(_0886_));
 sg13g2_o21ai_1 _4403_ (.B1(_0927_),
    .Y(_0928_),
    .A1(_0781_),
    .A2(_0884_));
 sg13g2_nand2_1 _4404_ (.Y(_0929_),
    .A(_0775_),
    .B(net853));
 sg13g2_o21ai_1 _4405_ (.B1(_0926_),
    .Y(_0930_),
    .A1(_0928_),
    .A2(_0929_));
 sg13g2_a21o_1 _4406_ (.A2(_0788_),
    .A1(net896),
    .B1(_0596_),
    .X(_0931_));
 sg13g2_a21oi_1 _4407_ (.A1(_0055_),
    .A2(net908),
    .Y(_0932_),
    .B1(_0931_));
 sg13g2_mux2_2 _4408_ (.A0(net858),
    .A1(_0932_),
    .S(_0930_),
    .X(_0933_));
 sg13g2_xnor2_1 _4409_ (.Y(_0934_),
    .A(_0917_),
    .B(_0924_));
 sg13g2_nand2_1 _4410_ (.Y(_0935_),
    .A(_0933_),
    .B(_0934_));
 sg13g2_a21oi_1 _4411_ (.A1(_0933_),
    .A2(_0934_),
    .Y(_0936_),
    .B1(_0925_));
 sg13g2_xnor2_1 _4412_ (.Y(_0937_),
    .A(_0905_),
    .B(_0914_));
 sg13g2_or2_1 _4413_ (.X(_0938_),
    .B(_0937_),
    .A(_0936_));
 sg13g2_o21ai_1 _4414_ (.B1(_0915_),
    .Y(_0939_),
    .A1(_0936_),
    .A2(_0937_));
 sg13g2_or2_1 _4415_ (.X(_0940_),
    .B(_0902_),
    .A(_0893_));
 sg13g2_nand2b_1 _4416_ (.Y(_0941_),
    .B(_0940_),
    .A_N(_0903_));
 sg13g2_nor2b_1 _4417_ (.A(_0941_),
    .B_N(_0939_),
    .Y(_0942_));
 sg13g2_a21oi_1 _4418_ (.A1(_0939_),
    .A2(_0940_),
    .Y(_0943_),
    .B1(_0903_));
 sg13g2_xor2_1 _4419_ (.B(_0890_),
    .A(_0881_),
    .X(_0944_));
 sg13g2_or2_1 _4420_ (.X(_0945_),
    .B(_0944_),
    .A(_0943_));
 sg13g2_o21ai_1 _4421_ (.B1(_0891_),
    .Y(_0946_),
    .A1(_0943_),
    .A2(_0944_));
 sg13g2_xnor2_1 _4422_ (.Y(_0947_),
    .A(_0862_),
    .B(_0878_));
 sg13g2_a21oi_2 _4423_ (.B1(_0879_),
    .Y(_0948_),
    .A2(_0947_),
    .A1(_0946_));
 sg13g2_nor2_1 _4424_ (.A(_0849_),
    .B(_0858_),
    .Y(_0949_));
 sg13g2_nor2_1 _4425_ (.A(_0859_),
    .B(_0949_),
    .Y(_0950_));
 sg13g2_o21ai_1 _4426_ (.B1(_0860_),
    .Y(_0951_),
    .A1(_0948_),
    .A2(_0949_));
 sg13g2_a21o_1 _4427_ (.A2(_0704_),
    .A1(_0703_),
    .B1(_0846_),
    .X(_0952_));
 sg13g2_nor2b_1 _4428_ (.A(_0847_),
    .B_N(_0952_),
    .Y(_0953_));
 sg13g2_nand2_1 _4429_ (.Y(_0954_),
    .A(_0951_),
    .B(_0953_));
 sg13g2_a21oi_1 _4430_ (.A1(_0951_),
    .A2(_0952_),
    .Y(_0955_),
    .B1(_0847_));
 sg13g2_nand2_1 _4431_ (.Y(_0956_),
    .A(_0032_),
    .B(net908));
 sg13g2_a21oi_1 _4432_ (.A1(net896),
    .A2(_0746_),
    .Y(_0957_),
    .B1(net886));
 sg13g2_nand2_1 _4433_ (.Y(_0958_),
    .A(net851),
    .B(_0928_));
 sg13g2_a21oi_1 _4434_ (.A1(net887),
    .A2(_0622_),
    .Y(_0959_),
    .B1(_0775_));
 sg13g2_a21oi_1 _4435_ (.A1(net853),
    .A2(_0885_),
    .Y(_0960_),
    .B1(_0959_));
 sg13g2_nand3_1 _4436_ (.B(_0958_),
    .C(_0960_),
    .A(_0806_),
    .Y(_0961_));
 sg13g2_xnor2_1 _4437_ (.Y(_0962_),
    .A(net858),
    .B(_0961_));
 sg13g2_a21oi_1 _4438_ (.A1(_0956_),
    .A2(_0957_),
    .Y(_0963_),
    .B1(_0962_));
 sg13g2_nand3_1 _4439_ (.B(_0957_),
    .C(_0962_),
    .A(_0956_),
    .Y(_0964_));
 sg13g2_nor2b_1 _4440_ (.A(_0963_),
    .B_N(_0964_),
    .Y(_0965_));
 sg13g2_xor2_1 _4441_ (.B(_0965_),
    .A(_0955_),
    .X(_0966_));
 sg13g2_or2_1 _4442_ (.X(_0967_),
    .B(_0966_),
    .A(_0677_));
 sg13g2_o21ai_1 _4443_ (.B1(_0696_),
    .Y(_0132_),
    .A1(net878),
    .A2(_0967_));
 sg13g2_o21ai_1 _4444_ (.B1(_0964_),
    .Y(_0968_),
    .A1(_0955_),
    .A2(_0963_));
 sg13g2_a21oi_1 _4445_ (.A1(net896),
    .A2(_0758_),
    .Y(_0969_),
    .B1(net886));
 sg13g2_o21ai_1 _4446_ (.B1(_0969_),
    .Y(_0970_),
    .A1(_2874_),
    .A2(net896));
 sg13g2_nor2_1 _4447_ (.A(net853),
    .B(_0918_),
    .Y(_0971_));
 sg13g2_a22oi_1 _4448_ (.Y(_0972_),
    .B1(_0921_),
    .B2(net851),
    .A2(_0873_),
    .A1(_0865_));
 sg13g2_nor2_1 _4449_ (.A(_0971_),
    .B(_0972_),
    .Y(_0973_));
 sg13g2_xnor2_1 _4450_ (.Y(_0974_),
    .A(_0730_),
    .B(_0973_));
 sg13g2_nor2b_1 _4451_ (.A(_0970_),
    .B_N(_0974_),
    .Y(_0975_));
 sg13g2_xnor2_1 _4452_ (.Y(_0976_),
    .A(_0970_),
    .B(_0974_));
 sg13g2_xnor2_1 _4453_ (.Y(_0977_),
    .A(_0968_),
    .B(_0976_));
 sg13g2_nor2_1 _4454_ (.A(_0677_),
    .B(_0977_),
    .Y(_0978_));
 sg13g2_nor2_1 _4455_ (.A(_0733_),
    .B(_0967_),
    .Y(_0979_));
 sg13g2_a21oi_1 _4456_ (.A1(_0733_),
    .A2(_0978_),
    .Y(_0980_),
    .B1(_0979_));
 sg13g2_nor2_1 _4457_ (.A(net700),
    .B(_0459_),
    .Y(_0981_));
 sg13g2_a21oi_1 _4458_ (.A1(_0459_),
    .A2(_0980_),
    .Y(_0133_),
    .B1(_0981_));
 sg13g2_a21oi_1 _4459_ (.A1(_0968_),
    .A2(_0976_),
    .Y(_0982_),
    .B1(_0975_));
 sg13g2_o21ai_1 _4460_ (.B1(_0595_),
    .Y(_0983_),
    .A1(net908),
    .A2(_0769_));
 sg13g2_a21oi_2 _4461_ (.B1(_0983_),
    .Y(_0984_),
    .A2(net908),
    .A1(_0031_));
 sg13g2_o21ai_1 _4462_ (.B1(_0737_),
    .Y(_0985_),
    .A1(net852),
    .A2(_0911_));
 sg13g2_nor2_1 _4463_ (.A(net852),
    .B(_0907_),
    .Y(_0986_));
 sg13g2_a21oi_1 _4464_ (.A1(net887),
    .A2(net852),
    .Y(_0987_),
    .B1(_0986_));
 sg13g2_a21o_1 _4465_ (.A2(_0853_),
    .A1(net852),
    .B1(_0987_),
    .X(_0988_));
 sg13g2_nor2_1 _4466_ (.A(_0464_),
    .B(_0577_),
    .Y(_0989_));
 sg13g2_nor2_1 _4467_ (.A(_0737_),
    .B(_0989_),
    .Y(_0990_));
 sg13g2_o21ai_1 _4468_ (.B1(_0990_),
    .Y(_0991_),
    .A1(_2913_),
    .A2(net909));
 sg13g2_o21ai_1 _4469_ (.B1(_0991_),
    .Y(_0992_),
    .A1(_0985_),
    .A2(_0988_));
 sg13g2_xnor2_1 _4470_ (.Y(_0993_),
    .A(net858),
    .B(_0992_));
 sg13g2_nand2b_1 _4471_ (.Y(_0994_),
    .B(_0984_),
    .A_N(_0993_));
 sg13g2_xor2_1 _4472_ (.B(_0993_),
    .A(_0984_),
    .X(_0995_));
 sg13g2_xnor2_1 _4473_ (.Y(_0996_),
    .A(_0982_),
    .B(_0995_));
 sg13g2_o21ai_1 _4474_ (.B1(_0733_),
    .Y(_0997_),
    .A1(_0677_),
    .A2(_0996_));
 sg13g2_nand2b_1 _4475_ (.Y(_0998_),
    .B(_0997_),
    .A_N(_0979_));
 sg13g2_o21ai_1 _4476_ (.B1(_0998_),
    .Y(_0999_),
    .A1(_3036_),
    .A2(net966));
 sg13g2_nand4_1 _4477_ (.B(net999),
    .C(net970),
    .A(_3033_),
    .Y(_1000_),
    .D(_0978_));
 sg13g2_and3_1 _4478_ (.X(_1001_),
    .A(_0459_),
    .B(_0999_),
    .C(_1000_));
 sg13g2_a21o_1 _4479_ (.A2(net878),
    .A1(net668),
    .B1(_1001_),
    .X(_0134_));
 sg13g2_o21ai_1 _4480_ (.B1(_0994_),
    .Y(_1002_),
    .A1(_0982_),
    .A2(_0995_));
 sg13g2_nor3_1 _4481_ (.A(_0617_),
    .B(_0636_),
    .C(_0647_),
    .Y(_1003_));
 sg13g2_nand4_1 _4482_ (.B(_0563_),
    .C(_0603_),
    .A(_0447_),
    .Y(_1004_),
    .D(_1003_));
 sg13g2_a21oi_1 _4483_ (.A1(_0446_),
    .A2(_0726_),
    .Y(_1005_),
    .B1(net886));
 sg13g2_nand2_2 _4484_ (.Y(_1006_),
    .A(_1004_),
    .B(_1005_));
 sg13g2_mux2_1 _4485_ (.A0(_0805_),
    .A1(_0895_),
    .S(net851),
    .X(_1007_));
 sg13g2_nand2_1 _4486_ (.Y(_1008_),
    .A(_0739_),
    .B(_0987_));
 sg13g2_nand4_1 _4487_ (.B(_0735_),
    .C(_0737_),
    .A(_0732_),
    .Y(_1009_),
    .D(_1008_));
 sg13g2_nor2_1 _4488_ (.A(_1007_),
    .B(_1009_),
    .Y(_1010_));
 sg13g2_xnor2_1 _4489_ (.Y(_1011_),
    .A(_0730_),
    .B(_1010_));
 sg13g2_nand2b_1 _4490_ (.Y(_1012_),
    .B(_1011_),
    .A_N(_1006_));
 sg13g2_xnor2_1 _4491_ (.Y(_1013_),
    .A(_1006_),
    .B(_1011_));
 sg13g2_nand2_1 _4492_ (.Y(_1014_),
    .A(_1002_),
    .B(_1013_));
 sg13g2_xor2_1 _4493_ (.B(_1013_),
    .A(_1002_),
    .X(_1015_));
 sg13g2_o21ai_1 _4494_ (.B1(_0457_),
    .Y(_1016_),
    .A1(_0053_),
    .A2(net909));
 sg13g2_a21oi_1 _4495_ (.A1(_0455_),
    .A2(_0725_),
    .Y(_1017_),
    .B1(_1016_));
 sg13g2_a22oi_1 _4496_ (.Y(_1018_),
    .B1(_1015_),
    .B2(_0446_),
    .A2(_0727_),
    .A1(net911));
 sg13g2_nand4_1 _4497_ (.B(_3046_),
    .C(_3054_),
    .A(_3036_),
    .Y(_1019_),
    .D(net970));
 sg13g2_nand2_1 _4498_ (.Y(_1020_),
    .A(_3046_),
    .B(net971));
 sg13g2_o21ai_1 _4499_ (.B1(_3110_),
    .Y(_1021_),
    .A1(_0502_),
    .A2(_1019_));
 sg13g2_o21ai_1 _4500_ (.B1(_1021_),
    .Y(_1022_),
    .A1(_0457_),
    .A2(_0728_));
 sg13g2_a21oi_1 _4501_ (.A1(_1017_),
    .A2(_1018_),
    .Y(_1023_),
    .B1(_1022_));
 sg13g2_nand3_1 _4502_ (.B(_3095_),
    .C(_0708_),
    .A(net970),
    .Y(_1024_));
 sg13g2_nand3_1 _4503_ (.B(_0709_),
    .C(_1024_),
    .A(net909),
    .Y(_1025_));
 sg13g2_xor2_1 _4504_ (.B(_1025_),
    .A(_1023_),
    .X(_1026_));
 sg13g2_nand2_1 _4505_ (.Y(_1027_),
    .A(net642),
    .B(net878));
 sg13g2_o21ai_1 _4506_ (.B1(_1027_),
    .Y(_0135_),
    .A1(net878),
    .A2(_1026_));
 sg13g2_a21oi_2 _4507_ (.B1(net930),
    .Y(_1028_),
    .A2(_2993_),
    .A1(_2947_));
 sg13g2_nand2_1 _4508_ (.Y(_1029_),
    .A(net451),
    .B(net904));
 sg13g2_nand2_1 _4509_ (.Y(_1030_),
    .A(_0109_),
    .B(net957));
 sg13g2_a21oi_1 _4510_ (.A1(_0109_),
    .A2(_2947_),
    .Y(_1031_),
    .B1(net1034));
 sg13g2_nand2b_1 _4511_ (.Y(_1032_),
    .B(_1030_),
    .A_N(net1034));
 sg13g2_o21ai_1 _4512_ (.B1(_1030_),
    .Y(_1033_),
    .A1(_2869_),
    .A2(net957));
 sg13g2_mux2_1 _4513_ (.A0(_0018_),
    .A1(_0016_),
    .S(net958),
    .X(_1034_));
 sg13g2_nand2b_1 _4514_ (.Y(_1035_),
    .B(_1033_),
    .A_N(_1034_));
 sg13g2_o21ai_1 _4515_ (.B1(_0009_),
    .Y(_1036_),
    .A1(_0014_),
    .A2(_2948_));
 sg13g2_mux2_2 _4516_ (.A0(_0019_),
    .A1(_0015_),
    .S(net957),
    .X(_1037_));
 sg13g2_nor2b_1 _4517_ (.A(_1037_),
    .B_N(_1036_),
    .Y(_1038_));
 sg13g2_nand2b_1 _4518_ (.Y(_1039_),
    .B(_1038_),
    .A_N(_1035_));
 sg13g2_nand2b_1 _4519_ (.Y(_1040_),
    .B(_1034_),
    .A_N(_1033_));
 sg13g2_nor2b_1 _4520_ (.A(_1036_),
    .B_N(_1037_),
    .Y(_1041_));
 sg13g2_nor2b_1 _4521_ (.A(_1040_),
    .B_N(_1041_),
    .Y(_1042_));
 sg13g2_nor2_1 _4522_ (.A(net948),
    .B(_1042_),
    .Y(_1043_));
 sg13g2_a21oi_1 _4523_ (.A1(net948),
    .A2(_1039_),
    .Y(_1044_),
    .B1(_1043_));
 sg13g2_and2_1 _4524_ (.A(_1036_),
    .B(_1037_),
    .X(_1045_));
 sg13g2_nor2_1 _4525_ (.A(net948),
    .B(_1040_),
    .Y(_1046_));
 sg13g2_nor2_2 _4526_ (.A(_1036_),
    .B(_1037_),
    .Y(_1047_));
 sg13g2_nor2b_1 _4527_ (.A(_1035_),
    .B_N(_1047_),
    .Y(_1048_));
 sg13g2_a221oi_1 _4528_ (.B2(net948),
    .C1(_1044_),
    .B1(_1048_),
    .A1(_1045_),
    .Y(_1049_),
    .A2(_1046_));
 sg13g2_nor2b_1 _4529_ (.A(net956),
    .B_N(_0070_),
    .Y(_1050_));
 sg13g2_a21oi_1 _4530_ (.A1(_0071_),
    .A2(net956),
    .Y(_1051_),
    .B1(_1050_));
 sg13g2_nand2_1 _4531_ (.Y(_1052_),
    .A(_1049_),
    .B(_1051_));
 sg13g2_nor3_1 _4532_ (.A(_1032_),
    .B(_1033_),
    .C(_1034_),
    .Y(_1053_));
 sg13g2_and3_1 _4533_ (.X(_1054_),
    .A(_1032_),
    .B(_1033_),
    .C(_1034_));
 sg13g2_a22oi_1 _4534_ (.Y(_1055_),
    .B1(_1054_),
    .B2(_1047_),
    .A2(_1053_),
    .A1(_1045_));
 sg13g2_nor2_1 _4535_ (.A(_1032_),
    .B(_1040_),
    .Y(_1056_));
 sg13g2_nor2_1 _4536_ (.A(_1031_),
    .B(_1035_),
    .Y(_1057_));
 sg13g2_a22oi_1 _4537_ (.Y(_1058_),
    .B1(_1057_),
    .B2(_1041_),
    .A2(_1056_),
    .A1(_1038_));
 sg13g2_and2_1 _4538_ (.A(_1055_),
    .B(_1058_),
    .X(_1059_));
 sg13g2_a22oi_1 _4539_ (.Y(_1060_),
    .B1(_1057_),
    .B2(_1047_),
    .A2(_1056_),
    .A1(_1045_));
 sg13g2_nor2_1 _4540_ (.A(net948),
    .B(_1039_),
    .Y(_1061_));
 sg13g2_a21oi_1 _4541_ (.A1(net948),
    .A2(_1042_),
    .Y(_1062_),
    .B1(_1061_));
 sg13g2_a22oi_1 _4542_ (.Y(_1063_),
    .B1(_1047_),
    .B2(net948),
    .A2(_1045_),
    .A1(_1033_));
 sg13g2_a21oi_2 _4543_ (.B1(_1063_),
    .Y(_1064_),
    .A2(_1033_),
    .A1(net948));
 sg13g2_a22oi_1 _4544_ (.Y(_1065_),
    .B1(_1054_),
    .B2(_1038_),
    .A2(_1053_),
    .A1(_1041_));
 sg13g2_and2_1 _4545_ (.A(_1049_),
    .B(_1065_),
    .X(_1066_));
 sg13g2_nand2b_1 _4546_ (.Y(_1067_),
    .B(_1066_),
    .A_N(_1064_));
 sg13g2_inv_1 _4547_ (.Y(_1068_),
    .A(_1067_));
 sg13g2_nand4_1 _4548_ (.B(_1060_),
    .C(_1062_),
    .A(_1059_),
    .Y(_1069_),
    .D(_1068_));
 sg13g2_nand3_1 _4549_ (.B(_1040_),
    .C(_1064_),
    .A(_1035_),
    .Y(_1070_));
 sg13g2_nand4_1 _4550_ (.B(_1066_),
    .C(_1069_),
    .A(_1059_),
    .Y(_1071_),
    .D(_1070_));
 sg13g2_mux2_1 _4551_ (.A0(_0064_),
    .A1(_0065_),
    .S(net956),
    .X(_1072_));
 sg13g2_nor2b_1 _4552_ (.A(_1072_),
    .B_N(_1071_),
    .Y(_1073_));
 sg13g2_nor2_1 _4553_ (.A(_1044_),
    .B(_1064_),
    .Y(_1074_));
 sg13g2_nand2_1 _4554_ (.Y(_1075_),
    .A(_1065_),
    .B(_1074_));
 sg13g2_nor2b_1 _4555_ (.A(net957),
    .B_N(_0068_),
    .Y(_1076_));
 sg13g2_a21oi_1 _4556_ (.A1(_0069_),
    .A2(net957),
    .Y(_1077_),
    .B1(_1076_));
 sg13g2_nand4_1 _4557_ (.B(_1060_),
    .C(_1062_),
    .A(_1059_),
    .Y(_1078_),
    .D(_1077_));
 sg13g2_a221oi_1 _4558_ (.B2(_1078_),
    .C1(_0008_),
    .B1(_1075_),
    .A1(_0012_),
    .Y(_1079_),
    .A2(net957));
 sg13g2_nand2b_1 _4559_ (.Y(_1080_),
    .B(_1062_),
    .A_N(_1064_));
 sg13g2_o21ai_1 _4560_ (.B1(net1054),
    .Y(_1081_),
    .A1(\dtop.field_top.alt_osc[3] ),
    .A2(_2948_));
 sg13g2_or2_1 _4561_ (.X(_1082_),
    .B(_1081_),
    .A(_1080_));
 sg13g2_o21ai_1 _4562_ (.B1(_1082_),
    .Y(_1083_),
    .A1(_1075_),
    .A2(_1078_));
 sg13g2_nand2_1 _4563_ (.Y(_1084_),
    .A(_1059_),
    .B(_1074_));
 sg13g2_mux2_1 _4564_ (.A0(_0067_),
    .A1(_0011_),
    .S(net957),
    .X(_1085_));
 sg13g2_a22oi_1 _4565_ (.Y(_1086_),
    .B1(_1084_),
    .B2(_1085_),
    .A2(_1081_),
    .A1(_1080_));
 sg13g2_o21ai_1 _4566_ (.B1(_1086_),
    .Y(_1087_),
    .A1(_1079_),
    .A2(_1083_));
 sg13g2_nor2_1 _4567_ (.A(_0066_),
    .B(net958),
    .Y(_1088_));
 sg13g2_nor2_1 _4568_ (.A(net683),
    .B(_2971_),
    .Y(_1089_));
 sg13g2_and3_1 _4569_ (.X(_1090_),
    .A(_1055_),
    .B(_1060_),
    .C(_1068_));
 sg13g2_o21ai_1 _4570_ (.B1(_1090_),
    .Y(_1091_),
    .A1(_1088_),
    .A2(_1089_));
 sg13g2_o21ai_1 _4571_ (.B1(_1087_),
    .Y(_1092_),
    .A1(_1084_),
    .A2(_1085_));
 sg13g2_nand2b_1 _4572_ (.Y(_1093_),
    .B(_1091_),
    .A_N(_1092_));
 sg13g2_or3_1 _4573_ (.A(_1088_),
    .B(_1089_),
    .C(_1090_),
    .X(_1094_));
 sg13g2_and2_1 _4574_ (.A(_1069_),
    .B(_1094_),
    .X(_1095_));
 sg13g2_xor2_1 _4575_ (.B(_1072_),
    .A(_1071_),
    .X(_1096_));
 sg13g2_a21oi_1 _4576_ (.A1(_1093_),
    .A2(_1095_),
    .Y(_1097_),
    .B1(_1096_));
 sg13g2_xor2_1 _4577_ (.B(_1051_),
    .A(_1049_),
    .X(_1098_));
 sg13g2_o21ai_1 _4578_ (.B1(_1098_),
    .Y(_1099_),
    .A1(_1073_),
    .A2(_1097_));
 sg13g2_nand2_1 _4579_ (.Y(_1100_),
    .A(_1052_),
    .B(_1099_));
 sg13g2_nor2b_1 _4580_ (.A(net956),
    .B_N(_0072_),
    .Y(_1101_));
 sg13g2_a21oi_1 _4581_ (.A1(_0073_),
    .A2(net956),
    .Y(_1102_),
    .B1(_1101_));
 sg13g2_and2_1 _4582_ (.A(_1100_),
    .B(_1102_),
    .X(_1103_));
 sg13g2_nor2b_1 _4583_ (.A(net953),
    .B_N(_0074_),
    .Y(_1104_));
 sg13g2_a21oi_1 _4584_ (.A1(_0026_),
    .A2(net953),
    .Y(_1105_),
    .B1(_1104_));
 sg13g2_and2_1 _4585_ (.A(_1103_),
    .B(_1105_),
    .X(_1106_));
 sg13g2_nor2b_1 _4586_ (.A(net953),
    .B_N(_0025_),
    .Y(_1107_));
 sg13g2_a21oi_1 _4587_ (.A1(_0099_),
    .A2(net953),
    .Y(_1108_),
    .B1(_1107_));
 sg13g2_and2_1 _4588_ (.A(_1106_),
    .B(_1108_),
    .X(_1109_));
 sg13g2_nor2b_1 _4589_ (.A(net955),
    .B_N(_0096_),
    .Y(_1110_));
 sg13g2_a21oi_2 _4590_ (.B1(_1110_),
    .Y(_1111_),
    .A2(net955),
    .A1(_0098_));
 sg13g2_nand2_1 _4591_ (.Y(_1112_),
    .A(_1109_),
    .B(_1111_));
 sg13g2_nor2b_1 _4592_ (.A(net954),
    .B_N(_0094_),
    .Y(_1113_));
 sg13g2_a21oi_1 _4593_ (.A1(_0093_),
    .A2(net954),
    .Y(_1114_),
    .B1(_1113_));
 sg13g2_nand3_1 _4594_ (.B(_1111_),
    .C(_1114_),
    .A(_1109_),
    .Y(_1115_));
 sg13g2_mux2_1 _4595_ (.A0(_0091_),
    .A1(_0106_),
    .S(net954),
    .X(_1116_));
 sg13g2_or2_1 _4596_ (.X(_1117_),
    .B(_1116_),
    .A(_1115_));
 sg13g2_mux2_1 _4597_ (.A0(_0103_),
    .A1(_0104_),
    .S(net953),
    .X(_1118_));
 sg13g2_mux2_1 _4598_ (.A0(_0101_),
    .A1(_0024_),
    .S(net953),
    .X(_1119_));
 sg13g2_nor3_1 _4599_ (.A(_1117_),
    .B(_1118_),
    .C(_1119_),
    .Y(_1120_));
 sg13g2_o21ai_1 _4600_ (.B1(_1119_),
    .Y(_1121_),
    .A1(_1117_),
    .A2(_1118_));
 sg13g2_nand2b_1 _4601_ (.Y(_1122_),
    .B(_1121_),
    .A_N(_1120_));
 sg13g2_o21ai_1 _4602_ (.B1(_1029_),
    .Y(_0136_),
    .A1(net913),
    .A2(_1122_));
 sg13g2_nand2_1 _4603_ (.Y(_1123_),
    .A(net398),
    .B(net904));
 sg13g2_mux2_1 _4604_ (.A0(net355),
    .A1(\dtop.field_top.fy[10] ),
    .S(net953),
    .X(_1124_));
 sg13g2_xnor2_1 _4605_ (.Y(_1125_),
    .A(_1120_),
    .B(_1124_));
 sg13g2_o21ai_1 _4606_ (.B1(_1123_),
    .Y(_0137_),
    .A1(net913),
    .A2(_1125_));
 sg13g2_a22oi_1 _4607_ (.Y(_1126_),
    .B1(_1028_),
    .B2(\dtop.field_top.fy[0] ),
    .A2(net930),
    .A1(net570));
 sg13g2_nand3_1 _4608_ (.B(_1095_),
    .C(_1096_),
    .A(_1093_),
    .Y(_1127_));
 sg13g2_nor2b_1 _4609_ (.A(_1097_),
    .B_N(_1127_),
    .Y(_1128_));
 sg13g2_inv_1 _4610_ (.Y(_1129_),
    .A(_1128_));
 sg13g2_o21ai_1 _4611_ (.B1(net571),
    .Y(_0138_),
    .A1(net914),
    .A2(_1129_));
 sg13g2_a22oi_1 _4612_ (.Y(_1130_),
    .B1(_1028_),
    .B2(\dtop.field_top.fy[1] ),
    .A2(net930),
    .A1(net305));
 sg13g2_or3_1 _4613_ (.A(_1073_),
    .B(_1097_),
    .C(_1098_),
    .X(_1131_));
 sg13g2_nand2_1 _4614_ (.Y(_1132_),
    .A(_1099_),
    .B(_1131_));
 sg13g2_o21ai_1 _4615_ (.B1(net306),
    .Y(_0139_),
    .A1(net913),
    .A2(_1132_));
 sg13g2_a22oi_1 _4616_ (.Y(_1133_),
    .B1(_1028_),
    .B2(\dtop.field_top.fy[2] ),
    .A2(net929),
    .A1(net322));
 sg13g2_xor2_1 _4617_ (.B(_1102_),
    .A(_1100_),
    .X(_1134_));
 sg13g2_inv_1 _4618_ (.Y(_1135_),
    .A(_1134_));
 sg13g2_o21ai_1 _4619_ (.B1(net323),
    .Y(_0140_),
    .A1(net914),
    .A2(_1135_));
 sg13g2_a22oi_1 _4620_ (.Y(_1136_),
    .B1(net904),
    .B2(\dtop.field_top.fy[3] ),
    .A2(net929),
    .A1(net353));
 sg13g2_xnor2_1 _4621_ (.Y(_1137_),
    .A(_1103_),
    .B(_1105_));
 sg13g2_o21ai_1 _4622_ (.B1(net354),
    .Y(_0141_),
    .A1(net914),
    .A2(_1137_));
 sg13g2_a22oi_1 _4623_ (.Y(_1138_),
    .B1(net904),
    .B2(net362),
    .A2(net928),
    .A1(_0021_));
 sg13g2_xnor2_1 _4624_ (.Y(_1139_),
    .A(_1106_),
    .B(_1108_));
 sg13g2_o21ai_1 _4625_ (.B1(net363),
    .Y(_0142_),
    .A1(net913),
    .A2(_1139_));
 sg13g2_a22oi_1 _4626_ (.Y(_1140_),
    .B1(net904),
    .B2(net412),
    .A2(net928),
    .A1(_0020_));
 sg13g2_xnor2_1 _4627_ (.Y(_1141_),
    .A(_1109_),
    .B(_1111_));
 sg13g2_o21ai_1 _4628_ (.B1(net413),
    .Y(_0143_),
    .A1(net913),
    .A2(_1141_));
 sg13g2_a22oi_1 _4629_ (.Y(_1142_),
    .B1(net904),
    .B2(\dtop.field_top.fy[6] ),
    .A2(net928),
    .A1(net314));
 sg13g2_xor2_1 _4630_ (.B(_1114_),
    .A(_1112_),
    .X(_1143_));
 sg13g2_o21ai_1 _4631_ (.B1(net315),
    .Y(_0144_),
    .A1(net913),
    .A2(_1143_));
 sg13g2_a22oi_1 _4632_ (.Y(_1144_),
    .B1(net904),
    .B2(\dtop.field_top.fy[7] ),
    .A2(net928),
    .A1(net307));
 sg13g2_xnor2_1 _4633_ (.Y(_1145_),
    .A(_1115_),
    .B(_1116_));
 sg13g2_o21ai_1 _4634_ (.B1(net308),
    .Y(_0145_),
    .A1(net913),
    .A2(_1145_));
 sg13g2_a22oi_1 _4635_ (.Y(_1146_),
    .B1(net904),
    .B2(net350),
    .A2(net928),
    .A1(_0079_));
 sg13g2_xnor2_1 _4636_ (.Y(_1147_),
    .A(_1117_),
    .B(_1118_));
 sg13g2_o21ai_1 _4637_ (.B1(net351),
    .Y(_0146_),
    .A1(net913),
    .A2(_1147_));
 sg13g2_nor2_2 _4638_ (.A(net304),
    .B(_2929_),
    .Y(_1148_));
 sg13g2_inv_2 _4639_ (.Y(_1149_),
    .A(_1148_));
 sg13g2_nor2_2 _4640_ (.A(_2947_),
    .B(_1148_),
    .Y(_1150_));
 sg13g2_a22oi_1 _4641_ (.Y(_1151_),
    .B1(_1150_),
    .B2(net487),
    .A2(net956),
    .A1(net477));
 sg13g2_o21ai_1 _4642_ (.B1(_1151_),
    .Y(_0147_),
    .A1(_1129_),
    .A2(_1149_));
 sg13g2_a22oi_1 _4643_ (.Y(_1152_),
    .B1(net947),
    .B2(net463),
    .A2(net956),
    .A1(\dtop.field_top.controller.timer[2] ));
 sg13g2_o21ai_1 _4644_ (.B1(net464),
    .Y(_0148_),
    .A1(_1132_),
    .A2(_1149_));
 sg13g2_a22oi_1 _4645_ (.Y(_1153_),
    .B1(_1150_),
    .B2(net613),
    .A2(net958),
    .A1(\dtop.field_top.controller.ppos[0] ));
 sg13g2_o21ai_1 _4646_ (.B1(net614),
    .Y(_0149_),
    .A1(_1135_),
    .A2(net979));
 sg13g2_a22oi_1 _4647_ (.Y(_1154_),
    .B1(_1150_),
    .B2(net497),
    .A2(net953),
    .A1(\dtop.field_top.controller.ppos[1] ));
 sg13g2_o21ai_1 _4648_ (.B1(net498),
    .Y(_0150_),
    .A1(_1137_),
    .A2(_1149_));
 sg13g2_a22oi_1 _4649_ (.Y(_1155_),
    .B1(net947),
    .B2(net484),
    .A2(net955),
    .A1(\dtop.field_top.controller.ppos[2] ));
 sg13g2_o21ai_1 _4650_ (.B1(net485),
    .Y(_0151_),
    .A1(_1139_),
    .A2(net979));
 sg13g2_a22oi_1 _4651_ (.Y(_1156_),
    .B1(net947),
    .B2(net379),
    .A2(net954),
    .A1(\dtop.field_top.controller.ppos[3] ));
 sg13g2_o21ai_1 _4652_ (.B1(net380),
    .Y(_0152_),
    .A1(_1141_),
    .A2(net979));
 sg13g2_a22oi_1 _4653_ (.Y(_1157_),
    .B1(net947),
    .B2(net407),
    .A2(net954),
    .A1(\dtop.field_top.controller.ppos[4] ));
 sg13g2_o21ai_1 _4654_ (.B1(net408),
    .Y(_0153_),
    .A1(_1143_),
    .A2(net979));
 sg13g2_a22oi_1 _4655_ (.Y(_1158_),
    .B1(net947),
    .B2(net377),
    .A2(net954),
    .A1(net1033));
 sg13g2_o21ai_1 _4656_ (.B1(_1158_),
    .Y(_0154_),
    .A1(_1145_),
    .A2(net979));
 sg13g2_a22oi_1 _4657_ (.Y(_1159_),
    .B1(net947),
    .B2(net511),
    .A2(net954),
    .A1(net1032));
 sg13g2_o21ai_1 _4658_ (.B1(net512),
    .Y(_0155_),
    .A1(_1147_),
    .A2(net979));
 sg13g2_a22oi_1 _4659_ (.Y(_1160_),
    .B1(net947),
    .B2(net369),
    .A2(net954),
    .A1(\dtop.field_top.controller.pattern0[0] ));
 sg13g2_o21ai_1 _4660_ (.B1(net370),
    .Y(_0156_),
    .A1(_1122_),
    .A2(net979));
 sg13g2_nor2b_1 _4661_ (.A(_2929_),
    .B_N(_2993_),
    .Y(_1161_));
 sg13g2_nand2b_1 _4662_ (.Y(_1162_),
    .B(_2993_),
    .A_N(net630));
 sg13g2_nand2b_1 _4663_ (.Y(_1163_),
    .B(net1057),
    .A_N(\dtop.field_top.alt_osc[2] ));
 sg13g2_and3_1 _4664_ (.X(_1164_),
    .A(net1008),
    .B(\dtop.field_top.alt_osc[1] ),
    .C(_1163_));
 sg13g2_a221oi_1 _4665_ (.B2(net1006),
    .C1(_1164_),
    .B1(\dtop.field_top.alt_osc[3] ),
    .A1(net1007),
    .Y(_1165_),
    .A2(\dtop.field_top.alt_osc[2] ));
 sg13g2_nand2b_1 _4666_ (.Y(_1166_),
    .B(net1050),
    .A_N(\dtop.field_top.alt_osc[4] ));
 sg13g2_o21ai_1 _4667_ (.B1(_1166_),
    .Y(_1167_),
    .A1(net1006),
    .A2(\dtop.field_top.alt_osc[3] ));
 sg13g2_a22oi_1 _4668_ (.Y(_1168_),
    .B1(\dtop.field_top.alt_osc[5] ),
    .B2(net1015),
    .A2(\dtop.field_top.alt_osc[4] ),
    .A1(net1004));
 sg13g2_o21ai_1 _4669_ (.B1(_1168_),
    .Y(_1169_),
    .A1(_1165_),
    .A2(_1167_));
 sg13g2_o21ai_1 _4670_ (.B1(_1169_),
    .Y(_1170_),
    .A1(net1015),
    .A2(\dtop.field_top.alt_osc[5] ));
 sg13g2_inv_1 _4671_ (.Y(_1171_),
    .A(_1170_));
 sg13g2_nor2_1 _4672_ (.A(_0014_),
    .B(_1170_),
    .Y(_1172_));
 sg13g2_o21ai_1 _4673_ (.B1(_0015_),
    .Y(_1173_),
    .A1(_0014_),
    .A2(_1170_));
 sg13g2_nor2_1 _4674_ (.A(\dtop.field_top.alt_osc[6] ),
    .B(\dtop.field_top.alt_osc[7] ),
    .Y(_1174_));
 sg13g2_a21oi_1 _4675_ (.A1(_2868_),
    .A2(_1174_),
    .Y(_1175_),
    .B1(_3047_));
 sg13g2_o21ai_1 _4676_ (.B1(_1175_),
    .Y(_1176_),
    .A1(_2868_),
    .A2(_1173_));
 sg13g2_nand2_1 _4677_ (.Y(_1177_),
    .A(net1046),
    .B(_1173_));
 sg13g2_nor2b_1 _4678_ (.A(\dtop.field_top.alt_osc[7] ),
    .B_N(_0014_),
    .Y(_1178_));
 sg13g2_nor2_1 _4679_ (.A(net1045),
    .B(_1178_),
    .Y(_1179_));
 sg13g2_nand2_1 _4680_ (.Y(_1180_),
    .A(\dtop.field_top.alt_osc[7] ),
    .B(_1171_));
 sg13g2_o21ai_1 _4681_ (.B1(_1179_),
    .Y(_1181_),
    .A1(\dtop.field_top.alt_osc[6] ),
    .A2(_1180_));
 sg13g2_nand2_1 _4682_ (.Y(_1182_),
    .A(_1177_),
    .B(_1181_));
 sg13g2_nand3_1 _4683_ (.B(_0016_),
    .C(_1182_),
    .A(net1014),
    .Y(_1183_));
 sg13g2_a21oi_1 _4684_ (.A1(_1176_),
    .A2(_1183_),
    .Y(_1184_),
    .B1(_0109_));
 sg13g2_nand2_1 _4685_ (.Y(_1185_),
    .A(net1013),
    .B(net1060));
 sg13g2_nand3_1 _4686_ (.B(_1170_),
    .C(_1185_),
    .A(\dtop.field_top.alt_osc[6] ),
    .Y(_1186_));
 sg13g2_a21oi_1 _4687_ (.A1(net1044),
    .A2(_2868_),
    .Y(_1187_),
    .B1(_1174_));
 sg13g2_nand3_1 _4688_ (.B(_1186_),
    .C(_1187_),
    .A(net1045),
    .Y(_1188_));
 sg13g2_nand2_1 _4689_ (.Y(_1189_),
    .A(net1042),
    .B(_0016_));
 sg13g2_nand4_1 _4690_ (.B(_1180_),
    .C(_1185_),
    .A(_1179_),
    .Y(_1190_),
    .D(_1189_));
 sg13g2_nand2_1 _4691_ (.Y(_1191_),
    .A(_1188_),
    .B(_1190_));
 sg13g2_nor2_1 _4692_ (.A(net1013),
    .B(_1177_),
    .Y(_1192_));
 sg13g2_a21oi_1 _4693_ (.A1(\dtop.field_top.rs.scan_y.pos[8] ),
    .A2(net1060),
    .Y(_1193_),
    .B1(_2953_));
 sg13g2_a221oi_1 _4694_ (.B2(_1193_),
    .C1(_2844_),
    .B1(_1192_),
    .A1(\dtop.field_top.rs.scan_y.pos[8] ),
    .Y(_1194_),
    .A2(_1191_));
 sg13g2_o21ai_1 _4695_ (.B1(net1039),
    .Y(_1195_),
    .A1(net1041),
    .A2(_1184_));
 sg13g2_a21o_1 _4696_ (.A2(_1172_),
    .A1(\dtop.field_top.alt_osc[7] ),
    .B1(_1178_),
    .X(_1196_));
 sg13g2_nor4_1 _4697_ (.A(_0109_),
    .B(net1060),
    .C(_3026_),
    .D(_1196_),
    .Y(_1197_));
 sg13g2_nor2_1 _4698_ (.A(_2843_),
    .B(_1197_),
    .Y(_1198_));
 sg13g2_o21ai_1 _4699_ (.B1(_1198_),
    .Y(_1199_),
    .A1(_1194_),
    .A2(_1195_));
 sg13g2_nor3_1 _4700_ (.A(net1042),
    .B(_0009_),
    .C(_1196_),
    .Y(_1200_));
 sg13g2_a21oi_1 _4701_ (.A1(net1042),
    .A2(_1182_),
    .Y(_1201_),
    .B1(_1200_));
 sg13g2_nand2_1 _4702_ (.Y(_1202_),
    .A(_2844_),
    .B(_1201_));
 sg13g2_xnor2_1 _4703_ (.Y(_1203_),
    .A(\dtop.field_top.alt_osc[7] ),
    .B(_1172_));
 sg13g2_nor3_1 _4704_ (.A(net1042),
    .B(_0009_),
    .C(_1174_),
    .Y(_1204_));
 sg13g2_nor3_1 _4705_ (.A(net1018),
    .B(_1192_),
    .C(_1204_),
    .Y(_1205_));
 sg13g2_o21ai_1 _4706_ (.B1(_1205_),
    .Y(_1206_),
    .A1(_3039_),
    .A2(_1203_));
 sg13g2_nand3_1 _4707_ (.B(_1202_),
    .C(_1206_),
    .A(net532),
    .Y(_1207_));
 sg13g2_nor2b_1 _4708_ (.A(\dtop.field_top.controller.ppos[4] ),
    .B_N(_0005_),
    .Y(_1208_));
 sg13g2_nand2_2 _4709_ (.Y(_1209_),
    .A(\dtop.field_top.controller.ppos[5] ),
    .B(\dtop.field_top.controller.ppos[6] ));
 sg13g2_nand3_1 _4710_ (.B(net1031),
    .C(_0108_),
    .A(\dtop.field_top.controller.pattern0[0] ),
    .Y(_1210_));
 sg13g2_and2_1 _4711_ (.A(net1031),
    .B(_1210_),
    .X(_1211_));
 sg13g2_nor2_2 _4712_ (.A(net1030),
    .B(_3061_),
    .Y(_1212_));
 sg13g2_nand3b_1 _4713_ (.B(\dtop.field_top.controller.pattern0[0] ),
    .C(net1031),
    .Y(_1213_),
    .A_N(\dtop.field_top.controller.pattern0[2] ));
 sg13g2_o21ai_1 _4714_ (.B1(_1211_),
    .Y(_1214_),
    .A1(_3063_),
    .A2(_1212_));
 sg13g2_xnor2_1 _4715_ (.Y(_1215_),
    .A(_0004_),
    .B(_1214_));
 sg13g2_mux4_1 _4716_ (.S0(net1033),
    .A0(_1208_),
    .A1(_0399_),
    .A2(_0398_),
    .A3(_1215_),
    .S1(net1032),
    .X(_1216_));
 sg13g2_mux4_1 _4717_ (.S0(net1033),
    .A0(_2871_),
    .A1(_0397_),
    .A2(_0396_),
    .A3(_0395_),
    .S1(net1032),
    .X(_1217_));
 sg13g2_and2_1 _4718_ (.A(\dtop.field_top.rs.scan_y.pos[8] ),
    .B(_1217_),
    .X(_1218_));
 sg13g2_nor4_1 _4719_ (.A(_2868_),
    .B(_0016_),
    .C(_1216_),
    .D(_1218_),
    .Y(_1219_));
 sg13g2_nand2_1 _4720_ (.Y(_1220_),
    .A(net1060),
    .B(\dtop.field_top.controller.ppos[0] ));
 sg13g2_a21oi_1 _4721_ (.A1(_1217_),
    .A2(_1220_),
    .Y(_1221_),
    .B1(\dtop.field_top.rs.scan_y.pos[8] ));
 sg13g2_nand2_1 _4722_ (.Y(_1222_),
    .A(\dtop.field_top.controller.pattern0[0] ),
    .B(_2850_));
 sg13g2_xnor2_1 _4723_ (.Y(_1223_),
    .A(\dtop.field_top.controller.pattern0[0] ),
    .B(\dtop.field_top.controller.pattern0[1] ));
 sg13g2_nor4_2 _4724_ (.A(\dtop.field_top.controller.ppos[4] ),
    .B(net1033),
    .C(net1032),
    .Y(_1224_),
    .D(_0006_));
 sg13g2_a221oi_1 _4725_ (.B2(net1030),
    .C1(_1224_),
    .B1(_1223_),
    .A1(_0108_),
    .Y(_1225_),
    .A2(_1222_));
 sg13g2_a21oi_1 _4726_ (.A1(_0395_),
    .A2(_1215_),
    .Y(_1226_),
    .B1(_1209_));
 sg13g2_nor2b_1 _4727_ (.A(net1033),
    .B_N(_0400_),
    .Y(_1227_));
 sg13g2_a21oi_1 _4728_ (.A1(net1033),
    .A2(_2870_),
    .Y(_1228_),
    .B1(net1032));
 sg13g2_or3_2 _4729_ (.A(_1226_),
    .B(_1227_),
    .C(_1228_),
    .X(_1229_));
 sg13g2_nor2_1 _4730_ (.A(_1219_),
    .B(_1221_),
    .Y(_1230_));
 sg13g2_nand4_1 _4731_ (.B(_1225_),
    .C(_1229_),
    .A(_1199_),
    .Y(_1231_),
    .D(_1230_));
 sg13g2_a21oi_2 _4732_ (.B1(_1231_),
    .Y(_1232_),
    .A2(_1207_),
    .A1(_2843_));
 sg13g2_nor2_1 _4733_ (.A(_1162_),
    .B(_1232_),
    .Y(_1233_));
 sg13g2_nand2b_1 _4734_ (.Y(_1234_),
    .B(_3066_),
    .A_N(\dtop.field_top.rside ));
 sg13g2_nand2_1 _4735_ (.Y(_1235_),
    .A(net1031),
    .B(_3063_));
 sg13g2_nand3_1 _4736_ (.B(_3063_),
    .C(_1209_),
    .A(net1031),
    .Y(_1236_));
 sg13g2_nor2_1 _4737_ (.A(net1030),
    .B(net1031),
    .Y(_1237_));
 sg13g2_o21ai_1 _4738_ (.B1(_1210_),
    .Y(_1238_),
    .A1(net1030),
    .A2(\dtop.field_top.controller.pattern0[1] ));
 sg13g2_o21ai_1 _4739_ (.B1(_1235_),
    .Y(_1239_),
    .A1(_2849_),
    .A2(_0079_));
 sg13g2_o21ai_1 _4740_ (.B1(_1236_),
    .Y(_1240_),
    .A1(_1238_),
    .A2(_1239_));
 sg13g2_nand2b_1 _4741_ (.Y(_1241_),
    .B(net1041),
    .A_N(\dtop.field_top.comp_value0_1[8] ));
 sg13g2_nor2_1 _4742_ (.A(net1042),
    .B(_2908_),
    .Y(_1242_));
 sg13g2_a22oi_1 _4743_ (.Y(_1243_),
    .B1(\dtop.field_top.comp_value0_1[2] ),
    .B2(net1007),
    .A2(\dtop.field_top.comp_value0_1[1] ),
    .A1(net1008));
 sg13g2_a221oi_1 _4744_ (.B2(net1054),
    .C1(_1243_),
    .B1(_2888_),
    .A1(net1057),
    .Y(_1244_),
    .A2(_2884_));
 sg13g2_a221oi_1 _4745_ (.B2(net1004),
    .C1(_1244_),
    .B1(\dtop.field_top.comp_value0_1[4] ),
    .A1(net1006),
    .Y(_1245_),
    .A2(\dtop.field_top.comp_value0_1[3] ));
 sg13g2_a221oi_1 _4746_ (.B2(net1049),
    .C1(_1245_),
    .B1(_2898_),
    .A1(net1050),
    .Y(_1246_),
    .A2(_2893_));
 sg13g2_a221oi_1 _4747_ (.B2(_2846_),
    .C1(_1246_),
    .B1(\dtop.field_top.comp_value0_1[6] ),
    .A1(net1015),
    .Y(_1247_),
    .A2(\dtop.field_top.comp_value0_1[5] ));
 sg13g2_a221oi_1 _4748_ (.B2(net1042),
    .C1(_1247_),
    .B1(_2908_),
    .A1(net1045),
    .Y(_1248_),
    .A2(_2903_));
 sg13g2_o21ai_1 _4749_ (.B1(_1241_),
    .Y(_1249_),
    .A1(_1242_),
    .A2(_1248_));
 sg13g2_a22oi_1 _4750_ (.Y(_1250_),
    .B1(\dtop.field_top.comp_value0_1[8] ),
    .B2(net1018),
    .A2(\dtop.field_top.comp_value0_1[9] ),
    .A1(net1017));
 sg13g2_or2_1 _4751_ (.X(_1251_),
    .B(\dtop.field_top.comp_value0_1[10] ),
    .A(net1035));
 sg13g2_o21ai_1 _4752_ (.B1(_1251_),
    .Y(_1252_),
    .A1(net1017),
    .A2(\dtop.field_top.comp_value0_1[9] ));
 sg13g2_a21oi_1 _4753_ (.A1(_1249_),
    .A2(_1250_),
    .Y(_1253_),
    .B1(_1252_));
 sg13g2_a21o_2 _4754_ (.A2(\dtop.field_top.comp_value0_1[10] ),
    .A1(net1035),
    .B1(_1253_),
    .X(_1254_));
 sg13g2_nand2b_1 _4755_ (.Y(_1255_),
    .B(net1041),
    .A_N(\dtop.field_top.comp_values0[4][8] ));
 sg13g2_nor2_1 _4756_ (.A(net1013),
    .B(\dtop.field_top.comp_values0[4][7] ),
    .Y(_1256_));
 sg13g2_nor2_1 _4757_ (.A(net1004),
    .B(\dtop.field_top.comp_values0[4][4] ),
    .Y(_1257_));
 sg13g2_a22oi_1 _4758_ (.Y(_1258_),
    .B1(\dtop.field_top.comp_values0[4][2] ),
    .B2(net1007),
    .A2(\dtop.field_top.comp_values0[4][1] ),
    .A1(net1008));
 sg13g2_a221oi_1 _4759_ (.B2(net1054),
    .C1(_1258_),
    .B1(_2889_),
    .A1(net1057),
    .Y(_1259_),
    .A2(_2885_));
 sg13g2_a21oi_1 _4760_ (.A1(net1006),
    .A2(\dtop.field_top.comp_values0[4][3] ),
    .Y(_1260_),
    .B1(_1259_));
 sg13g2_a22oi_1 _4761_ (.Y(_1261_),
    .B1(\dtop.field_top.comp_values0[4][5] ),
    .B2(net1015),
    .A2(\dtop.field_top.comp_values0[4][4] ),
    .A1(net1004));
 sg13g2_o21ai_1 _4762_ (.B1(_1261_),
    .Y(_1262_),
    .A1(_1257_),
    .A2(_1260_));
 sg13g2_a22oi_1 _4763_ (.Y(_1263_),
    .B1(_2904_),
    .B2(net1045),
    .A2(_2899_),
    .A1(net1049));
 sg13g2_a22oi_1 _4764_ (.Y(_1264_),
    .B1(_1262_),
    .B2(_1263_),
    .A2(\dtop.field_top.comp_values0[4][6] ),
    .A1(_2846_));
 sg13g2_a22oi_1 _4765_ (.Y(_1265_),
    .B1(\dtop.field_top.comp_values0[4][8] ),
    .B2(net1018),
    .A2(\dtop.field_top.comp_values0[4][7] ),
    .A1(net1013));
 sg13g2_o21ai_1 _4766_ (.B1(_1265_),
    .Y(_1266_),
    .A1(_1256_),
    .A2(_1264_));
 sg13g2_a22oi_1 _4767_ (.Y(_1267_),
    .B1(_1255_),
    .B2(_1266_),
    .A2(\dtop.field_top.comp_values0[4][9] ),
    .A1(net1017));
 sg13g2_a21oi_1 _4768_ (.A1(net1039),
    .A2(_2872_),
    .Y(_1268_),
    .B1(_1267_));
 sg13g2_o21ai_1 _4769_ (.B1(_1268_),
    .Y(_1269_),
    .A1(net1036),
    .A2(\dtop.field_top.comp_values0[4][10] ));
 sg13g2_nand2_1 _4770_ (.Y(_1270_),
    .A(net969),
    .B(_1269_));
 sg13g2_a21oi_2 _4771_ (.B1(_1270_),
    .Y(_1271_),
    .A2(\dtop.field_top.comp_values0[4][10] ),
    .A1(net1035));
 sg13g2_nand2_1 _4772_ (.Y(_1272_),
    .A(net1035),
    .B(\dtop.field_top.comp_values0[2][10] ));
 sg13g2_nand2_1 _4773_ (.Y(_1273_),
    .A(net1006),
    .B(\dtop.field_top.comp_values0[2][3] ));
 sg13g2_a22oi_1 _4774_ (.Y(_1274_),
    .B1(\dtop.field_top.comp_values0[2][2] ),
    .B2(net1007),
    .A2(\dtop.field_top.comp_values0[2][1] ),
    .A1(net1008));
 sg13g2_nor2_1 _4775_ (.A(net1007),
    .B(\dtop.field_top.comp_values0[2][2] ),
    .Y(_1275_));
 sg13g2_o21ai_1 _4776_ (.B1(_1273_),
    .Y(_1276_),
    .A1(_1274_),
    .A2(_1275_));
 sg13g2_a22oi_1 _4777_ (.Y(_1277_),
    .B1(_2895_),
    .B2(net1050),
    .A2(_2891_),
    .A1(net1054));
 sg13g2_nor2_1 _4778_ (.A(net1050),
    .B(_2895_),
    .Y(_1278_));
 sg13g2_a221oi_1 _4779_ (.B2(_1277_),
    .C1(_1278_),
    .B1(_1276_),
    .A1(net1015),
    .Y(_1279_),
    .A2(\dtop.field_top.comp_values0[2][5] ));
 sg13g2_a221oi_1 _4780_ (.B2(net1045),
    .C1(_1279_),
    .B1(_2906_),
    .A1(net1049),
    .Y(_1280_),
    .A2(_2901_));
 sg13g2_a221oi_1 _4781_ (.B2(net1013),
    .C1(_1280_),
    .B1(\dtop.field_top.comp_values0[2][7] ),
    .A1(_2846_),
    .Y(_1281_),
    .A2(\dtop.field_top.comp_values0[2][6] ));
 sg13g2_nand2b_1 _4782_ (.Y(_1282_),
    .B(net1041),
    .A_N(\dtop.field_top.comp_values0[2][8] ));
 sg13g2_o21ai_1 _4783_ (.B1(_1282_),
    .Y(_1283_),
    .A1(net1013),
    .A2(\dtop.field_top.comp_values0[2][7] ));
 sg13g2_nor2_1 _4784_ (.A(_1281_),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_a221oi_1 _4785_ (.B2(net1018),
    .C1(_1284_),
    .B1(\dtop.field_top.comp_values0[2][8] ),
    .A1(net1017),
    .Y(_1285_),
    .A2(\dtop.field_top.comp_values0[2][9] ));
 sg13g2_or2_1 _4786_ (.X(_1286_),
    .B(\dtop.field_top.comp_values0[2][10] ),
    .A(net1035));
 sg13g2_o21ai_1 _4787_ (.B1(_1286_),
    .Y(_1287_),
    .A1(net1017),
    .A2(\dtop.field_top.comp_values0[2][9] ));
 sg13g2_o21ai_1 _4788_ (.B1(_1272_),
    .Y(_1288_),
    .A1(_1285_),
    .A2(_1287_));
 sg13g2_nor3_1 _4789_ (.A(\dtop.field_top.sflag2 ),
    .B(net971),
    .C(_1288_),
    .Y(_1289_));
 sg13g2_o21ai_1 _4790_ (.B1(_1254_),
    .Y(_1290_),
    .A1(_1271_),
    .A2(_1289_));
 sg13g2_nand2b_1 _4791_ (.Y(_1291_),
    .B(net1045),
    .A_N(\dtop.field_top.comp_value0[5] ));
 sg13g2_a22oi_1 _4792_ (.Y(_1292_),
    .B1(\dtop.field_top.comp_value0[0] ),
    .B2(net1008),
    .A2(\dtop.field_top.comp_value0[1] ),
    .A1(net1007));
 sg13g2_a221oi_1 _4793_ (.B2(net1057),
    .C1(_1292_),
    .B1(_2924_),
    .A1(net1054),
    .Y(_1293_),
    .A2(_2923_));
 sg13g2_a21o_1 _4794_ (.A2(\dtop.field_top.comp_value0[2] ),
    .A1(net1006),
    .B1(_1293_),
    .X(_1294_));
 sg13g2_o21ai_1 _4795_ (.B1(_1294_),
    .Y(_1295_),
    .A1(net1004),
    .A2(\dtop.field_top.comp_value0[3] ));
 sg13g2_a22oi_1 _4796_ (.Y(_1296_),
    .B1(\dtop.field_top.comp_value0[3] ),
    .B2(net1004),
    .A2(\dtop.field_top.comp_value0[4] ),
    .A1(net1015));
 sg13g2_o21ai_1 _4797_ (.B1(_1291_),
    .Y(_1297_),
    .A1(net1015),
    .A2(\dtop.field_top.comp_value0[4] ));
 sg13g2_a21oi_1 _4798_ (.A1(_1295_),
    .A2(_1296_),
    .Y(_1298_),
    .B1(_1297_));
 sg13g2_a221oi_1 _4799_ (.B2(_2846_),
    .C1(_1298_),
    .B1(\dtop.field_top.comp_value0[5] ),
    .A1(net1013),
    .Y(_1299_),
    .A2(\dtop.field_top.comp_value0[6] ));
 sg13g2_a221oi_1 _4800_ (.B2(net1042),
    .C1(_1299_),
    .B1(_2922_),
    .A1(net1041),
    .Y(_1300_),
    .A2(_2921_));
 sg13g2_a221oi_1 _4801_ (.B2(net1018),
    .C1(_1300_),
    .B1(\dtop.field_top.comp_value0[7] ),
    .A1(net1017),
    .Y(_1301_),
    .A2(\dtop.field_top.comp_value0[8] ));
 sg13g2_or2_1 _4802_ (.X(_1302_),
    .B(\dtop.field_top.comp_value0_0[10] ),
    .A(net1035));
 sg13g2_o21ai_1 _4803_ (.B1(_1302_),
    .Y(_1303_),
    .A1(net1017),
    .A2(\dtop.field_top.comp_value0[8] ));
 sg13g2_nor2_1 _4804_ (.A(_1301_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_a21oi_2 _4805_ (.B1(_1304_),
    .Y(_1305_),
    .A2(\dtop.field_top.comp_value0_0[10] ),
    .A1(net1035));
 sg13g2_nand3_1 _4806_ (.B(_1288_),
    .C(_1305_),
    .A(\dtop.field_top.sflag2 ),
    .Y(_1306_));
 sg13g2_o21ai_1 _4807_ (.B1(_1290_),
    .Y(_1307_),
    .A1(net971),
    .A2(_1306_));
 sg13g2_nand2_1 _4808_ (.Y(_1308_),
    .A(\dtop.field_top.lside ),
    .B(_1307_));
 sg13g2_nor2_1 _4809_ (.A(net1018),
    .B(\dtop.field_top.comp_values0[3][8] ),
    .Y(_1309_));
 sg13g2_a22oi_1 _4810_ (.Y(_1310_),
    .B1(\dtop.field_top.comp_values0[3][2] ),
    .B2(net1007),
    .A2(\dtop.field_top.comp_values0[3][1] ),
    .A1(net1008));
 sg13g2_a221oi_1 _4811_ (.B2(net1054),
    .C1(_1310_),
    .B1(_2890_),
    .A1(net1057),
    .Y(_1311_),
    .A2(_2886_));
 sg13g2_a221oi_1 _4812_ (.B2(net1004),
    .C1(_1311_),
    .B1(\dtop.field_top.comp_values0[3][4] ),
    .A1(net1006),
    .Y(_1312_),
    .A2(\dtop.field_top.comp_values0[3][3] ));
 sg13g2_a221oi_1 _4813_ (.B2(net1049),
    .C1(_1312_),
    .B1(_2900_),
    .A1(net1050),
    .Y(_1313_),
    .A2(_2894_));
 sg13g2_a221oi_1 _4814_ (.B2(_2846_),
    .C1(_1313_),
    .B1(\dtop.field_top.comp_values0[3][6] ),
    .A1(net1015),
    .Y(_1314_),
    .A2(\dtop.field_top.comp_values0[3][5] ));
 sg13g2_a221oi_1 _4815_ (.B2(net1042),
    .C1(_1314_),
    .B1(_2909_),
    .A1(net1045),
    .Y(_1315_),
    .A2(_2905_));
 sg13g2_a221oi_1 _4816_ (.B2(net1018),
    .C1(_1315_),
    .B1(\dtop.field_top.comp_values0[3][8] ),
    .A1(net1013),
    .Y(_1316_),
    .A2(\dtop.field_top.comp_values0[3][7] ));
 sg13g2_nand2_1 _4817_ (.Y(_1317_),
    .A(net1017),
    .B(\dtop.field_top.comp_values0[3][9] ));
 sg13g2_o21ai_1 _4818_ (.B1(_1317_),
    .Y(_1318_),
    .A1(_1309_),
    .A2(_1316_));
 sg13g2_a22oi_1 _4819_ (.Y(_1319_),
    .B1(_2897_),
    .B2(_2843_),
    .A2(_2873_),
    .A1(net1039));
 sg13g2_a22oi_1 _4820_ (.Y(_1320_),
    .B1(_1318_),
    .B2(_1319_),
    .A2(\dtop.field_top.comp_values0[3][10] ),
    .A1(net1035));
 sg13g2_nor3_1 _4821_ (.A(\dtop.field_top.lside ),
    .B(_1254_),
    .C(_1320_),
    .Y(_1321_));
 sg13g2_nor3_1 _4822_ (.A(\dtop.field_top.rside ),
    .B(_1288_),
    .C(_1305_),
    .Y(_1322_));
 sg13g2_nand3_1 _4823_ (.B(_1288_),
    .C(_1320_),
    .A(\dtop.field_top.rside ),
    .Y(_1323_));
 sg13g2_nand2b_1 _4824_ (.Y(_1324_),
    .B(_1323_),
    .A_N(_1321_));
 sg13g2_o21ai_1 _4825_ (.B1(net971),
    .Y(_1325_),
    .A1(_1322_),
    .A2(_1324_));
 sg13g2_nand2_1 _4826_ (.Y(_1326_),
    .A(_1308_),
    .B(_1325_));
 sg13g2_nand2_1 _4827_ (.Y(_1327_),
    .A(_1240_),
    .B(_1326_));
 sg13g2_inv_1 _4828_ (.Y(_1328_),
    .A(_1327_));
 sg13g2_nand3b_1 _4829_ (.B(_3066_),
    .C(_1254_),
    .Y(_1329_),
    .A_N(_0082_));
 sg13g2_o21ai_1 _4830_ (.B1(_1240_),
    .Y(_1330_),
    .A1(_1271_),
    .A2(_1305_));
 sg13g2_a21o_1 _4831_ (.A2(_1329_),
    .A1(_1305_),
    .B1(_1330_),
    .X(_1331_));
 sg13g2_nand2_1 _4832_ (.Y(_1332_),
    .A(_1327_),
    .B(_1331_));
 sg13g2_nand2_1 _4833_ (.Y(_1333_),
    .A(net1032),
    .B(_2849_));
 sg13g2_and3_2 _4834_ (.X(_1334_),
    .A(_1211_),
    .B(_1236_),
    .C(_1333_));
 sg13g2_a21oi_1 _4835_ (.A1(net1030),
    .A2(_1223_),
    .Y(_1335_),
    .B1(_1237_));
 sg13g2_a21o_1 _4836_ (.A2(_1223_),
    .A1(net1030),
    .B1(_1237_),
    .X(_1336_));
 sg13g2_nand3b_1 _4837_ (.B(\dtop.field_top.controller.ppos[4] ),
    .C(\dtop.field_top.controller.ppos[3] ),
    .Y(_1337_),
    .A_N(net1033));
 sg13g2_a21oi_2 _4838_ (.B1(_1336_),
    .Y(_1338_),
    .A2(_1337_),
    .A1(_1212_));
 sg13g2_nand2_1 _4839_ (.Y(_1339_),
    .A(net1040),
    .B(_1338_));
 sg13g2_nand2_1 _4840_ (.Y(_1340_),
    .A(_0107_),
    .B(_1338_));
 sg13g2_xnor2_1 _4841_ (.Y(_1341_),
    .A(_2869_),
    .B(_1340_));
 sg13g2_nor2b_1 _4842_ (.A(_1339_),
    .B_N(_1341_),
    .Y(_1342_));
 sg13g2_nand3_1 _4843_ (.B(_0107_),
    .C(_1338_),
    .A(net1037),
    .Y(_1343_));
 sg13g2_o21ai_1 _4844_ (.B1(_1343_),
    .Y(_1344_),
    .A1(net1036),
    .A2(_1338_));
 sg13g2_nor2_2 _4845_ (.A(_1342_),
    .B(_1344_),
    .Y(_1345_));
 sg13g2_xor2_1 _4846_ (.B(_1341_),
    .A(_1339_),
    .X(_1346_));
 sg13g2_nand2b_1 _4847_ (.Y(_1347_),
    .B(_1346_),
    .A_N(\dtop.field_top.last_wave[7] ));
 sg13g2_a22oi_1 _4848_ (.Y(_1348_),
    .B1(_1347_),
    .B2(_1345_),
    .A2(_1346_),
    .A1(_0081_));
 sg13g2_nor2_1 _4849_ (.A(net1014),
    .B(\dtop.field_top.last_wave[6] ),
    .Y(_1349_));
 sg13g2_nand2b_1 _4850_ (.Y(_1350_),
    .B(net1046),
    .A_N(\dtop.field_top.last_wave[5] ));
 sg13g2_a22oi_1 _4851_ (.Y(_1351_),
    .B1(_2919_),
    .B2(net1056),
    .A2(_2918_),
    .A1(\dtop.field_top.afl_sub_pc[1] ));
 sg13g2_nand2_1 _4852_ (.Y(_1352_),
    .A(_2846_),
    .B(\dtop.field_top.last_wave[5] ));
 sg13g2_o21ai_1 _4853_ (.B1(_1352_),
    .Y(_1353_),
    .A1(net1048),
    .A2(_2920_));
 sg13g2_a22oi_1 _4854_ (.Y(_1354_),
    .B1(\dtop.field_top.last_wave[2] ),
    .B2(net1006),
    .A2(\dtop.field_top.last_wave[3] ),
    .A1(net1005));
 sg13g2_inv_1 _4855_ (.Y(_1355_),
    .A(_1354_));
 sg13g2_nor2_1 _4856_ (.A(_2863_),
    .B(\dtop.field_top.last_wave[2] ),
    .Y(_1356_));
 sg13g2_nor2_1 _4857_ (.A(net1005),
    .B(\dtop.field_top.last_wave[3] ),
    .Y(_1357_));
 sg13g2_nor3_1 _4858_ (.A(_1355_),
    .B(_1356_),
    .C(_1357_),
    .Y(_1358_));
 sg13g2_nor2_1 _4859_ (.A(net1056),
    .B(_2919_),
    .Y(_1359_));
 sg13g2_a221oi_1 _4860_ (.B2(_2862_),
    .C1(_1349_),
    .B1(\dtop.field_top.last_wave[1] ),
    .A1(net1008),
    .Y(_1360_),
    .A2(\dtop.field_top.last_wave[0] ));
 sg13g2_o21ai_1 _4861_ (.B1(_1350_),
    .Y(_1361_),
    .A1(net1016),
    .A2(\dtop.field_top.last_wave[4] ));
 sg13g2_nor2_1 _4862_ (.A(_1353_),
    .B(_1361_),
    .Y(_1362_));
 sg13g2_nand4_1 _4863_ (.B(_1358_),
    .C(_1360_),
    .A(_1351_),
    .Y(_1363_),
    .D(_1362_));
 sg13g2_a21o_1 _4864_ (.A2(_1363_),
    .A1(\dtop.field_top.last_wave[7] ),
    .B1(_1345_),
    .X(_1364_));
 sg13g2_o21ai_1 _4865_ (.B1(_1364_),
    .Y(_1365_),
    .A1(_0081_),
    .A2(_1346_));
 sg13g2_xnor2_1 _4866_ (.Y(_1366_),
    .A(net1040),
    .B(_1338_));
 sg13g2_o21ai_1 _4867_ (.B1(_1358_),
    .Y(_1367_),
    .A1(_1351_),
    .A2(_1359_));
 sg13g2_o21ai_1 _4868_ (.B1(_1367_),
    .Y(_1368_),
    .A1(_1354_),
    .A2(_1357_));
 sg13g2_a22oi_1 _4869_ (.Y(_1369_),
    .B1(_1362_),
    .B2(_1368_),
    .A2(_1353_),
    .A1(_1350_));
 sg13g2_nand2b_1 _4870_ (.Y(_1370_),
    .B(_1363_),
    .A_N(_1349_));
 sg13g2_a22oi_1 _4871_ (.Y(_1371_),
    .B1(_1366_),
    .B2(\dtop.field_top.last_wave[7] ),
    .A2(\dtop.field_top.last_wave[6] ),
    .A1(net1014));
 sg13g2_o21ai_1 _4872_ (.B1(_1371_),
    .Y(_1372_),
    .A1(_1369_),
    .A2(_1370_));
 sg13g2_o21ai_1 _4873_ (.B1(_1372_),
    .Y(_1373_),
    .A1(\dtop.field_top.last_wave[7] ),
    .A2(_1366_));
 sg13g2_a21oi_1 _4874_ (.A1(_1365_),
    .A2(_1373_),
    .Y(_1374_),
    .B1(_1348_));
 sg13g2_nand2b_1 _4875_ (.Y(_1375_),
    .B(_1346_),
    .A_N(_0080_));
 sg13g2_nor2_1 _4876_ (.A(\dtop.field_top.wave[7] ),
    .B(_1366_),
    .Y(_1376_));
 sg13g2_nand2_1 _4877_ (.Y(_1377_),
    .A(\dtop.field_top.wave[7] ),
    .B(_1366_));
 sg13g2_o21ai_1 _4878_ (.B1(_1377_),
    .Y(_1378_),
    .A1(net1044),
    .A2(_2917_));
 sg13g2_a22oi_1 _4879_ (.Y(_1379_),
    .B1(_2917_),
    .B2(net1044),
    .A2(_2916_),
    .A1(net1046));
 sg13g2_a22oi_1 _4880_ (.Y(_1380_),
    .B1(\dtop.field_top.wave[5] ),
    .B2(_2846_),
    .A2(\dtop.field_top.wave[4] ),
    .A1(net1016));
 sg13g2_nor2_1 _4881_ (.A(net1016),
    .B(\dtop.field_top.wave[4] ),
    .Y(_1381_));
 sg13g2_nand2_1 _4882_ (.Y(_1382_),
    .A(_2863_),
    .B(\dtop.field_top.wave[2] ));
 sg13g2_nand2_1 _4883_ (.Y(_1383_),
    .A(net1005),
    .B(\dtop.field_top.wave[3] ));
 sg13g2_nand2b_1 _4884_ (.Y(_1384_),
    .B(net1051),
    .A_N(\dtop.field_top.wave[3] ));
 sg13g2_nand2b_1 _4885_ (.Y(_1385_),
    .B(net1053),
    .A_N(\dtop.field_top.wave[2] ));
 sg13g2_nand4_1 _4886_ (.B(_1383_),
    .C(_1384_),
    .A(_1382_),
    .Y(_1386_),
    .D(_1385_));
 sg13g2_a22oi_1 _4887_ (.Y(_1387_),
    .B1(_2915_),
    .B2(net1056),
    .A2(_2914_),
    .A1(\dtop.field_top.afl_sub_pc[1] ));
 sg13g2_nand2_1 _4888_ (.Y(_1388_),
    .A(_2862_),
    .B(\dtop.field_top.wave[1] ));
 sg13g2_nor2b_1 _4889_ (.A(_1387_),
    .B_N(_1388_),
    .Y(_1389_));
 sg13g2_nor2b_1 _4890_ (.A(_1382_),
    .B_N(_1384_),
    .Y(_1390_));
 sg13g2_o21ai_1 _4891_ (.B1(_1383_),
    .Y(_1391_),
    .A1(_1386_),
    .A2(_1389_));
 sg13g2_nor2_1 _4892_ (.A(_1390_),
    .B(_1391_),
    .Y(_1392_));
 sg13g2_o21ai_1 _4893_ (.B1(_1380_),
    .Y(_1393_),
    .A1(_1381_),
    .A2(_1392_));
 sg13g2_a21oi_1 _4894_ (.A1(_1379_),
    .A2(_1393_),
    .Y(_1394_),
    .B1(_1378_));
 sg13g2_nor2_1 _4895_ (.A(_1376_),
    .B(_1394_),
    .Y(_1395_));
 sg13g2_nand2_1 _4896_ (.Y(_1396_),
    .A(\dtop.field_top.wave[7] ),
    .B(_1346_));
 sg13g2_nand2_1 _4897_ (.Y(_1397_),
    .A(_0080_),
    .B(_1345_));
 sg13g2_a22oi_1 _4898_ (.Y(_1398_),
    .B1(_1375_),
    .B2(_1395_),
    .A2(_1345_),
    .A1(_0080_));
 sg13g2_nor2_1 _4899_ (.A(_1345_),
    .B(_1346_),
    .Y(_1399_));
 sg13g2_a21oi_1 _4900_ (.A1(_0080_),
    .A2(_1346_),
    .Y(_1400_),
    .B1(_1345_));
 sg13g2_a21oi_1 _4901_ (.A1(_1396_),
    .A2(_1398_),
    .Y(_1401_),
    .B1(_1400_));
 sg13g2_o21ai_1 _4902_ (.B1(_1388_),
    .Y(_1402_),
    .A1(\dtop.field_top.afl_sub_pc[1] ),
    .A2(_2914_));
 sg13g2_nor3_1 _4903_ (.A(_1381_),
    .B(_1386_),
    .C(_1402_),
    .Y(_1403_));
 sg13g2_nand4_1 _4904_ (.B(_1380_),
    .C(_1387_),
    .A(_1379_),
    .Y(_1404_),
    .D(_1403_));
 sg13g2_xnor2_1 _4905_ (.Y(_1405_),
    .A(_1374_),
    .B(_1401_));
 sg13g2_nor4_1 _4906_ (.A(_1376_),
    .B(_1378_),
    .C(_1399_),
    .D(_1404_),
    .Y(_1406_));
 sg13g2_nand3_1 _4907_ (.B(_1397_),
    .C(_1406_),
    .A(_1375_),
    .Y(_1407_));
 sg13g2_a221oi_1 _4908_ (.B2(_1407_),
    .C1(_1334_),
    .B1(_1405_),
    .A1(_1234_),
    .Y(_1408_),
    .A2(_1332_));
 sg13g2_and2_1 _4909_ (.A(net966),
    .B(_1408_),
    .X(_1409_));
 sg13g2_nor2_2 _4910_ (.A(\dtop.field_top.fx[3] ),
    .B(\dtop.field_top.fx[2] ),
    .Y(_1410_));
 sg13g2_inv_1 _4911_ (.Y(_1411_),
    .A(net1003));
 sg13g2_mux2_1 _4912_ (.A0(_0023_),
    .A1(_0022_),
    .S(net1003),
    .X(_1412_));
 sg13g2_nor2_1 _4913_ (.A(_2838_),
    .B(_1412_),
    .Y(_1413_));
 sg13g2_mux2_1 _4914_ (.A0(_0105_),
    .A1(_0104_),
    .S(_1410_),
    .X(_1414_));
 sg13g2_nor2_1 _4915_ (.A(_0103_),
    .B(_1414_),
    .Y(_1415_));
 sg13g2_mux2_1 _4916_ (.A0(_0092_),
    .A1(_0091_),
    .S(net1003),
    .X(_1416_));
 sg13g2_nor2_1 _4917_ (.A(_0106_),
    .B(_1416_),
    .Y(_1417_));
 sg13g2_mux2_1 _4918_ (.A0(_0097_),
    .A1(_0096_),
    .S(net1003),
    .X(_1418_));
 sg13g2_nor2_1 _4919_ (.A(_2840_),
    .B(_1418_),
    .Y(_1419_));
 sg13g2_mux2_1 _4920_ (.A0(_0100_),
    .A1(_0099_),
    .S(net1003),
    .X(_1420_));
 sg13g2_nor2_1 _4921_ (.A(_2841_),
    .B(_1420_),
    .Y(_1421_));
 sg13g2_xor2_1 _4922_ (.B(_1418_),
    .A(_0098_),
    .X(_1422_));
 sg13g2_a21oi_1 _4923_ (.A1(_1421_),
    .A2(_1422_),
    .Y(_1423_),
    .B1(_1419_));
 sg13g2_mux2_1 _4924_ (.A0(_0095_),
    .A1(_0094_),
    .S(net1003),
    .X(_1424_));
 sg13g2_xor2_1 _4925_ (.B(_1424_),
    .A(\dtop.field_top.fy[6] ),
    .X(_1425_));
 sg13g2_nor2_1 _4926_ (.A(_1423_),
    .B(_1425_),
    .Y(_1426_));
 sg13g2_nor2_1 _4927_ (.A(_0093_),
    .B(_1424_),
    .Y(_1427_));
 sg13g2_nor2_1 _4928_ (.A(_1426_),
    .B(_1427_),
    .Y(_1428_));
 sg13g2_xor2_1 _4929_ (.B(_1416_),
    .A(\dtop.field_top.fy[7] ),
    .X(_1429_));
 sg13g2_nor2_1 _4930_ (.A(_1428_),
    .B(_1429_),
    .Y(_1430_));
 sg13g2_nor2_1 _4931_ (.A(_1417_),
    .B(_1430_),
    .Y(_1431_));
 sg13g2_xor2_1 _4932_ (.B(_1414_),
    .A(\dtop.field_top.fx[8] ),
    .X(_1432_));
 sg13g2_nor2_1 _4933_ (.A(_1431_),
    .B(_1432_),
    .Y(_1433_));
 sg13g2_mux2_1 _4934_ (.A0(_0102_),
    .A1(_0101_),
    .S(net1003),
    .X(_1434_));
 sg13g2_xnor2_1 _4935_ (.Y(_1435_),
    .A(\dtop.field_top.fy[9] ),
    .B(_1434_));
 sg13g2_o21ai_1 _4936_ (.B1(_1435_),
    .Y(_1436_),
    .A1(_1415_),
    .A2(_1433_));
 sg13g2_o21ai_1 _4937_ (.B1(_1436_),
    .Y(_1437_),
    .A1(_0024_),
    .A2(_1434_));
 sg13g2_nand2_1 _4938_ (.Y(_1438_),
    .A(_2838_),
    .B(_1412_));
 sg13g2_nand2b_1 _4939_ (.Y(_1439_),
    .B(_1438_),
    .A_N(_1413_));
 sg13g2_a21oi_1 _4940_ (.A1(_1437_),
    .A2(_1438_),
    .Y(_1440_),
    .B1(_1413_));
 sg13g2_nand2_1 _4941_ (.Y(_1441_),
    .A(\dtop.field_top.nsource.shuffle_state.in[1] ),
    .B(_1411_));
 sg13g2_xnor2_1 _4942_ (.Y(_1442_),
    .A(_0026_),
    .B(_1441_));
 sg13g2_xnor2_1 _4943_ (.Y(_1443_),
    .A(_1440_),
    .B(_1442_));
 sg13g2_xor2_1 _4944_ (.B(_1439_),
    .A(_1437_),
    .X(_1444_));
 sg13g2_xor2_1 _4945_ (.B(_1425_),
    .A(_1423_),
    .X(_1445_));
 sg13g2_nor4_2 _4946_ (.A(net1034),
    .B(_3028_),
    .C(_3039_),
    .Y(_1446_),
    .D(_3080_));
 sg13g2_xor2_1 _4947_ (.B(_1420_),
    .A(_0025_),
    .X(_1447_));
 sg13g2_nor4_1 _4948_ (.A(_0074_),
    .B(_1445_),
    .C(_1446_),
    .D(_1447_),
    .Y(_1448_));
 sg13g2_nand3_1 _4949_ (.B(_1444_),
    .C(_1448_),
    .A(_1443_),
    .Y(_1449_));
 sg13g2_xnor2_1 _4950_ (.Y(_1450_),
    .A(\dtop.field_top.fx[2] ),
    .B(\dtop.field_top.fx[1] ));
 sg13g2_xor2_1 _4951_ (.B(\dtop.field_top.fy[2] ),
    .A(\dtop.field_top.fy[1] ),
    .X(_1451_));
 sg13g2_inv_1 _4952_ (.Y(_1452_),
    .A(_1451_));
 sg13g2_nor3_1 _4953_ (.A(_1449_),
    .B(_1450_),
    .C(_1452_),
    .Y(_1453_));
 sg13g2_xnor2_1 _4954_ (.Y(_1454_),
    .A(_1428_),
    .B(_1429_));
 sg13g2_nor2_1 _4955_ (.A(_1450_),
    .B(_1451_),
    .Y(_1455_));
 sg13g2_xor2_1 _4956_ (.B(\dtop.field_top.fx[0] ),
    .A(\dtop.field_top.fx[2] ),
    .X(_1456_));
 sg13g2_nor2_1 _4957_ (.A(_1455_),
    .B(_1456_),
    .Y(_1457_));
 sg13g2_xor2_1 _4958_ (.B(\dtop.field_top.fy[2] ),
    .A(\dtop.field_top.fy[0] ),
    .X(_1458_));
 sg13g2_a21oi_1 _4959_ (.A1(_1450_),
    .A2(_1451_),
    .Y(_1459_),
    .B1(_1458_));
 sg13g2_nor4_2 _4960_ (.A(_1449_),
    .B(_1454_),
    .C(_1457_),
    .Y(_1460_),
    .D(_1459_));
 sg13g2_or3_1 _4961_ (.A(_1415_),
    .B(_1433_),
    .C(_1435_),
    .X(_1461_));
 sg13g2_nand2_1 _4962_ (.Y(_1462_),
    .A(_1436_),
    .B(_1461_));
 sg13g2_nor2_1 _4963_ (.A(_1454_),
    .B(_1462_),
    .Y(_1463_));
 sg13g2_nor2_1 _4964_ (.A(_1460_),
    .B(_1463_),
    .Y(_1464_));
 sg13g2_nor2b_2 _4965_ (.A(_1464_),
    .B_N(_1453_),
    .Y(_1465_));
 sg13g2_nor2_1 _4966_ (.A(_1332_),
    .B(_1408_),
    .Y(_1466_));
 sg13g2_inv_1 _4967_ (.Y(_1467_),
    .A(_1466_));
 sg13g2_a21oi_1 _4968_ (.A1(_1465_),
    .A2(_1466_),
    .Y(_1468_),
    .B1(_1409_));
 sg13g2_nor2b_2 _4969_ (.A(_1468_),
    .B_N(_1233_),
    .Y(_0286_));
 sg13g2_nor2b_1 _4970_ (.A(_1408_),
    .B_N(_1233_),
    .Y(_1469_));
 sg13g2_nand2_1 _4971_ (.Y(_1470_),
    .A(_1328_),
    .B(_1469_));
 sg13g2_nand3_1 _4972_ (.B(_1161_),
    .C(_1232_),
    .A(net341),
    .Y(_1471_));
 sg13g2_nand3b_1 _4973_ (.B(_1470_),
    .C(_1471_),
    .Y(_0157_),
    .A_N(_0286_));
 sg13g2_o21ai_1 _4974_ (.B1(_1233_),
    .Y(_1472_),
    .A1(_1465_),
    .A2(_1467_));
 sg13g2_nand2_1 _4975_ (.Y(_0158_),
    .A(_1471_),
    .B(_1472_));
 sg13g2_nand2b_1 _4976_ (.Y(_1473_),
    .B(_1453_),
    .A_N(_1463_));
 sg13g2_xnor2_1 _4977_ (.Y(_1474_),
    .A(_1460_),
    .B(_1473_));
 sg13g2_a21o_1 _4978_ (.A2(_1474_),
    .A1(_1331_),
    .B1(_1328_),
    .X(_1475_));
 sg13g2_nand2_1 _4979_ (.Y(_1476_),
    .A(_1469_),
    .B(_1475_));
 sg13g2_nand2_1 _4980_ (.Y(_0159_),
    .A(_1471_),
    .B(_1476_));
 sg13g2_nor2b_1 _4981_ (.A(_1474_),
    .B_N(_1331_),
    .Y(_1477_));
 sg13g2_or3_1 _4982_ (.A(_1328_),
    .B(_1408_),
    .C(_1477_),
    .X(_1478_));
 sg13g2_nor2_1 _4983_ (.A(_1232_),
    .B(_1409_),
    .Y(_1479_));
 sg13g2_a21oi_1 _4984_ (.A1(_1478_),
    .A2(_1479_),
    .Y(_0160_),
    .B1(_1162_));
 sg13g2_nor3_1 _4985_ (.A(_1232_),
    .B(_1408_),
    .C(_1475_),
    .Y(_1480_));
 sg13g2_a21oi_1 _4986_ (.A1(net372),
    .A2(_1161_),
    .Y(_1481_),
    .B1(_1233_));
 sg13g2_nor2_2 _4987_ (.A(_1480_),
    .B(_1481_),
    .Y(_0161_));
 sg13g2_nand3_1 _4988_ (.B(\dtop.field_top.channel[0] ),
    .C(\dtop.field_top.channel[3] ),
    .A(net1109),
    .Y(_1482_));
 sg13g2_inv_1 _4989_ (.Y(_1483_),
    .A(_1482_));
 sg13g2_nor2_1 _4990_ (.A(\dtop.field_top.channel[2] ),
    .B(_1482_),
    .Y(_1484_));
 sg13g2_or2_1 _4991_ (.X(_1485_),
    .B(_1482_),
    .A(\dtop.field_top.channel[2] ));
 sg13g2_or2_1 _4992_ (.X(_1486_),
    .B(net1032),
    .A(\dtop.field_top.controller.ppos[3] ));
 sg13g2_and2_1 _4993_ (.A(\dtop.field_top.controller.ppos[4] ),
    .B(\dtop.field_top.controller.ppos[5] ),
    .X(_1487_));
 sg13g2_a21o_1 _4994_ (.A2(_1487_),
    .A1(_1486_),
    .B1(_1213_),
    .X(_1488_));
 sg13g2_nand3_1 _4995_ (.B(net987),
    .C(_1488_),
    .A(_1335_),
    .Y(_1489_));
 sg13g2_and2_2 _4996_ (.A(\dtop.field_top.channel[3] ),
    .B(_1489_),
    .X(_1490_));
 sg13g2_and3_1 _4997_ (.X(_1491_),
    .A(_0109_),
    .B(_1213_),
    .C(_1335_));
 sg13g2_nand3_1 _4998_ (.B(_1213_),
    .C(_1335_),
    .A(_0109_),
    .Y(_1492_));
 sg13g2_nand2_1 _4999_ (.Y(_1493_),
    .A(_1483_),
    .B(_1491_));
 sg13g2_nand3b_1 _5000_ (.B(_1490_),
    .C(_1493_),
    .Y(_1494_),
    .A_N(\dtop.field_top.channel[2] ));
 sg13g2_inv_1 _5001_ (.Y(_1495_),
    .A(_1494_));
 sg13g2_and3_1 _5002_ (.X(_1496_),
    .A(\dtop.field_top.afl_pc[4] ),
    .B(net1047),
    .C(net1043));
 sg13g2_nor3_2 _5003_ (.A(net1037),
    .B(_3034_),
    .C(_1496_),
    .Y(_1497_));
 sg13g2_or4_1 _5004_ (.A(net1034),
    .B(_1212_),
    .C(_1336_),
    .D(_1497_),
    .X(_1498_));
 sg13g2_nor2_1 _5005_ (.A(_1213_),
    .B(_1337_),
    .Y(_1499_));
 sg13g2_o21ai_1 _5006_ (.B1(_1499_),
    .Y(_1500_),
    .A1(net1034),
    .A2(_1497_));
 sg13g2_nand3_1 _5007_ (.B(_1498_),
    .C(_1500_),
    .A(net987),
    .Y(_1501_));
 sg13g2_and2_1 _5008_ (.A(net1109),
    .B(_1501_),
    .X(_1502_));
 sg13g2_nor2b_1 _5009_ (.A(_1494_),
    .B_N(_1502_),
    .Y(_1503_));
 sg13g2_nand2_1 _5010_ (.Y(_1504_),
    .A(_1495_),
    .B(net964));
 sg13g2_nor2_1 _5011_ (.A(\dtop.field_top.player.osc0[21] ),
    .B(net1061),
    .Y(_1505_));
 sg13g2_and2_1 _5012_ (.A(\dtop.field_top.player.controller.pattern0[2] ),
    .B(_1505_),
    .X(_1506_));
 sg13g2_nor2_1 _5013_ (.A(net946),
    .B(_1506_),
    .Y(_1507_));
 sg13g2_nor2b_1 _5014_ (.A(net1061),
    .B_N(\dtop.field_top.player.osc0[21] ),
    .Y(_1508_));
 sg13g2_nand2b_1 _5015_ (.Y(_1509_),
    .B(\dtop.field_top.player.osc0[21] ),
    .A_N(net1061));
 sg13g2_nor2_2 _5016_ (.A(net1064),
    .B(net1069),
    .Y(_1510_));
 sg13g2_or2_2 _5017_ (.X(_1511_),
    .B(net1068),
    .A(net1064));
 sg13g2_nor2_1 _5018_ (.A(net1075),
    .B(_1511_),
    .Y(_1512_));
 sg13g2_nand2_2 _5019_ (.Y(_1513_),
    .A(net1020),
    .B(_1510_));
 sg13g2_nor2_2 _5020_ (.A(net1075),
    .B(net1083),
    .Y(_1514_));
 sg13g2_nand2_1 _5021_ (.Y(_1515_),
    .A(net1020),
    .B(_2834_));
 sg13g2_nor4_1 _5022_ (.A(net1083),
    .B(\dtop.field_top.player.controller.pattern0[2] ),
    .C(_1509_),
    .D(_1513_),
    .Y(_1516_));
 sg13g2_nand2_1 _5023_ (.Y(_1517_),
    .A(_2830_),
    .B(_1508_));
 sg13g2_nand2b_1 _5024_ (.Y(_1518_),
    .B(net1061),
    .A_N(\dtop.field_top.player.osc0[21] ));
 sg13g2_o21ai_1 _5025_ (.B1(_1517_),
    .Y(_1519_),
    .A1(_2830_),
    .A2(_1518_));
 sg13g2_and2_1 _5026_ (.A(\dtop.field_top.player.osc0[21] ),
    .B(net1061),
    .X(_1520_));
 sg13g2_nand3_1 _5027_ (.B(net1061),
    .C(\dtop.field_top.player.controller.pattern0[2] ),
    .A(\dtop.field_top.player.osc0[21] ),
    .Y(_1521_));
 sg13g2_or2_1 _5028_ (.X(_1522_),
    .B(_1520_),
    .A(_1505_));
 sg13g2_and2_1 _5029_ (.A(\dtop.field_top.player.controller.pattern0[2] ),
    .B(_1522_),
    .X(_1523_));
 sg13g2_nand2b_2 _5030_ (.Y(_1524_),
    .B(_2830_),
    .A_N(_1518_));
 sg13g2_nor2_1 _5031_ (.A(net1022),
    .B(net1067),
    .Y(_1525_));
 sg13g2_nand2_2 _5032_ (.Y(_1526_),
    .A(net1064),
    .B(net1021));
 sg13g2_nand4_1 _5033_ (.B(_1505_),
    .C(_1514_),
    .A(net1029),
    .Y(_1527_),
    .D(_1526_));
 sg13g2_o21ai_1 _5034_ (.B1(_1527_),
    .Y(_1528_),
    .A1(_1510_),
    .A2(_1524_));
 sg13g2_nor4_1 _5035_ (.A(_1516_),
    .B(_1519_),
    .C(_1523_),
    .D(_1528_),
    .Y(_1529_));
 sg13g2_nand2_1 _5036_ (.Y(_1530_),
    .A(net1094),
    .B(\dtop.field_top.player.osc0[12] ));
 sg13g2_o21ai_1 _5037_ (.B1(net940),
    .Y(_1531_),
    .A1(_1529_),
    .A2(_1530_));
 sg13g2_a221oi_1 _5038_ (.B2(_1483_),
    .C1(\dtop.field_top.channel[2] ),
    .B1(_1491_),
    .A1(\dtop.field_top.channel[3] ),
    .Y(_1532_),
    .A2(_1489_));
 sg13g2_and3_2 _5039_ (.X(_1533_),
    .A(net1109),
    .B(_1501_),
    .C(_1532_));
 sg13g2_nand3_1 _5040_ (.B(_1501_),
    .C(_1532_),
    .A(net1109),
    .Y(_1534_));
 sg13g2_and2_1 _5041_ (.A(_0110_),
    .B(net985),
    .X(_1535_));
 sg13g2_a21o_1 _5042_ (.A2(_1492_),
    .A1(net988),
    .B1(_1535_),
    .X(_1536_));
 sg13g2_a221oi_1 _5043_ (.B2(net987),
    .C1(_1535_),
    .B1(_1492_),
    .A1(\dtop.field_top.channel[3] ),
    .Y(_1537_),
    .A2(_1489_));
 sg13g2_or2_1 _5044_ (.X(_1538_),
    .B(_1536_),
    .A(_1490_));
 sg13g2_nor2_2 _5045_ (.A(_1533_),
    .B(_1537_),
    .Y(_1539_));
 sg13g2_nand2_2 _5046_ (.Y(_1540_),
    .A(_1534_),
    .B(_1538_));
 sg13g2_mux2_1 _5047_ (.A0(_1509_),
    .A1(_1518_),
    .S(_2830_),
    .X(_1541_));
 sg13g2_mux2_1 _5048_ (.A0(\dtop.field_top.player.controller.pattern0[1] ),
    .A1(net1029),
    .S(net1061),
    .X(_1542_));
 sg13g2_a21oi_1 _5049_ (.A1(_1521_),
    .A2(_1541_),
    .Y(_1543_),
    .B1(_1542_));
 sg13g2_a21o_1 _5050_ (.A2(_1541_),
    .A1(_1521_),
    .B1(_1542_),
    .X(_1544_));
 sg13g2_nand2_1 _5051_ (.Y(_1545_),
    .A(\dtop.field_top.player.controller.ppos[4] ),
    .B(net972));
 sg13g2_nor2_2 _5052_ (.A(net1084),
    .B(net1089),
    .Y(_1546_));
 sg13g2_or2_2 _5053_ (.X(_1547_),
    .B(net1089),
    .A(net1084));
 sg13g2_and2_2 _5054_ (.A(net1076),
    .B(_1546_),
    .X(_1548_));
 sg13g2_nand2_1 _5055_ (.Y(_1549_),
    .A(net1076),
    .B(_1546_));
 sg13g2_nand2b_1 _5056_ (.Y(_1550_),
    .B(net1093),
    .A_N(net1090));
 sg13g2_nand3_1 _5057_ (.B(_1525_),
    .C(_1548_),
    .A(net1093),
    .Y(_1551_));
 sg13g2_nor2_2 _5058_ (.A(net1062),
    .B(net1021),
    .Y(_1552_));
 sg13g2_nand2b_1 _5059_ (.Y(_1553_),
    .B(net1068),
    .A_N(net1064));
 sg13g2_a21oi_1 _5060_ (.A1(_1548_),
    .A2(_1552_),
    .Y(_1554_),
    .B1(_1545_));
 sg13g2_nor2_2 _5061_ (.A(net1083),
    .B(net1088),
    .Y(_1555_));
 sg13g2_nand2_2 _5062_ (.Y(_1556_),
    .A(_2834_),
    .B(_2835_));
 sg13g2_nand2_1 _5063_ (.Y(_1557_),
    .A(\dtop.field_top.player.controller.ppos[4] ),
    .B(_1556_));
 sg13g2_a21oi_1 _5064_ (.A1(net1067),
    .A2(\dtop.field_top.player.controller.ppos[4] ),
    .Y(_1558_),
    .B1(net1063));
 sg13g2_and2_1 _5065_ (.A(_1557_),
    .B(_1558_),
    .X(_1559_));
 sg13g2_nor2_1 _5066_ (.A(net1067),
    .B(net1012),
    .Y(_1560_));
 sg13g2_a21oi_1 _5067_ (.A1(net1066),
    .A2(_1548_),
    .Y(_1561_),
    .B1(net1012));
 sg13g2_or3_2 _5068_ (.A(net1080),
    .B(net1084),
    .C(net1089),
    .X(_1562_));
 sg13g2_o21ai_1 _5069_ (.B1(net1063),
    .Y(_1563_),
    .A1(net1066),
    .A2(_1562_));
 sg13g2_o21ai_1 _5070_ (.B1(net976),
    .Y(_1564_),
    .A1(_1561_),
    .A2(_1563_));
 sg13g2_o21ai_1 _5071_ (.B1(_1539_),
    .Y(_1565_),
    .A1(_1559_),
    .A2(_1564_));
 sg13g2_a21oi_1 _5072_ (.A1(_1551_),
    .A2(_1554_),
    .Y(_1566_),
    .B1(_1565_));
 sg13g2_nor3_2 _5073_ (.A(_2835_),
    .B(_2836_),
    .C(net1076),
    .Y(_1567_));
 sg13g2_nand3b_1 _5074_ (.B(net1089),
    .C(net1084),
    .Y(_1568_),
    .A_N(net1076));
 sg13g2_nand3_1 _5075_ (.B(net1084),
    .C(net1089),
    .A(net1080),
    .Y(_1569_));
 sg13g2_nor2_1 _5076_ (.A(net1073),
    .B(_1555_),
    .Y(_1570_));
 sg13g2_nor2_1 _5077_ (.A(net1079),
    .B(_2835_),
    .Y(_1571_));
 sg13g2_a22oi_1 _5078_ (.Y(_1572_),
    .B1(_1569_),
    .B2(_1570_),
    .A2(_1567_),
    .A1(net1073));
 sg13g2_or2_1 _5079_ (.X(_1573_),
    .B(_1572_),
    .A(net1067));
 sg13g2_nor2_2 _5080_ (.A(net1021),
    .B(net1070),
    .Y(_1574_));
 sg13g2_nand2_2 _5081_ (.Y(_1575_),
    .A(net1066),
    .B(net1012));
 sg13g2_nor2_2 _5082_ (.A(net1091),
    .B(net1093),
    .Y(_1576_));
 sg13g2_nand2_2 _5083_ (.Y(_1577_),
    .A(_1555_),
    .B(_1576_));
 sg13g2_nand2_1 _5084_ (.Y(_1578_),
    .A(_1569_),
    .B(_1577_));
 sg13g2_nand2_1 _5085_ (.Y(_1579_),
    .A(_1574_),
    .B(_1578_));
 sg13g2_a21oi_1 _5086_ (.A1(_1573_),
    .A2(_1579_),
    .Y(_1580_),
    .B1(net1062));
 sg13g2_nor2_1 _5087_ (.A(net1067),
    .B(net1070),
    .Y(_1581_));
 sg13g2_nand2_1 _5088_ (.Y(_1582_),
    .A(net1021),
    .B(net1012));
 sg13g2_nor2b_2 _5089_ (.A(net1090),
    .B_N(net1086),
    .Y(_1583_));
 sg13g2_nor2b_2 _5090_ (.A(net1084),
    .B_N(net1090),
    .Y(_1584_));
 sg13g2_nor3_1 _5091_ (.A(_2837_),
    .B(_1583_),
    .C(_1584_),
    .Y(_1585_));
 sg13g2_o21ai_1 _5092_ (.B1(_1581_),
    .Y(_1586_),
    .A1(net1081),
    .A2(_1585_));
 sg13g2_xnor2_1 _5093_ (.Y(_1587_),
    .A(net1073),
    .B(_1568_));
 sg13g2_nand2_2 _5094_ (.Y(_1588_),
    .A(net1066),
    .B(_1587_));
 sg13g2_nand3_1 _5095_ (.B(_1586_),
    .C(_1588_),
    .A(net1062),
    .Y(_1589_));
 sg13g2_nand2b_1 _5096_ (.Y(_1590_),
    .B(_1589_),
    .A_N(_1580_));
 sg13g2_a21oi_2 _5097_ (.B1(net1073),
    .Y(_1591_),
    .A2(net1085),
    .A1(net1080));
 sg13g2_a21o_2 _5098_ (.A2(net1085),
    .A1(net1079),
    .B1(net1071),
    .X(_1592_));
 sg13g2_nor3_1 _5099_ (.A(net1069),
    .B(_1550_),
    .C(_1591_),
    .Y(_1593_));
 sg13g2_nor2_1 _5100_ (.A(net1019),
    .B(_2834_),
    .Y(_1594_));
 sg13g2_nand2_2 _5101_ (.Y(_1595_),
    .A(net1072),
    .B(net1079));
 sg13g2_and3_1 _5102_ (.X(_1596_),
    .A(net1071),
    .B(net1079),
    .C(net1084));
 sg13g2_nand3_1 _5103_ (.B(net1082),
    .C(net1087),
    .A(net1071),
    .Y(_1597_));
 sg13g2_nor2_1 _5104_ (.A(net1068),
    .B(_1596_),
    .Y(_1598_));
 sg13g2_nand2_1 _5105_ (.Y(_1599_),
    .A(_1592_),
    .B(_1597_));
 sg13g2_nor3_2 _5106_ (.A(net1066),
    .B(_1591_),
    .C(_1596_),
    .Y(_1600_));
 sg13g2_nor2_2 _5107_ (.A(_1593_),
    .B(_1600_),
    .Y(_1601_));
 sg13g2_nand3_1 _5108_ (.B(_1588_),
    .C(_1601_),
    .A(net973),
    .Y(_1602_));
 sg13g2_nand2_1 _5109_ (.Y(_1603_),
    .A(_1533_),
    .B(_1602_));
 sg13g2_a21oi_1 _5110_ (.A1(net977),
    .A2(_1590_),
    .Y(_1604_),
    .B1(_1603_));
 sg13g2_and3_2 _5111_ (.X(_1605_),
    .A(net1109),
    .B(_1501_),
    .C(_1537_));
 sg13g2_nor2_2 _5112_ (.A(net1063),
    .B(net974),
    .Y(_1606_));
 sg13g2_nand2_2 _5113_ (.Y(_1607_),
    .A(net1022),
    .B(net976));
 sg13g2_nor2_1 _5114_ (.A(_2836_),
    .B(net1093),
    .Y(_1608_));
 sg13g2_a21oi_2 _5115_ (.B1(net1080),
    .Y(_1609_),
    .A2(net1089),
    .A1(net1084));
 sg13g2_and2_1 _5116_ (.A(_1547_),
    .B(_1609_),
    .X(_1610_));
 sg13g2_nand2b_2 _5117_ (.Y(_1611_),
    .B(_1610_),
    .A_N(_1608_));
 sg13g2_nand2b_1 _5118_ (.Y(_1612_),
    .B(_2837_),
    .A_N(_1569_));
 sg13g2_a21oi_1 _5119_ (.A1(_1595_),
    .A2(_1612_),
    .Y(_1613_),
    .B1(net1068));
 sg13g2_a21oi_1 _5120_ (.A1(_1574_),
    .A2(_1611_),
    .Y(_1614_),
    .B1(_1613_));
 sg13g2_nor2_1 _5121_ (.A(_1607_),
    .B(_1614_),
    .Y(_1615_));
 sg13g2_nor2_2 _5122_ (.A(net1022),
    .B(net972),
    .Y(_1616_));
 sg13g2_nand3_1 _5123_ (.B(net1085),
    .C(_1581_),
    .A(net1081),
    .Y(_1617_));
 sg13g2_nand2_1 _5124_ (.Y(_1618_),
    .A(net1067),
    .B(net1074));
 sg13g2_o21ai_1 _5125_ (.B1(_1617_),
    .Y(_1619_),
    .A1(_1555_),
    .A2(_1618_));
 sg13g2_nor2_2 _5126_ (.A(net1065),
    .B(\dtop.field_top.player.controller.ppos[6] ),
    .Y(_1620_));
 sg13g2_o21ai_1 _5127_ (.B1(_1620_),
    .Y(_1621_),
    .A1(net1070),
    .A2(_1609_));
 sg13g2_a221oi_1 _5128_ (.B2(net972),
    .C1(_1615_),
    .B1(_1621_),
    .A1(_1616_),
    .Y(_1622_),
    .A2(_1619_));
 sg13g2_and2_1 _5129_ (.A(_1605_),
    .B(_1622_),
    .X(_1623_));
 sg13g2_a221oi_1 _5130_ (.B2(net1109),
    .C1(_1536_),
    .B1(_1501_),
    .A1(\dtop.field_top.channel[3] ),
    .Y(_1624_),
    .A2(_1489_));
 sg13g2_nand2b_1 _5131_ (.Y(_1625_),
    .B(_1537_),
    .A_N(net964));
 sg13g2_a21oi_1 _5132_ (.A1(_1592_),
    .A2(_1597_),
    .Y(_1626_),
    .B1(net1068));
 sg13g2_or2_2 _5133_ (.X(_1627_),
    .B(_1576_),
    .A(net1088));
 sg13g2_nor2_1 _5134_ (.A(net1077),
    .B(_1618_),
    .Y(_1628_));
 sg13g2_nor2_1 _5135_ (.A(_2832_),
    .B(net1075),
    .Y(_1629_));
 sg13g2_a221oi_1 _5136_ (.B2(net1077),
    .C1(_1626_),
    .B1(_1629_),
    .A1(_1627_),
    .Y(_1630_),
    .A2(_1628_));
 sg13g2_nand2_1 _5137_ (.Y(_1631_),
    .A(net1089),
    .B(_1595_));
 sg13g2_nor2_1 _5138_ (.A(_2835_),
    .B(_1511_),
    .Y(_1632_));
 sg13g2_a21oi_1 _5139_ (.A1(_1592_),
    .A2(_1597_),
    .Y(_1633_),
    .B1(_1553_));
 sg13g2_a21oi_1 _5140_ (.A1(_1631_),
    .A2(_1632_),
    .Y(_1634_),
    .B1(_1633_));
 sg13g2_o21ai_1 _5141_ (.B1(_1634_),
    .Y(_1635_),
    .A1(net1023),
    .A2(_1630_));
 sg13g2_and2_1 _5142_ (.A(net974),
    .B(_1635_),
    .X(_1636_));
 sg13g2_nand2_1 _5143_ (.Y(_1637_),
    .A(_1599_),
    .B(_1616_));
 sg13g2_o21ai_1 _5144_ (.B1(net1079),
    .Y(_1638_),
    .A1(_2855_),
    .A2(_1608_));
 sg13g2_nor2_2 _5145_ (.A(net1071),
    .B(net1076),
    .Y(_1639_));
 sg13g2_nand2_2 _5146_ (.Y(_1640_),
    .A(_1547_),
    .B(_1639_));
 sg13g2_nand2_1 _5147_ (.Y(_1641_),
    .A(net1068),
    .B(_1640_));
 sg13g2_a21o_1 _5148_ (.A2(_1638_),
    .A1(net1072),
    .B1(_1641_),
    .X(_1642_));
 sg13g2_nand2b_1 _5149_ (.Y(_1643_),
    .B(_1642_),
    .A_N(_1626_));
 sg13g2_nand2_1 _5150_ (.Y(_1644_),
    .A(_1606_),
    .B(_1643_));
 sg13g2_a21oi_1 _5151_ (.A1(_1555_),
    .A2(_1642_),
    .Y(_1645_),
    .B1(_1644_));
 sg13g2_o21ai_1 _5152_ (.B1(_1624_),
    .Y(_1646_),
    .A1(_1593_),
    .A2(_1637_));
 sg13g2_nor3_1 _5153_ (.A(_1636_),
    .B(_1645_),
    .C(_1646_),
    .Y(_1647_));
 sg13g2_nor4_2 _5154_ (.A(_1566_),
    .B(_1604_),
    .C(_1623_),
    .Y(_1648_),
    .D(_1647_));
 sg13g2_nor2b_1 _5155_ (.A(net964),
    .B_N(_1532_),
    .Y(_1649_));
 sg13g2_a21oi_1 _5156_ (.A1(net1029),
    .A2(\dtop.field_top.player.controller.pattern0[2] ),
    .Y(_1650_),
    .B1(_1509_));
 sg13g2_a221oi_1 _5157_ (.B2(_1522_),
    .C1(_1650_),
    .B1(\dtop.field_top.player.controller.pattern0[2] ),
    .A1(net1029),
    .Y(_1651_),
    .A2(net1061));
 sg13g2_o21ai_1 _5158_ (.B1(_1513_),
    .Y(_1652_),
    .A1(net1069),
    .A2(_1515_));
 sg13g2_and4_2 _5159_ (.A(_1541_),
    .B(_1649_),
    .C(_1651_),
    .D(_1652_),
    .X(_1653_));
 sg13g2_nand4_1 _5160_ (.B(_1649_),
    .C(_1651_),
    .A(_1541_),
    .Y(_1654_),
    .D(_1652_));
 sg13g2_nor3_1 _5161_ (.A(_1513_),
    .B(_1524_),
    .C(_1577_),
    .Y(_1655_));
 sg13g2_o21ai_1 _5162_ (.B1(_1522_),
    .Y(_1656_),
    .A1(net1029),
    .A2(_1506_));
 sg13g2_inv_1 _5163_ (.Y(_1657_),
    .A(_1656_));
 sg13g2_nor4_1 _5164_ (.A(_1648_),
    .B(_1653_),
    .C(_1655_),
    .D(_1657_),
    .Y(_1658_));
 sg13g2_nor2_2 _5165_ (.A(_1494_),
    .B(net964),
    .Y(_1659_));
 sg13g2_nand2_1 _5166_ (.Y(_1660_),
    .A(net1024),
    .B(_1514_));
 sg13g2_a21oi_1 _5167_ (.A1(_1576_),
    .A2(_1660_),
    .Y(_1661_),
    .B1(_1654_));
 sg13g2_nor3_1 _5168_ (.A(_1658_),
    .B(_1659_),
    .C(_1661_),
    .Y(_1662_));
 sg13g2_nor4_2 _5169_ (.A(net1034),
    .B(_1213_),
    .C(_1337_),
    .Y(_1663_),
    .D(_1497_));
 sg13g2_o21ai_1 _5170_ (.B1(\dtop.field_top.channel[0] ),
    .Y(_1664_),
    .A1(net986),
    .A2(_1663_));
 sg13g2_nand2_1 _5171_ (.Y(_1665_),
    .A(_1659_),
    .B(_1664_));
 sg13g2_a21oi_1 _5172_ (.A1(_1510_),
    .A2(_1522_),
    .Y(_1666_),
    .B1(_1506_));
 sg13g2_nor4_1 _5173_ (.A(\dtop.field_top.player.osc0[22] ),
    .B(net988),
    .C(net942),
    .D(_1666_),
    .Y(_1667_));
 sg13g2_nor3_2 _5174_ (.A(_1494_),
    .B(net964),
    .C(_1664_),
    .Y(_1668_));
 sg13g2_nand2_2 _5175_ (.Y(_1669_),
    .A(_1659_),
    .B(net942));
 sg13g2_nand4_1 _5176_ (.B(_1524_),
    .C(_1526_),
    .A(_1514_),
    .Y(_1670_),
    .D(_1651_));
 sg13g2_a22oi_1 _5177_ (.Y(_1671_),
    .B1(_1520_),
    .B2(\dtop.field_top.player.controller.pattern0[2] ),
    .A2(_1508_),
    .A1(_2830_));
 sg13g2_o21ai_1 _5178_ (.B1(_1521_),
    .Y(_1672_),
    .A1(net1029),
    .A2(_1509_));
 sg13g2_o21ai_1 _5179_ (.B1(_1670_),
    .Y(_1673_),
    .A1(net1024),
    .A2(_1524_));
 sg13g2_nor3_1 _5180_ (.A(net938),
    .B(_1672_),
    .C(_1673_),
    .Y(_1674_));
 sg13g2_nor3_1 _5181_ (.A(_1662_),
    .B(_1667_),
    .C(_1674_),
    .Y(_1675_));
 sg13g2_o21ai_1 _5182_ (.B1(_1531_),
    .Y(_1676_),
    .A1(net951),
    .A2(_1675_));
 sg13g2_nor2_2 _5183_ (.A(net2),
    .B(_3002_),
    .Y(_1677_));
 sg13g2_or2_1 _5184_ (.X(_1678_),
    .B(_3002_),
    .A(net2));
 sg13g2_a21oi_2 _5185_ (.B1(net965),
    .Y(_1679_),
    .A2(_1664_),
    .A1(_1659_));
 sg13g2_nand2_2 _5186_ (.Y(_1680_),
    .A(net941),
    .B(_1677_));
 sg13g2_a21oi_2 _5187_ (.B1(_1651_),
    .Y(_1681_),
    .A2(_1649_),
    .A1(_1519_));
 sg13g2_nor2_2 _5188_ (.A(net1104),
    .B(net1100),
    .Y(_1682_));
 sg13g2_or2_2 _5189_ (.X(_1683_),
    .B(net1101),
    .A(net1103));
 sg13g2_nand2_1 _5190_ (.Y(_1684_),
    .A(net1107),
    .B(_1682_));
 sg13g2_nand3_1 _5191_ (.B(net1009),
    .C(_1682_),
    .A(net1107),
    .Y(_1685_));
 sg13g2_nand2_1 _5192_ (.Y(_1686_),
    .A(net1100),
    .B(_3020_));
 sg13g2_nand2_1 _5193_ (.Y(_1687_),
    .A(_1685_),
    .B(_1686_));
 sg13g2_nand2_1 _5194_ (.Y(_1688_),
    .A(_3016_),
    .B(_1682_));
 sg13g2_nor2_1 _5195_ (.A(_2856_),
    .B(net1100),
    .Y(_1689_));
 sg13g2_nand2b_1 _5196_ (.Y(_1690_),
    .B(net1103),
    .A_N(net1099));
 sg13g2_nor2_1 _5197_ (.A(net1105),
    .B(_1690_),
    .Y(_1691_));
 sg13g2_nand2_1 _5198_ (.Y(_1692_),
    .A(net1009),
    .B(_1689_));
 sg13g2_nand3_1 _5199_ (.B(_1686_),
    .C(_1692_),
    .A(_1684_),
    .Y(_1693_));
 sg13g2_nor2_2 _5200_ (.A(net1108),
    .B(net1105),
    .Y(_1694_));
 sg13g2_nand2_2 _5201_ (.Y(_1695_),
    .A(_2839_),
    .B(net1009));
 sg13g2_nor2_2 _5202_ (.A(_1683_),
    .B(_1694_),
    .Y(_1696_));
 sg13g2_nor2b_1 _5203_ (.A(_0111_),
    .B_N(_0113_),
    .Y(_1697_));
 sg13g2_o21ai_1 _5204_ (.B1(_1683_),
    .Y(_1698_),
    .A1(_0114_),
    .A2(_3018_));
 sg13g2_a21oi_2 _5205_ (.B1(_1693_),
    .Y(_1699_),
    .A2(_1696_),
    .A1(_3017_));
 sg13g2_o21ai_1 _5206_ (.B1(net1097),
    .Y(_1700_),
    .A1(_1696_),
    .A2(_1699_));
 sg13g2_o21ai_1 _5207_ (.B1(_1700_),
    .Y(_1701_),
    .A1(net1098),
    .A2(_1698_));
 sg13g2_nand4_1 _5208_ (.B(_1681_),
    .C(_1697_),
    .A(_1494_),
    .Y(_1702_),
    .D(_1701_));
 sg13g2_nor4_1 _5209_ (.A(net1099),
    .B(_0111_),
    .C(_0112_),
    .D(_3015_),
    .Y(_1703_));
 sg13g2_nand2_1 _5210_ (.Y(_1704_),
    .A(_1677_),
    .B(_1703_));
 sg13g2_nand2b_1 _5211_ (.Y(_1705_),
    .B(net1107),
    .A_N(net1095));
 sg13g2_a21o_1 _5212_ (.A2(_1682_),
    .A1(net1009),
    .B1(_1705_),
    .X(_1706_));
 sg13g2_a21oi_2 _5213_ (.B1(net1100),
    .Y(_1707_),
    .A2(net1105),
    .A1(net1103));
 sg13g2_nand2_1 _5214_ (.Y(_1708_),
    .A(net1095),
    .B(_1707_));
 sg13g2_nand2_1 _5215_ (.Y(_1709_),
    .A(net1026),
    .B(_1695_));
 sg13g2_a221oi_1 _5216_ (.B2(_1708_),
    .C1(_1709_),
    .B1(_1706_),
    .A1(\dtop.field_top.player.sched.alu.p0 ),
    .Y(_1710_),
    .A2(_1704_));
 sg13g2_o21ai_1 _5217_ (.B1(_1710_),
    .Y(_1711_),
    .A1(\dtop.field_top.player.sched.alu.p0 ),
    .A2(_1704_));
 sg13g2_nand3_1 _5218_ (.B(_3024_),
    .C(net944),
    .A(net1010),
    .Y(_1712_));
 sg13g2_o21ai_1 _5219_ (.B1(_1711_),
    .Y(_1713_),
    .A1(net1028),
    .A2(_1712_));
 sg13g2_nand2b_1 _5220_ (.Y(_1714_),
    .B(_1702_),
    .A_N(_1713_));
 sg13g2_a22oi_1 _5221_ (.Y(_1715_),
    .B1(_1679_),
    .B2(_1714_),
    .A2(_1676_),
    .A1(_3003_));
 sg13g2_nand2b_2 _5222_ (.Y(_1716_),
    .B(net1120),
    .A_N(_1715_));
 sg13g2_nor2_1 _5223_ (.A(net1117),
    .B(net1),
    .Y(_1717_));
 sg13g2_a21oi_1 _5224_ (.A1(net1117),
    .A2(_3015_),
    .Y(_1718_),
    .B1(_1717_));
 sg13g2_and2_1 _5225_ (.A(net965),
    .B(_1718_),
    .X(_1719_));
 sg13g2_inv_1 _5226_ (.Y(_1720_),
    .A(_1719_));
 sg13g2_nand2_1 _5227_ (.Y(_1721_),
    .A(_1716_),
    .B(_1719_));
 sg13g2_nor2_2 _5228_ (.A(net1099),
    .B(net1096),
    .Y(_1722_));
 sg13g2_and2_1 _5229_ (.A(_0111_),
    .B(_1722_),
    .X(_1723_));
 sg13g2_nand2_1 _5230_ (.Y(_1724_),
    .A(_0111_),
    .B(_1722_));
 sg13g2_nor2_2 _5231_ (.A(net1009),
    .B(_3001_),
    .Y(_1725_));
 sg13g2_nor2_2 _5232_ (.A(net1108),
    .B(_1725_),
    .Y(_1726_));
 sg13g2_o21ai_1 _5233_ (.B1(_1668_),
    .Y(_1727_),
    .A1(_1723_),
    .A2(_1726_));
 sg13g2_or2_1 _5234_ (.X(_1728_),
    .B(_1727_),
    .A(_3022_));
 sg13g2_nand3b_1 _5235_ (.B(net1011),
    .C(_1677_),
    .Y(_1729_),
    .A_N(_1728_));
 sg13g2_nor2_1 _5236_ (.A(_1511_),
    .B(net982),
    .Y(_1730_));
 sg13g2_a21o_1 _5237_ (.A2(_1730_),
    .A1(_1557_),
    .B1(net975),
    .X(_1731_));
 sg13g2_nand3_1 _5238_ (.B(_1548_),
    .C(_1560_),
    .A(net1093),
    .Y(_1732_));
 sg13g2_o21ai_1 _5239_ (.B1(net972),
    .Y(_1733_),
    .A1(\dtop.field_top.player.controller.ppos[6] ),
    .A2(_1732_));
 sg13g2_nand2_1 _5240_ (.Y(_1734_),
    .A(_1731_),
    .B(_1733_));
 sg13g2_nand3_1 _5241_ (.B(_1538_),
    .C(_1734_),
    .A(_1534_),
    .Y(_1735_));
 sg13g2_a21oi_2 _5242_ (.B1(_1582_),
    .Y(_1736_),
    .A2(_1547_),
    .A1(net1081));
 sg13g2_a21oi_2 _5243_ (.B1(_1586_),
    .Y(_1737_),
    .A2(_1547_),
    .A1(net1081));
 sg13g2_a22oi_1 _5244_ (.Y(_1738_),
    .B1(_1737_),
    .B2(_1616_),
    .A2(_1629_),
    .A1(_1606_));
 sg13g2_a221oi_1 _5245_ (.B2(net1087),
    .C1(net1069),
    .B1(_1594_),
    .A1(_1556_),
    .Y(_1739_),
    .A2(_1591_));
 sg13g2_or2_1 _5246_ (.X(_1740_),
    .B(_1739_),
    .A(net1063));
 sg13g2_nand2_1 _5247_ (.Y(_1741_),
    .A(net1089),
    .B(net1093));
 sg13g2_or2_1 _5248_ (.X(_1742_),
    .B(net1070),
    .A(net1076));
 sg13g2_nor4_1 _5249_ (.A(_2832_),
    .B(net1087),
    .C(_1741_),
    .D(_1742_),
    .Y(_1743_));
 sg13g2_o21ai_1 _5250_ (.B1(net1064),
    .Y(_1744_),
    .A1(net1065),
    .A2(_1599_));
 sg13g2_or3_1 _5251_ (.A(net974),
    .B(_1740_),
    .C(_1743_),
    .X(_1745_));
 sg13g2_o21ai_1 _5252_ (.B1(_1745_),
    .Y(_1746_),
    .A1(net974),
    .A2(_1744_));
 sg13g2_nor3_1 _5253_ (.A(_1625_),
    .B(_1636_),
    .C(_1746_),
    .Y(_1747_));
 sg13g2_o21ai_1 _5254_ (.B1(_1540_),
    .Y(_1748_),
    .A1(_1534_),
    .A2(_1738_));
 sg13g2_or2_1 _5255_ (.X(_1749_),
    .B(_1748_),
    .A(_1605_));
 sg13g2_o21ai_1 _5256_ (.B1(_1735_),
    .Y(_1750_),
    .A1(_1747_),
    .A2(_1749_));
 sg13g2_o21ai_1 _5257_ (.B1(net1073),
    .Y(_1751_),
    .A1(net1076),
    .A2(_1546_));
 sg13g2_a21o_1 _5258_ (.A2(_1751_),
    .A1(_1640_),
    .B1(net1065),
    .X(_1752_));
 sg13g2_mux2_1 _5259_ (.A0(_1601_),
    .A1(_1752_),
    .S(net1023),
    .X(_1753_));
 sg13g2_nor3_1 _5260_ (.A(net964),
    .B(_1538_),
    .C(_1753_),
    .Y(_1754_));
 sg13g2_nor3_2 _5261_ (.A(net1019),
    .B(_1555_),
    .C(net983),
    .Y(_1755_));
 sg13g2_nand2_1 _5262_ (.Y(_1756_),
    .A(_1510_),
    .B(_1595_));
 sg13g2_nand3_1 _5263_ (.B(net1088),
    .C(_1741_),
    .A(net1083),
    .Y(_1757_));
 sg13g2_nand2b_1 _5264_ (.Y(_1758_),
    .B(_1757_),
    .A_N(_1756_));
 sg13g2_nor2_1 _5265_ (.A(_1755_),
    .B(_1758_),
    .Y(_1759_));
 sg13g2_a21oi_1 _5266_ (.A1(_1605_),
    .A2(_1759_),
    .Y(_1760_),
    .B1(_1754_));
 sg13g2_nor3_1 _5267_ (.A(net1081),
    .B(\dtop.field_top.player.controller.ppos[6] ),
    .C(_1582_),
    .Y(_1761_));
 sg13g2_o21ai_1 _5268_ (.B1(_1601_),
    .Y(_1762_),
    .A1(net1062),
    .A2(_1588_));
 sg13g2_nand2_1 _5269_ (.Y(_1763_),
    .A(net973),
    .B(_1762_));
 sg13g2_nand3_1 _5270_ (.B(_1585_),
    .C(_1761_),
    .A(net976),
    .Y(_1764_));
 sg13g2_nand2_1 _5271_ (.Y(_1765_),
    .A(_1763_),
    .B(_1764_));
 sg13g2_a21oi_1 _5272_ (.A1(_1533_),
    .A2(_1765_),
    .Y(_1766_),
    .B1(_1539_));
 sg13g2_o21ai_1 _5273_ (.B1(_1766_),
    .Y(_1767_),
    .A1(net974),
    .A2(_1760_));
 sg13g2_and2_1 _5274_ (.A(_1735_),
    .B(_1767_),
    .X(_1768_));
 sg13g2_nor2_1 _5275_ (.A(net1029),
    .B(_1523_),
    .Y(_1769_));
 sg13g2_nand2b_2 _5276_ (.Y(_1770_),
    .B(_2830_),
    .A_N(_1523_));
 sg13g2_nand3_1 _5277_ (.B(net976),
    .C(_1588_),
    .A(net1062),
    .Y(_1771_));
 sg13g2_a21oi_1 _5278_ (.A1(_2832_),
    .A2(_1594_),
    .Y(_1772_),
    .B1(_1771_));
 sg13g2_nand2_1 _5279_ (.Y(_1773_),
    .A(_2853_),
    .B(_1587_));
 sg13g2_nand2_1 _5280_ (.Y(_1774_),
    .A(_1587_),
    .B(_1620_));
 sg13g2_and2_1 _5281_ (.A(net973),
    .B(_1774_),
    .X(_1775_));
 sg13g2_nor3_1 _5282_ (.A(_1534_),
    .B(_1772_),
    .C(_1775_),
    .Y(_1776_));
 sg13g2_a21oi_1 _5283_ (.A1(_1525_),
    .A2(_1547_),
    .Y(_1777_),
    .B1(_1580_));
 sg13g2_o21ai_1 _5284_ (.B1(_1776_),
    .Y(_1778_),
    .A1(net973),
    .A2(_1777_));
 sg13g2_nand4_1 _5285_ (.B(_1597_),
    .C(_1620_),
    .A(_1592_),
    .Y(_1779_),
    .D(net984));
 sg13g2_nand3_1 _5286_ (.B(_1740_),
    .C(_1744_),
    .A(net983),
    .Y(_1780_));
 sg13g2_nand3_1 _5287_ (.B(_1779_),
    .C(_1780_),
    .A(net978),
    .Y(_1781_));
 sg13g2_nand2_1 _5288_ (.Y(_1782_),
    .A(net975),
    .B(net984));
 sg13g2_nor3_1 _5289_ (.A(net1065),
    .B(_1627_),
    .C(_1742_),
    .Y(_1783_));
 sg13g2_nand2b_1 _5290_ (.Y(_1784_),
    .B(net1063),
    .A_N(_1783_));
 sg13g2_a21o_2 _5291_ (.A2(net1085),
    .A1(net1080),
    .B1(_1609_),
    .X(_1785_));
 sg13g2_nor2_1 _5292_ (.A(net1019),
    .B(_1511_),
    .Y(_1786_));
 sg13g2_nand2_1 _5293_ (.Y(_1787_),
    .A(net1075),
    .B(_1510_));
 sg13g2_o21ai_1 _5294_ (.B1(net1087),
    .Y(_1788_),
    .A1(net1079),
    .A2(\dtop.field_top.player.controller.ppos[1] ));
 sg13g2_o21ai_1 _5295_ (.B1(_1788_),
    .Y(_1789_),
    .A1(_1550_),
    .A2(_1556_));
 sg13g2_a221oi_1 _5296_ (.B2(_1512_),
    .C1(_1633_),
    .B1(_1789_),
    .A1(_1785_),
    .Y(_1790_),
    .A2(_1786_));
 sg13g2_nor2_2 _5297_ (.A(net978),
    .B(net984),
    .Y(_1791_));
 sg13g2_inv_1 _5298_ (.Y(_1792_),
    .A(_1791_));
 sg13g2_nand3_1 _5299_ (.B(_1784_),
    .C(_1790_),
    .A(net983),
    .Y(_1793_));
 sg13g2_o21ai_1 _5300_ (.B1(_1793_),
    .Y(_1794_),
    .A1(_1636_),
    .A2(_1791_));
 sg13g2_nand3_1 _5301_ (.B(_1781_),
    .C(_1794_),
    .A(_1624_),
    .Y(_1795_));
 sg13g2_and2_2 _5302_ (.A(net978),
    .B(_1605_),
    .X(_1796_));
 sg13g2_a22oi_1 _5303_ (.Y(_1797_),
    .B1(_1611_),
    .B2(net1071),
    .A2(_1584_),
    .A1(net1080));
 sg13g2_nand2b_1 _5304_ (.Y(_1798_),
    .B(_1552_),
    .A_N(_1797_));
 sg13g2_o21ai_1 _5305_ (.B1(_1574_),
    .Y(_1799_),
    .A1(net1080),
    .A2(_1627_));
 sg13g2_a21oi_1 _5306_ (.A1(_1617_),
    .A2(_1799_),
    .Y(_1800_),
    .B1(net1022));
 sg13g2_nand2_1 _5307_ (.Y(_1801_),
    .A(_1583_),
    .B(_1639_));
 sg13g2_a21oi_1 _5308_ (.A1(net1071),
    .A2(_1571_),
    .Y(_1802_),
    .B1(_1511_));
 sg13g2_a221oi_1 _5309_ (.B2(_1802_),
    .C1(_1800_),
    .B1(_1801_),
    .A1(net982),
    .Y(_1803_),
    .A2(_1786_));
 sg13g2_nand3_1 _5310_ (.B(_1798_),
    .C(_1803_),
    .A(_1796_),
    .Y(_1804_));
 sg13g2_nand3_1 _5311_ (.B(_1795_),
    .C(_1804_),
    .A(_1778_),
    .Y(_1805_));
 sg13g2_a21oi_1 _5312_ (.A1(\dtop.field_top.player.controller.ppos[2] ),
    .A2(_1514_),
    .Y(_1806_),
    .B1(_1756_));
 sg13g2_o21ai_1 _5313_ (.B1(_1806_),
    .Y(_1807_),
    .A1(net1075),
    .A2(_1569_));
 sg13g2_a21oi_1 _5314_ (.A1(net1075),
    .A2(_1546_),
    .Y(_1808_),
    .B1(_1807_));
 sg13g2_nor2_1 _5315_ (.A(net983),
    .B(_1758_),
    .Y(_1809_));
 sg13g2_o21ai_1 _5316_ (.B1(_1796_),
    .Y(_1810_),
    .A1(_1808_),
    .A2(_1809_));
 sg13g2_a221oi_1 _5317_ (.B2(_1570_),
    .C1(net1066),
    .B1(_1569_),
    .A1(net1073),
    .Y(_1811_),
    .A2(_1567_));
 sg13g2_nand2_1 _5318_ (.Y(_1812_),
    .A(_1562_),
    .B(_1569_));
 sg13g2_nor2_1 _5319_ (.A(_1575_),
    .B(_1812_),
    .Y(_1813_));
 sg13g2_nor3_2 _5320_ (.A(net1062),
    .B(_1811_),
    .C(_1813_),
    .Y(_1814_));
 sg13g2_o21ai_1 _5321_ (.B1(net977),
    .Y(_1815_),
    .A1(_1730_),
    .A2(_1814_));
 sg13g2_or2_1 _5322_ (.X(_1816_),
    .B(_1771_),
    .A(_1737_));
 sg13g2_and4_1 _5323_ (.A(net973),
    .B(_1588_),
    .C(_1601_),
    .D(net984),
    .X(_1817_));
 sg13g2_a21oi_1 _5324_ (.A1(_1774_),
    .A2(_1791_),
    .Y(_1818_),
    .B1(_1817_));
 sg13g2_and4_1 _5325_ (.A(_1533_),
    .B(_1815_),
    .C(_1816_),
    .D(_1818_),
    .X(_1819_));
 sg13g2_a21o_1 _5326_ (.A2(_1790_),
    .A1(_1784_),
    .B1(_1782_),
    .X(_1820_));
 sg13g2_a22oi_1 _5327_ (.Y(_1821_),
    .B1(_1791_),
    .B2(_1635_),
    .A2(_1753_),
    .A1(net978));
 sg13g2_and3_1 _5328_ (.X(_1822_),
    .A(_1624_),
    .B(_1820_),
    .C(_1821_));
 sg13g2_nor3_1 _5329_ (.A(_1539_),
    .B(_1819_),
    .C(_1822_),
    .Y(_1823_));
 sg13g2_o21ai_1 _5330_ (.B1(_1735_),
    .Y(_1824_),
    .A1(_1540_),
    .A2(_1792_));
 sg13g2_a21oi_1 _5331_ (.A1(_1810_),
    .A2(_1823_),
    .Y(_1825_),
    .B1(_1824_));
 sg13g2_nand2_1 _5332_ (.Y(_1826_),
    .A(net974),
    .B(_1787_));
 sg13g2_nand3_1 _5333_ (.B(_1731_),
    .C(_1826_),
    .A(_1539_),
    .Y(_1827_));
 sg13g2_or3_1 _5334_ (.A(\dtop.field_top.player.controller.ppos[2] ),
    .B(_1608_),
    .C(net984),
    .X(_1828_));
 sg13g2_a21oi_1 _5335_ (.A1(_1583_),
    .A2(net984),
    .Y(_1829_),
    .B1(_2834_));
 sg13g2_a22oi_1 _5336_ (.Y(_1830_),
    .B1(_1828_),
    .B2(_1829_),
    .A2(_1571_),
    .A1(net1019));
 sg13g2_a22oi_1 _5337_ (.Y(_1831_),
    .B1(_1639_),
    .B2(_1584_),
    .A2(_1595_),
    .A1(net1021));
 sg13g2_nor3_1 _5338_ (.A(net1019),
    .B(net1086),
    .C(net982),
    .Y(_1832_));
 sg13g2_nor2_1 _5339_ (.A(_1831_),
    .B(_1832_),
    .Y(_1833_));
 sg13g2_o21ai_1 _5340_ (.B1(_1833_),
    .Y(_1834_),
    .A1(net1068),
    .A2(_1830_));
 sg13g2_nor2_1 _5341_ (.A(net1070),
    .B(_1577_),
    .Y(_1835_));
 sg13g2_o21ai_1 _5342_ (.B1(_1617_),
    .Y(_1836_),
    .A1(net1021),
    .A2(_1835_));
 sg13g2_o21ai_1 _5343_ (.B1(_1620_),
    .Y(_1837_),
    .A1(net1070),
    .A2(_1610_));
 sg13g2_and2_1 _5344_ (.A(net972),
    .B(_1837_),
    .X(_1838_));
 sg13g2_a221oi_1 _5345_ (.B2(_1616_),
    .C1(_1838_),
    .B1(_1836_),
    .A1(_1606_),
    .Y(_1839_),
    .A2(_1834_));
 sg13g2_a21oi_1 _5346_ (.A1(_1640_),
    .A2(_1751_),
    .Y(_1840_),
    .B1(net1021));
 sg13g2_nor2_1 _5347_ (.A(_1739_),
    .B(_1840_),
    .Y(_1841_));
 sg13g2_mux2_1 _5348_ (.A0(_1752_),
    .A1(_1841_),
    .S(_1671_),
    .X(_1842_));
 sg13g2_nand2b_1 _5349_ (.Y(_1843_),
    .B(net1087),
    .A_N(\dtop.field_top.player.controller.ppos[1] ));
 sg13g2_a21oi_1 _5350_ (.A1(net1093),
    .A2(_1546_),
    .Y(_1844_),
    .B1(net1079));
 sg13g2_o21ai_1 _5351_ (.B1(_2834_),
    .Y(_1845_),
    .A1(_2837_),
    .A2(_1547_));
 sg13g2_a221oi_1 _5352_ (.B2(_1844_),
    .C1(_1513_),
    .B1(_1843_),
    .A1(net1079),
    .Y(_1846_),
    .A2(_1583_));
 sg13g2_nand3_1 _5353_ (.B(_1515_),
    .C(_1595_),
    .A(net1064),
    .Y(_1847_));
 sg13g2_a21oi_1 _5354_ (.A1(_1526_),
    .A2(_1847_),
    .Y(_1848_),
    .B1(_1626_));
 sg13g2_o21ai_1 _5355_ (.B1(net982),
    .Y(_1849_),
    .A1(_1846_),
    .A2(_1848_));
 sg13g2_nand2_1 _5356_ (.Y(_1850_),
    .A(net1022),
    .B(net1065));
 sg13g2_nor4_1 _5357_ (.A(net1012),
    .B(net983),
    .C(_1785_),
    .D(_1850_),
    .Y(_1851_));
 sg13g2_nor3_1 _5358_ (.A(_1556_),
    .B(_1671_),
    .C(_1787_),
    .Y(_1852_));
 sg13g2_nor3_1 _5359_ (.A(net977),
    .B(_1851_),
    .C(_1852_),
    .Y(_1853_));
 sg13g2_a221oi_1 _5360_ (.B2(_1853_),
    .C1(_1616_),
    .B1(_1849_),
    .A1(net977),
    .Y(_1854_),
    .A2(_1842_));
 sg13g2_nand2_1 _5361_ (.Y(_1855_),
    .A(_1574_),
    .B(_1812_));
 sg13g2_a21oi_2 _5362_ (.B1(_1607_),
    .Y(_1856_),
    .A2(_1855_),
    .A1(_1573_));
 sg13g2_nor4_1 _5363_ (.A(_1534_),
    .B(_1772_),
    .C(_1775_),
    .D(_1856_),
    .Y(_1857_));
 sg13g2_a221oi_1 _5364_ (.B2(_1624_),
    .C1(_1857_),
    .B1(_1854_),
    .A1(_1605_),
    .Y(_1858_),
    .A2(_1839_));
 sg13g2_nand2_1 _5365_ (.Y(_1859_),
    .A(_1827_),
    .B(_1858_));
 sg13g2_a221oi_1 _5366_ (.B2(_1858_),
    .C1(_1824_),
    .B1(_1827_),
    .A1(_1810_),
    .Y(_1860_),
    .A2(_1823_));
 sg13g2_nand2_1 _5367_ (.Y(_1861_),
    .A(_1805_),
    .B(_1860_));
 sg13g2_nand2_1 _5368_ (.Y(_1862_),
    .A(_1769_),
    .B(_1861_));
 sg13g2_a221oi_1 _5369_ (.B2(_1860_),
    .C1(_1770_),
    .B1(_1805_),
    .A1(_1735_),
    .Y(_1863_),
    .A2(_1767_));
 sg13g2_xor2_1 _5370_ (.B(_1863_),
    .A(_1750_),
    .X(_1864_));
 sg13g2_nand2_1 _5371_ (.Y(_1865_),
    .A(net943),
    .B(net938));
 sg13g2_nor2_2 _5372_ (.A(net951),
    .B(net950),
    .Y(_1866_));
 sg13g2_nand2_2 _5373_ (.Y(_1867_),
    .A(net946),
    .B(net938));
 sg13g2_a21oi_1 _5374_ (.A1(net1092),
    .A2(net950),
    .Y(_1868_),
    .B1(net951));
 sg13g2_o21ai_1 _5375_ (.B1(_1868_),
    .Y(_1869_),
    .A1(_1864_),
    .A2(_1865_));
 sg13g2_or2_2 _5376_ (.X(_1870_),
    .B(_1869_),
    .A(_0007_));
 sg13g2_nand3_1 _5377_ (.B(_1552_),
    .C(net984),
    .A(net1073),
    .Y(_1871_));
 sg13g2_a21oi_1 _5378_ (.A1(_1559_),
    .A2(net982),
    .Y(_1872_),
    .B1(_1564_));
 sg13g2_nand2_1 _5379_ (.Y(_1873_),
    .A(_1871_),
    .B(_1872_));
 sg13g2_a21oi_1 _5380_ (.A1(net1062),
    .A2(net1073),
    .Y(_1874_),
    .B1(net976));
 sg13g2_o21ai_1 _5381_ (.B1(_1874_),
    .Y(_1875_),
    .A1(net1063),
    .A2(_1561_));
 sg13g2_a21oi_2 _5382_ (.B1(_1540_),
    .Y(_1876_),
    .A2(_1875_),
    .A1(_1873_));
 sg13g2_nand3_1 _5383_ (.B(_1863_),
    .C(_1876_),
    .A(_1750_),
    .Y(_1877_));
 sg13g2_a21o_1 _5384_ (.A2(_1863_),
    .A1(_1750_),
    .B1(_1876_),
    .X(_1878_));
 sg13g2_nand3_1 _5385_ (.B(_1877_),
    .C(_1878_),
    .A(net943),
    .Y(_1879_));
 sg13g2_a21oi_2 _5386_ (.B1(net951),
    .Y(_1880_),
    .A2(_1879_),
    .A1(net938));
 sg13g2_xnor2_1 _5387_ (.Y(_1881_),
    .A(net1104),
    .B(_1880_));
 sg13g2_a221oi_1 _5388_ (.B2(_1879_),
    .C1(_0115_),
    .B1(_1669_),
    .A1(_1495_),
    .Y(_1882_),
    .A2(net964));
 sg13g2_o21ai_1 _5389_ (.B1(_1866_),
    .Y(_1883_),
    .A1(_1653_),
    .A2(_1877_));
 sg13g2_xnor2_1 _5390_ (.Y(_1884_),
    .A(net1102),
    .B(_1883_));
 sg13g2_nor2b_1 _5391_ (.A(_1884_),
    .B_N(_1882_),
    .Y(_1885_));
 sg13g2_xor2_1 _5392_ (.B(_1884_),
    .A(_1882_),
    .X(_1886_));
 sg13g2_o21ai_1 _5393_ (.B1(_1886_),
    .Y(_1887_),
    .A1(_1870_),
    .A2(_1881_));
 sg13g2_nor3_1 _5394_ (.A(_1870_),
    .B(_1881_),
    .C(_1886_),
    .Y(_1888_));
 sg13g2_nor2_1 _5395_ (.A(net981),
    .B(_1888_),
    .Y(_1889_));
 sg13g2_o21ai_1 _5396_ (.B1(net945),
    .Y(_1890_),
    .A1(_1723_),
    .A2(_1726_));
 sg13g2_nor3_1 _5397_ (.A(net1027),
    .B(net937),
    .C(_1890_),
    .Y(_1891_));
 sg13g2_a21oi_1 _5398_ (.A1(_3022_),
    .A2(net981),
    .Y(_1892_),
    .B1(_1890_));
 sg13g2_nand2_1 _5399_ (.Y(_1893_),
    .A(net1011),
    .B(_1892_));
 sg13g2_nor2_2 _5400_ (.A(net937),
    .B(_1893_),
    .Y(_1894_));
 sg13g2_nand3_1 _5401_ (.B(_1679_),
    .C(_1892_),
    .A(net1011),
    .Y(_1895_));
 sg13g2_o21ai_1 _5402_ (.B1(_1894_),
    .Y(_1896_),
    .A1(_2856_),
    .A2(net980));
 sg13g2_a21o_1 _5403_ (.A2(_1889_),
    .A1(_1887_),
    .B1(_1896_),
    .X(_1897_));
 sg13g2_inv_1 _5404_ (.Y(_1898_),
    .A(_1897_));
 sg13g2_nand2_1 _5405_ (.Y(_1899_),
    .A(_0114_),
    .B(_1883_));
 sg13g2_xor2_1 _5406_ (.B(_1899_),
    .A(_0112_),
    .X(_1900_));
 sg13g2_or3_1 _5407_ (.A(_1885_),
    .B(_1888_),
    .C(_1900_),
    .X(_1901_));
 sg13g2_o21ai_1 _5408_ (.B1(_1900_),
    .Y(_1902_),
    .A1(_1885_),
    .A2(_1888_));
 sg13g2_and3_1 _5409_ (.X(_1903_),
    .A(net980),
    .B(_1901_),
    .C(_1902_));
 sg13g2_nand3_1 _5410_ (.B(_1901_),
    .C(_1902_),
    .A(net980),
    .Y(_1904_));
 sg13g2_nor2_1 _5411_ (.A(_1895_),
    .B(_1903_),
    .Y(_1905_));
 sg13g2_nand2_1 _5412_ (.Y(_1906_),
    .A(_1894_),
    .B(_1904_));
 sg13g2_nor2_1 _5413_ (.A(_1898_),
    .B(_1905_),
    .Y(_1907_));
 sg13g2_a21oi_1 _5414_ (.A1(_0007_),
    .A2(_1869_),
    .Y(_1908_),
    .B1(net981));
 sg13g2_o21ai_1 _5415_ (.B1(_1891_),
    .Y(_1909_),
    .A1(_2839_),
    .A2(net980));
 sg13g2_a21oi_2 _5416_ (.B1(_1909_),
    .Y(_1910_),
    .A2(_1908_),
    .A1(_1870_));
 sg13g2_inv_1 _5417_ (.Y(_1911_),
    .A(_1910_));
 sg13g2_xnor2_1 _5418_ (.Y(_1912_),
    .A(_1870_),
    .B(_1881_));
 sg13g2_nand2_1 _5419_ (.Y(_1913_),
    .A(net1106),
    .B(net981));
 sg13g2_and2_1 _5420_ (.A(_1891_),
    .B(_1913_),
    .X(_1914_));
 sg13g2_o21ai_1 _5421_ (.B1(_1914_),
    .Y(_1915_),
    .A1(net981),
    .A2(_1912_));
 sg13g2_and2_2 _5422_ (.A(_1910_),
    .B(net869),
    .X(_1916_));
 sg13g2_nand2_1 _5423_ (.Y(_1917_),
    .A(_1907_),
    .B(_1916_));
 sg13g2_and2_2 _5424_ (.A(_1911_),
    .B(net869),
    .X(_1918_));
 sg13g2_nand2_1 _5425_ (.Y(_1919_),
    .A(net1078),
    .B(_1910_));
 sg13g2_o21ai_1 _5426_ (.B1(_1919_),
    .Y(_1920_),
    .A1(_2852_),
    .A2(_1910_));
 sg13g2_o21ai_1 _5427_ (.B1(_1898_),
    .Y(_1921_),
    .A1(net869),
    .A2(_1920_));
 sg13g2_a221oi_1 _5428_ (.B2(_2854_),
    .C1(_1921_),
    .B1(_1918_),
    .A1(_2853_),
    .Y(_1922_),
    .A2(_1916_));
 sg13g2_o21ai_1 _5429_ (.B1(_1902_),
    .Y(_1923_),
    .A1(net1098),
    .A2(_1899_));
 sg13g2_o21ai_1 _5430_ (.B1(net980),
    .Y(_1924_),
    .A1(net1098),
    .A2(_1902_));
 sg13g2_nand2b_1 _5431_ (.Y(_1925_),
    .B(_1923_),
    .A_N(_1924_));
 sg13g2_nand2_1 _5432_ (.Y(_1926_),
    .A(\dtop.field_top.player.controller.pattern0[1] ),
    .B(_1911_));
 sg13g2_a21oi_1 _5433_ (.A1(\dtop.field_top.player.controller.pattern0[0] ),
    .A2(_1910_),
    .Y(_1927_),
    .B1(net869));
 sg13g2_a221oi_1 _5434_ (.B2(_1927_),
    .C1(_1898_),
    .B1(_1926_),
    .A1(_2851_),
    .Y(_1928_),
    .A2(_1916_));
 sg13g2_or4_1 _5435_ (.A(net988),
    .B(_1906_),
    .C(_1925_),
    .D(_1928_),
    .X(_1929_));
 sg13g2_mux4_1 _5436_ (.S0(_1911_),
    .A0(\dtop.field_top.player.osc0[12] ),
    .A1(net1094),
    .A2(net1092),
    .A3(\dtop.field_top.player.osc0[15] ),
    .S1(net869),
    .X(_1930_));
 sg13g2_a21oi_1 _5437_ (.A1(_1894_),
    .A2(_1904_),
    .Y(_1931_),
    .B1(net988));
 sg13g2_mux2_1 _5438_ (.A0(_0015_),
    .A1(_0088_),
    .S(net985),
    .X(_1932_));
 sg13g2_and2_1 _5439_ (.A(_0085_),
    .B(net985),
    .X(_1933_));
 sg13g2_a21oi_1 _5440_ (.A1(_0012_),
    .A2(net987),
    .Y(_1934_),
    .B1(_1933_));
 sg13g2_and2_1 _5441_ (.A(_0086_),
    .B(net985),
    .X(_1935_));
 sg13g2_a21oi_1 _5442_ (.A1(_0069_),
    .A2(net987),
    .Y(_1936_),
    .B1(_1935_));
 sg13g2_mux2_1 _5443_ (.A0(_1936_),
    .A1(_1934_),
    .S(_1910_),
    .X(_1937_));
 sg13g2_nor2_1 _5444_ (.A(_1915_),
    .B(_1937_),
    .Y(_1938_));
 sg13g2_mux2_1 _5445_ (.A0(_0014_),
    .A1(_0087_),
    .S(net985),
    .X(_1939_));
 sg13g2_a221oi_1 _5446_ (.B2(_1916_),
    .C1(_1938_),
    .B1(_1939_),
    .A1(_1918_),
    .Y(_1940_),
    .A2(_1932_));
 sg13g2_a221oi_1 _5447_ (.B2(_1905_),
    .C1(_1898_),
    .B1(_1940_),
    .A1(_1930_),
    .Y(_1941_),
    .A2(_1931_));
 sg13g2_nand2_1 _5448_ (.Y(_1942_),
    .A(_1894_),
    .B(_1925_));
 sg13g2_nor2_1 _5449_ (.A(_2823_),
    .B(_1484_),
    .Y(_1943_));
 sg13g2_nand2_1 _5450_ (.Y(_1944_),
    .A(\dtop.field_top.player.osc0[10] ),
    .B(net985));
 sg13g2_nand2_1 _5451_ (.Y(_1945_),
    .A(\dtop.field_top.player.osc0[11] ),
    .B(net986));
 sg13g2_nor2_1 _5452_ (.A(_2824_),
    .B(net987),
    .Y(_1946_));
 sg13g2_and2_1 _5453_ (.A(_0089_),
    .B(net985),
    .X(_1947_));
 sg13g2_a21oi_1 _5454_ (.A1(_0016_),
    .A2(net987),
    .Y(_1948_),
    .B1(_1947_));
 sg13g2_mux2_1 _5455_ (.A0(_1946_),
    .A1(_1948_),
    .S(_1910_),
    .X(_1949_));
 sg13g2_nor2_1 _5456_ (.A(net869),
    .B(_1949_),
    .Y(_1950_));
 sg13g2_a221oi_1 _5457_ (.B2(_1918_),
    .C1(_1950_),
    .B1(_1945_),
    .A1(_1916_),
    .Y(_1951_),
    .A2(_1944_));
 sg13g2_mux2_1 _5458_ (.A0(_0013_),
    .A1(_0084_),
    .S(net985),
    .X(_1952_));
 sg13g2_nor2_1 _5459_ (.A(_2826_),
    .B(net989),
    .Y(_1953_));
 sg13g2_a21oi_2 _5460_ (.B1(_1953_),
    .Y(_1954_),
    .A2(net989),
    .A1(\dtop.field_top.alt_osc[2] ));
 sg13g2_and2_1 _5461_ (.A(\dtop.field_top.player.osc0[0] ),
    .B(net986),
    .X(_1955_));
 sg13g2_mux2_1 _5462_ (.A0(\dtop.field_top.player.osc0[1] ),
    .A1(\dtop.field_top.alt_osc[1] ),
    .S(net987),
    .X(_1956_));
 sg13g2_mux2_1 _5463_ (.A0(_1956_),
    .A1(_1955_),
    .S(_1910_),
    .X(_1957_));
 sg13g2_nor2_1 _5464_ (.A(net869),
    .B(_1957_),
    .Y(_1958_));
 sg13g2_a22oi_1 _5465_ (.Y(_1959_),
    .B1(_1954_),
    .B2(_1916_),
    .A2(_1952_),
    .A1(_1918_));
 sg13g2_nor3_1 _5466_ (.A(_1895_),
    .B(_1903_),
    .C(_1958_),
    .Y(_1960_));
 sg13g2_a221oi_1 _5467_ (.B2(_1960_),
    .C1(_1897_),
    .B1(_1959_),
    .A1(_1906_),
    .Y(_1961_),
    .A2(_1951_));
 sg13g2_or3_1 _5468_ (.A(_1941_),
    .B(_1942_),
    .C(_1961_),
    .X(_1962_));
 sg13g2_o21ai_1 _5469_ (.B1(_1962_),
    .Y(_1963_),
    .A1(_1922_),
    .A2(_1929_));
 sg13g2_or2_1 _5470_ (.X(_1964_),
    .B(_1918_),
    .A(_1897_));
 sg13g2_inv_1 _5471_ (.Y(_1965_),
    .A(_1964_));
 sg13g2_and3_1 _5472_ (.X(_1966_),
    .A(_1906_),
    .B(_1962_),
    .C(_1964_));
 sg13g2_nand2_1 _5473_ (.Y(_1967_),
    .A(_1907_),
    .B(_1918_));
 sg13g2_o21ai_1 _5474_ (.B1(_0113_),
    .Y(_1968_),
    .A1(_1905_),
    .A2(_1965_));
 sg13g2_nand2_1 _5475_ (.Y(_1969_),
    .A(_1967_),
    .B(_1968_));
 sg13g2_o21ai_1 _5476_ (.B1(_1917_),
    .Y(_1970_),
    .A1(_1966_),
    .A2(_1969_));
 sg13g2_nor4_1 _5477_ (.A(_1897_),
    .B(_1906_),
    .C(_1911_),
    .D(net869),
    .Y(_1971_));
 sg13g2_nor3_1 _5478_ (.A(_1729_),
    .B(_1942_),
    .C(_1971_),
    .Y(_1972_));
 sg13g2_nor2b_1 _5479_ (.A(_1967_),
    .B_N(_1942_),
    .Y(_1973_));
 sg13g2_a21o_1 _5480_ (.A2(_1963_),
    .A1(_1729_),
    .B1(_1973_),
    .X(_1974_));
 sg13g2_a221oi_1 _5481_ (.B2(_1972_),
    .C1(_1973_),
    .B1(_1970_),
    .A1(_1729_),
    .Y(_1975_),
    .A2(_1963_));
 sg13g2_a21o_2 _5482_ (.A2(_1972_),
    .A1(_1970_),
    .B1(_1974_),
    .X(_1976_));
 sg13g2_a21oi_1 _5483_ (.A1(_2928_),
    .A2(_1976_),
    .Y(_1977_),
    .B1(_1729_));
 sg13g2_nor3_1 _5484_ (.A(_1490_),
    .B(_1664_),
    .C(_1895_),
    .Y(_1978_));
 sg13g2_nor2_1 _5485_ (.A(_1690_),
    .B(_1695_),
    .Y(_1979_));
 sg13g2_o21ai_1 _5486_ (.B1(net1095),
    .Y(_1980_),
    .A1(_1690_),
    .A2(_1695_));
 sg13g2_nor2_1 _5487_ (.A(_1699_),
    .B(_1980_),
    .Y(_1981_));
 sg13g2_nor2_1 _5488_ (.A(net1097),
    .B(_1683_),
    .Y(_1982_));
 sg13g2_nand2_1 _5489_ (.Y(_1983_),
    .A(_2856_),
    .B(_1722_));
 sg13g2_a21oi_2 _5490_ (.B1(net1097),
    .Y(_1984_),
    .A2(_1683_),
    .A1(_2860_));
 sg13g2_inv_1 _5491_ (.Y(_1985_),
    .A(_1984_));
 sg13g2_a22oi_1 _5492_ (.Y(_1986_),
    .B1(_1984_),
    .B2(_1685_),
    .A2(_1981_),
    .A1(_1688_));
 sg13g2_nand2_1 _5493_ (.Y(_1987_),
    .A(net1025),
    .B(_1986_));
 sg13g2_nand2_1 _5494_ (.Y(_1988_),
    .A(net1095),
    .B(_1687_));
 sg13g2_a21o_1 _5495_ (.A2(_1987_),
    .A1(_1712_),
    .B1(_1680_),
    .X(_1989_));
 sg13g2_nor2_2 _5496_ (.A(_0111_),
    .B(net937),
    .Y(_1990_));
 sg13g2_nand4_1 _5497_ (.B(_1985_),
    .C(_1988_),
    .A(net1028),
    .Y(_1991_),
    .D(_1990_));
 sg13g2_xnor2_1 _5498_ (.Y(_1992_),
    .A(_1989_),
    .B(_1991_));
 sg13g2_o21ai_1 _5499_ (.B1(_1729_),
    .Y(_1993_),
    .A1(_1894_),
    .A2(_1992_));
 sg13g2_a21oi_1 _5500_ (.A1(_1976_),
    .A2(_1978_),
    .Y(_1994_),
    .B1(_1993_));
 sg13g2_o21ai_1 _5501_ (.B1(_1720_),
    .Y(_1995_),
    .A1(_1977_),
    .A2(_1994_));
 sg13g2_a21oi_1 _5502_ (.A1(_0113_),
    .A2(_1719_),
    .Y(_1996_),
    .B1(net1));
 sg13g2_and2_1 _5503_ (.A(_1995_),
    .B(_1996_),
    .X(_1997_));
 sg13g2_nor2_2 _5504_ (.A(net1096),
    .B(net1026),
    .Y(_1998_));
 sg13g2_nor2b_1 _5505_ (.A(net1097),
    .B_N(net1099),
    .Y(_1999_));
 sg13g2_nand4_1 _5506_ (.B(_0117_),
    .C(net952),
    .A(net1099),
    .Y(_2000_),
    .D(_1998_));
 sg13g2_nand2_1 _5507_ (.Y(_2001_),
    .A(_3009_),
    .B(_2000_));
 sg13g2_nor2_2 _5508_ (.A(net942),
    .B(_1678_),
    .Y(_2002_));
 sg13g2_nand3_1 _5509_ (.B(_3000_),
    .C(_1689_),
    .A(_2995_),
    .Y(_2003_));
 sg13g2_nand3b_1 _5510_ (.B(_3019_),
    .C(_1998_),
    .Y(_2004_),
    .A_N(net1100));
 sg13g2_nand2_1 _5511_ (.Y(_2005_),
    .A(_2003_),
    .B(_2004_));
 sg13g2_a22oi_1 _5512_ (.Y(_2006_),
    .B1(_2002_),
    .B2(_2005_),
    .A2(_2001_),
    .A1(_1679_));
 sg13g2_nand4_1 _5513_ (.B(net1099),
    .C(_1694_),
    .A(_2856_),
    .Y(_2007_),
    .D(_1998_));
 sg13g2_nand2_1 _5514_ (.Y(_2008_),
    .A(_2004_),
    .B(_2007_));
 sg13g2_nor2_1 _5515_ (.A(net1026),
    .B(_1708_),
    .Y(_2009_));
 sg13g2_o21ai_1 _5516_ (.B1(_2003_),
    .Y(_2010_),
    .A1(net1025),
    .A2(_1708_));
 sg13g2_nor2_1 _5517_ (.A(_2008_),
    .B(_2009_),
    .Y(_2011_));
 sg13g2_nor2_1 _5518_ (.A(_2008_),
    .B(_2010_),
    .Y(_2012_));
 sg13g2_o21ai_1 _5519_ (.B1(_2002_),
    .Y(_2013_),
    .A1(_1722_),
    .A2(_2012_));
 sg13g2_nand3_1 _5520_ (.B(_2995_),
    .C(net965),
    .A(net1120),
    .Y(_2014_));
 sg13g2_nand4_1 _5521_ (.B(_2860_),
    .C(net944),
    .A(net1010),
    .Y(_2015_),
    .D(_1724_));
 sg13g2_nand3_1 _5522_ (.B(net1095),
    .C(_3020_),
    .A(net1099),
    .Y(_2016_));
 sg13g2_or2_1 _5523_ (.X(_2017_),
    .B(_2016_),
    .A(net1010));
 sg13g2_nand3_1 _5524_ (.B(_2015_),
    .C(_2017_),
    .A(_1679_),
    .Y(_2018_));
 sg13g2_nand3_1 _5525_ (.B(_2014_),
    .C(_2018_),
    .A(_2013_),
    .Y(_2019_));
 sg13g2_and2_1 _5526_ (.A(_2002_),
    .B(_2010_),
    .X(_2020_));
 sg13g2_nor2_1 _5527_ (.A(net945),
    .B(_1999_),
    .Y(_2021_));
 sg13g2_a21oi_1 _5528_ (.A1(net1107),
    .A2(_1999_),
    .Y(_2022_),
    .B1(net944));
 sg13g2_a21oi_1 _5529_ (.A1(_0115_),
    .A2(_1694_),
    .Y(_2023_),
    .B1(_1724_));
 sg13g2_o21ai_1 _5530_ (.B1(net1010),
    .Y(_2024_),
    .A1(net952),
    .A2(_2023_));
 sg13g2_o21ai_1 _5531_ (.B1(_2017_),
    .Y(_2025_),
    .A1(_2022_),
    .A2(_2024_));
 sg13g2_a21o_1 _5532_ (.A2(_2025_),
    .A1(_1679_),
    .B1(_2020_),
    .X(_2026_));
 sg13g2_nand2b_1 _5533_ (.Y(_2027_),
    .B(_2019_),
    .A_N(_2026_));
 sg13g2_nor2_1 _5534_ (.A(_2006_),
    .B(_2027_),
    .Y(_2028_));
 sg13g2_a21oi_1 _5535_ (.A1(_2860_),
    .A2(_1725_),
    .Y(_2029_),
    .B1(net981));
 sg13g2_nor3_1 _5536_ (.A(net952),
    .B(_2023_),
    .C(_2029_),
    .Y(_2030_));
 sg13g2_or3_1 _5537_ (.A(net1025),
    .B(_2021_),
    .C(_2030_),
    .X(_2031_));
 sg13g2_nor2_1 _5538_ (.A(_3015_),
    .B(_1690_),
    .Y(_2032_));
 sg13g2_nand2_1 _5539_ (.Y(_2033_),
    .A(net1107),
    .B(_1691_));
 sg13g2_nand4_1 _5540_ (.B(_1688_),
    .C(_1706_),
    .A(net1025),
    .Y(_2034_),
    .D(_2033_));
 sg13g2_nand3_1 _5541_ (.B(_2031_),
    .C(_2034_),
    .A(net941),
    .Y(_2035_));
 sg13g2_nand3_1 _5542_ (.B(_1694_),
    .C(_1998_),
    .A(_1682_),
    .Y(_2036_));
 sg13g2_nand3_1 _5543_ (.B(_1689_),
    .C(_1998_),
    .A(_2995_),
    .Y(_2037_));
 sg13g2_nand2_1 _5544_ (.Y(_2038_),
    .A(_1998_),
    .B(_2032_));
 sg13g2_nand2_1 _5545_ (.Y(_2039_),
    .A(_2037_),
    .B(_2038_));
 sg13g2_nor2b_1 _5546_ (.A(_2039_),
    .B_N(_2036_),
    .Y(_2040_));
 sg13g2_o21ai_1 _5547_ (.B1(_2035_),
    .Y(_2041_),
    .A1(net941),
    .A2(_2040_));
 sg13g2_nor2_1 _5548_ (.A(net965),
    .B(_2041_),
    .Y(_2042_));
 sg13g2_nor2_1 _5549_ (.A(_2019_),
    .B(_2026_),
    .Y(_2043_));
 sg13g2_nand2b_1 _5550_ (.Y(_2044_),
    .B(_2043_),
    .A_N(_2042_));
 sg13g2_and2_1 _5551_ (.A(_2006_),
    .B(_2042_),
    .X(_2045_));
 sg13g2_nor2b_1 _5552_ (.A(_2027_),
    .B_N(_2045_),
    .Y(_2046_));
 sg13g2_and2_1 _5553_ (.A(_2027_),
    .B(_2045_),
    .X(_2047_));
 sg13g2_nand2b_1 _5554_ (.Y(_2048_),
    .B(_2026_),
    .A_N(_2019_));
 sg13g2_nor2_1 _5555_ (.A(_2006_),
    .B(_2048_),
    .Y(_2049_));
 sg13g2_a22oi_1 _5556_ (.Y(_2050_),
    .B1(net873),
    .B2(\dtop.field_top.channel_output[1] ),
    .A2(net881),
    .A1(\dtop.field_top.channel_output[10] ));
 sg13g2_a22oi_1 _5557_ (.Y(_2051_),
    .B1(_2049_),
    .B2(\dtop.field_top.player.out_acc[0] ),
    .A2(net874),
    .A1(\dtop.field_top.channel_output[0] ));
 sg13g2_and3_1 _5558_ (.X(_2052_),
    .A(net876),
    .B(_2050_),
    .C(_2051_));
 sg13g2_o21ai_1 _5559_ (.B1(_1728_),
    .Y(_2053_),
    .A1(net1107),
    .A2(net944));
 sg13g2_nand2_1 _5560_ (.Y(_2054_),
    .A(net1010),
    .B(_2053_));
 sg13g2_a21oi_1 _5561_ (.A1(_1684_),
    .A2(_1686_),
    .Y(_2055_),
    .B1(_1691_));
 sg13g2_nor3_1 _5562_ (.A(net1010),
    .B(_0112_),
    .C(_2055_),
    .Y(_2056_));
 sg13g2_nor2_1 _5563_ (.A(net937),
    .B(_2056_),
    .Y(_2057_));
 sg13g2_o21ai_1 _5564_ (.B1(_1998_),
    .Y(_2058_),
    .A1(_1696_),
    .A2(_1979_));
 sg13g2_nand3_1 _5565_ (.B(_2007_),
    .C(_2058_),
    .A(_2003_),
    .Y(_2059_));
 sg13g2_nand3_1 _5566_ (.B(_2038_),
    .C(_2058_),
    .A(_2012_),
    .Y(_2060_));
 sg13g2_a22oi_1 _5567_ (.Y(_2061_),
    .B1(_2060_),
    .B2(_2002_),
    .A2(_2057_),
    .A1(_2054_));
 sg13g2_and2_2 _5568_ (.A(_2014_),
    .B(_2061_),
    .X(_2062_));
 sg13g2_inv_1 _5569_ (.Y(_2063_),
    .A(_2062_));
 sg13g2_nor2_2 _5570_ (.A(_1975_),
    .B(_2063_),
    .Y(_2064_));
 sg13g2_nand2_2 _5571_ (.Y(_2065_),
    .A(_1976_),
    .B(_2062_));
 sg13g2_nand3_1 _5572_ (.B(_1688_),
    .C(_1692_),
    .A(net1095),
    .Y(_2066_));
 sg13g2_a21oi_1 _5573_ (.A1(_1684_),
    .A2(_1984_),
    .Y(_2067_),
    .B1(net1010));
 sg13g2_nand2_1 _5574_ (.Y(_2068_),
    .A(_2066_),
    .B(_2067_));
 sg13g2_nand4_1 _5575_ (.B(_1893_),
    .C(_2000_),
    .A(net941),
    .Y(_2069_),
    .D(_2068_));
 sg13g2_nor2_1 _5576_ (.A(net941),
    .B(_2039_),
    .Y(_2070_));
 sg13g2_nor2_1 _5577_ (.A(net965),
    .B(_2070_),
    .Y(_2071_));
 sg13g2_a21oi_2 _5578_ (.B1(_1719_),
    .Y(_2072_),
    .A2(_2071_),
    .A1(_2069_));
 sg13g2_nor2_2 _5579_ (.A(_1975_),
    .B(_2072_),
    .Y(_2073_));
 sg13g2_or2_2 _5580_ (.X(_2074_),
    .B(_2072_),
    .A(_1975_));
 sg13g2_a21oi_2 _5581_ (.B1(_1975_),
    .Y(_2075_),
    .A2(_2072_),
    .A1(_2063_));
 sg13g2_nand2_1 _5582_ (.Y(_2076_),
    .A(_0117_),
    .B(_1669_));
 sg13g2_o21ai_1 _5583_ (.B1(_2029_),
    .Y(_2077_),
    .A1(_1725_),
    .A2(_2076_));
 sg13g2_o21ai_1 _5584_ (.B1(net981),
    .Y(_2078_),
    .A1(_3022_),
    .A2(_1668_));
 sg13g2_a21oi_1 _5585_ (.A1(_2077_),
    .A2(_2078_),
    .Y(_2079_),
    .B1(net952));
 sg13g2_nor3_1 _5586_ (.A(net1027),
    .B(_2022_),
    .C(_2079_),
    .Y(_2080_));
 sg13g2_nand4_1 _5587_ (.B(_3008_),
    .C(_1685_),
    .A(net1095),
    .Y(_2081_),
    .D(_2055_));
 sg13g2_nand2_1 _5588_ (.Y(_2082_),
    .A(net1025),
    .B(_1705_));
 sg13g2_a21oi_1 _5589_ (.A1(net1105),
    .A2(_1982_),
    .Y(_2083_),
    .B1(_2082_));
 sg13g2_a21oi_1 _5590_ (.A1(_2081_),
    .A2(_2083_),
    .Y(_2084_),
    .B1(_2080_));
 sg13g2_nand2_1 _5591_ (.Y(_2085_),
    .A(_2002_),
    .B(_2059_));
 sg13g2_o21ai_1 _5592_ (.B1(_2085_),
    .Y(_2086_),
    .A1(net937),
    .A2(_2084_));
 sg13g2_or2_1 _5593_ (.X(_2087_),
    .B(_1681_),
    .A(_1490_));
 sg13g2_or2_1 _5594_ (.X(_2088_),
    .B(_2087_),
    .A(_2086_));
 sg13g2_nor4_2 _5595_ (.A(_0111_),
    .B(_2996_),
    .C(net937),
    .Y(_2089_),
    .D(_1983_));
 sg13g2_nand3_1 _5596_ (.B(_1982_),
    .C(_1990_),
    .A(_2995_),
    .Y(_2090_));
 sg13g2_or4_2 _5597_ (.A(_1975_),
    .B(_2075_),
    .C(_2088_),
    .D(_2090_),
    .X(_2091_));
 sg13g2_nand2b_2 _5598_ (.Y(_2092_),
    .B(_2836_),
    .A_N(_2091_));
 sg13g2_o21ai_1 _5599_ (.B1(_1976_),
    .Y(_2093_),
    .A1(_2086_),
    .A2(_2089_));
 sg13g2_and3_1 _5600_ (.X(_2094_),
    .A(_2064_),
    .B(_2073_),
    .C(_2093_));
 sg13g2_nand3_1 _5601_ (.B(_2073_),
    .C(_2093_),
    .A(_2064_),
    .Y(_2095_));
 sg13g2_and2_2 _5602_ (.A(_1729_),
    .B(_2094_),
    .X(_2096_));
 sg13g2_nand3_1 _5603_ (.B(_2062_),
    .C(_2072_),
    .A(_1976_),
    .Y(_2097_));
 sg13g2_and3_1 _5604_ (.X(_2098_),
    .A(_2064_),
    .B(_2074_),
    .C(_2093_));
 sg13g2_nand3_1 _5605_ (.B(_2086_),
    .C(_2090_),
    .A(_1976_),
    .Y(_2099_));
 sg13g2_nor2_1 _5606_ (.A(_2075_),
    .B(net850),
    .Y(_2100_));
 sg13g2_a22oi_1 _5607_ (.Y(_2101_),
    .B1(_2100_),
    .B2(net1028),
    .A2(_2098_),
    .A1(_1943_));
 sg13g2_nand3b_1 _5608_ (.B(_2089_),
    .C(_1976_),
    .Y(_2102_),
    .A_N(_2086_));
 sg13g2_nand2_1 _5609_ (.Y(_2103_),
    .A(_2092_),
    .B(_2101_));
 sg13g2_nand4_1 _5610_ (.B(_2063_),
    .C(_2072_),
    .A(_1976_),
    .Y(_2104_),
    .D(_2089_));
 sg13g2_nor2_2 _5611_ (.A(_2088_),
    .B(_2104_),
    .Y(_2105_));
 sg13g2_a21oi_1 _5612_ (.A1(\dtop.field_top.player.osc0[21] ),
    .A2(_2096_),
    .Y(_2106_),
    .B1(_2103_));
 sg13g2_nand2_2 _5613_ (.Y(_2107_),
    .A(_1992_),
    .B(_2092_));
 sg13g2_and4_1 _5614_ (.A(_1955_),
    .B(_2064_),
    .C(_2074_),
    .D(_2093_),
    .X(_2108_));
 sg13g2_nor3_1 _5615_ (.A(_2822_),
    .B(_2075_),
    .C(_2099_),
    .Y(_2109_));
 sg13g2_nor2_2 _5616_ (.A(_2097_),
    .B(net850),
    .Y(_2110_));
 sg13g2_nand2_1 _5617_ (.Y(_2111_),
    .A(net938),
    .B(_2110_));
 sg13g2_nor4_1 _5618_ (.A(_0087_),
    .B(net949),
    .C(_2097_),
    .D(_2099_),
    .Y(_2112_));
 sg13g2_and4_1 _5619_ (.A(_2927_),
    .B(_2064_),
    .C(_2073_),
    .D(_2093_),
    .X(_2113_));
 sg13g2_and3_2 _5620_ (.X(_2114_),
    .A(_2065_),
    .B(_2073_),
    .C(_2093_));
 sg13g2_inv_1 _5621_ (.Y(_2115_),
    .A(_2114_));
 sg13g2_nor3_2 _5622_ (.A(_2065_),
    .B(_2074_),
    .C(net850),
    .Y(_2116_));
 sg13g2_or3_1 _5623_ (.A(_2065_),
    .B(_2074_),
    .C(net850),
    .X(_2117_));
 sg13g2_nand2_1 _5624_ (.Y(_2118_),
    .A(_0084_),
    .B(net940));
 sg13g2_nor2_1 _5625_ (.A(_0086_),
    .B(net938),
    .Y(_2119_));
 sg13g2_o21ai_1 _5626_ (.B1(net946),
    .Y(_2120_),
    .A1(_0088_),
    .A2(net949));
 sg13g2_o21ai_1 _5627_ (.B1(_2118_),
    .Y(_2121_),
    .A1(_2119_),
    .A2(_2120_));
 sg13g2_nor4_1 _5628_ (.A(_2065_),
    .B(_2074_),
    .C(net850),
    .D(_2121_),
    .Y(_2122_));
 sg13g2_nor3_2 _5629_ (.A(_2064_),
    .B(_2074_),
    .C(net850),
    .Y(_2123_));
 sg13g2_nand3b_1 _5630_ (.B(_2065_),
    .C(_2073_),
    .Y(_2124_),
    .A_N(net850));
 sg13g2_or2_1 _5631_ (.X(_2125_),
    .B(_1860_),
    .A(_1805_));
 sg13g2_or2_1 _5632_ (.X(_2126_),
    .B(_2125_),
    .A(_1768_));
 sg13g2_nand3_1 _5633_ (.B(_1861_),
    .C(_2125_),
    .A(_1768_),
    .Y(_2127_));
 sg13g2_a21oi_1 _5634_ (.A1(_2126_),
    .A2(_2127_),
    .Y(_2128_),
    .B1(_1770_));
 sg13g2_a21o_1 _5635_ (.A2(_1805_),
    .A1(_1770_),
    .B1(_1653_),
    .X(_2129_));
 sg13g2_nor2_2 _5636_ (.A(_2835_),
    .B(net943),
    .Y(_2130_));
 sg13g2_nor2_1 _5637_ (.A(_1867_),
    .B(_2130_),
    .Y(_2131_));
 sg13g2_o21ai_1 _5638_ (.B1(_2131_),
    .Y(_2132_),
    .A1(_2128_),
    .A2(_2129_));
 sg13g2_nand2_1 _5639_ (.Y(_2133_),
    .A(_1769_),
    .B(_1825_));
 sg13g2_or2_1 _5640_ (.X(_2134_),
    .B(_2133_),
    .A(_1859_));
 sg13g2_a21oi_1 _5641_ (.A1(_1859_),
    .A2(_2133_),
    .Y(_2135_),
    .B1(_1653_));
 sg13g2_a221oi_1 _5642_ (.B2(_2135_),
    .C1(_1867_),
    .B1(_2134_),
    .A1(_1660_),
    .Y(_2136_),
    .A2(_2130_));
 sg13g2_xor2_1 _5643_ (.B(_2136_),
    .A(_2132_),
    .X(_2137_));
 sg13g2_xnor2_1 _5644_ (.Y(_2138_),
    .A(_1768_),
    .B(_1862_));
 sg13g2_nand4_1 _5645_ (.B(_1866_),
    .C(_2126_),
    .A(net943),
    .Y(_2139_),
    .D(_2138_));
 sg13g2_inv_1 _5646_ (.Y(_2140_),
    .A(_2139_));
 sg13g2_xnor2_1 _5647_ (.Y(_2141_),
    .A(_1770_),
    .B(_1825_));
 sg13g2_nor2_1 _5648_ (.A(_2855_),
    .B(_1654_),
    .Y(_2142_));
 sg13g2_a22oi_1 _5649_ (.Y(_2143_),
    .B1(_2142_),
    .B2(_1660_),
    .A2(_2141_),
    .A1(net943));
 sg13g2_nor2_2 _5650_ (.A(_1867_),
    .B(_2143_),
    .Y(_2144_));
 sg13g2_nand2b_1 _5651_ (.Y(_2145_),
    .B(_1866_),
    .A_N(_2143_));
 sg13g2_nand2_1 _5652_ (.Y(_2146_),
    .A(_2139_),
    .B(_2145_));
 sg13g2_nand2b_1 _5653_ (.Y(_2147_),
    .B(_2145_),
    .A_N(_2136_));
 sg13g2_nand2_2 _5654_ (.Y(_2148_),
    .A(_2140_),
    .B(_2144_));
 sg13g2_o21ai_1 _5655_ (.B1(_2148_),
    .Y(_2149_),
    .A1(_2137_),
    .A2(_2146_));
 sg13g2_nor4_1 _5656_ (.A(_2064_),
    .B(_2074_),
    .C(net850),
    .D(_2149_),
    .Y(_2150_));
 sg13g2_nor4_2 _5657_ (.A(_2108_),
    .B(_2109_),
    .C(_2113_),
    .Y(_2151_),
    .D(_2122_));
 sg13g2_nor4_1 _5658_ (.A(\dtop.field_top.player.osc0[4] ),
    .B(_2075_),
    .C(_2087_),
    .D(_2102_),
    .Y(_2152_));
 sg13g2_nor4_2 _5659_ (.A(_2112_),
    .B(_2114_),
    .C(_2150_),
    .Y(_2153_),
    .D(_2152_));
 sg13g2_and4_1 _5660_ (.A(_1992_),
    .B(_2092_),
    .C(_2151_),
    .D(_2153_),
    .X(_2154_));
 sg13g2_a22oi_1 _5661_ (.Y(_2155_),
    .B1(_2151_),
    .B2(_2153_),
    .A2(_2092_),
    .A1(_1992_));
 sg13g2_nor3_1 _5662_ (.A(_2052_),
    .B(_2154_),
    .C(_2155_),
    .Y(_2156_));
 sg13g2_o21ai_1 _5663_ (.B1(_2052_),
    .Y(_2157_),
    .A1(_2154_),
    .A2(_2155_));
 sg13g2_nand2b_1 _5664_ (.Y(_2158_),
    .B(_2157_),
    .A_N(_2156_));
 sg13g2_xor2_1 _5665_ (.B(_2158_),
    .A(_1997_),
    .X(_2159_));
 sg13g2_nor3_1 _5666_ (.A(net1120),
    .B(net2),
    .C(net1),
    .Y(_2160_));
 sg13g2_a21oi_1 _5667_ (.A1(net612),
    .A2(net868),
    .Y(_2161_),
    .B1(net1113));
 sg13g2_o21ai_1 _5668_ (.B1(_2161_),
    .Y(_0164_),
    .A1(net868),
    .A2(_2159_));
 sg13g2_a21oi_1 _5669_ (.A1(_1997_),
    .A2(_2157_),
    .Y(_2162_),
    .B1(_2156_));
 sg13g2_a22oi_1 _5670_ (.Y(_2163_),
    .B1(net880),
    .B2(\dtop.field_top.player.out_acc[1] ),
    .A2(net874),
    .A1(\dtop.field_top.channel_output[1] ));
 sg13g2_nand2_1 _5671_ (.Y(_2164_),
    .A(net876),
    .B(_2163_));
 sg13g2_a221oi_1 _5672_ (.B2(\dtop.field_top.channel_output[2] ),
    .C1(_2164_),
    .B1(net873),
    .A1(\dtop.field_top.channel_output[0] ),
    .Y(_2165_),
    .A2(net881));
 sg13g2_nor3_1 _5673_ (.A(\dtop.field_top.player.osc0[5] ),
    .B(_2088_),
    .C(_2104_),
    .Y(_2166_));
 sg13g2_a221oi_1 _5674_ (.B2(\dtop.field_top.channel_output[1] ),
    .C1(_2166_),
    .B1(_2100_),
    .A1(_1956_),
    .Y(_2167_),
    .A2(net849));
 sg13g2_mux2_1 _5675_ (.A0(_2144_),
    .A1(_2143_),
    .S(_2136_),
    .X(_2168_));
 sg13g2_nand2b_1 _5676_ (.Y(_2169_),
    .B(_2168_),
    .A_N(_2132_));
 sg13g2_nand2_1 _5677_ (.Y(_2170_),
    .A(_2139_),
    .B(_2169_));
 sg13g2_nand2_1 _5678_ (.Y(_2171_),
    .A(_2136_),
    .B(_2140_));
 sg13g2_nand3_1 _5679_ (.B(_2170_),
    .C(_2171_),
    .A(_2148_),
    .Y(_2172_));
 sg13g2_mux2_1 _5680_ (.A0(_0089_),
    .A1(_0087_),
    .S(net949),
    .X(_2173_));
 sg13g2_a22oi_1 _5681_ (.Y(_2174_),
    .B1(_2173_),
    .B2(net946),
    .A2(net939),
    .A1(_0085_));
 sg13g2_a22oi_1 _5682_ (.Y(_2175_),
    .B1(_2123_),
    .B2(_2172_),
    .A2(_2094_),
    .A1(_2926_));
 sg13g2_a21oi_1 _5683_ (.A1(_2116_),
    .A2(_2174_),
    .Y(_2176_),
    .B1(_2114_));
 sg13g2_nand3b_1 _5684_ (.B(net938),
    .C(_2110_),
    .Y(_2177_),
    .A_N(_0088_));
 sg13g2_nand4_1 _5685_ (.B(_2175_),
    .C(_2176_),
    .A(_2167_),
    .Y(_2178_),
    .D(_2177_));
 sg13g2_xor2_1 _5686_ (.B(_2178_),
    .A(_2107_),
    .X(_2179_));
 sg13g2_nand2b_1 _5687_ (.Y(_2180_),
    .B(_2179_),
    .A_N(_2165_));
 sg13g2_xnor2_1 _5688_ (.Y(_2181_),
    .A(_2165_),
    .B(_2179_));
 sg13g2_nand2b_1 _5689_ (.Y(_2182_),
    .B(_2181_),
    .A_N(_2162_));
 sg13g2_xor2_1 _5690_ (.B(_2181_),
    .A(_2162_),
    .X(_2183_));
 sg13g2_a21oi_1 _5691_ (.A1(net654),
    .A2(_1721_),
    .Y(_2184_),
    .B1(net1112));
 sg13g2_o21ai_1 _5692_ (.B1(_2184_),
    .Y(_0165_),
    .A1(net868),
    .A2(_2183_));
 sg13g2_a22oi_1 _5693_ (.Y(_2185_),
    .B1(net873),
    .B2(\dtop.field_top.channel_output[3] ),
    .A2(net881),
    .A1(\dtop.field_top.channel_output[5] ));
 sg13g2_a22oi_1 _5694_ (.Y(_2186_),
    .B1(net880),
    .B2(\dtop.field_top.player.out_acc[2] ),
    .A2(net874),
    .A1(\dtop.field_top.channel_output[2] ));
 sg13g2_and3_1 _5695_ (.X(_2187_),
    .A(net876),
    .B(_2185_),
    .C(_2186_));
 sg13g2_o21ai_1 _5696_ (.B1(_2171_),
    .Y(_2188_),
    .A1(_2132_),
    .A2(_2144_));
 sg13g2_o21ai_1 _5697_ (.B1(_2188_),
    .Y(_2189_),
    .A1(_2139_),
    .A2(_2144_));
 sg13g2_and2_1 _5698_ (.A(_2123_),
    .B(_2189_),
    .X(_2190_));
 sg13g2_nor2_1 _5699_ (.A(\dtop.field_top.player.controller.ppos[0] ),
    .B(_2095_),
    .Y(_2191_));
 sg13g2_mux2_1 _5700_ (.A0(_0090_),
    .A1(_0088_),
    .S(net949),
    .X(_2192_));
 sg13g2_a221oi_1 _5701_ (.B2(net946),
    .C1(_2117_),
    .B1(_2192_),
    .A1(_0086_),
    .Y(_2193_),
    .A2(net939));
 sg13g2_nor2_1 _5702_ (.A(\dtop.field_top.player.osc0[6] ),
    .B(_2091_),
    .Y(_2194_));
 sg13g2_nor4_1 _5703_ (.A(_2190_),
    .B(_2191_),
    .C(_2193_),
    .D(_2194_),
    .Y(_2195_));
 sg13g2_a21oi_1 _5704_ (.A1(\dtop.field_top.channel_output[2] ),
    .A2(net848),
    .Y(_2196_),
    .B1(_2114_));
 sg13g2_nand2b_1 _5705_ (.Y(_2197_),
    .B(_2098_),
    .A_N(_1954_));
 sg13g2_or2_1 _5706_ (.X(_2198_),
    .B(_2111_),
    .A(_0089_));
 sg13g2_nand4_1 _5707_ (.B(_2196_),
    .C(_2197_),
    .A(_2195_),
    .Y(_2199_),
    .D(_2198_));
 sg13g2_xor2_1 _5708_ (.B(_2199_),
    .A(net847),
    .X(_2200_));
 sg13g2_nor2b_1 _5709_ (.A(_2187_),
    .B_N(_2200_),
    .Y(_2201_));
 sg13g2_xor2_1 _5710_ (.B(_2200_),
    .A(_2187_),
    .X(_2202_));
 sg13g2_a21oi_2 _5711_ (.B1(_2202_),
    .Y(_2203_),
    .A2(_2182_),
    .A1(_2180_));
 sg13g2_nand3_1 _5712_ (.B(_2182_),
    .C(_2202_),
    .A(_2180_),
    .Y(_2204_));
 sg13g2_nor2b_2 _5713_ (.A(_2203_),
    .B_N(_2204_),
    .Y(_2205_));
 sg13g2_nand2b_1 _5714_ (.Y(_2206_),
    .B(_2205_),
    .A_N(net868));
 sg13g2_a21oi_1 _5715_ (.A1(net1094),
    .A2(net868),
    .Y(_2207_),
    .B1(net1111));
 sg13g2_nand2_1 _5716_ (.Y(_0166_),
    .A(_2206_),
    .B(_2207_));
 sg13g2_nor2_1 _5717_ (.A(_2201_),
    .B(_2203_),
    .Y(_2208_));
 sg13g2_a22oi_1 _5718_ (.Y(_2209_),
    .B1(net873),
    .B2(\dtop.field_top.channel_output[4] ),
    .A2(net881),
    .A1(\dtop.field_top.channel_output[1] ));
 sg13g2_a22oi_1 _5719_ (.Y(_2210_),
    .B1(net880),
    .B2(\dtop.field_top.player.out_acc[3] ),
    .A2(net875),
    .A1(\dtop.field_top.channel_output[3] ));
 sg13g2_nand3_1 _5720_ (.B(_2209_),
    .C(_2210_),
    .A(net876),
    .Y(_2211_));
 sg13g2_o21ai_1 _5721_ (.B1(_2139_),
    .Y(_2212_),
    .A1(_2132_),
    .A2(_2136_));
 sg13g2_o21ai_1 _5722_ (.B1(_2212_),
    .Y(_2213_),
    .A1(_2136_),
    .A2(_2148_));
 sg13g2_nor2_1 _5723_ (.A(\dtop.field_top.player.controller.timer[0] ),
    .B(net949),
    .Y(_2214_));
 sg13g2_o21ai_1 _5724_ (.B1(net946),
    .Y(_2215_),
    .A1(_0089_),
    .A2(net938));
 sg13g2_nor2_1 _5725_ (.A(_2214_),
    .B(_2215_),
    .Y(_2216_));
 sg13g2_a21oi_1 _5726_ (.A1(_0087_),
    .A2(net939),
    .Y(_2217_),
    .B1(_2216_));
 sg13g2_a21o_1 _5727_ (.A2(_1729_),
    .A1(\dtop.field_top.player.controller.ppos[1] ),
    .B1(_2095_),
    .X(_2218_));
 sg13g2_nand2_1 _5728_ (.Y(_2219_),
    .A(\dtop.field_top.channel_output[3] ),
    .B(net848));
 sg13g2_nand2b_1 _5729_ (.Y(_2220_),
    .B(net849),
    .A_N(_1952_));
 sg13g2_nor3_1 _5730_ (.A(\dtop.field_top.player.osc0[7] ),
    .B(_2088_),
    .C(_2104_),
    .Y(_2221_));
 sg13g2_o21ai_1 _5731_ (.B1(_2219_),
    .Y(_2222_),
    .A1(_0090_),
    .A2(_2111_));
 sg13g2_a22oi_1 _5732_ (.Y(_2223_),
    .B1(_2217_),
    .B2(_2116_),
    .A2(_2213_),
    .A1(_2123_));
 sg13g2_nand3_1 _5733_ (.B(_2220_),
    .C(_2223_),
    .A(_2218_),
    .Y(_2224_));
 sg13g2_nor4_2 _5734_ (.A(_2114_),
    .B(_2221_),
    .C(_2222_),
    .Y(_2225_),
    .D(_2224_));
 sg13g2_xnor2_1 _5735_ (.Y(_2226_),
    .A(net847),
    .B(_2225_));
 sg13g2_and2_1 _5736_ (.A(_2211_),
    .B(_2226_),
    .X(_2227_));
 sg13g2_xor2_1 _5737_ (.B(_2226_),
    .A(_2211_),
    .X(_2228_));
 sg13g2_o21ai_1 _5738_ (.B1(_2228_),
    .Y(_2229_),
    .A1(_2201_),
    .A2(_2203_));
 sg13g2_xor2_1 _5739_ (.B(_2228_),
    .A(_2208_),
    .X(_2230_));
 sg13g2_inv_1 _5740_ (.Y(_2231_),
    .A(_2230_));
 sg13g2_a21oi_1 _5741_ (.A1(net1092),
    .A2(net868),
    .Y(_2232_),
    .B1(net1111));
 sg13g2_o21ai_1 _5742_ (.B1(_2232_),
    .Y(_0167_),
    .A1(net867),
    .A2(_2230_));
 sg13g2_nand2b_1 _5743_ (.Y(_2233_),
    .B(_2229_),
    .A_N(_2227_));
 sg13g2_a22oi_1 _5744_ (.Y(_2234_),
    .B1(net880),
    .B2(\dtop.field_top.player.out_acc[4] ),
    .A2(net874),
    .A1(\dtop.field_top.channel_output[4] ));
 sg13g2_nand2_1 _5745_ (.Y(_2235_),
    .A(net876),
    .B(_2234_));
 sg13g2_a221oi_1 _5746_ (.B2(\dtop.field_top.channel_output[5] ),
    .C1(_2235_),
    .B1(net873),
    .A1(\dtop.field_top.channel_output[6] ),
    .Y(_2236_),
    .A2(net881));
 sg13g2_nand2_1 _5747_ (.Y(_2237_),
    .A(_2855_),
    .B(_2096_));
 sg13g2_nor2_1 _5748_ (.A(_2927_),
    .B(_1867_),
    .Y(_2238_));
 sg13g2_a221oi_1 _5749_ (.B2(_0090_),
    .C1(_2238_),
    .B1(net949),
    .A1(_0088_),
    .Y(_2239_),
    .A2(net939));
 sg13g2_xnor2_1 _5750_ (.Y(_2240_),
    .A(_2132_),
    .B(_2144_));
 sg13g2_nand2_1 _5751_ (.Y(_2241_),
    .A(_2139_),
    .B(_2240_));
 sg13g2_and4_1 _5752_ (.A(_2123_),
    .B(_2148_),
    .C(_2171_),
    .D(_2241_),
    .X(_2242_));
 sg13g2_nand2b_1 _5753_ (.Y(_2243_),
    .B(_2105_),
    .A_N(\dtop.field_top.player.osc0[8] ));
 sg13g2_a221oi_1 _5754_ (.B2(_2239_),
    .C1(_2242_),
    .B1(_2116_),
    .A1(\dtop.field_top.channel_output[4] ),
    .Y(_2244_),
    .A2(net848));
 sg13g2_a221oi_1 _5755_ (.B2(_2214_),
    .C1(_2114_),
    .B1(_2110_),
    .A1(_1934_),
    .Y(_2245_),
    .A2(net849));
 sg13g2_nand4_1 _5756_ (.B(_2243_),
    .C(_2244_),
    .A(_2237_),
    .Y(_2246_),
    .D(_2245_));
 sg13g2_xnor2_1 _5757_ (.Y(_2247_),
    .A(net847),
    .B(_2246_));
 sg13g2_nor2_1 _5758_ (.A(_2236_),
    .B(_2247_),
    .Y(_2248_));
 sg13g2_xnor2_1 _5759_ (.Y(_2249_),
    .A(_2236_),
    .B(_2247_));
 sg13g2_xnor2_1 _5760_ (.Y(_2250_),
    .A(_2233_),
    .B(_2249_));
 sg13g2_nand2b_1 _5761_ (.Y(_2251_),
    .B(_2250_),
    .A_N(net867));
 sg13g2_a21oi_1 _5762_ (.A1(net1088),
    .A2(net866),
    .Y(_2252_),
    .B1(net1110));
 sg13g2_nand2_1 _5763_ (.Y(_0168_),
    .A(_2251_),
    .B(_2252_));
 sg13g2_a22oi_1 _5764_ (.Y(_2253_),
    .B1(net880),
    .B2(\dtop.field_top.player.out_acc[5] ),
    .A2(net874),
    .A1(\dtop.field_top.channel_output[5] ));
 sg13g2_nand2_1 _5765_ (.Y(_2254_),
    .A(net876),
    .B(_2253_));
 sg13g2_a221oi_1 _5766_ (.B2(\dtop.field_top.channel_output[6] ),
    .C1(_2254_),
    .B1(net873),
    .A1(\dtop.field_top.channel_output[7] ),
    .Y(_2255_),
    .A2(net881));
 sg13g2_a22oi_1 _5767_ (.Y(_2256_),
    .B1(net848),
    .B2(\dtop.field_top.channel_output[5] ),
    .A2(net849),
    .A1(_1936_));
 sg13g2_and2_1 _5768_ (.A(_2132_),
    .B(_2168_),
    .X(_2257_));
 sg13g2_o21ai_1 _5769_ (.B1(_2148_),
    .Y(_2258_),
    .A1(_2212_),
    .A2(_2257_));
 sg13g2_nand2_1 _5770_ (.Y(_2259_),
    .A(\dtop.field_top.player.controller.timer[2] ),
    .B(_1866_));
 sg13g2_a22oi_1 _5771_ (.Y(_2260_),
    .B1(net949),
    .B2(\dtop.field_top.player.controller.timer[0] ),
    .A2(net939),
    .A1(_0089_));
 sg13g2_nand3_1 _5772_ (.B(_2259_),
    .C(_2260_),
    .A(_2116_),
    .Y(_2261_));
 sg13g2_nand2b_1 _5773_ (.Y(_2262_),
    .B(_2096_),
    .A_N(net1078));
 sg13g2_a21oi_1 _5774_ (.A1(_2123_),
    .A2(_2258_),
    .Y(_2263_),
    .B1(_2114_));
 sg13g2_nand4_1 _5775_ (.B(_2261_),
    .C(_2262_),
    .A(_2256_),
    .Y(_2264_),
    .D(_2263_));
 sg13g2_a21oi_1 _5776_ (.A1(_2824_),
    .A2(_2105_),
    .Y(_2265_),
    .B1(_2264_));
 sg13g2_o21ai_1 _5777_ (.B1(_2265_),
    .Y(_2266_),
    .A1(\dtop.field_top.player.controller.timer[1] ),
    .A2(_2111_));
 sg13g2_xor2_1 _5778_ (.B(_2266_),
    .A(net847),
    .X(_2267_));
 sg13g2_nor2b_1 _5779_ (.A(_2255_),
    .B_N(_2267_),
    .Y(_2268_));
 sg13g2_xor2_1 _5780_ (.B(_2267_),
    .A(_2255_),
    .X(_2269_));
 sg13g2_nor2_1 _5781_ (.A(_2227_),
    .B(_2248_),
    .Y(_2270_));
 sg13g2_a22oi_1 _5782_ (.Y(_2271_),
    .B1(_2270_),
    .B2(_2229_),
    .A2(_2247_),
    .A1(_2236_));
 sg13g2_a221oi_1 _5783_ (.B2(_2229_),
    .C1(_2269_),
    .B1(_2270_),
    .A1(_2236_),
    .Y(_2272_),
    .A2(_2247_));
 sg13g2_xor2_1 _5784_ (.B(_2271_),
    .A(_2269_),
    .X(_2273_));
 sg13g2_a21oi_1 _5785_ (.A1(net1083),
    .A2(net867),
    .Y(_2274_),
    .B1(net1110));
 sg13g2_o21ai_1 _5786_ (.B1(_2274_),
    .Y(_0169_),
    .A1(net866),
    .A2(_2273_));
 sg13g2_a22oi_1 _5787_ (.Y(_2275_),
    .B1(net880),
    .B2(\dtop.field_top.player.out_acc[6] ),
    .A2(net874),
    .A1(\dtop.field_top.channel_output[6] ));
 sg13g2_nand2_1 _5788_ (.Y(_2276_),
    .A(net876),
    .B(_2275_));
 sg13g2_a221oi_1 _5789_ (.B2(\dtop.field_top.channel_output[7] ),
    .C1(_2276_),
    .B1(net873),
    .A1(\dtop.field_top.channel_output[2] ),
    .Y(_2277_),
    .A2(net881));
 sg13g2_a21o_1 _5790_ (.A2(_2147_),
    .A1(_2132_),
    .B1(_2140_),
    .X(_2278_));
 sg13g2_a21oi_1 _5791_ (.A1(_2171_),
    .A2(_2278_),
    .Y(_2279_),
    .B1(_2124_));
 sg13g2_nand3_1 _5792_ (.B(_1796_),
    .C(_1835_),
    .A(_1620_),
    .Y(_2280_));
 sg13g2_or4_1 _5793_ (.A(_1513_),
    .B(net978),
    .C(_1577_),
    .D(_1625_),
    .X(_2281_));
 sg13g2_a21oi_2 _5794_ (.B1(_1653_),
    .Y(_2282_),
    .A2(_2281_),
    .A1(_2280_));
 sg13g2_nor2_1 _5795_ (.A(net1094),
    .B(_2282_),
    .Y(_2283_));
 sg13g2_nor2_1 _5796_ (.A(net950),
    .B(_2283_),
    .Y(_2284_));
 sg13g2_a221oi_1 _5797_ (.B2(_2927_),
    .C1(_2284_),
    .B1(net950),
    .A1(_1495_),
    .Y(_2285_),
    .A2(net964));
 sg13g2_a21oi_1 _5798_ (.A1(_0090_),
    .A2(net939),
    .Y(_2286_),
    .B1(_2285_));
 sg13g2_nand2_1 _5799_ (.Y(_2287_),
    .A(net1012),
    .B(_2096_));
 sg13g2_nand2b_1 _5800_ (.Y(_2288_),
    .B(net849),
    .A_N(_1939_));
 sg13g2_a221oi_1 _5801_ (.B2(_2286_),
    .C1(_2279_),
    .B1(_2116_),
    .A1(\dtop.field_top.channel_output[6] ),
    .Y(_2289_),
    .A2(net848));
 sg13g2_nand4_1 _5802_ (.B(_2287_),
    .C(_2288_),
    .A(_2115_),
    .Y(_2290_),
    .D(_2289_));
 sg13g2_a21oi_1 _5803_ (.A1(_2823_),
    .A2(_2105_),
    .Y(_2291_),
    .B1(_2290_));
 sg13g2_o21ai_1 _5804_ (.B1(_2291_),
    .Y(_2292_),
    .A1(\dtop.field_top.player.controller.timer[2] ),
    .A2(_2111_));
 sg13g2_xor2_1 _5805_ (.B(_2292_),
    .A(net847),
    .X(_2293_));
 sg13g2_nand2b_1 _5806_ (.Y(_2294_),
    .B(_2293_),
    .A_N(_2277_));
 sg13g2_xor2_1 _5807_ (.B(_2293_),
    .A(_2277_),
    .X(_2295_));
 sg13g2_inv_1 _5808_ (.Y(_2296_),
    .A(_2295_));
 sg13g2_nor3_1 _5809_ (.A(_2268_),
    .B(_2272_),
    .C(_2296_),
    .Y(_2297_));
 sg13g2_o21ai_1 _5810_ (.B1(_2296_),
    .Y(_2298_),
    .A1(_2268_),
    .A2(_2272_));
 sg13g2_nand2b_2 _5811_ (.Y(_2299_),
    .B(_2298_),
    .A_N(_2297_));
 sg13g2_a21oi_1 _5812_ (.A1(net1075),
    .A2(net866),
    .Y(_2300_),
    .B1(net1110));
 sg13g2_o21ai_1 _5813_ (.B1(_2300_),
    .Y(_0170_),
    .A1(net866),
    .A2(_2299_));
 sg13g2_a22oi_1 _5814_ (.Y(_2301_),
    .B1(net880),
    .B2(\dtop.field_top.player.out_acc[7] ),
    .A2(net874),
    .A1(\dtop.field_top.channel_output[7] ));
 sg13g2_nand2_1 _5815_ (.Y(_2302_),
    .A(net876),
    .B(_2301_));
 sg13g2_a221oi_1 _5816_ (.B2(\dtop.field_top.channel_output[8] ),
    .C1(_2302_),
    .B1(_2047_),
    .A1(\dtop.field_top.channel_output[9] ),
    .Y(_2303_),
    .A2(net882));
 sg13g2_nand2_1 _5817_ (.Y(_2304_),
    .A(_2110_),
    .B(_2284_));
 sg13g2_nand2_1 _5818_ (.Y(_2305_),
    .A(\dtop.field_top.channel_output[7] ),
    .B(net848));
 sg13g2_nand2b_1 _5819_ (.Y(_2306_),
    .B(net849),
    .A_N(_1932_));
 sg13g2_nor2b_1 _5820_ (.A(net1065),
    .B_N(_2096_),
    .Y(_2307_));
 sg13g2_o21ai_1 _5821_ (.B1(_2115_),
    .Y(_2308_),
    .A1(\dtop.field_top.player.osc0[11] ),
    .A2(_2091_));
 sg13g2_nand2_1 _5822_ (.Y(_2309_),
    .A(\dtop.field_top.player.controller.ppos[0] ),
    .B(_2282_));
 sg13g2_and2_1 _5823_ (.A(net1021),
    .B(_1587_),
    .X(_2310_));
 sg13g2_nor2_1 _5824_ (.A(_1607_),
    .B(_2310_),
    .Y(_2311_));
 sg13g2_o21ai_1 _5825_ (.B1(_2311_),
    .Y(_2312_),
    .A1(_1575_),
    .A2(_1578_));
 sg13g2_nor4_2 _5826_ (.A(net1067),
    .B(\dtop.field_top.player.controller.ppos[2] ),
    .C(_1550_),
    .Y(_2313_),
    .D(_1742_));
 sg13g2_nor2_1 _5827_ (.A(net976),
    .B(_2313_),
    .Y(_2314_));
 sg13g2_a21oi_1 _5828_ (.A1(_1736_),
    .A2(_1845_),
    .Y(_2315_),
    .B1(_1771_));
 sg13g2_a21oi_1 _5829_ (.A1(_1588_),
    .A2(_2314_),
    .Y(_2316_),
    .B1(_2315_));
 sg13g2_nand3_1 _5830_ (.B(_2312_),
    .C(_2316_),
    .A(_1533_),
    .Y(_2317_));
 sg13g2_a21oi_1 _5831_ (.A1(net1072),
    .A2(_1611_),
    .Y(_2318_),
    .B1(_1641_));
 sg13g2_or3_1 _5832_ (.A(net1077),
    .B(\dtop.field_top.player.controller.ppos[2] ),
    .C(_1608_),
    .X(_2319_));
 sg13g2_nand3_1 _5833_ (.B(net982),
    .C(_2319_),
    .A(net1019),
    .Y(_2320_));
 sg13g2_a221oi_1 _5834_ (.B2(_1801_),
    .C1(net1068),
    .B1(net984),
    .A1(net1071),
    .Y(_2321_),
    .A2(_1549_));
 sg13g2_a21oi_1 _5835_ (.A1(_2320_),
    .A2(_2321_),
    .Y(_2322_),
    .B1(_2318_));
 sg13g2_nand2_1 _5836_ (.Y(_2323_),
    .A(net972),
    .B(_1620_));
 sg13g2_o21ai_1 _5837_ (.B1(_2323_),
    .Y(_2324_),
    .A1(_1526_),
    .A2(net972));
 sg13g2_nand3_1 _5838_ (.B(_1609_),
    .C(_2324_),
    .A(net1012),
    .Y(_2325_));
 sg13g2_o21ai_1 _5839_ (.B1(_2325_),
    .Y(_2326_),
    .A1(_1607_),
    .A2(_2322_));
 sg13g2_nand2_1 _5840_ (.Y(_2327_),
    .A(net977),
    .B(_2313_));
 sg13g2_and3_1 _5841_ (.X(_2328_),
    .A(net1022),
    .B(net976),
    .C(_1752_));
 sg13g2_a221oi_1 _5842_ (.B2(net1063),
    .C1(_2328_),
    .B1(_2327_),
    .A1(net973),
    .Y(_2329_),
    .A2(_1732_));
 sg13g2_a221oi_1 _5843_ (.B2(_1624_),
    .C1(_1539_),
    .B1(_2329_),
    .A1(_1605_),
    .Y(_2330_),
    .A2(_2326_));
 sg13g2_a22oi_1 _5844_ (.Y(_2331_),
    .B1(_1562_),
    .B2(_1581_),
    .A2(_1548_),
    .A1(net1066));
 sg13g2_nor3_1 _5845_ (.A(\dtop.field_top.player.controller.ppos[6] ),
    .B(_1574_),
    .C(_2331_),
    .Y(_2332_));
 sg13g2_or3_1 _5846_ (.A(net1064),
    .B(net1065),
    .C(_1549_),
    .X(_2333_));
 sg13g2_a21oi_1 _5847_ (.A1(_1551_),
    .A2(_2333_),
    .Y(_2334_),
    .B1(_1545_));
 sg13g2_a21oi_1 _5848_ (.A1(net976),
    .A2(_2332_),
    .Y(_2335_),
    .B1(_2334_));
 sg13g2_a22oi_1 _5849_ (.Y(_2336_),
    .B1(_2335_),
    .B2(_1539_),
    .A2(_2330_),
    .A1(_2317_));
 sg13g2_mux2_1 _5850_ (.A0(_2836_),
    .A1(_2336_),
    .S(net943),
    .X(_2337_));
 sg13g2_nand2_1 _5851_ (.Y(_2338_),
    .A(_2836_),
    .B(_2337_));
 sg13g2_xnor2_1 _5852_ (.Y(_2339_),
    .A(net1091),
    .B(_2337_));
 sg13g2_xnor2_1 _5853_ (.Y(_2340_),
    .A(_2309_),
    .B(_2339_));
 sg13g2_nor2_1 _5854_ (.A(net950),
    .B(_2340_),
    .Y(_2341_));
 sg13g2_a21oi_1 _5855_ (.A1(_2926_),
    .A2(net949),
    .Y(_2342_),
    .B1(_2341_));
 sg13g2_a221oi_1 _5856_ (.B2(net946),
    .C1(_2117_),
    .B1(_2342_),
    .A1(\dtop.field_top.player.controller.timer[0] ),
    .Y(_2343_),
    .A2(net939));
 sg13g2_nand2b_1 _5857_ (.Y(_2344_),
    .B(_2132_),
    .A_N(_2147_));
 sg13g2_a21oi_1 _5858_ (.A1(_2139_),
    .A2(_2344_),
    .Y(_2345_),
    .B1(_2124_));
 sg13g2_nor4_1 _5859_ (.A(_2307_),
    .B(_2308_),
    .C(_2343_),
    .D(_2345_),
    .Y(_2346_));
 sg13g2_nand4_1 _5860_ (.B(_2305_),
    .C(_2306_),
    .A(_2304_),
    .Y(_2347_),
    .D(_2346_));
 sg13g2_xor2_1 _5861_ (.B(_2347_),
    .A(_2107_),
    .X(_2348_));
 sg13g2_nor2b_1 _5862_ (.A(_2303_),
    .B_N(_2348_),
    .Y(_2349_));
 sg13g2_xor2_1 _5863_ (.B(_2348_),
    .A(_2303_),
    .X(_2350_));
 sg13g2_a21oi_1 _5864_ (.A1(_2294_),
    .A2(_2298_),
    .Y(_2351_),
    .B1(_2350_));
 sg13g2_nand3_1 _5865_ (.B(_2298_),
    .C(_2350_),
    .A(_2294_),
    .Y(_2352_));
 sg13g2_nand2b_2 _5866_ (.Y(_2353_),
    .B(_2352_),
    .A_N(_2351_));
 sg13g2_a21oi_1 _5867_ (.A1(net1069),
    .A2(net866),
    .Y(_2354_),
    .B1(net1110));
 sg13g2_o21ai_1 _5868_ (.B1(_2354_),
    .Y(_0171_),
    .A1(net866),
    .A2(_2353_));
 sg13g2_a22oi_1 _5869_ (.Y(_2355_),
    .B1(_2049_),
    .B2(\dtop.field_top.player.out_acc[8] ),
    .A2(net874),
    .A1(\dtop.field_top.channel_output[8] ));
 sg13g2_nand2_1 _5870_ (.Y(_2356_),
    .A(_2044_),
    .B(_2355_));
 sg13g2_a221oi_1 _5871_ (.B2(\dtop.field_top.channel_output[9] ),
    .C1(_2356_),
    .B1(net873),
    .A1(\dtop.field_top.channel_output[4] ),
    .Y(_2357_),
    .A2(net881));
 sg13g2_nand2b_1 _5872_ (.Y(_2358_),
    .B(_2139_),
    .A_N(_2344_));
 sg13g2_a21oi_1 _5873_ (.A1(_2123_),
    .A2(_2358_),
    .Y(_2359_),
    .B1(_2114_));
 sg13g2_nor2_1 _5874_ (.A(net1070),
    .B(_2323_),
    .Y(_2360_));
 sg13g2_nand3_1 _5875_ (.B(_1610_),
    .C(_2360_),
    .A(_1605_),
    .Y(_2361_));
 sg13g2_nor3_1 _5876_ (.A(net1076),
    .B(_1575_),
    .C(_1627_),
    .Y(_2362_));
 sg13g2_nor3_1 _5877_ (.A(net1022),
    .B(_1600_),
    .C(_2362_),
    .Y(_2363_));
 sg13g2_nor3_1 _5878_ (.A(net1083),
    .B(net1091),
    .C(_1513_),
    .Y(_2364_));
 sg13g2_nand2b_1 _5879_ (.Y(_2365_),
    .B(_1634_),
    .A_N(_2364_));
 sg13g2_o21ai_1 _5880_ (.B1(net972),
    .Y(_2366_),
    .A1(_2363_),
    .A2(_2365_));
 sg13g2_nand3b_1 _5881_ (.B(_1745_),
    .C(_2366_),
    .Y(_2367_),
    .A_N(_1646_));
 sg13g2_o21ai_1 _5882_ (.B1(net982),
    .Y(_2368_),
    .A1(net1072),
    .A2(_1567_));
 sg13g2_o21ai_1 _5883_ (.B1(_2368_),
    .Y(_2369_),
    .A1(_1612_),
    .A2(net982));
 sg13g2_o21ai_1 _5884_ (.B1(_1510_),
    .Y(_2370_),
    .A1(_1755_),
    .A2(_2369_));
 sg13g2_a21oi_1 _5885_ (.A1(_1584_),
    .A2(_1639_),
    .Y(_2371_),
    .B1(_1553_));
 sg13g2_o21ai_1 _5886_ (.B1(_2371_),
    .Y(_2372_),
    .A1(net1019),
    .A2(_1611_));
 sg13g2_nor3_1 _5887_ (.A(net1080),
    .B(_1575_),
    .C(_1627_),
    .Y(_2373_));
 sg13g2_a21oi_1 _5888_ (.A1(_1598_),
    .A2(_1640_),
    .Y(_2374_),
    .B1(net1023));
 sg13g2_nand2b_1 _5889_ (.Y(_2375_),
    .B(_2374_),
    .A_N(_2373_));
 sg13g2_nand4_1 _5890_ (.B(_2370_),
    .C(_2372_),
    .A(_1796_),
    .Y(_2376_),
    .D(_2375_));
 sg13g2_nand4_1 _5891_ (.B(_2361_),
    .C(_2367_),
    .A(net943),
    .Y(_2377_),
    .D(_2376_));
 sg13g2_a221oi_1 _5892_ (.B2(net977),
    .C1(_1603_),
    .B1(_1814_),
    .A1(_1616_),
    .Y(_2378_),
    .A2(_1773_));
 sg13g2_nand3_1 _5893_ (.B(_1555_),
    .C(_1560_),
    .A(\dtop.field_top.player.controller.ppos[6] ),
    .Y(_2379_));
 sg13g2_nor3_1 _5894_ (.A(_1540_),
    .B(net974),
    .C(_2379_),
    .Y(_2380_));
 sg13g2_nor3_1 _5895_ (.A(_2377_),
    .B(_2378_),
    .C(_2380_),
    .Y(_2381_));
 sg13g2_nor2_1 _5896_ (.A(_2130_),
    .B(_2381_),
    .Y(_2382_));
 sg13g2_xnor2_1 _5897_ (.Y(_2383_),
    .A(\dtop.field_top.player.controller.ppos[2] ),
    .B(_2382_));
 sg13g2_and3_1 _5898_ (.X(_2384_),
    .A(_2309_),
    .B(_2338_),
    .C(_2383_));
 sg13g2_a21oi_1 _5899_ (.A1(_2309_),
    .A2(_2338_),
    .Y(_2385_),
    .B1(_2383_));
 sg13g2_nor2_2 _5900_ (.A(_2384_),
    .B(_2385_),
    .Y(_2386_));
 sg13g2_nand2b_1 _5901_ (.Y(_2387_),
    .B(_2386_),
    .A_N(_1659_));
 sg13g2_nor2_1 _5902_ (.A(_1664_),
    .B(_2283_),
    .Y(_2388_));
 sg13g2_nor2_2 _5903_ (.A(net950),
    .B(_2386_),
    .Y(_2389_));
 sg13g2_a21oi_1 _5904_ (.A1(_2387_),
    .A2(_2388_),
    .Y(_2390_),
    .B1(_2389_));
 sg13g2_a22oi_1 _5905_ (.Y(_2391_),
    .B1(_2390_),
    .B2(net946),
    .A2(net940),
    .A1(\dtop.field_top.player.controller.timer[1] ));
 sg13g2_a22oi_1 _5906_ (.Y(_2392_),
    .B1(_2116_),
    .B2(_2391_),
    .A2(net848),
    .A1(\dtop.field_top.channel_output[8] ));
 sg13g2_a22oi_1 _5907_ (.Y(_2393_),
    .B1(_2110_),
    .B2(_2341_),
    .A2(net849),
    .A1(_1948_));
 sg13g2_nand2b_1 _5908_ (.Y(_2394_),
    .B(_2105_),
    .A_N(\dtop.field_top.player.osc0[12] ));
 sg13g2_nand4_1 _5909_ (.B(_2392_),
    .C(_2393_),
    .A(_2359_),
    .Y(_2395_),
    .D(_2394_));
 sg13g2_a21oi_2 _5910_ (.B1(_2395_),
    .Y(_2396_),
    .A2(_2096_),
    .A1(_2854_));
 sg13g2_xnor2_1 _5911_ (.Y(_2397_),
    .A(net847),
    .B(_2396_));
 sg13g2_nor2b_1 _5912_ (.A(_2357_),
    .B_N(_2397_),
    .Y(_2398_));
 sg13g2_inv_1 _5913_ (.Y(_2399_),
    .A(_2398_));
 sg13g2_xor2_1 _5914_ (.B(_2397_),
    .A(_2357_),
    .X(_2400_));
 sg13g2_inv_1 _5915_ (.Y(_2401_),
    .A(_2400_));
 sg13g2_nor3_1 _5916_ (.A(_2349_),
    .B(_2351_),
    .C(_2401_),
    .Y(_2402_));
 sg13g2_o21ai_1 _5917_ (.B1(_2401_),
    .Y(_2403_),
    .A1(_2349_),
    .A2(_2351_));
 sg13g2_nand2b_2 _5918_ (.Y(_2404_),
    .B(_2403_),
    .A_N(_2402_));
 sg13g2_nand2b_1 _5919_ (.Y(_2405_),
    .B(_2404_),
    .A_N(net866));
 sg13g2_a21oi_1 _5920_ (.A1(net1024),
    .A2(net866),
    .Y(_2406_),
    .B1(net1110));
 sg13g2_and2_1 _5921_ (.A(_2405_),
    .B(_2406_),
    .X(_0172_));
 sg13g2_nand2_1 _5922_ (.Y(_2407_),
    .A(net1028),
    .B(_2045_));
 sg13g2_o21ai_1 _5923_ (.B1(_2044_),
    .Y(_2408_),
    .A1(_2048_),
    .A2(_2407_));
 sg13g2_a21oi_1 _5924_ (.A1(\dtop.field_top.player.out_acc[9] ),
    .A2(net880),
    .Y(_2409_),
    .B1(_2408_));
 sg13g2_a22oi_1 _5925_ (.Y(_2410_),
    .B1(net875),
    .B2(\dtop.field_top.channel_output[9] ),
    .A2(net882),
    .A1(\dtop.field_top.channel_output[3] ));
 sg13g2_nand3_1 _5926_ (.B(_2047_),
    .C(_2048_),
    .A(net1028),
    .Y(_2411_));
 sg13g2_nand3_1 _5927_ (.B(_2410_),
    .C(_2411_),
    .A(_2409_),
    .Y(_2412_));
 sg13g2_a21oi_2 _5928_ (.B1(_2385_),
    .Y(_2413_),
    .A2(_2382_),
    .A1(_2835_));
 sg13g2_o21ai_1 _5929_ (.B1(_2834_),
    .Y(_2414_),
    .A1(\dtop.field_top.player.controller.ppos[2] ),
    .A2(_1741_));
 sg13g2_a21oi_1 _5930_ (.A1(_1736_),
    .A2(_2414_),
    .Y(_2415_),
    .B1(_1771_));
 sg13g2_nor3_1 _5931_ (.A(_1607_),
    .B(_1813_),
    .C(_2310_),
    .Y(_2416_));
 sg13g2_nor3_1 _5932_ (.A(_1603_),
    .B(_2415_),
    .C(_2416_),
    .Y(_2417_));
 sg13g2_nor2_1 _5933_ (.A(net1019),
    .B(net1087),
    .Y(_2418_));
 sg13g2_a21oi_1 _5934_ (.A1(net1074),
    .A2(_1785_),
    .Y(_2419_),
    .B1(_1526_));
 sg13g2_a22oi_1 _5935_ (.Y(_2420_),
    .B1(_1640_),
    .B2(_2419_),
    .A2(_1591_),
    .A1(_1552_));
 sg13g2_o21ai_1 _5936_ (.B1(_2420_),
    .Y(_2421_),
    .A1(_1807_),
    .A2(_2418_));
 sg13g2_a21oi_1 _5937_ (.A1(net983),
    .A2(_1808_),
    .Y(_2422_),
    .B1(_2421_));
 sg13g2_nor2b_1 _5938_ (.A(_2422_),
    .B_N(_1796_),
    .Y(_2423_));
 sg13g2_a21oi_1 _5939_ (.A1(_1510_),
    .A2(_1785_),
    .Y(_2424_),
    .B1(_1633_));
 sg13g2_o21ai_1 _5940_ (.B1(_2424_),
    .Y(_2425_),
    .A1(net1022),
    .A2(_1630_));
 sg13g2_a221oi_1 _5941_ (.B2(net974),
    .C1(_1646_),
    .B1(_2425_),
    .A1(_1606_),
    .Y(_2426_),
    .A2(_1643_));
 sg13g2_or4_1 _5942_ (.A(_1653_),
    .B(_2417_),
    .C(_2423_),
    .D(_2426_),
    .X(_2427_));
 sg13g2_o21ai_1 _5943_ (.B1(_2427_),
    .Y(_2428_),
    .A1(_2834_),
    .A2(net943));
 sg13g2_xnor2_1 _5944_ (.Y(_2429_),
    .A(net1078),
    .B(_2428_));
 sg13g2_a21oi_1 _5945_ (.A1(_2413_),
    .A2(_2429_),
    .Y(_2430_),
    .B1(net950));
 sg13g2_o21ai_1 _5946_ (.B1(_2430_),
    .Y(_2431_),
    .A1(_2413_),
    .A2(_2429_));
 sg13g2_nor2_1 _5947_ (.A(_1669_),
    .B(_2340_),
    .Y(_2432_));
 sg13g2_nor2_1 _5948_ (.A(net951),
    .B(_2432_),
    .Y(_2433_));
 sg13g2_a221oi_1 _5949_ (.B2(_2433_),
    .C1(_2117_),
    .B1(_2431_),
    .A1(\dtop.field_top.player.controller.timer[2] ),
    .Y(_2434_),
    .A2(net939));
 sg13g2_a221oi_1 _5950_ (.B2(\dtop.field_top.channel_output[9] ),
    .C1(_2434_),
    .B1(net848),
    .A1(_1946_),
    .Y(_2435_),
    .A2(net849));
 sg13g2_o21ai_1 _5951_ (.B1(_2115_),
    .Y(_2436_),
    .A1(net1094),
    .A2(_2091_));
 sg13g2_a21oi_1 _5952_ (.A1(_2925_),
    .A2(_2096_),
    .Y(_2437_),
    .B1(_2436_));
 sg13g2_and2_1 _5953_ (.A(_2435_),
    .B(_2437_),
    .X(_2438_));
 sg13g2_xnor2_1 _5954_ (.Y(_2439_),
    .A(net847),
    .B(_2438_));
 sg13g2_nand2_1 _5955_ (.Y(_2440_),
    .A(_2412_),
    .B(_2439_));
 sg13g2_inv_1 _5956_ (.Y(_2441_),
    .A(_2440_));
 sg13g2_xor2_1 _5957_ (.B(_2439_),
    .A(_2412_),
    .X(_2442_));
 sg13g2_inv_1 _5958_ (.Y(_2443_),
    .A(_2442_));
 sg13g2_a21oi_2 _5959_ (.B1(_2443_),
    .Y(_2444_),
    .A2(_2403_),
    .A1(_2399_));
 sg13g2_nand3_1 _5960_ (.B(_2403_),
    .C(_2443_),
    .A(_2399_),
    .Y(_2445_));
 sg13g2_nand2b_2 _5961_ (.Y(_2446_),
    .B(_2445_),
    .A_N(_2444_));
 sg13g2_a21oi_1 _5962_ (.A1(net509),
    .A2(net867),
    .Y(_2447_),
    .B1(net1111));
 sg13g2_o21ai_1 _5963_ (.B1(_2447_),
    .Y(_0173_),
    .A1(net867),
    .A2(_2446_));
 sg13g2_nor2_1 _5964_ (.A(_2441_),
    .B(_2444_),
    .Y(_2448_));
 sg13g2_and3_1 _5965_ (.X(_2449_),
    .A(\dtop.field_top.channel_output[0] ),
    .B(_2043_),
    .C(_2045_));
 sg13g2_a221oi_1 _5966_ (.B2(net1028),
    .C1(_2449_),
    .B1(net875),
    .A1(\dtop.field_top.channel_output[8] ),
    .Y(_2450_),
    .A2(net882));
 sg13g2_nand2_1 _5967_ (.Y(_2451_),
    .A(_2409_),
    .B(_2450_));
 sg13g2_mux2_1 _5968_ (.A0(net847),
    .A1(_1992_),
    .S(_2106_),
    .X(_2452_));
 sg13g2_nand2b_1 _5969_ (.Y(_2453_),
    .B(_2452_),
    .A_N(_2451_));
 sg13g2_inv_1 _5970_ (.Y(_2454_),
    .A(_2453_));
 sg13g2_nand2b_1 _5971_ (.Y(_2455_),
    .B(_2451_),
    .A_N(_2452_));
 sg13g2_nand2_1 _5972_ (.Y(_2456_),
    .A(_2453_),
    .B(_2455_));
 sg13g2_inv_1 _5973_ (.Y(_2457_),
    .A(_2456_));
 sg13g2_nor3_1 _5974_ (.A(_2441_),
    .B(_2444_),
    .C(_2457_),
    .Y(_2458_));
 sg13g2_o21ai_1 _5975_ (.B1(_2457_),
    .Y(_2459_),
    .A1(_2441_),
    .A2(_2444_));
 sg13g2_nand2b_2 _5976_ (.Y(_2460_),
    .B(_2459_),
    .A_N(_2458_));
 sg13g2_a21oi_1 _5977_ (.A1(net690),
    .A2(net867),
    .Y(_2461_),
    .B1(net1110));
 sg13g2_o21ai_1 _5978_ (.B1(_2461_),
    .Y(_0174_),
    .A1(net867),
    .A2(_2460_));
 sg13g2_nor2_1 _5979_ (.A(_1125_),
    .B(net979),
    .Y(_2462_));
 sg13g2_a21oi_1 _5980_ (.A1(net355),
    .A2(net947),
    .Y(_2463_),
    .B1(_2462_));
 sg13g2_inv_1 _5981_ (.Y(_0175_),
    .A(_2463_));
 sg13g2_mux2_1 _5982_ (.A0(net372),
    .A1(_1232_),
    .S(net1059),
    .X(_0176_));
 sg13g2_nor2_1 _5983_ (.A(_0966_),
    .B(_0977_),
    .Y(_2464_));
 sg13g2_xnor2_1 _5984_ (.Y(_2465_),
    .A(_0966_),
    .B(_0977_));
 sg13g2_nand2_1 _5985_ (.Y(_2466_),
    .A(net622),
    .B(_0735_));
 sg13g2_o21ai_1 _5986_ (.B1(_2466_),
    .Y(_0177_),
    .A1(_0735_),
    .A2(_2465_));
 sg13g2_xnor2_1 _5987_ (.Y(_2467_),
    .A(_0996_),
    .B(_2464_));
 sg13g2_mux2_1 _5988_ (.A0(_2467_),
    .A1(net662),
    .S(_0735_),
    .X(_0178_));
 sg13g2_nand2_1 _5989_ (.Y(_2468_),
    .A(_3050_),
    .B(net970));
 sg13g2_o21ai_1 _5990_ (.B1(_2468_),
    .Y(_2469_),
    .A1(_3052_),
    .A2(net971));
 sg13g2_nand2_1 _5991_ (.Y(_2470_),
    .A(_0734_),
    .B(_2469_));
 sg13g2_xnor2_1 _5992_ (.Y(_2471_),
    .A(_0996_),
    .B(_1015_));
 sg13g2_mux2_1 _5993_ (.A0(_2471_),
    .A1(net701),
    .S(_2470_),
    .X(_0179_));
 sg13g2_nor2_1 _5994_ (.A(net971),
    .B(_3106_),
    .Y(_2472_));
 sg13g2_o21ai_1 _5995_ (.B1(_2468_),
    .Y(_2473_),
    .A1(net970),
    .A2(_3106_));
 sg13g2_o21ai_1 _5996_ (.B1(_3052_),
    .Y(_2474_),
    .A1(_3056_),
    .A2(_3107_));
 sg13g2_o21ai_1 _5997_ (.B1(_0734_),
    .Y(_2475_),
    .A1(_2473_),
    .A2(_2474_));
 sg13g2_mux2_1 _5998_ (.A0(_1015_),
    .A1(net696),
    .S(_2475_),
    .X(_0180_));
 sg13g2_nor2_2 _5999_ (.A(_3009_),
    .B(net986),
    .Y(_2476_));
 sg13g2_nand2_2 _6000_ (.Y(_2477_),
    .A(_3010_),
    .B(net989));
 sg13g2_nand2_1 _6001_ (.Y(_2478_),
    .A(net365),
    .B(net959));
 sg13g2_o21ai_1 _6002_ (.B1(_2478_),
    .Y(_0181_),
    .A1(_2918_),
    .A2(net959));
 sg13g2_nand2_1 _6003_ (.Y(_2479_),
    .A(net331),
    .B(net959));
 sg13g2_o21ai_1 _6004_ (.B1(_2479_),
    .Y(_0182_),
    .A1(_2919_),
    .A2(net959));
 sg13g2_mux2_1 _6005_ (.A0(net422),
    .A1(net418),
    .S(net959),
    .X(_0183_));
 sg13g2_mux2_1 _6006_ (.A0(net403),
    .A1(net400),
    .S(net959),
    .X(_0184_));
 sg13g2_nand2_1 _6007_ (.Y(_2480_),
    .A(net302),
    .B(net960));
 sg13g2_o21ai_1 _6008_ (.B1(_2480_),
    .Y(_0185_),
    .A1(_2920_),
    .A2(net960));
 sg13g2_mux2_1 _6009_ (.A0(net569),
    .A1(net416),
    .S(net960),
    .X(_0186_));
 sg13g2_mux2_1 _6010_ (.A0(net481),
    .A1(net404),
    .S(net963),
    .X(_0187_));
 sg13g2_mux2_1 _6011_ (.A0(\dtop.field_top.last_wave[7] ),
    .A1(net312),
    .S(net962),
    .X(_0188_));
 sg13g2_nor2_1 _6012_ (.A(net365),
    .B(net960),
    .Y(_2481_));
 sg13g2_a21oi_1 _6013_ (.A1(_2914_),
    .A2(net961),
    .Y(_0189_),
    .B1(_2481_));
 sg13g2_nor2_1 _6014_ (.A(net331),
    .B(net960),
    .Y(_2482_));
 sg13g2_a21oi_1 _6015_ (.A1(_2915_),
    .A2(net959),
    .Y(_0190_),
    .B1(_2482_));
 sg13g2_mux2_1 _6016_ (.A0(net418),
    .A1(\dtop.field_top.wave[2] ),
    .S(net959),
    .X(_0191_));
 sg13g2_mux2_1 _6017_ (.A0(net400),
    .A1(\dtop.field_top.wave[3] ),
    .S(net960),
    .X(_0192_));
 sg13g2_mux2_1 _6018_ (.A0(net302),
    .A1(net389),
    .S(net961),
    .X(_0193_));
 sg13g2_nor2_1 _6019_ (.A(net416),
    .B(net961),
    .Y(_2483_));
 sg13g2_a21oi_1 _6020_ (.A1(_2916_),
    .A2(net960),
    .Y(_0194_),
    .B1(_2483_));
 sg13g2_nor2_1 _6021_ (.A(net404),
    .B(net963),
    .Y(_2484_));
 sg13g2_a21oi_1 _6022_ (.A1(_2917_),
    .A2(net963),
    .Y(_0195_),
    .B1(_2484_));
 sg13g2_mux2_1 _6023_ (.A0(net312),
    .A1(net386),
    .S(net962),
    .X(_0196_));
 sg13g2_nand2_1 _6024_ (.Y(_2485_),
    .A(_3096_),
    .B(_0433_));
 sg13g2_o21ai_1 _6025_ (.B1(net992),
    .Y(_2486_),
    .A1(_3051_),
    .A2(_3068_));
 sg13g2_nor2b_1 _6026_ (.A(_2485_),
    .B_N(_2486_),
    .Y(_2487_));
 sg13g2_a22oi_1 _6027_ (.Y(_2488_),
    .B1(net990),
    .B2(_3083_),
    .A2(_3078_),
    .A1(net996));
 sg13g2_nand3_1 _6028_ (.B(_3106_),
    .C(_2488_),
    .A(_3094_),
    .Y(_2489_));
 sg13g2_a21oi_1 _6029_ (.A1(_3078_),
    .A2(net990),
    .Y(_2490_),
    .B1(_3108_));
 sg13g2_nand4_1 _6030_ (.B(_3095_),
    .C(_2487_),
    .A(net968),
    .Y(_2491_),
    .D(_2490_));
 sg13g2_or2_1 _6031_ (.X(_2492_),
    .B(_2491_),
    .A(_2489_));
 sg13g2_a221oi_1 _6032_ (.B2(net992),
    .C1(net968),
    .B1(_3070_),
    .A1(net997),
    .Y(_2493_),
    .A2(_3068_));
 sg13g2_o21ai_1 _6033_ (.B1(net993),
    .Y(_2494_),
    .A1(_3070_),
    .A2(_3078_));
 sg13g2_nand4_1 _6034_ (.B(_0433_),
    .C(_2493_),
    .A(_3099_),
    .Y(_2495_),
    .D(_2494_));
 sg13g2_nand3_1 _6035_ (.B(_2492_),
    .C(_2495_),
    .A(_0442_),
    .Y(_2496_));
 sg13g2_inv_1 _6036_ (.Y(_2497_),
    .A(_2496_));
 sg13g2_nand2_1 _6037_ (.Y(_2498_),
    .A(_3033_),
    .B(_2497_));
 sg13g2_nand2_1 _6038_ (.Y(_2499_),
    .A(net367),
    .B(net901));
 sg13g2_nand3_1 _6039_ (.B(_2492_),
    .C(_2495_),
    .A(_0442_),
    .Y(_2500_));
 sg13g2_o21ai_1 _6040_ (.B1(_2499_),
    .Y(_0197_),
    .A1(_2875_),
    .A2(net901));
 sg13g2_mux2_1 _6041_ (.A0(\dtop.field_top.acc[2] ),
    .A1(net541),
    .S(net901),
    .X(_0198_));
 sg13g2_nor2_1 _6042_ (.A(\dtop.field_top.acc[3] ),
    .B(net901),
    .Y(_2501_));
 sg13g2_a21oi_1 _6043_ (.A1(_2923_),
    .A2(net901),
    .Y(_0199_),
    .B1(_2501_));
 sg13g2_nand2_1 _6044_ (.Y(_2502_),
    .A(net432),
    .B(net901));
 sg13g2_o21ai_1 _6045_ (.B1(_2502_),
    .Y(_0200_),
    .A1(_2877_),
    .A2(net902));
 sg13g2_mux2_1 _6046_ (.A0(\dtop.field_top.acc[5] ),
    .A1(net545),
    .S(net901),
    .X(_0201_));
 sg13g2_mux2_1 _6047_ (.A0(\dtop.field_top.acc[6] ),
    .A1(net533),
    .S(net901),
    .X(_0202_));
 sg13g2_nor2_1 _6048_ (.A(\dtop.field_top.acc[7] ),
    .B(net902),
    .Y(_2503_));
 sg13g2_a21oi_1 _6049_ (.A1(_2922_),
    .A2(net902),
    .Y(_0203_),
    .B1(_2503_));
 sg13g2_nor2_1 _6050_ (.A(\dtop.field_top.acc[8] ),
    .B(net903),
    .Y(_2504_));
 sg13g2_a21oi_1 _6051_ (.A1(_2921_),
    .A2(net903),
    .Y(_0204_),
    .B1(_2504_));
 sg13g2_mux2_1 _6052_ (.A0(\dtop.field_top.acc[9] ),
    .A1(net562),
    .S(net903),
    .X(_0205_));
 sg13g2_mux2_1 _6053_ (.A0(\dtop.field_top.acc[10] ),
    .A1(net556),
    .S(net903),
    .X(_0206_));
 sg13g2_nand2_1 _6054_ (.Y(_2505_),
    .A(net333),
    .B(_2477_));
 sg13g2_nand2_1 _6055_ (.Y(_2506_),
    .A(\dtop.field_top.channel_output[3] ),
    .B(net963));
 sg13g2_o21ai_1 _6056_ (.B1(_2505_),
    .Y(_0207_),
    .A1(net877),
    .A2(_2506_));
 sg13g2_nand2_1 _6057_ (.Y(_2507_),
    .A(net375),
    .B(_2477_));
 sg13g2_nand2_1 _6058_ (.Y(_2508_),
    .A(\dtop.field_top.channel_output[4] ),
    .B(net963));
 sg13g2_o21ai_1 _6059_ (.B1(_2507_),
    .Y(_0208_),
    .A1(net877),
    .A2(_2508_));
 sg13g2_nand2_1 _6060_ (.Y(_2509_),
    .A(net537),
    .B(_2477_));
 sg13g2_nand2_1 _6061_ (.Y(_2510_),
    .A(\dtop.field_top.channel_output[5] ),
    .B(net962));
 sg13g2_o21ai_1 _6062_ (.B1(_2509_),
    .Y(_0209_),
    .A1(net877),
    .A2(_2510_));
 sg13g2_nand2_1 _6063_ (.Y(_2511_),
    .A(net616),
    .B(_2477_));
 sg13g2_nand2_1 _6064_ (.Y(_2512_),
    .A(\dtop.field_top.channel_output[6] ),
    .B(net962));
 sg13g2_o21ai_1 _6065_ (.B1(_2511_),
    .Y(_0210_),
    .A1(net877),
    .A2(_2512_));
 sg13g2_nand2_1 _6066_ (.Y(_2513_),
    .A(net389),
    .B(_2477_));
 sg13g2_nand2_1 _6067_ (.Y(_2514_),
    .A(net586),
    .B(net962));
 sg13g2_o21ai_1 _6068_ (.B1(_2513_),
    .Y(_0211_),
    .A1(net877),
    .A2(_2514_));
 sg13g2_nand2_1 _6069_ (.Y(_2515_),
    .A(net438),
    .B(_2477_));
 sg13g2_nand2_1 _6070_ (.Y(_2516_),
    .A(\dtop.field_top.channel_output[8] ),
    .B(net962));
 sg13g2_o21ai_1 _6071_ (.B1(_2515_),
    .Y(_0212_),
    .A1(net877),
    .A2(_2516_));
 sg13g2_nand2_1 _6072_ (.Y(_2517_),
    .A(net342),
    .B(_2477_));
 sg13g2_nand2_1 _6073_ (.Y(_2518_),
    .A(\dtop.field_top.channel_output[9] ),
    .B(net962));
 sg13g2_o21ai_1 _6074_ (.B1(_2517_),
    .Y(_0213_),
    .A1(net877),
    .A2(_2518_));
 sg13g2_nand2_1 _6075_ (.Y(_2519_),
    .A(\dtop.field_top.wave[7] ),
    .B(_2477_));
 sg13g2_nand2_1 _6076_ (.Y(_2520_),
    .A(net327),
    .B(net962));
 sg13g2_o21ai_1 _6077_ (.B1(_2519_),
    .Y(_0214_),
    .A1(net877),
    .A2(_2520_));
 sg13g2_and2_1 _6078_ (.A(net967),
    .B(_2494_),
    .X(_2521_));
 sg13g2_a21oi_1 _6079_ (.A1(net968),
    .A2(_2487_),
    .Y(_2522_),
    .B1(_2521_));
 sg13g2_nand2_1 _6080_ (.Y(_2523_),
    .A(_2497_),
    .B(_2522_));
 sg13g2_nor3_1 _6081_ (.A(net967),
    .B(_2485_),
    .C(_2489_),
    .Y(_2524_));
 sg13g2_a21o_1 _6082_ (.A2(_2493_),
    .A1(_3071_),
    .B1(_2524_),
    .X(_2525_));
 sg13g2_nand3_1 _6083_ (.B(_2522_),
    .C(_2525_),
    .A(_2497_),
    .Y(_2526_));
 sg13g2_mux2_1 _6084_ (.A0(\dtop.field_top.acc[0] ),
    .A1(net390),
    .S(net897),
    .X(_0215_));
 sg13g2_nand2_1 _6085_ (.Y(_2527_),
    .A(net329),
    .B(net897));
 sg13g2_o21ai_1 _6086_ (.B1(_2527_),
    .Y(_0216_),
    .A1(_2875_),
    .A2(net897));
 sg13g2_nand2_1 _6087_ (.Y(_2528_),
    .A(net360),
    .B(net897));
 sg13g2_o21ai_1 _6088_ (.B1(_2528_),
    .Y(_0217_),
    .A1(_2878_),
    .A2(net897));
 sg13g2_nor2_1 _6089_ (.A(\dtop.field_top.acc[3] ),
    .B(net898),
    .Y(_2529_));
 sg13g2_a21oi_1 _6090_ (.A1(_2888_),
    .A2(net898),
    .Y(_0218_),
    .B1(_2529_));
 sg13g2_nand2_1 _6091_ (.Y(_2530_),
    .A(net420),
    .B(net898));
 sg13g2_o21ai_1 _6092_ (.B1(_2530_),
    .Y(_0219_),
    .A1(_2877_),
    .A2(net898));
 sg13g2_nor2_1 _6093_ (.A(\dtop.field_top.acc[5] ),
    .B(net898),
    .Y(_2531_));
 sg13g2_a21oi_1 _6094_ (.A1(_2898_),
    .A2(net898),
    .Y(_0220_),
    .B1(_2531_));
 sg13g2_nor2_1 _6095_ (.A(\dtop.field_top.acc[6] ),
    .B(net897),
    .Y(_2532_));
 sg13g2_a21oi_1 _6096_ (.A1(_2903_),
    .A2(net898),
    .Y(_0221_),
    .B1(_2532_));
 sg13g2_nor2_1 _6097_ (.A(\dtop.field_top.acc[7] ),
    .B(net900),
    .Y(_2533_));
 sg13g2_a21oi_1 _6098_ (.A1(_2908_),
    .A2(net900),
    .Y(_0222_),
    .B1(_2533_));
 sg13g2_mux2_1 _6099_ (.A0(\dtop.field_top.acc[8] ),
    .A1(net495),
    .S(net899),
    .X(_0223_));
 sg13g2_mux2_1 _6100_ (.A0(\dtop.field_top.acc[9] ),
    .A1(net558),
    .S(net899),
    .X(_0224_));
 sg13g2_mux2_1 _6101_ (.A0(\dtop.field_top.acc[10] ),
    .A1(net503),
    .S(net899),
    .X(_0225_));
 sg13g2_mux2_1 _6102_ (.A0(\dtop.field_top.acc[11] ),
    .A1(net392),
    .S(net899),
    .X(_0226_));
 sg13g2_mux2_1 _6103_ (.A0(\dtop.field_top.acc[12] ),
    .A1(net382),
    .S(net899),
    .X(_0227_));
 sg13g2_mux2_1 _6104_ (.A0(\dtop.field_top.acc[13] ),
    .A1(net410),
    .S(net897),
    .X(_0228_));
 sg13g2_mux2_1 _6105_ (.A0(\dtop.field_top.acc[14] ),
    .A1(net387),
    .S(net899),
    .X(_0229_));
 sg13g2_nand2_1 _6106_ (.Y(_2534_),
    .A(net310),
    .B(net899));
 sg13g2_o21ai_1 _6107_ (.B1(_2534_),
    .Y(_0230_),
    .A1(_2881_),
    .A2(net899));
 sg13g2_mux2_1 _6108_ (.A0(\dtop.field_top.acc[16] ),
    .A1(net394),
    .S(net897),
    .X(_0231_));
 sg13g2_or3_1 _6109_ (.A(_2500_),
    .B(_2522_),
    .C(_2525_),
    .X(_2535_));
 sg13g2_mux2_1 _6110_ (.A0(\dtop.field_top.acc[0] ),
    .A1(net457),
    .S(net918),
    .X(_0232_));
 sg13g2_mux2_1 _6111_ (.A0(\dtop.field_top.acc[1] ),
    .A1(net543),
    .S(net918),
    .X(_0233_));
 sg13g2_nand2_1 _6112_ (.Y(_2536_),
    .A(net499),
    .B(net918));
 sg13g2_o21ai_1 _6113_ (.B1(_2536_),
    .Y(_0234_),
    .A1(_2878_),
    .A2(net918));
 sg13g2_mux2_1 _6114_ (.A0(\dtop.field_top.acc[3] ),
    .A1(net593),
    .S(net918),
    .X(_0235_));
 sg13g2_nor2_1 _6115_ (.A(\dtop.field_top.acc[4] ),
    .B(net919),
    .Y(_2537_));
 sg13g2_a21oi_1 _6116_ (.A1(_2895_),
    .A2(net919),
    .Y(_0236_),
    .B1(_2537_));
 sg13g2_mux2_1 _6117_ (.A0(\dtop.field_top.acc[5] ),
    .A1(net623),
    .S(net919),
    .X(_0237_));
 sg13g2_nor2_1 _6118_ (.A(\dtop.field_top.acc[6] ),
    .B(net919),
    .Y(_2538_));
 sg13g2_a21oi_1 _6119_ (.A1(_2906_),
    .A2(net919),
    .Y(_0238_),
    .B1(_2538_));
 sg13g2_mux2_1 _6120_ (.A0(\dtop.field_top.acc[7] ),
    .A1(net605),
    .S(net920),
    .X(_0239_));
 sg13g2_mux2_1 _6121_ (.A0(\dtop.field_top.acc[8] ),
    .A1(net606),
    .S(net920),
    .X(_0240_));
 sg13g2_mux2_1 _6122_ (.A0(\dtop.field_top.acc[9] ),
    .A1(net646),
    .S(net920),
    .X(_0241_));
 sg13g2_mux2_1 _6123_ (.A0(\dtop.field_top.acc[10] ),
    .A1(net577),
    .S(net920),
    .X(_0242_));
 sg13g2_mux2_1 _6124_ (.A0(\dtop.field_top.acc[11] ),
    .A1(net491),
    .S(net918),
    .X(_0243_));
 sg13g2_mux2_1 _6125_ (.A0(\dtop.field_top.acc[12] ),
    .A1(net453),
    .S(_2535_),
    .X(_0244_));
 sg13g2_mux2_1 _6126_ (.A0(\dtop.field_top.acc[13] ),
    .A1(net461),
    .S(net920),
    .X(_0245_));
 sg13g2_mux2_1 _6127_ (.A0(\dtop.field_top.acc[14] ),
    .A1(net449),
    .S(net918),
    .X(_0246_));
 sg13g2_mux2_1 _6128_ (.A0(\dtop.field_top.acc[15] ),
    .A1(net505),
    .S(net920),
    .X(_0247_));
 sg13g2_mux2_1 _6129_ (.A0(\dtop.field_top.acc[16] ),
    .A1(net535),
    .S(net918),
    .X(_0248_));
 sg13g2_or2_2 _6130_ (.X(_2539_),
    .B(_2525_),
    .A(_2523_));
 sg13g2_mux2_1 _6131_ (.A0(\dtop.field_top.acc[0] ),
    .A1(net479),
    .S(net884),
    .X(_0249_));
 sg13g2_nand2_1 _6132_ (.Y(_2540_),
    .A(net356),
    .B(net884));
 sg13g2_o21ai_1 _6133_ (.B1(_2540_),
    .Y(_0250_),
    .A1(_2875_),
    .A2(net884));
 sg13g2_nand2_1 _6134_ (.Y(_2541_),
    .A(net429),
    .B(net884));
 sg13g2_o21ai_1 _6135_ (.B1(_2541_),
    .Y(_0251_),
    .A1(_2878_),
    .A2(net884));
 sg13g2_nor2_1 _6136_ (.A(\dtop.field_top.acc[3] ),
    .B(net883),
    .Y(_2542_));
 sg13g2_a21oi_1 _6137_ (.A1(_2890_),
    .A2(net883),
    .Y(_0252_),
    .B1(_2542_));
 sg13g2_nand2_1 _6138_ (.Y(_2543_),
    .A(net514),
    .B(net883));
 sg13g2_o21ai_1 _6139_ (.B1(_2543_),
    .Y(_0253_),
    .A1(_2877_),
    .A2(net883));
 sg13g2_nor2_1 _6140_ (.A(\dtop.field_top.acc[5] ),
    .B(net883),
    .Y(_2544_));
 sg13g2_a21oi_1 _6141_ (.A1(_2900_),
    .A2(net883),
    .Y(_0254_),
    .B1(_2544_));
 sg13g2_nor2_1 _6142_ (.A(\dtop.field_top.acc[6] ),
    .B(net883),
    .Y(_2545_));
 sg13g2_a21oi_1 _6143_ (.A1(_2905_),
    .A2(net885),
    .Y(_0255_),
    .B1(_2545_));
 sg13g2_nor2_1 _6144_ (.A(\dtop.field_top.acc[7] ),
    .B(_2539_),
    .Y(_2546_));
 sg13g2_a21oi_1 _6145_ (.A1(_2909_),
    .A2(net883),
    .Y(_0256_),
    .B1(_2546_));
 sg13g2_mux2_1 _6146_ (.A0(\dtop.field_top.acc[8] ),
    .A1(net554),
    .S(_2539_),
    .X(_0257_));
 sg13g2_mux2_1 _6147_ (.A0(\dtop.field_top.acc[9] ),
    .A1(net625),
    .S(_2539_),
    .X(_0258_));
 sg13g2_mux2_1 _6148_ (.A0(\dtop.field_top.acc[10] ),
    .A1(net573),
    .S(net885),
    .X(_0259_));
 sg13g2_mux2_1 _6149_ (.A0(\dtop.field_top.acc[11] ),
    .A1(net475),
    .S(net885),
    .X(_0260_));
 sg13g2_mux2_1 _6150_ (.A0(\dtop.field_top.acc[12] ),
    .A1(net443),
    .S(net885),
    .X(_0261_));
 sg13g2_mux2_1 _6151_ (.A0(\dtop.field_top.acc[13] ),
    .A1(net445),
    .S(net884),
    .X(_0262_));
 sg13g2_mux2_1 _6152_ (.A0(\dtop.field_top.acc[14] ),
    .A1(net516),
    .S(net884),
    .X(_0263_));
 sg13g2_nand2_1 _6153_ (.Y(_2547_),
    .A(net337),
    .B(net885));
 sg13g2_o21ai_1 _6154_ (.B1(_2547_),
    .Y(_0264_),
    .A1(_2881_),
    .A2(net885));
 sg13g2_mux2_1 _6155_ (.A0(\dtop.field_top.acc[16] ),
    .A1(net467),
    .S(net884),
    .X(_0265_));
 sg13g2_mux2_1 _6156_ (.A0(_0433_),
    .A1(_2490_),
    .S(net968),
    .X(_2548_));
 sg13g2_or2_2 _6157_ (.X(_2549_),
    .B(_2548_),
    .A(_2496_));
 sg13g2_mux2_1 _6158_ (.A0(\dtop.field_top.acc[0] ),
    .A1(net518),
    .S(net915),
    .X(_0266_));
 sg13g2_nand2_1 _6159_ (.Y(_2550_),
    .A(net489),
    .B(net916));
 sg13g2_o21ai_1 _6160_ (.B1(_2550_),
    .Y(_0267_),
    .A1(_2875_),
    .A2(net916));
 sg13g2_nor2_1 _6161_ (.A(\dtop.field_top.acc[2] ),
    .B(net916),
    .Y(_2551_));
 sg13g2_a21oi_1 _6162_ (.A1(_2885_),
    .A2(net916),
    .Y(_0268_),
    .B1(_2551_));
 sg13g2_nor2_1 _6163_ (.A(\dtop.field_top.acc[3] ),
    .B(net915),
    .Y(_2552_));
 sg13g2_a21oi_1 _6164_ (.A1(_2889_),
    .A2(net915),
    .Y(_0269_),
    .B1(_2552_));
 sg13g2_nand2_1 _6165_ (.Y(_2553_),
    .A(net528),
    .B(net916));
 sg13g2_o21ai_1 _6166_ (.B1(_2553_),
    .Y(_0270_),
    .A1(_2877_),
    .A2(net916));
 sg13g2_nor2_1 _6167_ (.A(\dtop.field_top.acc[5] ),
    .B(net915),
    .Y(_2554_));
 sg13g2_a21oi_1 _6168_ (.A1(_2899_),
    .A2(net915),
    .Y(_0271_),
    .B1(_2554_));
 sg13g2_mux2_1 _6169_ (.A0(\dtop.field_top.acc[6] ),
    .A1(net631),
    .S(net916),
    .X(_0272_));
 sg13g2_mux2_1 _6170_ (.A0(\dtop.field_top.acc[7] ),
    .A1(net611),
    .S(net917),
    .X(_0273_));
 sg13g2_mux2_1 _6171_ (.A0(\dtop.field_top.acc[8] ),
    .A1(net595),
    .S(net917),
    .X(_0274_));
 sg13g2_nor2_1 _6172_ (.A(\dtop.field_top.acc[9] ),
    .B(net917),
    .Y(_2555_));
 sg13g2_a21oi_1 _6173_ (.A1(_2872_),
    .A2(net917),
    .Y(_0275_),
    .B1(_2555_));
 sg13g2_mux2_1 _6174_ (.A0(\dtop.field_top.acc[10] ),
    .A1(net608),
    .S(net917),
    .X(_0276_));
 sg13g2_mux2_1 _6175_ (.A0(\dtop.field_top.acc[11] ),
    .A1(net469),
    .S(net915),
    .X(_0277_));
 sg13g2_mux2_1 _6176_ (.A0(\dtop.field_top.acc[12] ),
    .A1(net465),
    .S(_2549_),
    .X(_0278_));
 sg13g2_mux2_1 _6177_ (.A0(\dtop.field_top.acc[13] ),
    .A1(net447),
    .S(net917),
    .X(_0279_));
 sg13g2_mux2_1 _6178_ (.A0(\dtop.field_top.acc[14] ),
    .A1(net547),
    .S(net915),
    .X(_0280_));
 sg13g2_nand2_1 _6179_ (.Y(_2556_),
    .A(net348),
    .B(_2549_));
 sg13g2_o21ai_1 _6180_ (.B1(_2556_),
    .Y(_0281_),
    .A1(_2881_),
    .A2(net917));
 sg13g2_mux2_1 _6181_ (.A0(\dtop.field_top.acc[16] ),
    .A1(net455),
    .S(net915),
    .X(_0282_));
 sg13g2_nand3_1 _6182_ (.B(_0734_),
    .C(_1020_),
    .A(_0438_),
    .Y(_2557_));
 sg13g2_mux2_1 _6183_ (.A0(_0053_),
    .A1(_2471_),
    .S(_2473_),
    .X(_2558_));
 sg13g2_mux2_1 _6184_ (.A0(_2558_),
    .A1(net560),
    .S(_2557_),
    .X(_0283_));
 sg13g2_nor2_1 _6185_ (.A(_3049_),
    .B(net966),
    .Y(_2559_));
 sg13g2_o21ai_1 _6186_ (.B1(_0734_),
    .Y(_2560_),
    .A1(_2472_),
    .A2(_2559_));
 sg13g2_mux2_1 _6187_ (.A0(_2558_),
    .A1(net584),
    .S(_2560_),
    .X(_0284_));
 sg13g2_and2_1 _6188_ (.A(_0001_),
    .B(_2989_),
    .X(_0287_));
 sg13g2_o21ai_1 _6189_ (.B1(net1117),
    .Y(_2561_),
    .A1(net629),
    .A2(_2946_));
 sg13g2_a21oi_1 _6190_ (.A1(net629),
    .A2(_2967_),
    .Y(_0288_),
    .B1(_2561_));
 sg13g2_nand2b_2 _6191_ (.Y(_2562_),
    .B(_2967_),
    .A_N(_2929_));
 sg13g2_nand2_1 _6192_ (.Y(_2563_),
    .A(net1116),
    .B(_2562_));
 sg13g2_a21oi_1 _6193_ (.A1(_2865_),
    .A2(_2971_),
    .Y(_0289_),
    .B1(net936));
 sg13g2_xnor2_1 _6194_ (.Y(_2564_),
    .A(net693),
    .B(net957));
 sg13g2_nand2_1 _6195_ (.Y(_0290_),
    .A(net935),
    .B(_2564_));
 sg13g2_xnor2_1 _6196_ (.Y(_2565_),
    .A(\dtop.field_top.alt_osc[2] ),
    .B(_1089_));
 sg13g2_nand2_1 _6197_ (.Y(_0291_),
    .A(net935),
    .B(net684));
 sg13g2_nor3_2 _6198_ (.A(_0011_),
    .B(_0010_),
    .C(_2971_),
    .Y(_2566_));
 sg13g2_xnor2_1 _6199_ (.Y(_2567_),
    .A(net676),
    .B(_2566_));
 sg13g2_nand2_1 _6200_ (.Y(_0292_),
    .A(net935),
    .B(net677));
 sg13g2_nand2b_1 _6201_ (.Y(_2568_),
    .B(_2566_),
    .A_N(_0013_));
 sg13g2_a21oi_1 _6202_ (.A1(net591),
    .A2(_2568_),
    .Y(_2569_),
    .B1(net931));
 sg13g2_o21ai_1 _6203_ (.B1(_2569_),
    .Y(_0293_),
    .A1(net591),
    .A2(_2568_));
 sg13g2_nand3_1 _6204_ (.B(\dtop.field_top.alt_osc[3] ),
    .C(_2566_),
    .A(net591),
    .Y(_2570_));
 sg13g2_xnor2_1 _6205_ (.Y(_2571_),
    .A(_2866_),
    .B(_2570_));
 sg13g2_nor2_1 _6206_ (.A(net931),
    .B(_2571_),
    .Y(_0294_));
 sg13g2_o21ai_1 _6207_ (.B1(\dtop.field_top.alt_osc[6] ),
    .Y(_2572_),
    .A1(net619),
    .A2(_2570_));
 sg13g2_or3_1 _6208_ (.A(\dtop.field_top.alt_osc[6] ),
    .B(net619),
    .C(_2570_),
    .X(_2573_));
 sg13g2_nand3_1 _6209_ (.B(net620),
    .C(_2573_),
    .A(net934),
    .Y(_0295_));
 sg13g2_or3_2 _6210_ (.A(_2866_),
    .B(_2867_),
    .C(_2570_),
    .X(_2574_));
 sg13g2_inv_1 _6211_ (.Y(_2575_),
    .A(_2574_));
 sg13g2_xor2_1 _6212_ (.B(_2574_),
    .A(net707),
    .X(_2576_));
 sg13g2_nand2_1 _6213_ (.Y(_0296_),
    .A(net934),
    .B(_2576_));
 sg13g2_o21ai_1 _6214_ (.B1(net1060),
    .Y(_2577_),
    .A1(net666),
    .A2(_2574_));
 sg13g2_or3_1 _6215_ (.A(net666),
    .B(net1060),
    .C(_2574_),
    .X(_2578_));
 sg13g2_nand3_1 _6216_ (.B(net667),
    .C(_2578_),
    .A(net934),
    .Y(_0297_));
 sg13g2_nand3_1 _6217_ (.B(net1060),
    .C(_2575_),
    .A(\dtop.field_top.alt_osc[7] ),
    .Y(_2579_));
 sg13g2_xor2_1 _6218_ (.B(_2579_),
    .A(net672),
    .X(_2580_));
 sg13g2_nor2_1 _6219_ (.A(net931),
    .B(_2580_),
    .Y(_0298_));
 sg13g2_o21ai_1 _6220_ (.B1(net601),
    .Y(_2581_),
    .A1(_0109_),
    .A2(_2579_));
 sg13g2_or3_1 _6221_ (.A(_0109_),
    .B(net601),
    .C(_2579_),
    .X(_2582_));
 sg13g2_nand3_1 _6222_ (.B(_2581_),
    .C(_2582_),
    .A(net934),
    .Y(_0299_));
 sg13g2_a21oi_1 _6223_ (.A1(net1108),
    .A2(_0007_),
    .Y(_2583_),
    .B1(_2076_));
 sg13g2_nand2_1 _6224_ (.Y(_2584_),
    .A(net1009),
    .B(_2583_));
 sg13g2_a21oi_2 _6225_ (.B1(net989),
    .Y(_2585_),
    .A2(_2584_),
    .A1(_2859_));
 sg13g2_nand2b_1 _6226_ (.Y(_2586_),
    .B(_3018_),
    .A_N(_0114_));
 sg13g2_o21ai_1 _6227_ (.B1(net1097),
    .Y(_2587_),
    .A1(_2585_),
    .A2(_2586_));
 sg13g2_nand2_1 _6228_ (.Y(_2588_),
    .A(net1106),
    .B(_0007_));
 sg13g2_mux2_1 _6229_ (.A0(_0007_),
    .A1(_2588_),
    .S(_2389_),
    .X(_2589_));
 sg13g2_nand2_1 _6230_ (.Y(_2590_),
    .A(_0115_),
    .B(_2589_));
 sg13g2_o21ai_1 _6231_ (.B1(_0114_),
    .Y(_2591_),
    .A1(_0115_),
    .A2(_2589_));
 sg13g2_a21oi_2 _6232_ (.B1(_2591_),
    .Y(_2592_),
    .A2(_2590_),
    .A1(_2431_));
 sg13g2_o21ai_1 _6233_ (.B1(net945),
    .Y(_2593_),
    .A1(_1698_),
    .A2(_2592_));
 sg13g2_nor2_1 _6234_ (.A(net1098),
    .B(_2593_),
    .Y(_2594_));
 sg13g2_o21ai_1 _6235_ (.B1(_2594_),
    .Y(_2595_),
    .A1(net1105),
    .A2(_1683_));
 sg13g2_nor3_1 _6236_ (.A(net1108),
    .B(net952),
    .C(_1683_),
    .Y(_2596_));
 sg13g2_or2_1 _6237_ (.X(_2597_),
    .B(_2596_),
    .A(_1980_));
 sg13g2_nand4_1 _6238_ (.B(_1716_),
    .C(_1990_),
    .A(_1705_),
    .Y(_2598_),
    .D(_2597_));
 sg13g2_a21oi_2 _6239_ (.B1(_2598_),
    .Y(_2599_),
    .A2(_2595_),
    .A1(_2587_));
 sg13g2_o21ai_1 _6240_ (.B1(net965),
    .Y(_2600_),
    .A1(net1115),
    .A2(_2996_));
 sg13g2_xor2_1 _6241_ (.B(_2600_),
    .A(_2448_),
    .X(_2601_));
 sg13g2_a21oi_1 _6242_ (.A1(_2455_),
    .A2(_2601_),
    .Y(_2602_),
    .B1(_2454_));
 sg13g2_a221oi_1 _6243_ (.B2(_2455_),
    .C1(_2454_),
    .B1(_2601_),
    .A1(_2090_),
    .Y(_2603_),
    .A2(_2600_));
 sg13g2_nand3b_1 _6244_ (.B(_2459_),
    .C(_2600_),
    .Y(_2604_),
    .A_N(_2458_));
 sg13g2_nand3_1 _6245_ (.B(_1699_),
    .C(_1990_),
    .A(net1096),
    .Y(_2605_));
 sg13g2_nand4_1 _6246_ (.B(_1983_),
    .C(_1990_),
    .A(net1028),
    .Y(_2606_),
    .D(_2016_));
 sg13g2_xnor2_1 _6247_ (.Y(_2607_),
    .A(_2605_),
    .B(_2606_));
 sg13g2_xnor2_1 _6248_ (.Y(_2608_),
    .A(_2604_),
    .B(_2607_));
 sg13g2_xnor2_1 _6249_ (.Y(_2609_),
    .A(_2603_),
    .B(_2608_));
 sg13g2_mux2_1 _6250_ (.A0(net440),
    .A1(_2609_),
    .S(_2599_),
    .X(_0300_));
 sg13g2_and3_1 _6251_ (.X(_0301_),
    .A(net1116),
    .B(net304),
    .C(_2562_));
 sg13g2_a21oi_1 _6252_ (.A1(_0443_),
    .A2(_0449_),
    .Y(_0302_),
    .B1(net936));
 sg13g2_xnor2_1 _6253_ (.Y(_2610_),
    .A(net1007),
    .B(_2941_));
 sg13g2_nor2_1 _6254_ (.A(_2563_),
    .B(_2610_),
    .Y(_0303_));
 sg13g2_nor2_1 _6255_ (.A(net659),
    .B(_2941_),
    .Y(_2611_));
 sg13g2_xnor2_1 _6256_ (.Y(_2612_),
    .A(net1053),
    .B(_2611_));
 sg13g2_nor2_1 _6257_ (.A(net936),
    .B(_2612_),
    .Y(_0304_));
 sg13g2_xnor2_1 _6258_ (.Y(_2613_),
    .A(net1004),
    .B(_2943_));
 sg13g2_nor2_1 _6259_ (.A(net936),
    .B(_2613_),
    .Y(_0305_));
 sg13g2_xnor2_1 _6260_ (.Y(_2614_),
    .A(net1047),
    .B(_2944_));
 sg13g2_nor2_1 _6261_ (.A(net936),
    .B(_2614_),
    .Y(_0306_));
 sg13g2_or2_2 _6262_ (.X(_2615_),
    .B(_3044_),
    .A(_2943_));
 sg13g2_xnor2_1 _6263_ (.Y(_2616_),
    .A(_2846_),
    .B(_2615_));
 sg13g2_nand3_1 _6264_ (.B(_2562_),
    .C(_2616_),
    .A(net1116),
    .Y(_0307_));
 sg13g2_nor2_1 _6265_ (.A(net713),
    .B(_2615_),
    .Y(_2617_));
 sg13g2_xnor2_1 _6266_ (.Y(_2618_),
    .A(net1043),
    .B(_2617_));
 sg13g2_nor2_1 _6267_ (.A(net936),
    .B(_2618_),
    .Y(_0308_));
 sg13g2_nor2_1 _6268_ (.A(_3047_),
    .B(_2615_),
    .Y(_2619_));
 sg13g2_xnor2_1 _6269_ (.Y(_2620_),
    .A(net1040),
    .B(_2619_));
 sg13g2_nor2_1 _6270_ (.A(net936),
    .B(_2620_),
    .Y(_0309_));
 sg13g2_nor3_1 _6271_ (.A(net599),
    .B(_3047_),
    .C(_2615_),
    .Y(_2621_));
 sg13g2_xnor2_1 _6272_ (.Y(_2622_),
    .A(net1038),
    .B(net600));
 sg13g2_nor2_1 _6273_ (.A(net936),
    .B(_2622_),
    .Y(_0310_));
 sg13g2_nand3_1 _6274_ (.B(net1038),
    .C(_2619_),
    .A(net1040),
    .Y(_2623_));
 sg13g2_xnor2_1 _6275_ (.Y(_2624_),
    .A(_2843_),
    .B(_2623_));
 sg13g2_nand3_1 _6276_ (.B(_2562_),
    .C(_2624_),
    .A(net1116),
    .Y(_0311_));
 sg13g2_nand2b_1 _6277_ (.Y(_2625_),
    .B(net358),
    .A_N(net318));
 sg13g2_nor2_1 _6278_ (.A(net346),
    .B(net1001),
    .Y(_2626_));
 sg13g2_a21oi_1 _6279_ (.A1(_1444_),
    .A2(net1001),
    .Y(_0312_),
    .B1(_2626_));
 sg13g2_mux2_1 _6280_ (.A0(net415),
    .A1(_1445_),
    .S(net1001),
    .X(_0313_));
 sg13g2_mux2_1 _6281_ (.A0(net339),
    .A1(_1447_),
    .S(net1001),
    .X(_0314_));
 sg13g2_nor2_1 _6282_ (.A(net325),
    .B(net1001),
    .Y(_2627_));
 sg13g2_a21oi_1 _6283_ (.A1(_1443_),
    .A2(net1001),
    .Y(_0315_),
    .B1(_2627_));
 sg13g2_nor2_1 _6284_ (.A(net320),
    .B(net1002),
    .Y(_2628_));
 sg13g2_a21oi_1 _6285_ (.A1(_1462_),
    .A2(net1001),
    .Y(_0316_),
    .B1(_2628_));
 sg13g2_nor2_1 _6286_ (.A(net359),
    .B(net1002),
    .Y(_2629_));
 sg13g2_a21oi_1 _6287_ (.A1(_1454_),
    .A2(net1001),
    .Y(_0317_),
    .B1(_2629_));
 sg13g2_xnor2_1 _6288_ (.Y(_2630_),
    .A(_1421_),
    .B(_1422_));
 sg13g2_nor2_1 _6289_ (.A(net344),
    .B(net1002),
    .Y(_2631_));
 sg13g2_a21oi_1 _6290_ (.A1(net1002),
    .A2(_2630_),
    .Y(_0318_),
    .B1(_2631_));
 sg13g2_nor2_1 _6291_ (.A(net335),
    .B(net1002),
    .Y(_2632_));
 sg13g2_xnor2_1 _6292_ (.Y(_2633_),
    .A(_1431_),
    .B(_1432_));
 sg13g2_a21oi_1 _6293_ (.A1(net1002),
    .A2(_2633_),
    .Y(_0319_),
    .B1(_2632_));
 sg13g2_mux2_1 _6294_ (.A0(net618),
    .A1(_1015_),
    .S(net912),
    .X(_0320_));
 sg13g2_nor2_1 _6295_ (.A(net643),
    .B(net912),
    .Y(_2634_));
 sg13g2_nand2_1 _6296_ (.Y(_2635_),
    .A(_1012_),
    .B(_1014_));
 sg13g2_xnor2_1 _6297_ (.Y(_2636_),
    .A(net858),
    .B(_2635_));
 sg13g2_a21oi_1 _6298_ (.A1(net912),
    .A2(_2636_),
    .Y(_0321_),
    .B1(_2634_));
 sg13g2_a21oi_1 _6299_ (.A1(_0445_),
    .A2(_0705_),
    .Y(_2637_),
    .B1(_0457_));
 sg13g2_nor2_1 _6300_ (.A(net402),
    .B(_2637_),
    .Y(_2638_));
 sg13g2_or3_1 _6301_ (.A(_0590_),
    .B(_0680_),
    .C(_0689_),
    .X(_2639_));
 sg13g2_o21ai_1 _6302_ (.B1(_0705_),
    .Y(_2640_),
    .A1(_0773_),
    .A2(_2639_));
 sg13g2_a22oi_1 _6303_ (.Y(_2641_),
    .B1(_1015_),
    .B2(_2640_),
    .A2(_0705_),
    .A1(_0678_));
 sg13g2_a21oi_1 _6304_ (.A1(_2637_),
    .A2(_2641_),
    .Y(_0322_),
    .B1(_2638_));
 sg13g2_xor2_1 _6305_ (.B(_0932_),
    .A(_0930_),
    .X(_2642_));
 sg13g2_nor2_2 _6306_ (.A(net878),
    .B(_0677_),
    .Y(_2643_));
 sg13g2_a22oi_1 _6307_ (.Y(_2644_),
    .B1(_2642_),
    .B2(_2643_),
    .A2(net879),
    .A1(net679));
 sg13g2_inv_1 _6308_ (.Y(_0323_),
    .A(net680));
 sg13g2_or2_1 _6309_ (.X(_2645_),
    .B(_0934_),
    .A(_0933_));
 sg13g2_nand3_1 _6310_ (.B(_2643_),
    .C(_2645_),
    .A(_0935_),
    .Y(_2646_));
 sg13g2_o21ai_1 _6311_ (.B1(_2646_),
    .Y(_0324_),
    .A1(_2875_),
    .A2(_0459_));
 sg13g2_nand2_1 _6312_ (.Y(_2647_),
    .A(_0936_),
    .B(_0937_));
 sg13g2_nand3_1 _6313_ (.B(_2643_),
    .C(_2647_),
    .A(_0938_),
    .Y(_2648_));
 sg13g2_o21ai_1 _6314_ (.B1(_2648_),
    .Y(_0325_),
    .A1(_2878_),
    .A2(_0459_));
 sg13g2_nand2_1 _6315_ (.Y(_2649_),
    .A(net681),
    .B(net879));
 sg13g2_nand2b_1 _6316_ (.Y(_2650_),
    .B(_0941_),
    .A_N(_0939_));
 sg13g2_nand2_1 _6317_ (.Y(_2651_),
    .A(_2643_),
    .B(_2650_));
 sg13g2_o21ai_1 _6318_ (.B1(_2649_),
    .Y(_0326_),
    .A1(_0942_),
    .A2(_2651_));
 sg13g2_nand2_1 _6319_ (.Y(_2652_),
    .A(_0943_),
    .B(_0944_));
 sg13g2_nand3_1 _6320_ (.B(_2643_),
    .C(_2652_),
    .A(_0945_),
    .Y(_2653_));
 sg13g2_o21ai_1 _6321_ (.B1(_2653_),
    .Y(_0327_),
    .A1(_2877_),
    .A2(_0459_));
 sg13g2_xnor2_1 _6322_ (.Y(_2654_),
    .A(_0946_),
    .B(_0947_));
 sg13g2_nor3_1 _6323_ (.A(net879),
    .B(_0677_),
    .C(_2654_),
    .Y(_2655_));
 sg13g2_a21oi_1 _6324_ (.A1(net697),
    .A2(net879),
    .Y(_2656_),
    .B1(_2655_));
 sg13g2_inv_1 _6325_ (.Y(_0328_),
    .A(_2656_));
 sg13g2_xnor2_1 _6326_ (.Y(_2657_),
    .A(_0948_),
    .B(_0950_));
 sg13g2_a22oi_1 _6327_ (.Y(_2658_),
    .B1(_2643_),
    .B2(_2657_),
    .A2(net879),
    .A1(net703));
 sg13g2_inv_1 _6328_ (.Y(_0329_),
    .A(_2658_));
 sg13g2_nand2_1 _6329_ (.Y(_2659_),
    .A(net709),
    .B(net878));
 sg13g2_nor2_1 _6330_ (.A(_0951_),
    .B(_0953_),
    .Y(_2660_));
 sg13g2_nand2_1 _6331_ (.Y(_2661_),
    .A(_0954_),
    .B(_2643_));
 sg13g2_o21ai_1 _6332_ (.B1(_2659_),
    .Y(_0330_),
    .A1(_2660_),
    .A2(_2661_));
 sg13g2_nand2_1 _6333_ (.Y(_2662_),
    .A(net434),
    .B(net933));
 sg13g2_o21ai_1 _6334_ (.B1(_2662_),
    .Y(_0331_),
    .A1(_2928_),
    .A2(net933));
 sg13g2_nand2_1 _6335_ (.Y(_2663_),
    .A(net477),
    .B(net934));
 sg13g2_o21ai_1 _6336_ (.B1(_2663_),
    .Y(_0332_),
    .A1(_2927_),
    .A2(net933));
 sg13g2_nand2_1 _6337_ (.Y(_2664_),
    .A(net471),
    .B(net933));
 sg13g2_o21ai_1 _6338_ (.B1(_2664_),
    .Y(_0333_),
    .A1(_2926_),
    .A2(net934));
 sg13g2_mux2_1 _6339_ (.A0(net649),
    .A1(\dtop.field_top.controller.ppos[0] ),
    .S(net934),
    .X(_0334_));
 sg13g2_mux2_1 _6340_ (.A0(\dtop.field_top.player.controller.ppos[1] ),
    .A1(net644),
    .S(net932),
    .X(_0335_));
 sg13g2_nand2_1 _6341_ (.Y(_2665_),
    .A(net627),
    .B(net932));
 sg13g2_o21ai_1 _6342_ (.B1(_2665_),
    .Y(_0336_),
    .A1(_2855_),
    .A2(net932));
 sg13g2_mux2_1 _6343_ (.A0(net678),
    .A1(net1077),
    .S(net929),
    .X(_0337_));
 sg13g2_nor2_1 _6344_ (.A(net653),
    .B(net928),
    .Y(_2666_));
 sg13g2_a21oi_1 _6345_ (.A1(net1012),
    .A2(net928),
    .Y(_0338_),
    .B1(_2666_));
 sg13g2_mux2_1 _6346_ (.A0(net1033),
    .A1(net1065),
    .S(net929),
    .X(_0339_));
 sg13g2_nor2_1 _6347_ (.A(net1032),
    .B(net928),
    .Y(_2667_));
 sg13g2_a21oi_1 _6348_ (.A1(_2854_),
    .A2(net929),
    .Y(_0340_),
    .B1(_2667_));
 sg13g2_nor2_1 _6349_ (.A(\dtop.field_top.controller.pattern0[0] ),
    .B(net930),
    .Y(_2668_));
 sg13g2_a21oi_1 _6350_ (.A1(_2925_),
    .A2(net930),
    .Y(_0341_),
    .B1(_2668_));
 sg13g2_nand2_1 _6351_ (.Y(_2669_),
    .A(net423),
    .B(net930));
 sg13g2_o21ai_1 _6352_ (.B1(_2669_),
    .Y(_0342_),
    .A1(_2850_),
    .A2(net930));
 sg13g2_nor2_1 _6353_ (.A(net1030),
    .B(net930),
    .Y(_2670_));
 sg13g2_a21oi_1 _6354_ (.A1(_2851_),
    .A2(net931),
    .Y(_0343_),
    .B1(_2670_));
 sg13g2_or2_2 _6355_ (.X(_2671_),
    .B(_2602_),
    .A(net868));
 sg13g2_a21oi_1 _6356_ (.A1(net425),
    .A2(_2671_),
    .Y(_2672_),
    .B1(net1110));
 sg13g2_o21ai_1 _6357_ (.B1(_2672_),
    .Y(_0344_),
    .A1(net425),
    .A2(_2671_));
 sg13g2_nor2_1 _6358_ (.A(_2975_),
    .B(_2989_),
    .Y(_0345_));
 sg13g2_nand2_1 _6359_ (.Y(_0346_),
    .A(_2975_),
    .B(_2988_));
 sg13g2_o21ai_1 _6360_ (.B1(_2002_),
    .Y(_2673_),
    .A1(net989),
    .A2(_2003_));
 sg13g2_nor4_1 _6361_ (.A(_0111_),
    .B(_0112_),
    .C(_3008_),
    .D(net989),
    .Y(_2674_));
 sg13g2_nand2b_1 _6362_ (.Y(_2675_),
    .B(_1679_),
    .A_N(_2674_));
 sg13g2_and4_1 _6363_ (.A(_1716_),
    .B(_2600_),
    .C(_2673_),
    .D(_2675_),
    .X(_2676_));
 sg13g2_o21ai_1 _6364_ (.B1(net1119),
    .Y(_2677_),
    .A1(net580),
    .A2(net864));
 sg13g2_a21oi_1 _6365_ (.A1(_2159_),
    .A2(net864),
    .Y(_0347_),
    .B1(_2677_));
 sg13g2_o21ai_1 _6366_ (.B1(net1118),
    .Y(_2678_),
    .A1(net603),
    .A2(net862));
 sg13g2_a21oi_1 _6367_ (.A1(_2183_),
    .A2(net862),
    .Y(_0348_),
    .B1(_2678_));
 sg13g2_nor2b_1 _6368_ (.A(_2205_),
    .B_N(net863),
    .Y(_2679_));
 sg13g2_o21ai_1 _6369_ (.B1(net1118),
    .Y(_2680_),
    .A1(net582),
    .A2(net862));
 sg13g2_nor2_1 _6370_ (.A(_2679_),
    .B(_2680_),
    .Y(_0349_));
 sg13g2_o21ai_1 _6371_ (.B1(net1118),
    .Y(_2681_),
    .A1(net522),
    .A2(net862));
 sg13g2_a21oi_1 _6372_ (.A1(_2230_),
    .A2(net862),
    .Y(_0350_),
    .B1(_2681_));
 sg13g2_nor2b_1 _6373_ (.A(_2250_),
    .B_N(net863),
    .Y(_2682_));
 sg13g2_o21ai_1 _6374_ (.B1(net1118),
    .Y(_2683_),
    .A1(net564),
    .A2(net864));
 sg13g2_nor2_1 _6375_ (.A(_2682_),
    .B(_2683_),
    .Y(_0351_));
 sg13g2_o21ai_1 _6376_ (.B1(net1118),
    .Y(_2684_),
    .A1(net549),
    .A2(net862));
 sg13g2_a21oi_1 _6377_ (.A1(_2273_),
    .A2(net862),
    .Y(_0352_),
    .B1(_2684_));
 sg13g2_o21ai_1 _6378_ (.B1(net1119),
    .Y(_2685_),
    .A1(net610),
    .A2(net862));
 sg13g2_a21oi_1 _6379_ (.A1(_2299_),
    .A2(net863),
    .Y(_0353_),
    .B1(_2685_));
 sg13g2_o21ai_1 _6380_ (.B1(net1119),
    .Y(_2686_),
    .A1(net575),
    .A2(net864));
 sg13g2_a21oi_1 _6381_ (.A1(_2353_),
    .A2(net863),
    .Y(_0354_),
    .B1(_2686_));
 sg13g2_o21ai_1 _6382_ (.B1(net1118),
    .Y(_2687_),
    .A1(net520),
    .A2(net865));
 sg13g2_a21oi_1 _6383_ (.A1(_2404_),
    .A2(net865),
    .Y(_0355_),
    .B1(_2687_));
 sg13g2_o21ai_1 _6384_ (.B1(net1118),
    .Y(_2688_),
    .A1(net526),
    .A2(net865));
 sg13g2_a21oi_1 _6385_ (.A1(_2446_),
    .A2(net865),
    .Y(_0356_),
    .B1(_2688_));
 sg13g2_a21o_1 _6386_ (.A2(_1694_),
    .A1(net1117),
    .B1(_1717_),
    .X(_2689_));
 sg13g2_nand3_1 _6387_ (.B(_1716_),
    .C(_2689_),
    .A(net965),
    .Y(_2690_));
 sg13g2_inv_2 _6388_ (.Y(_2691_),
    .A(net860));
 sg13g2_a21oi_1 _6389_ (.A1(net572),
    .A2(net860),
    .Y(_2692_),
    .B1(net1112));
 sg13g2_o21ai_1 _6390_ (.B1(_2692_),
    .Y(_0357_),
    .A1(_2159_),
    .A2(net860));
 sg13g2_a21oi_1 _6391_ (.A1(net579),
    .A2(net861),
    .Y(_2693_),
    .B1(net1112));
 sg13g2_o21ai_1 _6392_ (.B1(_2693_),
    .Y(_0358_),
    .A1(_2183_),
    .A2(net861));
 sg13g2_a21oi_1 _6393_ (.A1(_2205_),
    .A2(_2691_),
    .Y(_2694_),
    .B1(net1112));
 sg13g2_o21ai_1 _6394_ (.B1(_2694_),
    .Y(_0359_),
    .A1(_2826_),
    .A2(_2691_));
 sg13g2_a21oi_1 _6395_ (.A1(net431),
    .A2(net859),
    .Y(_2695_),
    .B1(net1110));
 sg13g2_o21ai_1 _6396_ (.B1(_2695_),
    .Y(_0360_),
    .A1(_2230_),
    .A2(net859));
 sg13g2_a21oi_1 _6397_ (.A1(_2250_),
    .A2(_2691_),
    .Y(_2696_),
    .B1(net1113));
 sg13g2_o21ai_1 _6398_ (.B1(_2696_),
    .Y(_0361_),
    .A1(_2825_),
    .A2(_2691_));
 sg13g2_a21oi_1 _6399_ (.A1(net483),
    .A2(net860),
    .Y(_2697_),
    .B1(net1112));
 sg13g2_o21ai_1 _6400_ (.B1(_2697_),
    .Y(_0362_),
    .A1(_2273_),
    .A2(net860));
 sg13g2_a21oi_1 _6401_ (.A1(net566),
    .A2(net860),
    .Y(_2698_),
    .B1(net1113));
 sg13g2_o21ai_1 _6402_ (.B1(_2698_),
    .Y(_0363_),
    .A1(_2299_),
    .A2(net860));
 sg13g2_a21oi_1 _6403_ (.A1(net482),
    .A2(net860),
    .Y(_2699_),
    .B1(net1112));
 sg13g2_o21ai_1 _6404_ (.B1(_2699_),
    .Y(_0364_),
    .A1(_2353_),
    .A2(net861));
 sg13g2_a21oi_1 _6405_ (.A1(net488),
    .A2(net859),
    .Y(_2700_),
    .B1(net1112));
 sg13g2_o21ai_1 _6406_ (.B1(_2700_),
    .Y(_0365_),
    .A1(_2404_),
    .A2(net859));
 sg13g2_a21oi_1 _6407_ (.A1(net510),
    .A2(net859),
    .Y(_2701_),
    .B1(net1112));
 sg13g2_o21ai_1 _6408_ (.B1(_2701_),
    .Y(_0366_),
    .A1(_2446_),
    .A2(net859));
 sg13g2_a21oi_1 _6409_ (.A1(net621),
    .A2(net859),
    .Y(_2702_),
    .B1(net1111));
 sg13g2_o21ai_1 _6410_ (.B1(_2702_),
    .Y(_0367_),
    .A1(_2460_),
    .A2(net859));
 sg13g2_a221oi_1 _6411_ (.B2(_1714_),
    .C1(_2014_),
    .B1(_1679_),
    .A1(_3003_),
    .Y(_2703_),
    .A2(_1676_));
 sg13g2_nor2b_1 _6412_ (.A(net580),
    .B_N(net870),
    .Y(_2704_));
 sg13g2_and2_1 _6413_ (.A(\dtop.field_top.player.out_pw[0] ),
    .B(_2980_),
    .X(_2705_));
 sg13g2_nor2b_1 _6414_ (.A(net871),
    .B_N(_2705_),
    .Y(_2706_));
 sg13g2_nor3_1 _6415_ (.A(net1115),
    .B(_2704_),
    .C(_2706_),
    .Y(_0368_));
 sg13g2_xor2_1 _6416_ (.B(_2705_),
    .A(\dtop.field_top.player.out_pw[1] ),
    .X(_2707_));
 sg13g2_nor2_1 _6417_ (.A(net871),
    .B(_2707_),
    .Y(_2708_));
 sg13g2_nor2b_1 _6418_ (.A(net603),
    .B_N(net870),
    .Y(_2709_));
 sg13g2_nor3_1 _6419_ (.A(net1115),
    .B(_2708_),
    .C(_2709_),
    .Y(_0369_));
 sg13g2_and3_1 _6420_ (.X(_2710_),
    .A(\dtop.field_top.player.out_pw[1] ),
    .B(\dtop.field_top.player.out_pw[2] ),
    .C(_2705_));
 sg13g2_a21oi_1 _6421_ (.A1(\dtop.field_top.player.out_pw[1] ),
    .A2(net384),
    .Y(_2711_),
    .B1(\dtop.field_top.player.out_pw[2] ));
 sg13g2_nor2_1 _6422_ (.A(_2710_),
    .B(_2711_),
    .Y(_2712_));
 sg13g2_nor2_1 _6423_ (.A(net871),
    .B(_2712_),
    .Y(_2713_));
 sg13g2_nor2b_1 _6424_ (.A(net582),
    .B_N(net870),
    .Y(_2714_));
 sg13g2_nor3_1 _6425_ (.A(net1114),
    .B(_2713_),
    .C(_2714_),
    .Y(_0370_));
 sg13g2_xor2_1 _6426_ (.B(_2710_),
    .A(\dtop.field_top.player.out_pw[3] ),
    .X(_2715_));
 sg13g2_nor2_1 _6427_ (.A(net871),
    .B(_2715_),
    .Y(_2716_));
 sg13g2_nor2b_1 _6428_ (.A(net522),
    .B_N(net870),
    .Y(_2717_));
 sg13g2_nor3_1 _6429_ (.A(net1114),
    .B(_2716_),
    .C(_2717_),
    .Y(_0371_));
 sg13g2_nand3_1 _6430_ (.B(\dtop.field_top.player.out_pw[4] ),
    .C(_2710_),
    .A(\dtop.field_top.player.out_pw[3] ),
    .Y(_2718_));
 sg13g2_a21o_1 _6431_ (.A2(_2710_),
    .A1(\dtop.field_top.player.out_pw[3] ),
    .B1(\dtop.field_top.player.out_pw[4] ),
    .X(_2719_));
 sg13g2_a21oi_1 _6432_ (.A1(_2718_),
    .A2(_2719_),
    .Y(_2720_),
    .B1(net870));
 sg13g2_nor2b_1 _6433_ (.A(net564),
    .B_N(net870),
    .Y(_2721_));
 sg13g2_nor3_1 _6434_ (.A(net1114),
    .B(_2720_),
    .C(_2721_),
    .Y(_0372_));
 sg13g2_nor2_1 _6435_ (.A(_2912_),
    .B(_2718_),
    .Y(_2722_));
 sg13g2_xnor2_1 _6436_ (.Y(_2723_),
    .A(\dtop.field_top.player.out_pw[5] ),
    .B(_2718_));
 sg13g2_nor2_1 _6437_ (.A(net871),
    .B(_2723_),
    .Y(_2724_));
 sg13g2_nor2b_1 _6438_ (.A(net549),
    .B_N(net870),
    .Y(_2725_));
 sg13g2_nor3_1 _6439_ (.A(net1114),
    .B(_2724_),
    .C(_2725_),
    .Y(_0373_));
 sg13g2_and2_1 _6440_ (.A(\dtop.field_top.player.out_pw[6] ),
    .B(_2722_),
    .X(_2726_));
 sg13g2_xnor2_1 _6441_ (.Y(_2727_),
    .A(net628),
    .B(_2722_));
 sg13g2_mux2_1 _6442_ (.A0(_2727_),
    .A1(_2829_),
    .S(net870),
    .X(_2728_));
 sg13g2_nor2_1 _6443_ (.A(net1114),
    .B(_2728_),
    .Y(_0374_));
 sg13g2_xor2_1 _6444_ (.B(_2726_),
    .A(\dtop.field_top.player.out_pw[7] ),
    .X(_2729_));
 sg13g2_o21ai_1 _6445_ (.B1(net1119),
    .Y(_2730_),
    .A1(net872),
    .A2(_2729_));
 sg13g2_a21oi_1 _6446_ (.A1(_2828_),
    .A2(net872),
    .Y(_0375_),
    .B1(_2730_));
 sg13g2_a21o_1 _6447_ (.A2(_2726_),
    .A1(\dtop.field_top.player.out_pw[7] ),
    .B1(\dtop.field_top.player.out_pw[8] ),
    .X(_2731_));
 sg13g2_nand2b_1 _6448_ (.Y(_2732_),
    .B(_2726_),
    .A_N(_2976_));
 sg13g2_a21oi_1 _6449_ (.A1(_2731_),
    .A2(_2732_),
    .Y(_2733_),
    .B1(net872));
 sg13g2_nor2b_1 _6450_ (.A(net520),
    .B_N(net872),
    .Y(_2734_));
 sg13g2_nor3_1 _6451_ (.A(net1114),
    .B(_2733_),
    .C(_2734_),
    .Y(_0376_));
 sg13g2_xnor2_1 _6452_ (.Y(_2735_),
    .A(\dtop.field_top.player.out_pw[9] ),
    .B(_2732_));
 sg13g2_o21ai_1 _6453_ (.B1(net1119),
    .Y(_2736_),
    .A1(net872),
    .A2(_2735_));
 sg13g2_a21oi_1 _6454_ (.A1(_2827_),
    .A2(net872),
    .Y(_0377_),
    .B1(_2736_));
 sg13g2_nand2_1 _6455_ (.Y(_2737_),
    .A(net1027),
    .B(_2587_));
 sg13g2_a22oi_1 _6456_ (.Y(_2738_),
    .B1(net945),
    .B2(_1696_),
    .A2(_3018_),
    .A1(net1101));
 sg13g2_nand3_1 _6457_ (.B(_2033_),
    .C(_2738_),
    .A(net1027),
    .Y(_2739_));
 sg13g2_a21oi_1 _6458_ (.A1(_2737_),
    .A2(_2739_),
    .Y(_2740_),
    .B1(_2594_));
 sg13g2_nand3b_1 _6459_ (.B(_2839_),
    .C(_0117_),
    .Y(_2741_),
    .A_N(_1869_));
 sg13g2_nor2_1 _6460_ (.A(_0007_),
    .B(_1880_),
    .Y(_2742_));
 sg13g2_xnor2_1 _6461_ (.Y(_2743_),
    .A(net1106),
    .B(_1880_));
 sg13g2_a221oi_1 _6462_ (.B2(_2743_),
    .C1(_2742_),
    .B1(_2741_),
    .A1(net1104),
    .Y(_2744_),
    .A2(_1883_));
 sg13g2_nor2_1 _6463_ (.A(net1104),
    .B(_1883_),
    .Y(_2745_));
 sg13g2_nor4_1 _6464_ (.A(_3022_),
    .B(net980),
    .C(_2744_),
    .D(_2745_),
    .Y(_2746_));
 sg13g2_nor3_1 _6465_ (.A(_2996_),
    .B(_3001_),
    .C(net981),
    .Y(_2747_));
 sg13g2_nor3_1 _6466_ (.A(net951),
    .B(_2746_),
    .C(_2747_),
    .Y(_2748_));
 sg13g2_nor3_1 _6467_ (.A(net1097),
    .B(net945),
    .C(_1707_),
    .Y(_2749_));
 sg13g2_nor3_1 _6468_ (.A(net1027),
    .B(_2748_),
    .C(_2749_),
    .Y(_2750_));
 sg13g2_o21ai_1 _6469_ (.B1(net941),
    .Y(_2751_),
    .A1(_2740_),
    .A2(_2750_));
 sg13g2_nor2b_1 _6470_ (.A(_2585_),
    .B_N(_2009_),
    .Y(_2752_));
 sg13g2_and3_1 _6471_ (.X(_2753_),
    .A(_2011_),
    .B(_2040_),
    .C(_2058_));
 sg13g2_nor3_1 _6472_ (.A(net965),
    .B(_2752_),
    .C(_2753_),
    .Y(_2754_));
 sg13g2_o21ai_1 _6473_ (.B1(_2751_),
    .Y(_2755_),
    .A1(_1679_),
    .A2(_2754_));
 sg13g2_nand2b_2 _6474_ (.Y(_2756_),
    .B(_1716_),
    .A_N(_2755_));
 sg13g2_and3_1 _6475_ (.X(_2757_),
    .A(_2995_),
    .B(_3001_),
    .C(net980));
 sg13g2_a22oi_1 _6476_ (.Y(_2758_),
    .B1(_2757_),
    .B2(net944),
    .A2(_2021_),
    .A1(net1107));
 sg13g2_nor3_1 _6477_ (.A(net1025),
    .B(net937),
    .C(_2758_),
    .Y(_2759_));
 sg13g2_nor2_1 _6478_ (.A(_3016_),
    .B(_1683_),
    .Y(_2760_));
 sg13g2_a22oi_1 _6479_ (.Y(_2761_),
    .B1(_2760_),
    .B2(_1998_),
    .A2(_2032_),
    .A1(_3000_));
 sg13g2_nand3_1 _6480_ (.B(_2012_),
    .C(_2761_),
    .A(_1677_),
    .Y(_2762_));
 sg13g2_o21ai_1 _6481_ (.B1(_2038_),
    .Y(_2763_),
    .A1(_1514_),
    .A2(_2037_));
 sg13g2_nor3_1 _6482_ (.A(net942),
    .B(_2762_),
    .C(_2763_),
    .Y(_2764_));
 sg13g2_or2_1 _6483_ (.X(_2765_),
    .B(_2764_),
    .A(_2759_));
 sg13g2_nor2_1 _6484_ (.A(_0117_),
    .B(_1999_),
    .Y(_2766_));
 sg13g2_o21ai_1 _6485_ (.B1(net1010),
    .Y(_2767_),
    .A1(net944),
    .A2(_2766_));
 sg13g2_nand3_1 _6486_ (.B(net980),
    .C(_1726_),
    .A(net1104),
    .Y(_2768_));
 sg13g2_a21o_1 _6487_ (.A2(_2768_),
    .A1(net944),
    .B1(_2767_),
    .X(_2769_));
 sg13g2_a21oi_2 _6488_ (.B1(_2070_),
    .Y(_2770_),
    .A2(_2769_),
    .A1(net941));
 sg13g2_nand2_1 _6489_ (.Y(_2771_),
    .A(_1680_),
    .B(_2762_));
 sg13g2_a21oi_1 _6490_ (.A1(net1096),
    .A2(_1726_),
    .Y(_2772_),
    .B1(net951));
 sg13g2_o21ai_1 _6491_ (.B1(net941),
    .Y(_2773_),
    .A1(_2767_),
    .A2(_2772_));
 sg13g2_nand2_1 _6492_ (.Y(_2774_),
    .A(_2771_),
    .B(_2773_));
 sg13g2_inv_1 _6493_ (.Y(_2775_),
    .A(_2774_));
 sg13g2_a21oi_1 _6494_ (.A1(net1099),
    .A2(_1726_),
    .Y(_2776_),
    .B1(net951));
 sg13g2_nor3_2 _6495_ (.A(_1680_),
    .B(_2767_),
    .C(_2776_),
    .Y(_2777_));
 sg13g2_nand2_1 _6496_ (.Y(_2778_),
    .A(_2770_),
    .B(_2777_));
 sg13g2_nand2b_1 _6497_ (.Y(_2779_),
    .B(_2765_),
    .A_N(_2778_));
 sg13g2_nor2_1 _6498_ (.A(_2774_),
    .B(_2779_),
    .Y(_2780_));
 sg13g2_nor2_2 _6499_ (.A(_2756_),
    .B(_2775_),
    .Y(_2781_));
 sg13g2_inv_1 _6500_ (.Y(_2782_),
    .A(_2781_));
 sg13g2_nor2_1 _6501_ (.A(_2756_),
    .B(_2780_),
    .Y(_2783_));
 sg13g2_o21ai_1 _6502_ (.B1(net1118),
    .Y(_2784_),
    .A1(net637),
    .A2(_2783_));
 sg13g2_a21oi_1 _6503_ (.A1(_2159_),
    .A2(_2783_),
    .Y(_0378_),
    .B1(_2784_));
 sg13g2_a21o_2 _6504_ (.A2(_2777_),
    .A1(_2775_),
    .B1(_2756_),
    .X(_2785_));
 sg13g2_o21ai_1 _6505_ (.B1(_2785_),
    .Y(_2786_),
    .A1(_2756_),
    .A2(_2770_));
 sg13g2_o21ai_1 _6506_ (.B1(net1121),
    .Y(_2787_),
    .A1(net656),
    .A2(_2786_));
 sg13g2_a21oi_1 _6507_ (.A1(_2183_),
    .A2(_2786_),
    .Y(_0379_),
    .B1(_2787_));
 sg13g2_a21o_1 _6508_ (.A2(_2771_),
    .A1(_2770_),
    .B1(_2765_),
    .X(_2788_));
 sg13g2_o21ai_1 _6509_ (.B1(_2785_),
    .Y(_2789_),
    .A1(_2756_),
    .A2(_2788_));
 sg13g2_nor2b_1 _6510_ (.A(_2205_),
    .B_N(_2789_),
    .Y(_2790_));
 sg13g2_o21ai_1 _6511_ (.B1(net1121),
    .Y(_2791_),
    .A1(net661),
    .A2(_2789_));
 sg13g2_nor2_1 _6512_ (.A(_2790_),
    .B(_2791_),
    .Y(_0380_));
 sg13g2_o21ai_1 _6513_ (.B1(net1121),
    .Y(_2792_),
    .A1(_2231_),
    .A2(_2785_));
 sg13g2_a21oi_1 _6514_ (.A1(_2821_),
    .A2(_2785_),
    .Y(_0381_),
    .B1(_2792_));
 sg13g2_a21oi_2 _6515_ (.B1(_2785_),
    .Y(_2793_),
    .A2(_2775_),
    .A1(_2770_));
 sg13g2_inv_1 _6516_ (.Y(_2794_),
    .A(_2793_));
 sg13g2_o21ai_1 _6517_ (.B1(_2794_),
    .Y(_2795_),
    .A1(_2765_),
    .A2(_2785_));
 sg13g2_nor2b_1 _6518_ (.A(_2250_),
    .B_N(_2795_),
    .Y(_2796_));
 sg13g2_o21ai_1 _6519_ (.B1(net1121),
    .Y(_2797_),
    .A1(net704),
    .A2(_2795_));
 sg13g2_nor2_1 _6520_ (.A(_2796_),
    .B(_2797_),
    .Y(_0382_));
 sg13g2_o21ai_1 _6521_ (.B1(net1121),
    .Y(_2798_),
    .A1(net706),
    .A2(_2793_));
 sg13g2_a21oi_1 _6522_ (.A1(_2273_),
    .A2(_2793_),
    .Y(_0383_),
    .B1(_2798_));
 sg13g2_a21oi_1 _6523_ (.A1(_2775_),
    .A2(_2788_),
    .Y(_2799_),
    .B1(_2785_));
 sg13g2_o21ai_1 _6524_ (.B1(net1121),
    .Y(_2800_),
    .A1(net694),
    .A2(_2799_));
 sg13g2_a21oi_1 _6525_ (.A1(_2299_),
    .A2(_2799_),
    .Y(_0384_),
    .B1(_2800_));
 sg13g2_o21ai_1 _6526_ (.B1(net1121),
    .Y(_2801_),
    .A1(net586),
    .A2(_2781_));
 sg13g2_a21oi_1 _6527_ (.A1(_2353_),
    .A2(_2781_),
    .Y(_0385_),
    .B1(_2801_));
 sg13g2_and3_1 _6528_ (.X(_2802_),
    .A(_2404_),
    .B(_2779_),
    .C(_2781_));
 sg13g2_a21oi_1 _6529_ (.A1(_2779_),
    .A2(_2781_),
    .Y(_2803_),
    .B1(net664));
 sg13g2_nor3_1 _6530_ (.A(net1114),
    .B(_2802_),
    .C(_2803_),
    .Y(_0386_));
 sg13g2_and3_1 _6531_ (.X(_2804_),
    .A(_2446_),
    .B(_2778_),
    .C(_2781_));
 sg13g2_a21oi_1 _6532_ (.A1(_2778_),
    .A2(_2781_),
    .Y(_2805_),
    .B1(net652));
 sg13g2_nor3_1 _6533_ (.A(net1114),
    .B(_2804_),
    .C(_2805_),
    .Y(_0387_));
 sg13g2_a21oi_1 _6534_ (.A1(_2777_),
    .A2(_2788_),
    .Y(_2806_),
    .B1(_2782_));
 sg13g2_o21ai_1 _6535_ (.B1(net1120),
    .Y(_2807_),
    .A1(net1028),
    .A2(_2806_));
 sg13g2_a21oi_1 _6536_ (.A1(_2460_),
    .A2(_2806_),
    .Y(_0388_),
    .B1(_2807_));
 sg13g2_or2_1 _6537_ (.X(_2808_),
    .B(_2755_),
    .A(_1729_));
 sg13g2_nand4_1 _6538_ (.B(_0117_),
    .C(net944),
    .A(_0111_),
    .Y(_2809_),
    .D(_1725_));
 sg13g2_o21ai_1 _6539_ (.B1(_2808_),
    .Y(_2810_),
    .A1(net937),
    .A2(_2809_));
 sg13g2_a21oi_1 _6540_ (.A1(_1716_),
    .A2(_2810_),
    .Y(_2811_),
    .B1(_2691_));
 sg13g2_nand2_1 _6541_ (.Y(_2812_),
    .A(net317),
    .B(_2811_));
 sg13g2_nor2b_1 _6542_ (.A(_2808_),
    .B_N(_1963_),
    .Y(_2813_));
 sg13g2_a21oi_1 _6543_ (.A1(_2609_),
    .A2(_2808_),
    .Y(_2814_),
    .B1(_2813_));
 sg13g2_o21ai_1 _6544_ (.B1(_2812_),
    .Y(_0389_),
    .A1(_2811_),
    .A2(_2814_));
 sg13g2_nor3_1 _6545_ (.A(net318),
    .B(\dtop.field_top.nsource.num_iter[1] ),
    .C(net1003),
    .Y(_0390_));
 sg13g2_o21ai_1 _6546_ (.B1(_1411_),
    .Y(_2815_),
    .A1(net318),
    .A2(net358));
 sg13g2_a21oi_1 _6547_ (.A1(net318),
    .A2(net358),
    .Y(_0391_),
    .B1(_2815_));
 sg13g2_nor3_1 _6548_ (.A(_0112_),
    .B(_2999_),
    .C(_3017_),
    .Y(_2816_));
 sg13g2_xnor2_1 _6549_ (.Y(_2817_),
    .A(net1025),
    .B(_2816_));
 sg13g2_a21oi_1 _6550_ (.A1(_3004_),
    .A2(_2817_),
    .Y(_0392_),
    .B1(net1115));
 sg13g2_xor2_1 _6551_ (.B(_3009_),
    .A(net633),
    .X(_2818_));
 sg13g2_nand2_1 _6552_ (.Y(_0393_),
    .A(net1117),
    .B(_2818_));
 sg13g2_nor3_1 _6553_ (.A(net710),
    .B(_3009_),
    .C(_3011_),
    .Y(_2819_));
 sg13g2_xor2_1 _6554_ (.B(_2819_),
    .A(\dtop.field_top.channel[3] ),
    .X(_2820_));
 sg13g2_a21o_1 _6555_ (.A2(_2820_),
    .A1(_3004_),
    .B1(net1115),
    .X(_0394_));
 sg13g2_dfrbp_1 _6556_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net88),
    .D(_0118_),
    .Q_N(_3269_),
    .Q(\dtop.field_top.rs.scan_y.state[0] ));
 sg13g2_dfrbp_1 _6557_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net285),
    .D(net641),
    .Q_N(_3268_),
    .Q(\dtop.field_top.rs.scan_y.state[1] ));
 sg13g2_dfrbp_1 _6558_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net284),
    .D(_0120_),
    .Q_N(_3267_),
    .Q(\dtop.field_top.channel[1] ));
 sg13g2_dfrbp_1 _6559_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net283),
    .D(_0121_),
    .Q_N(_0110_),
    .Q(\dtop.field_top.channel[2] ));
 sg13g2_dfrbp_1 _6560_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net282),
    .D(_0122_),
    .Q_N(_0117_),
    .Q(\dtop.field_top.player.chan_timer[0] ));
 sg13g2_dfrbp_1 _6561_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net281),
    .D(_0123_),
    .Q_N(_0007_),
    .Q(\dtop.field_top.player.chan_timer[1] ));
 sg13g2_dfrbp_1 _6562_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net280),
    .D(_0124_),
    .Q_N(_0115_),
    .Q(\dtop.field_top.player.chan_timer[2] ));
 sg13g2_dfrbp_1 _6563_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net279),
    .D(_0125_),
    .Q_N(_0114_),
    .Q(\dtop.field_top.player.chan_timer[3] ));
 sg13g2_dfrbp_1 _6564_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net278),
    .D(_0126_),
    .Q_N(_0112_),
    .Q(\dtop.field_top.player.chan_timer[4] ));
 sg13g2_dfrbp_1 _6565_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net277),
    .D(_0127_),
    .Q_N(_0046_),
    .Q(\dtop.field_top.acc[11] ));
 sg13g2_dfrbp_1 _6566_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net275),
    .D(_0128_),
    .Q_N(_0044_),
    .Q(\dtop.field_top.acc[12] ));
 sg13g2_dfrbp_1 _6567_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net273),
    .D(_0129_),
    .Q_N(_0042_),
    .Q(\dtop.field_top.acc[13] ));
 sg13g2_dfrbp_1 _6568_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net271),
    .D(_0130_),
    .Q_N(_0040_),
    .Q(\dtop.field_top.acc[14] ));
 sg13g2_dfrbp_1 _6569_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net269),
    .D(_0131_),
    .Q_N(_0038_),
    .Q(\dtop.field_top.acc[15] ));
 sg13g2_dfrbp_1 _6570_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net267),
    .D(_0132_),
    .Q_N(_0032_),
    .Q(\dtop.field_top.acc[8] ));
 sg13g2_dfrbp_1 _6571_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net266),
    .D(_0133_),
    .Q_N(_0027_),
    .Q(\dtop.field_top.acc[9] ));
 sg13g2_dfrbp_1 _6572_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net265),
    .D(_0134_),
    .Q_N(_0031_),
    .Q(\dtop.field_top.acc[10] ));
 sg13g2_dfrbp_1 _6573_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net264),
    .D(_0135_),
    .Q_N(_0053_),
    .Q(\dtop.field_top.acc[16] ));
 sg13g2_dfrbp_1 _6574_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net263),
    .D(net452),
    .Q_N(_0024_),
    .Q(\dtop.field_top.fy[9] ));
 sg13g2_dfrbp_1 _6575_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net261),
    .D(net399),
    .Q_N(_3266_),
    .Q(\dtop.field_top.fy[10] ));
 sg13g2_dfrbp_1 _6576_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net259),
    .D(_0138_),
    .Q_N(_0065_),
    .Q(\dtop.field_top.fy[0] ));
 sg13g2_dfrbp_1 _6577_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net258),
    .D(_0139_),
    .Q_N(_0071_),
    .Q(\dtop.field_top.fy[1] ));
 sg13g2_dfrbp_1 _6578_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net257),
    .D(net324),
    .Q_N(_0073_),
    .Q(\dtop.field_top.fy[2] ));
 sg13g2_dfrbp_1 _6579_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net256),
    .D(_0141_),
    .Q_N(_0026_),
    .Q(\dtop.field_top.fy[3] ));
 sg13g2_dfrbp_1 _6580_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net255),
    .D(net364),
    .Q_N(_0099_),
    .Q(\dtop.field_top.fy[4] ));
 sg13g2_dfrbp_1 _6581_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net254),
    .D(net414),
    .Q_N(_0098_),
    .Q(\dtop.field_top.fy[5] ));
 sg13g2_dfrbp_1 _6582_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net253),
    .D(net316),
    .Q_N(_0093_),
    .Q(\dtop.field_top.fy[6] ));
 sg13g2_dfrbp_1 _6583_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net252),
    .D(net309),
    .Q_N(_0106_),
    .Q(\dtop.field_top.fy[7] ));
 sg13g2_dfrbp_1 _6584_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net251),
    .D(net352),
    .Q_N(_0104_),
    .Q(\dtop.field_top.fy[8] ));
 sg13g2_dfrbp_1 _6585_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net248),
    .D(_0147_),
    .Q_N(_0064_),
    .Q(\dtop.field_top.fx[0] ));
 sg13g2_dfrbp_1 _6586_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net247),
    .D(_0148_),
    .Q_N(_0070_),
    .Q(\dtop.field_top.fx[1] ));
 sg13g2_dfrbp_1 _6587_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net246),
    .D(net615),
    .Q_N(_0072_),
    .Q(\dtop.field_top.fx[2] ));
 sg13g2_dfrbp_1 _6588_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net244),
    .D(_0150_),
    .Q_N(_0074_),
    .Q(\dtop.field_top.fx[3] ));
 sg13g2_dfrbp_1 _6589_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net243),
    .D(net486),
    .Q_N(_0025_),
    .Q(\dtop.field_top.fx[4] ));
 sg13g2_dfrbp_1 _6590_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net242),
    .D(net381),
    .Q_N(_0096_),
    .Q(\dtop.field_top.fx[5] ));
 sg13g2_dfrbp_1 _6591_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net241),
    .D(net409),
    .Q_N(_0094_),
    .Q(\dtop.field_top.fx[6] ));
 sg13g2_dfrbp_1 _6592_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net240),
    .D(net378),
    .Q_N(_0091_),
    .Q(\dtop.field_top.fx[7] ));
 sg13g2_dfrbp_1 _6593_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net239),
    .D(net513),
    .Q_N(_0103_),
    .Q(\dtop.field_top.fx[8] ));
 sg13g2_dfrbp_1 _6594_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net238),
    .D(net371),
    .Q_N(_0101_),
    .Q(\dtop.field_top.fx[9] ));
 sg13g2_dfrbp_1 _6595_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net237),
    .D(_0157_),
    .Q_N(_3265_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _6596_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net236),
    .D(_0158_),
    .Q_N(_3264_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _6597_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net235),
    .D(_0159_),
    .Q_N(_3263_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _6598_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net234),
    .D(_0160_),
    .Q_N(_3262_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _6599_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net233),
    .D(_0161_),
    .Q_N(_3261_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _6600_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net232),
    .D(_0162_),
    .Q_N(_3260_),
    .Q(_0006_));
 sg13g2_dfrbp_1 _6601_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net231),
    .D(_0163_),
    .Q_N(_3259_),
    .Q(_0005_));
 sg13g2_dfrbp_1 _6602_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net230),
    .D(_0164_),
    .Q_N(\dtop.field_top.player.controller.timer[1] ),
    .Q(\dtop.field_top.player.osc0[11] ));
 sg13g2_dfrbp_1 _6603_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net228),
    .D(_0165_),
    .Q_N(\dtop.field_top.player.controller.timer[2] ),
    .Q(\dtop.field_top.player.osc0[12] ));
 sg13g2_dfrbp_1 _6604_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net226),
    .D(_0166_),
    .Q_N(\dtop.field_top.player.controller.ppos[0] ),
    .Q(\dtop.field_top.player.osc0[13] ));
 sg13g2_dfrbp_1 _6605_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net224),
    .D(_0167_),
    .Q_N(\dtop.field_top.player.controller.ppos[1] ),
    .Q(\dtop.field_top.player.osc0[14] ));
 sg13g2_dfrbp_1 _6606_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net222),
    .D(_0168_),
    .Q_N(\dtop.field_top.player.controller.ppos[2] ),
    .Q(\dtop.field_top.player.osc0[15] ));
 sg13g2_dfrbp_1 _6607_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net220),
    .D(_0169_),
    .Q_N(\dtop.field_top.player.controller.ppos[3] ),
    .Q(\dtop.field_top.player.osc0[16] ));
 sg13g2_dfrbp_1 _6608_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net218),
    .D(_0170_),
    .Q_N(\dtop.field_top.player.controller.ppos[4] ),
    .Q(\dtop.field_top.player.osc0[17] ));
 sg13g2_dfrbp_1 _6609_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net216),
    .D(_0171_),
    .Q_N(\dtop.field_top.player.controller.ppos[5] ),
    .Q(\dtop.field_top.player.osc0[18] ));
 sg13g2_dfrbp_1 _6610_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net214),
    .D(_0172_),
    .Q_N(\dtop.field_top.player.controller.ppos[6] ),
    .Q(\dtop.field_top.player.osc0[19] ));
 sg13g2_dfrbp_1 _6611_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net212),
    .D(_0173_),
    .Q_N(\dtop.field_top.player.controller.pattern0[0] ),
    .Q(\dtop.field_top.player.osc0[20] ));
 sg13g2_dfrbp_1 _6612_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net210),
    .D(_0174_),
    .Q_N(\dtop.field_top.player.controller.pattern0[1] ),
    .Q(\dtop.field_top.player.osc0[21] ));
 sg13g2_dfrbp_1 _6613_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net208),
    .D(_0175_),
    .Q_N(_0022_),
    .Q(\dtop.field_top.fx[10] ));
 sg13g2_dfrbp_1 _6614_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net206),
    .D(net373),
    .Q_N(_0083_),
    .Q(\dtop.field_top.logo_prev_pixel ));
 sg13g2_dfrbp_1 _6615_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net205),
    .D(_0177_),
    .Q_N(_3258_),
    .Q(\dtop.field_top.masked_bits[0] ));
 sg13g2_dfrbp_1 _6616_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net204),
    .D(_0178_),
    .Q_N(_3257_),
    .Q(\dtop.field_top.masked_bits[1] ));
 sg13g2_dfrbp_1 _6617_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net203),
    .D(_0179_),
    .Q_N(_3256_),
    .Q(\dtop.field_top.sflag2 ));
 sg13g2_dfrbp_1 _6618_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net202),
    .D(_0180_),
    .Q_N(_3255_),
    .Q(\dtop.field_top.sflag ));
 sg13g2_dfrbp_1 _6619_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net201),
    .D(net366),
    .Q_N(_3254_),
    .Q(\dtop.field_top.last_wave[0] ));
 sg13g2_dfrbp_1 _6620_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net200),
    .D(net332),
    .Q_N(_3253_),
    .Q(\dtop.field_top.last_wave[1] ));
 sg13g2_dfrbp_1 _6621_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net199),
    .D(_0183_),
    .Q_N(_3252_),
    .Q(\dtop.field_top.last_wave[2] ));
 sg13g2_dfrbp_1 _6622_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net198),
    .D(_0184_),
    .Q_N(_3251_),
    .Q(\dtop.field_top.last_wave[3] ));
 sg13g2_dfrbp_1 _6623_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net197),
    .D(net303),
    .Q_N(_3250_),
    .Q(\dtop.field_top.last_wave[4] ));
 sg13g2_dfrbp_1 _6624_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net196),
    .D(_0186_),
    .Q_N(_3249_),
    .Q(\dtop.field_top.last_wave[5] ));
 sg13g2_dfrbp_1 _6625_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net195),
    .D(_0187_),
    .Q_N(_3248_),
    .Q(\dtop.field_top.last_wave[6] ));
 sg13g2_dfrbp_1 _6626_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net89),
    .D(net313),
    .Q_N(_0081_),
    .Q(\dtop.field_top.last_wave[7] ));
 sg13g2_dfrbp_1 _6627_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net245),
    .D(_0000_),
    .Q_N(_3270_),
    .Q(_0399_));
 sg13g2_dfrbp_1 _6628_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net194),
    .D(_0001_),
    .Q_N(_3247_),
    .Q(_0397_));
 sg13g2_dfrbp_1 _6629_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net193),
    .D(_0189_),
    .Q_N(_3246_),
    .Q(\dtop.field_top.prev_wave[0] ));
 sg13g2_dfrbp_1 _6630_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net192),
    .D(_0190_),
    .Q_N(_3245_),
    .Q(\dtop.field_top.prev_wave[1] ));
 sg13g2_dfrbp_1 _6631_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net191),
    .D(net419),
    .Q_N(_3244_),
    .Q(\dtop.field_top.prev_wave[2] ));
 sg13g2_dfrbp_1 _6632_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net190),
    .D(net401),
    .Q_N(_3243_),
    .Q(\dtop.field_top.prev_wave[3] ));
 sg13g2_dfrbp_1 _6633_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net189),
    .D(_0193_),
    .Q_N(_3242_),
    .Q(\dtop.field_top.prev_wave[4] ));
 sg13g2_dfrbp_1 _6634_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net188),
    .D(net417),
    .Q_N(_3241_),
    .Q(\dtop.field_top.prev_wave[5] ));
 sg13g2_dfrbp_1 _6635_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net187),
    .D(_0195_),
    .Q_N(_3240_),
    .Q(\dtop.field_top.prev_wave[6] ));
 sg13g2_dfrbp_1 _6636_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net186),
    .D(_0196_),
    .Q_N(_3239_),
    .Q(\dtop.field_top.prev_wave[7] ));
 sg13g2_dfrbp_1 _6637_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net185),
    .D(net368),
    .Q_N(_3238_),
    .Q(\dtop.field_top.comp_value0[0] ));
 sg13g2_dfrbp_1 _6638_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net184),
    .D(net542),
    .Q_N(_3237_),
    .Q(\dtop.field_top.comp_value0[1] ));
 sg13g2_dfrbp_1 _6639_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net183),
    .D(net442),
    .Q_N(_3236_),
    .Q(\dtop.field_top.comp_value0[2] ));
 sg13g2_dfrbp_1 _6640_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net182),
    .D(net433),
    .Q_N(_3235_),
    .Q(\dtop.field_top.comp_value0[3] ));
 sg13g2_dfrbp_1 _6641_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net181),
    .D(net546),
    .Q_N(_3234_),
    .Q(\dtop.field_top.comp_value0[4] ));
 sg13g2_dfrbp_1 _6642_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net180),
    .D(net534),
    .Q_N(_3233_),
    .Q(\dtop.field_top.comp_value0[5] ));
 sg13g2_dfrbp_1 _6643_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net179),
    .D(net406),
    .Q_N(_3232_),
    .Q(\dtop.field_top.comp_value0[6] ));
 sg13g2_dfrbp_1 _6644_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net178),
    .D(net397),
    .Q_N(_3231_),
    .Q(\dtop.field_top.comp_value0[7] ));
 sg13g2_dfrbp_1 _6645_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net177),
    .D(net563),
    .Q_N(_3230_),
    .Q(\dtop.field_top.comp_value0[8] ));
 sg13g2_dfrbp_1 _6646_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net176),
    .D(net557),
    .Q_N(_3229_),
    .Q(\dtop.field_top.comp_value0_0[10] ));
 sg13g2_dfrbp_1 _6647_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net175),
    .D(net334),
    .Q_N(_3228_),
    .Q(\dtop.field_top.wave[0] ));
 sg13g2_dfrbp_1 _6648_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net173),
    .D(net376),
    .Q_N(_3227_),
    .Q(\dtop.field_top.wave[1] ));
 sg13g2_dfrbp_1 _6649_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net171),
    .D(net538),
    .Q_N(_3226_),
    .Q(\dtop.field_top.wave[2] ));
 sg13g2_dfrbp_1 _6650_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net169),
    .D(net617),
    .Q_N(_3225_),
    .Q(\dtop.field_top.wave[3] ));
 sg13g2_dfrbp_1 _6651_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net167),
    .D(_0211_),
    .Q_N(_3224_),
    .Q(\dtop.field_top.wave[4] ));
 sg13g2_dfrbp_1 _6652_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net165),
    .D(net439),
    .Q_N(_3223_),
    .Q(\dtop.field_top.wave[5] ));
 sg13g2_dfrbp_1 _6653_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net163),
    .D(net343),
    .Q_N(_3222_),
    .Q(\dtop.field_top.wave[6] ));
 sg13g2_dfrbp_1 _6654_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net161),
    .D(net328),
    .Q_N(_0080_),
    .Q(\dtop.field_top.wave[7] ));
 sg13g2_dfrbp_1 _6655_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net159),
    .D(net391),
    .Q_N(_0056_),
    .Q(\dtop.field_top.comp_value0_1[0] ));
 sg13g2_dfrbp_1 _6656_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net158),
    .D(net330),
    .Q_N(_0030_),
    .Q(\dtop.field_top.comp_value0_1[1] ));
 sg13g2_dfrbp_1 _6657_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net157),
    .D(net361),
    .Q_N(_0049_),
    .Q(\dtop.field_top.comp_value0_1[2] ));
 sg13g2_dfrbp_1 _6658_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net156),
    .D(net460),
    .Q_N(_0050_),
    .Q(\dtop.field_top.comp_value0_1[3] ));
 sg13g2_dfrbp_1 _6659_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net155),
    .D(net421),
    .Q_N(_0051_),
    .Q(\dtop.field_top.comp_value0_1[4] ));
 sg13g2_dfrbp_1 _6660_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net154),
    .D(net427),
    .Q_N(_0057_),
    .Q(\dtop.field_top.comp_value0_1[5] ));
 sg13g2_dfrbp_1 _6661_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net153),
    .D(net474),
    .Q_N(_0058_),
    .Q(\dtop.field_top.comp_value0_1[6] ));
 sg13g2_dfrbp_1 _6662_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net152),
    .D(net437),
    .Q_N(_0059_),
    .Q(\dtop.field_top.comp_value0_1[7] ));
 sg13g2_dfrbp_1 _6663_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net151),
    .D(net496),
    .Q_N(_0060_),
    .Q(\dtop.field_top.comp_value0_1[8] ));
 sg13g2_dfrbp_1 _6664_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net150),
    .D(net559),
    .Q_N(_0028_),
    .Q(\dtop.field_top.comp_value0_1[9] ));
 sg13g2_dfrbp_1 _6665_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net149),
    .D(net504),
    .Q_N(_0052_),
    .Q(\dtop.field_top.comp_value0_1[10] ));
 sg13g2_dfrbp_1 _6666_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net148),
    .D(net393),
    .Q_N(_0047_),
    .Q(\dtop.field_top.reg1[11] ));
 sg13g2_dfrbp_1 _6667_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net147),
    .D(net383),
    .Q_N(_0045_),
    .Q(\dtop.field_top.reg1[12] ));
 sg13g2_dfrbp_1 _6668_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net146),
    .D(net411),
    .Q_N(_0043_),
    .Q(\dtop.field_top.reg1[13] ));
 sg13g2_dfrbp_1 _6669_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net145),
    .D(net388),
    .Q_N(_0041_),
    .Q(\dtop.field_top.reg1[14] ));
 sg13g2_dfrbp_1 _6670_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net144),
    .D(net311),
    .Q_N(_0039_),
    .Q(\dtop.field_top.reg1[15] ));
 sg13g2_dfrbp_1 _6671_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net143),
    .D(net395),
    .Q_N(_0054_),
    .Q(\dtop.field_top.reg1[16] ));
 sg13g2_dfrbp_1 _6672_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net142),
    .D(net458),
    .Q_N(_3221_),
    .Q(\dtop.field_top.comp_values0[2][0] ));
 sg13g2_dfrbp_1 _6673_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net141),
    .D(net544),
    .Q_N(_3220_),
    .Q(\dtop.field_top.comp_values0[2][1] ));
 sg13g2_dfrbp_1 _6674_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net140),
    .D(net500),
    .Q_N(_3219_),
    .Q(\dtop.field_top.comp_values0[2][2] ));
 sg13g2_dfrbp_1 _6675_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net139),
    .D(net594),
    .Q_N(_3218_),
    .Q(\dtop.field_top.comp_values0[2][3] ));
 sg13g2_dfrbp_1 _6676_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net138),
    .D(net552),
    .Q_N(_3217_),
    .Q(\dtop.field_top.comp_values0[2][4] ));
 sg13g2_dfrbp_1 _6677_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net137),
    .D(net624),
    .Q_N(_3216_),
    .Q(\dtop.field_top.comp_values0[2][5] ));
 sg13g2_dfrbp_1 _6678_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net136),
    .D(net598),
    .Q_N(_3215_),
    .Q(\dtop.field_top.comp_values0[2][6] ));
 sg13g2_dfrbp_1 _6679_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net135),
    .D(_0239_),
    .Q_N(_3214_),
    .Q(\dtop.field_top.comp_values0[2][7] ));
 sg13g2_dfrbp_1 _6680_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net134),
    .D(net607),
    .Q_N(_3213_),
    .Q(\dtop.field_top.comp_values0[2][8] ));
 sg13g2_dfrbp_1 _6681_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net133),
    .D(net647),
    .Q_N(_3212_),
    .Q(\dtop.field_top.comp_values0[2][9] ));
 sg13g2_dfrbp_1 _6682_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net132),
    .D(net578),
    .Q_N(_3211_),
    .Q(\dtop.field_top.comp_values0[2][10] ));
 sg13g2_dfrbp_1 _6683_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net131),
    .D(net492),
    .Q_N(_3210_),
    .Q(\dtop.field_top.reg2[11] ));
 sg13g2_dfrbp_1 _6684_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net130),
    .D(net454),
    .Q_N(_3209_),
    .Q(\dtop.field_top.reg2[12] ));
 sg13g2_dfrbp_1 _6685_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net129),
    .D(net462),
    .Q_N(_3208_),
    .Q(\dtop.field_top.reg2[13] ));
 sg13g2_dfrbp_1 _6686_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net128),
    .D(net450),
    .Q_N(_3207_),
    .Q(\dtop.field_top.reg2[14] ));
 sg13g2_dfrbp_1 _6687_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net127),
    .D(net506),
    .Q_N(_3206_),
    .Q(\dtop.field_top.reg2[15] ));
 sg13g2_dfrbp_1 _6688_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net126),
    .D(net536),
    .Q_N(_3205_),
    .Q(\dtop.field_top.reg2[16] ));
 sg13g2_dfrbp_1 _6689_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net125),
    .D(net480),
    .Q_N(_3204_),
    .Q(\dtop.field_top.comp_values0[3][0] ));
 sg13g2_dfrbp_1 _6690_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net124),
    .D(net357),
    .Q_N(_3203_),
    .Q(\dtop.field_top.comp_values0[3][1] ));
 sg13g2_dfrbp_1 _6691_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net123),
    .D(net430),
    .Q_N(_3202_),
    .Q(\dtop.field_top.comp_values0[3][2] ));
 sg13g2_dfrbp_1 _6692_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net122),
    .D(net531),
    .Q_N(_3201_),
    .Q(\dtop.field_top.comp_values0[3][3] ));
 sg13g2_dfrbp_1 _6693_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net121),
    .D(net515),
    .Q_N(_3200_),
    .Q(\dtop.field_top.comp_values0[3][4] ));
 sg13g2_dfrbp_1 _6694_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net120),
    .D(net540),
    .Q_N(_3199_),
    .Q(\dtop.field_top.comp_values0[3][5] ));
 sg13g2_dfrbp_1 _6695_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net119),
    .D(net502),
    .Q_N(_3198_),
    .Q(\dtop.field_top.comp_values0[3][6] ));
 sg13g2_dfrbp_1 _6696_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net118),
    .D(net494),
    .Q_N(_3197_),
    .Q(\dtop.field_top.comp_values0[3][7] ));
 sg13g2_dfrbp_1 _6697_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net117),
    .D(net555),
    .Q_N(_3196_),
    .Q(\dtop.field_top.comp_values0[3][8] ));
 sg13g2_dfrbp_1 _6698_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net116),
    .D(net626),
    .Q_N(_3195_),
    .Q(\dtop.field_top.comp_values0[3][9] ));
 sg13g2_dfrbp_1 _6699_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net115),
    .D(net574),
    .Q_N(_3194_),
    .Q(\dtop.field_top.comp_values0[3][10] ));
 sg13g2_dfrbp_1 _6700_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net114),
    .D(net476),
    .Q_N(_3193_),
    .Q(\dtop.field_top.reg3[11] ));
 sg13g2_dfrbp_1 _6701_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net113),
    .D(net444),
    .Q_N(_3192_),
    .Q(\dtop.field_top.reg3[12] ));
 sg13g2_dfrbp_1 _6702_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net112),
    .D(net446),
    .Q_N(_3191_),
    .Q(\dtop.field_top.reg3[13] ));
 sg13g2_dfrbp_1 _6703_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net111),
    .D(net517),
    .Q_N(_3190_),
    .Q(\dtop.field_top.reg3[14] ));
 sg13g2_dfrbp_1 _6704_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net110),
    .D(net338),
    .Q_N(_3189_),
    .Q(\dtop.field_top.reg3[15] ));
 sg13g2_dfrbp_1 _6705_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net109),
    .D(net468),
    .Q_N(_3188_),
    .Q(\dtop.field_top.reg3[16] ));
 sg13g2_dfrbp_1 _6706_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net108),
    .D(net519),
    .Q_N(_3187_),
    .Q(\dtop.field_top.comp_values0[4][0] ));
 sg13g2_dfrbp_1 _6707_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net107),
    .D(net490),
    .Q_N(_3186_),
    .Q(\dtop.field_top.comp_values0[4][1] ));
 sg13g2_dfrbp_1 _6708_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net106),
    .D(net525),
    .Q_N(_3185_),
    .Q(\dtop.field_top.comp_values0[4][2] ));
 sg13g2_dfrbp_1 _6709_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net105),
    .D(net568),
    .Q_N(_3184_),
    .Q(\dtop.field_top.comp_values0[4][3] ));
 sg13g2_dfrbp_1 _6710_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net104),
    .D(net529),
    .Q_N(_3183_),
    .Q(\dtop.field_top.comp_values0[4][4] ));
 sg13g2_dfrbp_1 _6711_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net103),
    .D(net590),
    .Q_N(_3182_),
    .Q(\dtop.field_top.comp_values0[4][5] ));
 sg13g2_dfrbp_1 _6712_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net102),
    .D(net632),
    .Q_N(_3181_),
    .Q(\dtop.field_top.comp_values0[4][6] ));
 sg13g2_dfrbp_1 _6713_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net101),
    .D(_0273_),
    .Q_N(_3180_),
    .Q(\dtop.field_top.comp_values0[4][7] ));
 sg13g2_dfrbp_1 _6714_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net100),
    .D(net596),
    .Q_N(_3179_),
    .Q(\dtop.field_top.comp_values0[4][8] ));
 sg13g2_dfrbp_1 _6715_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net99),
    .D(net508),
    .Q_N(_3178_),
    .Q(\dtop.field_top.comp_values0[4][9] ));
 sg13g2_dfrbp_1 _6716_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net98),
    .D(net609),
    .Q_N(_3177_),
    .Q(\dtop.field_top.comp_values0[4][10] ));
 sg13g2_dfrbp_1 _6717_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net97),
    .D(net470),
    .Q_N(_3176_),
    .Q(\dtop.field_top.reg4[11] ));
 sg13g2_dfrbp_1 _6718_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net96),
    .D(net466),
    .Q_N(_3175_),
    .Q(\dtop.field_top.reg4[12] ));
 sg13g2_dfrbp_1 _6719_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net95),
    .D(net448),
    .Q_N(_3174_),
    .Q(\dtop.field_top.reg4[13] ));
 sg13g2_dfrbp_1 _6720_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net94),
    .D(net548),
    .Q_N(_3173_),
    .Q(\dtop.field_top.reg4[14] ));
 sg13g2_dfrbp_1 _6721_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net93),
    .D(net349),
    .Q_N(_3172_),
    .Q(\dtop.field_top.reg4[15] ));
 sg13g2_dfrbp_1 _6722_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net92),
    .D(net456),
    .Q_N(_3171_),
    .Q(\dtop.field_top.reg4[16] ));
 sg13g2_dfrbp_1 _6723_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net91),
    .D(net561),
    .Q_N(_0082_),
    .Q(\dtop.field_top.lside ));
 sg13g2_dfrbp_1 _6724_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net90),
    .D(net585),
    .Q_N(_3170_),
    .Q(\dtop.field_top.rside ));
 sg13g2_dfrbp_1 _6725_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net87),
    .D(_0285_),
    .Q_N(_3169_),
    .Q(_0400_));
 sg13g2_dfrbp_1 _6726_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net86),
    .D(_0286_),
    .Q_N(_3168_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _6727_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net85),
    .D(_0287_),
    .Q_N(_3167_),
    .Q(_0396_));
 sg13g2_dfrbp_1 _6728_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net84),
    .D(_0288_),
    .Q_N(_3166_),
    .Q(\dtop.field_top.rs.scan_x.state[0] ));
 sg13g2_dfrbp_1 _6729_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net83),
    .D(_0289_),
    .Q_N(_3165_),
    .Q(\dtop.field_top.rs.scan_x.state[1] ));
 sg13g2_dfrbp_1 _6730_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net82),
    .D(_0290_),
    .Q_N(_0010_),
    .Q(\dtop.field_top.alt_osc[1] ));
 sg13g2_dfrbp_1 _6731_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net81),
    .D(_0291_),
    .Q_N(_0011_),
    .Q(\dtop.field_top.alt_osc[2] ));
 sg13g2_dfrbp_1 _6732_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net80),
    .D(_0292_),
    .Q_N(_0013_),
    .Q(\dtop.field_top.alt_osc[3] ));
 sg13g2_dfrbp_1 _6733_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net79),
    .D(net592),
    .Q_N(_0012_),
    .Q(\dtop.field_top.alt_osc[4] ));
 sg13g2_dfrbp_1 _6734_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net78),
    .D(_0294_),
    .Q_N(_0069_),
    .Q(\dtop.field_top.alt_osc[5] ));
 sg13g2_dfrbp_1 _6735_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net77),
    .D(_0295_),
    .Q_N(_0014_),
    .Q(\dtop.field_top.alt_osc[6] ));
 sg13g2_dfrbp_1 _6736_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net76),
    .D(_0296_),
    .Q_N(_0015_),
    .Q(\dtop.field_top.alt_osc[7] ));
 sg13g2_dfrbp_1 _6737_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net75),
    .D(_0297_),
    .Q_N(_0016_),
    .Q(\dtop.field_top.alt_osc[8] ));
 sg13g2_dfrbp_1 _6738_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net74),
    .D(_0298_),
    .Q_N(_0109_),
    .Q(\dtop.field_top.rs.scan_y.pos[8] ));
 sg13g2_dfrbp_1 _6739_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net73),
    .D(_0299_),
    .Q_N(_3164_),
    .Q(\dtop.field_top.rs.scan_y.pos[9] ));
 sg13g2_dfrbp_1 _6740_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net72),
    .D(_0300_),
    .Q_N(_3163_),
    .Q(\dtop.field_top.player.sched.alu.p0 ));
 sg13g2_dfrbp_1 _6741_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net71),
    .D(_0301_),
    .Q_N(_0116_),
    .Q(\dtop.field_top.afl_sub_pc[0] ));
 sg13g2_dfrbp_1 _6742_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net70),
    .D(net687),
    .Q_N(_0066_),
    .Q(\dtop.field_top.afl_sub_pc[1] ));
 sg13g2_dfrbp_1 _6743_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net69),
    .D(_0303_),
    .Q_N(_0067_),
    .Q(\dtop.field_top.afl_pc[0] ));
 sg13g2_dfrbp_1 _6744_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net68),
    .D(_0304_),
    .Q_N(_3162_),
    .Q(\dtop.field_top.afl_pc[1] ));
 sg13g2_dfrbp_1 _6745_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net67),
    .D(_0305_),
    .Q_N(_0008_),
    .Q(\dtop.field_top.afl_pc[2] ));
 sg13g2_dfrbp_1 _6746_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net66),
    .D(_0306_),
    .Q_N(_0068_),
    .Q(\dtop.field_top.afl_pc[3] ));
 sg13g2_dfrbp_1 _6747_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net65),
    .D(_0307_),
    .Q_N(_0009_),
    .Q(\dtop.field_top.afl_pc[4] ));
 sg13g2_dfrbp_1 _6748_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net64),
    .D(_0308_),
    .Q_N(_0019_),
    .Q(\dtop.field_top.afl_pc[5] ));
 sg13g2_dfrbp_1 _6749_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net63),
    .D(_0309_),
    .Q_N(_0018_),
    .Q(\dtop.field_top.afl_pc[6] ));
 sg13g2_dfrbp_1 _6750_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net62),
    .D(_0310_),
    .Q_N(_0017_),
    .Q(\dtop.field_top.afl_pc[7] ));
 sg13g2_dfrbp_1 _6751_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net61),
    .D(_0311_),
    .Q_N(_0107_),
    .Q(\dtop.field_top.afl_pc[8] ));
 sg13g2_dfrbp_1 _6752_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net60),
    .D(net347),
    .Q_N(_0100_),
    .Q(\dtop.field_top.nsource.shuffle_state.in[0] ));
 sg13g2_dfrbp_1 _6753_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net59),
    .D(_0313_),
    .Q_N(_3161_),
    .Q(\dtop.field_top.nsource.shuffle_state.in[1] ));
 sg13g2_dfrbp_1 _6754_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net58),
    .D(net340),
    .Q_N(_0023_),
    .Q(\dtop.field_top.nsource.shuffle_state.in[2] ));
 sg13g2_dfrbp_1 _6755_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net57),
    .D(net326),
    .Q_N(_0102_),
    .Q(\dtop.field_top.nsource.shuffle_state.in[3] ));
 sg13g2_dfrbp_1 _6756_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net56),
    .D(net321),
    .Q_N(_0097_),
    .Q(\dtop.field_top.nsource.shuffle_state.in[4] ));
 sg13g2_dfrbp_1 _6757_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net55),
    .D(_0317_),
    .Q_N(_0095_),
    .Q(\dtop.field_top.nsource.shuffle_state.in[5] ));
 sg13g2_dfrbp_1 _6758_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net54),
    .D(net345),
    .Q_N(_0092_),
    .Q(\dtop.field_top.nsource.shuffle_state.in[6] ));
 sg13g2_dfrbp_1 _6759_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net53),
    .D(net336),
    .Q_N(_0105_),
    .Q(\dtop.field_top.nsource.shuffle_state.in[7] ));
 sg13g2_dfrbp_1 _6760_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net52),
    .D(_0320_),
    .Q_N(_0063_),
    .Q(\dtop.field_top.afl_alu.last_r_sum_msbs[0] ));
 sg13g2_dfrbp_1 _6761_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net51),
    .D(_0321_),
    .Q_N(_3160_),
    .Q(\dtop.field_top.afl_alu.last_r_sum_msbs[1] ));
 sg13g2_dfrbp_1 _6762_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net50),
    .D(_0322_),
    .Q_N(_3159_),
    .Q(\dtop.field_top.afl_alu.p ));
 sg13g2_dfrbp_1 _6763_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net49),
    .D(_0323_),
    .Q_N(_0055_),
    .Q(\dtop.field_top.acc[0] ));
 sg13g2_dfrbp_1 _6764_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net47),
    .D(_0324_),
    .Q_N(_0029_),
    .Q(\dtop.field_top.acc[1] ));
 sg13g2_dfrbp_1 _6765_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net45),
    .D(_0325_),
    .Q_N(_0048_),
    .Q(\dtop.field_top.acc[2] ));
 sg13g2_dfrbp_1 _6766_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net43),
    .D(_0326_),
    .Q_N(_0037_),
    .Q(\dtop.field_top.acc[3] ));
 sg13g2_dfrbp_1 _6767_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net41),
    .D(_0327_),
    .Q_N(_0036_),
    .Q(\dtop.field_top.acc[4] ));
 sg13g2_dfrbp_1 _6768_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net39),
    .D(_0328_),
    .Q_N(_0035_),
    .Q(\dtop.field_top.acc[5] ));
 sg13g2_dfrbp_1 _6769_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net37),
    .D(_0329_),
    .Q_N(_0034_),
    .Q(\dtop.field_top.acc[6] ));
 sg13g2_dfrbp_1 _6770_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net35),
    .D(_0330_),
    .Q_N(_0033_),
    .Q(\dtop.field_top.acc[7] ));
 sg13g2_dfrbp_1 _6771_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net33),
    .D(net435),
    .Q_N(_3158_),
    .Q(\dtop.field_top.controller.timer[0] ));
 sg13g2_dfrbp_1 _6772_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net32),
    .D(net478),
    .Q_N(_3157_),
    .Q(\dtop.field_top.controller.timer[1] ));
 sg13g2_dfrbp_1 _6773_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net31),
    .D(net472),
    .Q_N(_0075_),
    .Q(\dtop.field_top.controller.timer[2] ));
 sg13g2_dfrbp_1 _6774_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net30),
    .D(net650),
    .Q_N(_0076_),
    .Q(\dtop.field_top.controller.ppos[0] ));
 sg13g2_dfrbp_1 _6775_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net29),
    .D(net645),
    .Q_N(_0062_),
    .Q(\dtop.field_top.controller.ppos[1] ));
 sg13g2_dfrbp_1 _6776_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net28),
    .D(_0336_),
    .Q_N(_0061_),
    .Q(\dtop.field_top.controller.ppos[2] ));
 sg13g2_dfrbp_1 _6777_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net27),
    .D(_0337_),
    .Q_N(_0021_),
    .Q(\dtop.field_top.controller.ppos[3] ));
 sg13g2_dfrbp_1 _6778_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net26),
    .D(_0338_),
    .Q_N(_0020_),
    .Q(\dtop.field_top.controller.ppos[4] ));
 sg13g2_dfrbp_1 _6779_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net25),
    .D(_0339_),
    .Q_N(_0077_),
    .Q(\dtop.field_top.controller.ppos[5] ));
 sg13g2_dfrbp_1 _6780_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net24),
    .D(net689),
    .Q_N(_0078_),
    .Q(\dtop.field_top.controller.ppos[6] ));
 sg13g2_dfrbp_1 _6781_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net23),
    .D(net588),
    .Q_N(_0079_),
    .Q(\dtop.field_top.controller.pattern0[0] ));
 sg13g2_dfrbp_1 _6782_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net22),
    .D(net424),
    .Q_N(_3156_),
    .Q(\dtop.field_top.controller.pattern0[1] ));
 sg13g2_dfrbp_1 _6783_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net249),
    .D(net675),
    .Q_N(_0108_),
    .Q(\dtop.field_top.controller.pattern0[2] ));
 sg13g2_dfrbp_1 _6784_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net21),
    .D(\dtop.field_top.player.out_pw_high ),
    .Q_N(_3155_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _6785_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net20),
    .D(_0344_),
    .Q_N(\dtop.field_top.player.controller.pattern0[2] ),
    .Q(\dtop.field_top.player.osc0[22] ));
 sg13g2_dfrbp_1 _6786_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net18),
    .D(_0345_),
    .Q_N(_3154_),
    .Q(_0398_));
 sg13g2_dfrbp_1 _6787_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net250),
    .D(_0346_),
    .Q_N(_3271_),
    .Q(_0401_));
 sg13g2_dfrbp_1 _6788_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net293),
    .D(\dtop.field_top.rs.vsync ),
    .Q_N(_3272_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _6789_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net17),
    .D(\dtop.field_top.hsync ),
    .Q_N(_3153_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _6790_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net300),
    .D(_0347_),
    .Q_N(_3152_),
    .Q(\dtop.field_top.player.out_acc[0] ));
 sg13g2_dfrbp_1 _6791_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net298),
    .D(_0348_),
    .Q_N(_3151_),
    .Q(\dtop.field_top.player.out_acc[1] ));
 sg13g2_dfrbp_1 _6792_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net296),
    .D(_0349_),
    .Q_N(_3150_),
    .Q(\dtop.field_top.player.out_acc[2] ));
 sg13g2_dfrbp_1 _6793_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net292),
    .D(_0350_),
    .Q_N(_3149_),
    .Q(\dtop.field_top.player.out_acc[3] ));
 sg13g2_dfrbp_1 _6794_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net290),
    .D(_0351_),
    .Q_N(_3148_),
    .Q(\dtop.field_top.player.out_acc[4] ));
 sg13g2_dfrbp_1 _6795_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net288),
    .D(_0352_),
    .Q_N(_3147_),
    .Q(\dtop.field_top.player.out_acc[5] ));
 sg13g2_dfrbp_1 _6796_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net286),
    .D(_0353_),
    .Q_N(_3146_),
    .Q(\dtop.field_top.player.out_acc[6] ));
 sg13g2_dfrbp_1 _6797_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net274),
    .D(_0354_),
    .Q_N(_3145_),
    .Q(\dtop.field_top.player.out_acc[7] ));
 sg13g2_dfrbp_1 _6798_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net270),
    .D(_0355_),
    .Q_N(_3144_),
    .Q(\dtop.field_top.player.out_acc[8] ));
 sg13g2_dfrbp_1 _6799_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net262),
    .D(_0356_),
    .Q_N(_3143_),
    .Q(\dtop.field_top.player.out_acc[9] ));
 sg13g2_dfrbp_1 _6800_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net229),
    .D(_0357_),
    .Q_N(_3142_),
    .Q(\dtop.field_top.player.osc0[0] ));
 sg13g2_dfrbp_1 _6801_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net225),
    .D(_0358_),
    .Q_N(_3141_),
    .Q(\dtop.field_top.player.osc0[1] ));
 sg13g2_dfrbp_1 _6802_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net221),
    .D(_0359_),
    .Q_N(_3140_),
    .Q(\dtop.field_top.player.osc0[2] ));
 sg13g2_dfrbp_1 _6803_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net217),
    .D(_0360_),
    .Q_N(_0084_),
    .Q(\dtop.field_top.player.osc0[3] ));
 sg13g2_dfrbp_1 _6804_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net213),
    .D(_0361_),
    .Q_N(_0085_),
    .Q(\dtop.field_top.player.osc0[4] ));
 sg13g2_dfrbp_1 _6805_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net209),
    .D(_0362_),
    .Q_N(_0086_),
    .Q(\dtop.field_top.player.osc0[5] ));
 sg13g2_dfrbp_1 _6806_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net174),
    .D(_0363_),
    .Q_N(_0087_),
    .Q(\dtop.field_top.player.osc0[6] ));
 sg13g2_dfrbp_1 _6807_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net170),
    .D(_0364_),
    .Q_N(_0088_),
    .Q(\dtop.field_top.player.osc0[7] ));
 sg13g2_dfrbp_1 _6808_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net166),
    .D(_0365_),
    .Q_N(_0089_),
    .Q(\dtop.field_top.player.osc0[8] ));
 sg13g2_dfrbp_1 _6809_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net162),
    .D(_0366_),
    .Q_N(_0090_),
    .Q(\dtop.field_top.player.osc0[9] ));
 sg13g2_dfrbp_1 _6810_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net48),
    .D(_0367_),
    .Q_N(\dtop.field_top.player.controller.timer[0] ),
    .Q(\dtop.field_top.player.osc0[10] ));
 sg13g2_dfrbp_1 _6811_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net44),
    .D(net581),
    .Q_N(_3139_),
    .Q(\dtop.field_top.player.out_pw[0] ));
 sg13g2_dfrbp_1 _6812_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net42),
    .D(net604),
    .Q_N(_3138_),
    .Q(\dtop.field_top.player.out_pw[1] ));
 sg13g2_dfrbp_1 _6813_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net40),
    .D(net583),
    .Q_N(_3137_),
    .Q(\dtop.field_top.player.out_pw[2] ));
 sg13g2_dfrbp_1 _6814_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net38),
    .D(net523),
    .Q_N(_3136_),
    .Q(\dtop.field_top.player.out_pw[3] ));
 sg13g2_dfrbp_1 _6815_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net36),
    .D(net565),
    .Q_N(_3135_),
    .Q(\dtop.field_top.player.out_pw[4] ));
 sg13g2_dfrbp_1 _6816_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net34),
    .D(net550),
    .Q_N(_3134_),
    .Q(\dtop.field_top.player.out_pw[5] ));
 sg13g2_dfrbp_1 _6817_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net19),
    .D(_0374_),
    .Q_N(_3133_),
    .Q(\dtop.field_top.player.out_pw[6] ));
 sg13g2_dfrbp_1 _6818_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net299),
    .D(net576),
    .Q_N(_3132_),
    .Q(\dtop.field_top.player.out_pw[7] ));
 sg13g2_dfrbp_1 _6819_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net297),
    .D(net521),
    .Q_N(_3131_),
    .Q(\dtop.field_top.player.out_pw[8] ));
 sg13g2_dfrbp_1 _6820_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net295),
    .D(net527),
    .Q_N(_3130_),
    .Q(\dtop.field_top.player.out_pw[9] ));
 sg13g2_dfrbp_1 _6821_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net291),
    .D(_0378_),
    .Q_N(_3129_),
    .Q(\dtop.field_top.channel_output[0] ));
 sg13g2_dfrbp_1 _6822_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net287),
    .D(_0379_),
    .Q_N(_3128_),
    .Q(\dtop.field_top.channel_output[1] ));
 sg13g2_dfrbp_1 _6823_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net272),
    .D(_0380_),
    .Q_N(_3127_),
    .Q(\dtop.field_top.channel_output[2] ));
 sg13g2_dfrbp_1 _6824_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net260),
    .D(_0381_),
    .Q_N(_3126_),
    .Q(\dtop.field_top.channel_output[3] ));
 sg13g2_dfrbp_1 _6825_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net223),
    .D(_0382_),
    .Q_N(_3125_),
    .Q(\dtop.field_top.channel_output[4] ));
 sg13g2_dfrbp_1 _6826_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net215),
    .D(_0383_),
    .Q_N(_3124_),
    .Q(\dtop.field_top.channel_output[5] ));
 sg13g2_dfrbp_1 _6827_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net207),
    .D(_0384_),
    .Q_N(_3123_),
    .Q(\dtop.field_top.channel_output[6] ));
 sg13g2_dfrbp_1 _6828_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net168),
    .D(_0385_),
    .Q_N(_3122_),
    .Q(\dtop.field_top.channel_output[7] ));
 sg13g2_dfrbp_1 _6829_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net160),
    .D(_0386_),
    .Q_N(_3121_),
    .Q(\dtop.field_top.channel_output[8] ));
 sg13g2_dfrbp_1 _6830_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net289),
    .D(_0387_),
    .Q_N(_3120_),
    .Q(\dtop.field_top.channel_output[9] ));
 sg13g2_dfrbp_1 _6831_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net294),
    .D(_0388_),
    .Q_N(_3273_),
    .Q(\dtop.field_top.channel_output[10] ));
 sg13g2_dfrbp_1 _6832_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net227),
    .D(_0002_),
    .Q_N(_3274_),
    .Q(_0004_));
 sg13g2_dfrbp_1 _6833_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net268),
    .D(_0003_),
    .Q_N(_3119_),
    .Q(_0395_));
 sg13g2_dfrbp_1 _6834_ (.CLK(clknet_3_6__leaf_clk),
    .RESET_B(net219),
    .D(_0389_),
    .Q_N(_0113_),
    .Q(\dtop.field_top.player.sched.alu.p1 ));
 sg13g2_dfrbp_1 _6835_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net211),
    .D(net319),
    .Q_N(_3118_),
    .Q(\dtop.field_top.nsource.num_iter[0] ));
 sg13g2_dfrbp_1 _6836_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net172),
    .D(_0391_),
    .Q_N(_3117_),
    .Q(\dtop.field_top.nsource.num_iter[1] ));
 sg13g2_dfrbp_1 _6837_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net164),
    .D(_0392_),
    .Q_N(_0111_),
    .Q(\dtop.field_top.player.chan_timer[5] ));
 sg13g2_dfrbp_1 _6838_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net46),
    .D(_0393_),
    .Q_N(_3116_),
    .Q(\dtop.field_top.channel[0] ));
 sg13g2_dfrbp_1 _6839_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net276),
    .D(_0394_),
    .Q_N(_3115_),
    .Q(\dtop.field_top.channel[3] ));
 sg13g2_tiehi _6786__18 (.L_HI(net18));
 sg13g2_tiehi _6817__19 (.L_HI(net19));
 sg13g2_tiehi _6785__20 (.L_HI(net20));
 sg13g2_tiehi _6784__21 (.L_HI(net21));
 sg13g2_tiehi _6782__22 (.L_HI(net22));
 sg13g2_tiehi _6781__23 (.L_HI(net23));
 sg13g2_tiehi _6780__24 (.L_HI(net24));
 sg13g2_tiehi _6779__25 (.L_HI(net25));
 sg13g2_tiehi _6778__26 (.L_HI(net26));
 sg13g2_tiehi _6777__27 (.L_HI(net27));
 sg13g2_tiehi _6776__28 (.L_HI(net28));
 sg13g2_tiehi _6775__29 (.L_HI(net29));
 sg13g2_tiehi _6774__30 (.L_HI(net30));
 sg13g2_tiehi _6773__31 (.L_HI(net31));
 sg13g2_tiehi _6772__32 (.L_HI(net32));
 sg13g2_tiehi _6771__33 (.L_HI(net33));
 sg13g2_tiehi _6816__34 (.L_HI(net34));
 sg13g2_tiehi _6770__35 (.L_HI(net35));
 sg13g2_tiehi _6815__36 (.L_HI(net36));
 sg13g2_tiehi _6769__37 (.L_HI(net37));
 sg13g2_tiehi _6814__38 (.L_HI(net38));
 sg13g2_tiehi _6768__39 (.L_HI(net39));
 sg13g2_tiehi _6813__40 (.L_HI(net40));
 sg13g2_tiehi _6767__41 (.L_HI(net41));
 sg13g2_tiehi _6812__42 (.L_HI(net42));
 sg13g2_tiehi _6766__43 (.L_HI(net43));
 sg13g2_tiehi _6811__44 (.L_HI(net44));
 sg13g2_tiehi _6765__45 (.L_HI(net45));
 sg13g2_tiehi _6838__46 (.L_HI(net46));
 sg13g2_tiehi _6764__47 (.L_HI(net47));
 sg13g2_tiehi _6810__48 (.L_HI(net48));
 sg13g2_tiehi _6763__49 (.L_HI(net49));
 sg13g2_tiehi _6762__50 (.L_HI(net50));
 sg13g2_tiehi _6761__51 (.L_HI(net51));
 sg13g2_tiehi _6760__52 (.L_HI(net52));
 sg13g2_tiehi _6759__53 (.L_HI(net53));
 sg13g2_tiehi _6758__54 (.L_HI(net54));
 sg13g2_tiehi _6757__55 (.L_HI(net55));
 sg13g2_tiehi _6756__56 (.L_HI(net56));
 sg13g2_tiehi _6755__57 (.L_HI(net57));
 sg13g2_tiehi _6754__58 (.L_HI(net58));
 sg13g2_tiehi _6753__59 (.L_HI(net59));
 sg13g2_tiehi _6752__60 (.L_HI(net60));
 sg13g2_tiehi _6751__61 (.L_HI(net61));
 sg13g2_tiehi _6750__62 (.L_HI(net62));
 sg13g2_tiehi _6749__63 (.L_HI(net63));
 sg13g2_tiehi _6748__64 (.L_HI(net64));
 sg13g2_tiehi _6747__65 (.L_HI(net65));
 sg13g2_tiehi _6746__66 (.L_HI(net66));
 sg13g2_tiehi _6745__67 (.L_HI(net67));
 sg13g2_tiehi _6744__68 (.L_HI(net68));
 sg13g2_tiehi _6743__69 (.L_HI(net69));
 sg13g2_tiehi _6742__70 (.L_HI(net70));
 sg13g2_tiehi _6741__71 (.L_HI(net71));
 sg13g2_tiehi _6740__72 (.L_HI(net72));
 sg13g2_tiehi _6739__73 (.L_HI(net73));
 sg13g2_tiehi _6738__74 (.L_HI(net74));
 sg13g2_tiehi _6737__75 (.L_HI(net75));
 sg13g2_tiehi _6736__76 (.L_HI(net76));
 sg13g2_tiehi _6735__77 (.L_HI(net77));
 sg13g2_tiehi _6734__78 (.L_HI(net78));
 sg13g2_tiehi _6733__79 (.L_HI(net79));
 sg13g2_tiehi _6732__80 (.L_HI(net80));
 sg13g2_tiehi _6731__81 (.L_HI(net81));
 sg13g2_tiehi _6730__82 (.L_HI(net82));
 sg13g2_tiehi _6729__83 (.L_HI(net83));
 sg13g2_tiehi _6728__84 (.L_HI(net84));
 sg13g2_tiehi _6727__85 (.L_HI(net85));
 sg13g2_tiehi _6726__86 (.L_HI(net86));
 sg13g2_tiehi _6725__87 (.L_HI(net87));
 sg13g2_tiehi _6556__88 (.L_HI(net88));
 sg13g2_tiehi _6626__89 (.L_HI(net89));
 sg13g2_tiehi _6724__90 (.L_HI(net90));
 sg13g2_tiehi _6723__91 (.L_HI(net91));
 sg13g2_tiehi _6722__92 (.L_HI(net92));
 sg13g2_tiehi _6721__93 (.L_HI(net93));
 sg13g2_tiehi _6720__94 (.L_HI(net94));
 sg13g2_tiehi _6719__95 (.L_HI(net95));
 sg13g2_tiehi _6718__96 (.L_HI(net96));
 sg13g2_tiehi _6717__97 (.L_HI(net97));
 sg13g2_tiehi _6716__98 (.L_HI(net98));
 sg13g2_tiehi _6715__99 (.L_HI(net99));
 sg13g2_tiehi _6714__100 (.L_HI(net100));
 sg13g2_tiehi _6713__101 (.L_HI(net101));
 sg13g2_tiehi _6712__102 (.L_HI(net102));
 sg13g2_tiehi _6711__103 (.L_HI(net103));
 sg13g2_tiehi _6710__104 (.L_HI(net104));
 sg13g2_tiehi _6709__105 (.L_HI(net105));
 sg13g2_tiehi _6708__106 (.L_HI(net106));
 sg13g2_tiehi _6707__107 (.L_HI(net107));
 sg13g2_tiehi _6706__108 (.L_HI(net108));
 sg13g2_tiehi _6705__109 (.L_HI(net109));
 sg13g2_tiehi _6704__110 (.L_HI(net110));
 sg13g2_tiehi _6703__111 (.L_HI(net111));
 sg13g2_tiehi _6702__112 (.L_HI(net112));
 sg13g2_tiehi _6701__113 (.L_HI(net113));
 sg13g2_tiehi _6700__114 (.L_HI(net114));
 sg13g2_tiehi _6699__115 (.L_HI(net115));
 sg13g2_tiehi _6698__116 (.L_HI(net116));
 sg13g2_tiehi _6697__117 (.L_HI(net117));
 sg13g2_tiehi _6696__118 (.L_HI(net118));
 sg13g2_tiehi _6695__119 (.L_HI(net119));
 sg13g2_tiehi _6694__120 (.L_HI(net120));
 sg13g2_tiehi _6693__121 (.L_HI(net121));
 sg13g2_tiehi _6692__122 (.L_HI(net122));
 sg13g2_tiehi _6691__123 (.L_HI(net123));
 sg13g2_tiehi _6690__124 (.L_HI(net124));
 sg13g2_tiehi _6689__125 (.L_HI(net125));
 sg13g2_tiehi _6688__126 (.L_HI(net126));
 sg13g2_tiehi _6687__127 (.L_HI(net127));
 sg13g2_tiehi _6686__128 (.L_HI(net128));
 sg13g2_tiehi _6685__129 (.L_HI(net129));
 sg13g2_tiehi _6684__130 (.L_HI(net130));
 sg13g2_tiehi _6683__131 (.L_HI(net131));
 sg13g2_tiehi _6682__132 (.L_HI(net132));
 sg13g2_tiehi _6681__133 (.L_HI(net133));
 sg13g2_tiehi _6680__134 (.L_HI(net134));
 sg13g2_tiehi _6679__135 (.L_HI(net135));
 sg13g2_tiehi _6678__136 (.L_HI(net136));
 sg13g2_tiehi _6677__137 (.L_HI(net137));
 sg13g2_tiehi _6676__138 (.L_HI(net138));
 sg13g2_tiehi _6675__139 (.L_HI(net139));
 sg13g2_tiehi _6674__140 (.L_HI(net140));
 sg13g2_tiehi _6673__141 (.L_HI(net141));
 sg13g2_tiehi _6672__142 (.L_HI(net142));
 sg13g2_tiehi _6671__143 (.L_HI(net143));
 sg13g2_tiehi _6670__144 (.L_HI(net144));
 sg13g2_tiehi _6669__145 (.L_HI(net145));
 sg13g2_tiehi _6668__146 (.L_HI(net146));
 sg13g2_tiehi _6667__147 (.L_HI(net147));
 sg13g2_tiehi _6666__148 (.L_HI(net148));
 sg13g2_tiehi _6665__149 (.L_HI(net149));
 sg13g2_tiehi _6664__150 (.L_HI(net150));
 sg13g2_tiehi _6663__151 (.L_HI(net151));
 sg13g2_tiehi _6662__152 (.L_HI(net152));
 sg13g2_tiehi _6661__153 (.L_HI(net153));
 sg13g2_tiehi _6660__154 (.L_HI(net154));
 sg13g2_tiehi _6659__155 (.L_HI(net155));
 sg13g2_tiehi _6658__156 (.L_HI(net156));
 sg13g2_tiehi _6657__157 (.L_HI(net157));
 sg13g2_tiehi _6656__158 (.L_HI(net158));
 sg13g2_tiehi _6655__159 (.L_HI(net159));
 sg13g2_tiehi _6829__160 (.L_HI(net160));
 sg13g2_tiehi _6654__161 (.L_HI(net161));
 sg13g2_tiehi _6809__162 (.L_HI(net162));
 sg13g2_tiehi _6653__163 (.L_HI(net163));
 sg13g2_tiehi _6837__164 (.L_HI(net164));
 sg13g2_tiehi _6652__165 (.L_HI(net165));
 sg13g2_tiehi _6808__166 (.L_HI(net166));
 sg13g2_tiehi _6651__167 (.L_HI(net167));
 sg13g2_tiehi _6828__168 (.L_HI(net168));
 sg13g2_tiehi _6650__169 (.L_HI(net169));
 sg13g2_tiehi _6807__170 (.L_HI(net170));
 sg13g2_tiehi _6649__171 (.L_HI(net171));
 sg13g2_tiehi _6836__172 (.L_HI(net172));
 sg13g2_tiehi _6648__173 (.L_HI(net173));
 sg13g2_tiehi _6806__174 (.L_HI(net174));
 sg13g2_tiehi _6647__175 (.L_HI(net175));
 sg13g2_tiehi _6646__176 (.L_HI(net176));
 sg13g2_tiehi _6645__177 (.L_HI(net177));
 sg13g2_tiehi _6644__178 (.L_HI(net178));
 sg13g2_tiehi _6643__179 (.L_HI(net179));
 sg13g2_tiehi _6642__180 (.L_HI(net180));
 sg13g2_tiehi _6641__181 (.L_HI(net181));
 sg13g2_tiehi _6640__182 (.L_HI(net182));
 sg13g2_tiehi _6639__183 (.L_HI(net183));
 sg13g2_tiehi _6638__184 (.L_HI(net184));
 sg13g2_tiehi _6637__185 (.L_HI(net185));
 sg13g2_tiehi _6636__186 (.L_HI(net186));
 sg13g2_tiehi _6635__187 (.L_HI(net187));
 sg13g2_tiehi _6634__188 (.L_HI(net188));
 sg13g2_tiehi _6633__189 (.L_HI(net189));
 sg13g2_tiehi _6632__190 (.L_HI(net190));
 sg13g2_tiehi _6631__191 (.L_HI(net191));
 sg13g2_tiehi _6630__192 (.L_HI(net192));
 sg13g2_tiehi _6629__193 (.L_HI(net193));
 sg13g2_tiehi _6628__194 (.L_HI(net194));
 sg13g2_tiehi _6625__195 (.L_HI(net195));
 sg13g2_tiehi _6624__196 (.L_HI(net196));
 sg13g2_tiehi _6623__197 (.L_HI(net197));
 sg13g2_tiehi _6622__198 (.L_HI(net198));
 sg13g2_tiehi _6621__199 (.L_HI(net199));
 sg13g2_tiehi _6620__200 (.L_HI(net200));
 sg13g2_tiehi _6619__201 (.L_HI(net201));
 sg13g2_tiehi _6618__202 (.L_HI(net202));
 sg13g2_tiehi _6617__203 (.L_HI(net203));
 sg13g2_tiehi _6616__204 (.L_HI(net204));
 sg13g2_tiehi _6615__205 (.L_HI(net205));
 sg13g2_tiehi _6614__206 (.L_HI(net206));
 sg13g2_tiehi _6827__207 (.L_HI(net207));
 sg13g2_tiehi _6613__208 (.L_HI(net208));
 sg13g2_tiehi _6805__209 (.L_HI(net209));
 sg13g2_tiehi _6612__210 (.L_HI(net210));
 sg13g2_tiehi _6835__211 (.L_HI(net211));
 sg13g2_tiehi _6611__212 (.L_HI(net212));
 sg13g2_tiehi _6804__213 (.L_HI(net213));
 sg13g2_tiehi _6610__214 (.L_HI(net214));
 sg13g2_tiehi _6826__215 (.L_HI(net215));
 sg13g2_tiehi _6609__216 (.L_HI(net216));
 sg13g2_tiehi _6803__217 (.L_HI(net217));
 sg13g2_tiehi _6608__218 (.L_HI(net218));
 sg13g2_tiehi _6834__219 (.L_HI(net219));
 sg13g2_tiehi _6607__220 (.L_HI(net220));
 sg13g2_tiehi _6802__221 (.L_HI(net221));
 sg13g2_tiehi _6606__222 (.L_HI(net222));
 sg13g2_tiehi _6825__223 (.L_HI(net223));
 sg13g2_tiehi _6605__224 (.L_HI(net224));
 sg13g2_tiehi _6801__225 (.L_HI(net225));
 sg13g2_tiehi _6604__226 (.L_HI(net226));
 sg13g2_tiehi _6832__227 (.L_HI(net227));
 sg13g2_tiehi _6603__228 (.L_HI(net228));
 sg13g2_tiehi _6800__229 (.L_HI(net229));
 sg13g2_tiehi _6602__230 (.L_HI(net230));
 sg13g2_tiehi _6601__231 (.L_HI(net231));
 sg13g2_tiehi _6600__232 (.L_HI(net232));
 sg13g2_tiehi _6599__233 (.L_HI(net233));
 sg13g2_tiehi _6598__234 (.L_HI(net234));
 sg13g2_tiehi _6597__235 (.L_HI(net235));
 sg13g2_tiehi _6596__236 (.L_HI(net236));
 sg13g2_tiehi _6595__237 (.L_HI(net237));
 sg13g2_tiehi _6594__238 (.L_HI(net238));
 sg13g2_tiehi _6593__239 (.L_HI(net239));
 sg13g2_tiehi _6592__240 (.L_HI(net240));
 sg13g2_tiehi _6591__241 (.L_HI(net241));
 sg13g2_tiehi _6590__242 (.L_HI(net242));
 sg13g2_tiehi _6589__243 (.L_HI(net243));
 sg13g2_tiehi _6588__244 (.L_HI(net244));
 sg13g2_tiehi _6627__245 (.L_HI(net245));
 sg13g2_tiehi _6587__246 (.L_HI(net246));
 sg13g2_tiehi _6586__247 (.L_HI(net247));
 sg13g2_tiehi _6585__248 (.L_HI(net248));
 sg13g2_tiehi _6783__249 (.L_HI(net249));
 sg13g2_tiehi _6787__250 (.L_HI(net250));
 sg13g2_tiehi _6584__251 (.L_HI(net251));
 sg13g2_tiehi _6583__252 (.L_HI(net252));
 sg13g2_tiehi _6582__253 (.L_HI(net253));
 sg13g2_tiehi _6581__254 (.L_HI(net254));
 sg13g2_tiehi _6580__255 (.L_HI(net255));
 sg13g2_tiehi _6579__256 (.L_HI(net256));
 sg13g2_tiehi _6578__257 (.L_HI(net257));
 sg13g2_tiehi _6577__258 (.L_HI(net258));
 sg13g2_tiehi _6576__259 (.L_HI(net259));
 sg13g2_tiehi _6824__260 (.L_HI(net260));
 sg13g2_tiehi _6575__261 (.L_HI(net261));
 sg13g2_tiehi _6799__262 (.L_HI(net262));
 sg13g2_tiehi _6574__263 (.L_HI(net263));
 sg13g2_tiehi _6573__264 (.L_HI(net264));
 sg13g2_tiehi _6572__265 (.L_HI(net265));
 sg13g2_tiehi _6571__266 (.L_HI(net266));
 sg13g2_tiehi _6570__267 (.L_HI(net267));
 sg13g2_tiehi _6833__268 (.L_HI(net268));
 sg13g2_tiehi _6569__269 (.L_HI(net269));
 sg13g2_tiehi _6798__270 (.L_HI(net270));
 sg13g2_tiehi _6568__271 (.L_HI(net271));
 sg13g2_tiehi _6823__272 (.L_HI(net272));
 sg13g2_tiehi _6567__273 (.L_HI(net273));
 sg13g2_tiehi _6797__274 (.L_HI(net274));
 sg13g2_tiehi _6566__275 (.L_HI(net275));
 sg13g2_tiehi _6839__276 (.L_HI(net276));
 sg13g2_tiehi _6565__277 (.L_HI(net277));
 sg13g2_tiehi _6564__278 (.L_HI(net278));
 sg13g2_tiehi _6563__279 (.L_HI(net279));
 sg13g2_tiehi _6562__280 (.L_HI(net280));
 sg13g2_tiehi _6561__281 (.L_HI(net281));
 sg13g2_tiehi _6560__282 (.L_HI(net282));
 sg13g2_tiehi _6559__283 (.L_HI(net283));
 sg13g2_tiehi _6558__284 (.L_HI(net284));
 sg13g2_tiehi _6557__285 (.L_HI(net285));
 sg13g2_tiehi _6796__286 (.L_HI(net286));
 sg13g2_tiehi _6822__287 (.L_HI(net287));
 sg13g2_tiehi _6795__288 (.L_HI(net288));
 sg13g2_tiehi _6830__289 (.L_HI(net289));
 sg13g2_tiehi _6794__290 (.L_HI(net290));
 sg13g2_tiehi _6821__291 (.L_HI(net291));
 sg13g2_tiehi _6793__292 (.L_HI(net292));
 sg13g2_tiehi _6788__293 (.L_HI(net293));
 sg13g2_tiehi _6831__294 (.L_HI(net294));
 sg13g2_tiehi _6820__295 (.L_HI(net295));
 sg13g2_tiehi _6792__296 (.L_HI(net296));
 sg13g2_tiehi _6819__297 (.L_HI(net297));
 sg13g2_tiehi _6791__298 (.L_HI(net298));
 sg13g2_tiehi _6818__299 (.L_HI(net299));
 sg13g2_tiehi _6790__300 (.L_HI(net300));
 sg13g2_tiehi tt_um_toivoh_demo_tt10_301 (.L_HI(net301));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_toivoh_demo_tt10_4 (.L_LO(net4));
 sg13g2_tielo tt_um_toivoh_demo_tt10_5 (.L_LO(net5));
 sg13g2_tielo tt_um_toivoh_demo_tt10_6 (.L_LO(net6));
 sg13g2_tielo tt_um_toivoh_demo_tt10_7 (.L_LO(net7));
 sg13g2_tielo tt_um_toivoh_demo_tt10_8 (.L_LO(net8));
 sg13g2_tielo tt_um_toivoh_demo_tt10_9 (.L_LO(net9));
 sg13g2_tielo tt_um_toivoh_demo_tt10_10 (.L_LO(net10));
 sg13g2_tielo tt_um_toivoh_demo_tt10_11 (.L_LO(net11));
 sg13g2_tielo tt_um_toivoh_demo_tt10_12 (.L_LO(net12));
 sg13g2_tielo tt_um_toivoh_demo_tt10_13 (.L_LO(net13));
 sg13g2_tielo tt_um_toivoh_demo_tt10_14 (.L_LO(net14));
 sg13g2_tielo tt_um_toivoh_demo_tt10_15 (.L_LO(net15));
 sg13g2_tielo tt_um_toivoh_demo_tt10_16 (.L_LO(net16));
 sg13g2_tiehi _6789__17 (.L_HI(net17));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(_2107_));
 sg13g2_buf_2 fanout848 (.A(_2100_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_2098_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_2099_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_0810_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_0808_),
    .X(net853));
 sg13g2_buf_4 fanout854 (.X(net854),
    .A(net855));
 sg13g2_buf_4 fanout855 (.X(net855),
    .A(_0751_));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(_0740_));
 sg13g2_buf_2 fanout857 (.A(_0740_),
    .X(net857));
 sg13g2_buf_4 fanout858 (.X(net858),
    .A(_0731_));
 sg13g2_buf_2 fanout859 (.A(net861),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(net861),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_2690_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(net863),
    .X(net862));
 sg13g2_buf_1 fanout863 (.A(net864),
    .X(net863));
 sg13g2_buf_1 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_1 fanout865 (.A(_2676_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(net867),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net868),
    .X(net867));
 sg13g2_buf_4 fanout868 (.X(net868),
    .A(_1721_));
 sg13g2_buf_2 fanout869 (.A(_1915_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(net872),
    .X(net870));
 sg13g2_buf_1 fanout871 (.A(net872),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_2703_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_2047_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_1 fanout875 (.A(_2046_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_2044_),
    .X(net876));
 sg13g2_buf_4 fanout877 (.X(net877),
    .A(_1676_));
 sg13g2_buf_4 fanout878 (.X(net878),
    .A(net879));
 sg13g2_buf_4 fanout879 (.X(net879),
    .A(_0458_));
 sg13g2_buf_2 fanout880 (.A(_2049_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(net882),
    .X(net881));
 sg13g2_buf_1 fanout882 (.A(_2028_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(net885),
    .X(net883));
 sg13g2_buf_4 fanout884 (.X(net884),
    .A(net885));
 sg13g2_buf_4 fanout885 (.X(net885),
    .A(_2539_));
 sg13g2_buf_4 fanout886 (.X(net886),
    .A(_0596_));
 sg13g2_buf_2 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_4 fanout888 (.X(net888),
    .A(_0593_));
 sg13g2_buf_4 fanout889 (.X(net889),
    .A(_0578_));
 sg13g2_buf_2 fanout890 (.A(_0578_),
    .X(net890));
 sg13g2_buf_4 fanout891 (.X(net891),
    .A(net892));
 sg13g2_buf_2 fanout892 (.A(_0575_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(net894),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_0575_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_0474_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_0474_),
    .X(net896));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(net900));
 sg13g2_buf_2 fanout898 (.A(net900),
    .X(net898));
 sg13g2_buf_4 fanout899 (.X(net899),
    .A(net900));
 sg13g2_buf_2 fanout900 (.A(_2526_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(net902),
    .X(net901));
 sg13g2_buf_1 fanout902 (.A(net903),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(_2498_),
    .X(net903));
 sg13g2_buf_4 fanout904 (.X(net904),
    .A(_1028_));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(_0697_));
 sg13g2_buf_2 fanout906 (.A(net907),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(net908),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_0473_),
    .X(net908));
 sg13g2_buf_4 fanout909 (.X(net909),
    .A(_0465_));
 sg13g2_buf_2 fanout910 (.A(net911),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(net912),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_0462_),
    .X(net912));
 sg13g2_buf_4 fanout913 (.X(net913),
    .A(net914));
 sg13g2_buf_2 fanout914 (.A(_2994_),
    .X(net914));
 sg13g2_buf_4 fanout915 (.X(net915),
    .A(net916));
 sg13g2_buf_2 fanout916 (.A(net917),
    .X(net916));
 sg13g2_buf_4 fanout917 (.X(net917),
    .A(_2549_));
 sg13g2_buf_4 fanout918 (.X(net918),
    .A(net920));
 sg13g2_buf_2 fanout919 (.A(net920),
    .X(net919));
 sg13g2_buf_4 fanout920 (.X(net920),
    .A(_2535_));
 sg13g2_buf_4 fanout921 (.X(net921),
    .A(net922));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(_0540_));
 sg13g2_buf_2 fanout923 (.A(_0540_),
    .X(net923));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(net925));
 sg13g2_buf_4 fanout925 (.X(net925),
    .A(_0529_));
 sg13g2_buf_4 fanout926 (.X(net926),
    .A(net927));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(_0527_));
 sg13g2_buf_2 fanout928 (.A(net929),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_2973_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_2973_),
    .X(net930));
 sg13g2_buf_1 fanout931 (.A(_2973_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(net933),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(net934),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_2972_),
    .X(net934));
 sg13g2_buf_1 fanout935 (.A(_2972_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_2563_),
    .X(net936));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(_1680_));
 sg13g2_buf_4 fanout938 (.X(net938),
    .A(_1669_));
 sg13g2_buf_2 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_1 fanout940 (.A(_1507_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(net942),
    .X(net941));
 sg13g2_buf_4 fanout942 (.X(net942),
    .A(_1665_));
 sg13g2_buf_4 fanout943 (.X(net943),
    .A(_1654_));
 sg13g2_buf_2 fanout944 (.A(net945),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_1504_),
    .X(net945));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(_1504_));
 sg13g2_buf_4 fanout947 (.X(net947),
    .A(_1150_));
 sg13g2_buf_2 fanout948 (.A(_1031_),
    .X(net948));
 sg13g2_buf_4 fanout949 (.X(net949),
    .A(net950));
 sg13g2_buf_2 fanout950 (.A(_1668_),
    .X(net950));
 sg13g2_buf_4 fanout951 (.X(net951),
    .A(_1503_));
 sg13g2_buf_2 fanout952 (.A(_1503_),
    .X(net952));
 sg13g2_buf_4 fanout953 (.X(net953),
    .A(net955));
 sg13g2_buf_2 fanout954 (.A(net955),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(net956),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(net958),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(net958),
    .X(net957));
 sg13g2_buf_4 fanout958 (.X(net958),
    .A(_2970_));
 sg13g2_buf_2 fanout959 (.A(net960),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(net961),
    .X(net960));
 sg13g2_buf_1 fanout961 (.A(_2476_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_2476_),
    .X(net962));
 sg13g2_buf_1 fanout963 (.A(_2476_),
    .X(net963));
 sg13g2_buf_4 fanout964 (.X(net964),
    .A(_1502_));
 sg13g2_buf_2 fanout965 (.A(_1678_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(net967),
    .X(net966));
 sg13g2_buf_4 fanout967 (.X(net967),
    .A(_3066_));
 sg13g2_buf_2 fanout968 (.A(net969),
    .X(net968));
 sg13g2_buf_1 fanout969 (.A(_3065_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(net971),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_3065_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(net975),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(net975),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(net975),
    .X(net974));
 sg13g2_buf_1 fanout975 (.A(_1544_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(net977),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(net978),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_1543_),
    .X(net978));
 sg13g2_buf_4 fanout979 (.X(net979),
    .A(_1149_));
 sg13g2_buf_2 fanout980 (.A(_1724_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_1723_),
    .X(net981));
 sg13g2_buf_4 fanout982 (.X(net982),
    .A(_1672_));
 sg13g2_buf_2 fanout983 (.A(_1672_),
    .X(net983));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(_1671_));
 sg13g2_buf_2 fanout985 (.A(net986),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_1485_),
    .X(net986));
 sg13g2_buf_4 fanout987 (.X(net987),
    .A(net989));
 sg13g2_buf_2 fanout988 (.A(net989),
    .X(net988));
 sg13g2_buf_4 fanout989 (.X(net989),
    .A(_1484_));
 sg13g2_buf_2 fanout990 (.A(_3081_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(net992),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_3048_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(net996),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(net995),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(net996),
    .X(net995));
 sg13g2_buf_1 fanout996 (.A(_3040_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(net1000),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(net999),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(net1000),
    .X(net999));
 sg13g2_buf_1 fanout1000 (.A(_3035_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_2625_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_2625_),
    .X(net1002));
 sg13g2_buf_4 fanout1003 (.X(net1003),
    .A(_1410_));
 sg13g2_buf_4 fanout1004 (.X(net1004),
    .A(_2864_));
 sg13g2_buf_2 fanout1005 (.A(_2864_),
    .X(net1005));
 sg13g2_buf_4 fanout1006 (.X(net1006),
    .A(_2863_));
 sg13g2_buf_4 fanout1007 (.X(net1007),
    .A(_2862_));
 sg13g2_buf_4 fanout1008 (.X(net1008),
    .A(_2861_));
 sg13g2_buf_4 fanout1009 (.X(net1009),
    .A(_2858_));
 sg13g2_buf_2 fanout1010 (.A(net1011),
    .X(net1010));
 sg13g2_buf_1 fanout1011 (.A(_2857_),
    .X(net1011));
 sg13g2_buf_4 fanout1012 (.X(net1012),
    .A(_2852_));
 sg13g2_buf_2 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_4 fanout1014 (.X(net1014),
    .A(_2848_));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(_2847_));
 sg13g2_buf_2 fanout1016 (.A(_2847_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_2845_),
    .X(net1017));
 sg13g2_buf_4 fanout1018 (.X(net1018),
    .A(_2844_));
 sg13g2_buf_2 fanout1019 (.A(net1020),
    .X(net1019));
 sg13g2_buf_1 fanout1020 (.A(_2833_),
    .X(net1020));
 sg13g2_buf_4 fanout1021 (.X(net1021),
    .A(_2832_));
 sg13g2_buf_4 fanout1022 (.X(net1022),
    .A(net1023));
 sg13g2_buf_2 fanout1023 (.A(net1024),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_2831_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(\dtop.field_top.player.chan_timer[5] ),
    .X(net1025));
 sg13g2_buf_1 fanout1026 (.A(net1027),
    .X(net1026));
 sg13g2_buf_4 fanout1027 (.X(net1027),
    .A(\dtop.field_top.player.chan_timer[5] ));
 sg13g2_buf_4 fanout1028 (.X(net1028),
    .A(net327));
 sg13g2_buf_2 fanout1029 (.A(\dtop.field_top.player.osc0[22] ),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(net674),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(\dtop.field_top.controller.pattern0[1] ),
    .X(net1031));
 sg13g2_buf_4 fanout1032 (.X(net1032),
    .A(net688));
 sg13g2_buf_4 fanout1033 (.X(net1033),
    .A(\dtop.field_top.controller.ppos[5] ));
 sg13g2_buf_4 fanout1034 (.X(net1034),
    .A(_0107_));
 sg13g2_buf_2 fanout1035 (.A(net1036),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(\dtop.field_top.afl_pc[8] ),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(net1039),
    .X(net1037));
 sg13g2_buf_1 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(\dtop.field_top.afl_pc[7] ),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(net1041),
    .X(net1040));
 sg13g2_buf_4 fanout1041 (.X(net1041),
    .A(\dtop.field_top.afl_pc[6] ));
 sg13g2_buf_2 fanout1042 (.A(net1044),
    .X(net1042));
 sg13g2_buf_4 fanout1043 (.X(net1043),
    .A(net1044));
 sg13g2_buf_4 fanout1044 (.X(net1044),
    .A(\dtop.field_top.afl_pc[5] ));
 sg13g2_buf_4 fanout1045 (.X(net1045),
    .A(net1046));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(\dtop.field_top.afl_pc[4] ));
 sg13g2_buf_4 fanout1047 (.X(net1047),
    .A(net1048));
 sg13g2_buf_4 fanout1048 (.X(net1048),
    .A(net1049));
 sg13g2_buf_2 fanout1049 (.A(\dtop.field_top.afl_pc[3] ),
    .X(net1049));
 sg13g2_buf_4 fanout1050 (.X(net1050),
    .A(\dtop.field_top.afl_pc[2] ));
 sg13g2_buf_2 fanout1051 (.A(\dtop.field_top.afl_pc[2] ),
    .X(net1051));
 sg13g2_buf_4 fanout1052 (.X(net1052),
    .A(net1053));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(net1054));
 sg13g2_buf_4 fanout1054 (.X(net1054),
    .A(\dtop.field_top.afl_pc[1] ));
 sg13g2_buf_4 fanout1055 (.X(net1055),
    .A(net1056));
 sg13g2_buf_4 fanout1056 (.X(net1056),
    .A(net1057));
 sg13g2_buf_4 fanout1057 (.X(net1057),
    .A(\dtop.field_top.afl_pc[0] ));
 sg13g2_buf_4 fanout1058 (.X(net1058),
    .A(\dtop.field_top.afl_sub_pc[0] ));
 sg13g2_buf_1 fanout1059 (.A(\dtop.field_top.afl_sub_pc[0] ),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(\dtop.field_top.alt_osc[8] ),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(\dtop.field_top.player.osc0[20] ),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(net1063),
    .X(net1062));
 sg13g2_buf_4 fanout1063 (.X(net1063),
    .A(net1064));
 sg13g2_buf_2 fanout1064 (.A(\dtop.field_top.player.osc0[19] ),
    .X(net1064));
 sg13g2_buf_4 fanout1065 (.X(net1065),
    .A(net695));
 sg13g2_buf_4 fanout1066 (.X(net1066),
    .A(net1067));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(net1069));
 sg13g2_buf_2 fanout1068 (.A(net1069),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(net698),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(\dtop.field_top.player.controller.ppos[4] ),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(net1074),
    .X(net1071));
 sg13g2_buf_1 fanout1072 (.A(net1074),
    .X(net1072));
 sg13g2_buf_4 fanout1073 (.X(net1073),
    .A(net1074));
 sg13g2_buf_2 fanout1074 (.A(net1075),
    .X(net1074));
 sg13g2_buf_4 fanout1075 (.X(net1075),
    .A(net702));
 sg13g2_buf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(net1078),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(\dtop.field_top.player.controller.ppos[3] ),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(net1082),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(net1082),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(net1082),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(net1083),
    .X(net1082));
 sg13g2_buf_4 fanout1083 (.X(net1083),
    .A(net685));
 sg13g2_buf_2 fanout1084 (.A(net1086),
    .X(net1084));
 sg13g2_buf_1 fanout1085 (.A(net1086),
    .X(net1085));
 sg13g2_buf_1 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(net1088),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(\dtop.field_top.player.osc0[15] ),
    .X(net1088));
 sg13g2_buf_4 fanout1089 (.X(net1089),
    .A(net1090));
 sg13g2_buf_2 fanout1090 (.A(net1091),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(net1092),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(net682),
    .X(net1092));
 sg13g2_buf_4 fanout1093 (.X(net1093),
    .A(\dtop.field_top.player.osc0[13] ));
 sg13g2_buf_2 fanout1094 (.A(net705),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(net1096),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(net1097),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(net1098),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(net669),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(net1101),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(net1101),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(net1102),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(net691),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(net1104),
    .X(net1103));
 sg13g2_buf_4 fanout1104 (.X(net1104),
    .A(\dtop.field_top.player.chan_timer[2] ));
 sg13g2_buf_4 fanout1105 (.X(net1105),
    .A(net1106));
 sg13g2_buf_2 fanout1106 (.A(\dtop.field_top.player.chan_timer[1] ),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_4 fanout1108 (.X(net1108),
    .A(\dtop.field_top.player.chan_timer[0] ));
 sg13g2_buf_2 fanout1109 (.A(\dtop.field_top.channel[1] ),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(net1113),
    .X(net1110));
 sg13g2_buf_1 fanout1111 (.A(net1113),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(_2160_),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(net1115),
    .X(net1114));
 sg13g2_buf_4 fanout1115 (.X(net1115),
    .A(_2842_));
 sg13g2_buf_2 fanout1116 (.A(net1117),
    .X(net1116));
 sg13g2_buf_4 fanout1117 (.X(net1117),
    .A(rst_n));
 sg13g2_buf_2 fanout1118 (.A(net1119),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(net1120),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(net1121),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(rst_n),
    .X(net1121));
 sg13g2_buf_2 input1 (.A(ui_in[6]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[7]),
    .X(net2));
 sg13g2_tielo tt_um_toivoh_demo_tt10_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_5_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_25_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_26_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_6_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_7_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_13_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_22_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_32_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_21_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\dtop.field_top.prev_wave[4] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0185_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0116_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0076_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold5 (.A(_1130_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0078_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold7 (.A(_1144_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0145_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold9 (.A(\dtop.field_top.reg1[15] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0230_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold11 (.A(\dtop.field_top.prev_wave[7] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0188_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0077_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold14 (.A(_1142_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0144_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold16 (.A(\dtop.field_top.player.sched.alu.p1 ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold17 (.A(\dtop.field_top.nsource.num_iter[0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0390_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold19 (.A(\dtop.field_top.nsource.shuffle_state.in[4] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0316_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0062_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold22 (.A(_1133_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0140_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold24 (.A(\dtop.field_top.nsource.shuffle_state.in[3] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0315_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold26 (.A(\dtop.field_top.channel_output[10] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0214_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold28 (.A(\dtop.field_top.comp_value0_1[1] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0216_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold30 (.A(\dtop.field_top.prev_wave[1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0182_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold32 (.A(\dtop.field_top.wave[0] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0207_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold34 (.A(\dtop.field_top.nsource.shuffle_state.in[7] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0319_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold36 (.A(\dtop.field_top.reg3[15] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0264_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold38 (.A(\dtop.field_top.nsource.shuffle_state.in[2] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0314_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0083_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold41 (.A(\dtop.field_top.wave[6] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0213_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold43 (.A(\dtop.field_top.nsource.shuffle_state.in[6] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0318_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold45 (.A(\dtop.field_top.nsource.shuffle_state.in[0] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0312_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold47 (.A(\dtop.field_top.reg4[15] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0281_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold49 (.A(\dtop.field_top.fy[8] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold50 (.A(_1146_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0146_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0061_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold53 (.A(_1136_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold54 (.A(\dtop.field_top.fx[10] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold55 (.A(\dtop.field_top.comp_values0[3][1] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0250_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold57 (.A(\dtop.field_top.nsource.num_iter[1] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold58 (.A(\dtop.field_top.nsource.shuffle_state.in[5] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold59 (.A(\dtop.field_top.comp_value0_1[2] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0217_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold61 (.A(\dtop.field_top.fy[4] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold62 (.A(_1138_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0142_),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold64 (.A(\dtop.field_top.prev_wave[0] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0181_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold66 (.A(\dtop.field_top.comp_value0[0] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0197_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold68 (.A(\dtop.field_top.fx[9] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold69 (.A(_1160_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0156_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold71 (.A(\dtop.field_top.logo_prev_pixel ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0176_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold73 (.A(\dtop.field_top.player.osc0[2] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold74 (.A(\dtop.field_top.wave[1] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0208_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold76 (.A(\dtop.field_top.fx[7] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0154_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold78 (.A(\dtop.field_top.fx[5] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold79 (.A(_1156_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0152_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold81 (.A(\dtop.field_top.reg1[12] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0227_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold83 (.A(\dtop.field_top.player.out_pw[0] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold84 (.A(_2980_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold85 (.A(\dtop.field_top.wave[7] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold86 (.A(\dtop.field_top.reg1[14] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0229_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold88 (.A(\dtop.field_top.wave[4] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold89 (.A(\dtop.field_top.comp_value0_1[0] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0215_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold91 (.A(\dtop.field_top.reg1[11] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0226_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold93 (.A(\dtop.field_top.reg1[16] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0231_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold95 (.A(\dtop.field_top.comp_value0[7] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0204_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold97 (.A(\dtop.field_top.fy[10] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0137_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold99 (.A(\dtop.field_top.prev_wave[3] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0192_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold101 (.A(\dtop.field_top.afl_alu.p ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold102 (.A(\dtop.field_top.last_wave[3] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold103 (.A(\dtop.field_top.prev_wave[6] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold104 (.A(\dtop.field_top.comp_value0[6] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0203_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold106 (.A(\dtop.field_top.fx[6] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold107 (.A(_1157_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0153_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold109 (.A(\dtop.field_top.reg1[13] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0228_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold111 (.A(\dtop.field_top.fy[5] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold112 (.A(_1140_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0143_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold114 (.A(\dtop.field_top.nsource.shuffle_state.in[1] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold115 (.A(\dtop.field_top.prev_wave[5] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0194_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold117 (.A(\dtop.field_top.prev_wave[2] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0191_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold119 (.A(\dtop.field_top.comp_value0_1[4] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0219_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold121 (.A(\dtop.field_top.last_wave[2] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold122 (.A(\dtop.field_top.player.controller.pattern0[1] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0342_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold124 (.A(\dtop.field_top.player.osc0[22] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold125 (.A(\dtop.field_top.comp_value0_1[5] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0220_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold127 (.A(\dtop.field_top.player.osc0[4] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold128 (.A(\dtop.field_top.comp_values0[3][2] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0251_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold130 (.A(\dtop.field_top.player.osc0[3] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold131 (.A(\dtop.field_top.comp_value0[3] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0200_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold133 (.A(\dtop.field_top.controller.timer[0] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0331_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold135 (.A(\dtop.field_top.comp_value0_1[7] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0222_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold137 (.A(\dtop.field_top.wave[5] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0212_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold139 (.A(\dtop.field_top.player.sched.alu.p0 ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold140 (.A(\dtop.field_top.comp_value0[2] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0199_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold142 (.A(\dtop.field_top.reg3[12] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0261_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold144 (.A(\dtop.field_top.reg3[13] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0262_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold146 (.A(\dtop.field_top.reg4[13] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0279_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold148 (.A(\dtop.field_top.reg2[14] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0246_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold150 (.A(\dtop.field_top.fy[9] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0136_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold152 (.A(\dtop.field_top.reg2[12] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0244_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold154 (.A(\dtop.field_top.reg4[16] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0282_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold156 (.A(\dtop.field_top.comp_values0[2][0] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0232_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold158 (.A(\dtop.field_top.comp_value0_1[3] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0218_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold160 (.A(\dtop.field_top.reg2[13] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0245_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold162 (.A(\dtop.field_top.fx[1] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold163 (.A(_1152_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold164 (.A(\dtop.field_top.reg4[12] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0278_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold166 (.A(\dtop.field_top.reg3[16] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0265_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold168 (.A(\dtop.field_top.reg4[11] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0277_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold170 (.A(\dtop.field_top.controller.timer[2] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0333_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold172 (.A(\dtop.field_top.comp_value0_1[6] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0221_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold174 (.A(\dtop.field_top.reg3[11] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0260_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold176 (.A(\dtop.field_top.controller.timer[1] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0332_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold178 (.A(\dtop.field_top.comp_values0[3][0] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0249_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold180 (.A(\dtop.field_top.last_wave[6] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold181 (.A(\dtop.field_top.player.osc0[7] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold182 (.A(\dtop.field_top.player.osc0[5] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold183 (.A(\dtop.field_top.fx[4] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold184 (.A(_1155_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0151_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold186 (.A(\dtop.field_top.fx[0] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold187 (.A(\dtop.field_top.player.osc0[8] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold188 (.A(\dtop.field_top.comp_values0[4][1] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0267_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold190 (.A(\dtop.field_top.reg2[11] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0243_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold192 (.A(\dtop.field_top.comp_values0[3][7] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0256_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold194 (.A(\dtop.field_top.comp_value0_1[8] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0223_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold196 (.A(\dtop.field_top.fx[3] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold197 (.A(_1154_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold198 (.A(\dtop.field_top.comp_values0[2][2] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0234_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold200 (.A(\dtop.field_top.comp_values0[3][6] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0255_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold202 (.A(\dtop.field_top.comp_value0_1[10] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0225_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold204 (.A(\dtop.field_top.reg2[15] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0247_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold206 (.A(\dtop.field_top.comp_values0[4][9] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0275_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold208 (.A(\dtop.field_top.player.osc0[20] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold209 (.A(\dtop.field_top.player.osc0[9] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold210 (.A(\dtop.field_top.fx[8] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold211 (.A(_1159_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0155_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold213 (.A(\dtop.field_top.comp_values0[3][4] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0253_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold215 (.A(\dtop.field_top.reg3[14] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0263_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold217 (.A(\dtop.field_top.comp_values0[4][0] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0266_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold219 (.A(\dtop.field_top.player.out_acc[8] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0376_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold221 (.A(\dtop.field_top.player.out_acc[3] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0371_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold223 (.A(\dtop.field_top.comp_values0[4][2] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0268_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold225 (.A(\dtop.field_top.player.out_acc[9] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0377_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold227 (.A(\dtop.field_top.comp_values0[4][4] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0270_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold229 (.A(\dtop.field_top.comp_values0[3][3] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0252_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0017_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold232 (.A(\dtop.field_top.comp_value0[5] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0202_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold234 (.A(\dtop.field_top.reg2[16] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0248_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold236 (.A(\dtop.field_top.wave[2] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0209_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold238 (.A(\dtop.field_top.comp_values0[3][5] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0254_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold240 (.A(\dtop.field_top.comp_value0[1] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0198_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold242 (.A(\dtop.field_top.comp_values0[2][1] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0233_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold244 (.A(\dtop.field_top.comp_value0[4] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0201_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold246 (.A(\dtop.field_top.reg4[14] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0280_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold248 (.A(\dtop.field_top.player.out_acc[5] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0373_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold250 (.A(\dtop.field_top.comp_values0[2][4] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0236_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold252 (.A(\dtop.field_top.acc[12] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold253 (.A(\dtop.field_top.comp_values0[3][8] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0257_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold255 (.A(\dtop.field_top.comp_value0_0[10] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0206_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold257 (.A(\dtop.field_top.comp_value0_1[9] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0224_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold259 (.A(\dtop.field_top.lside ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0283_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold261 (.A(\dtop.field_top.comp_value0[8] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0205_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold263 (.A(\dtop.field_top.player.out_acc[4] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0372_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold265 (.A(\dtop.field_top.player.osc0[6] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold266 (.A(\dtop.field_top.comp_values0[4][3] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0269_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold268 (.A(\dtop.field_top.last_wave[5] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0075_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold270 (.A(_1126_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold271 (.A(\dtop.field_top.player.osc0[0] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold272 (.A(\dtop.field_top.comp_values0[3][10] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0259_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold274 (.A(\dtop.field_top.player.out_acc[7] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0375_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold276 (.A(\dtop.field_top.comp_values0[2][10] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0242_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold278 (.A(\dtop.field_top.player.osc0[1] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold279 (.A(\dtop.field_top.player.out_acc[0] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0368_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold281 (.A(\dtop.field_top.player.out_acc[2] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0370_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold283 (.A(\dtop.field_top.rside ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0284_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold285 (.A(\dtop.field_top.channel_output[7] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold286 (.A(\dtop.field_top.player.controller.pattern0[0] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0341_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold288 (.A(\dtop.field_top.comp_values0[4][5] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0271_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold290 (.A(\dtop.field_top.alt_osc[4] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0293_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold292 (.A(\dtop.field_top.comp_values0[2][3] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0235_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold294 (.A(\dtop.field_top.comp_values0[4][8] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0274_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold296 (.A(\dtop.field_top.comp_values0[2][6] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0238_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0018_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold299 (.A(_2621_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold300 (.A(\dtop.field_top.rs.scan_y.pos[9] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold301 (.A(\dtop.field_top.rs.scan_x.state[1] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold302 (.A(\dtop.field_top.player.out_acc[1] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0369_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold304 (.A(\dtop.field_top.comp_values0[2][7] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold305 (.A(\dtop.field_top.comp_values0[2][8] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0240_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold307 (.A(\dtop.field_top.comp_values0[4][10] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0276_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold309 (.A(\dtop.field_top.player.out_acc[6] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold310 (.A(\dtop.field_top.comp_values0[4][7] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold311 (.A(\dtop.field_top.player.osc0[11] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold312 (.A(\dtop.field_top.fx[2] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold313 (.A(_1153_),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0149_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold315 (.A(\dtop.field_top.wave[3] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0210_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold317 (.A(\dtop.field_top.afl_alu.last_r_sum_msbs[0] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0069_),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold319 (.A(_2572_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold320 (.A(\dtop.field_top.player.osc0[10] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold321 (.A(\dtop.field_top.masked_bits[0] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold322 (.A(\dtop.field_top.comp_values0[2][5] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0237_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold324 (.A(\dtop.field_top.comp_values0[3][9] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0258_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold326 (.A(\dtop.field_top.controller.ppos[2] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold327 (.A(\dtop.field_top.player.out_pw[6] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold328 (.A(\dtop.field_top.rs.scan_x.state[0] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold329 (.A(_2929_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold330 (.A(\dtop.field_top.comp_values0[4][6] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0272_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold332 (.A(\dtop.field_top.channel[0] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold333 (.A(_3013_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold334 (.A(\dtop.field_top.channel[2] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold335 (.A(_3014_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold336 (.A(\dtop.field_top.channel_output[0] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold337 (.A(\dtop.field_top.acc[13] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold338 (.A(\dtop.field_top.rs.scan_y.state[1] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold339 (.A(_2992_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0119_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold341 (.A(\dtop.field_top.acc[16] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold342 (.A(\dtop.field_top.afl_alu.last_r_sum_msbs[1] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold343 (.A(\dtop.field_top.controller.ppos[1] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0335_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold345 (.A(\dtop.field_top.comp_values0[2][9] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0241_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0008_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold348 (.A(\dtop.field_top.player.controller.ppos[0] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0334_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold350 (.A(\dtop.field_top.acc[15] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold351 (.A(\dtop.field_top.channel_output[9] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold352 (.A(\dtop.field_top.controller.ppos[4] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold353 (.A(\dtop.field_top.player.osc0[12] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold354 (.A(\dtop.field_top.acc[11] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold355 (.A(\dtop.field_top.channel_output[1] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold356 (.A(\dtop.field_top.channel_output[3] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold357 (.A(\dtop.field_top.acc[14] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0067_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0021_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold360 (.A(\dtop.field_top.channel_output[2] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold361 (.A(\dtop.field_top.masked_bits[1] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0117_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold363 (.A(\dtop.field_top.channel_output[8] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0020_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0015_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold366 (.A(_2577_),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold367 (.A(\dtop.field_top.acc[10] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold368 (.A(\dtop.field_top.player.chan_timer[4] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold369 (.A(_3025_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold370 (.A(\dtop.field_top.acc[8] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold371 (.A(\dtop.field_top.rs.scan_y.pos[8] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold372 (.A(\dtop.field_top.acc[4] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold373 (.A(\dtop.field_top.controller.pattern0[2] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0343_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold375 (.A(\dtop.field_top.alt_osc[3] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold376 (.A(_2567_),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold377 (.A(\dtop.field_top.controller.ppos[3] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold378 (.A(\dtop.field_top.acc[0] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold379 (.A(_2644_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold380 (.A(\dtop.field_top.acc[3] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold381 (.A(\dtop.field_top.player.osc0[14] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0010_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold383 (.A(_2565_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold384 (.A(\dtop.field_top.player.osc0[16] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold385 (.A(\dtop.field_top.afl_sub_pc[1] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0302_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold387 (.A(\dtop.field_top.controller.ppos[6] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0340_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold389 (.A(\dtop.field_top.player.osc0[21] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold390 (.A(\dtop.field_top.player.chan_timer[3] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold391 (.A(\dtop.field_top.rs.scan_x.state[0] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold392 (.A(\dtop.field_top.alt_osc[1] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold393 (.A(\dtop.field_top.channel_output[6] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold394 (.A(\dtop.field_top.player.controller.ppos[5] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold395 (.A(\dtop.field_top.sflag ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold396 (.A(\dtop.field_top.acc[5] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold397 (.A(\dtop.field_top.player.osc0[18] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold398 (.A(\dtop.field_top.rs.scan_y.state[0] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold399 (.A(\dtop.field_top.acc[9] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold400 (.A(\dtop.field_top.sflag2 ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold401 (.A(\dtop.field_top.player.osc0[17] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold402 (.A(\dtop.field_top.acc[6] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold403 (.A(\dtop.field_top.channel_output[4] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold404 (.A(\dtop.field_top.player.osc0[13] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold405 (.A(\dtop.field_top.channel_output[5] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold406 (.A(\dtop.field_top.alt_osc[7] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold407 (.A(\dtop.field_top.acc[1] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold408 (.A(\dtop.field_top.acc[7] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0110_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold410 (.A(\dtop.field_top.acc[2] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold411 (.A(\dtop.field_top.alt_osc[5] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0009_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold413 (.A(\dtop.field_top.afl_pc[4] ),
    .X(net714));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_fill_1 FILLER_0_0 ();
 sg13g2_fill_2 FILLER_0_129 ();
 sg13g2_fill_2 FILLER_0_140 ();
 sg13g2_fill_2 FILLER_0_233 ();
 sg13g2_fill_1 FILLER_0_235 ();
 sg13g2_fill_1 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_fill_2 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_fill_1 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_5 ();
 sg13g2_fill_2 FILLER_1_87 ();
 sg13g2_fill_2 FILLER_1_255 ();
 sg13g2_fill_1 FILLER_1_311 ();
 sg13g2_fill_2 FILLER_1_328 ();
 sg13g2_fill_1 FILLER_1_330 ();
 sg13g2_fill_2 FILLER_1_336 ();
 sg13g2_fill_1 FILLER_1_338 ();
 sg13g2_fill_2 FILLER_1_351 ();
 sg13g2_fill_2 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_fill_2 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_35 ();
 sg13g2_fill_1 FILLER_2_50 ();
 sg13g2_fill_1 FILLER_2_174 ();
 sg13g2_fill_2 FILLER_2_320 ();
 sg13g2_fill_1 FILLER_2_322 ();
 sg13g2_fill_2 FILLER_2_336 ();
 sg13g2_fill_1 FILLER_2_338 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_2 ();
 sg13g2_fill_2 FILLER_3_12 ();
 sg13g2_fill_2 FILLER_3_86 ();
 sg13g2_fill_1 FILLER_3_119 ();
 sg13g2_fill_1 FILLER_3_135 ();
 sg13g2_fill_1 FILLER_3_319 ();
 sg13g2_fill_2 FILLER_3_325 ();
 sg13g2_fill_1 FILLER_3_327 ();
 sg13g2_fill_2 FILLER_3_350 ();
 sg13g2_fill_1 FILLER_4_55 ();
 sg13g2_fill_1 FILLER_4_112 ();
 sg13g2_fill_1 FILLER_4_122 ();
 sg13g2_fill_2 FILLER_4_153 ();
 sg13g2_fill_1 FILLER_4_210 ();
 sg13g2_fill_1 FILLER_4_229 ();
 sg13g2_fill_2 FILLER_4_253 ();
 sg13g2_fill_1 FILLER_4_344 ();
 sg13g2_fill_1 FILLER_4_350 ();
 sg13g2_fill_1 FILLER_4_374 ();
 sg13g2_fill_2 FILLER_4_379 ();
 sg13g2_fill_1 FILLER_4_381 ();
 sg13g2_fill_2 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_213 ();
 sg13g2_fill_1 FILLER_5_215 ();
 sg13g2_fill_1 FILLER_5_233 ();
 sg13g2_fill_1 FILLER_5_240 ();
 sg13g2_fill_1 FILLER_5_282 ();
 sg13g2_fill_1 FILLER_5_321 ();
 sg13g2_fill_2 FILLER_5_370 ();
 sg13g2_fill_2 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_403 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_11 ();
 sg13g2_fill_1 FILLER_6_173 ();
 sg13g2_fill_2 FILLER_6_197 ();
 sg13g2_fill_1 FILLER_6_199 ();
 sg13g2_fill_1 FILLER_6_272 ();
 sg13g2_fill_2 FILLER_6_321 ();
 sg13g2_fill_1 FILLER_6_323 ();
 sg13g2_fill_1 FILLER_6_329 ();
 sg13g2_fill_2 FILLER_6_368 ();
 sg13g2_fill_2 FILLER_6_384 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_39 ();
 sg13g2_fill_1 FILLER_7_133 ();
 sg13g2_fill_2 FILLER_7_189 ();
 sg13g2_fill_2 FILLER_7_305 ();
 sg13g2_fill_1 FILLER_7_322 ();
 sg13g2_fill_2 FILLER_7_348 ();
 sg13g2_fill_1 FILLER_7_366 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_fill_1 FILLER_7_380 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_111 ();
 sg13g2_fill_2 FILLER_8_201 ();
 sg13g2_fill_1 FILLER_8_313 ();
 sg13g2_fill_2 FILLER_8_335 ();
 sg13g2_fill_1 FILLER_8_337 ();
 sg13g2_fill_2 FILLER_8_381 ();
 sg13g2_fill_1 FILLER_8_383 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_fill_2 FILLER_9_26 ();
 sg13g2_fill_1 FILLER_9_209 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_48 ();
 sg13g2_fill_1 FILLER_10_96 ();
 sg13g2_fill_1 FILLER_10_121 ();
 sg13g2_fill_2 FILLER_10_131 ();
 sg13g2_fill_2 FILLER_10_263 ();
 sg13g2_fill_2 FILLER_10_273 ();
 sg13g2_fill_1 FILLER_10_275 ();
 sg13g2_fill_2 FILLER_10_326 ();
 sg13g2_fill_2 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_365 ();
 sg13g2_fill_1 FILLER_10_367 ();
 sg13g2_fill_1 FILLER_10_386 ();
 sg13g2_fill_2 FILLER_10_392 ();
 sg13g2_fill_1 FILLER_11_40 ();
 sg13g2_fill_1 FILLER_11_123 ();
 sg13g2_fill_1 FILLER_11_187 ();
 sg13g2_fill_1 FILLER_11_210 ();
 sg13g2_fill_2 FILLER_11_276 ();
 sg13g2_fill_2 FILLER_11_332 ();
 sg13g2_fill_1 FILLER_11_367 ();
 sg13g2_fill_1 FILLER_11_376 ();
 sg13g2_fill_2 FILLER_11_388 ();
 sg13g2_fill_2 FILLER_12_40 ();
 sg13g2_fill_1 FILLER_12_230 ();
 sg13g2_fill_2 FILLER_12_321 ();
 sg13g2_fill_1 FILLER_12_344 ();
 sg13g2_fill_2 FILLER_12_350 ();
 sg13g2_fill_1 FILLER_12_360 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_fill_1 FILLER_12_397 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_13_26 ();
 sg13g2_fill_2 FILLER_13_106 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_258 ();
 sg13g2_fill_2 FILLER_13_286 ();
 sg13g2_fill_1 FILLER_13_288 ();
 sg13g2_fill_1 FILLER_13_378 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_85 ();
 sg13g2_fill_1 FILLER_14_123 ();
 sg13g2_fill_1 FILLER_14_138 ();
 sg13g2_fill_2 FILLER_14_148 ();
 sg13g2_fill_2 FILLER_14_271 ();
 sg13g2_fill_2 FILLER_14_305 ();
 sg13g2_fill_2 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_337 ();
 sg13g2_fill_2 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_385 ();
 sg13g2_fill_1 FILLER_14_387 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_50 ();
 sg13g2_fill_2 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_293 ();
 sg13g2_fill_2 FILLER_15_359 ();
 sg13g2_fill_1 FILLER_15_361 ();
 sg13g2_fill_2 FILLER_15_373 ();
 sg13g2_fill_1 FILLER_15_375 ();
 sg13g2_fill_2 FILLER_15_382 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_94 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_fill_2 FILLER_16_210 ();
 sg13g2_fill_2 FILLER_16_238 ();
 sg13g2_fill_1 FILLER_16_240 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_fill_1 FILLER_16_332 ();
 sg13g2_fill_1 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_385 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_1 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_166 ();
 sg13g2_fill_2 FILLER_17_325 ();
 sg13g2_fill_1 FILLER_17_327 ();
 sg13g2_fill_2 FILLER_17_351 ();
 sg13g2_fill_1 FILLER_17_353 ();
 sg13g2_fill_1 FILLER_17_363 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_372 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_18_310 ();
 sg13g2_fill_2 FILLER_18_336 ();
 sg13g2_fill_1 FILLER_18_338 ();
 sg13g2_fill_2 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_18_378 ();
 sg13g2_fill_1 FILLER_19_12 ();
 sg13g2_fill_1 FILLER_19_40 ();
 sg13g2_fill_2 FILLER_19_96 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_1 FILLER_19_263 ();
 sg13g2_fill_2 FILLER_19_295 ();
 sg13g2_fill_1 FILLER_19_308 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_fill_1 FILLER_19_325 ();
 sg13g2_fill_2 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_334 ();
 sg13g2_fill_2 FILLER_19_341 ();
 sg13g2_fill_1 FILLER_19_343 ();
 sg13g2_fill_2 FILLER_19_363 ();
 sg13g2_fill_1 FILLER_19_365 ();
 sg13g2_fill_1 FILLER_19_378 ();
 sg13g2_fill_2 FILLER_19_388 ();
 sg13g2_fill_2 FILLER_20_129 ();
 sg13g2_fill_1 FILLER_20_149 ();
 sg13g2_fill_2 FILLER_20_270 ();
 sg13g2_fill_1 FILLER_20_272 ();
 sg13g2_fill_2 FILLER_20_287 ();
 sg13g2_fill_1 FILLER_20_289 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_fill_2 FILLER_20_336 ();
 sg13g2_fill_2 FILLER_20_357 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_1 FILLER_21_79 ();
 sg13g2_fill_2 FILLER_21_90 ();
 sg13g2_fill_2 FILLER_21_127 ();
 sg13g2_fill_1 FILLER_21_139 ();
 sg13g2_fill_2 FILLER_21_185 ();
 sg13g2_fill_1 FILLER_21_209 ();
 sg13g2_fill_1 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_282 ();
 sg13g2_fill_2 FILLER_21_307 ();
 sg13g2_fill_1 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_328 ();
 sg13g2_fill_2 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_385 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_2 FILLER_22_43 ();
 sg13g2_fill_1 FILLER_22_54 ();
 sg13g2_fill_2 FILLER_22_69 ();
 sg13g2_fill_1 FILLER_22_79 ();
 sg13g2_fill_2 FILLER_22_124 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_164 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_fill_2 FILLER_22_195 ();
 sg13g2_fill_2 FILLER_22_212 ();
 sg13g2_fill_1 FILLER_22_258 ();
 sg13g2_fill_1 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_339 ();
 sg13g2_fill_1 FILLER_22_341 ();
 sg13g2_fill_1 FILLER_22_347 ();
 sg13g2_fill_2 FILLER_22_391 ();
 sg13g2_fill_1 FILLER_23_72 ();
 sg13g2_fill_2 FILLER_23_91 ();
 sg13g2_fill_1 FILLER_23_110 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_fill_1 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_fill_2 FILLER_23_350 ();
 sg13g2_fill_1 FILLER_23_352 ();
 sg13g2_fill_1 FILLER_23_363 ();
 sg13g2_fill_1 FILLER_23_380 ();
 sg13g2_fill_2 FILLER_23_388 ();
 sg13g2_fill_1 FILLER_23_390 ();
 sg13g2_fill_1 FILLER_24_19 ();
 sg13g2_fill_1 FILLER_24_52 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_fill_1 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_243 ();
 sg13g2_fill_2 FILLER_24_267 ();
 sg13g2_fill_2 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_376 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_73 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_302 ();
 sg13g2_fill_2 FILLER_25_343 ();
 sg13g2_fill_2 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_fill_1 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_fill_1 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_101 ();
 sg13g2_fill_1 FILLER_27_116 ();
 sg13g2_fill_2 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_fill_2 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_2 FILLER_27_290 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_fill_2 FILLER_27_344 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_decap_4 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_fill_2 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_fill_2 FILLER_28_19 ();
 sg13g2_fill_2 FILLER_28_74 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_decap_4 FILLER_28_365 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_decap_4 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_29_17 ();
 sg13g2_fill_1 FILLER_29_179 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_fill_2 FILLER_29_195 ();
 sg13g2_fill_1 FILLER_29_197 ();
 sg13g2_fill_2 FILLER_29_220 ();
 sg13g2_fill_2 FILLER_29_290 ();
 sg13g2_fill_2 FILLER_29_323 ();
 sg13g2_fill_1 FILLER_29_325 ();
 sg13g2_fill_1 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_15 ();
 sg13g2_fill_2 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_152 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_194 ();
 sg13g2_fill_2 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_279 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_354 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_fill_2 FILLER_30_364 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_fill_1 FILLER_31_39 ();
 sg13g2_fill_2 FILLER_31_93 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_fill_2 FILLER_31_159 ();
 sg13g2_fill_2 FILLER_31_206 ();
 sg13g2_fill_2 FILLER_31_264 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_361 ();
 sg13g2_fill_1 FILLER_31_391 ();
 sg13g2_fill_1 FILLER_31_402 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_36 ();
 sg13g2_fill_1 FILLER_32_47 ();
 sg13g2_fill_1 FILLER_32_75 ();
 sg13g2_fill_2 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_176 ();
 sg13g2_fill_1 FILLER_32_288 ();
 sg13g2_fill_2 FILLER_32_327 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_349 ();
 sg13g2_fill_2 FILLER_32_361 ();
 sg13g2_fill_2 FILLER_32_380 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_fill_2 FILLER_33_26 ();
 sg13g2_fill_1 FILLER_33_46 ();
 sg13g2_fill_2 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_116 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_281 ();
 sg13g2_fill_2 FILLER_33_330 ();
 sg13g2_fill_2 FILLER_33_348 ();
 sg13g2_fill_1 FILLER_33_350 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_fill_1 FILLER_33_383 ();
 sg13g2_fill_2 FILLER_33_397 ();
 sg13g2_fill_1 FILLER_33_399 ();
 sg13g2_fill_1 FILLER_34_73 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_fill_1 FILLER_34_133 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_174 ();
 sg13g2_fill_2 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_237 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_346 ();
 sg13g2_fill_2 FILLER_34_354 ();
 sg13g2_fill_1 FILLER_34_374 ();
 sg13g2_fill_2 FILLER_34_380 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_fill_2 FILLER_35_26 ();
 sg13g2_fill_1 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_145 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_275 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_fill_2 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_326 ();
 sg13g2_fill_2 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_334 ();
 sg13g2_fill_1 FILLER_35_350 ();
 sg13g2_fill_2 FILLER_35_390 ();
 sg13g2_fill_1 FILLER_35_392 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_fill_2 FILLER_36_85 ();
 sg13g2_fill_2 FILLER_36_93 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_fill_1 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_289 ();
 sg13g2_decap_4 FILLER_36_313 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_37_44 ();
 sg13g2_fill_2 FILLER_37_55 ();
 sg13g2_fill_2 FILLER_37_106 ();
 sg13g2_fill_2 FILLER_37_113 ();
 sg13g2_fill_1 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_fill_2 FILLER_37_265 ();
 sg13g2_fill_1 FILLER_37_267 ();
 sg13g2_fill_1 FILLER_37_310 ();
 sg13g2_fill_1 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_320 ();
 sg13g2_fill_1 FILLER_37_327 ();
 sg13g2_decap_4 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_fill_1 FILLER_38_45 ();
 sg13g2_fill_1 FILLER_38_55 ();
 sg13g2_fill_2 FILLER_38_73 ();
 sg13g2_fill_1 FILLER_38_75 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_fill_2 FILLER_38_114 ();
 sg13g2_fill_1 FILLER_38_116 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_fill_2 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_decap_4 FILLER_38_255 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_338 ();
 sg13g2_fill_1 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_365 ();
 sg13g2_fill_2 FILLER_38_390 ();
 sg13g2_fill_1 FILLER_38_392 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_fill_1 FILLER_39_31 ();
 sg13g2_fill_2 FILLER_39_66 ();
 sg13g2_fill_1 FILLER_39_68 ();
 sg13g2_fill_2 FILLER_39_113 ();
 sg13g2_fill_2 FILLER_39_169 ();
 sg13g2_fill_1 FILLER_39_183 ();
 sg13g2_fill_2 FILLER_39_205 ();
 sg13g2_fill_1 FILLER_39_207 ();
 sg13g2_fill_1 FILLER_39_215 ();
 sg13g2_fill_1 FILLER_39_254 ();
 sg13g2_fill_2 FILLER_39_321 ();
 sg13g2_fill_2 FILLER_39_339 ();
 sg13g2_fill_1 FILLER_39_341 ();
 sg13g2_fill_1 FILLER_39_395 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_21 ();
 sg13g2_fill_1 FILLER_40_42 ();
 sg13g2_fill_2 FILLER_40_64 ();
 sg13g2_fill_1 FILLER_40_113 ();
 sg13g2_fill_1 FILLER_40_126 ();
 sg13g2_fill_1 FILLER_40_133 ();
 sg13g2_fill_1 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_171 ();
 sg13g2_fill_2 FILLER_40_251 ();
 sg13g2_fill_1 FILLER_40_253 ();
 sg13g2_fill_2 FILLER_40_264 ();
 sg13g2_fill_1 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_358 ();
 sg13g2_fill_1 FILLER_40_365 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_fill_2 FILLER_40_385 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_fill_2 FILLER_41_30 ();
 sg13g2_fill_1 FILLER_41_58 ();
 sg13g2_fill_1 FILLER_41_68 ();
 sg13g2_fill_1 FILLER_41_201 ();
 sg13g2_fill_2 FILLER_41_206 ();
 sg13g2_decap_4 FILLER_41_225 ();
 sg13g2_fill_1 FILLER_41_238 ();
 sg13g2_fill_2 FILLER_41_308 ();
 sg13g2_fill_1 FILLER_41_310 ();
 sg13g2_fill_2 FILLER_41_363 ();
 sg13g2_fill_2 FILLER_41_379 ();
 sg13g2_fill_1 FILLER_41_381 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_fill_1 FILLER_42_26 ();
 sg13g2_fill_1 FILLER_42_54 ();
 sg13g2_fill_2 FILLER_42_81 ();
 sg13g2_fill_2 FILLER_42_95 ();
 sg13g2_fill_1 FILLER_42_97 ();
 sg13g2_fill_1 FILLER_42_104 ();
 sg13g2_decap_4 FILLER_42_184 ();
 sg13g2_fill_1 FILLER_42_202 ();
 sg13g2_fill_1 FILLER_42_262 ();
 sg13g2_fill_2 FILLER_42_276 ();
 sg13g2_fill_1 FILLER_42_294 ();
 sg13g2_fill_1 FILLER_42_314 ();
 sg13g2_fill_1 FILLER_42_332 ();
 sg13g2_fill_2 FILLER_42_341 ();
 sg13g2_fill_2 FILLER_42_357 ();
 sg13g2_fill_1 FILLER_42_359 ();
 sg13g2_fill_2 FILLER_42_384 ();
 sg13g2_fill_1 FILLER_42_386 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_fill_2 FILLER_43_26 ();
 sg13g2_fill_1 FILLER_43_102 ();
 sg13g2_fill_2 FILLER_43_158 ();
 sg13g2_fill_2 FILLER_43_206 ();
 sg13g2_fill_1 FILLER_43_208 ();
 sg13g2_fill_2 FILLER_43_214 ();
 sg13g2_fill_1 FILLER_43_216 ();
 sg13g2_decap_4 FILLER_43_243 ();
 sg13g2_fill_2 FILLER_43_257 ();
 sg13g2_fill_1 FILLER_43_274 ();
 sg13g2_fill_1 FILLER_43_305 ();
 sg13g2_fill_1 FILLER_43_347 ();
 sg13g2_fill_2 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_48 ();
 sg13g2_fill_1 FILLER_44_77 ();
 sg13g2_fill_1 FILLER_44_94 ();
 sg13g2_fill_1 FILLER_44_118 ();
 sg13g2_fill_1 FILLER_44_185 ();
 sg13g2_fill_1 FILLER_44_195 ();
 sg13g2_fill_1 FILLER_44_236 ();
 sg13g2_fill_1 FILLER_44_268 ();
 sg13g2_fill_1 FILLER_44_278 ();
 sg13g2_fill_1 FILLER_44_289 ();
 sg13g2_decap_8 FILLER_44_304 ();
 sg13g2_fill_2 FILLER_44_311 ();
 sg13g2_fill_1 FILLER_44_313 ();
 sg13g2_fill_1 FILLER_44_352 ();
 sg13g2_fill_1 FILLER_44_365 ();
 sg13g2_fill_1 FILLER_44_394 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_94 ();
 sg13g2_fill_1 FILLER_45_125 ();
 sg13g2_fill_2 FILLER_45_149 ();
 sg13g2_fill_1 FILLER_45_151 ();
 sg13g2_fill_1 FILLER_45_180 ();
 sg13g2_decap_8 FILLER_45_226 ();
 sg13g2_decap_8 FILLER_45_233 ();
 sg13g2_decap_8 FILLER_45_240 ();
 sg13g2_decap_4 FILLER_45_247 ();
 sg13g2_fill_1 FILLER_45_251 ();
 sg13g2_fill_2 FILLER_45_261 ();
 sg13g2_fill_2 FILLER_45_288 ();
 sg13g2_fill_1 FILLER_45_290 ();
 sg13g2_fill_2 FILLER_45_298 ();
 sg13g2_fill_1 FILLER_45_300 ();
 sg13g2_decap_4 FILLER_45_314 ();
 sg13g2_fill_1 FILLER_45_347 ();
 sg13g2_fill_1 FILLER_45_360 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_78 ();
 sg13g2_fill_1 FILLER_46_83 ();
 sg13g2_fill_1 FILLER_46_93 ();
 sg13g2_fill_2 FILLER_46_122 ();
 sg13g2_fill_1 FILLER_46_147 ();
 sg13g2_fill_2 FILLER_46_192 ();
 sg13g2_fill_2 FILLER_46_235 ();
 sg13g2_fill_1 FILLER_46_237 ();
 sg13g2_decap_4 FILLER_46_323 ();
 sg13g2_fill_2 FILLER_46_327 ();
 sg13g2_fill_2 FILLER_46_352 ();
 sg13g2_fill_1 FILLER_46_377 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_27 ();
 sg13g2_fill_1 FILLER_47_29 ();
 sg13g2_fill_1 FILLER_47_39 ();
 sg13g2_fill_2 FILLER_47_57 ();
 sg13g2_fill_2 FILLER_47_80 ();
 sg13g2_fill_2 FILLER_47_88 ();
 sg13g2_fill_1 FILLER_47_129 ();
 sg13g2_fill_1 FILLER_47_140 ();
 sg13g2_fill_1 FILLER_47_151 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_fill_2 FILLER_47_206 ();
 sg13g2_fill_2 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_348 ();
 sg13g2_fill_2 FILLER_47_355 ();
 sg13g2_fill_2 FILLER_47_375 ();
 sg13g2_fill_1 FILLER_47_377 ();
 sg13g2_fill_2 FILLER_47_386 ();
 sg13g2_fill_2 FILLER_47_398 ();
 sg13g2_fill_1 FILLER_48_26 ();
 sg13g2_fill_2 FILLER_48_42 ();
 sg13g2_fill_1 FILLER_48_44 ();
 sg13g2_fill_1 FILLER_48_91 ();
 sg13g2_fill_1 FILLER_48_102 ();
 sg13g2_fill_1 FILLER_48_121 ();
 sg13g2_fill_1 FILLER_48_129 ();
 sg13g2_fill_1 FILLER_48_135 ();
 sg13g2_fill_2 FILLER_48_142 ();
 sg13g2_fill_1 FILLER_48_144 ();
 sg13g2_fill_1 FILLER_48_153 ();
 sg13g2_fill_2 FILLER_48_172 ();
 sg13g2_fill_1 FILLER_48_205 ();
 sg13g2_fill_1 FILLER_48_215 ();
 sg13g2_fill_2 FILLER_48_225 ();
 sg13g2_fill_2 FILLER_48_245 ();
 sg13g2_fill_1 FILLER_48_247 ();
 sg13g2_fill_2 FILLER_48_271 ();
 sg13g2_fill_1 FILLER_48_273 ();
 sg13g2_fill_1 FILLER_48_296 ();
 sg13g2_decap_8 FILLER_48_340 ();
 sg13g2_decap_8 FILLER_48_347 ();
 sg13g2_fill_1 FILLER_48_354 ();
 sg13g2_fill_1 FILLER_48_370 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_116 ();
 sg13g2_fill_1 FILLER_49_146 ();
 sg13g2_decap_8 FILLER_49_152 ();
 sg13g2_decap_8 FILLER_49_162 ();
 sg13g2_fill_2 FILLER_49_169 ();
 sg13g2_fill_1 FILLER_49_171 ();
 sg13g2_fill_1 FILLER_49_218 ();
 sg13g2_fill_2 FILLER_49_264 ();
 sg13g2_fill_1 FILLER_49_266 ();
 sg13g2_fill_2 FILLER_49_292 ();
 sg13g2_fill_1 FILLER_49_294 ();
 sg13g2_fill_1 FILLER_49_302 ();
 sg13g2_fill_2 FILLER_49_309 ();
 sg13g2_fill_2 FILLER_49_332 ();
 sg13g2_fill_2 FILLER_49_375 ();
 sg13g2_fill_2 FILLER_50_26 ();
 sg13g2_fill_2 FILLER_50_61 ();
 sg13g2_fill_1 FILLER_50_76 ();
 sg13g2_fill_2 FILLER_50_86 ();
 sg13g2_fill_1 FILLER_50_151 ();
 sg13g2_fill_1 FILLER_50_164 ();
 sg13g2_fill_1 FILLER_50_197 ();
 sg13g2_fill_1 FILLER_50_259 ();
 sg13g2_fill_2 FILLER_50_269 ();
 sg13g2_fill_1 FILLER_50_289 ();
 sg13g2_fill_2 FILLER_50_296 ();
 sg13g2_fill_1 FILLER_50_298 ();
 sg13g2_fill_2 FILLER_50_305 ();
 sg13g2_fill_2 FILLER_50_335 ();
 sg13g2_fill_2 FILLER_50_378 ();
 sg13g2_fill_1 FILLER_50_391 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_fill_1 FILLER_51_41 ();
 sg13g2_fill_2 FILLER_51_52 ();
 sg13g2_fill_2 FILLER_51_59 ();
 sg13g2_decap_4 FILLER_51_69 ();
 sg13g2_fill_1 FILLER_51_86 ();
 sg13g2_fill_2 FILLER_51_103 ();
 sg13g2_fill_1 FILLER_51_166 ();
 sg13g2_fill_1 FILLER_51_193 ();
 sg13g2_fill_2 FILLER_51_225 ();
 sg13g2_fill_1 FILLER_51_227 ();
 sg13g2_fill_2 FILLER_51_291 ();
 sg13g2_fill_1 FILLER_51_293 ();
 sg13g2_fill_1 FILLER_51_302 ();
 sg13g2_fill_2 FILLER_51_341 ();
 sg13g2_fill_1 FILLER_51_366 ();
 sg13g2_fill_2 FILLER_51_372 ();
 sg13g2_fill_1 FILLER_51_374 ();
 sg13g2_fill_1 FILLER_51_394 ();
 sg13g2_fill_1 FILLER_52_18 ();
 sg13g2_fill_2 FILLER_52_62 ();
 sg13g2_fill_2 FILLER_52_110 ();
 sg13g2_fill_2 FILLER_52_120 ();
 sg13g2_fill_1 FILLER_52_154 ();
 sg13g2_fill_1 FILLER_52_216 ();
 sg13g2_fill_2 FILLER_52_297 ();
 sg13g2_fill_1 FILLER_52_310 ();
 sg13g2_fill_2 FILLER_52_340 ();
 sg13g2_fill_1 FILLER_52_342 ();
 sg13g2_fill_2 FILLER_52_356 ();
 sg13g2_fill_1 FILLER_52_358 ();
 sg13g2_fill_2 FILLER_52_383 ();
 sg13g2_fill_1 FILLER_52_385 ();
 sg13g2_fill_1 FILLER_53_73 ();
 sg13g2_fill_1 FILLER_53_91 ();
 sg13g2_fill_2 FILLER_53_109 ();
 sg13g2_fill_2 FILLER_53_123 ();
 sg13g2_fill_1 FILLER_53_125 ();
 sg13g2_fill_2 FILLER_53_155 ();
 sg13g2_fill_2 FILLER_53_168 ();
 sg13g2_fill_2 FILLER_53_178 ();
 sg13g2_decap_8 FILLER_53_187 ();
 sg13g2_fill_2 FILLER_53_194 ();
 sg13g2_fill_1 FILLER_53_208 ();
 sg13g2_decap_8 FILLER_53_213 ();
 sg13g2_fill_1 FILLER_53_220 ();
 sg13g2_fill_1 FILLER_53_234 ();
 sg13g2_fill_1 FILLER_53_277 ();
 sg13g2_fill_2 FILLER_53_321 ();
 sg13g2_fill_2 FILLER_53_355 ();
 sg13g2_fill_2 FILLER_53_383 ();
 sg13g2_fill_2 FILLER_54_26 ();
 sg13g2_fill_2 FILLER_54_72 ();
 sg13g2_fill_1 FILLER_54_74 ();
 sg13g2_fill_2 FILLER_54_93 ();
 sg13g2_fill_1 FILLER_54_129 ();
 sg13g2_fill_2 FILLER_54_135 ();
 sg13g2_fill_1 FILLER_54_170 ();
 sg13g2_decap_4 FILLER_54_176 ();
 sg13g2_fill_1 FILLER_54_180 ();
 sg13g2_fill_1 FILLER_54_185 ();
 sg13g2_fill_1 FILLER_54_195 ();
 sg13g2_fill_2 FILLER_54_218 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_fill_2 FILLER_54_226 ();
 sg13g2_fill_1 FILLER_54_228 ();
 sg13g2_decap_4 FILLER_54_234 ();
 sg13g2_fill_1 FILLER_54_271 ();
 sg13g2_fill_1 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_299 ();
 sg13g2_fill_1 FILLER_54_319 ();
 sg13g2_fill_1 FILLER_54_346 ();
 sg13g2_fill_1 FILLER_54_388 ();
 sg13g2_fill_2 FILLER_55_54 ();
 sg13g2_decap_8 FILLER_55_78 ();
 sg13g2_decap_4 FILLER_55_91 ();
 sg13g2_fill_1 FILLER_55_95 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_fill_2 FILLER_55_118 ();
 sg13g2_fill_1 FILLER_55_120 ();
 sg13g2_fill_1 FILLER_55_169 ();
 sg13g2_fill_2 FILLER_55_178 ();
 sg13g2_fill_1 FILLER_55_180 ();
 sg13g2_fill_2 FILLER_55_301 ();
 sg13g2_fill_2 FILLER_55_336 ();
 sg13g2_fill_1 FILLER_55_348 ();
 sg13g2_fill_2 FILLER_55_357 ();
 sg13g2_fill_1 FILLER_56_57 ();
 sg13g2_fill_2 FILLER_56_67 ();
 sg13g2_fill_1 FILLER_56_69 ();
 sg13g2_fill_2 FILLER_56_74 ();
 sg13g2_fill_1 FILLER_56_76 ();
 sg13g2_fill_2 FILLER_56_95 ();
 sg13g2_fill_1 FILLER_56_97 ();
 sg13g2_fill_1 FILLER_56_120 ();
 sg13g2_fill_2 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_132 ();
 sg13g2_fill_2 FILLER_56_138 ();
 sg13g2_fill_1 FILLER_56_140 ();
 sg13g2_fill_1 FILLER_56_175 ();
 sg13g2_fill_2 FILLER_56_202 ();
 sg13g2_fill_2 FILLER_56_327 ();
 sg13g2_fill_1 FILLER_56_329 ();
 sg13g2_fill_2 FILLER_56_356 ();
 sg13g2_fill_2 FILLER_56_389 ();
 sg13g2_fill_1 FILLER_56_391 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_36 ();
 sg13g2_fill_1 FILLER_57_38 ();
 sg13g2_fill_2 FILLER_57_59 ();
 sg13g2_fill_1 FILLER_57_104 ();
 sg13g2_fill_2 FILLER_57_120 ();
 sg13g2_fill_2 FILLER_57_128 ();
 sg13g2_fill_1 FILLER_57_136 ();
 sg13g2_fill_2 FILLER_57_143 ();
 sg13g2_fill_2 FILLER_57_153 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_fill_1 FILLER_57_184 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_fill_2 FILLER_57_251 ();
 sg13g2_fill_1 FILLER_57_298 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_fill_2 FILLER_57_358 ();
 sg13g2_fill_1 FILLER_57_360 ();
 sg13g2_fill_2 FILLER_57_392 ();
 sg13g2_fill_1 FILLER_57_394 ();
 sg13g2_fill_2 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_fill_1 FILLER_58_47 ();
 sg13g2_fill_1 FILLER_58_64 ();
 sg13g2_fill_2 FILLER_58_71 ();
 sg13g2_fill_2 FILLER_58_94 ();
 sg13g2_fill_2 FILLER_58_101 ();
 sg13g2_fill_1 FILLER_58_103 ();
 sg13g2_fill_1 FILLER_58_131 ();
 sg13g2_fill_1 FILLER_58_138 ();
 sg13g2_fill_1 FILLER_58_144 ();
 sg13g2_decap_4 FILLER_58_154 ();
 sg13g2_fill_1 FILLER_58_158 ();
 sg13g2_fill_2 FILLER_58_202 ();
 sg13g2_fill_2 FILLER_58_244 ();
 sg13g2_fill_2 FILLER_58_251 ();
 sg13g2_fill_2 FILLER_58_266 ();
 sg13g2_fill_2 FILLER_58_276 ();
 sg13g2_fill_2 FILLER_58_290 ();
 sg13g2_fill_1 FILLER_58_292 ();
 sg13g2_fill_2 FILLER_58_323 ();
 sg13g2_fill_2 FILLER_58_354 ();
 sg13g2_fill_1 FILLER_58_356 ();
 sg13g2_fill_2 FILLER_58_380 ();
 sg13g2_fill_2 FILLER_58_388 ();
 sg13g2_fill_2 FILLER_59_26 ();
 sg13g2_fill_1 FILLER_59_28 ();
 sg13g2_fill_2 FILLER_59_57 ();
 sg13g2_fill_2 FILLER_59_90 ();
 sg13g2_fill_1 FILLER_59_143 ();
 sg13g2_fill_2 FILLER_59_168 ();
 sg13g2_fill_2 FILLER_59_195 ();
 sg13g2_fill_1 FILLER_59_197 ();
 sg13g2_fill_2 FILLER_59_221 ();
 sg13g2_fill_2 FILLER_59_253 ();
 sg13g2_fill_1 FILLER_59_255 ();
 sg13g2_fill_2 FILLER_59_282 ();
 sg13g2_fill_1 FILLER_59_284 ();
 sg13g2_fill_1 FILLER_59_295 ();
 sg13g2_fill_2 FILLER_59_301 ();
 sg13g2_fill_1 FILLER_59_303 ();
 sg13g2_fill_1 FILLER_59_341 ();
 sg13g2_fill_2 FILLER_59_355 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_2 ();
 sg13g2_fill_2 FILLER_60_37 ();
 sg13g2_fill_2 FILLER_60_47 ();
 sg13g2_fill_1 FILLER_60_49 ();
 sg13g2_fill_1 FILLER_60_126 ();
 sg13g2_fill_1 FILLER_60_143 ();
 sg13g2_fill_2 FILLER_60_154 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_fill_1 FILLER_60_212 ();
 sg13g2_fill_2 FILLER_60_220 ();
 sg13g2_fill_1 FILLER_60_254 ();
 sg13g2_fill_2 FILLER_60_304 ();
 sg13g2_fill_2 FILLER_60_347 ();
 sg13g2_fill_2 FILLER_60_371 ();
 sg13g2_fill_1 FILLER_60_383 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_7 ();
 sg13g2_fill_1 FILLER_61_17 ();
 sg13g2_fill_2 FILLER_61_39 ();
 sg13g2_decap_4 FILLER_61_60 ();
 sg13g2_fill_2 FILLER_61_96 ();
 sg13g2_fill_2 FILLER_61_110 ();
 sg13g2_fill_2 FILLER_61_123 ();
 sg13g2_fill_1 FILLER_61_125 ();
 sg13g2_decap_4 FILLER_61_140 ();
 sg13g2_fill_1 FILLER_61_144 ();
 sg13g2_fill_2 FILLER_61_167 ();
 sg13g2_fill_1 FILLER_61_195 ();
 sg13g2_fill_1 FILLER_61_216 ();
 sg13g2_fill_1 FILLER_61_367 ();
 sg13g2_fill_2 FILLER_61_382 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_9 ();
 sg13g2_fill_2 FILLER_62_38 ();
 sg13g2_fill_1 FILLER_62_40 ();
 sg13g2_fill_2 FILLER_62_45 ();
 sg13g2_fill_1 FILLER_62_47 ();
 sg13g2_fill_2 FILLER_62_60 ();
 sg13g2_fill_1 FILLER_62_78 ();
 sg13g2_fill_2 FILLER_62_100 ();
 sg13g2_fill_2 FILLER_62_111 ();
 sg13g2_decap_4 FILLER_62_136 ();
 sg13g2_fill_2 FILLER_62_140 ();
 sg13g2_fill_2 FILLER_62_182 ();
 sg13g2_fill_1 FILLER_62_184 ();
 sg13g2_fill_2 FILLER_62_197 ();
 sg13g2_fill_1 FILLER_62_228 ();
 sg13g2_fill_2 FILLER_62_237 ();
 sg13g2_fill_1 FILLER_62_239 ();
 sg13g2_fill_2 FILLER_62_279 ();
 sg13g2_fill_1 FILLER_62_281 ();
 sg13g2_fill_1 FILLER_62_292 ();
 sg13g2_fill_2 FILLER_62_329 ();
 sg13g2_fill_2 FILLER_62_349 ();
 sg13g2_fill_2 FILLER_62_362 ();
 sg13g2_fill_2 FILLER_62_403 ();
 sg13g2_fill_2 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_45 ();
 sg13g2_fill_1 FILLER_63_55 ();
 sg13g2_fill_2 FILLER_63_62 ();
 sg13g2_fill_2 FILLER_63_87 ();
 sg13g2_fill_1 FILLER_63_93 ();
 sg13g2_decap_4 FILLER_63_102 ();
 sg13g2_decap_4 FILLER_63_110 ();
 sg13g2_fill_2 FILLER_63_114 ();
 sg13g2_fill_2 FILLER_63_138 ();
 sg13g2_fill_1 FILLER_63_140 ();
 sg13g2_fill_1 FILLER_63_145 ();
 sg13g2_fill_2 FILLER_63_170 ();
 sg13g2_fill_1 FILLER_63_172 ();
 sg13g2_decap_4 FILLER_63_192 ();
 sg13g2_decap_4 FILLER_63_200 ();
 sg13g2_fill_2 FILLER_63_224 ();
 sg13g2_fill_1 FILLER_63_283 ();
 sg13g2_fill_1 FILLER_63_312 ();
 sg13g2_fill_2 FILLER_63_321 ();
 sg13g2_fill_2 FILLER_63_327 ();
 sg13g2_fill_2 FILLER_63_344 ();
 sg13g2_fill_1 FILLER_63_383 ();
 sg13g2_decap_4 FILLER_64_101 ();
 sg13g2_fill_1 FILLER_64_105 ();
 sg13g2_fill_1 FILLER_64_126 ();
 sg13g2_fill_1 FILLER_64_137 ();
 sg13g2_fill_2 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_157 ();
 sg13g2_decap_4 FILLER_64_164 ();
 sg13g2_fill_1 FILLER_64_168 ();
 sg13g2_fill_2 FILLER_64_173 ();
 sg13g2_fill_1 FILLER_64_185 ();
 sg13g2_fill_1 FILLER_64_189 ();
 sg13g2_fill_1 FILLER_64_208 ();
 sg13g2_fill_1 FILLER_64_253 ();
 sg13g2_fill_2 FILLER_64_264 ();
 sg13g2_fill_1 FILLER_64_266 ();
 sg13g2_fill_2 FILLER_64_302 ();
 sg13g2_fill_1 FILLER_64_336 ();
 sg13g2_fill_1 FILLER_64_348 ();
 sg13g2_fill_1 FILLER_64_359 ();
 sg13g2_fill_1 FILLER_64_385 ();
 sg13g2_fill_2 FILLER_64_392 ();
 sg13g2_fill_1 FILLER_64_394 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_78 ();
 sg13g2_fill_2 FILLER_65_104 ();
 sg13g2_fill_1 FILLER_65_106 ();
 sg13g2_fill_2 FILLER_65_164 ();
 sg13g2_fill_1 FILLER_65_166 ();
 sg13g2_fill_2 FILLER_65_172 ();
 sg13g2_fill_1 FILLER_65_174 ();
 sg13g2_fill_2 FILLER_65_199 ();
 sg13g2_fill_1 FILLER_65_221 ();
 sg13g2_fill_1 FILLER_65_265 ();
 sg13g2_fill_2 FILLER_65_364 ();
 sg13g2_fill_1 FILLER_65_380 ();
 sg13g2_fill_2 FILLER_65_387 ();
 sg13g2_fill_2 FILLER_65_394 ();
 sg13g2_fill_1 FILLER_65_396 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_28 ();
 sg13g2_fill_2 FILLER_66_41 ();
 sg13g2_fill_1 FILLER_66_43 ();
 sg13g2_fill_1 FILLER_66_57 ();
 sg13g2_fill_1 FILLER_66_66 ();
 sg13g2_fill_2 FILLER_66_106 ();
 sg13g2_fill_1 FILLER_66_176 ();
 sg13g2_fill_1 FILLER_66_210 ();
 sg13g2_fill_1 FILLER_66_290 ();
 sg13g2_fill_2 FILLER_66_325 ();
 sg13g2_fill_1 FILLER_66_335 ();
 sg13g2_fill_2 FILLER_66_350 ();
 sg13g2_fill_1 FILLER_66_389 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_35 ();
 sg13g2_fill_1 FILLER_67_37 ();
 sg13g2_fill_1 FILLER_67_43 ();
 sg13g2_fill_2 FILLER_67_73 ();
 sg13g2_fill_2 FILLER_67_118 ();
 sg13g2_fill_2 FILLER_67_130 ();
 sg13g2_fill_1 FILLER_67_132 ();
 sg13g2_fill_1 FILLER_67_147 ();
 sg13g2_fill_2 FILLER_67_267 ();
 sg13g2_fill_2 FILLER_67_359 ();
 sg13g2_fill_2 FILLER_67_377 ();
 sg13g2_fill_1 FILLER_67_392 ();
 sg13g2_fill_1 FILLER_67_402 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_39 ();
 sg13g2_fill_2 FILLER_68_56 ();
 sg13g2_fill_1 FILLER_68_97 ();
 sg13g2_fill_1 FILLER_68_173 ();
 sg13g2_fill_2 FILLER_68_276 ();
 sg13g2_fill_2 FILLER_68_325 ();
 sg13g2_fill_1 FILLER_68_327 ();
 sg13g2_fill_2 FILLER_68_351 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_51 ();
 sg13g2_fill_2 FILLER_69_60 ();
 sg13g2_fill_1 FILLER_69_76 ();
 sg13g2_fill_1 FILLER_69_85 ();
 sg13g2_fill_1 FILLER_69_93 ();
 sg13g2_fill_1 FILLER_69_115 ();
 sg13g2_fill_1 FILLER_69_151 ();
 sg13g2_fill_1 FILLER_69_157 ();
 sg13g2_fill_2 FILLER_69_194 ();
 sg13g2_fill_2 FILLER_69_212 ();
 sg13g2_fill_2 FILLER_69_240 ();
 sg13g2_fill_1 FILLER_69_287 ();
 sg13g2_fill_2 FILLER_69_306 ();
 sg13g2_fill_2 FILLER_69_313 ();
 sg13g2_fill_2 FILLER_69_336 ();
 sg13g2_fill_1 FILLER_69_338 ();
 sg13g2_fill_1 FILLER_69_382 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_33 ();
 sg13g2_fill_2 FILLER_70_54 ();
 sg13g2_fill_1 FILLER_70_56 ();
 sg13g2_fill_2 FILLER_70_63 ();
 sg13g2_fill_1 FILLER_70_65 ();
 sg13g2_fill_2 FILLER_70_86 ();
 sg13g2_fill_2 FILLER_70_147 ();
 sg13g2_fill_2 FILLER_70_172 ();
 sg13g2_fill_2 FILLER_70_220 ();
 sg13g2_fill_1 FILLER_70_282 ();
 sg13g2_fill_1 FILLER_70_352 ();
 sg13g2_fill_2 FILLER_70_362 ();
 sg13g2_fill_1 FILLER_70_364 ();
 sg13g2_fill_1 FILLER_70_393 ();
 sg13g2_fill_1 FILLER_70_398 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_decap_4 FILLER_71_5 ();
 sg13g2_decap_8 FILLER_71_18 ();
 sg13g2_fill_2 FILLER_71_25 ();
 sg13g2_fill_1 FILLER_71_44 ();
 sg13g2_fill_1 FILLER_71_49 ();
 sg13g2_fill_2 FILLER_71_69 ();
 sg13g2_fill_1 FILLER_71_71 ();
 sg13g2_fill_1 FILLER_71_180 ();
 sg13g2_fill_1 FILLER_71_200 ();
 sg13g2_fill_2 FILLER_71_241 ();
 sg13g2_fill_1 FILLER_71_279 ();
 sg13g2_fill_2 FILLER_71_348 ();
 sg13g2_fill_2 FILLER_71_381 ();
 sg13g2_fill_1 FILLER_71_396 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_30 ();
 sg13g2_fill_2 FILLER_72_53 ();
 sg13g2_fill_1 FILLER_72_55 ();
 sg13g2_fill_2 FILLER_72_78 ();
 sg13g2_fill_2 FILLER_72_89 ();
 sg13g2_fill_1 FILLER_72_197 ();
 sg13g2_fill_2 FILLER_72_251 ();
 sg13g2_fill_2 FILLER_72_258 ();
 sg13g2_fill_1 FILLER_72_260 ();
 sg13g2_fill_2 FILLER_72_345 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_45 ();
 sg13g2_fill_2 FILLER_73_55 ();
 sg13g2_fill_2 FILLER_73_77 ();
 sg13g2_fill_1 FILLER_73_109 ();
 sg13g2_fill_1 FILLER_73_136 ();
 sg13g2_fill_1 FILLER_73_160 ();
 sg13g2_fill_2 FILLER_73_175 ();
 sg13g2_fill_2 FILLER_73_252 ();
 sg13g2_fill_2 FILLER_73_269 ();
 sg13g2_fill_2 FILLER_73_327 ();
 sg13g2_fill_1 FILLER_73_339 ();
 sg13g2_fill_2 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_37 ();
 sg13g2_fill_1 FILLER_74_43 ();
 sg13g2_fill_2 FILLER_74_75 ();
 sg13g2_fill_1 FILLER_74_90 ();
 sg13g2_fill_2 FILLER_74_188 ();
 sg13g2_fill_2 FILLER_74_213 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_110 ();
 sg13g2_fill_2 FILLER_75_141 ();
 sg13g2_fill_1 FILLER_75_162 ();
 sg13g2_fill_2 FILLER_75_172 ();
 sg13g2_fill_1 FILLER_75_211 ();
 sg13g2_fill_1 FILLER_75_256 ();
 sg13g2_fill_1 FILLER_75_306 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_37 ();
 sg13g2_fill_2 FILLER_76_87 ();
 sg13g2_fill_1 FILLER_76_115 ();
 sg13g2_fill_1 FILLER_76_191 ();
 sg13g2_fill_1 FILLER_76_270 ();
 sg13g2_fill_1 FILLER_76_276 ();
 sg13g2_fill_2 FILLER_76_303 ();
 sg13g2_fill_1 FILLER_76_305 ();
 sg13g2_fill_2 FILLER_76_332 ();
 sg13g2_fill_2 FILLER_76_370 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_157 ();
 sg13g2_fill_1 FILLER_77_244 ();
 sg13g2_fill_2 FILLER_77_291 ();
 sg13g2_fill_1 FILLER_77_324 ();
 sg13g2_decap_4 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_34 ();
 sg13g2_fill_1 FILLER_78_48 ();
 sg13g2_fill_2 FILLER_78_65 ();
 sg13g2_fill_1 FILLER_78_99 ();
 sg13g2_fill_2 FILLER_78_209 ();
 sg13g2_fill_1 FILLER_78_245 ();
 sg13g2_fill_1 FILLER_78_277 ();
 sg13g2_fill_2 FILLER_78_288 ();
 sg13g2_fill_2 FILLER_78_321 ();
 sg13g2_fill_1 FILLER_78_323 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_11 ();
 sg13g2_fill_1 FILLER_79_40 ();
 sg13g2_fill_1 FILLER_79_46 ();
 sg13g2_fill_2 FILLER_79_106 ();
 sg13g2_fill_2 FILLER_79_121 ();
 sg13g2_fill_1 FILLER_79_123 ();
 sg13g2_fill_1 FILLER_79_214 ();
 sg13g2_fill_2 FILLER_79_323 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_39 ();
 sg13g2_fill_1 FILLER_80_41 ();
 sg13g2_fill_2 FILLER_80_92 ();
 sg13g2_fill_1 FILLER_80_165 ();
 sg13g2_fill_2 FILLER_80_260 ();
 sg13g2_fill_2 FILLER_80_286 ();
 sg13g2_fill_2 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_390 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net301;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
endmodule

module tt_um_zoom_zoom (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire clknet_leaf_0_clk;
 wire _06992_;
 wire _06993_;
 wire \cpu.ALU.a[0] ;
 wire \cpu.ALU.a[10] ;
 wire \cpu.ALU.a[11] ;
 wire \cpu.ALU.a[12] ;
 wire \cpu.ALU.a[13] ;
 wire \cpu.ALU.a[14] ;
 wire \cpu.ALU.a[15] ;
 wire \cpu.ALU.a[1] ;
 wire \cpu.ALU.a[2] ;
 wire \cpu.ALU.a[3] ;
 wire \cpu.ALU.a[4] ;
 wire \cpu.ALU.a[5] ;
 wire \cpu.ALU.a[6] ;
 wire \cpu.ALU.a[7] ;
 wire \cpu.ALU.a[8] ;
 wire \cpu.ALU.a[9] ;
 wire \cpu.ALU.b[0] ;
 wire \cpu.ALU.b[10] ;
 wire \cpu.ALU.b[11] ;
 wire \cpu.ALU.b[12] ;
 wire \cpu.ALU.b[13] ;
 wire \cpu.ALU.b[14] ;
 wire \cpu.ALU.b[15] ;
 wire \cpu.ALU.b[1] ;
 wire \cpu.ALU.b[2] ;
 wire \cpu.ALU.b[3] ;
 wire \cpu.ALU.b[4] ;
 wire \cpu.ALU.b[5] ;
 wire \cpu.ALU.b[6] ;
 wire \cpu.ALU.b[7] ;
 wire \cpu.ALU.b[8] ;
 wire \cpu.ALU.b[9] ;
 wire \cpu.ALU.mode[0] ;
 wire \cpu.ALU.mode[1] ;
 wire \cpu.ALU.mode[2] ;
 wire \cpu.current_address[0] ;
 wire \cpu.current_address[10] ;
 wire \cpu.current_address[11] ;
 wire \cpu.current_address[12] ;
 wire \cpu.current_address[13] ;
 wire \cpu.current_address[14] ;
 wire \cpu.current_address[15] ;
 wire \cpu.current_address[1] ;
 wire \cpu.current_address[2] ;
 wire \cpu.current_address[3] ;
 wire \cpu.current_address[4] ;
 wire \cpu.current_address[5] ;
 wire \cpu.current_address[6] ;
 wire \cpu.current_address[7] ;
 wire \cpu.current_address[8] ;
 wire \cpu.current_address[9] ;
 wire \cpu.current_instruction[0] ;
 wire \cpu.current_instruction[10] ;
 wire \cpu.current_instruction[11] ;
 wire \cpu.current_instruction[12] ;
 wire \cpu.current_instruction[13] ;
 wire \cpu.current_instruction[14] ;
 wire \cpu.current_instruction[15] ;
 wire \cpu.current_instruction[1] ;
 wire \cpu.current_instruction[2] ;
 wire \cpu.current_instruction[3] ;
 wire \cpu.current_instruction[4] ;
 wire \cpu.current_instruction[5] ;
 wire \cpu.current_instruction[6] ;
 wire \cpu.current_instruction[7] ;
 wire \cpu.current_instruction[8] ;
 wire \cpu.current_instruction[9] ;
 wire \cpu.data_out[0] ;
 wire \cpu.data_out[10] ;
 wire \cpu.data_out[11] ;
 wire \cpu.data_out[12] ;
 wire \cpu.data_out[13] ;
 wire \cpu.data_out[14] ;
 wire \cpu.data_out[15] ;
 wire \cpu.data_out[1] ;
 wire \cpu.data_out[2] ;
 wire \cpu.data_out[3] ;
 wire \cpu.data_out[4] ;
 wire \cpu.data_out[5] ;
 wire \cpu.data_out[6] ;
 wire \cpu.data_out[7] ;
 wire \cpu.data_out[8] ;
 wire \cpu.data_out[9] ;
 wire \cpu.execution_stage[0] ;
 wire \cpu.execution_stage[1] ;
 wire \cpu.execution_stage[2] ;
 wire \cpu.execution_stage[3] ;
 wire \cpu.execution_stage[4] ;
 wire \cpu.execution_stage[5] ;
 wire \cpu.jump_con ;
 wire \cpu.keccak_alu.registers[0] ;
 wire \cpu.keccak_alu.registers[100] ;
 wire \cpu.keccak_alu.registers[101] ;
 wire \cpu.keccak_alu.registers[102] ;
 wire \cpu.keccak_alu.registers[103] ;
 wire \cpu.keccak_alu.registers[104] ;
 wire \cpu.keccak_alu.registers[105] ;
 wire \cpu.keccak_alu.registers[106] ;
 wire \cpu.keccak_alu.registers[107] ;
 wire \cpu.keccak_alu.registers[108] ;
 wire \cpu.keccak_alu.registers[109] ;
 wire \cpu.keccak_alu.registers[10] ;
 wire \cpu.keccak_alu.registers[110] ;
 wire \cpu.keccak_alu.registers[111] ;
 wire \cpu.keccak_alu.registers[112] ;
 wire \cpu.keccak_alu.registers[113] ;
 wire \cpu.keccak_alu.registers[114] ;
 wire \cpu.keccak_alu.registers[115] ;
 wire \cpu.keccak_alu.registers[116] ;
 wire \cpu.keccak_alu.registers[117] ;
 wire \cpu.keccak_alu.registers[118] ;
 wire \cpu.keccak_alu.registers[119] ;
 wire \cpu.keccak_alu.registers[11] ;
 wire \cpu.keccak_alu.registers[120] ;
 wire \cpu.keccak_alu.registers[121] ;
 wire \cpu.keccak_alu.registers[122] ;
 wire \cpu.keccak_alu.registers[123] ;
 wire \cpu.keccak_alu.registers[124] ;
 wire \cpu.keccak_alu.registers[125] ;
 wire \cpu.keccak_alu.registers[126] ;
 wire \cpu.keccak_alu.registers[127] ;
 wire \cpu.keccak_alu.registers[128] ;
 wire \cpu.keccak_alu.registers[129] ;
 wire \cpu.keccak_alu.registers[12] ;
 wire \cpu.keccak_alu.registers[130] ;
 wire \cpu.keccak_alu.registers[131] ;
 wire \cpu.keccak_alu.registers[132] ;
 wire \cpu.keccak_alu.registers[133] ;
 wire \cpu.keccak_alu.registers[134] ;
 wire \cpu.keccak_alu.registers[135] ;
 wire \cpu.keccak_alu.registers[136] ;
 wire \cpu.keccak_alu.registers[137] ;
 wire \cpu.keccak_alu.registers[138] ;
 wire \cpu.keccak_alu.registers[139] ;
 wire \cpu.keccak_alu.registers[13] ;
 wire \cpu.keccak_alu.registers[140] ;
 wire \cpu.keccak_alu.registers[141] ;
 wire \cpu.keccak_alu.registers[142] ;
 wire \cpu.keccak_alu.registers[143] ;
 wire \cpu.keccak_alu.registers[144] ;
 wire \cpu.keccak_alu.registers[145] ;
 wire \cpu.keccak_alu.registers[146] ;
 wire \cpu.keccak_alu.registers[147] ;
 wire \cpu.keccak_alu.registers[148] ;
 wire \cpu.keccak_alu.registers[149] ;
 wire \cpu.keccak_alu.registers[14] ;
 wire \cpu.keccak_alu.registers[150] ;
 wire \cpu.keccak_alu.registers[151] ;
 wire \cpu.keccak_alu.registers[152] ;
 wire \cpu.keccak_alu.registers[153] ;
 wire \cpu.keccak_alu.registers[154] ;
 wire \cpu.keccak_alu.registers[155] ;
 wire \cpu.keccak_alu.registers[156] ;
 wire \cpu.keccak_alu.registers[157] ;
 wire \cpu.keccak_alu.registers[158] ;
 wire \cpu.keccak_alu.registers[159] ;
 wire \cpu.keccak_alu.registers[15] ;
 wire \cpu.keccak_alu.registers[160] ;
 wire \cpu.keccak_alu.registers[161] ;
 wire \cpu.keccak_alu.registers[162] ;
 wire \cpu.keccak_alu.registers[163] ;
 wire \cpu.keccak_alu.registers[164] ;
 wire \cpu.keccak_alu.registers[165] ;
 wire \cpu.keccak_alu.registers[166] ;
 wire \cpu.keccak_alu.registers[167] ;
 wire \cpu.keccak_alu.registers[168] ;
 wire \cpu.keccak_alu.registers[169] ;
 wire \cpu.keccak_alu.registers[16] ;
 wire \cpu.keccak_alu.registers[170] ;
 wire \cpu.keccak_alu.registers[171] ;
 wire \cpu.keccak_alu.registers[172] ;
 wire \cpu.keccak_alu.registers[173] ;
 wire \cpu.keccak_alu.registers[174] ;
 wire \cpu.keccak_alu.registers[175] ;
 wire \cpu.keccak_alu.registers[176] ;
 wire \cpu.keccak_alu.registers[177] ;
 wire \cpu.keccak_alu.registers[178] ;
 wire \cpu.keccak_alu.registers[179] ;
 wire \cpu.keccak_alu.registers[17] ;
 wire \cpu.keccak_alu.registers[180] ;
 wire \cpu.keccak_alu.registers[181] ;
 wire \cpu.keccak_alu.registers[182] ;
 wire \cpu.keccak_alu.registers[183] ;
 wire \cpu.keccak_alu.registers[184] ;
 wire \cpu.keccak_alu.registers[185] ;
 wire \cpu.keccak_alu.registers[186] ;
 wire \cpu.keccak_alu.registers[187] ;
 wire \cpu.keccak_alu.registers[188] ;
 wire \cpu.keccak_alu.registers[189] ;
 wire \cpu.keccak_alu.registers[18] ;
 wire \cpu.keccak_alu.registers[190] ;
 wire \cpu.keccak_alu.registers[191] ;
 wire \cpu.keccak_alu.registers[192] ;
 wire \cpu.keccak_alu.registers[193] ;
 wire \cpu.keccak_alu.registers[194] ;
 wire \cpu.keccak_alu.registers[195] ;
 wire \cpu.keccak_alu.registers[196] ;
 wire \cpu.keccak_alu.registers[197] ;
 wire \cpu.keccak_alu.registers[198] ;
 wire \cpu.keccak_alu.registers[199] ;
 wire \cpu.keccak_alu.registers[19] ;
 wire \cpu.keccak_alu.registers[1] ;
 wire \cpu.keccak_alu.registers[200] ;
 wire \cpu.keccak_alu.registers[201] ;
 wire \cpu.keccak_alu.registers[202] ;
 wire \cpu.keccak_alu.registers[203] ;
 wire \cpu.keccak_alu.registers[204] ;
 wire \cpu.keccak_alu.registers[205] ;
 wire \cpu.keccak_alu.registers[206] ;
 wire \cpu.keccak_alu.registers[207] ;
 wire \cpu.keccak_alu.registers[208] ;
 wire \cpu.keccak_alu.registers[209] ;
 wire \cpu.keccak_alu.registers[20] ;
 wire \cpu.keccak_alu.registers[210] ;
 wire \cpu.keccak_alu.registers[211] ;
 wire \cpu.keccak_alu.registers[212] ;
 wire \cpu.keccak_alu.registers[213] ;
 wire \cpu.keccak_alu.registers[214] ;
 wire \cpu.keccak_alu.registers[215] ;
 wire \cpu.keccak_alu.registers[216] ;
 wire \cpu.keccak_alu.registers[217] ;
 wire \cpu.keccak_alu.registers[218] ;
 wire \cpu.keccak_alu.registers[219] ;
 wire \cpu.keccak_alu.registers[21] ;
 wire \cpu.keccak_alu.registers[220] ;
 wire \cpu.keccak_alu.registers[221] ;
 wire \cpu.keccak_alu.registers[222] ;
 wire \cpu.keccak_alu.registers[223] ;
 wire \cpu.keccak_alu.registers[224] ;
 wire \cpu.keccak_alu.registers[225] ;
 wire \cpu.keccak_alu.registers[226] ;
 wire \cpu.keccak_alu.registers[227] ;
 wire \cpu.keccak_alu.registers[228] ;
 wire \cpu.keccak_alu.registers[229] ;
 wire \cpu.keccak_alu.registers[22] ;
 wire \cpu.keccak_alu.registers[230] ;
 wire \cpu.keccak_alu.registers[231] ;
 wire \cpu.keccak_alu.registers[232] ;
 wire \cpu.keccak_alu.registers[233] ;
 wire \cpu.keccak_alu.registers[234] ;
 wire \cpu.keccak_alu.registers[235] ;
 wire \cpu.keccak_alu.registers[236] ;
 wire \cpu.keccak_alu.registers[237] ;
 wire \cpu.keccak_alu.registers[238] ;
 wire \cpu.keccak_alu.registers[239] ;
 wire \cpu.keccak_alu.registers[23] ;
 wire \cpu.keccak_alu.registers[240] ;
 wire \cpu.keccak_alu.registers[241] ;
 wire \cpu.keccak_alu.registers[242] ;
 wire \cpu.keccak_alu.registers[243] ;
 wire \cpu.keccak_alu.registers[244] ;
 wire \cpu.keccak_alu.registers[245] ;
 wire \cpu.keccak_alu.registers[246] ;
 wire \cpu.keccak_alu.registers[247] ;
 wire \cpu.keccak_alu.registers[248] ;
 wire \cpu.keccak_alu.registers[249] ;
 wire \cpu.keccak_alu.registers[24] ;
 wire \cpu.keccak_alu.registers[250] ;
 wire \cpu.keccak_alu.registers[251] ;
 wire \cpu.keccak_alu.registers[252] ;
 wire \cpu.keccak_alu.registers[253] ;
 wire \cpu.keccak_alu.registers[254] ;
 wire \cpu.keccak_alu.registers[255] ;
 wire \cpu.keccak_alu.registers[256] ;
 wire \cpu.keccak_alu.registers[257] ;
 wire \cpu.keccak_alu.registers[258] ;
 wire \cpu.keccak_alu.registers[259] ;
 wire \cpu.keccak_alu.registers[25] ;
 wire \cpu.keccak_alu.registers[260] ;
 wire \cpu.keccak_alu.registers[261] ;
 wire \cpu.keccak_alu.registers[262] ;
 wire \cpu.keccak_alu.registers[263] ;
 wire \cpu.keccak_alu.registers[264] ;
 wire \cpu.keccak_alu.registers[265] ;
 wire \cpu.keccak_alu.registers[266] ;
 wire \cpu.keccak_alu.registers[267] ;
 wire \cpu.keccak_alu.registers[268] ;
 wire \cpu.keccak_alu.registers[269] ;
 wire \cpu.keccak_alu.registers[26] ;
 wire \cpu.keccak_alu.registers[270] ;
 wire \cpu.keccak_alu.registers[271] ;
 wire \cpu.keccak_alu.registers[272] ;
 wire \cpu.keccak_alu.registers[273] ;
 wire \cpu.keccak_alu.registers[274] ;
 wire \cpu.keccak_alu.registers[275] ;
 wire \cpu.keccak_alu.registers[276] ;
 wire \cpu.keccak_alu.registers[277] ;
 wire \cpu.keccak_alu.registers[278] ;
 wire \cpu.keccak_alu.registers[279] ;
 wire \cpu.keccak_alu.registers[27] ;
 wire \cpu.keccak_alu.registers[280] ;
 wire \cpu.keccak_alu.registers[281] ;
 wire \cpu.keccak_alu.registers[282] ;
 wire \cpu.keccak_alu.registers[283] ;
 wire \cpu.keccak_alu.registers[284] ;
 wire \cpu.keccak_alu.registers[285] ;
 wire \cpu.keccak_alu.registers[286] ;
 wire \cpu.keccak_alu.registers[287] ;
 wire \cpu.keccak_alu.registers[288] ;
 wire \cpu.keccak_alu.registers[289] ;
 wire \cpu.keccak_alu.registers[28] ;
 wire \cpu.keccak_alu.registers[290] ;
 wire \cpu.keccak_alu.registers[291] ;
 wire \cpu.keccak_alu.registers[292] ;
 wire \cpu.keccak_alu.registers[293] ;
 wire \cpu.keccak_alu.registers[294] ;
 wire \cpu.keccak_alu.registers[295] ;
 wire \cpu.keccak_alu.registers[296] ;
 wire \cpu.keccak_alu.registers[297] ;
 wire \cpu.keccak_alu.registers[298] ;
 wire \cpu.keccak_alu.registers[299] ;
 wire \cpu.keccak_alu.registers[29] ;
 wire \cpu.keccak_alu.registers[2] ;
 wire \cpu.keccak_alu.registers[300] ;
 wire \cpu.keccak_alu.registers[301] ;
 wire \cpu.keccak_alu.registers[302] ;
 wire \cpu.keccak_alu.registers[303] ;
 wire \cpu.keccak_alu.registers[304] ;
 wire \cpu.keccak_alu.registers[305] ;
 wire \cpu.keccak_alu.registers[306] ;
 wire \cpu.keccak_alu.registers[307] ;
 wire \cpu.keccak_alu.registers[308] ;
 wire \cpu.keccak_alu.registers[309] ;
 wire \cpu.keccak_alu.registers[30] ;
 wire \cpu.keccak_alu.registers[310] ;
 wire \cpu.keccak_alu.registers[311] ;
 wire \cpu.keccak_alu.registers[312] ;
 wire \cpu.keccak_alu.registers[313] ;
 wire \cpu.keccak_alu.registers[314] ;
 wire \cpu.keccak_alu.registers[315] ;
 wire \cpu.keccak_alu.registers[316] ;
 wire \cpu.keccak_alu.registers[317] ;
 wire \cpu.keccak_alu.registers[318] ;
 wire \cpu.keccak_alu.registers[319] ;
 wire \cpu.keccak_alu.registers[31] ;
 wire \cpu.keccak_alu.registers[32] ;
 wire \cpu.keccak_alu.registers[33] ;
 wire \cpu.keccak_alu.registers[34] ;
 wire \cpu.keccak_alu.registers[35] ;
 wire \cpu.keccak_alu.registers[36] ;
 wire \cpu.keccak_alu.registers[37] ;
 wire \cpu.keccak_alu.registers[38] ;
 wire \cpu.keccak_alu.registers[39] ;
 wire \cpu.keccak_alu.registers[3] ;
 wire \cpu.keccak_alu.registers[40] ;
 wire \cpu.keccak_alu.registers[41] ;
 wire \cpu.keccak_alu.registers[42] ;
 wire \cpu.keccak_alu.registers[43] ;
 wire \cpu.keccak_alu.registers[44] ;
 wire \cpu.keccak_alu.registers[45] ;
 wire \cpu.keccak_alu.registers[46] ;
 wire \cpu.keccak_alu.registers[47] ;
 wire \cpu.keccak_alu.registers[48] ;
 wire \cpu.keccak_alu.registers[49] ;
 wire \cpu.keccak_alu.registers[4] ;
 wire \cpu.keccak_alu.registers[50] ;
 wire \cpu.keccak_alu.registers[51] ;
 wire \cpu.keccak_alu.registers[52] ;
 wire \cpu.keccak_alu.registers[53] ;
 wire \cpu.keccak_alu.registers[54] ;
 wire \cpu.keccak_alu.registers[55] ;
 wire \cpu.keccak_alu.registers[56] ;
 wire \cpu.keccak_alu.registers[57] ;
 wire \cpu.keccak_alu.registers[58] ;
 wire \cpu.keccak_alu.registers[59] ;
 wire \cpu.keccak_alu.registers[5] ;
 wire \cpu.keccak_alu.registers[60] ;
 wire \cpu.keccak_alu.registers[61] ;
 wire \cpu.keccak_alu.registers[62] ;
 wire \cpu.keccak_alu.registers[63] ;
 wire \cpu.keccak_alu.registers[64] ;
 wire \cpu.keccak_alu.registers[65] ;
 wire \cpu.keccak_alu.registers[66] ;
 wire \cpu.keccak_alu.registers[67] ;
 wire \cpu.keccak_alu.registers[68] ;
 wire \cpu.keccak_alu.registers[69] ;
 wire \cpu.keccak_alu.registers[6] ;
 wire \cpu.keccak_alu.registers[70] ;
 wire \cpu.keccak_alu.registers[71] ;
 wire \cpu.keccak_alu.registers[72] ;
 wire \cpu.keccak_alu.registers[73] ;
 wire \cpu.keccak_alu.registers[74] ;
 wire \cpu.keccak_alu.registers[75] ;
 wire \cpu.keccak_alu.registers[76] ;
 wire \cpu.keccak_alu.registers[77] ;
 wire \cpu.keccak_alu.registers[78] ;
 wire \cpu.keccak_alu.registers[79] ;
 wire \cpu.keccak_alu.registers[7] ;
 wire \cpu.keccak_alu.registers[80] ;
 wire \cpu.keccak_alu.registers[81] ;
 wire \cpu.keccak_alu.registers[82] ;
 wire \cpu.keccak_alu.registers[83] ;
 wire \cpu.keccak_alu.registers[84] ;
 wire \cpu.keccak_alu.registers[85] ;
 wire \cpu.keccak_alu.registers[86] ;
 wire \cpu.keccak_alu.registers[87] ;
 wire \cpu.keccak_alu.registers[88] ;
 wire \cpu.keccak_alu.registers[89] ;
 wire \cpu.keccak_alu.registers[8] ;
 wire \cpu.keccak_alu.registers[90] ;
 wire \cpu.keccak_alu.registers[91] ;
 wire \cpu.keccak_alu.registers[92] ;
 wire \cpu.keccak_alu.registers[93] ;
 wire \cpu.keccak_alu.registers[94] ;
 wire \cpu.keccak_alu.registers[95] ;
 wire \cpu.keccak_alu.registers[96] ;
 wire \cpu.keccak_alu.registers[97] ;
 wire \cpu.keccak_alu.registers[98] ;
 wire \cpu.keccak_alu.registers[99] ;
 wire \cpu.keccak_alu.registers[9] ;
 wire \cpu.memory_in[0] ;
 wire \cpu.memory_in[10] ;
 wire \cpu.memory_in[11] ;
 wire \cpu.memory_in[12] ;
 wire \cpu.memory_in[13] ;
 wire \cpu.memory_in[14] ;
 wire \cpu.memory_in[15] ;
 wire \cpu.memory_in[1] ;
 wire \cpu.memory_in[2] ;
 wire \cpu.memory_in[3] ;
 wire \cpu.memory_in[4] ;
 wire \cpu.memory_in[5] ;
 wire \cpu.memory_in[6] ;
 wire \cpu.memory_in[7] ;
 wire \cpu.memory_in[8] ;
 wire \cpu.memory_in[9] ;
 wire \cpu.memory_ready ;
 wire \cpu.registers[1][0] ;
 wire \cpu.registers[1][10] ;
 wire \cpu.registers[1][11] ;
 wire \cpu.registers[1][12] ;
 wire \cpu.registers[1][13] ;
 wire \cpu.registers[1][14] ;
 wire \cpu.registers[1][15] ;
 wire \cpu.registers[1][1] ;
 wire \cpu.registers[1][2] ;
 wire \cpu.registers[1][3] ;
 wire \cpu.registers[1][4] ;
 wire \cpu.registers[1][5] ;
 wire \cpu.registers[1][6] ;
 wire \cpu.registers[1][7] ;
 wire \cpu.registers[1][8] ;
 wire \cpu.registers[1][9] ;
 wire \cpu.registers[2][0] ;
 wire \cpu.registers[2][10] ;
 wire \cpu.registers[2][11] ;
 wire \cpu.registers[2][12] ;
 wire \cpu.registers[2][13] ;
 wire \cpu.registers[2][14] ;
 wire \cpu.registers[2][15] ;
 wire \cpu.registers[2][1] ;
 wire \cpu.registers[2][2] ;
 wire \cpu.registers[2][3] ;
 wire \cpu.registers[2][4] ;
 wire \cpu.registers[2][5] ;
 wire \cpu.registers[2][6] ;
 wire \cpu.registers[2][7] ;
 wire \cpu.registers[2][8] ;
 wire \cpu.registers[2][9] ;
 wire \cpu.registers[3][0] ;
 wire \cpu.registers[3][10] ;
 wire \cpu.registers[3][11] ;
 wire \cpu.registers[3][12] ;
 wire \cpu.registers[3][13] ;
 wire \cpu.registers[3][14] ;
 wire \cpu.registers[3][15] ;
 wire \cpu.registers[3][1] ;
 wire \cpu.registers[3][2] ;
 wire \cpu.registers[3][3] ;
 wire \cpu.registers[3][4] ;
 wire \cpu.registers[3][5] ;
 wire \cpu.registers[3][6] ;
 wire \cpu.registers[3][7] ;
 wire \cpu.registers[3][8] ;
 wire \cpu.registers[3][9] ;
 wire \cpu.registers[4][0] ;
 wire \cpu.registers[4][10] ;
 wire \cpu.registers[4][11] ;
 wire \cpu.registers[4][12] ;
 wire \cpu.registers[4][13] ;
 wire \cpu.registers[4][14] ;
 wire \cpu.registers[4][15] ;
 wire \cpu.registers[4][1] ;
 wire \cpu.registers[4][2] ;
 wire \cpu.registers[4][3] ;
 wire \cpu.registers[4][4] ;
 wire \cpu.registers[4][5] ;
 wire \cpu.registers[4][6] ;
 wire \cpu.registers[4][7] ;
 wire \cpu.registers[4][8] ;
 wire \cpu.registers[4][9] ;
 wire \cpu.registers[5][0] ;
 wire \cpu.registers[5][10] ;
 wire \cpu.registers[5][11] ;
 wire \cpu.registers[5][12] ;
 wire \cpu.registers[5][13] ;
 wire \cpu.registers[5][14] ;
 wire \cpu.registers[5][15] ;
 wire \cpu.registers[5][1] ;
 wire \cpu.registers[5][2] ;
 wire \cpu.registers[5][3] ;
 wire \cpu.registers[5][4] ;
 wire \cpu.registers[5][5] ;
 wire \cpu.registers[5][6] ;
 wire \cpu.registers[5][7] ;
 wire \cpu.registers[5][8] ;
 wire \cpu.registers[5][9] ;
 wire \cpu.registers[6][0] ;
 wire \cpu.registers[6][10] ;
 wire \cpu.registers[6][11] ;
 wire \cpu.registers[6][12] ;
 wire \cpu.registers[6][13] ;
 wire \cpu.registers[6][14] ;
 wire \cpu.registers[6][15] ;
 wire \cpu.registers[6][1] ;
 wire \cpu.registers[6][2] ;
 wire \cpu.registers[6][3] ;
 wire \cpu.registers[6][4] ;
 wire \cpu.registers[6][5] ;
 wire \cpu.registers[6][6] ;
 wire \cpu.registers[6][7] ;
 wire \cpu.registers[6][8] ;
 wire \cpu.registers[6][9] ;
 wire \cpu.registers[7][0] ;
 wire \cpu.registers[7][10] ;
 wire \cpu.registers[7][11] ;
 wire \cpu.registers[7][12] ;
 wire \cpu.registers[7][13] ;
 wire \cpu.registers[7][14] ;
 wire \cpu.registers[7][15] ;
 wire \cpu.registers[7][1] ;
 wire \cpu.registers[7][2] ;
 wire \cpu.registers[7][3] ;
 wire \cpu.registers[7][4] ;
 wire \cpu.registers[7][5] ;
 wire \cpu.registers[7][6] ;
 wire \cpu.registers[7][7] ;
 wire \cpu.registers[7][8] ;
 wire \cpu.registers[7][9] ;
 wire \cpu.request ;
 wire \cpu.request_address[0] ;
 wire \cpu.request_address[10] ;
 wire \cpu.request_address[11] ;
 wire \cpu.request_address[12] ;
 wire \cpu.request_address[13] ;
 wire \cpu.request_address[14] ;
 wire \cpu.request_address[15] ;
 wire \cpu.request_address[1] ;
 wire \cpu.request_address[2] ;
 wire \cpu.request_address[3] ;
 wire \cpu.request_address[4] ;
 wire \cpu.request_address[5] ;
 wire \cpu.request_address[6] ;
 wire \cpu.request_address[7] ;
 wire \cpu.request_address[8] ;
 wire \cpu.request_address[9] ;
 wire \cpu.request_type ;
 wire \cpu.reset ;
 wire \cpu.rx_speed[0] ;
 wire \cpu.rx_speed[10] ;
 wire \cpu.rx_speed[11] ;
 wire \cpu.rx_speed[12] ;
 wire \cpu.rx_speed[1] ;
 wire \cpu.rx_speed[2] ;
 wire \cpu.rx_speed[3] ;
 wire \cpu.rx_speed[4] ;
 wire \cpu.rx_speed[5] ;
 wire \cpu.rx_speed[6] ;
 wire \cpu.rx_speed[7] ;
 wire \cpu.rx_speed[8] ;
 wire \cpu.rx_speed[9] ;
 wire \cpu.set_rx_speed ;
 wire \cpu.tx ;
 wire \cpu.uart.bit_counter[0] ;
 wire \cpu.uart.bit_counter[1] ;
 wire \cpu.uart.bit_counter[2] ;
 wire \cpu.uart.busy ;
 wire \cpu.uart.cycle_counter[0] ;
 wire \cpu.uart.cycle_counter[10] ;
 wire \cpu.uart.cycle_counter[11] ;
 wire \cpu.uart.cycle_counter[12] ;
 wire \cpu.uart.cycle_counter[1] ;
 wire \cpu.uart.cycle_counter[2] ;
 wire \cpu.uart.cycle_counter[3] ;
 wire \cpu.uart.cycle_counter[4] ;
 wire \cpu.uart.cycle_counter[5] ;
 wire \cpu.uart.cycle_counter[6] ;
 wire \cpu.uart.cycle_counter[7] ;
 wire \cpu.uart.cycle_counter[8] ;
 wire \cpu.uart.cycle_counter[9] ;
 wire \cpu.uart.cycles_per_bit[0] ;
 wire \cpu.uart.cycles_per_bit[10] ;
 wire \cpu.uart.cycles_per_bit[11] ;
 wire \cpu.uart.cycles_per_bit[12] ;
 wire \cpu.uart.cycles_per_bit[1] ;
 wire \cpu.uart.cycles_per_bit[2] ;
 wire \cpu.uart.cycles_per_bit[3] ;
 wire \cpu.uart.cycles_per_bit[4] ;
 wire \cpu.uart.cycles_per_bit[5] ;
 wire \cpu.uart.cycles_per_bit[6] ;
 wire \cpu.uart.cycles_per_bit[7] ;
 wire \cpu.uart.cycles_per_bit[8] ;
 wire \cpu.uart.cycles_per_bit[9] ;
 wire \cpu.uart.data_sending[0] ;
 wire \cpu.uart.data_sending[1] ;
 wire \cpu.uart.data_sending[2] ;
 wire \cpu.uart.data_sending[3] ;
 wire \cpu.uart.data_sending[4] ;
 wire \cpu.uart.data_sending[5] ;
 wire \cpu.uart.data_sending[6] ;
 wire \cpu.uart.data_sending[7] ;
 wire \cpu.uart.send ;
 wire \cpu.uart.stage[0] ;
 wire \cpu.uart.stage[1] ;
 wire \cpu.uart.stage[2] ;
 wire \cpu.uart_inbound ;
 wire \cpu.write_complete ;
 wire \data_received[0] ;
 wire \data_received[1] ;
 wire \data_received[2] ;
 wire \data_received[3] ;
 wire \data_received[4] ;
 wire \data_received[5] ;
 wire \data_received[6] ;
 wire \data_received[7] ;
 wire lower_bit;
 wire \memory_controller.next_state[0] ;
 wire \memory_controller.next_state[1] ;
 wire \memory_controller.next_state[2] ;
 wire \memory_controller.next_state[3] ;
 wire \memory_controller.next_state[4] ;
 wire \memory_controller.read_enable ;
 wire \memory_controller.register_enable ;
 wire \memory_controller.state[0] ;
 wire \memory_controller.state[1] ;
 wire \memory_controller.state[2] ;
 wire \memory_controller.state[3] ;
 wire \memory_controller.state[4] ;
 wire \memory_controller.uart_memory_address[10] ;
 wire \memory_controller.upper_bit ;
 wire \memory_controller.wait_counter[0] ;
 wire \memory_controller.wait_counter[1] ;
 wire \memory_controller.wait_counter[2] ;
 wire \memory_controller.wait_counter[3] ;
 wire \memory_controller.wait_counter[4] ;
 wire \memory_controller.wait_counter[5] ;
 wire \memory_controller.write_enable ;
 wire net13;
 wire net14;
 wire \uart_receiver/_000_ ;
 wire \uart_receiver/_001_ ;
 wire \uart_receiver/_002_ ;
 wire \uart_receiver/_003_ ;
 wire \uart_receiver/_004_ ;
 wire \uart_receiver/_005_ ;
 wire \uart_receiver/_006_ ;
 wire \uart_receiver/_007_ ;
 wire \uart_receiver/_008_ ;
 wire \uart_receiver/_009_ ;
 wire \uart_receiver/_010_ ;
 wire \uart_receiver/_011_ ;
 wire \uart_receiver/_012_ ;
 wire \uart_receiver/_013_ ;
 wire \uart_receiver/_014_ ;
 wire \uart_receiver/_015_ ;
 wire \uart_receiver/_016_ ;
 wire \uart_receiver/_017_ ;
 wire \uart_receiver/_018_ ;
 wire \uart_receiver/_019_ ;
 wire \uart_receiver/_020_ ;
 wire \uart_receiver/_021_ ;
 wire \uart_receiver/_022_ ;
 wire \uart_receiver/_023_ ;
 wire \uart_receiver/_024_ ;
 wire \uart_receiver/_025_ ;
 wire \uart_receiver/_026_ ;
 wire \uart_receiver/_027_ ;
 wire \uart_receiver/_028_ ;
 wire \uart_receiver/_029_ ;
 wire \uart_receiver/_030_ ;
 wire \uart_receiver/_031_ ;
 wire \uart_receiver/_032_ ;
 wire \uart_receiver/_033_ ;
 wire \uart_receiver/_034_ ;
 wire \uart_receiver/_035_ ;
 wire \uart_receiver/_036_ ;
 wire \uart_receiver/_037_ ;
 wire \uart_receiver/_038_ ;
 wire \uart_receiver/_039_ ;
 wire \uart_receiver/_040_ ;
 wire \uart_receiver/_041_ ;
 wire \uart_receiver/_042_ ;
 wire \uart_receiver/_043_ ;
 wire \uart_receiver/_044_ ;
 wire \uart_receiver/_045_ ;
 wire \uart_receiver/_046_ ;
 wire \uart_receiver/_047_ ;
 wire \uart_receiver/_048_ ;
 wire \uart_receiver/_049_ ;
 wire \uart_receiver/_050_ ;
 wire \uart_receiver/_051_ ;
 wire \uart_receiver/_052_ ;
 wire \uart_receiver/_053_ ;
 wire \uart_receiver/_054_ ;
 wire \uart_receiver/_055_ ;
 wire \uart_receiver/_056_ ;
 wire \uart_receiver/_057_ ;
 wire \uart_receiver/_058_ ;
 wire \uart_receiver/_059_ ;
 wire \uart_receiver/_060_ ;
 wire \uart_receiver/_061_ ;
 wire \uart_receiver/_062_ ;
 wire \uart_receiver/_063_ ;
 wire \uart_receiver/_064_ ;
 wire \uart_receiver/_065_ ;
 wire \uart_receiver/_066_ ;
 wire \uart_receiver/_067_ ;
 wire \uart_receiver/_068_ ;
 wire \uart_receiver/_069_ ;
 wire \uart_receiver/_070_ ;
 wire \uart_receiver/_071_ ;
 wire \uart_receiver/_072_ ;
 wire \uart_receiver/_073_ ;
 wire \uart_receiver/_074_ ;
 wire \uart_receiver/_075_ ;
 wire \uart_receiver/_076_ ;
 wire \uart_receiver/_077_ ;
 wire \uart_receiver/_078_ ;
 wire \uart_receiver/_079_ ;
 wire \uart_receiver/_080_ ;
 wire \uart_receiver/_081_ ;
 wire \uart_receiver/_082_ ;
 wire \uart_receiver/_083_ ;
 wire \uart_receiver/_084_ ;
 wire \uart_receiver/_085_ ;
 wire \uart_receiver/_086_ ;
 wire \uart_receiver/_087_ ;
 wire \uart_receiver/_088_ ;
 wire \uart_receiver/_089_ ;
 wire \uart_receiver/_090_ ;
 wire \uart_receiver/_091_ ;
 wire \uart_receiver/_092_ ;
 wire \uart_receiver/_093_ ;
 wire \uart_receiver/_094_ ;
 wire \uart_receiver/_095_ ;
 wire \uart_receiver/_096_ ;
 wire \uart_receiver/_097_ ;
 wire \uart_receiver/_098_ ;
 wire \uart_receiver/_099_ ;
 wire \uart_receiver/_100_ ;
 wire \uart_receiver/_101_ ;
 wire \uart_receiver/_102_ ;
 wire \uart_receiver/_103_ ;
 wire \uart_receiver/_104_ ;
 wire \uart_receiver/_105_ ;
 wire \uart_receiver/_106_ ;
 wire \uart_receiver/_107_ ;
 wire \uart_receiver/_108_ ;
 wire \uart_receiver/_109_ ;
 wire \uart_receiver/_110_ ;
 wire \uart_receiver/_111_ ;
 wire \uart_receiver/_112_ ;
 wire \uart_receiver/_113_ ;
 wire \uart_receiver/_114_ ;
 wire \uart_receiver/_115_ ;
 wire \uart_receiver/_116_ ;
 wire \uart_receiver/_117_ ;
 wire \uart_receiver/_118_ ;
 wire \uart_receiver/_119_ ;
 wire \uart_receiver/_120_ ;
 wire \uart_receiver/_121_ ;
 wire \uart_receiver/_122_ ;
 wire \uart_receiver/_123_ ;
 wire \uart_receiver/_124_ ;
 wire \uart_receiver/_125_ ;
 wire \uart_receiver/_126_ ;
 wire \uart_receiver/_127_ ;
 wire \uart_receiver/_128_ ;
 wire \uart_receiver/_129_ ;
 wire \uart_receiver/_130_ ;
 wire \uart_receiver/_131_ ;
 wire \uart_receiver/_132_ ;
 wire \uart_receiver/_133_ ;
 wire \uart_receiver/_134_ ;
 wire \uart_receiver/_135_ ;
 wire \uart_receiver/_136_ ;
 wire \uart_receiver/_137_ ;
 wire \uart_receiver/_138_ ;
 wire \uart_receiver/_139_ ;
 wire \uart_receiver/_140_ ;
 wire \uart_receiver/_141_ ;
 wire \uart_receiver/_142_ ;
 wire \uart_receiver/_143_ ;
 wire \uart_receiver/_144_ ;
 wire \uart_receiver/_145_ ;
 wire \uart_receiver/_146_ ;
 wire \uart_receiver/_147_ ;
 wire \uart_receiver/_148_ ;
 wire \uart_receiver/_149_ ;
 wire \uart_receiver/_150_ ;
 wire \uart_receiver/_151_ ;
 wire \uart_receiver/_152_ ;
 wire \uart_receiver/_153_ ;
 wire \uart_receiver/_154_ ;
 wire \uart_receiver/_155_ ;
 wire \uart_receiver/_156_ ;
 wire \uart_receiver/_157_ ;
 wire \uart_receiver/_158_ ;
 wire \uart_receiver/_159_ ;
 wire \uart_receiver/_160_ ;
 wire \uart_receiver/_161_ ;
 wire \uart_receiver/_162_ ;
 wire \uart_receiver/_163_ ;
 wire \uart_receiver/_164_ ;
 wire \uart_receiver/_165_ ;
 wire \uart_receiver/_166_ ;
 wire \uart_receiver/_167_ ;
 wire \uart_receiver/_168_ ;
 wire \uart_receiver/_169_ ;
 wire \uart_receiver/_170_ ;
 wire \uart_receiver/_171_ ;
 wire \uart_receiver/_172_ ;
 wire \uart_receiver/_173_ ;
 wire \uart_receiver/_174_ ;
 wire \uart_receiver/_175_ ;
 wire \uart_receiver/_176_ ;
 wire \uart_receiver/_177_ ;
 wire \uart_receiver/_178_ ;
 wire \uart_receiver/_179_ ;
 wire \uart_receiver/_180_ ;
 wire \uart_receiver/_181_ ;
 wire \uart_receiver/_182_ ;
 wire \uart_receiver/_183_ ;
 wire \uart_receiver/_184_ ;
 wire \uart_receiver/_185_ ;
 wire \uart_receiver/_186_ ;
 wire \uart_receiver/_187_ ;
 wire \uart_receiver/_188_ ;
 wire \uart_receiver/_189_ ;
 wire \uart_receiver/_190_ ;
 wire \uart_receiver/_191_ ;
 wire \uart_receiver/_192_ ;
 wire \uart_receiver/_193_ ;
 wire \uart_receiver/_194_ ;
 wire \uart_receiver/_195_ ;
 wire \uart_receiver/_196_ ;
 wire \uart_receiver/_197_ ;
 wire \uart_receiver/_198_ ;
 wire \uart_receiver/_199_ ;
 wire \uart_receiver/_200_ ;
 wire \uart_receiver/_201_ ;
 wire \uart_receiver/_202_ ;
 wire \uart_receiver/_203_ ;
 wire \uart_receiver/_204_ ;
 wire \uart_receiver/_205_ ;
 wire \uart_receiver/_206_ ;
 wire \uart_receiver/_207_ ;
 wire \uart_receiver/_208_ ;
 wire \uart_receiver/_209_ ;
 wire \uart_receiver/_210_ ;
 wire \uart_receiver/_211_ ;
 wire \uart_receiver/_212_ ;
 wire \uart_receiver/_213_ ;
 wire \uart_receiver/_214_ ;
 wire \uart_receiver/_215_ ;
 wire \uart_receiver/_216_ ;
 wire \uart_receiver/_217_ ;
 wire \uart_receiver/_218_ ;
 wire \uart_receiver/_219_ ;
 wire \uart_receiver/_220_ ;
 wire \uart_receiver/_221_ ;
 wire \uart_receiver/_222_ ;
 wire \uart_receiver/_223_ ;
 wire \uart_receiver/_224_ ;
 wire \uart_receiver/_225_ ;
 wire \uart_receiver/_226_ ;
 wire \uart_receiver/_227_ ;
 wire \uart_receiver/_228_ ;
 wire \uart_receiver/_229_ ;
 wire \uart_receiver/_230_ ;
 wire \uart_receiver/_231_ ;
 wire \uart_receiver/_232_ ;
 wire \uart_receiver/_233_ ;
 wire \uart_receiver/_234_ ;
 wire \uart_receiver/_235_ ;
 wire \uart_receiver/_236_ ;
 wire \uart_receiver/_237_ ;
 wire \uart_receiver/_238_ ;
 wire \uart_receiver/_239_ ;
 wire \uart_receiver/_240_ ;
 wire \uart_receiver/_241_ ;
 wire \uart_receiver/_242_ ;
 wire \uart_receiver/_243_ ;
 wire \uart_receiver/_244_ ;
 wire \uart_receiver/_245_ ;
 wire \uart_receiver/_246_ ;
 wire \uart_receiver/_247_ ;
 wire \uart_receiver/_248_ ;
 wire \uart_receiver/_249_ ;
 wire \uart_receiver/_250_ ;
 wire \uart_receiver/_251_ ;
 wire \uart_receiver/_252_ ;
 wire \uart_receiver/_253_ ;
 wire \uart_receiver/_254_ ;
 wire \uart_receiver/_255_ ;
 wire \uart_receiver/_256_ ;
 wire \uart_receiver/_257_ ;
 wire \uart_receiver/_258_ ;
 wire \uart_receiver/_259_ ;
 wire \uart_receiver/_260_ ;
 wire \uart_receiver/_261_ ;
 wire \uart_receiver/_262_ ;
 wire \uart_receiver/_263_ ;
 wire \uart_receiver/_264_ ;
 wire \uart_receiver/_265_ ;
 wire \uart_receiver/_266_ ;
 wire \uart_receiver/_267_ ;
 wire \uart_receiver/_268_ ;
 wire \uart_receiver/_269_ ;
 wire \uart_receiver/_270_ ;
 wire \uart_receiver/_271_ ;
 wire \uart_receiver/_272_ ;
 wire \uart_receiver/_273_ ;
 wire \uart_receiver/_274_ ;
 wire \uart_receiver/_275_ ;
 wire \uart_receiver/_276_ ;
 wire \uart_receiver/_277_ ;
 wire \uart_receiver/_278_ ;
 wire \uart_receiver/_279_ ;
 wire \uart_receiver/_280_ ;
 wire \uart_receiver/_281_ ;
 wire \uart_receiver/_282_ ;
 wire \uart_receiver/_283_ ;
 wire \uart_receiver/_284_ ;
 wire \uart_receiver/_285_ ;
 wire \uart_receiver/_286_ ;
 wire \uart_receiver/_287_ ;
 wire \uart_receiver/_288_ ;
 wire \uart_receiver/_289_ ;
 wire \uart_receiver/_290_ ;
 wire \uart_receiver/_291_ ;
 wire \uart_receiver/_292_ ;
 wire \uart_receiver/_293_ ;
 wire \uart_receiver/_294_ ;
 wire \uart_receiver/_295_ ;
 wire \uart_receiver/_296_ ;
 wire \uart_receiver/_297_ ;
 wire \uart_receiver/_298_ ;
 wire \uart_receiver/_299_ ;
 wire \uart_receiver/_300_ ;
 wire \uart_receiver/_301_ ;
 wire \uart_receiver/_302_ ;
 wire \uart_receiver/_303_ ;
 wire \uart_receiver/_304_ ;
 wire \uart_receiver/_305_ ;
 wire \uart_receiver/_306_ ;
 wire \uart_receiver/_307_ ;
 wire \uart_receiver/_308_ ;
 wire \uart_receiver/_309_ ;
 wire \uart_receiver/_310_ ;
 wire \uart_receiver/_311_ ;
 wire \uart_receiver/_312_ ;
 wire \uart_receiver/_313_ ;
 wire \uart_receiver/_314_ ;
 wire \uart_receiver/_315_ ;
 wire \uart_receiver/_316_ ;
 wire \uart_receiver/_317_ ;
 wire \uart_receiver/_318_ ;
 wire \uart_receiver/_319_ ;
 wire \uart_receiver/_320_ ;
 wire \uart_receiver/_321_ ;
 wire \uart_receiver/_322_ ;
 wire \uart_receiver/_323_ ;
 wire \uart_receiver/_324_ ;
 wire \uart_receiver/_325_ ;
 wire \uart_receiver/_326_ ;
 wire \uart_receiver/_327_ ;
 wire \uart_receiver/_328_ ;
 wire \uart_receiver/_329_ ;
 wire \uart_receiver/_330_ ;
 wire \uart_receiver/_331_ ;
 wire \uart_receiver/_332_ ;
 wire \uart_receiver/_333_ ;
 wire \uart_receiver/bit_counter[0] ;
 wire \uart_receiver/bit_counter[1] ;
 wire \uart_receiver/bit_counter[2] ;
 wire \uart_receiver/cycle_counter[0] ;
 wire \uart_receiver/cycle_counter[10] ;
 wire \uart_receiver/cycle_counter[11] ;
 wire \uart_receiver/cycle_counter[12] ;
 wire \uart_receiver/cycle_counter[1] ;
 wire \uart_receiver/cycle_counter[2] ;
 wire \uart_receiver/cycle_counter[3] ;
 wire \uart_receiver/cycle_counter[4] ;
 wire \uart_receiver/cycle_counter[5] ;
 wire \uart_receiver/cycle_counter[6] ;
 wire \uart_receiver/cycle_counter[7] ;
 wire \uart_receiver/cycle_counter[8] ;
 wire \uart_receiver/cycle_counter[9] ;
 wire \uart_receiver/cycles_per_bit[0] ;
 wire \uart_receiver/cycles_per_bit[10] ;
 wire \uart_receiver/cycles_per_bit[11] ;
 wire \uart_receiver/cycles_per_bit[12] ;
 wire \uart_receiver/cycles_per_bit[1] ;
 wire \uart_receiver/cycles_per_bit[2] ;
 wire \uart_receiver/cycles_per_bit[3] ;
 wire \uart_receiver/cycles_per_bit[4] ;
 wire \uart_receiver/cycles_per_bit[5] ;
 wire \uart_receiver/cycles_per_bit[6] ;
 wire \uart_receiver/cycles_per_bit[7] ;
 wire \uart_receiver/cycles_per_bit[8] ;
 wire \uart_receiver/cycles_per_bit[9] ;
 wire \uart_receiver/data[0] ;
 wire \uart_receiver/data[1] ;
 wire \uart_receiver/data[2] ;
 wire \uart_receiver/data[3] ;
 wire \uart_receiver/data[4] ;
 wire \uart_receiver/data[5] ;
 wire \uart_receiver/data[6] ;
 wire \uart_receiver/data[7] ;
 wire \uart_receiver/stage[0] ;
 wire \uart_receiver/stage[1] ;
 wire \uart_receiver/stage[2] ;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;

 sg13g2_inv_1 _06994_ (.Y(_00884_),
    .A(\cpu.uart.stage[1] ));
 sg13g2_inv_2 _06995_ (.Y(_00885_),
    .A(net4314));
 sg13g2_inv_1 _06996_ (.Y(_00886_),
    .A(net4327));
 sg13g2_inv_1 _06997_ (.Y(_00887_),
    .A(net4452));
 sg13g2_inv_2 _06998_ (.Y(_00888_),
    .A(net4302));
 sg13g2_inv_2 _06999_ (.Y(_00889_),
    .A(net4300));
 sg13g2_inv_1 _07000_ (.Y(_00890_),
    .A(_00018_));
 sg13g2_inv_1 _07001_ (.Y(_00891_),
    .A(\memory_controller.state[1] ));
 sg13g2_inv_2 _07002_ (.Y(_00892_),
    .A(net4376));
 sg13g2_inv_1 _07003_ (.Y(_00893_),
    .A(net4368));
 sg13g2_inv_1 _07004_ (.Y(_00894_),
    .A(\cpu.execution_stage[1] ));
 sg13g2_inv_2 _07005_ (.Y(_00895_),
    .A(net4334));
 sg13g2_inv_1 _07006_ (.Y(_00896_),
    .A(_00021_));
 sg13g2_inv_1 _07007_ (.Y(_00897_),
    .A(_00025_));
 sg13g2_inv_1 _07008_ (.Y(_00898_),
    .A(net80));
 sg13g2_inv_1 _07009_ (.Y(_00899_),
    .A(net785));
 sg13g2_inv_1 _07010_ (.Y(_00900_),
    .A(net184));
 sg13g2_inv_1 _07011_ (.Y(_00901_),
    .A(\cpu.uart.cycles_per_bit[5] ));
 sg13g2_inv_1 _07012_ (.Y(_00902_),
    .A(\cpu.uart.cycle_counter[7] ));
 sg13g2_inv_1 _07013_ (.Y(_00903_),
    .A(net229));
 sg13g2_inv_1 _07014_ (.Y(_00904_),
    .A(\cpu.uart.bit_counter[1] ));
 sg13g2_inv_1 _07015_ (.Y(_00905_),
    .A(_00007_));
 sg13g2_inv_4 _07016_ (.A(net4437),
    .Y(_00906_));
 sg13g2_inv_1 _07017_ (.Y(_00907_),
    .A(net619));
 sg13g2_inv_1 _07018_ (.Y(_00908_),
    .A(net50));
 sg13g2_inv_1 _07019_ (.Y(_00909_),
    .A(net160));
 sg13g2_inv_1 _07020_ (.Y(_00910_),
    .A(net422));
 sg13g2_inv_1 _07021_ (.Y(_00911_),
    .A(net432));
 sg13g2_inv_1 _07022_ (.Y(_00912_),
    .A(net534));
 sg13g2_inv_1 _07023_ (.Y(_00913_),
    .A(net56));
 sg13g2_inv_1 _07024_ (.Y(_00914_),
    .A(net162));
 sg13g2_inv_1 _07025_ (.Y(_00915_),
    .A(net447));
 sg13g2_inv_1 _07026_ (.Y(_00916_),
    .A(net200));
 sg13g2_inv_1 _07027_ (.Y(_00917_),
    .A(net485));
 sg13g2_inv_1 _07028_ (.Y(_00918_),
    .A(net321));
 sg13g2_inv_1 _07029_ (.Y(_00919_),
    .A(net491));
 sg13g2_inv_1 _07030_ (.Y(_00920_),
    .A(net47));
 sg13g2_inv_1 _07031_ (.Y(_00921_),
    .A(_00033_));
 sg13g2_inv_1 _07032_ (.Y(_00922_),
    .A(net219));
 sg13g2_inv_1 _07033_ (.Y(_00923_),
    .A(net726));
 sg13g2_inv_1 _07034_ (.Y(_00924_),
    .A(net271));
 sg13g2_inv_1 _07035_ (.Y(_00925_),
    .A(net629));
 sg13g2_inv_1 _07036_ (.Y(_00926_),
    .A(net752));
 sg13g2_inv_1 _07037_ (.Y(_00927_),
    .A(net100));
 sg13g2_inv_1 _07038_ (.Y(_00928_),
    .A(_00034_));
 sg13g2_inv_1 _07039_ (.Y(_00929_),
    .A(net298));
 sg13g2_inv_1 _07040_ (.Y(_00930_),
    .A(net595));
 sg13g2_inv_1 _07041_ (.Y(_00931_),
    .A(net360));
 sg13g2_inv_1 _07042_ (.Y(_00932_),
    .A(net593));
 sg13g2_inv_1 _07043_ (.Y(_00933_),
    .A(net350));
 sg13g2_inv_1 _07044_ (.Y(_00934_),
    .A(net90));
 sg13g2_inv_1 _07045_ (.Y(_00935_),
    .A(_00035_));
 sg13g2_inv_1 _07046_ (.Y(_00936_),
    .A(net364));
 sg13g2_inv_1 _07047_ (.Y(_00937_),
    .A(net508));
 sg13g2_inv_1 _07048_ (.Y(_00938_),
    .A(net292));
 sg13g2_inv_1 _07049_ (.Y(_00939_),
    .A(net500));
 sg13g2_inv_1 _07050_ (.Y(_00940_),
    .A(net570));
 sg13g2_inv_1 _07051_ (.Y(_00941_),
    .A(net239));
 sg13g2_inv_1 _07052_ (.Y(_00942_),
    .A(net93));
 sg13g2_inv_1 _07053_ (.Y(_00943_),
    .A(net583));
 sg13g2_inv_1 _07054_ (.Y(_00944_),
    .A(net471));
 sg13g2_inv_1 _07055_ (.Y(_00945_),
    .A(net250));
 sg13g2_inv_1 _07056_ (.Y(_00946_),
    .A(net475));
 sg13g2_inv_1 _07057_ (.Y(_00947_),
    .A(net626));
 sg13g2_inv_1 _07058_ (.Y(_00948_),
    .A(net255));
 sg13g2_inv_1 _07059_ (.Y(_00949_),
    .A(net95));
 sg13g2_inv_1 _07060_ (.Y(_00950_),
    .A(_00037_));
 sg13g2_inv_1 _07061_ (.Y(_00951_),
    .A(net372));
 sg13g2_inv_1 _07062_ (.Y(_00952_),
    .A(net591));
 sg13g2_inv_1 _07063_ (.Y(_00953_),
    .A(net274));
 sg13g2_inv_1 _07064_ (.Y(_00954_),
    .A(net526));
 sg13g2_inv_1 _07065_ (.Y(_00955_),
    .A(net576));
 sg13g2_inv_1 _07066_ (.Y(_00956_),
    .A(net290));
 sg13g2_inv_1 _07067_ (.Y(_00957_),
    .A(net84));
 sg13g2_inv_1 _07068_ (.Y(_00958_),
    .A(net334));
 sg13g2_inv_1 _07069_ (.Y(_00959_),
    .A(net730));
 sg13g2_inv_1 _07070_ (.Y(_00960_),
    .A(net402));
 sg13g2_inv_1 _07071_ (.Y(_00961_),
    .A(net797));
 sg13g2_inv_1 _07072_ (.Y(_00962_),
    .A(net530));
 sg13g2_inv_1 _07073_ (.Y(_00963_),
    .A(net353));
 sg13g2_inv_1 _07074_ (.Y(_00964_),
    .A(net96));
 sg13g2_inv_1 _07075_ (.Y(_00965_),
    .A(_00039_));
 sg13g2_inv_1 _07076_ (.Y(_00966_),
    .A(net243));
 sg13g2_inv_1 _07077_ (.Y(_00967_),
    .A(net524));
 sg13g2_inv_1 _07078_ (.Y(_00968_),
    .A(net222));
 sg13g2_inv_1 _07079_ (.Y(_00969_),
    .A(net686));
 sg13g2_inv_1 _07080_ (.Y(_00970_),
    .A(net462));
 sg13g2_inv_1 _07081_ (.Y(_00971_),
    .A(net227));
 sg13g2_inv_1 _07082_ (.Y(_00972_),
    .A(net89));
 sg13g2_inv_1 _07083_ (.Y(_00973_),
    .A(_00040_));
 sg13g2_inv_1 _07084_ (.Y(_00974_),
    .A(net482));
 sg13g2_inv_1 _07085_ (.Y(_00975_),
    .A(net771));
 sg13g2_inv_1 _07086_ (.Y(_00976_),
    .A(net312));
 sg13g2_inv_1 _07087_ (.Y(_00977_),
    .A(net703));
 sg13g2_inv_1 _07088_ (.Y(_00978_),
    .A(net480));
 sg13g2_inv_1 _07089_ (.Y(_00979_),
    .A(net302));
 sg13g2_inv_1 _07090_ (.Y(_00980_),
    .A(net106));
 sg13g2_inv_1 _07091_ (.Y(_00981_),
    .A(_00041_));
 sg13g2_inv_1 _07092_ (.Y(_00982_),
    .A(net366));
 sg13g2_inv_1 _07093_ (.Y(_00983_),
    .A(net713));
 sg13g2_inv_1 _07094_ (.Y(_00984_),
    .A(net340));
 sg13g2_inv_1 _07095_ (.Y(_00985_),
    .A(net601));
 sg13g2_inv_1 _07096_ (.Y(_00986_),
    .A(net553));
 sg13g2_inv_1 _07097_ (.Y(_00987_),
    .A(net286));
 sg13g2_inv_1 _07098_ (.Y(_00988_),
    .A(net109));
 sg13g2_inv_1 _07099_ (.Y(_00989_),
    .A(_00042_));
 sg13g2_inv_1 _07100_ (.Y(_00990_),
    .A(net336));
 sg13g2_inv_1 _07101_ (.Y(_00991_),
    .A(net668));
 sg13g2_inv_1 _07102_ (.Y(_00992_),
    .A(net294));
 sg13g2_inv_1 _07103_ (.Y(_00993_),
    .A(net646));
 sg13g2_inv_1 _07104_ (.Y(_00994_),
    .A(net544));
 sg13g2_inv_1 _07105_ (.Y(_00995_),
    .A(net370));
 sg13g2_inv_1 _07106_ (.Y(_00996_),
    .A(net757));
 sg13g2_inv_1 _07107_ (.Y(_00997_),
    .A(net267));
 sg13g2_inv_1 _07108_ (.Y(_00998_),
    .A(net254));
 sg13g2_inv_1 _07109_ (.Y(_00999_),
    .A(net153));
 sg13g2_inv_1 _07110_ (.Y(_01000_),
    .A(net172));
 sg13g2_inv_1 _07111_ (.Y(_01001_),
    .A(\cpu.keccak_alu.registers[1] ));
 sg13g2_inv_1 _07112_ (.Y(_01002_),
    .A(\cpu.keccak_alu.registers[97] ));
 sg13g2_inv_2 _07113_ (.Y(_01003_),
    .A(net4546));
 sg13g2_inv_1 _07114_ (.Y(_01004_),
    .A(\cpu.keccak_alu.registers[145] ));
 sg13g2_inv_1 _07115_ (.Y(_01005_),
    .A(net389));
 sg13g2_inv_1 _07116_ (.Y(_01006_),
    .A(net94));
 sg13g2_inv_1 _07117_ (.Y(_01007_),
    .A(net210));
 sg13g2_inv_1 _07118_ (.Y(_01008_),
    .A(net171));
 sg13g2_inv_1 _07119_ (.Y(_01009_),
    .A(\cpu.keccak_alu.registers[18] ));
 sg13g2_inv_1 _07120_ (.Y(_01010_),
    .A(\cpu.keccak_alu.registers[114] ));
 sg13g2_inv_1 _07121_ (.Y(_01011_),
    .A(net4532));
 sg13g2_inv_1 _07122_ (.Y(_01012_),
    .A(\cpu.keccak_alu.registers[146] ));
 sg13g2_inv_1 _07123_ (.Y(_01013_),
    .A(net282));
 sg13g2_inv_1 _07124_ (.Y(_01014_),
    .A(net231));
 sg13g2_inv_1 _07125_ (.Y(_01015_),
    .A(net193));
 sg13g2_inv_1 _07126_ (.Y(_01016_),
    .A(net132));
 sg13g2_inv_1 _07127_ (.Y(_01017_),
    .A(net685));
 sg13g2_inv_1 _07128_ (.Y(_01018_),
    .A(net719));
 sg13g2_inv_1 _07129_ (.Y(_01019_),
    .A(net4530));
 sg13g2_inv_1 _07130_ (.Y(_01020_),
    .A(\cpu.keccak_alu.registers[163] ));
 sg13g2_inv_2 _07131_ (.Y(_01021_),
    .A(\cpu.keccak_alu.registers[179] ));
 sg13g2_inv_1 _07132_ (.Y(_01022_),
    .A(net453));
 sg13g2_inv_1 _07133_ (.Y(_01023_),
    .A(net116));
 sg13g2_inv_1 _07134_ (.Y(_01024_),
    .A(net108));
 sg13g2_inv_1 _07135_ (.Y(_01025_),
    .A(net180));
 sg13g2_inv_1 _07136_ (.Y(_01026_),
    .A(net624));
 sg13g2_inv_1 _07137_ (.Y(_01027_),
    .A(net600));
 sg13g2_inv_1 _07138_ (.Y(_01028_),
    .A(net4523));
 sg13g2_inv_1 _07139_ (.Y(_01029_),
    .A(net4487));
 sg13g2_inv_1 _07140_ (.Y(_01030_),
    .A(net484));
 sg13g2_inv_1 _07141_ (.Y(_01031_),
    .A(net101));
 sg13g2_inv_1 _07142_ (.Y(_01032_),
    .A(net390));
 sg13g2_inv_1 _07143_ (.Y(_01033_),
    .A(net332));
 sg13g2_inv_1 _07144_ (.Y(_01034_),
    .A(\cpu.keccak_alu.registers[101] ));
 sg13g2_inv_1 _07145_ (.Y(_01035_),
    .A(\cpu.keccak_alu.registers[117] ));
 sg13g2_inv_1 _07146_ (.Y(_01036_),
    .A(net4517));
 sg13g2_inv_1 _07147_ (.Y(_01037_),
    .A(net897));
 sg13g2_inv_1 _07148_ (.Y(_01038_),
    .A(net181));
 sg13g2_inv_1 _07149_ (.Y(_01039_),
    .A(net221));
 sg13g2_inv_1 _07150_ (.Y(_01040_),
    .A(net218));
 sg13g2_inv_1 _07151_ (.Y(_01041_),
    .A(net164));
 sg13g2_inv_1 _07152_ (.Y(_01042_),
    .A(\cpu.keccak_alu.registers[22] ));
 sg13g2_inv_1 _07153_ (.Y(_01043_),
    .A(\cpu.keccak_alu.registers[70] ));
 sg13g2_inv_1 _07154_ (.Y(_01044_),
    .A(\cpu.keccak_alu.registers[102] ));
 sg13g2_inv_1 _07155_ (.Y(_01045_),
    .A(\cpu.keccak_alu.registers[118] ));
 sg13g2_inv_1 _07156_ (.Y(_01046_),
    .A(net4515));
 sg13g2_inv_1 _07157_ (.Y(_01047_),
    .A(net921));
 sg13g2_inv_1 _07158_ (.Y(_01048_),
    .A(net251));
 sg13g2_inv_1 _07159_ (.Y(_01049_),
    .A(net444));
 sg13g2_inv_1 _07160_ (.Y(_01050_),
    .A(net167));
 sg13g2_inv_1 _07161_ (.Y(_01051_),
    .A(net195));
 sg13g2_inv_1 _07162_ (.Y(_01052_),
    .A(net517));
 sg13g2_inv_1 _07163_ (.Y(_01053_),
    .A(\cpu.keccak_alu.registers[103] ));
 sg13g2_inv_1 _07164_ (.Y(_01054_),
    .A(\cpu.keccak_alu.registers[119] ));
 sg13g2_inv_2 _07165_ (.Y(_01055_),
    .A(net604));
 sg13g2_inv_1 _07166_ (.Y(_01056_),
    .A(net942));
 sg13g2_inv_1 _07167_ (.Y(_01057_),
    .A(net156));
 sg13g2_inv_1 _07168_ (.Y(_01058_),
    .A(net556));
 sg13g2_inv_1 _07169_ (.Y(_01059_),
    .A(net276));
 sg13g2_inv_1 _07170_ (.Y(_01060_),
    .A(net173));
 sg13g2_inv_1 _07171_ (.Y(_01061_),
    .A(\cpu.keccak_alu.registers[56] ));
 sg13g2_inv_1 _07172_ (.Y(_01062_),
    .A(\cpu.keccak_alu.registers[72] ));
 sg13g2_inv_1 _07173_ (.Y(_01063_),
    .A(\cpu.keccak_alu.registers[88] ));
 sg13g2_inv_1 _07174_ (.Y(_01064_),
    .A(net4511));
 sg13g2_inv_1 _07175_ (.Y(_01065_),
    .A(\cpu.keccak_alu.registers[184] ));
 sg13g2_inv_1 _07176_ (.Y(_01066_),
    .A(net454));
 sg13g2_inv_1 _07177_ (.Y(_01067_),
    .A(net346));
 sg13g2_inv_1 _07178_ (.Y(_01068_),
    .A(net125));
 sg13g2_inv_1 _07179_ (.Y(_01069_),
    .A(net157));
 sg13g2_inv_1 _07180_ (.Y(_01070_),
    .A(\cpu.keccak_alu.registers[25] ));
 sg13g2_inv_1 _07181_ (.Y(_01071_),
    .A(\cpu.keccak_alu.registers[57] ));
 sg13g2_inv_1 _07182_ (.Y(_01072_),
    .A(\cpu.keccak_alu.registers[73] ));
 sg13g2_inv_1 _07183_ (.Y(_01073_),
    .A(net734));
 sg13g2_inv_1 _07184_ (.Y(_01074_),
    .A(net310));
 sg13g2_inv_1 _07185_ (.Y(_01075_),
    .A(net562));
 sg13g2_inv_1 _07186_ (.Y(_01076_),
    .A(net209));
 sg13g2_inv_1 _07187_ (.Y(_01077_),
    .A(net237));
 sg13g2_inv_1 _07188_ (.Y(_01078_),
    .A(\cpu.keccak_alu.registers[74] ));
 sg13g2_inv_1 _07189_ (.Y(_01079_),
    .A(net261));
 sg13g2_inv_1 _07190_ (.Y(_01080_),
    .A(\cpu.keccak_alu.registers[106] ));
 sg13g2_inv_1 _07191_ (.Y(_01081_),
    .A(net338));
 sg13g2_inv_1 _07192_ (.Y(_01082_),
    .A(net697));
 sg13g2_inv_1 _07193_ (.Y(_01083_),
    .A(net129));
 sg13g2_inv_1 _07194_ (.Y(_01084_),
    .A(net128));
 sg13g2_inv_1 _07195_ (.Y(_01085_),
    .A(\cpu.keccak_alu.registers[27] ));
 sg13g2_inv_1 _07196_ (.Y(_01086_),
    .A(\cpu.keccak_alu.registers[59] ));
 sg13g2_inv_1 _07197_ (.Y(_01087_),
    .A(\cpu.keccak_alu.registers[107] ));
 sg13g2_inv_1 _07198_ (.Y(_01088_),
    .A(\cpu.keccak_alu.registers[139] ));
 sg13g2_inv_1 _07199_ (.Y(_01089_),
    .A(net4484));
 sg13g2_inv_1 _07200_ (.Y(_01090_),
    .A(net283));
 sg13g2_inv_1 _07201_ (.Y(_01091_),
    .A(net499));
 sg13g2_inv_1 _07202_ (.Y(_01092_),
    .A(net144));
 sg13g2_inv_1 _07203_ (.Y(_01093_),
    .A(net152));
 sg13g2_inv_1 _07204_ (.Y(_01094_),
    .A(\cpu.keccak_alu.registers[28] ));
 sg13g2_inv_1 _07205_ (.Y(_01095_),
    .A(\cpu.keccak_alu.registers[76] ));
 sg13g2_inv_1 _07206_ (.Y(_01096_),
    .A(\cpu.keccak_alu.registers[124] ));
 sg13g2_inv_1 _07207_ (.Y(_01097_),
    .A(\cpu.keccak_alu.registers[156] ));
 sg13g2_inv_1 _07208_ (.Y(_01098_),
    .A(net4489));
 sg13g2_inv_1 _07209_ (.Y(_01099_),
    .A(net608));
 sg13g2_inv_1 _07210_ (.Y(_01100_),
    .A(net546));
 sg13g2_inv_1 _07211_ (.Y(_01101_),
    .A(net672));
 sg13g2_inv_1 _07212_ (.Y(_01102_),
    .A(net189));
 sg13g2_inv_1 _07213_ (.Y(_01103_),
    .A(\cpu.keccak_alu.registers[77] ));
 sg13g2_inv_1 _07214_ (.Y(_01104_),
    .A(net408));
 sg13g2_inv_1 _07215_ (.Y(_01105_),
    .A(\cpu.keccak_alu.registers[125] ));
 sg13g2_inv_1 _07216_ (.Y(_01106_),
    .A(\cpu.keccak_alu.registers[189] ));
 sg13g2_inv_1 _07217_ (.Y(_01107_),
    .A(net386));
 sg13g2_inv_1 _07218_ (.Y(_01108_),
    .A(net165));
 sg13g2_inv_1 _07219_ (.Y(_01109_),
    .A(net269));
 sg13g2_inv_1 _07220_ (.Y(_01110_),
    .A(net122));
 sg13g2_inv_1 _07221_ (.Y(_01111_),
    .A(net104));
 sg13g2_inv_1 _07222_ (.Y(_01112_),
    .A(net406));
 sg13g2_inv_1 _07223_ (.Y(_01113_),
    .A(net732));
 sg13g2_inv_1 _07224_ (.Y(_01114_),
    .A(net396));
 sg13g2_inv_1 _07225_ (.Y(_01115_),
    .A(net652));
 sg13g2_inv_1 _07226_ (.Y(_01116_),
    .A(net514));
 sg13g2_inv_1 _07227_ (.Y(_01117_),
    .A(net362));
 sg13g2_inv_1 _07228_ (.Y(_01118_),
    .A(\cpu.keccak_alu.registers[78] ));
 sg13g2_inv_1 _07229_ (.Y(_01119_),
    .A(net425));
 sg13g2_inv_1 _07230_ (.Y(_01120_),
    .A(\cpu.keccak_alu.registers[110] ));
 sg13g2_inv_2 _07231_ (.Y(_01121_),
    .A(\cpu.keccak_alu.registers[158] ));
 sg13g2_inv_1 _07232_ (.Y(_01122_),
    .A(net277));
 sg13g2_inv_1 _07233_ (.Y(_01123_),
    .A(net511));
 sg13g2_inv_1 _07234_ (.Y(_01124_),
    .A(net138));
 sg13g2_inv_1 _07235_ (.Y(_01125_),
    .A(net166));
 sg13g2_inv_1 _07236_ (.Y(_01126_),
    .A(net133));
 sg13g2_inv_1 _07237_ (.Y(_01127_),
    .A(net512));
 sg13g2_inv_1 _07238_ (.Y(_01128_),
    .A(net691));
 sg13g2_inv_1 _07239_ (.Y(_01129_),
    .A(net329));
 sg13g2_inv_1 _07240_ (.Y(_01130_),
    .A(net622));
 sg13g2_inv_1 _07241_ (.Y(_01131_),
    .A(net536));
 sg13g2_inv_1 _07242_ (.Y(_01132_),
    .A(net284));
 sg13g2_inv_1 _07243_ (.Y(_01133_),
    .A(\cpu.keccak_alu.registers[79] ));
 sg13g2_inv_1 _07244_ (.Y(_01134_),
    .A(\cpu.keccak_alu.registers[111] ));
 sg13g2_inv_1 _07245_ (.Y(_01135_),
    .A(net606));
 sg13g2_inv_1 _07246_ (.Y(_01136_),
    .A(net196));
 sg13g2_inv_1 _07247_ (.Y(_01137_),
    .A(net296));
 sg13g2_inv_1 _07248_ (.Y(_01138_),
    .A(net431));
 sg13g2_inv_1 _07249_ (.Y(_01139_),
    .A(net126));
 sg13g2_inv_1 _07250_ (.Y(_01140_),
    .A(net439));
 sg13g2_inv_1 _07251_ (.Y(_01141_),
    .A(net656));
 sg13g2_inv_1 _07252_ (.Y(_01142_),
    .A(net399));
 sg13g2_inv_1 _07253_ (.Y(_01143_),
    .A(net711));
 sg13g2_inv_1 _07254_ (.Y(_01144_),
    .A(net326));
 sg13g2_inv_1 _07255_ (.Y(_01145_),
    .A(net445));
 sg13g2_inv_1 _07256_ (.Y(_01146_),
    .A(net875));
 sg13g2_inv_1 _07257_ (.Y(_01147_),
    .A(\cpu.request_address[3] ));
 sg13g2_inv_1 _07258_ (.Y(_01148_),
    .A(net913));
 sg13g2_inv_1 _07259_ (.Y(_01149_),
    .A(net904));
 sg13g2_inv_1 _07260_ (.Y(_01150_),
    .A(net929));
 sg13g2_inv_1 _07261_ (.Y(_01151_),
    .A(net541));
 sg13g2_inv_1 _07262_ (.Y(_01152_),
    .A(net877));
 sg13g2_inv_1 _07263_ (.Y(_01153_),
    .A(net235));
 sg13g2_inv_1 _07264_ (.Y(_01154_),
    .A(net743));
 sg13g2_inv_1 _07265_ (.Y(_01155_),
    .A(net355));
 sg13g2_inv_1 _07266_ (.Y(_01156_),
    .A(net717));
 sg13g2_inv_1 _07267_ (.Y(_01157_),
    .A(net319));
 sg13g2_inv_1 _07268_ (.Y(_01158_),
    .A(net584));
 sg13g2_inv_1 _07269_ (.Y(_01159_),
    .A(net317));
 sg13g2_inv_1 _07270_ (.Y(_01160_),
    .A(net611));
 sg13g2_inv_1 _07271_ (.Y(_01161_),
    .A(net324));
 sg13g2_inv_1 _07272_ (.Y(_01162_),
    .A(net763));
 sg13g2_inv_1 _07273_ (.Y(_01163_),
    .A(net805));
 sg13g2_inv_1 _07274_ (.Y(_01164_),
    .A(net470));
 sg13g2_inv_1 _07275_ (.Y(_01165_),
    .A(net357));
 sg13g2_inv_2 _07276_ (.Y(_01166_),
    .A(_00067_));
 sg13g2_inv_2 _07277_ (.Y(_01167_),
    .A(_00072_));
 sg13g2_inv_2 _07278_ (.Y(_01168_),
    .A(_00116_));
 sg13g2_inv_1 _07279_ (.Y(_01169_),
    .A(net4576));
 sg13g2_inv_4 _07280_ (.A(net4363),
    .Y(_01170_));
 sg13g2_inv_4 _07281_ (.A(net4351),
    .Y(_01171_));
 sg13g2_inv_1 _07282_ (.Y(_01172_),
    .A(net4348));
 sg13g2_inv_4 _07283_ (.A(net4344),
    .Y(_01173_));
 sg13g2_inv_1 _07284_ (.Y(_01174_),
    .A(net4339));
 sg13g2_inv_4 _07285_ (.A(net4338),
    .Y(_01175_));
 sg13g2_inv_2 _07286_ (.Y(_01176_),
    .A(net4293));
 sg13g2_inv_2 _07287_ (.Y(_01177_),
    .A(net4287));
 sg13g2_inv_2 _07288_ (.Y(_01178_),
    .A(net4275));
 sg13g2_inv_2 _07289_ (.Y(_01179_),
    .A(net4273));
 sg13g2_inv_1 _07290_ (.Y(_01180_),
    .A(\cpu.ALU.mode[0] ));
 sg13g2_inv_1 _07291_ (.Y(_01181_),
    .A(_00152_));
 sg13g2_inv_1 _07292_ (.Y(_01182_),
    .A(_00160_));
 sg13g2_inv_1 _07293_ (.Y(_01183_),
    .A(_00180_));
 sg13g2_inv_1 _07294_ (.Y(_01184_),
    .A(\cpu.ALU.b[9] ));
 sg13g2_inv_1 _07295_ (.Y(_01185_),
    .A(\cpu.ALU.a[11] ));
 sg13g2_inv_1 _07296_ (.Y(_01186_),
    .A(_00189_));
 sg13g2_inv_1 _07297_ (.Y(_01187_),
    .A(_00192_));
 sg13g2_inv_1 _07298_ (.Y(_01188_),
    .A(\cpu.ALU.a[12] ));
 sg13g2_inv_1 _07299_ (.Y(_01189_),
    .A(_00193_));
 sg13g2_inv_1 _07300_ (.Y(_01190_),
    .A(_00196_));
 sg13g2_inv_1 _07301_ (.Y(_01191_),
    .A(\cpu.ALU.a[15] ));
 sg13g2_inv_4 _07302_ (.A(net4630),
    .Y(\cpu.reset ));
 sg13g2_inv_1 _07303_ (.Y(_01192_),
    .A(net23));
 sg13g2_inv_1 _07304_ (.Y(_01193_),
    .A(net20));
 sg13g2_inv_1 _07305_ (.Y(_01194_),
    .A(net22));
 sg13g2_inv_1 _07306_ (.Y(_01195_),
    .A(net21));
 sg13g2_nand2b_1 _07307_ (.Y(_01196_),
    .B(\cpu.uart.send ),
    .A_N(net4475));
 sg13g2_xnor2_1 _07308_ (.Y(_01197_),
    .A(\cpu.uart.cycles_per_bit[1] ),
    .B(\cpu.uart.cycle_counter[1] ));
 sg13g2_nand2b_1 _07309_ (.Y(_01198_),
    .B(\cpu.uart.cycles_per_bit[0] ),
    .A_N(\cpu.uart.cycle_counter[0] ));
 sg13g2_nor2b_1 _07310_ (.A(\cpu.uart.cycle_counter[9] ),
    .B_N(\cpu.uart.cycles_per_bit[9] ),
    .Y(_01199_));
 sg13g2_nand2b_1 _07311_ (.Y(_01200_),
    .B(\cpu.uart.cycles_per_bit[8] ),
    .A_N(\cpu.uart.cycle_counter[8] ));
 sg13g2_xnor2_1 _07312_ (.Y(_01201_),
    .A(\cpu.uart.cycles_per_bit[12] ),
    .B(\cpu.uart.cycle_counter[12] ));
 sg13g2_nor2b_1 _07313_ (.A(\cpu.uart.cycle_counter[2] ),
    .B_N(\cpu.uart.cycles_per_bit[2] ),
    .Y(_01202_));
 sg13g2_nand2b_1 _07314_ (.Y(_01203_),
    .B(\cpu.uart.cycle_counter[2] ),
    .A_N(\cpu.uart.cycles_per_bit[2] ));
 sg13g2_nand2b_1 _07315_ (.Y(_01204_),
    .B(\cpu.uart.cycle_counter[9] ),
    .A_N(\cpu.uart.cycles_per_bit[9] ));
 sg13g2_nand2b_1 _07316_ (.Y(_01205_),
    .B(\cpu.uart.cycle_counter[6] ),
    .A_N(\cpu.uart.cycles_per_bit[6] ));
 sg13g2_nor2b_1 _07317_ (.A(\cpu.uart.cycle_counter[6] ),
    .B_N(\cpu.uart.cycles_per_bit[6] ),
    .Y(_01206_));
 sg13g2_nand3_1 _07318_ (.B(_01201_),
    .C(_01205_),
    .A(_01198_),
    .Y(_01207_));
 sg13g2_a22oi_1 _07319_ (.Y(_01208_),
    .B1(_00903_),
    .B2(\cpu.uart.cycle_counter[8] ),
    .A2(_00902_),
    .A1(\cpu.uart.cycles_per_bit[7] ));
 sg13g2_xnor2_1 _07320_ (.Y(_01209_),
    .A(\cpu.uart.cycles_per_bit[10] ),
    .B(\cpu.uart.cycle_counter[10] ));
 sg13g2_xnor2_1 _07321_ (.Y(_01210_),
    .A(\cpu.uart.cycles_per_bit[4] ),
    .B(\cpu.uart.cycle_counter[4] ));
 sg13g2_nand4_1 _07322_ (.B(_01208_),
    .C(_01209_),
    .A(_01200_),
    .Y(_01211_),
    .D(_01210_));
 sg13g2_nor4_1 _07323_ (.A(_01199_),
    .B(_01206_),
    .C(_01207_),
    .D(_01211_),
    .Y(_01212_));
 sg13g2_o21ai_1 _07324_ (.B1(_01203_),
    .Y(_01213_),
    .A1(\cpu.uart.cycles_per_bit[7] ),
    .A2(_00902_));
 sg13g2_xor2_1 _07325_ (.B(\cpu.uart.cycle_counter[11] ),
    .A(\cpu.uart.cycles_per_bit[11] ),
    .X(_01214_));
 sg13g2_o21ai_1 _07326_ (.B1(_01204_),
    .Y(_01215_),
    .A1(_00901_),
    .A2(\cpu.uart.cycle_counter[5] ));
 sg13g2_nor4_1 _07327_ (.A(_01202_),
    .B(_01213_),
    .C(_01214_),
    .D(_01215_),
    .Y(_01216_));
 sg13g2_xor2_1 _07328_ (.B(\cpu.uart.cycle_counter[3] ),
    .A(\cpu.uart.cycles_per_bit[3] ),
    .X(_01217_));
 sg13g2_a221oi_1 _07329_ (.B2(\cpu.uart.cycle_counter[5] ),
    .C1(_01217_),
    .B1(_00901_),
    .A1(_00900_),
    .Y(_01218_),
    .A2(\cpu.uart.cycle_counter[0] ));
 sg13g2_nand4_1 _07330_ (.B(_01212_),
    .C(_01216_),
    .A(_01197_),
    .Y(_01219_),
    .D(_01218_));
 sg13g2_nor2_1 _07331_ (.A(\cpu.uart.bit_counter[1] ),
    .B(net4267),
    .Y(_01220_));
 sg13g2_nand2_1 _07332_ (.Y(_01221_),
    .A(_00029_),
    .B(_01220_));
 sg13g2_inv_1 _07333_ (.Y(_01222_),
    .A(_01221_));
 sg13g2_nor4_1 _07334_ (.A(_00884_),
    .B(net4477),
    .C(_01219_),
    .D(_01221_),
    .Y(_01223_));
 sg13g2_a21oi_1 _07335_ (.A1(net30),
    .A2(_01196_),
    .Y(_00262_),
    .B1(_01223_));
 sg13g2_a21oi_1 _07336_ (.A1(net4243),
    .A2(net45),
    .Y(_00261_),
    .B1(\cpu.execution_stage[1] ));
 sg13g2_nand2b_2 _07337_ (.Y(_01224_),
    .B(\cpu.current_instruction[2] ),
    .A_N(\cpu.current_instruction[3] ));
 sg13g2_nor2_2 _07338_ (.A(\cpu.current_instruction[1] ),
    .B(_01224_),
    .Y(_01225_));
 sg13g2_nand2b_2 _07339_ (.Y(_01226_),
    .B(\cpu.current_instruction[1] ),
    .A_N(\cpu.current_instruction[0] ));
 sg13g2_nor2_2 _07340_ (.A(_01224_),
    .B(_01226_),
    .Y(_01227_));
 sg13g2_or2_1 _07341_ (.X(_01228_),
    .B(_01226_),
    .A(_01224_));
 sg13g2_nand2b_2 _07342_ (.Y(_01229_),
    .B(\cpu.current_instruction[0] ),
    .A_N(\cpu.current_instruction[1] ));
 sg13g2_nand2b_2 _07343_ (.Y(_01230_),
    .B(net208),
    .A_N(\cpu.current_instruction[2] ));
 sg13g2_nor2_2 _07344_ (.A(_01229_),
    .B(_01230_),
    .Y(_01231_));
 sg13g2_or2_1 _07345_ (.X(_01232_),
    .B(_01230_),
    .A(_01229_));
 sg13g2_nand2_2 _07346_ (.Y(_01233_),
    .A(net4078),
    .B(net4071));
 sg13g2_nor2_1 _07347_ (.A(_01225_),
    .B(_01233_),
    .Y(_01234_));
 sg13g2_nor3_2 _07348_ (.A(\cpu.current_instruction[0] ),
    .B(\cpu.current_instruction[1] ),
    .C(_01224_),
    .Y(_01235_));
 sg13g2_nand2_1 _07349_ (.Y(_01236_),
    .A(net4448),
    .B(\cpu.current_instruction[6] ));
 sg13g2_nor2_1 _07350_ (.A(net4450),
    .B(_01236_),
    .Y(_01237_));
 sg13g2_nand2b_1 _07351_ (.Y(_01238_),
    .B(net4239),
    .A_N(_01236_));
 sg13g2_nand2_1 _07352_ (.Y(_01239_),
    .A(_01235_),
    .B(net4065));
 sg13g2_nor2b_1 _07353_ (.A(_01234_),
    .B_N(net4306),
    .Y(_01240_));
 sg13g2_nand2_1 _07354_ (.Y(_01241_),
    .A(_01226_),
    .B(_01229_));
 sg13g2_nor2_1 _07355_ (.A(_01224_),
    .B(_01229_),
    .Y(_01242_));
 sg13g2_nand2_1 _07356_ (.Y(_01243_),
    .A(\cpu.current_instruction[0] ),
    .B(_01225_));
 sg13g2_nand2_2 _07357_ (.Y(_01244_),
    .A(net4079),
    .B(net3866));
 sg13g2_nand2_1 _07358_ (.Y(_01245_),
    .A(net4326),
    .B(net4239));
 sg13g2_nor2_1 _07359_ (.A(net4257),
    .B(_01245_),
    .Y(_01246_));
 sg13g2_nand2_2 _07360_ (.Y(_01247_),
    .A(net4238),
    .B(net4050));
 sg13g2_a221oi_1 _07361_ (.B2(_01246_),
    .C1(net809),
    .B1(_01244_),
    .A1(_01239_),
    .Y(_00260_),
    .A2(_01240_));
 sg13g2_nor2_1 _07362_ (.A(net4239),
    .B(net3865),
    .Y(_01248_));
 sg13g2_nand2_2 _07363_ (.Y(_01249_),
    .A(net4451),
    .B(net4049));
 sg13g2_nand2_2 _07364_ (.Y(_01250_),
    .A(net4217),
    .B(net4208));
 sg13g2_nor2_2 _07365_ (.A(net4071),
    .B(_01250_),
    .Y(_01251_));
 sg13g2_a21oi_1 _07366_ (.A1(_01235_),
    .A2(_01237_),
    .Y(_01252_),
    .B1(_01251_));
 sg13g2_a21oi_1 _07367_ (.A1(_01249_),
    .A2(_01252_),
    .Y(_01253_),
    .B1(_00022_));
 sg13g2_a22oi_1 _07368_ (.Y(_01254_),
    .B1(net4074),
    .B2(_01250_),
    .A2(_01227_),
    .A1(net4450));
 sg13g2_or2_1 _07369_ (.X(_01255_),
    .B(net3861),
    .A(_00020_));
 sg13g2_or2_2 _07370_ (.X(_01256_),
    .B(\cpu.current_instruction[2] ),
    .A(\cpu.current_instruction[3] ));
 sg13g2_nor2_2 _07371_ (.A(_01229_),
    .B(_01256_),
    .Y(_01257_));
 sg13g2_nor2_1 _07372_ (.A(_01226_),
    .B(_01256_),
    .Y(_01258_));
 sg13g2_or2_1 _07373_ (.X(_01259_),
    .B(_01256_),
    .A(_01226_));
 sg13g2_nor2_2 _07374_ (.A(_01257_),
    .B(net4038),
    .Y(_01260_));
 sg13g2_nand3_1 _07375_ (.B(_01255_),
    .C(_01260_),
    .A(_01239_),
    .Y(_01261_));
 sg13g2_o21ai_1 _07376_ (.B1(net4316),
    .Y(_01262_),
    .A1(_01253_),
    .A2(_01261_));
 sg13g2_nand2_2 _07377_ (.Y(_01263_),
    .A(\cpu.current_instruction[0] ),
    .B(\cpu.current_instruction[1] ));
 sg13g2_nor2_2 _07378_ (.A(_01224_),
    .B(_01263_),
    .Y(_01264_));
 sg13g2_or2_1 _07379_ (.X(_01265_),
    .B(_01263_),
    .A(_01224_));
 sg13g2_o21ai_1 _07380_ (.B1(net4032),
    .Y(_01266_),
    .A1(_01241_),
    .A2(_01256_));
 sg13g2_nor3_2 _07381_ (.A(\cpu.current_instruction[0] ),
    .B(\cpu.current_instruction[1] ),
    .C(_01230_),
    .Y(_01267_));
 sg13g2_nand2_1 _07382_ (.Y(_01268_),
    .A(net4311),
    .B(_01267_));
 sg13g2_nand3_1 _07383_ (.B(net933),
    .C(_01267_),
    .A(net4311),
    .Y(_01269_));
 sg13g2_nand2_1 _07384_ (.Y(_01270_),
    .A(net4325),
    .B(net4051));
 sg13g2_o21ai_1 _07385_ (.B1(_01270_),
    .Y(_01271_),
    .A1(_00020_),
    .A2(net4053));
 sg13g2_a22oi_1 _07386_ (.Y(_01272_),
    .B1(_01271_),
    .B2(net4301),
    .A2(_01266_),
    .A1(net4306));
 sg13g2_nand3_1 _07387_ (.B(_01269_),
    .C(_01272_),
    .A(_01262_),
    .Y(_00001_));
 sg13g2_nand2b_1 _07388_ (.Y(_01273_),
    .B(_01260_),
    .A_N(_01233_));
 sg13g2_o21ai_1 _07389_ (.B1(net4306),
    .Y(_01274_),
    .A1(_01225_),
    .A2(_01273_));
 sg13g2_nand2_1 _07390_ (.Y(_01275_),
    .A(_00017_),
    .B(_01227_));
 sg13g2_nand2b_1 _07391_ (.Y(_01276_),
    .B(_01275_),
    .A_N(_01251_));
 sg13g2_a21oi_1 _07392_ (.A1(_01252_),
    .A2(_01275_),
    .Y(_01277_),
    .B1(net4326));
 sg13g2_a22oi_1 _07393_ (.Y(_01278_),
    .B1(_01260_),
    .B2(_01234_),
    .A2(net4053),
    .A1(_00022_));
 sg13g2_o21ai_1 _07394_ (.B1(_01278_),
    .Y(_01279_),
    .A1(net4335),
    .A2(net3860));
 sg13g2_o21ai_1 _07395_ (.B1(net4316),
    .Y(_01280_),
    .A1(_01277_),
    .A2(_01279_));
 sg13g2_nand2_1 _07396_ (.Y(_00002_),
    .A(_01274_),
    .B(_01280_));
 sg13g2_nand3b_1 _07397_ (.B(net30),
    .C(\cpu.uart.send ),
    .Y(_01281_),
    .A_N(net4475));
 sg13g2_nand2_1 _07398_ (.Y(_01282_),
    .A(\cpu.uart.bit_counter[1] ),
    .B(net4267));
 sg13g2_nand3_1 _07399_ (.B(net4267),
    .C(net580),
    .A(\cpu.uart.bit_counter[1] ),
    .Y(_01283_));
 sg13g2_nor3_1 _07400_ (.A(net4477),
    .B(_01219_),
    .C(_01283_),
    .Y(_01284_));
 sg13g2_o21ai_1 _07401_ (.B1(net4150),
    .Y(_00006_),
    .A1(_00899_),
    .A2(_01284_));
 sg13g2_nand2_1 _07402_ (.Y(_01285_),
    .A(net817),
    .B(_01219_));
 sg13g2_o21ai_1 _07403_ (.B1(net817),
    .Y(_01286_),
    .A1(net4477),
    .A2(_01221_));
 sg13g2_nand2_1 _07404_ (.Y(_01287_),
    .A(net785),
    .B(_01284_));
 sg13g2_nand3_1 _07405_ (.B(_01286_),
    .C(_01287_),
    .A(_01285_),
    .Y(_00005_));
 sg13g2_nand2b_2 _07406_ (.Y(_01288_),
    .B(net4317),
    .A_N(_00022_));
 sg13g2_nand2_1 _07407_ (.Y(_01289_),
    .A(net831),
    .B(_01244_));
 sg13g2_nor2_2 _07408_ (.A(net4236),
    .B(net4055),
    .Y(_01290_));
 sg13g2_nand2_1 _07409_ (.Y(_01291_),
    .A(net4301),
    .B(net3866));
 sg13g2_nor2_1 _07410_ (.A(net4233),
    .B(net3865),
    .Y(_01292_));
 sg13g2_nand2_1 _07411_ (.Y(_01293_),
    .A(net4301),
    .B(net4051));
 sg13g2_a22oi_1 _07412_ (.Y(_01294_),
    .B1(_01292_),
    .B2(_00022_),
    .A2(_01290_),
    .A1(net4205));
 sg13g2_o21ai_1 _07413_ (.B1(_01294_),
    .Y(_00004_),
    .A1(_01288_),
    .A2(_01289_));
 sg13g2_nor2b_1 _07414_ (.A(_01267_),
    .B_N(net4306),
    .Y(_01295_));
 sg13g2_nand4_1 _07415_ (.B(_01256_),
    .C(net4033),
    .A(_01234_),
    .Y(_01296_),
    .D(_01295_));
 sg13g2_nand3_1 _07416_ (.B(net342),
    .C(_01267_),
    .A(net4310),
    .Y(_01297_));
 sg13g2_nand3_1 _07417_ (.B(_01296_),
    .C(_01297_),
    .A(_00888_),
    .Y(_00003_));
 sg13g2_nor2b_1 _07418_ (.A(\memory_controller.state[3] ),
    .B_N(\memory_controller.state[2] ),
    .Y(_01298_));
 sg13g2_nand2_2 _07419_ (.Y(_01299_),
    .A(net4331),
    .B(_01298_));
 sg13g2_nor2_1 _07420_ (.A(net4333),
    .B(_01299_),
    .Y(_01300_));
 sg13g2_nor2_2 _07421_ (.A(\memory_controller.state[3] ),
    .B(\memory_controller.state[2] ),
    .Y(_01301_));
 sg13g2_nand2b_2 _07422_ (.Y(_01302_),
    .B(\memory_controller.state[1] ),
    .A_N(net4333));
 sg13g2_nand3b_1 _07423_ (.B(_01301_),
    .C(\memory_controller.state[1] ),
    .Y(_01303_),
    .A_N(net4333));
 sg13g2_nor2_1 _07424_ (.A(net4332),
    .B(_01303_),
    .Y(_01304_));
 sg13g2_nor2b_2 _07425_ (.A(\memory_controller.state[2] ),
    .B_N(\memory_controller.state[3] ),
    .Y(_01305_));
 sg13g2_nand2_2 _07426_ (.Y(_01306_),
    .A(net4331),
    .B(_01305_));
 sg13g2_nor2_2 _07427_ (.A(\memory_controller.state[1] ),
    .B(net4333),
    .Y(_01307_));
 sg13g2_nor2b_1 _07428_ (.A(_01306_),
    .B_N(_01307_),
    .Y(_01308_));
 sg13g2_nor3_1 _07429_ (.A(_01300_),
    .B(_01304_),
    .C(_01308_),
    .Y(_01309_));
 sg13g2_nor2b_1 _07430_ (.A(\memory_controller.state[1] ),
    .B_N(net4333),
    .Y(_01310_));
 sg13g2_nand2_2 _07431_ (.Y(_01311_),
    .A(_00891_),
    .B(\memory_controller.state[0] ));
 sg13g2_nand2_2 _07432_ (.Y(_01312_),
    .A(net4332),
    .B(_01298_));
 sg13g2_nand3_1 _07433_ (.B(\memory_controller.state[2] ),
    .C(net4331),
    .A(\memory_controller.state[3] ),
    .Y(_01313_));
 sg13g2_a21oi_1 _07434_ (.A1(_01312_),
    .A2(_01313_),
    .Y(_01314_),
    .B1(_01311_));
 sg13g2_nand2_1 _07435_ (.Y(_01315_),
    .A(net4332),
    .B(_01305_));
 sg13g2_nor2_2 _07436_ (.A(_01311_),
    .B(_01315_),
    .Y(_01316_));
 sg13g2_nand3_1 _07437_ (.B(_01305_),
    .C(_01310_),
    .A(net4332),
    .Y(_01317_));
 sg13g2_and2_1 _07438_ (.A(\memory_controller.state[1] ),
    .B(net4333),
    .X(_01318_));
 sg13g2_nand2_2 _07439_ (.Y(_01319_),
    .A(\memory_controller.state[1] ),
    .B(net4333));
 sg13g2_nor2_2 _07440_ (.A(_01312_),
    .B(_01319_),
    .Y(_01320_));
 sg13g2_nor2_1 _07441_ (.A(_01316_),
    .B(_01320_),
    .Y(_01321_));
 sg13g2_nor2_1 _07442_ (.A(_01306_),
    .B(_01319_),
    .Y(_01322_));
 sg13g2_nor4_1 _07443_ (.A(_01314_),
    .B(_01316_),
    .C(_01320_),
    .D(_01322_),
    .Y(_01323_));
 sg13g2_and2_2 _07444_ (.A(_01309_),
    .B(_01323_),
    .X(_01324_));
 sg13g2_nor2_1 _07445_ (.A(net55),
    .B(_01324_),
    .Y(_00010_));
 sg13g2_xnor2_1 _07446_ (.Y(_01325_),
    .A(net450),
    .B(net55));
 sg13g2_nor2_1 _07447_ (.A(_01324_),
    .B(_01325_),
    .Y(_00011_));
 sg13g2_and3_1 _07448_ (.X(_01326_),
    .A(net168),
    .B(\memory_controller.wait_counter[1] ),
    .C(net55));
 sg13g2_a21oi_1 _07449_ (.A1(\memory_controller.wait_counter[1] ),
    .A2(net55),
    .Y(_01327_),
    .B1(net168));
 sg13g2_nor3_1 _07450_ (.A(_01324_),
    .B(_01326_),
    .C(net169),
    .Y(_00012_));
 sg13g2_and2_1 _07451_ (.A(net379),
    .B(_01326_),
    .X(_01328_));
 sg13g2_nor2_1 _07452_ (.A(net379),
    .B(_01326_),
    .Y(_01329_));
 sg13g2_nor3_1 _07453_ (.A(_01324_),
    .B(_01328_),
    .C(net380),
    .Y(_00013_));
 sg13g2_nand2_1 _07454_ (.Y(_01330_),
    .A(net566),
    .B(_01328_));
 sg13g2_xnor2_1 _07455_ (.Y(_01331_),
    .A(net566),
    .B(_01328_));
 sg13g2_nor2_1 _07456_ (.A(_01324_),
    .B(_01331_),
    .Y(_00014_));
 sg13g2_xor2_1 _07457_ (.B(_01330_),
    .A(net667),
    .X(_01332_));
 sg13g2_nor2_1 _07458_ (.A(_01324_),
    .B(_01332_),
    .Y(_00015_));
 sg13g2_nor2_1 _07459_ (.A(\cpu.uart_inbound ),
    .B(net944),
    .Y(_01333_));
 sg13g2_or2_1 _07460_ (.X(_01334_),
    .B(\cpu.registers[1][0] ),
    .A(\cpu.uart_inbound ));
 sg13g2_nor3_1 _07461_ (.A(net4051),
    .B(_01257_),
    .C(net4038),
    .Y(_01335_));
 sg13g2_nor2b_1 _07462_ (.A(\cpu.current_instruction[6] ),
    .B_N(net4448),
    .Y(_01336_));
 sg13g2_nand2_2 _07463_ (.Y(_01337_),
    .A(_00024_),
    .B(_01336_));
 sg13g2_nor2_1 _07464_ (.A(net4380),
    .B(_00897_),
    .Y(_01338_));
 sg13g2_and2_2 _07465_ (.A(net4402),
    .B(_01338_),
    .X(_01339_));
 sg13g2_nand2_1 _07466_ (.Y(_01340_),
    .A(net4396),
    .B(_01338_));
 sg13g2_a221oi_1 _07467_ (.B2(_01257_),
    .C1(_01335_),
    .B1(net3853),
    .A1(net4038),
    .Y(_01341_),
    .A2(_01337_));
 sg13g2_a21oi_1 _07468_ (.A1(_01247_),
    .A2(_01341_),
    .Y(_01342_),
    .B1(_01333_));
 sg13g2_nor3_1 _07469_ (.A(\cpu.ALU.mode[1] ),
    .B(_01180_),
    .C(_00148_),
    .Y(_01343_));
 sg13g2_inv_1 _07470_ (.Y(_01344_),
    .A(net4029));
 sg13g2_nor2b_2 _07471_ (.A(\cpu.ALU.mode[1] ),
    .B_N(_00148_),
    .Y(_01345_));
 sg13g2_nand2b_1 _07472_ (.Y(_01346_),
    .B(net4474),
    .A_N(net4465));
 sg13g2_xor2_1 _07473_ (.B(net4474),
    .A(net4465),
    .X(_01347_));
 sg13g2_a22oi_1 _07474_ (.Y(_01348_),
    .B1(_01345_),
    .B2(_01347_),
    .A2(net4030),
    .A1(net4463));
 sg13g2_nand2_2 _07475_ (.Y(_01349_),
    .A(net4465),
    .B(net4474));
 sg13g2_nand2_1 _07476_ (.Y(_01350_),
    .A(\cpu.ALU.mode[1] ),
    .B(_00148_));
 sg13g2_nor2_2 _07477_ (.A(\cpu.ALU.mode[0] ),
    .B(_01350_),
    .Y(_01351_));
 sg13g2_nand2b_1 _07478_ (.Y(_01352_),
    .B(_01351_),
    .A_N(_01349_));
 sg13g2_nor2_1 _07479_ (.A(_01180_),
    .B(_01350_),
    .Y(_01353_));
 sg13g2_nand3_1 _07480_ (.B(\cpu.ALU.mode[0] ),
    .C(_00148_),
    .A(\cpu.ALU.mode[1] ),
    .Y(_01354_));
 sg13g2_nand2_1 _07481_ (.Y(_01355_),
    .A(_01349_),
    .B(_01353_));
 sg13g2_nand3_1 _07482_ (.B(_01352_),
    .C(_01355_),
    .A(_01348_),
    .Y(_01356_));
 sg13g2_inv_1 _07483_ (.Y(_01357_),
    .A(_01356_));
 sg13g2_nor2_1 _07484_ (.A(net4036),
    .B(_01337_),
    .Y(_01358_));
 sg13g2_a21oi_1 _07485_ (.A1(_01257_),
    .A2(net3854),
    .Y(_01359_),
    .B1(_01358_));
 sg13g2_inv_1 _07486_ (.Y(_01360_),
    .A(_01359_));
 sg13g2_a21oi_1 _07487_ (.A1(_01356_),
    .A2(_01360_),
    .Y(_01361_),
    .B1(_01342_));
 sg13g2_nand3b_1 _07488_ (.B(_00026_),
    .C(net4450),
    .Y(_01362_),
    .A_N(net4449));
 sg13g2_inv_4 _07489_ (.A(net4149),
    .Y(_01363_));
 sg13g2_nor2_1 _07490_ (.A(_01235_),
    .B(_01264_),
    .Y(_01364_));
 sg13g2_a21o_1 _07491_ (.A2(net4148),
    .A1(_01264_),
    .B1(_01364_),
    .X(_01365_));
 sg13g2_a21oi_1 _07492_ (.A1(_01235_),
    .A2(net3853),
    .Y(_01366_),
    .B1(_01365_));
 sg13g2_nand3_1 _07493_ (.B(_01235_),
    .C(net3854),
    .A(\cpu.current_address[0] ),
    .Y(_01367_));
 sg13g2_o21ai_1 _07494_ (.B1(_01367_),
    .Y(_01368_),
    .A1(_01333_),
    .A2(_01366_));
 sg13g2_nor2_2 _07495_ (.A(net4320),
    .B(net4299),
    .Y(_01369_));
 sg13g2_or2_1 _07496_ (.X(_01370_),
    .B(net4307),
    .A(net4316));
 sg13g2_nor2_2 _07497_ (.A(net4301),
    .B(_01370_),
    .Y(_01371_));
 sg13g2_or2_1 _07498_ (.X(_01372_),
    .B(_01371_),
    .A(_01290_));
 sg13g2_a21oi_1 _07499_ (.A1(net4326),
    .A2(net3854),
    .Y(_01373_),
    .B1(_01334_));
 sg13g2_nor3_1 _07500_ (.A(net4243),
    .B(_01170_),
    .C(net3852),
    .Y(_01374_));
 sg13g2_a21oi_1 _07501_ (.A1(net4317),
    .A2(_01245_),
    .Y(_01375_),
    .B1(net4301));
 sg13g2_nor4_1 _07502_ (.A(net3865),
    .B(_01373_),
    .C(_01374_),
    .D(_01375_),
    .Y(_01376_));
 sg13g2_a221oi_1 _07503_ (.B2(_01334_),
    .C1(_01376_),
    .B1(_01372_),
    .A1(net4309),
    .Y(_01377_),
    .A2(_01368_));
 sg13g2_o21ai_1 _07504_ (.B1(_01377_),
    .Y(_06992_),
    .A1(net4257),
    .A2(_01361_));
 sg13g2_a22oi_1 _07505_ (.Y(_01378_),
    .B1(net4472),
    .B2(net4465),
    .A2(net4474),
    .A1(net4463));
 sg13g2_nand2_2 _07506_ (.Y(_01379_),
    .A(net4463),
    .B(net4472));
 sg13g2_or2_1 _07507_ (.X(_01380_),
    .B(_01379_),
    .A(_01349_));
 sg13g2_nor3_1 _07508_ (.A(\cpu.ALU.mode[0] ),
    .B(_01350_),
    .C(_01378_),
    .Y(_01381_));
 sg13g2_nor3_1 _07509_ (.A(\cpu.ALU.mode[1] ),
    .B(\cpu.ALU.mode[0] ),
    .C(_00148_),
    .Y(_01382_));
 sg13g2_a22oi_1 _07510_ (.Y(_01383_),
    .B1(net4145),
    .B2(net4465),
    .A2(_01379_),
    .A1(net4028));
 sg13g2_a22oi_1 _07511_ (.Y(_01384_),
    .B1(_01380_),
    .B2(_01381_),
    .A2(net4029),
    .A1(net4461));
 sg13g2_xnor2_1 _07512_ (.Y(_01385_),
    .A(net4463),
    .B(net4472));
 sg13g2_and2_1 _07513_ (.A(_01180_),
    .B(_01345_),
    .X(_01386_));
 sg13g2_nand2_1 _07514_ (.Y(_01387_),
    .A(_01180_),
    .B(_01345_));
 sg13g2_a21oi_1 _07515_ (.A1(_01349_),
    .A2(_01385_),
    .Y(_01388_),
    .B1(_01387_));
 sg13g2_o21ai_1 _07516_ (.B1(_01388_),
    .Y(_01389_),
    .A1(_01349_),
    .A2(_01385_));
 sg13g2_and2_2 _07517_ (.A(\cpu.ALU.mode[0] ),
    .B(_01345_),
    .X(_01390_));
 sg13g2_nand2_1 _07518_ (.Y(_01391_),
    .A(\cpu.ALU.mode[0] ),
    .B(_01345_));
 sg13g2_xor2_1 _07519_ (.B(_01385_),
    .A(_01346_),
    .X(_01392_));
 sg13g2_nand2_1 _07520_ (.Y(_01393_),
    .A(_01390_),
    .B(_01392_));
 sg13g2_and4_2 _07521_ (.A(_01383_),
    .B(_01384_),
    .C(_01389_),
    .D(_01393_),
    .X(_01394_));
 sg13g2_inv_1 _07522_ (.Y(_01395_),
    .A(_01394_));
 sg13g2_nor2_1 _07523_ (.A(net4330),
    .B(\cpu.registers[1][1] ),
    .Y(_01396_));
 sg13g2_nor2_1 _07524_ (.A(_01341_),
    .B(_01396_),
    .Y(_01397_));
 sg13g2_a21oi_1 _07525_ (.A1(net4243),
    .A2(_00152_),
    .Y(_01398_),
    .B1(net3865));
 sg13g2_nand3_1 _07526_ (.B(net4362),
    .C(net3854),
    .A(net4326),
    .Y(_01399_));
 sg13g2_o21ai_1 _07527_ (.B1(_01398_),
    .Y(_01400_),
    .A1(net4240),
    .A2(_01399_));
 sg13g2_o21ai_1 _07528_ (.B1(_01400_),
    .Y(_01401_),
    .A1(_01359_),
    .A2(_01394_));
 sg13g2_o21ai_1 _07529_ (.B1(net4317),
    .Y(_01402_),
    .A1(_01397_),
    .A2(_01401_));
 sg13g2_nand3_1 _07530_ (.B(_01398_),
    .C(_01399_),
    .A(net4301),
    .Y(_01403_));
 sg13g2_o21ai_1 _07531_ (.B1(_01372_),
    .Y(_01404_),
    .A1(net4326),
    .A2(net878));
 sg13g2_nand3_1 _07532_ (.B(_01235_),
    .C(net3854),
    .A(\cpu.current_address[1] ),
    .Y(_01405_));
 sg13g2_o21ai_1 _07533_ (.B1(_01405_),
    .Y(_01406_),
    .A1(_01366_),
    .A2(_01396_));
 sg13g2_nand2_1 _07534_ (.Y(_01407_),
    .A(net4309),
    .B(_01406_));
 sg13g2_nand4_1 _07535_ (.B(_01403_),
    .C(_01404_),
    .A(_01402_),
    .Y(_06993_),
    .D(_01407_));
 sg13g2_nor3_1 _07536_ (.A(net4452),
    .B(net342),
    .C(_01268_),
    .Y(_00008_));
 sg13g2_nor3_1 _07537_ (.A(net4241),
    .B(net342),
    .C(_01268_),
    .Y(_00009_));
 sg13g2_nand2_2 _07538_ (.Y(_01408_),
    .A(net4330),
    .B(net45));
 sg13g2_inv_1 _07539_ (.Y(_00000_),
    .A(net4140));
 sg13g2_o21ai_1 _07540_ (.B1(net4317),
    .Y(_01409_),
    .A1(net4051),
    .A2(_01356_));
 sg13g2_and2_2 _07541_ (.A(net4233),
    .B(_01409_),
    .X(_01410_));
 sg13g2_nor2_1 _07542_ (.A(net4385),
    .B(net4210),
    .Y(_01411_));
 sg13g2_nand2_2 _07543_ (.Y(_01412_),
    .A(net4213),
    .B(net4367));
 sg13g2_nor2_2 _07544_ (.A(net4392),
    .B(net4002),
    .Y(_01413_));
 sg13g2_nor2_1 _07545_ (.A(_00147_),
    .B(net3851),
    .Y(_01414_));
 sg13g2_a21oi_1 _07546_ (.A1(_01170_),
    .A2(net3851),
    .Y(_01415_),
    .B1(_01414_));
 sg13g2_nor3_2 _07547_ (.A(net4380),
    .B(net4396),
    .C(_00897_),
    .Y(_01416_));
 sg13g2_nor3_2 _07548_ (.A(_00016_),
    .B(_01229_),
    .C(_01256_),
    .Y(_01417_));
 sg13g2_and2_1 _07549_ (.A(_00890_),
    .B(_01235_),
    .X(_01418_));
 sg13g2_nor2_1 _07550_ (.A(_01417_),
    .B(_01418_),
    .Y(_01419_));
 sg13g2_nor2_2 _07551_ (.A(_01416_),
    .B(_01419_),
    .Y(_01420_));
 sg13g2_nand2b_1 _07552_ (.Y(_01421_),
    .B(_01420_),
    .A_N(net3849));
 sg13g2_a21o_1 _07553_ (.A2(_01416_),
    .A1(_01235_),
    .B1(_01364_),
    .X(_01422_));
 sg13g2_a22oi_1 _07554_ (.Y(_01423_),
    .B1(_01422_),
    .B2(_00890_),
    .A2(_01270_),
    .A1(_00896_));
 sg13g2_a21oi_1 _07555_ (.A1(net4316),
    .A2(_01335_),
    .Y(_01424_),
    .B1(_01371_));
 sg13g2_nor2_1 _07556_ (.A(net4312),
    .B(net3864),
    .Y(_01425_));
 sg13g2_nand2_1 _07557_ (.Y(_01426_),
    .A(net4326),
    .B(net4451));
 sg13g2_and2_1 _07558_ (.A(_01425_),
    .B(_01426_),
    .X(_01427_));
 sg13g2_nor2_1 _07559_ (.A(net4448),
    .B(\cpu.current_instruction[6] ),
    .Y(_01428_));
 sg13g2_nand2_1 _07560_ (.Y(_01429_),
    .A(_00024_),
    .B(_01428_));
 sg13g2_nor2_1 _07561_ (.A(net4312),
    .B(_01429_),
    .Y(_01430_));
 sg13g2_a221oi_1 _07562_ (.B2(net4038),
    .C1(_01427_),
    .B1(_01430_),
    .A1(_01416_),
    .Y(_01431_),
    .A2(_01417_));
 sg13g2_and2_2 _07563_ (.A(_01424_),
    .B(_01431_),
    .X(_01432_));
 sg13g2_nor2b_1 _07564_ (.A(net4448),
    .B_N(\cpu.current_instruction[6] ),
    .Y(_01433_));
 sg13g2_nor2_1 _07565_ (.A(net4450),
    .B(net4448),
    .Y(_01434_));
 sg13g2_nand2_1 _07566_ (.Y(_01435_),
    .A(net4239),
    .B(_01433_));
 sg13g2_nor2_1 _07567_ (.A(_00018_),
    .B(net4032),
    .Y(_01436_));
 sg13g2_and2_1 _07568_ (.A(net4038),
    .B(_01429_),
    .X(_01437_));
 sg13g2_a21oi_1 _07569_ (.A1(net4445),
    .A2(_01428_),
    .Y(_01438_),
    .B1(net4257));
 sg13g2_a22oi_1 _07570_ (.Y(_01439_),
    .B1(_01437_),
    .B2(_01438_),
    .A2(_01436_),
    .A1(net3999));
 sg13g2_nand4_1 _07571_ (.B(_01423_),
    .C(_01432_),
    .A(_01421_),
    .Y(_01440_),
    .D(_01439_));
 sg13g2_nand3_1 _07572_ (.B(net4033),
    .C(net4147),
    .A(\cpu.current_address[0] ),
    .Y(_01441_));
 sg13g2_o21ai_1 _07573_ (.B1(_01441_),
    .Y(_01442_),
    .A1(net4051),
    .A2(_01409_));
 sg13g2_inv_2 _07574_ (.Y(_01443_),
    .A(_01442_));
 sg13g2_o21ai_1 _07575_ (.B1(_01443_),
    .Y(_01444_),
    .A1(_01410_),
    .A2(_01415_));
 sg13g2_mux2_1 _07576_ (.A0(_01444_),
    .A1(net418),
    .S(net3626),
    .X(_00263_));
 sg13g2_nand3_1 _07577_ (.B(net4033),
    .C(net4147),
    .A(\cpu.current_address[1] ),
    .Y(_01445_));
 sg13g2_a21oi_1 _07578_ (.A1(net3867),
    .A2(_01394_),
    .Y(_01446_),
    .B1(net4261));
 sg13g2_nand2_1 _07579_ (.Y(_01447_),
    .A(net3867),
    .B(_01446_));
 sg13g2_nand2_2 _07580_ (.Y(_01448_),
    .A(_01445_),
    .B(_01447_));
 sg13g2_nor2b_1 _07581_ (.A(net3851),
    .B_N(_00151_),
    .Y(_01449_));
 sg13g2_a21oi_1 _07582_ (.A1(net4362),
    .A2(net3850),
    .Y(_01450_),
    .B1(_01449_));
 sg13g2_nor2_2 _07583_ (.A(\cpu.execution_stage[5] ),
    .B(_01446_),
    .Y(_01451_));
 sg13g2_a21oi_1 _07584_ (.A1(_01445_),
    .A2(_01451_),
    .Y(_01452_),
    .B1(net3625));
 sg13g2_o21ai_1 _07585_ (.B1(_01452_),
    .Y(_01453_),
    .A1(_01448_),
    .A2(_01450_));
 sg13g2_nand2_1 _07586_ (.Y(_01454_),
    .A(net224),
    .B(net3625));
 sg13g2_nand2_1 _07587_ (.Y(_00264_),
    .A(_01453_),
    .B(_01454_));
 sg13g2_nand2_1 _07588_ (.Y(_01455_),
    .A(net4465),
    .B(net4470));
 sg13g2_nand2_1 _07589_ (.Y(_01456_),
    .A(net4473),
    .B(net4461));
 sg13g2_xor2_1 _07590_ (.B(_01456_),
    .A(_01379_),
    .X(_01457_));
 sg13g2_nand2b_1 _07591_ (.Y(_01458_),
    .B(_01457_),
    .A_N(_01455_));
 sg13g2_xor2_1 _07592_ (.B(_01457_),
    .A(_01455_),
    .X(_01459_));
 sg13g2_nand2_1 _07593_ (.Y(_01460_),
    .A(_01380_),
    .B(_01459_));
 sg13g2_or2_1 _07594_ (.X(_01461_),
    .B(_01459_),
    .A(_01380_));
 sg13g2_nand3_1 _07595_ (.B(_01460_),
    .C(_01461_),
    .A(_01351_),
    .Y(_01462_));
 sg13g2_nand2_1 _07596_ (.Y(_01463_),
    .A(net4461),
    .B(\cpu.ALU.b[2] ));
 sg13g2_inv_1 _07597_ (.Y(_01464_),
    .A(_01463_));
 sg13g2_xor2_1 _07598_ (.B(net4470),
    .A(net4461),
    .X(_01465_));
 sg13g2_o21ai_1 _07599_ (.B1(_01379_),
    .Y(_01466_),
    .A1(_01349_),
    .A2(_01385_));
 sg13g2_o21ai_1 _07600_ (.B1(net4027),
    .Y(_01467_),
    .A1(_01465_),
    .A2(_01466_));
 sg13g2_a21o_1 _07601_ (.A2(_01466_),
    .A1(_01465_),
    .B1(_01467_),
    .X(_01468_));
 sg13g2_nor2b_1 _07602_ (.A(net4472),
    .B_N(net4463),
    .Y(_01469_));
 sg13g2_a21oi_1 _07603_ (.A1(_01346_),
    .A2(_01385_),
    .Y(_01470_),
    .B1(_01469_));
 sg13g2_a21oi_1 _07604_ (.A1(_01465_),
    .A2(_01470_),
    .Y(_01471_),
    .B1(_01391_));
 sg13g2_o21ai_1 _07605_ (.B1(_01471_),
    .Y(_01472_),
    .A1(_01465_),
    .A2(_01470_));
 sg13g2_nor2_1 _07606_ (.A(_01354_),
    .B(_01464_),
    .Y(_01473_));
 sg13g2_a221oi_1 _07607_ (.B2(net4463),
    .C1(_01473_),
    .B1(net4145),
    .A1(net4459),
    .Y(_01474_),
    .A2(net4030));
 sg13g2_nand4_1 _07608_ (.B(_01468_),
    .C(_01472_),
    .A(_01462_),
    .Y(_01475_),
    .D(_01474_));
 sg13g2_o21ai_1 _07609_ (.B1(net4319),
    .Y(_01476_),
    .A1(net4052),
    .A2(_01475_));
 sg13g2_and2_1 _07610_ (.A(net4231),
    .B(_01476_),
    .X(_01477_));
 sg13g2_nor2b_1 _07611_ (.A(net3851),
    .B_N(_00155_),
    .Y(_01478_));
 sg13g2_a221oi_1 _07612_ (.B2(net4231),
    .C1(_01478_),
    .B1(_01476_),
    .A1(net4353),
    .Y(_01479_),
    .A2(net3851));
 sg13g2_nand3_1 _07613_ (.B(net4033),
    .C(net4147),
    .A(net466),
    .Y(_01480_));
 sg13g2_o21ai_1 _07614_ (.B1(_01480_),
    .Y(_01481_),
    .A1(net4052),
    .A2(_01476_));
 sg13g2_nor3_1 _07615_ (.A(net3626),
    .B(_01479_),
    .C(_01481_),
    .Y(_01482_));
 sg13g2_a21oi_1 _07616_ (.A1(_00916_),
    .A2(net3626),
    .Y(_00265_),
    .B1(_01482_));
 sg13g2_nand2_2 _07617_ (.Y(_01483_),
    .A(net4466),
    .B(net4469));
 sg13g2_o21ai_1 _07618_ (.B1(_01458_),
    .Y(_01484_),
    .A1(_01379_),
    .A2(_01456_));
 sg13g2_nand2_1 _07619_ (.Y(_01485_),
    .A(net4464),
    .B(net4470));
 sg13g2_and4_1 _07620_ (.A(net4473),
    .B(net4461),
    .C(net4471),
    .D(net4459),
    .X(_01486_));
 sg13g2_a22oi_1 _07621_ (.Y(_01487_),
    .B1(net4459),
    .B2(net4473),
    .A2(net4471),
    .A1(net4461));
 sg13g2_nor3_1 _07622_ (.A(_01485_),
    .B(_01486_),
    .C(_01487_),
    .Y(_01488_));
 sg13g2_o21ai_1 _07623_ (.B1(_01485_),
    .Y(_01489_),
    .A1(_01486_),
    .A2(_01487_));
 sg13g2_nor2b_1 _07624_ (.A(_01488_),
    .B_N(_01489_),
    .Y(_01490_));
 sg13g2_nand2_1 _07625_ (.Y(_01491_),
    .A(_01484_),
    .B(_01490_));
 sg13g2_xnor2_1 _07626_ (.Y(_01492_),
    .A(_01484_),
    .B(_01490_));
 sg13g2_xnor2_1 _07627_ (.Y(_01493_),
    .A(_01483_),
    .B(_01492_));
 sg13g2_or2_1 _07628_ (.X(_01494_),
    .B(_01493_),
    .A(_01461_));
 sg13g2_nand2_1 _07629_ (.Y(_01495_),
    .A(_01461_),
    .B(_01493_));
 sg13g2_nand3_1 _07630_ (.B(_01494_),
    .C(_01495_),
    .A(_01351_),
    .Y(_01496_));
 sg13g2_and2_1 _07631_ (.A(net4459),
    .B(\cpu.ALU.b[3] ),
    .X(_01497_));
 sg13g2_nand2_2 _07632_ (.Y(_01498_),
    .A(net4460),
    .B(\cpu.ALU.b[3] ));
 sg13g2_xnor2_1 _07633_ (.Y(_01499_),
    .A(net4459),
    .B(net4469));
 sg13g2_nand2b_1 _07634_ (.Y(_01500_),
    .B(net4461),
    .A_N(net4470));
 sg13g2_o21ai_1 _07635_ (.B1(_01500_),
    .Y(_01501_),
    .A1(_01465_),
    .A2(_01470_));
 sg13g2_a21oi_1 _07636_ (.A1(_01499_),
    .A2(_01501_),
    .Y(_01502_),
    .B1(net4025));
 sg13g2_o21ai_1 _07637_ (.B1(_01502_),
    .Y(_01503_),
    .A1(_01499_),
    .A2(_01501_));
 sg13g2_nor2_1 _07638_ (.A(_01354_),
    .B(_01497_),
    .Y(_01504_));
 sg13g2_a221oi_1 _07639_ (.B2(net4462),
    .C1(_01504_),
    .B1(net4145),
    .A1(net4457),
    .Y(_01505_),
    .A2(net4030));
 sg13g2_a21oi_1 _07640_ (.A1(_01465_),
    .A2(_01466_),
    .Y(_01506_),
    .B1(_01464_));
 sg13g2_a21oi_1 _07641_ (.A1(_01499_),
    .A2(_01506_),
    .Y(_01507_),
    .B1(_01387_));
 sg13g2_o21ai_1 _07642_ (.B1(_01507_),
    .Y(_01508_),
    .A1(_01499_),
    .A2(_01506_));
 sg13g2_nand4_1 _07643_ (.B(_01503_),
    .C(_01505_),
    .A(_01496_),
    .Y(_01509_),
    .D(_01508_));
 sg13g2_nor2_1 _07644_ (.A(net4057),
    .B(_01509_),
    .Y(_01510_));
 sg13g2_nor2_2 _07645_ (.A(net4262),
    .B(_01510_),
    .Y(_01511_));
 sg13g2_o21ai_1 _07646_ (.B1(net4319),
    .Y(_01512_),
    .A1(net4057),
    .A2(_01509_));
 sg13g2_nand2_1 _07647_ (.Y(_01513_),
    .A(_01171_),
    .B(net3850));
 sg13g2_o21ai_1 _07648_ (.B1(_01513_),
    .Y(_01514_),
    .A1(_00159_),
    .A2(net3850));
 sg13g2_o21ai_1 _07649_ (.B1(_01511_),
    .Y(_01515_),
    .A1(net3868),
    .A2(_01514_));
 sg13g2_and3_2 _07650_ (.X(_01516_),
    .A(\cpu.current_address[3] ),
    .B(net4033),
    .C(net4147));
 sg13g2_a21oi_1 _07651_ (.A1(net4300),
    .A2(_01514_),
    .Y(_01517_),
    .B1(_01516_));
 sg13g2_nor2b_1 _07652_ (.A(net3626),
    .B_N(_01517_),
    .Y(_01518_));
 sg13g2_a22oi_1 _07653_ (.Y(_00266_),
    .B1(_01515_),
    .B2(_01518_),
    .A2(net3625),
    .A1(_00924_));
 sg13g2_a22oi_1 _07654_ (.Y(_01519_),
    .B1(\cpu.ALU.b[4] ),
    .B2(net4466),
    .A2(net4469),
    .A1(net4464));
 sg13g2_nand2_1 _07655_ (.Y(_01520_),
    .A(net4464),
    .B(net4468));
 sg13g2_or2_1 _07656_ (.X(_01521_),
    .B(_01520_),
    .A(_01483_));
 sg13g2_nand2b_1 _07657_ (.Y(_01522_),
    .B(_01521_),
    .A_N(_01519_));
 sg13g2_or2_1 _07658_ (.X(_01523_),
    .B(_01488_),
    .A(_01486_));
 sg13g2_and4_1 _07659_ (.A(net4474),
    .B(net4471),
    .C(net4460),
    .D(net4458),
    .X(_01524_));
 sg13g2_a22oi_1 _07660_ (.Y(_01525_),
    .B1(net4458),
    .B2(net4473),
    .A2(net4460),
    .A1(net4472));
 sg13g2_nor2_1 _07661_ (.A(_01524_),
    .B(_01525_),
    .Y(_01526_));
 sg13g2_xnor2_1 _07662_ (.Y(_01527_),
    .A(_01463_),
    .B(_01526_));
 sg13g2_nand2_1 _07663_ (.Y(_01528_),
    .A(_01523_),
    .B(_01527_));
 sg13g2_nor2_1 _07664_ (.A(_01523_),
    .B(_01527_),
    .Y(_01529_));
 sg13g2_xor2_1 _07665_ (.B(_01527_),
    .A(_01523_),
    .X(_01530_));
 sg13g2_xnor2_1 _07666_ (.Y(_01531_),
    .A(_01522_),
    .B(_01530_));
 sg13g2_o21ai_1 _07667_ (.B1(_01491_),
    .Y(_01532_),
    .A1(_01483_),
    .A2(_01492_));
 sg13g2_nand2_1 _07668_ (.Y(_01533_),
    .A(_01531_),
    .B(_01532_));
 sg13g2_xnor2_1 _07669_ (.Y(_01534_),
    .A(_01531_),
    .B(_01532_));
 sg13g2_nor2_1 _07670_ (.A(_01494_),
    .B(_01534_),
    .Y(_01535_));
 sg13g2_xor2_1 _07671_ (.B(_01534_),
    .A(_01494_),
    .X(_01536_));
 sg13g2_nand2_2 _07672_ (.Y(_01537_),
    .A(net4457),
    .B(net4468));
 sg13g2_inv_1 _07673_ (.Y(_01538_),
    .A(_01537_));
 sg13g2_xor2_1 _07674_ (.B(net4468),
    .A(net4457),
    .X(_01539_));
 sg13g2_xnor2_1 _07675_ (.Y(_01540_),
    .A(net4457),
    .B(net4468));
 sg13g2_nor2b_1 _07676_ (.A(net4469),
    .B_N(net4459),
    .Y(_01541_));
 sg13g2_a21oi_1 _07677_ (.A1(_01499_),
    .A2(_01501_),
    .Y(_01542_),
    .B1(_01541_));
 sg13g2_a21oi_1 _07678_ (.A1(_01539_),
    .A2(_01542_),
    .Y(_01543_),
    .B1(net4025));
 sg13g2_o21ai_1 _07679_ (.B1(_01543_),
    .Y(_01544_),
    .A1(_01539_),
    .A2(_01542_));
 sg13g2_o21ai_1 _07680_ (.B1(_01498_),
    .Y(_01545_),
    .A1(_01499_),
    .A2(_01506_));
 sg13g2_o21ai_1 _07681_ (.B1(net4027),
    .Y(_01546_),
    .A1(_01539_),
    .A2(_01545_));
 sg13g2_a21o_1 _07682_ (.A2(_01545_),
    .A1(_01539_),
    .B1(_01546_),
    .X(_01547_));
 sg13g2_nand2_1 _07683_ (.Y(_01548_),
    .A(net4459),
    .B(net4145));
 sg13g2_a22oi_1 _07684_ (.Y(_01549_),
    .B1(net4028),
    .B2(_01537_),
    .A2(net4030),
    .A1(net4455));
 sg13g2_nand4_1 _07685_ (.B(_01547_),
    .C(_01548_),
    .A(_01544_),
    .Y(_01550_),
    .D(_01549_));
 sg13g2_a21oi_2 _07686_ (.B1(_01550_),
    .Y(_01551_),
    .A2(_01536_),
    .A1(_01351_));
 sg13g2_a21o_2 _07687_ (.A2(_01551_),
    .A1(net3869),
    .B1(net4266),
    .X(_01552_));
 sg13g2_nand2_1 _07688_ (.Y(_01553_),
    .A(_01172_),
    .B(_01413_));
 sg13g2_o21ai_1 _07689_ (.B1(_01553_),
    .Y(_01554_),
    .A1(_00163_),
    .A2(net3850));
 sg13g2_nor2_1 _07690_ (.A(net3869),
    .B(_01554_),
    .Y(_01555_));
 sg13g2_and3_2 _07691_ (.X(_01556_),
    .A(\cpu.current_address[4] ),
    .B(net4033),
    .C(net4147));
 sg13g2_a21oi_1 _07692_ (.A1(net4300),
    .A2(_01554_),
    .Y(_01557_),
    .B1(_01556_));
 sg13g2_o21ai_1 _07693_ (.B1(_01557_),
    .Y(_01558_),
    .A1(_01552_),
    .A2(_01555_));
 sg13g2_mux2_1 _07694_ (.A0(_01558_),
    .A1(net410),
    .S(net3625),
    .X(_00267_));
 sg13g2_o21ai_1 _07695_ (.B1(_01528_),
    .Y(_01559_),
    .A1(_01522_),
    .A2(_01529_));
 sg13g2_nand2_1 _07696_ (.Y(_01560_),
    .A(net4466),
    .B(\cpu.ALU.b[5] ));
 sg13g2_nand2_1 _07697_ (.Y(_01561_),
    .A(net4462),
    .B(net4468));
 sg13g2_nand2_1 _07698_ (.Y(_01562_),
    .A(net4462),
    .B(net4469));
 sg13g2_xor2_1 _07699_ (.B(_01562_),
    .A(_01520_),
    .X(_01563_));
 sg13g2_nand2b_1 _07700_ (.Y(_01564_),
    .B(_01563_),
    .A_N(_01560_));
 sg13g2_xor2_1 _07701_ (.B(_01563_),
    .A(_01560_),
    .X(_01565_));
 sg13g2_a21o_1 _07702_ (.A2(_01526_),
    .A1(_01464_),
    .B1(_01524_),
    .X(_01566_));
 sg13g2_nand2_1 _07703_ (.Y(_01567_),
    .A(net4460),
    .B(net4470));
 sg13g2_nand2_1 _07704_ (.Y(_01568_),
    .A(net4471),
    .B(net4456));
 sg13g2_and4_1 _07705_ (.A(net4473),
    .B(net4471),
    .C(net4458),
    .D(net4456),
    .X(_01569_));
 sg13g2_a22oi_1 _07706_ (.Y(_01570_),
    .B1(net4456),
    .B2(net4473),
    .A2(net4458),
    .A1(net4471));
 sg13g2_nor3_1 _07707_ (.A(_01567_),
    .B(_01569_),
    .C(_01570_),
    .Y(_01571_));
 sg13g2_o21ai_1 _07708_ (.B1(_01567_),
    .Y(_01572_),
    .A1(_01569_),
    .A2(_01570_));
 sg13g2_nor2b_1 _07709_ (.A(_01571_),
    .B_N(_01572_),
    .Y(_01573_));
 sg13g2_nand2_1 _07710_ (.Y(_01574_),
    .A(_01566_),
    .B(_01573_));
 sg13g2_xnor2_1 _07711_ (.Y(_01575_),
    .A(_01566_),
    .B(_01573_));
 sg13g2_xnor2_1 _07712_ (.Y(_01576_),
    .A(_01565_),
    .B(_01575_));
 sg13g2_nand2b_1 _07713_ (.Y(_01577_),
    .B(_01559_),
    .A_N(_01576_));
 sg13g2_xor2_1 _07714_ (.B(_01576_),
    .A(_01559_),
    .X(_01578_));
 sg13g2_xor2_1 _07715_ (.B(_01578_),
    .A(_01521_),
    .X(_01579_));
 sg13g2_nand2b_1 _07716_ (.Y(_01580_),
    .B(_01579_),
    .A_N(_01533_));
 sg13g2_xnor2_1 _07717_ (.Y(_01581_),
    .A(_01533_),
    .B(_01579_));
 sg13g2_and2_1 _07718_ (.A(_01535_),
    .B(_01581_),
    .X(_01582_));
 sg13g2_xor2_1 _07719_ (.B(_01581_),
    .A(_01535_),
    .X(_01583_));
 sg13g2_nor2_1 _07720_ (.A(net4455),
    .B(net4467),
    .Y(_01584_));
 sg13g2_xnor2_1 _07721_ (.Y(_01585_),
    .A(net4455),
    .B(net4467));
 sg13g2_nand2b_1 _07722_ (.Y(_01586_),
    .B(net4457),
    .A_N(net4468));
 sg13g2_o21ai_1 _07723_ (.B1(_01586_),
    .Y(_01587_),
    .A1(_01539_),
    .A2(_01542_));
 sg13g2_and2_1 _07724_ (.A(_01585_),
    .B(_01587_),
    .X(_01588_));
 sg13g2_o21ai_1 _07725_ (.B1(_01390_),
    .Y(_01589_),
    .A1(_01585_),
    .A2(_01587_));
 sg13g2_a21oi_1 _07726_ (.A1(_01539_),
    .A2(_01545_),
    .Y(_01590_),
    .B1(_01538_));
 sg13g2_xor2_1 _07727_ (.B(_01590_),
    .A(_01585_),
    .X(_01591_));
 sg13g2_a21oi_1 _07728_ (.A1(net4455),
    .A2(net4467),
    .Y(_01592_),
    .B1(_01354_));
 sg13g2_a221oi_1 _07729_ (.B2(net4457),
    .C1(_01592_),
    .B1(net4145),
    .A1(net4454),
    .Y(_01593_),
    .A2(net4030));
 sg13g2_o21ai_1 _07730_ (.B1(_01593_),
    .Y(_01594_),
    .A1(_01588_),
    .A2(_01589_));
 sg13g2_a221oi_1 _07731_ (.B2(net4027),
    .C1(_01594_),
    .B1(_01591_),
    .A1(_01351_),
    .Y(_01595_),
    .A2(_01583_));
 sg13g2_nand2_2 _07732_ (.Y(_01596_),
    .A(net3867),
    .B(_01595_));
 sg13g2_nor2_1 _07733_ (.A(_00167_),
    .B(net3850),
    .Y(_01597_));
 sg13g2_a21oi_1 _07734_ (.A1(_01173_),
    .A2(net3850),
    .Y(_01598_),
    .B1(_01597_));
 sg13g2_a21oi_1 _07735_ (.A1(net4054),
    .A2(_01598_),
    .Y(_01599_),
    .B1(net4260));
 sg13g2_nand2_1 _07736_ (.Y(_01600_),
    .A(_01596_),
    .B(_01599_));
 sg13g2_and3_2 _07737_ (.X(_01601_),
    .A(\cpu.current_address[5] ),
    .B(net4034),
    .C(net4147));
 sg13g2_nor2_1 _07738_ (.A(net4234),
    .B(_01598_),
    .Y(_01602_));
 sg13g2_nor3_1 _07739_ (.A(net3625),
    .B(_01601_),
    .C(_01602_),
    .Y(_01603_));
 sg13g2_a22oi_1 _07740_ (.Y(_00268_),
    .B1(_01600_),
    .B2(_01603_),
    .A2(net3625),
    .A1(_00938_));
 sg13g2_o21ai_1 _07741_ (.B1(_01577_),
    .Y(_01604_),
    .A1(_01521_),
    .A2(_01578_));
 sg13g2_o21ai_1 _07742_ (.B1(_01564_),
    .Y(_01605_),
    .A1(_01520_),
    .A2(_01562_));
 sg13g2_nand2_2 _07743_ (.Y(_01606_),
    .A(net4465),
    .B(\cpu.ALU.b[6] ));
 sg13g2_nand2b_1 _07744_ (.Y(_01607_),
    .B(_01605_),
    .A_N(_01606_));
 sg13g2_xnor2_1 _07745_ (.Y(_01608_),
    .A(_01605_),
    .B(_01606_));
 sg13g2_inv_1 _07746_ (.Y(_01609_),
    .A(_01608_));
 sg13g2_o21ai_1 _07747_ (.B1(_01574_),
    .Y(_01610_),
    .A1(_01565_),
    .A2(_01575_));
 sg13g2_nand2_1 _07748_ (.Y(_01611_),
    .A(net4463),
    .B(net4467));
 sg13g2_xnor2_1 _07749_ (.Y(_01612_),
    .A(_01497_),
    .B(_01561_));
 sg13g2_nand2b_1 _07750_ (.Y(_01613_),
    .B(_01612_),
    .A_N(_01611_));
 sg13g2_xor2_1 _07751_ (.B(_01612_),
    .A(_01611_),
    .X(_01614_));
 sg13g2_or2_1 _07752_ (.X(_01615_),
    .B(_01571_),
    .A(_01569_));
 sg13g2_nand2_1 _07753_ (.Y(_01616_),
    .A(net4470),
    .B(net4457));
 sg13g2_nand2_1 _07754_ (.Y(_01617_),
    .A(net4473),
    .B(\cpu.ALU.a[6] ));
 sg13g2_or2_1 _07755_ (.X(_01618_),
    .B(_01617_),
    .A(_01568_));
 sg13g2_and2_1 _07756_ (.A(_01568_),
    .B(_01617_),
    .X(_01619_));
 sg13g2_xor2_1 _07757_ (.B(_01617_),
    .A(_01568_),
    .X(_01620_));
 sg13g2_xnor2_1 _07758_ (.Y(_01621_),
    .A(_01616_),
    .B(_01620_));
 sg13g2_nand2_1 _07759_ (.Y(_01622_),
    .A(_01615_),
    .B(_01621_));
 sg13g2_xnor2_1 _07760_ (.Y(_01623_),
    .A(_01615_),
    .B(_01621_));
 sg13g2_xor2_1 _07761_ (.B(_01623_),
    .A(_01614_),
    .X(_01624_));
 sg13g2_nand2_1 _07762_ (.Y(_01625_),
    .A(_01610_),
    .B(_01624_));
 sg13g2_xnor2_1 _07763_ (.Y(_01626_),
    .A(_01610_),
    .B(_01624_));
 sg13g2_xnor2_1 _07764_ (.Y(_01627_),
    .A(_01609_),
    .B(_01626_));
 sg13g2_nand2b_1 _07765_ (.Y(_01628_),
    .B(_01604_),
    .A_N(_01627_));
 sg13g2_xnor2_1 _07766_ (.Y(_01629_),
    .A(_01604_),
    .B(_01627_));
 sg13g2_nor2b_1 _07767_ (.A(_01580_),
    .B_N(_01629_),
    .Y(_01630_));
 sg13g2_xnor2_1 _07768_ (.Y(_01631_),
    .A(_01580_),
    .B(_01629_));
 sg13g2_o21ai_1 _07769_ (.B1(_01351_),
    .Y(_01632_),
    .A1(_01582_),
    .A2(_01631_));
 sg13g2_a21oi_1 _07770_ (.A1(_01582_),
    .A2(_01631_),
    .Y(_01633_),
    .B1(_01632_));
 sg13g2_and2_1 _07771_ (.A(net4454),
    .B(\cpu.ALU.b[6] ),
    .X(_01634_));
 sg13g2_xor2_1 _07772_ (.B(\cpu.ALU.b[6] ),
    .A(net4454),
    .X(_01635_));
 sg13g2_xnor2_1 _07773_ (.Y(_01636_),
    .A(net4454),
    .B(\cpu.ALU.b[6] ));
 sg13g2_a221oi_1 _07774_ (.B2(_01545_),
    .C1(_01538_),
    .B1(_01539_),
    .A1(net4455),
    .Y(_01637_),
    .A2(net4467));
 sg13g2_nor3_2 _07775_ (.A(_01584_),
    .B(_01636_),
    .C(_01637_),
    .Y(_01638_));
 sg13g2_o21ai_1 _07776_ (.B1(_01636_),
    .Y(_01639_),
    .A1(_01584_),
    .A2(_01637_));
 sg13g2_nand2_1 _07777_ (.Y(_01640_),
    .A(net4027),
    .B(_01639_));
 sg13g2_nor2_1 _07778_ (.A(_01638_),
    .B(_01640_),
    .Y(_01641_));
 sg13g2_a22oi_1 _07779_ (.Y(_01642_),
    .B1(net4145),
    .B2(net4455),
    .A2(net4030),
    .A1(net4453));
 sg13g2_o21ai_1 _07780_ (.B1(_01642_),
    .Y(_01643_),
    .A1(_01354_),
    .A2(_01634_));
 sg13g2_nor2b_1 _07781_ (.A(net4467),
    .B_N(net4455),
    .Y(_01644_));
 sg13g2_a21oi_1 _07782_ (.A1(_01585_),
    .A2(_01587_),
    .Y(_01645_),
    .B1(_01644_));
 sg13g2_o21ai_1 _07783_ (.B1(_01390_),
    .Y(_01646_),
    .A1(_01635_),
    .A2(_01645_));
 sg13g2_a21oi_1 _07784_ (.A1(_01635_),
    .A2(_01645_),
    .Y(_01647_),
    .B1(_01646_));
 sg13g2_nor4_2 _07785_ (.A(_01633_),
    .B(_01641_),
    .C(_01643_),
    .Y(_01648_),
    .D(_01647_));
 sg13g2_nand2_2 _07786_ (.Y(_01649_),
    .A(net3867),
    .B(_01648_));
 sg13g2_nor2b_1 _07787_ (.A(net3850),
    .B_N(_00171_),
    .Y(_01650_));
 sg13g2_a21oi_1 _07788_ (.A1(net4341),
    .A2(net3850),
    .Y(_01651_),
    .B1(_01650_));
 sg13g2_o21ai_1 _07789_ (.B1(net4319),
    .Y(_01652_),
    .A1(net3868),
    .A2(_01651_));
 sg13g2_inv_1 _07790_ (.Y(_01653_),
    .A(_01652_));
 sg13g2_nand3_1 _07791_ (.B(net4033),
    .C(net4147),
    .A(net142),
    .Y(_01654_));
 sg13g2_a221oi_1 _07792_ (.B2(_01649_),
    .C1(net3625),
    .B1(_01653_),
    .A1(net4299),
    .Y(_01655_),
    .A2(_01651_));
 sg13g2_a22oi_1 _07793_ (.Y(_00269_),
    .B1(_01654_),
    .B2(_01655_),
    .A2(net3625),
    .A1(_00945_));
 sg13g2_a21oi_2 _07794_ (.B1(_01630_),
    .Y(_01656_),
    .A2(_01631_),
    .A1(_01582_));
 sg13g2_o21ai_1 _07795_ (.B1(_01625_),
    .Y(_01657_),
    .A1(_01609_),
    .A2(_01626_));
 sg13g2_nand2_1 _07796_ (.Y(_01658_),
    .A(net4466),
    .B(\cpu.ALU.b[7] ));
 sg13g2_o21ai_1 _07797_ (.B1(_01613_),
    .Y(_01659_),
    .A1(_01498_),
    .A2(_01561_));
 sg13g2_nand2_1 _07798_ (.Y(_01660_),
    .A(net4464),
    .B(\cpu.ALU.b[6] ));
 sg13g2_nand2b_1 _07799_ (.Y(_01661_),
    .B(_01659_),
    .A_N(_01660_));
 sg13g2_xnor2_1 _07800_ (.Y(_01662_),
    .A(_01659_),
    .B(_01660_));
 sg13g2_nand2b_1 _07801_ (.Y(_01663_),
    .B(_01662_),
    .A_N(_01658_));
 sg13g2_xnor2_1 _07802_ (.Y(_01664_),
    .A(_01658_),
    .B(_01662_));
 sg13g2_o21ai_1 _07803_ (.B1(_01622_),
    .Y(_01665_),
    .A1(_01614_),
    .A2(_01623_));
 sg13g2_nand2_1 _07804_ (.Y(_01666_),
    .A(net4462),
    .B(\cpu.ALU.b[5] ));
 sg13g2_a22oi_1 _07805_ (.Y(_01667_),
    .B1(net4468),
    .B2(net4459),
    .A2(net4469),
    .A1(net4457));
 sg13g2_a21oi_1 _07806_ (.A1(_01497_),
    .A2(_01538_),
    .Y(_01668_),
    .B1(_01667_));
 sg13g2_nand2b_1 _07807_ (.Y(_01669_),
    .B(_01668_),
    .A_N(_01666_));
 sg13g2_xor2_1 _07808_ (.B(_01668_),
    .A(_01666_),
    .X(_01670_));
 sg13g2_o21ai_1 _07809_ (.B1(_01618_),
    .Y(_01671_),
    .A1(_01616_),
    .A2(_01619_));
 sg13g2_nand2_1 _07810_ (.Y(_01672_),
    .A(net4470),
    .B(net4456));
 sg13g2_nand2_1 _07811_ (.Y(_01673_),
    .A(net4471),
    .B(\cpu.ALU.a[7] ));
 sg13g2_and4_1 _07812_ (.A(net4473),
    .B(net4472),
    .C(\cpu.ALU.a[6] ),
    .D(net4453),
    .X(_01674_));
 sg13g2_a22oi_1 _07813_ (.Y(_01675_),
    .B1(net4453),
    .B2(net4474),
    .A2(net4454),
    .A1(net4471));
 sg13g2_nor3_1 _07814_ (.A(_01672_),
    .B(_01674_),
    .C(_01675_),
    .Y(_01676_));
 sg13g2_o21ai_1 _07815_ (.B1(_01672_),
    .Y(_01677_),
    .A1(_01674_),
    .A2(_01675_));
 sg13g2_nor2b_1 _07816_ (.A(_01676_),
    .B_N(_01677_),
    .Y(_01678_));
 sg13g2_nand2_1 _07817_ (.Y(_01679_),
    .A(_01671_),
    .B(_01678_));
 sg13g2_xnor2_1 _07818_ (.Y(_01680_),
    .A(_01671_),
    .B(_01678_));
 sg13g2_xor2_1 _07819_ (.B(_01680_),
    .A(_01670_),
    .X(_01681_));
 sg13g2_and2_1 _07820_ (.A(_01665_),
    .B(_01681_),
    .X(_01682_));
 sg13g2_or2_1 _07821_ (.X(_01683_),
    .B(_01681_),
    .A(_01665_));
 sg13g2_xnor2_1 _07822_ (.Y(_01684_),
    .A(_01665_),
    .B(_01681_));
 sg13g2_xnor2_1 _07823_ (.Y(_01685_),
    .A(_01664_),
    .B(_01684_));
 sg13g2_nand2_1 _07824_ (.Y(_01686_),
    .A(_01657_),
    .B(_01685_));
 sg13g2_xnor2_1 _07825_ (.Y(_01687_),
    .A(_01657_),
    .B(_01685_));
 sg13g2_xor2_1 _07826_ (.B(_01687_),
    .A(_01607_),
    .X(_01688_));
 sg13g2_nor2b_1 _07827_ (.A(_01628_),
    .B_N(_01688_),
    .Y(_01689_));
 sg13g2_xnor2_1 _07828_ (.Y(_01690_),
    .A(_01628_),
    .B(_01688_));
 sg13g2_nor2b_1 _07829_ (.A(_01656_),
    .B_N(_01690_),
    .Y(_01691_));
 sg13g2_xnor2_1 _07830_ (.Y(_01692_),
    .A(_01656_),
    .B(_01690_));
 sg13g2_nand2_1 _07831_ (.Y(_01693_),
    .A(net4453),
    .B(\cpu.ALU.b[7] ));
 sg13g2_xnor2_1 _07832_ (.Y(_01694_),
    .A(net4453),
    .B(\cpu.ALU.b[7] ));
 sg13g2_inv_1 _07833_ (.Y(_01695_),
    .A(_01694_));
 sg13g2_nand2b_1 _07834_ (.Y(_01696_),
    .B(net4454),
    .A_N(\cpu.ALU.b[6] ));
 sg13g2_o21ai_1 _07835_ (.B1(_01696_),
    .Y(_01697_),
    .A1(_01635_),
    .A2(_01645_));
 sg13g2_a21oi_1 _07836_ (.A1(_01694_),
    .A2(_01697_),
    .Y(_01698_),
    .B1(net4025));
 sg13g2_o21ai_1 _07837_ (.B1(_01698_),
    .Y(_01699_),
    .A1(_01694_),
    .A2(_01697_));
 sg13g2_o21ai_1 _07838_ (.B1(_01695_),
    .Y(_01700_),
    .A1(_01634_),
    .A2(_01638_));
 sg13g2_nor3_1 _07839_ (.A(_01634_),
    .B(_01638_),
    .C(_01695_),
    .Y(_01701_));
 sg13g2_nand3b_1 _07840_ (.B(net4026),
    .C(_01700_),
    .Y(_01702_),
    .A_N(_01701_));
 sg13g2_nand2_1 _07841_ (.Y(_01703_),
    .A(\cpu.ALU.a[8] ),
    .B(net4029));
 sg13g2_a22oi_1 _07842_ (.Y(_01704_),
    .B1(_01693_),
    .B2(net4028),
    .A2(net4145),
    .A1(net4454));
 sg13g2_nand4_1 _07843_ (.B(_01702_),
    .C(_01703_),
    .A(_01699_),
    .Y(_01705_),
    .D(_01704_));
 sg13g2_a21oi_2 _07844_ (.B1(_01705_),
    .Y(_01706_),
    .A2(_01692_),
    .A1(_01351_));
 sg13g2_nand2_2 _07845_ (.Y(_01707_),
    .A(net3866),
    .B(_01706_));
 sg13g2_nor2_1 _07846_ (.A(_00175_),
    .B(net3851),
    .Y(_01708_));
 sg13g2_a21oi_1 _07847_ (.A1(_01175_),
    .A2(net3851),
    .Y(_01709_),
    .B1(_01708_));
 sg13g2_a21oi_1 _07848_ (.A1(net4052),
    .A2(_01709_),
    .Y(_01710_),
    .B1(net4259));
 sg13g2_nand2_1 _07849_ (.Y(_01711_),
    .A(_01707_),
    .B(_01710_));
 sg13g2_o21ai_1 _07850_ (.B1(net4147),
    .Y(_01712_),
    .A1(net4446),
    .A2(net4034));
 sg13g2_a21oi_2 _07851_ (.B1(_01712_),
    .Y(_01713_),
    .A2(net4033),
    .A1(_01151_));
 sg13g2_nor2_1 _07852_ (.A(net4231),
    .B(_01709_),
    .Y(_01714_));
 sg13g2_nor3_1 _07853_ (.A(net3626),
    .B(_01713_),
    .C(_01714_),
    .Y(_01715_));
 sg13g2_a22oi_1 _07854_ (.Y(_00270_),
    .B1(_01711_),
    .B2(_01715_),
    .A2(net3626),
    .A1(_00953_));
 sg13g2_nor2_1 _07855_ (.A(_01689_),
    .B(_01691_),
    .Y(_01716_));
 sg13g2_o21ai_1 _07856_ (.B1(_01686_),
    .Y(_01717_),
    .A1(_01607_),
    .A2(_01687_));
 sg13g2_nand2_1 _07857_ (.Y(_01718_),
    .A(_01661_),
    .B(_01663_));
 sg13g2_a21oi_1 _07858_ (.A1(_01664_),
    .A2(_01683_),
    .Y(_01719_),
    .B1(_01682_));
 sg13g2_nor2_1 _07859_ (.A(_01674_),
    .B(_01676_),
    .Y(_01720_));
 sg13g2_nand2_1 _07860_ (.Y(_01721_),
    .A(net4460),
    .B(net4467));
 sg13g2_xnor2_1 _07861_ (.Y(_01722_),
    .A(_01720_),
    .B(_01721_));
 sg13g2_nand2_1 _07862_ (.Y(_01723_),
    .A(net4464),
    .B(\cpu.ALU.b[7] ));
 sg13g2_nand2_1 _07863_ (.Y(_01724_),
    .A(net4462),
    .B(\cpu.ALU.b[6] ));
 sg13g2_xor2_1 _07864_ (.B(_01724_),
    .A(_01723_),
    .X(_01725_));
 sg13g2_nand2_1 _07865_ (.Y(_01726_),
    .A(\cpu.ALU.b[2] ),
    .B(net4454));
 sg13g2_xnor2_1 _07866_ (.Y(_01727_),
    .A(_01673_),
    .B(_01726_));
 sg13g2_xnor2_1 _07867_ (.Y(_01728_),
    .A(_01725_),
    .B(_01727_));
 sg13g2_nand2_1 _07868_ (.Y(_01729_),
    .A(net4469),
    .B(net4456));
 sg13g2_xor2_1 _07869_ (.B(_01729_),
    .A(_01537_),
    .X(_01730_));
 sg13g2_xnor2_1 _07870_ (.Y(_01731_),
    .A(_01728_),
    .B(_01730_));
 sg13g2_xnor2_1 _07871_ (.Y(_01732_),
    .A(_01722_),
    .B(_01731_));
 sg13g2_o21ai_1 _07872_ (.B1(_01669_),
    .Y(_01733_),
    .A1(_01498_),
    .A2(_01537_));
 sg13g2_o21ai_1 _07873_ (.B1(_01679_),
    .Y(_01734_),
    .A1(_01670_),
    .A2(_01680_));
 sg13g2_xnor2_1 _07874_ (.Y(_01735_),
    .A(_01733_),
    .B(_01734_));
 sg13g2_xnor2_1 _07875_ (.Y(_01736_),
    .A(_01732_),
    .B(_01735_));
 sg13g2_xor2_1 _07876_ (.B(_01736_),
    .A(_01719_),
    .X(_01737_));
 sg13g2_xnor2_1 _07877_ (.Y(_01738_),
    .A(_01718_),
    .B(_01737_));
 sg13g2_xnor2_1 _07878_ (.Y(_01739_),
    .A(_01717_),
    .B(_01738_));
 sg13g2_xnor2_1 _07879_ (.Y(_01740_),
    .A(_01716_),
    .B(_01739_));
 sg13g2_nand2_1 _07880_ (.Y(_01741_),
    .A(\cpu.ALU.a[8] ),
    .B(\cpu.ALU.b[8] ));
 sg13g2_xor2_1 _07881_ (.B(\cpu.ALU.b[8] ),
    .A(\cpu.ALU.a[8] ),
    .X(_01742_));
 sg13g2_xnor2_1 _07882_ (.Y(_01743_),
    .A(\cpu.ALU.a[8] ),
    .B(\cpu.ALU.b[8] ));
 sg13g2_nand3_1 _07883_ (.B(_01700_),
    .C(_01743_),
    .A(_01693_),
    .Y(_01744_));
 sg13g2_a21o_1 _07884_ (.A2(_01700_),
    .A1(_01693_),
    .B1(_01743_),
    .X(_01745_));
 sg13g2_nand3_1 _07885_ (.B(_01744_),
    .C(_01745_),
    .A(net4027),
    .Y(_01746_));
 sg13g2_nor2b_1 _07886_ (.A(\cpu.ALU.b[7] ),
    .B_N(net4453),
    .Y(_01747_));
 sg13g2_a21oi_1 _07887_ (.A1(_01694_),
    .A2(_01697_),
    .Y(_01748_),
    .B1(_01747_));
 sg13g2_or2_1 _07888_ (.X(_01749_),
    .B(_01748_),
    .A(_01742_));
 sg13g2_a21oi_1 _07889_ (.A1(_01742_),
    .A2(_01748_),
    .Y(_01750_),
    .B1(net4025));
 sg13g2_nand2_1 _07890_ (.Y(_01751_),
    .A(_01749_),
    .B(_01750_));
 sg13g2_nand2_1 _07891_ (.Y(_01752_),
    .A(\cpu.ALU.a[9] ),
    .B(net4029));
 sg13g2_a22oi_1 _07892_ (.Y(_01753_),
    .B1(_01741_),
    .B2(net4028),
    .A2(net4144),
    .A1(net4453));
 sg13g2_nand4_1 _07893_ (.B(_01751_),
    .C(_01752_),
    .A(_01746_),
    .Y(_01754_),
    .D(_01753_));
 sg13g2_a21o_2 _07894_ (.A2(_01740_),
    .A1(_01351_),
    .B1(_01754_),
    .X(_01755_));
 sg13g2_nand2b_2 _07895_ (.Y(_01756_),
    .B(net3865),
    .A_N(_01755_));
 sg13g2_mux2_1 _07896_ (.A0(_00179_),
    .A1(net4297),
    .S(net3849),
    .X(_01757_));
 sg13g2_a21oi_1 _07897_ (.A1(net4045),
    .A2(_01757_),
    .Y(_01758_),
    .B1(net4251));
 sg13g2_nand2_1 _07898_ (.Y(_01759_),
    .A(_01756_),
    .B(_01758_));
 sg13g2_o21ai_1 _07899_ (.B1(net4146),
    .Y(_01760_),
    .A1(net4440),
    .A2(net4031));
 sg13g2_a21oi_2 _07900_ (.B1(_01760_),
    .Y(_01761_),
    .A2(net4031),
    .A1(_01153_));
 sg13g2_nor2_1 _07901_ (.A(net4225),
    .B(_01757_),
    .Y(_01762_));
 sg13g2_nor3_1 _07902_ (.A(net3623),
    .B(_01761_),
    .C(_01762_),
    .Y(_01763_));
 sg13g2_a22oi_1 _07903_ (.Y(_00271_),
    .B1(_01759_),
    .B2(_01763_),
    .A2(net3623),
    .A1(_00960_));
 sg13g2_nand2_1 _07904_ (.Y(_01764_),
    .A(\cpu.ALU.a[9] ),
    .B(\cpu.ALU.b[9] ));
 sg13g2_xor2_1 _07905_ (.B(\cpu.ALU.b[9] ),
    .A(\cpu.ALU.a[9] ),
    .X(_01765_));
 sg13g2_xnor2_1 _07906_ (.Y(_01766_),
    .A(\cpu.ALU.a[9] ),
    .B(\cpu.ALU.b[9] ));
 sg13g2_nand2b_1 _07907_ (.Y(_01767_),
    .B(\cpu.ALU.a[8] ),
    .A_N(\cpu.ALU.b[8] ));
 sg13g2_nand3_1 _07908_ (.B(_01765_),
    .C(_01767_),
    .A(_01749_),
    .Y(_01768_));
 sg13g2_or3_1 _07909_ (.A(_01742_),
    .B(_01748_),
    .C(_01765_),
    .X(_01769_));
 sg13g2_nor2_1 _07910_ (.A(_01765_),
    .B(_01767_),
    .Y(_01770_));
 sg13g2_nor2_1 _07911_ (.A(net4025),
    .B(_01770_),
    .Y(_01771_));
 sg13g2_nand3_1 _07912_ (.B(_01769_),
    .C(_01771_),
    .A(_01768_),
    .Y(_01772_));
 sg13g2_nand3_1 _07913_ (.B(_01745_),
    .C(_01766_),
    .A(_01741_),
    .Y(_01773_));
 sg13g2_nand2b_1 _07914_ (.Y(_01774_),
    .B(_01765_),
    .A_N(_01745_));
 sg13g2_nand2b_1 _07915_ (.Y(_01775_),
    .B(_01765_),
    .A_N(_01741_));
 sg13g2_nand4_1 _07916_ (.B(_01773_),
    .C(_01774_),
    .A(net4026),
    .Y(_01776_),
    .D(_01775_));
 sg13g2_nand2_1 _07917_ (.Y(_01777_),
    .A(\cpu.ALU.a[10] ),
    .B(net4029));
 sg13g2_a22oi_1 _07918_ (.Y(_01778_),
    .B1(_01764_),
    .B2(net4028),
    .A2(net4144),
    .A1(\cpu.ALU.a[8] ));
 sg13g2_and4_2 _07919_ (.A(_01772_),
    .B(_01776_),
    .C(_01777_),
    .D(_01778_),
    .X(_01779_));
 sg13g2_nand2_2 _07920_ (.Y(_01780_),
    .A(net3864),
    .B(_01779_));
 sg13g2_nor2_1 _07921_ (.A(_00183_),
    .B(net3849),
    .Y(_01781_));
 sg13g2_a21oi_1 _07922_ (.A1(_01176_),
    .A2(net3849),
    .Y(_01782_),
    .B1(_01781_));
 sg13g2_a21oi_1 _07923_ (.A1(net4048),
    .A2(_01782_),
    .Y(_01783_),
    .B1(net4256));
 sg13g2_nand2_1 _07924_ (.Y(_01784_),
    .A(_01780_),
    .B(_01783_));
 sg13g2_o21ai_1 _07925_ (.B1(net4146),
    .Y(_01785_),
    .A1(\cpu.current_address[9] ),
    .A2(_01264_));
 sg13g2_a21oi_2 _07926_ (.B1(_01785_),
    .Y(_01786_),
    .A2(_01264_),
    .A1(net4201));
 sg13g2_nor2_1 _07927_ (.A(net4227),
    .B(_01782_),
    .Y(_01787_));
 sg13g2_nor3_1 _07928_ (.A(net3624),
    .B(_01786_),
    .C(_01787_),
    .Y(_01788_));
 sg13g2_a22oi_1 _07929_ (.Y(_00272_),
    .B1(_01784_),
    .B2(_01788_),
    .A2(net3624),
    .A1(_00968_));
 sg13g2_nand2_1 _07930_ (.Y(_01789_),
    .A(\cpu.ALU.a[10] ),
    .B(\cpu.ALU.b[10] ));
 sg13g2_xor2_1 _07931_ (.B(\cpu.ALU.b[10] ),
    .A(\cpu.ALU.a[10] ),
    .X(_01790_));
 sg13g2_nand2_1 _07932_ (.Y(_01791_),
    .A(_01764_),
    .B(_01775_));
 sg13g2_inv_1 _07933_ (.Y(_01792_),
    .A(_01791_));
 sg13g2_o21ai_1 _07934_ (.B1(_01792_),
    .Y(_01793_),
    .A1(_01745_),
    .A2(_01766_));
 sg13g2_nand2_1 _07935_ (.Y(_01794_),
    .A(_01790_),
    .B(_01793_));
 sg13g2_xor2_1 _07936_ (.B(_01793_),
    .A(_01790_),
    .X(_01795_));
 sg13g2_a22oi_1 _07937_ (.Y(_01796_),
    .B1(_01789_),
    .B2(net4028),
    .A2(net4144),
    .A1(\cpu.ALU.a[9] ));
 sg13g2_o21ai_1 _07938_ (.B1(_01796_),
    .Y(_01797_),
    .A1(_01185_),
    .A2(_01344_));
 sg13g2_a21oi_1 _07939_ (.A1(\cpu.ALU.a[9] ),
    .A2(_01184_),
    .Y(_01798_),
    .B1(_01770_));
 sg13g2_nand3_1 _07940_ (.B(_01790_),
    .C(_01798_),
    .A(_01769_),
    .Y(_01799_));
 sg13g2_a21oi_1 _07941_ (.A1(_01769_),
    .A2(_01798_),
    .Y(_01800_),
    .B1(_01790_));
 sg13g2_nor2_1 _07942_ (.A(net4025),
    .B(_01800_),
    .Y(_01801_));
 sg13g2_a221oi_1 _07943_ (.B2(_01801_),
    .C1(_01797_),
    .B1(_01799_),
    .A1(net4026),
    .Y(_01802_),
    .A2(_01795_));
 sg13g2_nand2_2 _07944_ (.Y(_01803_),
    .A(net3862),
    .B(_01802_));
 sg13g2_nor2_1 _07945_ (.A(_00187_),
    .B(net3848),
    .Y(_01804_));
 sg13g2_a21oi_1 _07946_ (.A1(_01177_),
    .A2(net3848),
    .Y(_01805_),
    .B1(_01804_));
 sg13g2_a21oi_1 _07947_ (.A1(net4043),
    .A2(_01805_),
    .Y(_01806_),
    .B1(net4246));
 sg13g2_nand2_1 _07948_ (.Y(_01807_),
    .A(_01803_),
    .B(_01806_));
 sg13g2_o21ai_1 _07949_ (.B1(net4146),
    .Y(_01808_),
    .A1(net4432),
    .A2(net4032));
 sg13g2_a21oi_2 _07950_ (.B1(_01808_),
    .Y(_01809_),
    .A2(net4031),
    .A1(_01155_));
 sg13g2_nor2_1 _07951_ (.A(net4224),
    .B(_01805_),
    .Y(_01810_));
 sg13g2_nor3_1 _07952_ (.A(net3622),
    .B(_01809_),
    .C(_01810_),
    .Y(_01811_));
 sg13g2_a22oi_1 _07953_ (.Y(_00273_),
    .B1(_01807_),
    .B2(_01811_),
    .A2(net3622),
    .A1(_00976_));
 sg13g2_nand2_1 _07954_ (.Y(_01812_),
    .A(\cpu.ALU.a[11] ),
    .B(\cpu.ALU.b[11] ));
 sg13g2_xor2_1 _07955_ (.B(\cpu.ALU.b[11] ),
    .A(\cpu.ALU.a[11] ),
    .X(_01813_));
 sg13g2_xnor2_1 _07956_ (.Y(_01814_),
    .A(\cpu.ALU.a[11] ),
    .B(\cpu.ALU.b[11] ));
 sg13g2_nand2b_1 _07957_ (.Y(_01815_),
    .B(\cpu.ALU.a[10] ),
    .A_N(\cpu.ALU.b[10] ));
 sg13g2_nor2b_1 _07958_ (.A(_01800_),
    .B_N(_01815_),
    .Y(_01816_));
 sg13g2_a21oi_1 _07959_ (.A1(_01813_),
    .A2(_01816_),
    .Y(_01817_),
    .B1(net4025));
 sg13g2_o21ai_1 _07960_ (.B1(_01817_),
    .Y(_01818_),
    .A1(_01813_),
    .A2(_01816_));
 sg13g2_nand3_1 _07961_ (.B(_01794_),
    .C(_01814_),
    .A(_01789_),
    .Y(_01819_));
 sg13g2_nand2b_1 _07962_ (.Y(_01820_),
    .B(_01813_),
    .A_N(_01789_));
 sg13g2_nand3_1 _07963_ (.B(_01793_),
    .C(_01813_),
    .A(_01790_),
    .Y(_01821_));
 sg13g2_nand4_1 _07964_ (.B(_01819_),
    .C(_01820_),
    .A(net4026),
    .Y(_01822_),
    .D(_01821_));
 sg13g2_nand2_1 _07965_ (.Y(_01823_),
    .A(\cpu.ALU.a[10] ),
    .B(net4144));
 sg13g2_a22oi_1 _07966_ (.Y(_01824_),
    .B1(net4028),
    .B2(_01812_),
    .A2(net4029),
    .A1(\cpu.ALU.a[12] ));
 sg13g2_and4_2 _07967_ (.A(_01818_),
    .B(_01822_),
    .C(_01823_),
    .D(_01824_),
    .X(_01825_));
 sg13g2_nand2_2 _07968_ (.Y(_01826_),
    .A(net3863),
    .B(_01825_));
 sg13g2_mux2_1 _07969_ (.A0(_00191_),
    .A1(net4285),
    .S(net3848),
    .X(_01827_));
 sg13g2_a21oi_1 _07970_ (.A1(net4046),
    .A2(_01827_),
    .Y(_01828_),
    .B1(net4252));
 sg13g2_nand2_1 _07971_ (.Y(_01829_),
    .A(_01826_),
    .B(_01828_));
 sg13g2_o21ai_1 _07972_ (.B1(net4146),
    .Y(_01830_),
    .A1(net4431),
    .A2(net4032));
 sg13g2_a21oi_2 _07973_ (.B1(_01830_),
    .Y(_01831_),
    .A2(net4031),
    .A1(_01157_));
 sg13g2_nor2_1 _07974_ (.A(net4229),
    .B(_01827_),
    .Y(_01832_));
 sg13g2_nor3_1 _07975_ (.A(net3623),
    .B(_01831_),
    .C(_01832_),
    .Y(_01833_));
 sg13g2_a22oi_1 _07976_ (.Y(_00274_),
    .B1(_01829_),
    .B2(_01833_),
    .A2(net3623),
    .A1(_00984_));
 sg13g2_and2_1 _07977_ (.A(\cpu.ALU.a[12] ),
    .B(\cpu.ALU.b[12] ),
    .X(_01834_));
 sg13g2_xnor2_1 _07978_ (.Y(_01835_),
    .A(\cpu.ALU.a[12] ),
    .B(\cpu.ALU.b[12] ));
 sg13g2_and2_1 _07979_ (.A(_01812_),
    .B(_01820_),
    .X(_01836_));
 sg13g2_a21oi_1 _07980_ (.A1(_01821_),
    .A2(_01836_),
    .Y(_01837_),
    .B1(_01835_));
 sg13g2_nand3_1 _07981_ (.B(_01835_),
    .C(_01836_),
    .A(_01821_),
    .Y(_01838_));
 sg13g2_nand2_1 _07982_ (.Y(_01839_),
    .A(net4026),
    .B(_01838_));
 sg13g2_or3_1 _07983_ (.A(_01765_),
    .B(_01790_),
    .C(_01813_),
    .X(_01840_));
 sg13g2_o21ai_1 _07984_ (.B1(_01815_),
    .Y(_01841_),
    .A1(_01790_),
    .A2(_01798_));
 sg13g2_nor2_1 _07985_ (.A(_01185_),
    .B(\cpu.ALU.b[11] ),
    .Y(_01842_));
 sg13g2_a21oi_1 _07986_ (.A1(_01814_),
    .A2(_01841_),
    .Y(_01843_),
    .B1(_01842_));
 sg13g2_o21ai_1 _07987_ (.B1(_01843_),
    .Y(_01844_),
    .A1(_01749_),
    .A2(_01840_));
 sg13g2_nand2_1 _07988_ (.Y(_01845_),
    .A(_01835_),
    .B(_01844_));
 sg13g2_nor2_1 _07989_ (.A(_01835_),
    .B(_01844_),
    .Y(_01846_));
 sg13g2_nor2_1 _07990_ (.A(net4025),
    .B(_01846_),
    .Y(_01847_));
 sg13g2_a22oi_1 _07991_ (.Y(_01848_),
    .B1(net4144),
    .B2(\cpu.ALU.a[11] ),
    .A2(net4029),
    .A1(\cpu.ALU.a[13] ));
 sg13g2_o21ai_1 _07992_ (.B1(_01848_),
    .Y(_01849_),
    .A1(_01354_),
    .A2(_01834_));
 sg13g2_a21oi_1 _07993_ (.A1(_01845_),
    .A2(_01847_),
    .Y(_01850_),
    .B1(_01849_));
 sg13g2_o21ai_1 _07994_ (.B1(_01850_),
    .Y(_01851_),
    .A1(_01837_),
    .A2(_01839_));
 sg13g2_nand2b_2 _07995_ (.Y(_01852_),
    .B(net3864),
    .A_N(_01851_));
 sg13g2_mux2_1 _07996_ (.A0(_00195_),
    .A1(net4280),
    .S(net3849),
    .X(_01853_));
 sg13g2_a21oi_1 _07997_ (.A1(net4047),
    .A2(_01853_),
    .Y(_01854_),
    .B1(net4255));
 sg13g2_nor2_1 _07998_ (.A(net4227),
    .B(_01853_),
    .Y(_01855_));
 sg13g2_o21ai_1 _07999_ (.B1(net4146),
    .Y(_01856_),
    .A1(net4412),
    .A2(net4032));
 sg13g2_a21oi_2 _08000_ (.B1(_01856_),
    .Y(_01857_),
    .A2(net4032),
    .A1(_01159_));
 sg13g2_a21oi_1 _08001_ (.A1(_01852_),
    .A2(_01854_),
    .Y(_01858_),
    .B1(_01855_));
 sg13g2_nor2_1 _08002_ (.A(net3624),
    .B(_01857_),
    .Y(_01859_));
 sg13g2_a22oi_1 _08003_ (.Y(_00275_),
    .B1(_01858_),
    .B2(_01859_),
    .A2(net3624),
    .A1(_00992_));
 sg13g2_nand2_1 _08004_ (.Y(_01860_),
    .A(\cpu.ALU.a[13] ),
    .B(\cpu.ALU.b[13] ));
 sg13g2_xor2_1 _08005_ (.B(\cpu.ALU.b[13] ),
    .A(\cpu.ALU.a[13] ),
    .X(_01861_));
 sg13g2_xnor2_1 _08006_ (.Y(_01862_),
    .A(\cpu.ALU.a[13] ),
    .B(\cpu.ALU.b[13] ));
 sg13g2_o21ai_1 _08007_ (.B1(_01861_),
    .Y(_01863_),
    .A1(_01834_),
    .A2(_01837_));
 sg13g2_nor3_1 _08008_ (.A(_01834_),
    .B(_01837_),
    .C(_01861_),
    .Y(_01864_));
 sg13g2_nor2b_1 _08009_ (.A(_01864_),
    .B_N(net4026),
    .Y(_01865_));
 sg13g2_a22oi_1 _08010_ (.Y(_01866_),
    .B1(_01860_),
    .B2(net4028),
    .A2(net4144),
    .A1(\cpu.ALU.a[12] ));
 sg13g2_o21ai_1 _08011_ (.B1(_01866_),
    .Y(_01867_),
    .A1(_00201_),
    .A2(_01344_));
 sg13g2_o21ai_1 _08012_ (.B1(_01845_),
    .Y(_01868_),
    .A1(_01188_),
    .A2(\cpu.ALU.b[12] ));
 sg13g2_xnor2_1 _08013_ (.Y(_01869_),
    .A(_01861_),
    .B(_01868_));
 sg13g2_a221oi_1 _08014_ (.B2(_01390_),
    .C1(_01867_),
    .B1(_01869_),
    .A1(_01863_),
    .Y(_01870_),
    .A2(_01865_));
 sg13g2_nand2_2 _08015_ (.Y(_01871_),
    .A(net3862),
    .B(_01870_));
 sg13g2_nor2_1 _08016_ (.A(_00199_),
    .B(net3848),
    .Y(_01872_));
 sg13g2_a21oi_1 _08017_ (.A1(_01178_),
    .A2(net3848),
    .Y(_01873_),
    .B1(_01872_));
 sg13g2_a21oi_1 _08018_ (.A1(net4042),
    .A2(_01873_),
    .Y(_01874_),
    .B1(net4249));
 sg13g2_nand2_1 _08019_ (.Y(_01875_),
    .A(_01871_),
    .B(_01874_));
 sg13g2_o21ai_1 _08020_ (.B1(net4146),
    .Y(_01876_),
    .A1(net4396),
    .A2(net4031));
 sg13g2_a21oi_2 _08021_ (.B1(_01876_),
    .Y(_01877_),
    .A2(net4031),
    .A1(_01161_));
 sg13g2_nor2_1 _08022_ (.A(net4223),
    .B(_01873_),
    .Y(_01878_));
 sg13g2_nor3_1 _08023_ (.A(net3622),
    .B(_01877_),
    .C(_01878_),
    .Y(_01879_));
 sg13g2_a22oi_1 _08024_ (.Y(_00276_),
    .B1(_01875_),
    .B2(_01879_),
    .A2(net3622),
    .A1(_01114_));
 sg13g2_nand2_1 _08025_ (.Y(_01880_),
    .A(\cpu.ALU.a[14] ),
    .B(\cpu.ALU.b[14] ));
 sg13g2_inv_1 _08026_ (.Y(_01881_),
    .A(_01880_));
 sg13g2_nor2_1 _08027_ (.A(\cpu.ALU.a[14] ),
    .B(\cpu.ALU.b[14] ),
    .Y(_01882_));
 sg13g2_nor2_2 _08028_ (.A(_01881_),
    .B(_01882_),
    .Y(_01883_));
 sg13g2_and2_1 _08029_ (.A(_01860_),
    .B(_01863_),
    .X(_01884_));
 sg13g2_xnor2_1 _08030_ (.Y(_01885_),
    .A(_01883_),
    .B(_01884_));
 sg13g2_a22oi_1 _08031_ (.Y(_01886_),
    .B1(net4144),
    .B2(\cpu.ALU.a[13] ),
    .A2(net4029),
    .A1(\cpu.ALU.a[15] ));
 sg13g2_o21ai_1 _08032_ (.B1(_01886_),
    .Y(_01887_),
    .A1(_01354_),
    .A2(_01881_));
 sg13g2_nor2b_1 _08033_ (.A(\cpu.ALU.b[13] ),
    .B_N(\cpu.ALU.a[13] ),
    .Y(_01888_));
 sg13g2_a21oi_2 _08034_ (.B1(_01888_),
    .Y(_01889_),
    .A2(_01868_),
    .A1(_01862_));
 sg13g2_xor2_1 _08035_ (.B(_01889_),
    .A(_01883_),
    .X(_01890_));
 sg13g2_a221oi_1 _08036_ (.B2(_01390_),
    .C1(_01887_),
    .B1(_01890_),
    .A1(net4026),
    .Y(_01891_),
    .A2(_01885_));
 sg13g2_nand2_2 _08037_ (.Y(_01892_),
    .A(net3862),
    .B(_01891_));
 sg13g2_nor2_1 _08038_ (.A(_00204_),
    .B(net3848),
    .Y(_01893_));
 sg13g2_a21oi_1 _08039_ (.A1(_01179_),
    .A2(net3848),
    .Y(_01894_),
    .B1(_01893_));
 sg13g2_a21oi_1 _08040_ (.A1(net4043),
    .A2(_01894_),
    .Y(_01895_),
    .B1(net4246));
 sg13g2_nand2_1 _08041_ (.Y(_01896_),
    .A(_01892_),
    .B(_01895_));
 sg13g2_o21ai_1 _08042_ (.B1(net4146),
    .Y(_01897_),
    .A1(\cpu.current_address[14] ),
    .A2(_01264_));
 sg13g2_a21oi_2 _08043_ (.B1(_01897_),
    .Y(_01898_),
    .A2(_01264_),
    .A1(net4215));
 sg13g2_nor2_1 _08044_ (.A(net4221),
    .B(_01894_),
    .Y(_01899_));
 sg13g2_nor3_1 _08045_ (.A(net3622),
    .B(_01898_),
    .C(_01899_),
    .Y(_01900_));
 sg13g2_a22oi_1 _08046_ (.Y(_00277_),
    .B1(_01896_),
    .B2(_01900_),
    .A2(net3622),
    .A1(_01129_));
 sg13g2_nor2_1 _08047_ (.A(_01191_),
    .B(\cpu.ALU.b[15] ),
    .Y(_01901_));
 sg13g2_xnor2_1 _08048_ (.Y(_01902_),
    .A(\cpu.ALU.a[15] ),
    .B(\cpu.ALU.b[15] ));
 sg13g2_o21ai_1 _08049_ (.B1(_01880_),
    .Y(_01903_),
    .A1(_01882_),
    .A2(_01884_));
 sg13g2_xnor2_1 _08050_ (.Y(_01904_),
    .A(_01902_),
    .B(_01903_));
 sg13g2_nor2b_1 _08051_ (.A(_00201_),
    .B_N(net4144),
    .Y(_01905_));
 sg13g2_a21oi_1 _08052_ (.A1(\cpu.ALU.a[15] ),
    .A2(\cpu.ALU.b[15] ),
    .Y(_01906_),
    .B1(_01354_));
 sg13g2_or2_1 _08053_ (.X(_01907_),
    .B(_01906_),
    .A(_01905_));
 sg13g2_nand2b_1 _08054_ (.Y(_01908_),
    .B(\cpu.ALU.a[14] ),
    .A_N(\cpu.ALU.b[14] ));
 sg13g2_o21ai_1 _08055_ (.B1(_01908_),
    .Y(_01909_),
    .A1(_01883_),
    .A2(_01889_));
 sg13g2_xor2_1 _08056_ (.B(_01909_),
    .A(_01902_),
    .X(_01910_));
 sg13g2_a221oi_1 _08057_ (.B2(_01390_),
    .C1(_01907_),
    .B1(_01910_),
    .A1(net4026),
    .Y(_01911_),
    .A2(_01904_));
 sg13g2_nand2_2 _08058_ (.Y(_01912_),
    .A(net3862),
    .B(_01911_));
 sg13g2_mux2_1 _08059_ (.A0(_00208_),
    .A1(_00145_),
    .S(net3848),
    .X(_01913_));
 sg13g2_a21oi_1 _08060_ (.A1(net4042),
    .A2(_01913_),
    .Y(_01914_),
    .B1(net4248));
 sg13g2_nand2_1 _08061_ (.Y(_01915_),
    .A(_01912_),
    .B(_01914_));
 sg13g2_o21ai_1 _08062_ (.B1(net4146),
    .Y(_01916_),
    .A1(net4368),
    .A2(net4031));
 sg13g2_a21oi_2 _08063_ (.B1(_01916_),
    .Y(_01917_),
    .A2(net4031),
    .A1(_01164_));
 sg13g2_nor2_1 _08064_ (.A(net4223),
    .B(_01913_),
    .Y(_01918_));
 sg13g2_nor3_1 _08065_ (.A(net3622),
    .B(_01917_),
    .C(_01918_),
    .Y(_01919_));
 sg13g2_a22oi_1 _08066_ (.Y(_00278_),
    .B1(_01915_),
    .B2(_01919_),
    .A2(net3622),
    .A1(_01142_));
 sg13g2_nand3_1 _08067_ (.B(net4396),
    .C(_00025_),
    .A(net4380),
    .Y(_01920_));
 sg13g2_nand2_1 _08068_ (.Y(_01921_),
    .A(_01420_),
    .B(net4135));
 sg13g2_nand2_2 _08069_ (.Y(_01922_),
    .A(net4450),
    .B(net4448));
 sg13g2_inv_1 _08070_ (.Y(_01923_),
    .A(_01922_));
 sg13g2_nor2_2 _08071_ (.A(\cpu.current_instruction[6] ),
    .B(_01922_),
    .Y(_01924_));
 sg13g2_inv_1 _08072_ (.Y(_01925_),
    .A(net3996));
 sg13g2_and2_1 _08073_ (.A(net4308),
    .B(_01264_),
    .X(_01926_));
 sg13g2_nor2b_2 _08074_ (.A(net4312),
    .B_N(_01437_),
    .Y(_01927_));
 sg13g2_nand3_1 _08075_ (.B(\cpu.current_instruction[6] ),
    .C(_00024_),
    .A(net4448),
    .Y(_01928_));
 sg13g2_a22oi_1 _08076_ (.Y(_01929_),
    .B1(_01927_),
    .B2(_01928_),
    .A2(_01926_),
    .A1(_01925_));
 sg13g2_nand4_1 _08077_ (.B(_01432_),
    .C(_01921_),
    .A(_01423_),
    .Y(_01930_),
    .D(_01929_));
 sg13g2_nor2_1 _08078_ (.A(_01170_),
    .B(net4137),
    .Y(_01931_));
 sg13g2_a221oi_1 _08079_ (.B2(_00211_),
    .C1(_01931_),
    .B1(net4137),
    .A1(net4233),
    .Y(_01932_),
    .A2(_01409_));
 sg13g2_nor2_1 _08080_ (.A(net3620),
    .B(_01932_),
    .Y(_01933_));
 sg13g2_a22oi_1 _08081_ (.Y(_00279_),
    .B1(_01933_),
    .B2(_01443_),
    .A2(net3620),
    .A1(_00907_));
 sg13g2_mux2_1 _08082_ (.A0(net4361),
    .A1(_00212_),
    .S(net4137),
    .X(_01934_));
 sg13g2_nor2_1 _08083_ (.A(_01451_),
    .B(_01934_),
    .Y(_01935_));
 sg13g2_nor3_1 _08084_ (.A(_01448_),
    .B(net3621),
    .C(_01935_),
    .Y(_01936_));
 sg13g2_a21oi_1 _08085_ (.A1(_00911_),
    .A2(net3620),
    .Y(_00280_),
    .B1(_01936_));
 sg13g2_mux2_1 _08086_ (.A0(net4353),
    .A1(_00213_),
    .S(net4137),
    .X(_01937_));
 sg13g2_nor2_1 _08087_ (.A(_01477_),
    .B(_01937_),
    .Y(_01938_));
 sg13g2_nor3_1 _08088_ (.A(_01481_),
    .B(net3620),
    .C(_01938_),
    .Y(_01939_));
 sg13g2_a21oi_1 _08089_ (.A1(_00917_),
    .A2(net3620),
    .Y(_00281_),
    .B1(_01939_));
 sg13g2_nor2_1 _08090_ (.A(_01171_),
    .B(net4136),
    .Y(_01940_));
 sg13g2_a21oi_1 _08091_ (.A1(_00214_),
    .A2(net4136),
    .Y(_01941_),
    .B1(_01940_));
 sg13g2_o21ai_1 _08092_ (.B1(_01511_),
    .Y(_01942_),
    .A1(net3868),
    .A2(_01941_));
 sg13g2_a21oi_1 _08093_ (.A1(net4299),
    .A2(_01941_),
    .Y(_01943_),
    .B1(_01516_));
 sg13g2_nor2b_1 _08094_ (.A(net3619),
    .B_N(_01943_),
    .Y(_01944_));
 sg13g2_a22oi_1 _08095_ (.Y(_00282_),
    .B1(_01942_),
    .B2(_01944_),
    .A2(net3619),
    .A1(_00925_));
 sg13g2_nand2_1 _08096_ (.Y(_01945_),
    .A(_00215_),
    .B(net4136));
 sg13g2_o21ai_1 _08097_ (.B1(_01945_),
    .Y(_01946_),
    .A1(net4156),
    .A2(net4136));
 sg13g2_a21oi_1 _08098_ (.A1(net4056),
    .A2(_01946_),
    .Y(_01947_),
    .B1(_01552_));
 sg13g2_nor2_1 _08099_ (.A(net4235),
    .B(_01946_),
    .Y(_01948_));
 sg13g2_nor4_1 _08100_ (.A(_01556_),
    .B(net3619),
    .C(_01947_),
    .D(_01948_),
    .Y(_01949_));
 sg13g2_a21oi_1 _08101_ (.A1(_00931_),
    .A2(net3619),
    .Y(_00283_),
    .B1(_01949_));
 sg13g2_nand2_1 _08102_ (.Y(_01950_),
    .A(_00216_),
    .B(net4136));
 sg13g2_o21ai_1 _08103_ (.B1(_01950_),
    .Y(_01951_),
    .A1(_01173_),
    .A2(net4136));
 sg13g2_a21oi_1 _08104_ (.A1(net4054),
    .A2(_01951_),
    .Y(_01952_),
    .B1(net4260));
 sg13g2_nand2_1 _08105_ (.Y(_01953_),
    .A(_01596_),
    .B(_01952_));
 sg13g2_nor2_1 _08106_ (.A(net4234),
    .B(_01951_),
    .Y(_01954_));
 sg13g2_nor3_1 _08107_ (.A(_01601_),
    .B(net3619),
    .C(_01954_),
    .Y(_01955_));
 sg13g2_a22oi_1 _08108_ (.Y(_00284_),
    .B1(_01953_),
    .B2(_01955_),
    .A2(net3619),
    .A1(_00939_));
 sg13g2_nor2_1 _08109_ (.A(_01174_),
    .B(net4136),
    .Y(_01956_));
 sg13g2_a21oi_1 _08110_ (.A1(_00217_),
    .A2(net4136),
    .Y(_01957_),
    .B1(_01956_));
 sg13g2_o21ai_1 _08111_ (.B1(net4321),
    .Y(_01958_),
    .A1(net3868),
    .A2(_01957_));
 sg13g2_inv_1 _08112_ (.Y(_01959_),
    .A(_01958_));
 sg13g2_a221oi_1 _08113_ (.B2(_01649_),
    .C1(net3619),
    .B1(_01959_),
    .A1(net4299),
    .Y(_01960_),
    .A2(_01957_));
 sg13g2_a22oi_1 _08114_ (.Y(_00285_),
    .B1(_01960_),
    .B2(_01654_),
    .A2(net3619),
    .A1(_00946_));
 sg13g2_nand2_1 _08115_ (.Y(_01961_),
    .A(_00218_),
    .B(net4137));
 sg13g2_o21ai_1 _08116_ (.B1(_01961_),
    .Y(_01962_),
    .A1(_01175_),
    .A2(net4137));
 sg13g2_a21oi_1 _08117_ (.A1(net4052),
    .A2(_01962_),
    .Y(_01963_),
    .B1(net4259));
 sg13g2_nand2_1 _08118_ (.Y(_01964_),
    .A(_01707_),
    .B(_01963_));
 sg13g2_nor2_1 _08119_ (.A(net4231),
    .B(_01962_),
    .Y(_01965_));
 sg13g2_nor3_1 _08120_ (.A(_01713_),
    .B(net3620),
    .C(_01965_),
    .Y(_01966_));
 sg13g2_a22oi_1 _08121_ (.Y(_00286_),
    .B1(_01964_),
    .B2(_01966_),
    .A2(net3620),
    .A1(_00954_));
 sg13g2_mux2_1 _08122_ (.A0(net4298),
    .A1(_00219_),
    .S(net4134),
    .X(_01967_));
 sg13g2_a21oi_1 _08123_ (.A1(net4044),
    .A2(_01967_),
    .Y(_01968_),
    .B1(net4251));
 sg13g2_nand2_1 _08124_ (.Y(_01969_),
    .A(_01756_),
    .B(_01968_));
 sg13g2_nor2_1 _08125_ (.A(net4225),
    .B(_01967_),
    .Y(_01970_));
 sg13g2_nor3_1 _08126_ (.A(_01761_),
    .B(net3618),
    .C(_01970_),
    .Y(_01971_));
 sg13g2_a22oi_1 _08127_ (.Y(_00287_),
    .B1(_01969_),
    .B2(_01971_),
    .A2(net3618),
    .A1(_00961_));
 sg13g2_nand2_1 _08128_ (.Y(_01972_),
    .A(_00220_),
    .B(net4135));
 sg13g2_o21ai_1 _08129_ (.B1(_01972_),
    .Y(_01973_),
    .A1(net4154),
    .A2(net4135));
 sg13g2_a21oi_1 _08130_ (.A1(net4048),
    .A2(_01973_),
    .Y(_01974_),
    .B1(net4256));
 sg13g2_nand2_1 _08131_ (.Y(_01975_),
    .A(_01780_),
    .B(_01974_));
 sg13g2_nor2_1 _08132_ (.A(net4228),
    .B(_01973_),
    .Y(_01976_));
 sg13g2_nor3_1 _08133_ (.A(_01786_),
    .B(net3618),
    .C(_01976_),
    .Y(_01977_));
 sg13g2_a22oi_1 _08134_ (.Y(_00288_),
    .B1(_01975_),
    .B2(_01977_),
    .A2(net3618),
    .A1(_00969_));
 sg13g2_nand2_1 _08135_ (.Y(_01978_),
    .A(_00221_),
    .B(net4134));
 sg13g2_o21ai_1 _08136_ (.B1(_01978_),
    .Y(_01979_),
    .A1(net4153),
    .A2(net4134));
 sg13g2_a21oi_1 _08137_ (.A1(net4040),
    .A2(_01979_),
    .Y(_01980_),
    .B1(net4246));
 sg13g2_nand2_1 _08138_ (.Y(_01981_),
    .A(_01803_),
    .B(_01980_));
 sg13g2_nor2_1 _08139_ (.A(net4221),
    .B(_01979_),
    .Y(_01982_));
 sg13g2_nor3_1 _08140_ (.A(_01809_),
    .B(net3617),
    .C(_01982_),
    .Y(_01983_));
 sg13g2_a22oi_1 _08141_ (.Y(_00289_),
    .B1(_01981_),
    .B2(_01983_),
    .A2(net3617),
    .A1(_00977_));
 sg13g2_mux2_1 _08142_ (.A0(net4284),
    .A1(_00222_),
    .S(net4135),
    .X(_01984_));
 sg13g2_a21oi_1 _08143_ (.A1(net4046),
    .A2(_01984_),
    .Y(_01985_),
    .B1(net4252));
 sg13g2_nand2_1 _08144_ (.Y(_01986_),
    .A(_01826_),
    .B(_01985_));
 sg13g2_nor2_1 _08145_ (.A(net4229),
    .B(_01984_),
    .Y(_01987_));
 sg13g2_nor3_1 _08146_ (.A(_01831_),
    .B(net3621),
    .C(_01987_),
    .Y(_01988_));
 sg13g2_a22oi_1 _08147_ (.Y(_00290_),
    .B1(_01986_),
    .B2(_01988_),
    .A2(net3618),
    .A1(_00985_));
 sg13g2_mux2_1 _08148_ (.A0(net4280),
    .A1(_00223_),
    .S(net4135),
    .X(_01989_));
 sg13g2_a21oi_1 _08149_ (.A1(net4047),
    .A2(_01989_),
    .Y(_01990_),
    .B1(net4255));
 sg13g2_nand2_1 _08150_ (.Y(_01991_),
    .A(_01852_),
    .B(_01990_));
 sg13g2_nor2_1 _08151_ (.A(net4227),
    .B(_01989_),
    .Y(_01992_));
 sg13g2_nor3_1 _08152_ (.A(_01857_),
    .B(net3618),
    .C(_01992_),
    .Y(_01993_));
 sg13g2_a22oi_1 _08153_ (.Y(_00291_),
    .B1(_01991_),
    .B2(_01993_),
    .A2(net3618),
    .A1(_00993_));
 sg13g2_nand2_1 _08154_ (.Y(_01994_),
    .A(_00224_),
    .B(net4134));
 sg13g2_o21ai_1 _08155_ (.B1(_01994_),
    .Y(_01995_),
    .A1(_01178_),
    .A2(net4134));
 sg13g2_a21oi_1 _08156_ (.A1(net4041),
    .A2(_01995_),
    .Y(_01996_),
    .B1(net4247));
 sg13g2_nand2_1 _08157_ (.Y(_01997_),
    .A(_01871_),
    .B(_01996_));
 sg13g2_nor2_1 _08158_ (.A(net4222),
    .B(_01995_),
    .Y(_01998_));
 sg13g2_nor3_1 _08159_ (.A(_01877_),
    .B(net3617),
    .C(_01998_),
    .Y(_01999_));
 sg13g2_a22oi_1 _08160_ (.Y(_00292_),
    .B1(_01997_),
    .B2(_01999_),
    .A2(net3617),
    .A1(_01115_));
 sg13g2_nand2_1 _08161_ (.Y(_02000_),
    .A(_00225_),
    .B(net4134));
 sg13g2_o21ai_1 _08162_ (.B1(_02000_),
    .Y(_02001_),
    .A1(_01179_),
    .A2(net4134));
 sg13g2_a21oi_1 _08163_ (.A1(net4040),
    .A2(_02001_),
    .Y(_02002_),
    .B1(net4247));
 sg13g2_nand2_1 _08164_ (.Y(_02003_),
    .A(_01892_),
    .B(_02002_));
 sg13g2_nor2_1 _08165_ (.A(net4221),
    .B(_02001_),
    .Y(_02004_));
 sg13g2_nor3_1 _08166_ (.A(_01898_),
    .B(net3617),
    .C(_02004_),
    .Y(_02005_));
 sg13g2_a22oi_1 _08167_ (.Y(_00293_),
    .B1(_02003_),
    .B2(_02005_),
    .A2(net3617),
    .A1(_01130_));
 sg13g2_mux2_1 _08168_ (.A0(net4268),
    .A1(_00226_),
    .S(net4134),
    .X(_02006_));
 sg13g2_a21oi_1 _08169_ (.A1(net4041),
    .A2(_02006_),
    .Y(_02007_),
    .B1(net4248));
 sg13g2_nand2_1 _08170_ (.Y(_02008_),
    .A(_01912_),
    .B(_02007_));
 sg13g2_nor2_1 _08171_ (.A(net4222),
    .B(_02006_),
    .Y(_02009_));
 sg13g2_nor3_1 _08172_ (.A(_01917_),
    .B(net3617),
    .C(_02009_),
    .Y(_02010_));
 sg13g2_a22oi_1 _08173_ (.Y(_00294_),
    .B1(_02008_),
    .B2(_02010_),
    .A2(net3617),
    .A1(_01143_));
 sg13g2_nor3_2 _08174_ (.A(net4217),
    .B(net4396),
    .C(_00897_),
    .Y(_02011_));
 sg13g2_mux2_1 _08175_ (.A0(_00049_),
    .A1(net4365),
    .S(net3994),
    .X(_02012_));
 sg13g2_nand2b_1 _08176_ (.Y(_02013_),
    .B(_01420_),
    .A_N(net3992));
 sg13g2_nand2_1 _08177_ (.Y(_02014_),
    .A(_00024_),
    .B(_01433_));
 sg13g2_and2_1 _08178_ (.A(net4239),
    .B(_01336_),
    .X(_02015_));
 sg13g2_inv_1 _08179_ (.Y(_02016_),
    .A(net3988));
 sg13g2_a22oi_1 _08180_ (.Y(_02017_),
    .B1(_02016_),
    .B2(_01926_),
    .A2(_02014_),
    .A1(_01927_));
 sg13g2_nand4_1 _08181_ (.B(_01432_),
    .C(_02013_),
    .A(_01423_),
    .Y(_02018_),
    .D(_02017_));
 sg13g2_o21ai_1 _08182_ (.B1(_01443_),
    .Y(_02019_),
    .A1(_01410_),
    .A2(_02012_));
 sg13g2_mux2_1 _08183_ (.A0(_02019_),
    .A1(net518),
    .S(net3616),
    .X(_00295_));
 sg13g2_mux2_1 _08184_ (.A0(_00050_),
    .A1(net4362),
    .S(net3993),
    .X(_02020_));
 sg13g2_nor2_1 _08185_ (.A(_01451_),
    .B(_02020_),
    .Y(_02021_));
 sg13g2_nor3_1 _08186_ (.A(_01448_),
    .B(net3615),
    .C(_02021_),
    .Y(_02022_));
 sg13g2_a21oi_1 _08187_ (.A1(_00912_),
    .A2(net3615),
    .Y(_00296_),
    .B1(_02022_));
 sg13g2_nor2b_1 _08188_ (.A(net3994),
    .B_N(_00051_),
    .Y(_02023_));
 sg13g2_a221oi_1 _08189_ (.B2(net4353),
    .C1(_02023_),
    .B1(net3994),
    .A1(net4232),
    .Y(_02024_),
    .A2(_01476_));
 sg13g2_nor3_1 _08190_ (.A(_01481_),
    .B(net3616),
    .C(_02024_),
    .Y(_02025_));
 sg13g2_a21oi_1 _08191_ (.A1(_00918_),
    .A2(net3616),
    .Y(_00297_),
    .B1(_02025_));
 sg13g2_nor2b_1 _08192_ (.A(net3994),
    .B_N(_00052_),
    .Y(_02026_));
 sg13g2_a21oi_1 _08193_ (.A1(net4351),
    .A2(net3993),
    .Y(_02027_),
    .B1(_02026_));
 sg13g2_o21ai_1 _08194_ (.B1(_01511_),
    .Y(_02028_),
    .A1(net3868),
    .A2(_02027_));
 sg13g2_a21oi_1 _08195_ (.A1(net4300),
    .A2(_02027_),
    .Y(_02029_),
    .B1(_01516_));
 sg13g2_nor2b_1 _08196_ (.A(net3615),
    .B_N(_02029_),
    .Y(_02030_));
 sg13g2_a22oi_1 _08197_ (.Y(_00298_),
    .B1(_02028_),
    .B2(_02030_),
    .A2(net3615),
    .A1(_00926_));
 sg13g2_nor2_1 _08198_ (.A(_00053_),
    .B(net3993),
    .Y(_02031_));
 sg13g2_a21oi_1 _08199_ (.A1(_01172_),
    .A2(net3993),
    .Y(_02032_),
    .B1(_02031_));
 sg13g2_a21oi_1 _08200_ (.A1(net4057),
    .A2(_02032_),
    .Y(_02033_),
    .B1(_01552_));
 sg13g2_or2_1 _08201_ (.X(_02034_),
    .B(_02032_),
    .A(net4235));
 sg13g2_nor3_1 _08202_ (.A(_01556_),
    .B(net3615),
    .C(_02033_),
    .Y(_02035_));
 sg13g2_a22oi_1 _08203_ (.Y(_00299_),
    .B1(_02034_),
    .B2(_02035_),
    .A2(net3615),
    .A1(_00932_));
 sg13g2_nor2_1 _08204_ (.A(_00054_),
    .B(net3993),
    .Y(_02036_));
 sg13g2_a21oi_1 _08205_ (.A1(_01173_),
    .A2(net3993),
    .Y(_02037_),
    .B1(_02036_));
 sg13g2_a21oi_1 _08206_ (.A1(net4054),
    .A2(_02037_),
    .Y(_02038_),
    .B1(net4261));
 sg13g2_nand2_1 _08207_ (.Y(_02039_),
    .A(_01596_),
    .B(_02038_));
 sg13g2_nor2_1 _08208_ (.A(net4234),
    .B(_02037_),
    .Y(_02040_));
 sg13g2_nor3_1 _08209_ (.A(_01601_),
    .B(net3615),
    .C(_02040_),
    .Y(_02041_));
 sg13g2_a22oi_1 _08210_ (.Y(_00300_),
    .B1(_02039_),
    .B2(_02041_),
    .A2(net3615),
    .A1(_00940_));
 sg13g2_nor2_1 _08211_ (.A(_00055_),
    .B(net3993),
    .Y(_02042_));
 sg13g2_a21oi_1 _08212_ (.A1(net4155),
    .A2(net3993),
    .Y(_02043_),
    .B1(_02042_));
 sg13g2_a21oi_1 _08213_ (.A1(net4056),
    .A2(_02043_),
    .Y(_02044_),
    .B1(net4262));
 sg13g2_nand2_1 _08214_ (.Y(_02045_),
    .A(_01649_),
    .B(_02044_));
 sg13g2_o21ai_1 _08215_ (.B1(_01654_),
    .Y(_02046_),
    .A1(net4235),
    .A2(_02043_));
 sg13g2_nor2_1 _08216_ (.A(net3616),
    .B(_02046_),
    .Y(_02047_));
 sg13g2_a22oi_1 _08217_ (.Y(_00301_),
    .B1(_02045_),
    .B2(_02047_),
    .A2(net3616),
    .A1(_00947_));
 sg13g2_nor2_1 _08218_ (.A(_00056_),
    .B(net3994),
    .Y(_02048_));
 sg13g2_a21oi_1 _08219_ (.A1(_01175_),
    .A2(net3994),
    .Y(_02049_),
    .B1(_02048_));
 sg13g2_a21oi_1 _08220_ (.A1(net4052),
    .A2(_02049_),
    .Y(_02050_),
    .B1(net4259));
 sg13g2_nand2_1 _08221_ (.Y(_02051_),
    .A(_01707_),
    .B(_02050_));
 sg13g2_nor2_1 _08222_ (.A(net4232),
    .B(_02049_),
    .Y(_02052_));
 sg13g2_nor3_1 _08223_ (.A(_01713_),
    .B(net3616),
    .C(_02052_),
    .Y(_02053_));
 sg13g2_a22oi_1 _08224_ (.Y(_00302_),
    .B1(_02051_),
    .B2(_02053_),
    .A2(net3616),
    .A1(_00955_));
 sg13g2_mux2_1 _08225_ (.A0(_00057_),
    .A1(net4298),
    .S(net3991),
    .X(_02054_));
 sg13g2_a21oi_1 _08226_ (.A1(net4044),
    .A2(_02054_),
    .Y(_02055_),
    .B1(net4251));
 sg13g2_nand2_1 _08227_ (.Y(_02056_),
    .A(_01756_),
    .B(_02055_));
 sg13g2_nor2_1 _08228_ (.A(net4225),
    .B(_02054_),
    .Y(_02057_));
 sg13g2_nor3_1 _08229_ (.A(_01761_),
    .B(net3612),
    .C(_02057_),
    .Y(_02058_));
 sg13g2_a22oi_1 _08230_ (.Y(_00303_),
    .B1(_02056_),
    .B2(_02058_),
    .A2(net3612),
    .A1(_00962_));
 sg13g2_nor2_1 _08231_ (.A(_00058_),
    .B(net3992),
    .Y(_02059_));
 sg13g2_a21oi_1 _08232_ (.A1(net4154),
    .A2(net3992),
    .Y(_02060_),
    .B1(_02059_));
 sg13g2_a21oi_1 _08233_ (.A1(net4048),
    .A2(_02060_),
    .Y(_02061_),
    .B1(net4256));
 sg13g2_nand2_1 _08234_ (.Y(_02062_),
    .A(_01780_),
    .B(_02061_));
 sg13g2_nor2_1 _08235_ (.A(net4228),
    .B(_02060_),
    .Y(_02063_));
 sg13g2_nor3_1 _08236_ (.A(_01786_),
    .B(net3614),
    .C(_02063_),
    .Y(_02064_));
 sg13g2_a22oi_1 _08237_ (.Y(_00304_),
    .B1(_02062_),
    .B2(_02064_),
    .A2(net3614),
    .A1(_00970_));
 sg13g2_nor2_1 _08238_ (.A(_00059_),
    .B(net3991),
    .Y(_02065_));
 sg13g2_a21oi_1 _08239_ (.A1(net4153),
    .A2(net3991),
    .Y(_02066_),
    .B1(_02065_));
 sg13g2_a21oi_1 _08240_ (.A1(net4044),
    .A2(_02066_),
    .Y(_02067_),
    .B1(net4250));
 sg13g2_nand2_1 _08241_ (.Y(_02068_),
    .A(_01803_),
    .B(_02067_));
 sg13g2_nor2_1 _08242_ (.A(net4225),
    .B(_02066_),
    .Y(_02069_));
 sg13g2_nor3_1 _08243_ (.A(_01809_),
    .B(net3612),
    .C(_02069_),
    .Y(_02070_));
 sg13g2_a22oi_1 _08244_ (.Y(_00305_),
    .B1(_02068_),
    .B2(_02070_),
    .A2(net3612),
    .A1(_00978_));
 sg13g2_mux2_1 _08245_ (.A0(_00060_),
    .A1(net4285),
    .S(net3992),
    .X(_02071_));
 sg13g2_a21oi_1 _08246_ (.A1(net4046),
    .A2(_02071_),
    .Y(_02072_),
    .B1(net4251));
 sg13g2_nand2_1 _08247_ (.Y(_02073_),
    .A(_01826_),
    .B(_02072_));
 sg13g2_nor2_1 _08248_ (.A(net4229),
    .B(_02071_),
    .Y(_02074_));
 sg13g2_nor3_1 _08249_ (.A(_01831_),
    .B(net3613),
    .C(_02074_),
    .Y(_02075_));
 sg13g2_a22oi_1 _08250_ (.Y(_00306_),
    .B1(_02073_),
    .B2(_02075_),
    .A2(net3613),
    .A1(_00986_));
 sg13g2_mux2_1 _08251_ (.A0(_00061_),
    .A1(_00142_),
    .S(net3992),
    .X(_02076_));
 sg13g2_a21oi_1 _08252_ (.A1(net4047),
    .A2(_02076_),
    .Y(_02077_),
    .B1(net4256));
 sg13g2_nor2_1 _08253_ (.A(net4227),
    .B(_02076_),
    .Y(_02078_));
 sg13g2_a21oi_1 _08254_ (.A1(_01852_),
    .A2(_02077_),
    .Y(_02079_),
    .B1(_02078_));
 sg13g2_nor2_1 _08255_ (.A(_01857_),
    .B(net3614),
    .Y(_02080_));
 sg13g2_a22oi_1 _08256_ (.Y(_00307_),
    .B1(_02079_),
    .B2(_02080_),
    .A2(net3614),
    .A1(_00994_));
 sg13g2_nor2_1 _08257_ (.A(_00062_),
    .B(net3991),
    .Y(_02081_));
 sg13g2_a21oi_1 _08258_ (.A1(_01178_),
    .A2(net3991),
    .Y(_02082_),
    .B1(_02081_));
 sg13g2_a21oi_1 _08259_ (.A1(net4045),
    .A2(_02082_),
    .Y(_02083_),
    .B1(net4249));
 sg13g2_nand2_1 _08260_ (.Y(_02084_),
    .A(_01871_),
    .B(_02083_));
 sg13g2_nor2_1 _08261_ (.A(net4226),
    .B(_02082_),
    .Y(_02085_));
 sg13g2_nor3_1 _08262_ (.A(_01877_),
    .B(net3613),
    .C(_02085_),
    .Y(_02086_));
 sg13g2_a22oi_1 _08263_ (.Y(_00308_),
    .B1(_02084_),
    .B2(_02086_),
    .A2(net3613),
    .A1(_01116_));
 sg13g2_nor2_1 _08264_ (.A(_00063_),
    .B(net3991),
    .Y(_02087_));
 sg13g2_a21oi_1 _08265_ (.A1(net4151),
    .A2(net3991),
    .Y(_02088_),
    .B1(_02087_));
 sg13g2_a21oi_1 _08266_ (.A1(net4044),
    .A2(_02088_),
    .Y(_02089_),
    .B1(net4249));
 sg13g2_nand2_1 _08267_ (.Y(_02090_),
    .A(_01892_),
    .B(_02089_));
 sg13g2_nor2_1 _08268_ (.A(net4226),
    .B(_02088_),
    .Y(_02091_));
 sg13g2_nor3_1 _08269_ (.A(_01898_),
    .B(net3612),
    .C(_02091_),
    .Y(_02092_));
 sg13g2_a22oi_1 _08270_ (.Y(_00309_),
    .B1(_02090_),
    .B2(_02092_),
    .A2(net3612),
    .A1(_01131_));
 sg13g2_mux2_1 _08271_ (.A0(_00064_),
    .A1(net4268),
    .S(net3991),
    .X(_02093_));
 sg13g2_a21o_1 _08272_ (.A2(_02093_),
    .A1(net4045),
    .B1(net4249),
    .X(_02094_));
 sg13g2_a21oi_1 _08273_ (.A1(net3862),
    .A2(_01911_),
    .Y(_02095_),
    .B1(_02094_));
 sg13g2_nor2_1 _08274_ (.A(net4226),
    .B(_02093_),
    .Y(_02096_));
 sg13g2_nor4_1 _08275_ (.A(_01917_),
    .B(net3612),
    .C(_02095_),
    .D(_02096_),
    .Y(_02097_));
 sg13g2_a21oi_1 _08276_ (.A1(_01144_),
    .A2(net3612),
    .Y(_00310_),
    .B1(_02097_));
 sg13g2_a221oi_1 _08277_ (.B2(net4148),
    .C1(_01427_),
    .B1(_01436_),
    .A1(_01250_),
    .Y(_02098_),
    .A2(_01418_));
 sg13g2_nand3_1 _08278_ (.B(_01424_),
    .C(_02098_),
    .A(_01423_),
    .Y(_02099_));
 sg13g2_mux2_1 _08279_ (.A0(net4353),
    .A1(_00156_),
    .S(net3853),
    .X(_02100_));
 sg13g2_nor2_1 _08280_ (.A(net3865),
    .B(_02100_),
    .Y(_02101_));
 sg13g2_nand4_1 _08281_ (.B(_01540_),
    .C(_01585_),
    .A(_01499_),
    .Y(_02102_),
    .D(_01636_));
 sg13g2_nor3_1 _08282_ (.A(_01347_),
    .B(_01465_),
    .C(_02102_),
    .Y(_02103_));
 sg13g2_nand4_1 _08283_ (.B(_01743_),
    .C(_01835_),
    .A(_01694_),
    .Y(_02104_),
    .D(_01862_));
 sg13g2_nor3_1 _08284_ (.A(_01392_),
    .B(_01840_),
    .C(_02104_),
    .Y(_02105_));
 sg13g2_nand3b_1 _08285_ (.B(_02103_),
    .C(_02105_),
    .Y(_02106_),
    .A_N(_01890_));
 sg13g2_o21ai_1 _08286_ (.B1(net3865),
    .Y(_02107_),
    .A1(_01910_),
    .A2(_02106_));
 sg13g2_a21oi_1 _08287_ (.A1(_01191_),
    .A2(\cpu.ALU.b[15] ),
    .Y(_02108_),
    .B1(_01909_));
 sg13g2_nor3_2 _08288_ (.A(_01901_),
    .B(_02107_),
    .C(_02108_),
    .Y(_02109_));
 sg13g2_o21ai_1 _08289_ (.B1(net4317),
    .Y(_02110_),
    .A1(_02101_),
    .A2(_02109_));
 sg13g2_o21ai_1 _08290_ (.B1(_01480_),
    .Y(_02111_),
    .A1(net4232),
    .A2(_02100_));
 sg13g2_nor2_1 _08291_ (.A(_02099_),
    .B(_02111_),
    .Y(_02112_));
 sg13g2_a22oi_1 _08292_ (.Y(_00311_),
    .B1(_02110_),
    .B2(_02112_),
    .A2(_02099_),
    .A1(_00919_));
 sg13g2_nor2_1 _08293_ (.A(_00160_),
    .B(_01339_),
    .Y(_02113_));
 sg13g2_a21oi_1 _08294_ (.A1(_01171_),
    .A2(net3855),
    .Y(_02114_),
    .B1(_02113_));
 sg13g2_inv_1 _08295_ (.Y(_02115_),
    .A(_02114_));
 sg13g2_a21oi_1 _08296_ (.A1(net4056),
    .A2(_02114_),
    .Y(_02116_),
    .B1(net4263));
 sg13g2_nand2_1 _08297_ (.Y(_02117_),
    .A(net179),
    .B(_02099_));
 sg13g2_a221oi_1 _08298_ (.B2(_02107_),
    .C1(_01516_),
    .B1(_02116_),
    .A1(net4300),
    .Y(_02118_),
    .A2(_02115_));
 sg13g2_o21ai_1 _08299_ (.B1(_02117_),
    .Y(_00312_),
    .A1(_02099_),
    .A2(_02118_));
 sg13g2_nor2_1 _08300_ (.A(_00164_),
    .B(_01339_),
    .Y(_02119_));
 sg13g2_a21oi_1 _08301_ (.A1(net4156),
    .A2(net3854),
    .Y(_02120_),
    .B1(_02119_));
 sg13g2_nor2_1 _08302_ (.A(net3867),
    .B(_02120_),
    .Y(_02121_));
 sg13g2_nor4_1 _08303_ (.A(_01356_),
    .B(_01395_),
    .C(_01475_),
    .D(_01509_),
    .Y(_02122_));
 sg13g2_and3_1 _08304_ (.X(_02123_),
    .A(_01551_),
    .B(_01595_),
    .C(_02122_));
 sg13g2_and4_1 _08305_ (.A(_01648_),
    .B(_01706_),
    .C(_01779_),
    .D(_02123_),
    .X(_02124_));
 sg13g2_nand3_1 _08306_ (.B(_01825_),
    .C(_02124_),
    .A(_01802_),
    .Y(_02125_));
 sg13g2_nor3_1 _08307_ (.A(_01756_),
    .B(_01851_),
    .C(_02125_),
    .Y(_02126_));
 sg13g2_and4_2 _08308_ (.A(_01870_),
    .B(_01891_),
    .C(_01911_),
    .D(_02126_),
    .X(_02127_));
 sg13g2_o21ai_1 _08309_ (.B1(net4319),
    .Y(_02128_),
    .A1(_02121_),
    .A2(_02127_));
 sg13g2_nor2_1 _08310_ (.A(net4235),
    .B(_02120_),
    .Y(_02129_));
 sg13g2_nor3_1 _08311_ (.A(_01556_),
    .B(_02099_),
    .C(_02129_),
    .Y(_02130_));
 sg13g2_a22oi_1 _08312_ (.Y(_00313_),
    .B1(_02128_),
    .B2(_02130_),
    .A2(_02099_),
    .A1(_00933_));
 sg13g2_nand2_1 _08313_ (.Y(_02131_),
    .A(net4065),
    .B(_01418_));
 sg13g2_nor2_1 _08314_ (.A(_00152_),
    .B(net3998),
    .Y(_02132_));
 sg13g2_nor2_2 _08315_ (.A(_00026_),
    .B(_01922_),
    .Y(_02133_));
 sg13g2_or2_1 _08316_ (.X(_02134_),
    .B(_01922_),
    .A(_00026_));
 sg13g2_nand2_1 _08317_ (.Y(_02135_),
    .A(\cpu.registers[1][3] ),
    .B(_02133_));
 sg13g2_o21ai_1 _08318_ (.B1(_02135_),
    .Y(_02136_),
    .A1(_00164_),
    .A2(net4148));
 sg13g2_nor3_1 _08319_ (.A(net4239),
    .B(net4449),
    .C(_00026_),
    .Y(_02137_));
 sg13g2_inv_1 _08320_ (.Y(_02138_),
    .A(net3983));
 sg13g2_a221oi_1 _08321_ (.B2(_00156_),
    .C1(_02132_),
    .B1(net3995),
    .A1(_00026_),
    .Y(_02139_),
    .A2(_01434_));
 sg13g2_a221oi_1 _08322_ (.B2(\cpu.registers[1][0] ),
    .C1(_02136_),
    .B1(net3984),
    .A1(\cpu.registers[1][2] ),
    .Y(_02140_),
    .A2(net3989));
 sg13g2_a221oi_1 _08323_ (.B2(_02140_),
    .C1(_02131_),
    .B1(_02139_),
    .A1(_00017_),
    .Y(_02141_),
    .A2(_01923_));
 sg13g2_a21o_1 _08324_ (.A2(_02131_),
    .A1(net204),
    .B1(_02141_),
    .X(_00314_));
 sg13g2_and2_2 _08325_ (.A(net4444),
    .B(net4441),
    .X(_02142_));
 sg13g2_nand2b_1 _08326_ (.Y(_02143_),
    .B(net4132),
    .A_N(_00030_));
 sg13g2_inv_2 _08327_ (.Y(_02144_),
    .A(net3982));
 sg13g2_nand2_1 _08328_ (.Y(_02145_),
    .A(\cpu.registers[7][0] ),
    .B(_02144_));
 sg13g2_nor2b_1 _08329_ (.A(net4441),
    .B_N(net4444),
    .Y(_02146_));
 sg13g2_nand2b_1 _08330_ (.Y(_02147_),
    .B(net4446),
    .A_N(net4442));
 sg13g2_nor2_1 _08331_ (.A(net4436),
    .B(_02147_),
    .Y(_02148_));
 sg13g2_nor2_1 _08332_ (.A(_00030_),
    .B(_02147_),
    .Y(_02149_));
 sg13g2_a22oi_1 _08333_ (.Y(_02150_),
    .B1(net3978),
    .B2(\cpu.registers[5][0] ),
    .A2(net3980),
    .A1(\cpu.registers[1][0] ));
 sg13g2_nor2b_2 _08334_ (.A(net4444),
    .B_N(net4441),
    .Y(_02151_));
 sg13g2_nor2b_1 _08335_ (.A(_00030_),
    .B_N(net4128),
    .Y(_02152_));
 sg13g2_and2_2 _08336_ (.A(net4201),
    .B(net4133),
    .X(_02153_));
 sg13g2_a22oi_1 _08337_ (.Y(_02154_),
    .B1(net3973),
    .B2(\cpu.registers[3][0] ),
    .A2(net3976),
    .A1(\cpu.registers[6][0] ));
 sg13g2_nor2_1 _08338_ (.A(net4444),
    .B(net4441),
    .Y(_02155_));
 sg13g2_or2_1 _08339_ (.X(_02156_),
    .B(net4441),
    .A(net4444));
 sg13g2_nor2_1 _08340_ (.A(_00030_),
    .B(net4123),
    .Y(_02157_));
 sg13g2_and2_1 _08341_ (.A(net4201),
    .B(net4129),
    .X(_02158_));
 sg13g2_a22oi_1 _08342_ (.Y(_02159_),
    .B1(net3970),
    .B2(\cpu.registers[2][0] ),
    .A2(net3972),
    .A1(\cpu.registers[4][0] ));
 sg13g2_and4_2 _08343_ (.A(_02145_),
    .B(_02150_),
    .C(_02154_),
    .D(_02159_),
    .X(_02160_));
 sg13g2_inv_1 _08344_ (.Y(_02161_),
    .A(_02160_));
 sg13g2_nand2_1 _08345_ (.Y(_02162_),
    .A(net460),
    .B(net3859));
 sg13g2_o21ai_1 _08346_ (.B1(_02162_),
    .Y(_00315_),
    .A1(net3858),
    .A2(_02160_));
 sg13g2_nor2_1 _08347_ (.A(_00031_),
    .B(net3982),
    .Y(_02163_));
 sg13g2_a221oi_1 _08348_ (.B2(\cpu.registers[4][1] ),
    .C1(_02163_),
    .B1(net3972),
    .A1(\cpu.registers[1][1] ),
    .Y(_02164_),
    .A2(net3980));
 sg13g2_a22oi_1 _08349_ (.Y(_02165_),
    .B1(net3974),
    .B2(\cpu.registers[3][1] ),
    .A2(net3976),
    .A1(\cpu.registers[6][1] ));
 sg13g2_a22oi_1 _08350_ (.Y(_02166_),
    .B1(net3970),
    .B2(\cpu.registers[2][1] ),
    .A2(net3978),
    .A1(\cpu.registers[5][1] ));
 sg13g2_and3_2 _08351_ (.X(_02167_),
    .A(_02164_),
    .B(_02165_),
    .C(_02166_));
 sg13g2_inv_1 _08352_ (.Y(_02168_),
    .A(_02167_));
 sg13g2_nand2_1 _08353_ (.Y(_02169_),
    .A(net311),
    .B(net3858));
 sg13g2_o21ai_1 _08354_ (.B1(_02169_),
    .Y(_00316_),
    .A1(net3859),
    .A2(_02167_));
 sg13g2_nor3_1 _08355_ (.A(_00030_),
    .B(_00915_),
    .C(_02147_),
    .Y(_02170_));
 sg13g2_a221oi_1 _08356_ (.B2(\cpu.registers[3][2] ),
    .C1(_02170_),
    .B1(net3974),
    .A1(\cpu.registers[1][2] ),
    .Y(_02171_),
    .A2(net3980));
 sg13g2_nand2_1 _08357_ (.Y(_02172_),
    .A(\cpu.registers[4][2] ),
    .B(net3972));
 sg13g2_or2_1 _08358_ (.X(_02173_),
    .B(net3982),
    .A(_00032_));
 sg13g2_a22oi_1 _08359_ (.Y(_02174_),
    .B1(net3970),
    .B2(\cpu.registers[2][2] ),
    .A2(net3976),
    .A1(\cpu.registers[6][2] ));
 sg13g2_and4_2 _08360_ (.A(_02171_),
    .B(_02172_),
    .C(_02173_),
    .D(_02174_),
    .X(_02175_));
 sg13g2_nand4_1 _08361_ (.B(_02172_),
    .C(_02173_),
    .A(_02171_),
    .Y(_02176_),
    .D(_02174_));
 sg13g2_nand2_1 _08362_ (.Y(_02177_),
    .A(net633),
    .B(net3858));
 sg13g2_o21ai_1 _08363_ (.B1(_02177_),
    .Y(_00317_),
    .A1(net3858),
    .A2(_02175_));
 sg13g2_a22oi_1 _08364_ (.Y(_02178_),
    .B1(net3972),
    .B2(\cpu.registers[4][3] ),
    .A2(net3978),
    .A1(\cpu.registers[5][3] ));
 sg13g2_o21ai_1 _08365_ (.B1(_02178_),
    .Y(_02179_),
    .A1(_00033_),
    .A2(net3982));
 sg13g2_a22oi_1 _08366_ (.Y(_02180_),
    .B1(net3970),
    .B2(\cpu.registers[2][3] ),
    .A2(net3974),
    .A1(\cpu.registers[3][3] ));
 sg13g2_a22oi_1 _08367_ (.Y(_02181_),
    .B1(net3976),
    .B2(\cpu.registers[6][3] ),
    .A2(net3980),
    .A1(\cpu.registers[1][3] ));
 sg13g2_nand2_1 _08368_ (.Y(_02182_),
    .A(_02180_),
    .B(_02181_));
 sg13g2_nor2_2 _08369_ (.A(_02179_),
    .B(_02182_),
    .Y(_02183_));
 sg13g2_inv_1 _08370_ (.Y(_02184_),
    .A(_02183_));
 sg13g2_nand2_1 _08371_ (.Y(_02185_),
    .A(net631),
    .B(net3858));
 sg13g2_o21ai_1 _08372_ (.B1(_02185_),
    .Y(_00318_),
    .A1(net3859),
    .A2(_02183_));
 sg13g2_a22oi_1 _08373_ (.Y(_02186_),
    .B1(net3970),
    .B2(\cpu.registers[2][4] ),
    .A2(net3972),
    .A1(\cpu.registers[4][4] ));
 sg13g2_o21ai_1 _08374_ (.B1(_02186_),
    .Y(_02187_),
    .A1(_00034_),
    .A2(net3982));
 sg13g2_a22oi_1 _08375_ (.Y(_02188_),
    .B1(net3978),
    .B2(\cpu.registers[5][4] ),
    .A2(net3980),
    .A1(\cpu.registers[1][4] ));
 sg13g2_a22oi_1 _08376_ (.Y(_02189_),
    .B1(net3974),
    .B2(\cpu.registers[3][4] ),
    .A2(net3976),
    .A1(\cpu.registers[6][4] ));
 sg13g2_nand2_1 _08377_ (.Y(_02190_),
    .A(_02188_),
    .B(_02189_));
 sg13g2_nor2_2 _08378_ (.A(_02187_),
    .B(_02190_),
    .Y(_02191_));
 sg13g2_inv_1 _08379_ (.Y(_02192_),
    .A(_02191_));
 sg13g2_nand2_1 _08380_ (.Y(_02193_),
    .A(net578),
    .B(net3858));
 sg13g2_o21ai_1 _08381_ (.B1(_02193_),
    .Y(_00319_),
    .A1(net3857),
    .A2(_02191_));
 sg13g2_nand2_1 _08382_ (.Y(_02194_),
    .A(\cpu.registers[2][5] ),
    .B(net3970));
 sg13g2_a22oi_1 _08383_ (.Y(_02195_),
    .B1(net3972),
    .B2(\cpu.registers[4][5] ),
    .A2(net3978),
    .A1(\cpu.registers[5][5] ));
 sg13g2_a22oi_1 _08384_ (.Y(_02196_),
    .B1(_02153_),
    .B2(\cpu.registers[3][5] ),
    .A2(_02144_),
    .A1(_00935_));
 sg13g2_a22oi_1 _08385_ (.Y(_02197_),
    .B1(net3976),
    .B2(\cpu.registers[6][5] ),
    .A2(net3980),
    .A1(\cpu.registers[1][5] ));
 sg13g2_and4_2 _08386_ (.A(_02194_),
    .B(_02195_),
    .C(_02196_),
    .D(_02197_),
    .X(_02198_));
 sg13g2_inv_1 _08387_ (.Y(_02199_),
    .A(_02198_));
 sg13g2_nand2_1 _08388_ (.Y(_02200_),
    .A(net242),
    .B(net3858));
 sg13g2_o21ai_1 _08389_ (.B1(_02200_),
    .Y(_00320_),
    .A1(net3858),
    .A2(_02198_));
 sg13g2_a22oi_1 _08390_ (.Y(_02201_),
    .B1(net3976),
    .B2(\cpu.registers[6][6] ),
    .A2(net3980),
    .A1(\cpu.registers[1][6] ));
 sg13g2_o21ai_1 _08391_ (.B1(_02201_),
    .Y(_02202_),
    .A1(_00036_),
    .A2(net3981));
 sg13g2_a22oi_1 _08392_ (.Y(_02203_),
    .B1(net3972),
    .B2(\cpu.registers[4][6] ),
    .A2(net3974),
    .A1(\cpu.registers[3][6] ));
 sg13g2_inv_1 _08393_ (.Y(_02204_),
    .A(_02203_));
 sg13g2_a221oi_1 _08394_ (.B2(\cpu.registers[2][6] ),
    .C1(_02204_),
    .B1(net3970),
    .A1(\cpu.registers[5][6] ),
    .Y(_02205_),
    .A2(net3978));
 sg13g2_nor2b_2 _08395_ (.A(_02202_),
    .B_N(_02205_),
    .Y(_02206_));
 sg13g2_inv_1 _08396_ (.Y(_02207_),
    .A(_02206_));
 sg13g2_nand2_1 _08397_ (.Y(_02208_),
    .A(net405),
    .B(net3857));
 sg13g2_o21ai_1 _08398_ (.B1(_02208_),
    .Y(_00321_),
    .A1(net3857),
    .A2(_02206_));
 sg13g2_a22oi_1 _08399_ (.Y(_02209_),
    .B1(net3970),
    .B2(\cpu.registers[2][7] ),
    .A2(net3976),
    .A1(\cpu.registers[6][7] ));
 sg13g2_o21ai_1 _08400_ (.B1(_02209_),
    .Y(_02210_),
    .A1(_00037_),
    .A2(net3981));
 sg13g2_a22oi_1 _08401_ (.Y(_02211_),
    .B1(_02153_),
    .B2(\cpu.registers[3][7] ),
    .A2(net3978),
    .A1(\cpu.registers[5][7] ));
 sg13g2_inv_1 _08402_ (.Y(_02212_),
    .A(_02211_));
 sg13g2_a221oi_1 _08403_ (.B2(\cpu.registers[4][7] ),
    .C1(_02212_),
    .B1(net3972),
    .A1(\cpu.registers[1][7] ),
    .Y(_02213_),
    .A2(net3980));
 sg13g2_nor2b_2 _08404_ (.A(_02210_),
    .B_N(_02213_),
    .Y(_02214_));
 sg13g2_inv_1 _08405_ (.Y(_02215_),
    .A(_02214_));
 sg13g2_nand2_1 _08406_ (.Y(_02216_),
    .A(net681),
    .B(net3857));
 sg13g2_o21ai_1 _08407_ (.B1(_02216_),
    .Y(_00322_),
    .A1(net3856),
    .A2(_02214_));
 sg13g2_a22oi_1 _08408_ (.Y(_02217_),
    .B1(net3973),
    .B2(\cpu.registers[3][8] ),
    .A2(net3975),
    .A1(\cpu.registers[6][8] ));
 sg13g2_o21ai_1 _08409_ (.B1(_02217_),
    .Y(_02218_),
    .A1(_00038_),
    .A2(net3981));
 sg13g2_a22oi_1 _08410_ (.Y(_02219_),
    .B1(net3969),
    .B2(\cpu.registers[2][8] ),
    .A2(net3977),
    .A1(\cpu.registers[5][8] ));
 sg13g2_a22oi_1 _08411_ (.Y(_02220_),
    .B1(net3971),
    .B2(\cpu.registers[4][8] ),
    .A2(net3979),
    .A1(\cpu.registers[1][8] ));
 sg13g2_nand2_1 _08412_ (.Y(_02221_),
    .A(_02219_),
    .B(_02220_));
 sg13g2_nor2_2 _08413_ (.A(_02218_),
    .B(_02221_),
    .Y(_02222_));
 sg13g2_inv_1 _08414_ (.Y(_02223_),
    .A(_02222_));
 sg13g2_nand2_1 _08415_ (.Y(_02224_),
    .A(net270),
    .B(net3857));
 sg13g2_o21ai_1 _08416_ (.B1(_02224_),
    .Y(_00323_),
    .A1(net3857),
    .A2(_02222_));
 sg13g2_nand2_1 _08417_ (.Y(_02225_),
    .A(\cpu.registers[4][9] ),
    .B(net3971));
 sg13g2_a22oi_1 _08418_ (.Y(_02226_),
    .B1(net3975),
    .B2(\cpu.registers[6][9] ),
    .A2(_02144_),
    .A1(_00965_));
 sg13g2_a22oi_1 _08419_ (.Y(_02227_),
    .B1(net3974),
    .B2(\cpu.registers[3][9] ),
    .A2(net3979),
    .A1(\cpu.registers[1][9] ));
 sg13g2_a22oi_1 _08420_ (.Y(_02228_),
    .B1(net3969),
    .B2(\cpu.registers[2][9] ),
    .A2(net3977),
    .A1(\cpu.registers[5][9] ));
 sg13g2_and4_2 _08421_ (.A(_02225_),
    .B(_02226_),
    .C(_02227_),
    .D(_02228_),
    .X(_02229_));
 sg13g2_inv_1 _08422_ (.Y(_02230_),
    .A(_02229_));
 sg13g2_nand2_1 _08423_ (.Y(_02231_),
    .A(net248),
    .B(net3856));
 sg13g2_o21ai_1 _08424_ (.B1(_02231_),
    .Y(_00324_),
    .A1(_01269_),
    .A2(_02229_));
 sg13g2_nor2_1 _08425_ (.A(_00040_),
    .B(net3981),
    .Y(_02232_));
 sg13g2_a221oi_1 _08426_ (.B2(\cpu.registers[3][10] ),
    .C1(_02232_),
    .B1(net3973),
    .A1(\cpu.registers[5][10] ),
    .Y(_02233_),
    .A2(net3977));
 sg13g2_a22oi_1 _08427_ (.Y(_02234_),
    .B1(net3971),
    .B2(\cpu.registers[4][10] ),
    .A2(net3975),
    .A1(\cpu.registers[6][10] ));
 sg13g2_a22oi_1 _08428_ (.Y(_02235_),
    .B1(net3969),
    .B2(\cpu.registers[2][10] ),
    .A2(net3979),
    .A1(\cpu.registers[1][10] ));
 sg13g2_and3_2 _08429_ (.X(_02236_),
    .A(_02233_),
    .B(_02234_),
    .C(_02235_));
 sg13g2_inv_1 _08430_ (.Y(_02237_),
    .A(_02236_));
 sg13g2_nand2_1 _08431_ (.Y(_02238_),
    .A(net409),
    .B(net3856));
 sg13g2_o21ai_1 _08432_ (.B1(_02238_),
    .Y(_00325_),
    .A1(net3856),
    .A2(_02236_));
 sg13g2_nand2_1 _08433_ (.Y(_02239_),
    .A(\cpu.registers[4][11] ),
    .B(net3971));
 sg13g2_a22oi_1 _08434_ (.Y(_02240_),
    .B1(net3977),
    .B2(\cpu.registers[5][11] ),
    .A2(net3979),
    .A1(\cpu.registers[1][11] ));
 sg13g2_a22oi_1 _08435_ (.Y(_02241_),
    .B1(net3975),
    .B2(\cpu.registers[6][11] ),
    .A2(_02144_),
    .A1(_00981_));
 sg13g2_a22oi_1 _08436_ (.Y(_02242_),
    .B1(net3969),
    .B2(\cpu.registers[2][11] ),
    .A2(net3973),
    .A1(\cpu.registers[3][11] ));
 sg13g2_and4_2 _08437_ (.A(_02239_),
    .B(_02240_),
    .C(_02241_),
    .D(_02242_),
    .X(_02243_));
 sg13g2_inv_1 _08438_ (.Y(_02244_),
    .A(_02243_));
 sg13g2_nand2_1 _08439_ (.Y(_02245_),
    .A(net127),
    .B(net3856));
 sg13g2_o21ai_1 _08440_ (.B1(_02245_),
    .Y(_00326_),
    .A1(net3856),
    .A2(_02243_));
 sg13g2_nor2_1 _08441_ (.A(_00042_),
    .B(net3981),
    .Y(_02246_));
 sg13g2_a221oi_1 _08442_ (.B2(\cpu.registers[3][12] ),
    .C1(_02246_),
    .B1(net3973),
    .A1(\cpu.registers[5][12] ),
    .Y(_02247_),
    .A2(net3977));
 sg13g2_a22oi_1 _08443_ (.Y(_02248_),
    .B1(net3975),
    .B2(\cpu.registers[6][12] ),
    .A2(net3979),
    .A1(\cpu.registers[1][12] ));
 sg13g2_a22oi_1 _08444_ (.Y(_02249_),
    .B1(net3969),
    .B2(\cpu.registers[2][12] ),
    .A2(net3971),
    .A1(\cpu.registers[4][12] ));
 sg13g2_and3_2 _08445_ (.X(_02250_),
    .A(_02247_),
    .B(_02248_),
    .C(_02249_));
 sg13g2_inv_1 _08446_ (.Y(_02251_),
    .A(_02250_));
 sg13g2_nand2_1 _08447_ (.Y(_02252_),
    .A(net41),
    .B(net3856));
 sg13g2_o21ai_1 _08448_ (.B1(_02252_),
    .Y(_00327_),
    .A1(net3856),
    .A2(_02250_));
 sg13g2_nor2_2 _08449_ (.A(net4312),
    .B(net4071),
    .Y(_02253_));
 sg13g2_nand4_1 _08450_ (.B(net4217),
    .C(net4208),
    .A(net4325),
    .Y(_02254_),
    .D(_02253_));
 sg13g2_nor2_2 _08451_ (.A(net4394),
    .B(net4418),
    .Y(_02255_));
 sg13g2_nor3_2 _08452_ (.A(net4443),
    .B(net4395),
    .C(net4418),
    .Y(_02256_));
 sg13g2_nand2_1 _08453_ (.Y(_02257_),
    .A(net4125),
    .B(_02255_));
 sg13g2_nand3_1 _08454_ (.B(net4125),
    .C(_02255_),
    .A(net4201),
    .Y(_02258_));
 sg13g2_nor2_1 _08455_ (.A(net4430),
    .B(net4433),
    .Y(_02259_));
 sg13g2_nor2_1 _08456_ (.A(net4432),
    .B(_02258_),
    .Y(_02260_));
 sg13g2_or4_2 _08457_ (.A(net4430),
    .B(net4432),
    .C(_02254_),
    .D(_02258_),
    .X(_02261_));
 sg13g2_nand2_1 _08458_ (.Y(_02262_),
    .A(net665),
    .B(net3767));
 sg13g2_o21ai_1 _08459_ (.B1(_02262_),
    .Y(_00328_),
    .A1(net4364),
    .A2(net3767));
 sg13g2_nand2_1 _08460_ (.Y(_02263_),
    .A(net331),
    .B(net3767));
 sg13g2_o21ai_1 _08461_ (.B1(_02263_),
    .Y(_00329_),
    .A1(net4358),
    .A2(net3767));
 sg13g2_nand2_1 _08462_ (.Y(_02264_),
    .A(net523),
    .B(net3767));
 sg13g2_o21ai_1 _08463_ (.B1(_02264_),
    .Y(_00330_),
    .A1(net4355),
    .A2(net3766));
 sg13g2_nor2_1 _08464_ (.A(_01171_),
    .B(net3767),
    .Y(_02265_));
 sg13g2_a21oi_1 _08465_ (.A1(_01017_),
    .A2(net3766),
    .Y(_00331_),
    .B1(_02265_));
 sg13g2_nor2_1 _08466_ (.A(net4156),
    .B(net3766),
    .Y(_02266_));
 sg13g2_a21oi_1 _08467_ (.A1(_01026_),
    .A2(net3766),
    .Y(_00332_),
    .B1(_02266_));
 sg13g2_nand2_1 _08468_ (.Y(_02267_),
    .A(net416),
    .B(net3766));
 sg13g2_o21ai_1 _08469_ (.B1(_02267_),
    .Y(_00333_),
    .A1(net4343),
    .A2(net3766));
 sg13g2_nand2_1 _08470_ (.Y(_02268_),
    .A(net651),
    .B(net3766));
 sg13g2_o21ai_1 _08471_ (.B1(_02268_),
    .Y(_00334_),
    .A1(net4340),
    .A2(net3766));
 sg13g2_nand2_1 _08472_ (.Y(_02269_),
    .A(net574),
    .B(net3765));
 sg13g2_o21ai_1 _08473_ (.B1(_02269_),
    .Y(_00335_),
    .A1(net4337),
    .A2(net3765));
 sg13g2_nand2_1 _08474_ (.Y(_02270_),
    .A(net613),
    .B(net3765));
 sg13g2_o21ai_1 _08475_ (.B1(_02270_),
    .Y(_00336_),
    .A1(net4294),
    .A2(net3765));
 sg13g2_nand2_1 _08476_ (.Y(_02271_),
    .A(net585),
    .B(net3763));
 sg13g2_o21ai_1 _08477_ (.B1(_02271_),
    .Y(_00337_),
    .A1(net4290),
    .A2(net3763));
 sg13g2_nand2_1 _08478_ (.Y(_02272_),
    .A(net557),
    .B(net3763));
 sg13g2_o21ai_1 _08479_ (.B1(_02272_),
    .Y(_00338_),
    .A1(net4286),
    .A2(net3763));
 sg13g2_nand2_1 _08480_ (.Y(_02273_),
    .A(net441),
    .B(net3764));
 sg13g2_o21ai_1 _08481_ (.B1(_02273_),
    .Y(_00339_),
    .A1(net4282),
    .A2(net3764));
 sg13g2_nand2_1 _08482_ (.Y(_02274_),
    .A(net582),
    .B(net3765));
 sg13g2_o21ai_1 _08483_ (.B1(_02274_),
    .Y(_00340_),
    .A1(net4277),
    .A2(net3765));
 sg13g2_nand2_1 _08484_ (.Y(_02275_),
    .A(net612),
    .B(net3763));
 sg13g2_o21ai_1 _08485_ (.B1(_02275_),
    .Y(_00341_),
    .A1(net4275),
    .A2(net3763));
 sg13g2_nand2_1 _08486_ (.Y(_02276_),
    .A(net564),
    .B(net3763));
 sg13g2_o21ai_1 _08487_ (.B1(_02276_),
    .Y(_00342_),
    .A1(net4273),
    .A2(net3763));
 sg13g2_nand2_1 _08488_ (.Y(_02277_),
    .A(net684),
    .B(net3764));
 sg13g2_o21ai_1 _08489_ (.B1(_02277_),
    .Y(_00343_),
    .A1(net4269),
    .A2(net3764));
 sg13g2_nand2_1 _08490_ (.Y(_02278_),
    .A(net4431),
    .B(net4433));
 sg13g2_xnor2_1 _08491_ (.Y(_02279_),
    .A(net4430),
    .B(_02260_));
 sg13g2_nor2b_1 _08492_ (.A(_00044_),
    .B_N(_02279_),
    .Y(_02280_));
 sg13g2_and2_1 _08493_ (.A(net4391),
    .B(net4412),
    .X(_02281_));
 sg13g2_nor4_2 _08494_ (.A(net4430),
    .B(_00044_),
    .C(_02255_),
    .Y(_02282_),
    .D(net4115));
 sg13g2_or4_2 _08495_ (.A(net4430),
    .B(_00044_),
    .C(_02255_),
    .D(net4115),
    .X(_02283_));
 sg13g2_nor2_1 _08496_ (.A(net4443),
    .B(net3966),
    .Y(_02284_));
 sg13g2_nand2b_2 _08497_ (.Y(_02285_),
    .B(net3968),
    .A_N(net4446));
 sg13g2_a21oi_2 _08498_ (.B1(net4432),
    .Y(_02286_),
    .A2(_02257_),
    .A1(net4436));
 sg13g2_nand2_2 _08499_ (.Y(_02287_),
    .A(_02258_),
    .B(_02286_));
 sg13g2_nor2_1 _08500_ (.A(_02254_),
    .B(_02287_),
    .Y(_02288_));
 sg13g2_xnor2_1 _08501_ (.Y(_02289_),
    .A(net4439),
    .B(_02256_));
 sg13g2_and2_2 _08502_ (.A(net3761),
    .B(_02289_),
    .X(_02290_));
 sg13g2_nand2_2 _08503_ (.Y(_02291_),
    .A(net3761),
    .B(_02289_));
 sg13g2_nand2_1 _08504_ (.Y(_02292_),
    .A(_02284_),
    .B(net3711));
 sg13g2_nor2_1 _08505_ (.A(_01170_),
    .B(net3694),
    .Y(_02293_));
 sg13g2_a21oi_1 _08506_ (.A1(_00996_),
    .A2(net3693),
    .Y(_00344_),
    .B1(_02293_));
 sg13g2_nor2_1 _08507_ (.A(net4358),
    .B(_02285_),
    .Y(_02294_));
 sg13g2_a22oi_1 _08508_ (.Y(_02295_),
    .B1(_02294_),
    .B2(net3710),
    .A2(net3693),
    .A1(net639));
 sg13g2_inv_1 _08509_ (.Y(_00345_),
    .A(_02295_));
 sg13g2_nand2_1 _08510_ (.Y(_02296_),
    .A(net178),
    .B(net3693));
 sg13g2_o21ai_1 _08511_ (.B1(_02296_),
    .Y(_00346_),
    .A1(net4356),
    .A2(net3693));
 sg13g2_nor2_1 _08512_ (.A(net4350),
    .B(_02285_),
    .Y(_02297_));
 sg13g2_a22oi_1 _08513_ (.Y(_02298_),
    .B1(_02297_),
    .B2(_02290_),
    .A2(net3693),
    .A1(net784));
 sg13g2_inv_1 _08514_ (.Y(_00347_),
    .A(_02298_));
 sg13g2_nand2_1 _08515_ (.Y(_02299_),
    .A(net528),
    .B(net3693));
 sg13g2_xnor2_1 _08516_ (.Y(_02300_),
    .A(net4443),
    .B(_02255_));
 sg13g2_xor2_1 _08517_ (.B(_02255_),
    .A(net4443),
    .X(_02301_));
 sg13g2_nand3_1 _08518_ (.B(net3968),
    .C(net3965),
    .A(net4156),
    .Y(_02302_));
 sg13g2_o21ai_1 _08519_ (.B1(_02299_),
    .Y(_00348_),
    .A1(_02291_),
    .A2(_02302_));
 sg13g2_nor4_2 _08520_ (.A(net4442),
    .B(net4343),
    .C(_02283_),
    .Y(_02303_),
    .D(net3963));
 sg13g2_a22oi_1 _08521_ (.Y(_02304_),
    .B1(_02303_),
    .B2(_02288_),
    .A2(net3693),
    .A1(net786));
 sg13g2_inv_1 _08522_ (.Y(_00349_),
    .A(_02304_));
 sg13g2_nor4_2 _08523_ (.A(net4442),
    .B(net4342),
    .C(_02283_),
    .Y(_02305_),
    .D(net3963));
 sg13g2_a22oi_1 _08524_ (.Y(_02306_),
    .B1(_02305_),
    .B2(net3762),
    .A2(net3693),
    .A1(net437));
 sg13g2_inv_1 _08525_ (.Y(_00350_),
    .A(net438));
 sg13g2_nor4_2 _08526_ (.A(net4441),
    .B(net4337),
    .C(_02283_),
    .Y(_02307_),
    .D(net3962));
 sg13g2_a22oi_1 _08527_ (.Y(_02308_),
    .B1(_02307_),
    .B2(net3762),
    .A2(net3692),
    .A1(net636));
 sg13g2_inv_1 _08528_ (.Y(_00351_),
    .A(_02308_));
 sg13g2_nor4_2 _08529_ (.A(net4439),
    .B(net4296),
    .C(net3966),
    .Y(_02309_),
    .D(_02301_));
 sg13g2_a22oi_1 _08530_ (.Y(_02310_),
    .B1(_02309_),
    .B2(net3762),
    .A2(net3692),
    .A1(net725));
 sg13g2_inv_1 _08531_ (.Y(_00352_),
    .A(_02310_));
 sg13g2_nand2_1 _08532_ (.Y(_02311_),
    .A(net586),
    .B(net3692));
 sg13g2_nand3_1 _08533_ (.B(net3967),
    .C(net3964),
    .A(net4154),
    .Y(_02312_));
 sg13g2_o21ai_1 _08534_ (.B1(_02311_),
    .Y(_00353_),
    .A1(net3707),
    .A2(_02312_));
 sg13g2_nand2_1 _08535_ (.Y(_02313_),
    .A(net671),
    .B(net3692));
 sg13g2_nand3_1 _08536_ (.B(net3967),
    .C(net3964),
    .A(net4153),
    .Y(_02314_));
 sg13g2_o21ai_1 _08537_ (.B1(_02313_),
    .Y(_00354_),
    .A1(net3707),
    .A2(_02314_));
 sg13g2_nand2_1 _08538_ (.Y(_02315_),
    .A(net741),
    .B(net3692));
 sg13g2_nand3b_1 _08539_ (.B(net3967),
    .C(net3964),
    .Y(_02316_),
    .A_N(net4283));
 sg13g2_o21ai_1 _08540_ (.B1(_02315_),
    .Y(_00355_),
    .A1(net3707),
    .A2(_02316_));
 sg13g2_nand3b_1 _08541_ (.B(net3968),
    .C(net3965),
    .Y(_02317_),
    .A_N(net4279));
 sg13g2_nand2_1 _08542_ (.Y(_02318_),
    .A(net699),
    .B(net3694));
 sg13g2_o21ai_1 _08543_ (.B1(_02318_),
    .Y(_00356_),
    .A1(_02291_),
    .A2(_02317_));
 sg13g2_nand2_1 _08544_ (.Y(_02319_),
    .A(net493),
    .B(net3692));
 sg13g2_nand3_1 _08545_ (.B(net3967),
    .C(net3964),
    .A(net4152),
    .Y(_02320_));
 sg13g2_o21ai_1 _08546_ (.B1(_02319_),
    .Y(_00357_),
    .A1(net3707),
    .A2(_02320_));
 sg13g2_nand3_1 _08547_ (.B(net3967),
    .C(net3964),
    .A(net4151),
    .Y(_02321_));
 sg13g2_nand2_1 _08548_ (.Y(_02322_),
    .A(net599),
    .B(net3692));
 sg13g2_o21ai_1 _08549_ (.B1(_02322_),
    .Y(_00358_),
    .A1(net3707),
    .A2(_02321_));
 sg13g2_nand2_1 _08550_ (.Y(_02323_),
    .A(net558),
    .B(net3692));
 sg13g2_nand3b_1 _08551_ (.B(net3967),
    .C(net3964),
    .Y(_02324_),
    .A_N(net4270));
 sg13g2_o21ai_1 _08552_ (.B1(_02323_),
    .Y(_00359_),
    .A1(net3708),
    .A2(_02324_));
 sg13g2_nor2b_1 _08553_ (.A(net4412),
    .B_N(net4391),
    .Y(_02325_));
 sg13g2_and2_2 _08554_ (.A(_02279_),
    .B(net4103),
    .X(_02326_));
 sg13g2_nand2_1 _08555_ (.Y(_02327_),
    .A(_02279_),
    .B(net4103));
 sg13g2_nor2_2 _08556_ (.A(net4443),
    .B(net3759),
    .Y(_02328_));
 sg13g2_nand2_1 _08557_ (.Y(_02329_),
    .A(net3711),
    .B(_02328_));
 sg13g2_nor3_1 _08558_ (.A(net4447),
    .B(net4363),
    .C(net3760),
    .Y(_02330_));
 sg13g2_a22oi_1 _08559_ (.Y(_02331_),
    .B1(_02330_),
    .B2(net3710),
    .A2(net3691),
    .A1(net662));
 sg13g2_inv_1 _08560_ (.Y(_00360_),
    .A(_02331_));
 sg13g2_nand2_1 _08561_ (.Y(_02332_),
    .A(net464),
    .B(net3690));
 sg13g2_o21ai_1 _08562_ (.B1(_02332_),
    .Y(_00361_),
    .A1(net4358),
    .A2(net3690));
 sg13g2_nand2_1 _08563_ (.Y(_02333_),
    .A(net395),
    .B(net3690));
 sg13g2_o21ai_1 _08564_ (.B1(_02333_),
    .Y(_00362_),
    .A1(net4356),
    .A2(net3690));
 sg13g2_nor3_1 _08565_ (.A(net4447),
    .B(net4350),
    .C(net3760),
    .Y(_02334_));
 sg13g2_a22oi_1 _08566_ (.Y(_02335_),
    .B1(_02334_),
    .B2(net3711),
    .A2(net3690),
    .A1(net628));
 sg13g2_inv_1 _08567_ (.Y(_00363_),
    .A(_02335_));
 sg13g2_nor4_2 _08568_ (.A(net4441),
    .B(net4349),
    .C(net3963),
    .Y(_02336_),
    .D(net3760));
 sg13g2_a22oi_1 _08569_ (.Y(_02337_),
    .B1(_02336_),
    .B2(net3762),
    .A2(net3690),
    .A1(net689));
 sg13g2_inv_1 _08570_ (.Y(_00364_),
    .A(net690));
 sg13g2_nor4_2 _08571_ (.A(net4441),
    .B(net4343),
    .C(net3963),
    .Y(_02338_),
    .D(net3760));
 sg13g2_a22oi_1 _08572_ (.Y(_02339_),
    .B1(_02338_),
    .B2(net3762),
    .A2(net3690),
    .A1(net676));
 sg13g2_inv_1 _08573_ (.Y(_00365_),
    .A(_02339_));
 sg13g2_nor3_2 _08574_ (.A(net4342),
    .B(net3962),
    .C(net3759),
    .Y(_02340_));
 sg13g2_a22oi_1 _08575_ (.Y(_02341_),
    .B1(_02340_),
    .B2(net3711),
    .A2(net3690),
    .A1(net658));
 sg13g2_inv_1 _08576_ (.Y(_00366_),
    .A(net659));
 sg13g2_nor4_2 _08577_ (.A(net4442),
    .B(net4337),
    .C(net3963),
    .Y(_02342_),
    .D(net3759));
 sg13g2_a22oi_1 _08578_ (.Y(_02343_),
    .B1(_02342_),
    .B2(net3762),
    .A2(net3691),
    .A1(net774));
 sg13g2_inv_1 _08579_ (.Y(_00367_),
    .A(_02343_));
 sg13g2_nor4_2 _08580_ (.A(net4440),
    .B(net4296),
    .C(net3961),
    .Y(_02344_),
    .D(net3758));
 sg13g2_a22oi_1 _08581_ (.Y(_02345_),
    .B1(_02344_),
    .B2(net3762),
    .A2(net3689),
    .A1(net670));
 sg13g2_inv_1 _08582_ (.Y(_00368_),
    .A(_02345_));
 sg13g2_nor4_2 _08583_ (.A(net4439),
    .B(net4291),
    .C(net3959),
    .Y(_02346_),
    .D(net3756));
 sg13g2_a22oi_1 _08584_ (.Y(_02347_),
    .B1(_02346_),
    .B2(net3761),
    .A2(net3689),
    .A1(net801));
 sg13g2_inv_1 _08585_ (.Y(_00369_),
    .A(_02347_));
 sg13g2_nor4_2 _08586_ (.A(net4439),
    .B(net4288),
    .C(net3959),
    .Y(_02348_),
    .D(net3756));
 sg13g2_a22oi_1 _08587_ (.Y(_02349_),
    .B1(_02348_),
    .B2(net3761),
    .A2(net3689),
    .A1(net758));
 sg13g2_inv_1 _08588_ (.Y(_00370_),
    .A(_02349_));
 sg13g2_nor4_2 _08589_ (.A(net4439),
    .B(net4283),
    .C(net3960),
    .Y(_02350_),
    .D(net3757));
 sg13g2_a22oi_1 _08590_ (.Y(_02351_),
    .B1(_02350_),
    .B2(net3761),
    .A2(net3689),
    .A1(net755));
 sg13g2_inv_1 _08591_ (.Y(_00371_),
    .A(_02351_));
 sg13g2_nor3_2 _08592_ (.A(net4279),
    .B(net3962),
    .C(net3759),
    .Y(_02352_));
 sg13g2_a22oi_1 _08593_ (.Y(_02353_),
    .B1(_02352_),
    .B2(net3711),
    .A2(net3689),
    .A1(net825));
 sg13g2_inv_1 _08594_ (.Y(_00372_),
    .A(_02353_));
 sg13g2_nor4_2 _08595_ (.A(net4439),
    .B(net4276),
    .C(net3960),
    .Y(_02354_),
    .D(net3757));
 sg13g2_a22oi_1 _08596_ (.Y(_02355_),
    .B1(_02354_),
    .B2(net3761),
    .A2(net3689),
    .A1(net775));
 sg13g2_inv_1 _08597_ (.Y(_00373_),
    .A(_02355_));
 sg13g2_nor4_2 _08598_ (.A(net4439),
    .B(net4272),
    .C(net3959),
    .Y(_02356_),
    .D(net3756));
 sg13g2_a22oi_1 _08599_ (.Y(_02357_),
    .B1(_02356_),
    .B2(net3761),
    .A2(net3689),
    .A1(net688));
 sg13g2_inv_1 _08600_ (.Y(_00374_),
    .A(_02357_));
 sg13g2_nor4_2 _08601_ (.A(net4439),
    .B(net4269),
    .C(net3960),
    .Y(_02358_),
    .D(net3757));
 sg13g2_a22oi_1 _08602_ (.Y(_02359_),
    .B1(_02358_),
    .B2(net3761),
    .A2(net3689),
    .A1(net768));
 sg13g2_inv_1 _08603_ (.Y(_00375_),
    .A(_02359_));
 sg13g2_o21ai_1 _08604_ (.B1(_02280_),
    .Y(_02360_),
    .A1(_02255_),
    .A2(net4115));
 sg13g2_nor2_2 _08605_ (.A(net3962),
    .B(_02360_),
    .Y(_02361_));
 sg13g2_nor3_2 _08606_ (.A(net3708),
    .B(net3962),
    .C(_02360_),
    .Y(_02362_));
 sg13g2_nand2b_1 _08607_ (.Y(_02363_),
    .B(net575),
    .A_N(net3688));
 sg13g2_nand2_1 _08608_ (.Y(_02364_),
    .A(_01170_),
    .B(_02361_));
 sg13g2_o21ai_1 _08609_ (.B1(_02363_),
    .Y(_00376_),
    .A1(net3709),
    .A2(_02364_));
 sg13g2_nand2b_1 _08610_ (.Y(_02365_),
    .B(net660),
    .A_N(net3688));
 sg13g2_nand2b_1 _08611_ (.Y(_02366_),
    .B(_02361_),
    .A_N(net4360));
 sg13g2_o21ai_1 _08612_ (.B1(_02365_),
    .Y(_00377_),
    .A1(net3709),
    .A2(_02366_));
 sg13g2_nand2b_1 _08613_ (.Y(_02367_),
    .B(net551),
    .A_N(net3688));
 sg13g2_nand2b_1 _08614_ (.Y(_02368_),
    .B(_02361_),
    .A_N(net4356));
 sg13g2_o21ai_1 _08615_ (.B1(_02367_),
    .Y(_00378_),
    .A1(net3709),
    .A2(_02368_));
 sg13g2_nand2b_1 _08616_ (.Y(_02369_),
    .B(net559),
    .A_N(net3688));
 sg13g2_nand2_1 _08617_ (.Y(_02370_),
    .A(_01171_),
    .B(_02361_));
 sg13g2_o21ai_1 _08618_ (.B1(_02369_),
    .Y(_00379_),
    .A1(net3709),
    .A2(_02370_));
 sg13g2_nor2_1 _08619_ (.A(net644),
    .B(net3687),
    .Y(_02371_));
 sg13g2_a21oi_1 _08620_ (.A1(net4348),
    .A2(net3687),
    .Y(_00380_),
    .B1(_02371_));
 sg13g2_nor2_1 _08621_ (.A(net776),
    .B(net3687),
    .Y(_02372_));
 sg13g2_a21oi_1 _08622_ (.A1(net4343),
    .A2(net3687),
    .Y(_00381_),
    .B1(_02372_));
 sg13g2_nor2_1 _08623_ (.A(net609),
    .B(net3687),
    .Y(_02373_));
 sg13g2_a21oi_1 _08624_ (.A1(net4339),
    .A2(net3687),
    .Y(_00382_),
    .B1(_02373_));
 sg13g2_nor2_1 _08625_ (.A(net737),
    .B(net3687),
    .Y(_02374_));
 sg13g2_a21oi_1 _08626_ (.A1(net4336),
    .A2(net3687),
    .Y(_00383_),
    .B1(_02374_));
 sg13g2_nor2_1 _08627_ (.A(net770),
    .B(net3686),
    .Y(_02375_));
 sg13g2_a21oi_1 _08628_ (.A1(net4294),
    .A2(net3686),
    .Y(_00384_),
    .B1(_02375_));
 sg13g2_nor2_1 _08629_ (.A(net661),
    .B(net3684),
    .Y(_02376_));
 sg13g2_a21oi_1 _08630_ (.A1(net4291),
    .A2(net3684),
    .Y(_00385_),
    .B1(_02376_));
 sg13g2_nor2_1 _08631_ (.A(net742),
    .B(net3684),
    .Y(_02377_));
 sg13g2_a21oi_1 _08632_ (.A1(net4287),
    .A2(net3684),
    .Y(_00386_),
    .B1(_02377_));
 sg13g2_nor2_1 _08633_ (.A(net767),
    .B(net3684),
    .Y(_02378_));
 sg13g2_a21oi_1 _08634_ (.A1(net4281),
    .A2(net3684),
    .Y(_00387_),
    .B1(_02378_));
 sg13g2_nor2_1 _08635_ (.A(net716),
    .B(net3686),
    .Y(_02379_));
 sg13g2_a21oi_1 _08636_ (.A1(net4277),
    .A2(net3686),
    .Y(_00388_),
    .B1(_02379_));
 sg13g2_nor2_1 _08637_ (.A(net735),
    .B(net3685),
    .Y(_02380_));
 sg13g2_a21oi_1 _08638_ (.A1(net4275),
    .A2(net3685),
    .Y(_00389_),
    .B1(_02380_));
 sg13g2_nor2_1 _08639_ (.A(net783),
    .B(net3684),
    .Y(_02381_));
 sg13g2_a21oi_1 _08640_ (.A1(net4273),
    .A2(net3684),
    .Y(_00390_),
    .B1(_02381_));
 sg13g2_nor2_1 _08641_ (.A(net655),
    .B(net3685),
    .Y(_02382_));
 sg13g2_a21oi_1 _08642_ (.A1(net4269),
    .A2(net3685),
    .Y(_00391_),
    .B1(_02382_));
 sg13g2_nand3_1 _08643_ (.B(_02255_),
    .C(_02279_),
    .A(net4443),
    .Y(_02383_));
 sg13g2_nor2_1 _08644_ (.A(net3708),
    .B(_02383_),
    .Y(_02384_));
 sg13g2_nor2_1 _08645_ (.A(\cpu.keccak_alu.registers[64] ),
    .B(net3681),
    .Y(_02385_));
 sg13g2_a21oi_1 _08646_ (.A1(net4364),
    .A2(net3682),
    .Y(_00392_),
    .B1(_02385_));
 sg13g2_nor2_1 _08647_ (.A(net555),
    .B(net3682),
    .Y(_02386_));
 sg13g2_a21oi_1 _08648_ (.A1(net4358),
    .A2(net3681),
    .Y(_00393_),
    .B1(_02386_));
 sg13g2_nor2_1 _08649_ (.A(net610),
    .B(net3681),
    .Y(_02387_));
 sg13g2_a21oi_1 _08650_ (.A1(net4355),
    .A2(net3681),
    .Y(_00394_),
    .B1(_02387_));
 sg13g2_nor2_1 _08651_ (.A(net638),
    .B(net3681),
    .Y(_02388_));
 sg13g2_a21oi_1 _08652_ (.A1(net4350),
    .A2(net3681),
    .Y(_00395_),
    .B1(_02388_));
 sg13g2_nor2_1 _08653_ (.A(net635),
    .B(net3681),
    .Y(_02389_));
 sg13g2_a21oi_1 _08654_ (.A1(net4347),
    .A2(net3681),
    .Y(_00396_),
    .B1(_02389_));
 sg13g2_nor2_1 _08655_ (.A(net543),
    .B(net3682),
    .Y(_02390_));
 sg13g2_a21oi_1 _08656_ (.A1(net4344),
    .A2(net3682),
    .Y(_00397_),
    .B1(_02390_));
 sg13g2_nor2_1 _08657_ (.A(net769),
    .B(net3682),
    .Y(_02391_));
 sg13g2_a21oi_1 _08658_ (.A1(net4340),
    .A2(net3682),
    .Y(_00398_),
    .B1(_02391_));
 sg13g2_nor2_1 _08659_ (.A(net603),
    .B(net3680),
    .Y(_02392_));
 sg13g2_a21oi_1 _08660_ (.A1(net4336),
    .A2(net3680),
    .Y(_00399_),
    .B1(_02392_));
 sg13g2_nor2_1 _08661_ (.A(net226),
    .B(net3683),
    .Y(_02393_));
 sg13g2_a21oi_1 _08662_ (.A1(net4294),
    .A2(net3683),
    .Y(_00400_),
    .B1(_02393_));
 sg13g2_nor2_1 _08663_ (.A(net232),
    .B(net3679),
    .Y(_02394_));
 sg13g2_a21oi_1 _08664_ (.A1(net4290),
    .A2(net3679),
    .Y(_00401_),
    .B1(_02394_));
 sg13g2_nor2_1 _08665_ (.A(net333),
    .B(net3679),
    .Y(_02395_));
 sg13g2_a21oi_1 _08666_ (.A1(net4286),
    .A2(net3679),
    .Y(_00402_),
    .B1(_02395_));
 sg13g2_nor2_1 _08667_ (.A(net503),
    .B(net3680),
    .Y(_02396_));
 sg13g2_a21oi_1 _08668_ (.A1(net4281),
    .A2(net3680),
    .Y(_00403_),
    .B1(_02396_));
 sg13g2_nor2_1 _08669_ (.A(net520),
    .B(net3680),
    .Y(_02397_));
 sg13g2_a21oi_1 _08670_ (.A1(net4278),
    .A2(net3683),
    .Y(_00404_),
    .B1(_02397_));
 sg13g2_nor2_1 _08671_ (.A(net297),
    .B(net3679),
    .Y(_02398_));
 sg13g2_a21oi_1 _08672_ (.A1(net4275),
    .A2(net3679),
    .Y(_00405_),
    .B1(_02398_));
 sg13g2_nor2_1 _08673_ (.A(net262),
    .B(net3679),
    .Y(_02399_));
 sg13g2_a21oi_1 _08674_ (.A1(net4273),
    .A2(net3679),
    .Y(_00406_),
    .B1(_02399_));
 sg13g2_nor2_1 _08675_ (.A(net740),
    .B(net3680),
    .Y(_02400_));
 sg13g2_a21oi_1 _08676_ (.A1(net4270),
    .A2(net3680),
    .Y(_00407_),
    .B1(_02400_));
 sg13g2_nand3_1 _08677_ (.B(net3711),
    .C(net3961),
    .A(net3968),
    .Y(_02401_));
 sg13g2_nand2_1 _08678_ (.Y(_02402_),
    .A(net621),
    .B(net3678));
 sg13g2_o21ai_1 _08679_ (.B1(_02402_),
    .Y(_00408_),
    .A1(net4363),
    .A2(net3678));
 sg13g2_nand2_1 _08680_ (.Y(_02403_),
    .A(net477),
    .B(net3678));
 sg13g2_o21ai_1 _08681_ (.B1(_02403_),
    .Y(_00409_),
    .A1(net4358),
    .A2(net3678));
 sg13g2_nand2_1 _08682_ (.Y(_02404_),
    .A(net421),
    .B(net3677));
 sg13g2_o21ai_1 _08683_ (.B1(_02404_),
    .Y(_00410_),
    .A1(net4355),
    .A2(net3677));
 sg13g2_nor2_1 _08684_ (.A(_01171_),
    .B(net3678),
    .Y(_02405_));
 sg13g2_a21oi_1 _08685_ (.A1(_01018_),
    .A2(net3678),
    .Y(_00411_),
    .B1(_02405_));
 sg13g2_nor2_1 _08686_ (.A(net4156),
    .B(net3677),
    .Y(_02406_));
 sg13g2_a21oi_1 _08687_ (.A1(_01027_),
    .A2(net3677),
    .Y(_00412_),
    .B1(_02406_));
 sg13g2_nand2_1 _08688_ (.Y(_02407_),
    .A(net496),
    .B(net3677));
 sg13g2_o21ai_1 _08689_ (.B1(_02407_),
    .Y(_00413_),
    .A1(net4344),
    .A2(net3677));
 sg13g2_nand2_1 _08690_ (.Y(_02408_),
    .A(net618),
    .B(net3677));
 sg13g2_o21ai_1 _08691_ (.B1(_02408_),
    .Y(_00414_),
    .A1(net4340),
    .A2(net3677));
 sg13g2_nor2_1 _08692_ (.A(_01175_),
    .B(net3676),
    .Y(_02409_));
 sg13g2_a21oi_1 _08693_ (.A1(_01052_),
    .A2(net3676),
    .Y(_00415_),
    .B1(_02409_));
 sg13g2_nand2_1 _08694_ (.Y(_02410_),
    .A(net301),
    .B(net3676));
 sg13g2_o21ai_1 _08695_ (.B1(_02410_),
    .Y(_00416_),
    .A1(net4294),
    .A2(net3676));
 sg13g2_nor2_1 _08696_ (.A(net4154),
    .B(net3674),
    .Y(_02411_));
 sg13g2_a21oi_1 _08697_ (.A1(_01073_),
    .A2(net3674),
    .Y(_00417_),
    .B1(_02411_));
 sg13g2_nor2_1 _08698_ (.A(net4153),
    .B(net3674),
    .Y(_02412_));
 sg13g2_a21oi_1 _08699_ (.A1(_01079_),
    .A2(net3674),
    .Y(_00418_),
    .B1(_02412_));
 sg13g2_nand2_1 _08700_ (.Y(_02413_),
    .A(net257),
    .B(net3675));
 sg13g2_o21ai_1 _08701_ (.B1(_02413_),
    .Y(_00419_),
    .A1(net4281),
    .A2(net3675));
 sg13g2_nand2_1 _08702_ (.Y(_02414_),
    .A(net452),
    .B(net3676));
 sg13g2_o21ai_1 _08703_ (.B1(_02414_),
    .Y(_00420_),
    .A1(net4278),
    .A2(net3676));
 sg13g2_nor2_1 _08704_ (.A(net4152),
    .B(net3674),
    .Y(_02415_));
 sg13g2_a21oi_1 _08705_ (.A1(_01104_),
    .A2(net3674),
    .Y(_00421_),
    .B1(_02415_));
 sg13g2_nor2_1 _08706_ (.A(net4151),
    .B(net3674),
    .Y(_02416_));
 sg13g2_a21oi_1 _08707_ (.A1(_01119_),
    .A2(net3674),
    .Y(_00422_),
    .B1(_02416_));
 sg13g2_nand2_1 _08708_ (.Y(_02417_),
    .A(net304),
    .B(net3675));
 sg13g2_o21ai_1 _08709_ (.B1(_02417_),
    .Y(_00423_),
    .A1(net4270),
    .A2(net3675));
 sg13g2_nand2_2 _08710_ (.Y(_02418_),
    .A(net4446),
    .B(_02326_));
 sg13g2_nor2_1 _08711_ (.A(net3707),
    .B(_02418_),
    .Y(_02419_));
 sg13g2_nor2_1 _08712_ (.A(net754),
    .B(net3672),
    .Y(_02420_));
 sg13g2_a21oi_1 _08713_ (.A1(net4363),
    .A2(net3672),
    .Y(_00424_),
    .B1(_02420_));
 sg13g2_nor2_1 _08714_ (.A(net616),
    .B(net3671),
    .Y(_02421_));
 sg13g2_a21oi_1 _08715_ (.A1(net4360),
    .A2(net3671),
    .Y(_00425_),
    .B1(_02421_));
 sg13g2_nor2_1 _08716_ (.A(net561),
    .B(net3671),
    .Y(_02422_));
 sg13g2_a21oi_1 _08717_ (.A1(net4356),
    .A2(net3671),
    .Y(_00426_),
    .B1(_02422_));
 sg13g2_nor2_1 _08718_ (.A(net696),
    .B(net3671),
    .Y(_02423_));
 sg13g2_a21oi_1 _08719_ (.A1(net4351),
    .A2(net3671),
    .Y(_00427_),
    .B1(_02423_));
 sg13g2_nor2_1 _08720_ (.A(net808),
    .B(net3671),
    .Y(_02424_));
 sg13g2_a21oi_1 _08721_ (.A1(net4347),
    .A2(net3671),
    .Y(_00428_),
    .B1(_02424_));
 sg13g2_o21ai_1 _08722_ (.B1(net862),
    .Y(_02425_),
    .A1(net3709),
    .A2(_02418_));
 sg13g2_nand3_1 _08723_ (.B(net3963),
    .C(_02326_),
    .A(_01173_),
    .Y(_02426_));
 sg13g2_o21ai_1 _08724_ (.B1(_02425_),
    .Y(_00429_),
    .A1(net3709),
    .A2(_02426_));
 sg13g2_nor2_1 _08725_ (.A(net648),
    .B(net3672),
    .Y(_02427_));
 sg13g2_a21oi_1 _08726_ (.A1(net4339),
    .A2(net3672),
    .Y(_00430_),
    .B1(_02427_));
 sg13g2_nor2_1 _08727_ (.A(net590),
    .B(net3673),
    .Y(_02428_));
 sg13g2_a21oi_1 _08728_ (.A1(net4336),
    .A2(net3673),
    .Y(_00431_),
    .B1(_02428_));
 sg13g2_o21ai_1 _08729_ (.B1(net637),
    .Y(_02429_),
    .A1(net3708),
    .A2(_02418_));
 sg13g2_nand3b_1 _08730_ (.B(net3961),
    .C(_02326_),
    .Y(_02430_),
    .A_N(net4296));
 sg13g2_o21ai_1 _08731_ (.B1(_02429_),
    .Y(_00432_),
    .A1(net3708),
    .A2(_02430_));
 sg13g2_nor2_1 _08732_ (.A(net488),
    .B(net3669),
    .Y(_02431_));
 sg13g2_a21oi_1 _08733_ (.A1(net4292),
    .A2(net3669),
    .Y(_00433_),
    .B1(_02431_));
 sg13g2_nor2_1 _08734_ (.A(net549),
    .B(net3669),
    .Y(_02432_));
 sg13g2_a21oi_1 _08735_ (.A1(net4288),
    .A2(net3669),
    .Y(_00434_),
    .B1(_02432_));
 sg13g2_nor2_1 _08736_ (.A(net617),
    .B(net3669),
    .Y(_02433_));
 sg13g2_a21oi_1 _08737_ (.A1(net4281),
    .A2(net3669),
    .Y(_00435_),
    .B1(_02433_));
 sg13g2_nor2_1 _08738_ (.A(net434),
    .B(net3670),
    .Y(_02434_));
 sg13g2_a21oi_1 _08739_ (.A1(net4278),
    .A2(net3670),
    .Y(_00436_),
    .B1(_02434_));
 sg13g2_o21ai_1 _08740_ (.B1(net455),
    .Y(_02435_),
    .A1(net3707),
    .A2(_02418_));
 sg13g2_nand3_1 _08741_ (.B(net3959),
    .C(_02326_),
    .A(net4152),
    .Y(_02436_));
 sg13g2_o21ai_1 _08742_ (.B1(_02435_),
    .Y(_00437_),
    .A1(net3707),
    .A2(_02436_));
 sg13g2_nor2_1 _08743_ (.A(net572),
    .B(net3669),
    .Y(_02437_));
 sg13g2_a21oi_1 _08744_ (.A1(net4272),
    .A2(net3669),
    .Y(_00438_),
    .B1(_02437_));
 sg13g2_nor2_1 _08745_ (.A(net705),
    .B(net3670),
    .Y(_02438_));
 sg13g2_a21oi_1 _08746_ (.A1(net4269),
    .A2(net3670),
    .Y(_00439_),
    .B1(_02438_));
 sg13g2_nand2b_2 _08747_ (.Y(_02439_),
    .B(net3963),
    .A_N(_02360_));
 sg13g2_nor2_2 _08748_ (.A(net3708),
    .B(_02439_),
    .Y(_02440_));
 sg13g2_nor2_1 _08749_ (.A(net700),
    .B(_02440_),
    .Y(_02441_));
 sg13g2_a21oi_1 _08750_ (.A1(net4363),
    .A2(net3610),
    .Y(_00440_),
    .B1(_02441_));
 sg13g2_nor2_1 _08751_ (.A(net715),
    .B(net3610),
    .Y(_02442_));
 sg13g2_a21oi_1 _08752_ (.A1(net4360),
    .A2(net3610),
    .Y(_00441_),
    .B1(_02442_));
 sg13g2_nor2_1 _08753_ (.A(net607),
    .B(net3610),
    .Y(_02443_));
 sg13g2_a21oi_1 _08754_ (.A1(net4356),
    .A2(net3610),
    .Y(_00442_),
    .B1(_02443_));
 sg13g2_nor2_1 _08755_ (.A(net675),
    .B(net3610),
    .Y(_02444_));
 sg13g2_a21oi_1 _08756_ (.A1(net4351),
    .A2(net3610),
    .Y(_00443_),
    .B1(_02444_));
 sg13g2_nor2_1 _08757_ (.A(net728),
    .B(net3610),
    .Y(_02445_));
 sg13g2_a21oi_1 _08758_ (.A1(net4347),
    .A2(net3611),
    .Y(_00444_),
    .B1(_02445_));
 sg13g2_nor2_1 _08759_ (.A(net632),
    .B(net3611),
    .Y(_02446_));
 sg13g2_a21oi_1 _08760_ (.A1(net4343),
    .A2(net3611),
    .Y(_00445_),
    .B1(_02446_));
 sg13g2_nor2_1 _08761_ (.A(net552),
    .B(net3611),
    .Y(_02447_));
 sg13g2_a21oi_1 _08762_ (.A1(net4339),
    .A2(net3611),
    .Y(_00446_),
    .B1(_02447_));
 sg13g2_nor2_1 _08763_ (.A(net654),
    .B(net3611),
    .Y(_02448_));
 sg13g2_a21oi_1 _08764_ (.A1(net4336),
    .A2(net3611),
    .Y(_00447_),
    .B1(_02448_));
 sg13g2_nor2_1 _08765_ (.A(net548),
    .B(net3609),
    .Y(_02449_));
 sg13g2_a21oi_1 _08766_ (.A1(net4294),
    .A2(net3609),
    .Y(_00448_),
    .B1(_02449_));
 sg13g2_nor2_1 _08767_ (.A(net759),
    .B(net3607),
    .Y(_02450_));
 sg13g2_a21oi_1 _08768_ (.A1(net4292),
    .A2(net3607),
    .Y(_00449_),
    .B1(_02450_));
 sg13g2_nor2_1 _08769_ (.A(net799),
    .B(net3607),
    .Y(_02451_));
 sg13g2_a21oi_1 _08770_ (.A1(net4288),
    .A2(net3607),
    .Y(_00450_),
    .B1(_02451_));
 sg13g2_nor2_1 _08771_ (.A(net751),
    .B(net3607),
    .Y(_02452_));
 sg13g2_a21oi_1 _08772_ (.A1(net4281),
    .A2(net3607),
    .Y(_00451_),
    .B1(_02452_));
 sg13g2_nor2_1 _08773_ (.A(net666),
    .B(net3609),
    .Y(_02453_));
 sg13g2_a21oi_1 _08774_ (.A1(net4277),
    .A2(net3609),
    .Y(_00452_),
    .B1(_02453_));
 sg13g2_nor2_1 _08775_ (.A(net567),
    .B(net3608),
    .Y(_02454_));
 sg13g2_a21oi_1 _08776_ (.A1(net4276),
    .A2(net3608),
    .Y(_00453_),
    .B1(_02454_));
 sg13g2_nor2_1 _08777_ (.A(net729),
    .B(net3607),
    .Y(_02455_));
 sg13g2_a21oi_1 _08778_ (.A1(net4272),
    .A2(net3607),
    .Y(_00454_),
    .B1(_02455_));
 sg13g2_nor2_1 _08779_ (.A(net529),
    .B(net3608),
    .Y(_02456_));
 sg13g2_a21oi_1 _08780_ (.A1(net4269),
    .A2(net3608),
    .Y(_00455_),
    .B1(_02456_));
 sg13g2_nand2_2 _08781_ (.Y(_02457_),
    .A(_02256_),
    .B(_02279_));
 sg13g2_or2_1 _08782_ (.X(_02458_),
    .B(net3755),
    .A(net3708));
 sg13g2_nor2_1 _08783_ (.A(net4364),
    .B(_02457_),
    .Y(_02459_));
 sg13g2_a22oi_1 _08784_ (.Y(_02460_),
    .B1(_02459_),
    .B2(net3710),
    .A2(net3668),
    .A1(net4574));
 sg13g2_inv_1 _08785_ (.Y(_00456_),
    .A(_02460_));
 sg13g2_nor2_2 _08786_ (.A(net4359),
    .B(net3755),
    .Y(_02461_));
 sg13g2_a22oi_1 _08787_ (.Y(_02462_),
    .B1(_02461_),
    .B2(net3710),
    .A2(net3668),
    .A1(net4547));
 sg13g2_inv_1 _08788_ (.Y(_00457_),
    .A(_02462_));
 sg13g2_nor2_2 _08789_ (.A(net4355),
    .B(net3755),
    .Y(_02463_));
 sg13g2_a22oi_1 _08790_ (.Y(_02464_),
    .B1(_02463_),
    .B2(net3710),
    .A2(net3668),
    .A1(net4533));
 sg13g2_inv_1 _08791_ (.Y(_00458_),
    .A(_02464_));
 sg13g2_nor2_1 _08792_ (.A(net4350),
    .B(net3755),
    .Y(_02465_));
 sg13g2_a22oi_1 _08793_ (.Y(_02466_),
    .B1(_02465_),
    .B2(net3710),
    .A2(net3668),
    .A1(net4530));
 sg13g2_inv_1 _08794_ (.Y(_00459_),
    .A(_02466_));
 sg13g2_nor2_1 _08795_ (.A(net4347),
    .B(net3755),
    .Y(_02467_));
 sg13g2_a22oi_1 _08796_ (.Y(_02468_),
    .B1(_02467_),
    .B2(net3710),
    .A2(net3668),
    .A1(net4522));
 sg13g2_inv_1 _08797_ (.Y(_00460_),
    .A(_02468_));
 sg13g2_nor2_1 _08798_ (.A(_01173_),
    .B(net3667),
    .Y(_02469_));
 sg13g2_a21oi_1 _08799_ (.A1(net4161),
    .A2(net3667),
    .Y(_00461_),
    .B1(_02469_));
 sg13g2_nor2_2 _08800_ (.A(net4339),
    .B(net3755),
    .Y(_02470_));
 sg13g2_a22oi_1 _08801_ (.Y(_02471_),
    .B1(_02470_),
    .B2(net3710),
    .A2(net3668),
    .A1(net4515));
 sg13g2_inv_1 _08802_ (.Y(_00462_),
    .A(_02471_));
 sg13g2_nor2_1 _08803_ (.A(_01175_),
    .B(net3667),
    .Y(_02472_));
 sg13g2_a21oi_1 _08804_ (.A1(_01055_),
    .A2(net3667),
    .Y(_00463_),
    .B1(_02472_));
 sg13g2_nand2_1 _08805_ (.Y(_02473_),
    .A(net4510),
    .B(net3665));
 sg13g2_o21ai_1 _08806_ (.B1(_02473_),
    .Y(_00464_),
    .A1(net4294),
    .A2(net3665));
 sg13g2_nand2_1 _08807_ (.Y(_02474_),
    .A(net4509),
    .B(net3664));
 sg13g2_o21ai_1 _08808_ (.B1(_02474_),
    .Y(_00465_),
    .A1(net4292),
    .A2(net3664));
 sg13g2_nand2_1 _08809_ (.Y(_02475_),
    .A(net848),
    .B(net3664));
 sg13g2_o21ai_1 _08810_ (.B1(_02475_),
    .Y(_00466_),
    .A1(net4288),
    .A2(net3664));
 sg13g2_nand2_1 _08811_ (.Y(_02476_),
    .A(net861),
    .B(net3664));
 sg13g2_o21ai_1 _08812_ (.B1(_02476_),
    .Y(_00467_),
    .A1(net4282),
    .A2(net3664));
 sg13g2_nand2_1 _08813_ (.Y(_02477_),
    .A(net4507),
    .B(net3665));
 sg13g2_o21ai_1 _08814_ (.B1(_02477_),
    .Y(_00468_),
    .A1(net4279),
    .A2(net3665));
 sg13g2_nand2_1 _08815_ (.Y(_02478_),
    .A(net4506),
    .B(net3666));
 sg13g2_o21ai_1 _08816_ (.B1(_02478_),
    .Y(_00469_),
    .A1(net4276),
    .A2(net3666));
 sg13g2_nand2_1 _08817_ (.Y(_02479_),
    .A(net458),
    .B(net3664));
 sg13g2_o21ai_1 _08818_ (.B1(_02479_),
    .Y(_00470_),
    .A1(net4272),
    .A2(net3664));
 sg13g2_nor2_1 _08819_ (.A(net4270),
    .B(net3755),
    .Y(_02480_));
 sg13g2_a22oi_1 _08820_ (.Y(_02481_),
    .B1(_02480_),
    .B2(net3711),
    .A2(net3666),
    .A1(net4504));
 sg13g2_inv_1 _08821_ (.Y(_00471_),
    .A(_02481_));
 sg13g2_nor2_2 _08822_ (.A(_02287_),
    .B(_02289_),
    .Y(_02482_));
 sg13g2_nor3_2 _08823_ (.A(_02254_),
    .B(_02287_),
    .C(_02289_),
    .Y(_02483_));
 sg13g2_nand2b_1 _08824_ (.Y(_02484_),
    .B(net3754),
    .A_N(_02254_));
 sg13g2_nor2_2 _08825_ (.A(_02285_),
    .B(net3706),
    .Y(_02485_));
 sg13g2_nand2_1 _08826_ (.Y(_02486_),
    .A(_02284_),
    .B(_02483_));
 sg13g2_nor2_1 _08827_ (.A(net4503),
    .B(_02485_),
    .Y(_02487_));
 sg13g2_a21oi_1 _08828_ (.A1(net4365),
    .A2(_02485_),
    .Y(_00472_),
    .B1(_02487_));
 sg13g2_nand2_1 _08829_ (.Y(_02488_),
    .A(net924),
    .B(net3699));
 sg13g2_o21ai_1 _08830_ (.B1(_02488_),
    .Y(_00473_),
    .A1(net4362),
    .A2(net3699));
 sg13g2_nor2_1 _08831_ (.A(net940),
    .B(_02485_),
    .Y(_02489_));
 sg13g2_a21oi_1 _08832_ (.A1(net4354),
    .A2(_02485_),
    .Y(_00474_),
    .B1(_02489_));
 sg13g2_nand2_1 _08833_ (.Y(_02490_),
    .A(\cpu.keccak_alu.registers[147] ),
    .B(net3699));
 sg13g2_o21ai_1 _08834_ (.B1(_02490_),
    .Y(_00475_),
    .A1(net4352),
    .A2(net3699));
 sg13g2_nand2_1 _08835_ (.Y(_02491_),
    .A(net906),
    .B(net3699));
 sg13g2_o21ai_1 _08836_ (.B1(_02491_),
    .Y(_00476_),
    .A1(_02302_),
    .A2(_02484_));
 sg13g2_nand4_1 _08837_ (.B(net3968),
    .C(net3965),
    .A(_01173_),
    .Y(_02492_),
    .D(_02483_));
 sg13g2_o21ai_1 _08838_ (.B1(_02492_),
    .Y(_00477_),
    .A1(_01037_),
    .A2(_02485_));
 sg13g2_nand4_1 _08839_ (.B(net3967),
    .C(net3965),
    .A(net4155),
    .Y(_02493_),
    .D(_02483_));
 sg13g2_o21ai_1 _08840_ (.B1(_02493_),
    .Y(_00478_),
    .A1(_01047_),
    .A2(_02485_));
 sg13g2_nor4_1 _08841_ (.A(net4337),
    .B(net3966),
    .C(net3961),
    .D(net3704),
    .Y(_02494_));
 sg13g2_a21o_1 _08842_ (.A2(net3699),
    .A1(net4502),
    .B1(_02494_),
    .X(_00479_));
 sg13g2_nor4_1 _08843_ (.A(net4296),
    .B(net3966),
    .C(net3960),
    .D(net3703),
    .Y(_02495_));
 sg13g2_a21o_1 _08844_ (.A2(net3699),
    .A1(net4501),
    .B1(_02495_),
    .X(_00480_));
 sg13g2_nand2_1 _08845_ (.Y(_02496_),
    .A(net4500),
    .B(net3700));
 sg13g2_o21ai_1 _08846_ (.B1(_02496_),
    .Y(_00481_),
    .A1(_02312_),
    .A2(net3701));
 sg13g2_nand2_1 _08847_ (.Y(_02497_),
    .A(net882),
    .B(net3700));
 sg13g2_o21ai_1 _08848_ (.B1(_02497_),
    .Y(_00482_),
    .A1(_02314_),
    .A2(net3701));
 sg13g2_nand2_1 _08849_ (.Y(_02498_),
    .A(net4499),
    .B(net3700));
 sg13g2_o21ai_1 _08850_ (.B1(_02498_),
    .Y(_00483_),
    .A1(_02316_),
    .A2(net3701));
 sg13g2_nand2_1 _08851_ (.Y(_02499_),
    .A(net872),
    .B(net3700));
 sg13g2_o21ai_1 _08852_ (.B1(_02499_),
    .Y(_00484_),
    .A1(_02317_),
    .A2(net3704));
 sg13g2_nand2_1 _08853_ (.Y(_02500_),
    .A(net4498),
    .B(net3700));
 sg13g2_o21ai_1 _08854_ (.B1(_02500_),
    .Y(_00485_),
    .A1(_02320_),
    .A2(net3701));
 sg13g2_nand2_1 _08855_ (.Y(_02501_),
    .A(net911),
    .B(net3700));
 sg13g2_o21ai_1 _08856_ (.B1(_02501_),
    .Y(_00486_),
    .A1(_02321_),
    .A2(net3701));
 sg13g2_nand2_1 _08857_ (.Y(_02502_),
    .A(net880),
    .B(net3699));
 sg13g2_o21ai_1 _08858_ (.B1(_02502_),
    .Y(_00487_),
    .A1(_02324_),
    .A2(net3703));
 sg13g2_nor3_2 _08859_ (.A(net4443),
    .B(net3759),
    .C(net3704),
    .Y(_02503_));
 sg13g2_nand2_1 _08860_ (.Y(_02504_),
    .A(_02328_),
    .B(_02483_));
 sg13g2_nand2_1 _08861_ (.Y(_02505_),
    .A(net4497),
    .B(net3663));
 sg13g2_o21ai_1 _08862_ (.B1(_02505_),
    .Y(_00488_),
    .A1(net4365),
    .A2(net3663));
 sg13g2_nor2_1 _08863_ (.A(net4496),
    .B(_02503_),
    .Y(_02506_));
 sg13g2_a21oi_1 _08864_ (.A1(net4362),
    .A2(_02503_),
    .Y(_00489_),
    .B1(_02506_));
 sg13g2_nor2_1 _08865_ (.A(net926),
    .B(_02503_),
    .Y(_02507_));
 sg13g2_a21oi_1 _08866_ (.A1(net4353),
    .A2(_02503_),
    .Y(_00490_),
    .B1(_02507_));
 sg13g2_nand2_1 _08867_ (.Y(_02508_),
    .A(net4495),
    .B(net3663));
 sg13g2_o21ai_1 _08868_ (.B1(_02508_),
    .Y(_00491_),
    .A1(net4352),
    .A2(net3663));
 sg13g2_nor4_1 _08869_ (.A(net4349),
    .B(net3962),
    .C(net3759),
    .D(net3704),
    .Y(_02509_));
 sg13g2_a21o_1 _08870_ (.A2(net3663),
    .A1(net4494),
    .B1(_02509_),
    .X(_00492_));
 sg13g2_nor4_1 _08871_ (.A(net4346),
    .B(net3961),
    .C(net3759),
    .D(net3704),
    .Y(_02510_));
 sg13g2_a21o_1 _08872_ (.A2(net3663),
    .A1(net4493),
    .B1(_02510_),
    .X(_00493_));
 sg13g2_a22oi_1 _08873_ (.Y(_02511_),
    .B1(net3662),
    .B2(net916),
    .A2(_02483_),
    .A1(_02340_));
 sg13g2_inv_1 _08874_ (.Y(_00494_),
    .A(_02511_));
 sg13g2_nand4_1 _08875_ (.B(net3965),
    .C(_02326_),
    .A(_01175_),
    .Y(_02512_),
    .D(_02483_));
 sg13g2_o21ai_1 _08876_ (.B1(_02512_),
    .Y(_00495_),
    .A1(_01056_),
    .A2(_02503_));
 sg13g2_nor4_1 _08877_ (.A(net4296),
    .B(net3961),
    .C(net3758),
    .D(net3703),
    .Y(_02513_));
 sg13g2_a21o_1 _08878_ (.A2(net3662),
    .A1(net900),
    .B1(_02513_),
    .X(_00496_));
 sg13g2_nor4_1 _08879_ (.A(net4291),
    .B(net3959),
    .C(net3756),
    .D(net3702),
    .Y(_02514_));
 sg13g2_a21o_1 _08880_ (.A2(net3662),
    .A1(net920),
    .B1(_02514_),
    .X(_00497_));
 sg13g2_nor4_1 _08881_ (.A(net4288),
    .B(net3959),
    .C(net3756),
    .D(net3702),
    .Y(_02515_));
 sg13g2_a21o_1 _08882_ (.A2(net3662),
    .A1(net4492),
    .B1(_02515_),
    .X(_00498_));
 sg13g2_nor4_1 _08883_ (.A(net4283),
    .B(net3960),
    .C(net3756),
    .D(net3702),
    .Y(_02516_));
 sg13g2_a21o_1 _08884_ (.A2(net3662),
    .A1(net4490),
    .B1(_02516_),
    .X(_00499_));
 sg13g2_a22oi_1 _08885_ (.Y(_02517_),
    .B1(net3663),
    .B2(net247),
    .A2(_02483_),
    .A1(_02352_));
 sg13g2_inv_1 _08886_ (.Y(_00500_),
    .A(_02517_));
 sg13g2_nor4_1 _08887_ (.A(net4276),
    .B(net3959),
    .C(net3756),
    .D(net3702),
    .Y(_02518_));
 sg13g2_a21o_1 _08888_ (.A2(net3662),
    .A1(net4488),
    .B1(_02518_),
    .X(_00501_));
 sg13g2_nor4_1 _08889_ (.A(net4272),
    .B(net3959),
    .C(net3756),
    .D(net3702),
    .Y(_02519_));
 sg13g2_a21o_1 _08890_ (.A2(net3662),
    .A1(net912),
    .B1(_02519_),
    .X(_00502_));
 sg13g2_nor4_1 _08891_ (.A(net4270),
    .B(net3961),
    .C(net3758),
    .D(net3703),
    .Y(_02520_));
 sg13g2_a21o_1 _08892_ (.A2(net3662),
    .A1(net935),
    .B1(_02520_),
    .X(_00503_));
 sg13g2_nor3_2 _08893_ (.A(net3962),
    .B(_02360_),
    .C(net3704),
    .Y(_02521_));
 sg13g2_nand2b_1 _08894_ (.Y(_02522_),
    .B(\cpu.keccak_alu.registers[176] ),
    .A_N(_02521_));
 sg13g2_o21ai_1 _08895_ (.B1(_02522_),
    .Y(_00504_),
    .A1(_02364_),
    .A2(net3706));
 sg13g2_nand2b_1 _08896_ (.Y(_02523_),
    .B(net930),
    .A_N(net3661));
 sg13g2_o21ai_1 _08897_ (.B1(_02523_),
    .Y(_00505_),
    .A1(_02366_),
    .A2(net3706));
 sg13g2_nand2b_1 _08898_ (.Y(_02524_),
    .B(net910),
    .A_N(net3661));
 sg13g2_o21ai_1 _08899_ (.B1(_02524_),
    .Y(_00506_),
    .A1(_02368_),
    .A2(net3706));
 sg13g2_nand2b_1 _08900_ (.Y(_02525_),
    .B(net932),
    .A_N(net3661));
 sg13g2_o21ai_1 _08901_ (.B1(_02525_),
    .Y(_00507_),
    .A1(_02370_),
    .A2(net3706));
 sg13g2_nor2_1 _08902_ (.A(net4487),
    .B(net3660),
    .Y(_02526_));
 sg13g2_a21oi_1 _08903_ (.A1(net4349),
    .A2(net3660),
    .Y(_00508_),
    .B1(_02526_));
 sg13g2_nor2_1 _08904_ (.A(net123),
    .B(net3660),
    .Y(_02527_));
 sg13g2_a21oi_1 _08905_ (.A1(net4346),
    .A2(net3660),
    .Y(_00509_),
    .B1(_02527_));
 sg13g2_nor2_1 _08906_ (.A(net4485),
    .B(_02521_),
    .Y(_02528_));
 sg13g2_a21oi_1 _08907_ (.A1(net4342),
    .A2(_02521_),
    .Y(_00510_),
    .B1(_02528_));
 sg13g2_nor2_1 _08908_ (.A(net837),
    .B(net3661),
    .Y(_02529_));
 sg13g2_a21oi_1 _08909_ (.A1(net4336),
    .A2(net3661),
    .Y(_00511_),
    .B1(_02529_));
 sg13g2_nor2_1 _08910_ (.A(net828),
    .B(net3661),
    .Y(_02530_));
 sg13g2_a21oi_1 _08911_ (.A1(net4294),
    .A2(net3661),
    .Y(_00512_),
    .B1(_02530_));
 sg13g2_nor2_1 _08912_ (.A(net907),
    .B(net3658),
    .Y(_02531_));
 sg13g2_a21oi_1 _08913_ (.A1(net4291),
    .A2(net3658),
    .Y(_00513_),
    .B1(_02531_));
 sg13g2_nor2_1 _08914_ (.A(net915),
    .B(net3658),
    .Y(_02532_));
 sg13g2_a21oi_1 _08915_ (.A1(net4286),
    .A2(net3658),
    .Y(_00514_),
    .B1(_02532_));
 sg13g2_nor2_1 _08916_ (.A(net4484),
    .B(net3658),
    .Y(_02533_));
 sg13g2_a21oi_1 _08917_ (.A1(net4281),
    .A2(net3658),
    .Y(_00515_),
    .B1(_02533_));
 sg13g2_nor2_1 _08918_ (.A(net4483),
    .B(net3660),
    .Y(_02534_));
 sg13g2_a21oi_1 _08919_ (.A1(net4277),
    .A2(net3660),
    .Y(_00516_),
    .B1(_02534_));
 sg13g2_nor2_1 _08920_ (.A(net4482),
    .B(net3659),
    .Y(_02535_));
 sg13g2_a21oi_1 _08921_ (.A1(net4275),
    .A2(net3659),
    .Y(_00517_),
    .B1(_02535_));
 sg13g2_nor2_1 _08922_ (.A(net871),
    .B(net3658),
    .Y(_02536_));
 sg13g2_a21oi_1 _08923_ (.A1(net4272),
    .A2(net3658),
    .Y(_00518_),
    .B1(_02536_));
 sg13g2_nor2_1 _08924_ (.A(net885),
    .B(net3659),
    .Y(_02537_));
 sg13g2_a21oi_1 _08925_ (.A1(net4268),
    .A2(net3659),
    .Y(_00519_),
    .B1(_02537_));
 sg13g2_nor2_2 _08926_ (.A(_02383_),
    .B(net3704),
    .Y(_02538_));
 sg13g2_nor2_1 _08927_ (.A(net412),
    .B(net3657),
    .Y(_02539_));
 sg13g2_a21oi_1 _08928_ (.A1(net4364),
    .A2(net3657),
    .Y(_00520_),
    .B1(_02539_));
 sg13g2_nor2_1 _08929_ (.A(net260),
    .B(net3657),
    .Y(_02540_));
 sg13g2_a21oi_1 _08930_ (.A1(net4358),
    .A2(net3657),
    .Y(_00521_),
    .B1(_02540_));
 sg13g2_nor2_1 _08931_ (.A(net384),
    .B(net3657),
    .Y(_02541_));
 sg13g2_a21oi_1 _08932_ (.A1(net4355),
    .A2(net3657),
    .Y(_00522_),
    .B1(_02541_));
 sg13g2_nor2_1 _08933_ (.A(net443),
    .B(net3656),
    .Y(_02542_));
 sg13g2_a21oi_1 _08934_ (.A1(net4350),
    .A2(net3656),
    .Y(_00523_),
    .B1(_02542_));
 sg13g2_nor2_1 _08935_ (.A(net538),
    .B(net3656),
    .Y(_02543_));
 sg13g2_a21oi_1 _08936_ (.A1(net4347),
    .A2(net3656),
    .Y(_00524_),
    .B1(_02543_));
 sg13g2_nor2_1 _08937_ (.A(net479),
    .B(net3656),
    .Y(_02544_));
 sg13g2_a21oi_1 _08938_ (.A1(net4343),
    .A2(net3656),
    .Y(_00525_),
    .B1(_02544_));
 sg13g2_nor2_1 _08939_ (.A(net426),
    .B(net3656),
    .Y(_02545_));
 sg13g2_a21oi_1 _08940_ (.A1(net4340),
    .A2(net3656),
    .Y(_00526_),
    .B1(_02545_));
 sg13g2_nor2_1 _08941_ (.A(net323),
    .B(net3655),
    .Y(_02546_));
 sg13g2_a21oi_1 _08942_ (.A1(net4337),
    .A2(net3655),
    .Y(_00527_),
    .B1(_02546_));
 sg13g2_nor2_1 _08943_ (.A(net417),
    .B(net3655),
    .Y(_02547_));
 sg13g2_a21oi_1 _08944_ (.A1(net4295),
    .A2(net3655),
    .Y(_00528_),
    .B1(_02547_));
 sg13g2_nor2_1 _08945_ (.A(net573),
    .B(net3653),
    .Y(_02548_));
 sg13g2_a21oi_1 _08946_ (.A1(net4290),
    .A2(net3653),
    .Y(_00529_),
    .B1(_02548_));
 sg13g2_nor2_1 _08947_ (.A(net383),
    .B(net3653),
    .Y(_02549_));
 sg13g2_a21oi_1 _08948_ (.A1(net4286),
    .A2(net3653),
    .Y(_00530_),
    .B1(_02549_));
 sg13g2_nor2_1 _08949_ (.A(net505),
    .B(net3653),
    .Y(_02550_));
 sg13g2_a21oi_1 _08950_ (.A1(net4282),
    .A2(net3653),
    .Y(_00531_),
    .B1(_02550_));
 sg13g2_nor2_1 _08951_ (.A(net478),
    .B(net3655),
    .Y(_02551_));
 sg13g2_a21oi_1 _08952_ (.A1(net4277),
    .A2(net3655),
    .Y(_00532_),
    .B1(_02551_));
 sg13g2_nor2_1 _08953_ (.A(net649),
    .B(net3654),
    .Y(_02552_));
 sg13g2_a21oi_1 _08954_ (.A1(net4275),
    .A2(net3654),
    .Y(_00533_),
    .B1(_02552_));
 sg13g2_nor2_1 _08955_ (.A(net461),
    .B(net3653),
    .Y(_02553_));
 sg13g2_a21oi_1 _08956_ (.A1(net4273),
    .A2(net3653),
    .Y(_00534_),
    .B1(_02553_));
 sg13g2_nor2_1 _08957_ (.A(net540),
    .B(net3654),
    .Y(_02554_));
 sg13g2_a21oi_1 _08958_ (.A1(net4270),
    .A2(net3654),
    .Y(_00535_),
    .B1(_02554_));
 sg13g2_nor3_2 _08959_ (.A(net3966),
    .B(net3964),
    .C(net3703),
    .Y(_02555_));
 sg13g2_nand3_1 _08960_ (.B(net3967),
    .C(_02483_),
    .A(net4443),
    .Y(_02556_));
 sg13g2_nor2_1 _08961_ (.A(net387),
    .B(net3652),
    .Y(_02557_));
 sg13g2_a21oi_1 _08962_ (.A1(net4364),
    .A2(net3652),
    .Y(_00536_),
    .B1(_02557_));
 sg13g2_nor2_1 _08963_ (.A(net424),
    .B(net3652),
    .Y(_02558_));
 sg13g2_a21oi_1 _08964_ (.A1(net4359),
    .A2(net3652),
    .Y(_00537_),
    .B1(_02558_));
 sg13g2_nor2_1 _08965_ (.A(net300),
    .B(net3651),
    .Y(_02559_));
 sg13g2_a21oi_1 _08966_ (.A1(net4356),
    .A2(net3651),
    .Y(_00538_),
    .B1(_02559_));
 sg13g2_nor2_1 _08967_ (.A(net625),
    .B(net3651),
    .Y(_02560_));
 sg13g2_a21oi_1 _08968_ (.A1(net4351),
    .A2(net3651),
    .Y(_00539_),
    .B1(_02560_));
 sg13g2_nor2_1 _08969_ (.A(net415),
    .B(net3651),
    .Y(_02561_));
 sg13g2_a21oi_1 _08970_ (.A1(net4347),
    .A2(net3651),
    .Y(_00540_),
    .B1(_02561_));
 sg13g2_nor4_1 _08971_ (.A(net4346),
    .B(net3966),
    .C(net3965),
    .D(net3704),
    .Y(_02562_));
 sg13g2_a21o_1 _08972_ (.A2(_02556_),
    .A1(net778),
    .B1(_02562_),
    .X(_00541_));
 sg13g2_nor2_1 _08973_ (.A(net502),
    .B(net3651),
    .Y(_02563_));
 sg13g2_a21oi_1 _08974_ (.A1(net4340),
    .A2(net3651),
    .Y(_00542_),
    .B1(_02563_));
 sg13g2_nor2_1 _08975_ (.A(net281),
    .B(net3650),
    .Y(_02564_));
 sg13g2_a21oi_1 _08976_ (.A1(net4337),
    .A2(net3650),
    .Y(_00543_),
    .B1(_02564_));
 sg13g2_nor4_1 _08977_ (.A(net4296),
    .B(net3966),
    .C(net3964),
    .D(net3703),
    .Y(_02565_));
 sg13g2_a21o_1 _08978_ (.A2(_02556_),
    .A1(net773),
    .B1(_02565_),
    .X(_00544_));
 sg13g2_nor2_1 _08979_ (.A(net359),
    .B(net3649),
    .Y(_02566_));
 sg13g2_a21oi_1 _08980_ (.A1(net4290),
    .A2(net3649),
    .Y(_00545_),
    .B1(_02566_));
 sg13g2_nor2_1 _08981_ (.A(net487),
    .B(net3649),
    .Y(_02567_));
 sg13g2_a21oi_1 _08982_ (.A1(net4286),
    .A2(net3649),
    .Y(_00546_),
    .B1(_02567_));
 sg13g2_nor2_1 _08983_ (.A(net560),
    .B(net3650),
    .Y(_02568_));
 sg13g2_a21oi_1 _08984_ (.A1(net4282),
    .A2(net3650),
    .Y(_00547_),
    .B1(_02568_));
 sg13g2_nor2_1 _08985_ (.A(net473),
    .B(net3650),
    .Y(_02569_));
 sg13g2_a21oi_1 _08986_ (.A1(net4279),
    .A2(net3650),
    .Y(_00548_),
    .B1(_02569_));
 sg13g2_nor4_1 _08987_ (.A(net4276),
    .B(net3966),
    .C(net3965),
    .D(net3702),
    .Y(_02570_));
 sg13g2_a21o_1 _08988_ (.A2(_02556_),
    .A1(net615),
    .B1(_02570_),
    .X(_00549_));
 sg13g2_nor2_1 _08989_ (.A(net465),
    .B(net3649),
    .Y(_02571_));
 sg13g2_a21oi_1 _08990_ (.A1(net4273),
    .A2(net3649),
    .Y(_00550_),
    .B1(_02571_));
 sg13g2_nor2_1 _08991_ (.A(net442),
    .B(net3649),
    .Y(_02572_));
 sg13g2_a21oi_1 _08992_ (.A1(net4269),
    .A2(net3649),
    .Y(_00551_),
    .B1(_02572_));
 sg13g2_nor2_2 _08993_ (.A(_02418_),
    .B(net3701),
    .Y(_02573_));
 sg13g2_nor2_1 _08994_ (.A(net420),
    .B(net3648),
    .Y(_02574_));
 sg13g2_a21oi_1 _08995_ (.A1(net4363),
    .A2(net3648),
    .Y(_00552_),
    .B1(_02574_));
 sg13g2_nor2_1 _08996_ (.A(net328),
    .B(net3648),
    .Y(_02575_));
 sg13g2_a21oi_1 _08997_ (.A1(net4358),
    .A2(net3648),
    .Y(_00553_),
    .B1(_02575_));
 sg13g2_nor2_1 _08998_ (.A(net349),
    .B(net3647),
    .Y(_02576_));
 sg13g2_a21oi_1 _08999_ (.A1(net4356),
    .A2(net3647),
    .Y(_00554_),
    .B1(_02576_));
 sg13g2_nor2_1 _09000_ (.A(net414),
    .B(net3647),
    .Y(_02577_));
 sg13g2_a21oi_1 _09001_ (.A1(net4350),
    .A2(net3647),
    .Y(_00555_),
    .B1(_02577_));
 sg13g2_nor2_1 _09002_ (.A(net674),
    .B(net3647),
    .Y(_02578_));
 sg13g2_a21oi_1 _09003_ (.A1(net4348),
    .A2(net3647),
    .Y(_00556_),
    .B1(_02578_));
 sg13g2_o21ai_1 _09004_ (.B1(net273),
    .Y(_02579_),
    .A1(_02418_),
    .A2(net3706));
 sg13g2_o21ai_1 _09005_ (.B1(_02579_),
    .Y(_00557_),
    .A1(_02426_),
    .A2(net3706));
 sg13g2_nor2_1 _09006_ (.A(net375),
    .B(net3647),
    .Y(_02580_));
 sg13g2_a21oi_1 _09007_ (.A1(net4339),
    .A2(net3647),
    .Y(_00558_),
    .B1(_02580_));
 sg13g2_nor2_1 _09008_ (.A(net494),
    .B(net3646),
    .Y(_02581_));
 sg13g2_a21oi_1 _09009_ (.A1(net4336),
    .A2(net3646),
    .Y(_00559_),
    .B1(_02581_));
 sg13g2_o21ai_1 _09010_ (.B1(net539),
    .Y(_02582_),
    .A1(_02418_),
    .A2(net3703));
 sg13g2_o21ai_1 _09011_ (.B1(_02582_),
    .Y(_00560_),
    .A1(_02430_),
    .A2(net3703));
 sg13g2_nor2_1 _09012_ (.A(net547),
    .B(net3645),
    .Y(_02583_));
 sg13g2_a21oi_1 _09013_ (.A1(net4290),
    .A2(net3645),
    .Y(_00561_),
    .B1(_02583_));
 sg13g2_nor2_1 _09014_ (.A(net449),
    .B(net3645),
    .Y(_02584_));
 sg13g2_a21oi_1 _09015_ (.A1(net4287),
    .A2(net3645),
    .Y(_00562_),
    .B1(_02584_));
 sg13g2_nor2_1 _09016_ (.A(net683),
    .B(net3645),
    .Y(_02585_));
 sg13g2_a21oi_1 _09017_ (.A1(net4281),
    .A2(net3645),
    .Y(_00563_),
    .B1(_02585_));
 sg13g2_nor2_1 _09018_ (.A(net459),
    .B(net3646),
    .Y(_02586_));
 sg13g2_a21oi_1 _09019_ (.A1(net4277),
    .A2(net3646),
    .Y(_00564_),
    .B1(_02586_));
 sg13g2_o21ai_1 _09020_ (.B1(net401),
    .Y(_02587_),
    .A1(_02418_),
    .A2(net3701));
 sg13g2_o21ai_1 _09021_ (.B1(_02587_),
    .Y(_00565_),
    .A1(_02436_),
    .A2(net3701));
 sg13g2_nor2_1 _09022_ (.A(\cpu.keccak_alu.registers[238] ),
    .B(net3645),
    .Y(_02588_));
 sg13g2_a21oi_1 _09023_ (.A1(net4274),
    .A2(net3645),
    .Y(_00566_),
    .B1(_02588_));
 sg13g2_nor2_1 _09024_ (.A(net316),
    .B(net3646),
    .Y(_02589_));
 sg13g2_a21oi_1 _09025_ (.A1(net4269),
    .A2(net3646),
    .Y(_00567_),
    .B1(_02589_));
 sg13g2_nor4_2 _09026_ (.A(_02254_),
    .B(_02287_),
    .C(_02289_),
    .Y(_02590_),
    .D(_02439_));
 sg13g2_nor2_1 _09027_ (.A(net510),
    .B(net3605),
    .Y(_02591_));
 sg13g2_a21oi_1 _09028_ (.A1(net4363),
    .A2(net3605),
    .Y(_00568_),
    .B1(_02591_));
 sg13g2_nor2_1 _09029_ (.A(net597),
    .B(net3606),
    .Y(_02592_));
 sg13g2_a21oi_1 _09030_ (.A1(net4361),
    .A2(net3606),
    .Y(_00569_),
    .B1(_02592_));
 sg13g2_nor2_1 _09031_ (.A(net748),
    .B(net3605),
    .Y(_02593_));
 sg13g2_a21oi_1 _09032_ (.A1(net4356),
    .A2(net3605),
    .Y(_00570_),
    .B1(_02593_));
 sg13g2_nor2_1 _09033_ (.A(net532),
    .B(net3605),
    .Y(_02594_));
 sg13g2_a21oi_1 _09034_ (.A1(net4350),
    .A2(net3605),
    .Y(_00571_),
    .B1(_02594_));
 sg13g2_nor2_1 _09035_ (.A(net693),
    .B(net3605),
    .Y(_02595_));
 sg13g2_a21oi_1 _09036_ (.A1(net4347),
    .A2(net3605),
    .Y(_00572_),
    .B1(_02595_));
 sg13g2_nor2_1 _09037_ (.A(net504),
    .B(net3606),
    .Y(_02596_));
 sg13g2_a21oi_1 _09038_ (.A1(net4343),
    .A2(net3604),
    .Y(_00573_),
    .B1(_02596_));
 sg13g2_nor2_1 _09039_ (.A(net563),
    .B(net3606),
    .Y(_02597_));
 sg13g2_a21oi_1 _09040_ (.A1(net4339),
    .A2(net3606),
    .Y(_00574_),
    .B1(_02597_));
 sg13g2_nor2_1 _09041_ (.A(net358),
    .B(net3604),
    .Y(_02598_));
 sg13g2_a21oi_1 _09042_ (.A1(net4336),
    .A2(net3604),
    .Y(_00575_),
    .B1(_02598_));
 sg13g2_nor2_1 _09043_ (.A(net587),
    .B(net3604),
    .Y(_02599_));
 sg13g2_a21oi_1 _09044_ (.A1(net4294),
    .A2(net3602),
    .Y(_00576_),
    .B1(_02599_));
 sg13g2_nor2_1 _09045_ (.A(net490),
    .B(net3602),
    .Y(_02600_));
 sg13g2_a21oi_1 _09046_ (.A1(net4290),
    .A2(net3602),
    .Y(_00577_),
    .B1(_02600_));
 sg13g2_nor2_1 _09047_ (.A(net430),
    .B(net3602),
    .Y(_02601_));
 sg13g2_a21oi_1 _09048_ (.A1(net4286),
    .A2(net3602),
    .Y(_00578_),
    .B1(_02601_));
 sg13g2_nor2_1 _09049_ (.A(net614),
    .B(net3603),
    .Y(_02602_));
 sg13g2_a21oi_1 _09050_ (.A1(net4281),
    .A2(net3602),
    .Y(_00579_),
    .B1(_02602_));
 sg13g2_nor2_1 _09051_ (.A(net411),
    .B(net3604),
    .Y(_02603_));
 sg13g2_a21oi_1 _09052_ (.A1(net4277),
    .A2(net3604),
    .Y(_00580_),
    .B1(_02603_));
 sg13g2_nor2_1 _09053_ (.A(net404),
    .B(net3603),
    .Y(_02604_));
 sg13g2_a21oi_1 _09054_ (.A1(net4275),
    .A2(net3603),
    .Y(_00581_),
    .B1(_02604_));
 sg13g2_nor2_1 _09055_ (.A(net533),
    .B(net3602),
    .Y(_02605_));
 sg13g2_a21oi_1 _09056_ (.A1(net4272),
    .A2(net3602),
    .Y(_00582_),
    .B1(_02605_));
 sg13g2_nor2_1 _09057_ (.A(net435),
    .B(net3603),
    .Y(_02606_));
 sg13g2_a21oi_1 _09058_ (.A1(net4268),
    .A2(net3603),
    .Y(_00583_),
    .B1(_02606_));
 sg13g2_nor3_2 _09059_ (.A(net4430),
    .B(net4432),
    .C(_00044_),
    .Y(_02607_));
 sg13g2_and2_1 _09060_ (.A(\cpu.registers[4][0] ),
    .B(net4096),
    .X(_02608_));
 sg13g2_nand2b_1 _09061_ (.Y(_02609_),
    .B(net4430),
    .A_N(net4432));
 sg13g2_nor2_1 _09062_ (.A(net4418),
    .B(_02609_),
    .Y(_02610_));
 sg13g2_nand2b_1 _09063_ (.Y(_02611_),
    .B(net4432),
    .A_N(net4430));
 sg13g2_nor2_1 _09064_ (.A(net4418),
    .B(_02611_),
    .Y(_02612_));
 sg13g2_a221oi_1 _09065_ (.B2(\cpu.registers[1][0] ),
    .C1(_02608_),
    .B1(net3956),
    .A1(\cpu.registers[2][0] ),
    .Y(_02613_),
    .A2(net3958));
 sg13g2_nor2_1 _09066_ (.A(net4418),
    .B(_02278_),
    .Y(_02614_));
 sg13g2_nor2_1 _09067_ (.A(_00044_),
    .B(_02611_),
    .Y(_02615_));
 sg13g2_a22oi_1 _09068_ (.Y(_02616_),
    .B1(net3952),
    .B2(\cpu.registers[5][0] ),
    .A2(net3954),
    .A1(\cpu.registers[3][0] ));
 sg13g2_nor2_1 _09069_ (.A(_00044_),
    .B(_02609_),
    .Y(_02617_));
 sg13g2_or2_1 _09070_ (.X(_02618_),
    .B(_02278_),
    .A(_00044_));
 sg13g2_inv_4 _09071_ (.A(net3948),
    .Y(_02619_));
 sg13g2_a22oi_1 _09072_ (.Y(_02620_),
    .B1(_02619_),
    .B2(\cpu.registers[7][0] ),
    .A2(net3950),
    .A1(\cpu.registers[6][0] ));
 sg13g2_nand3_1 _09073_ (.B(_02616_),
    .C(_02620_),
    .A(_02613_),
    .Y(_02621_));
 sg13g2_nor2_1 _09074_ (.A(_01233_),
    .B(net4051),
    .Y(_02622_));
 sg13g2_nand2b_1 _09075_ (.Y(_02623_),
    .B(net3864),
    .A_N(_01233_));
 sg13g2_nor2_1 _09076_ (.A(_01258_),
    .B(net3798),
    .Y(_02624_));
 sg13g2_nand3_1 _09077_ (.B(net4078),
    .C(net3864),
    .A(net4306),
    .Y(_02625_));
 sg13g2_nand2b_1 _09078_ (.Y(_02626_),
    .B(net4307),
    .A_N(\cpu.execution_stage[0] ));
 sg13g2_nand2_1 _09079_ (.Y(_02627_),
    .A(net4143),
    .B(_02626_));
 sg13g2_o21ai_1 _09080_ (.B1(_02627_),
    .Y(_02628_),
    .A1(_01273_),
    .A2(_02625_));
 sg13g2_inv_1 _09081_ (.Y(_02629_),
    .A(net3748));
 sg13g2_nor2_1 _09082_ (.A(_00018_),
    .B(net4074),
    .Y(_02630_));
 sg13g2_o21ai_1 _09083_ (.B1(_02630_),
    .Y(_02631_),
    .A1(_00043_),
    .A2(net4037));
 sg13g2_a221oi_1 _09084_ (.B2(net3753),
    .C1(_02631_),
    .B1(_02621_),
    .A1(net4450),
    .Y(_02632_),
    .A2(_01244_));
 sg13g2_nor2_1 _09085_ (.A(net4474),
    .B(_02629_),
    .Y(_02633_));
 sg13g2_a21oi_1 _09086_ (.A1(_02629_),
    .A2(_02632_),
    .Y(_00584_),
    .B1(_02633_));
 sg13g2_nor2_1 _09087_ (.A(_00031_),
    .B(net3948),
    .Y(_02634_));
 sg13g2_a221oi_1 _09088_ (.B2(\cpu.registers[2][1] ),
    .C1(_02634_),
    .B1(net3958),
    .A1(\cpu.registers[4][1] ),
    .Y(_02635_),
    .A2(net4096));
 sg13g2_a22oi_1 _09089_ (.Y(_02636_),
    .B1(net3950),
    .B2(\cpu.registers[6][1] ),
    .A2(net3956),
    .A1(\cpu.registers[1][1] ));
 sg13g2_a22oi_1 _09090_ (.Y(_02637_),
    .B1(net3952),
    .B2(\cpu.registers[5][1] ),
    .A2(net3954),
    .A1(\cpu.registers[3][1] ));
 sg13g2_nand3_1 _09091_ (.B(_02636_),
    .C(_02637_),
    .A(_02635_),
    .Y(_02638_));
 sg13g2_nand2_2 _09092_ (.Y(_02639_),
    .A(net4306),
    .B(_02629_));
 sg13g2_nor3_2 _09093_ (.A(net4038),
    .B(net3797),
    .C(_02639_),
    .Y(_02640_));
 sg13g2_nand3_1 _09094_ (.B(net3753),
    .C(_02629_),
    .A(net4306),
    .Y(_02641_));
 sg13g2_nand2_1 _09095_ (.Y(_02642_),
    .A(net4472),
    .B(_02628_));
 sg13g2_nor2_1 _09096_ (.A(_00030_),
    .B(net4036),
    .Y(_02643_));
 sg13g2_a221oi_1 _09097_ (.B2(_02638_),
    .C1(_02643_),
    .B1(net3752),
    .A1(net4240),
    .Y(_02644_),
    .A2(_01244_));
 sg13g2_o21ai_1 _09098_ (.B1(_02642_),
    .Y(_00585_),
    .A1(_02639_),
    .A2(_02644_));
 sg13g2_nor2_1 _09099_ (.A(_00032_),
    .B(net3948),
    .Y(_02645_));
 sg13g2_a221oi_1 _09100_ (.B2(\cpu.registers[5][2] ),
    .C1(_02645_),
    .B1(net3952),
    .A1(\cpu.registers[1][2] ),
    .Y(_02646_),
    .A2(net3956));
 sg13g2_a22oi_1 _09101_ (.Y(_02647_),
    .B1(net3954),
    .B2(\cpu.registers[3][2] ),
    .A2(net4096),
    .A1(\cpu.registers[4][2] ));
 sg13g2_a22oi_1 _09102_ (.Y(_02648_),
    .B1(net3950),
    .B2(\cpu.registers[6][2] ),
    .A2(net3958),
    .A1(\cpu.registers[2][2] ));
 sg13g2_nand3_1 _09103_ (.B(_02647_),
    .C(_02648_),
    .A(_02646_),
    .Y(_02649_));
 sg13g2_nand2_1 _09104_ (.Y(_02650_),
    .A(net4470),
    .B(net3749));
 sg13g2_a22oi_1 _09105_ (.Y(_02651_),
    .B1(net3752),
    .B2(_02649_),
    .A2(net4039),
    .A1(net4433));
 sg13g2_o21ai_1 _09106_ (.B1(_02650_),
    .Y(_00586_),
    .A1(_02639_),
    .A2(_02651_));
 sg13g2_nand2_1 _09107_ (.Y(_02652_),
    .A(\cpu.registers[2][3] ),
    .B(net3958));
 sg13g2_a22oi_1 _09108_ (.Y(_02653_),
    .B1(net3952),
    .B2(\cpu.registers[5][3] ),
    .A2(net3956),
    .A1(\cpu.registers[1][3] ));
 sg13g2_a22oi_1 _09109_ (.Y(_02654_),
    .B1(_02619_),
    .B2(_00921_),
    .A2(net4096),
    .A1(\cpu.registers[4][3] ));
 sg13g2_a22oi_1 _09110_ (.Y(_02655_),
    .B1(net3950),
    .B2(\cpu.registers[6][3] ),
    .A2(net3954),
    .A1(\cpu.registers[3][3] ));
 sg13g2_nand4_1 _09111_ (.B(_02653_),
    .C(_02654_),
    .A(_02652_),
    .Y(_02656_),
    .D(_02655_));
 sg13g2_nand2_1 _09112_ (.Y(_02657_),
    .A(net4469),
    .B(net3749));
 sg13g2_a22oi_1 _09113_ (.Y(_02658_),
    .B1(net3751),
    .B2(_02656_),
    .A2(net4039),
    .A1(net194));
 sg13g2_o21ai_1 _09114_ (.B1(_02657_),
    .Y(_00587_),
    .A1(_02639_),
    .A2(_02658_));
 sg13g2_nand2_1 _09115_ (.Y(_02659_),
    .A(\cpu.registers[5][4] ),
    .B(net3952));
 sg13g2_a22oi_1 _09116_ (.Y(_02660_),
    .B1(net3950),
    .B2(\cpu.registers[6][4] ),
    .A2(net3954),
    .A1(\cpu.registers[3][4] ));
 sg13g2_a22oi_1 _09117_ (.Y(_02661_),
    .B1(_02619_),
    .B2(_00928_),
    .A2(net3956),
    .A1(\cpu.registers[1][4] ));
 sg13g2_a22oi_1 _09118_ (.Y(_02662_),
    .B1(net3958),
    .B2(\cpu.registers[2][4] ),
    .A2(net4096),
    .A1(\cpu.registers[4][4] ));
 sg13g2_nand4_1 _09119_ (.B(_02660_),
    .C(_02661_),
    .A(_02659_),
    .Y(_02663_),
    .D(_02662_));
 sg13g2_a22oi_1 _09120_ (.Y(_02664_),
    .B1(net3752),
    .B2(_02663_),
    .A2(net4039),
    .A1(net4422));
 sg13g2_nand2_1 _09121_ (.Y(_02665_),
    .A(net4468),
    .B(net3749));
 sg13g2_o21ai_1 _09122_ (.B1(_02665_),
    .Y(_00588_),
    .A1(_02639_),
    .A2(_02664_));
 sg13g2_nor2_1 _09123_ (.A(_00035_),
    .B(net3948),
    .Y(_02666_));
 sg13g2_a221oi_1 _09124_ (.B2(\cpu.registers[1][5] ),
    .C1(_02666_),
    .B1(net3956),
    .A1(\cpu.registers[4][5] ),
    .Y(_02667_),
    .A2(net4096));
 sg13g2_a22oi_1 _09125_ (.Y(_02668_),
    .B1(net3950),
    .B2(\cpu.registers[6][5] ),
    .A2(net3952),
    .A1(\cpu.registers[5][5] ));
 sg13g2_a22oi_1 _09126_ (.Y(_02669_),
    .B1(net3954),
    .B2(\cpu.registers[3][5] ),
    .A2(net3958),
    .A1(\cpu.registers[2][5] ));
 sg13g2_nand3_1 _09127_ (.B(_02668_),
    .C(_02669_),
    .A(_02667_),
    .Y(_02670_));
 sg13g2_a22oi_1 _09128_ (.Y(_02671_),
    .B1(net3751),
    .B2(_02670_),
    .A2(net4039),
    .A1(net4402));
 sg13g2_nand2_1 _09129_ (.Y(_02672_),
    .A(net4467),
    .B(net3749));
 sg13g2_o21ai_1 _09130_ (.B1(_02672_),
    .Y(_00589_),
    .A1(_02639_),
    .A2(_02671_));
 sg13g2_nand2_1 _09131_ (.Y(_02673_),
    .A(net901),
    .B(net3749));
 sg13g2_nor2_1 _09132_ (.A(_00036_),
    .B(net3947),
    .Y(_02674_));
 sg13g2_a221oi_1 _09133_ (.B2(\cpu.registers[6][6] ),
    .C1(_02674_),
    .B1(net3950),
    .A1(\cpu.registers[3][6] ),
    .Y(_02675_),
    .A2(net3954));
 sg13g2_a22oi_1 _09134_ (.Y(_02676_),
    .B1(net3952),
    .B2(\cpu.registers[5][6] ),
    .A2(net4096),
    .A1(\cpu.registers[4][6] ));
 sg13g2_a22oi_1 _09135_ (.Y(_02677_),
    .B1(net3956),
    .B2(\cpu.registers[1][6] ),
    .A2(net3958),
    .A1(\cpu.registers[2][6] ));
 sg13g2_nand3_1 _09136_ (.B(_02676_),
    .C(_02677_),
    .A(_02675_),
    .Y(_02678_));
 sg13g2_a22oi_1 _09137_ (.Y(_02679_),
    .B1(net3752),
    .B2(_02678_),
    .A2(net4039),
    .A1(net4382));
 sg13g2_o21ai_1 _09138_ (.B1(_02673_),
    .Y(_00590_),
    .A1(_02639_),
    .A2(_02679_));
 sg13g2_nand2_1 _09139_ (.Y(_02680_),
    .A(net811),
    .B(net3749));
 sg13g2_nand2_1 _09140_ (.Y(_02681_),
    .A(\cpu.registers[6][7] ),
    .B(net3950));
 sg13g2_a22oi_1 _09141_ (.Y(_02682_),
    .B1(net3954),
    .B2(\cpu.registers[3][7] ),
    .A2(net3956),
    .A1(\cpu.registers[1][7] ));
 sg13g2_a22oi_1 _09142_ (.Y(_02683_),
    .B1(_02619_),
    .B2(_00950_),
    .A2(net3958),
    .A1(\cpu.registers[2][7] ));
 sg13g2_a22oi_1 _09143_ (.Y(_02684_),
    .B1(net3952),
    .B2(\cpu.registers[5][7] ),
    .A2(net4096),
    .A1(\cpu.registers[4][7] ));
 sg13g2_nand4_1 _09144_ (.B(_02682_),
    .C(_02683_),
    .A(_02681_),
    .Y(_02685_),
    .D(_02684_));
 sg13g2_a22oi_1 _09145_ (.Y(_02686_),
    .B1(net3752),
    .B2(_02685_),
    .A2(net4039),
    .A1(\cpu.current_instruction[15] ));
 sg13g2_o21ai_1 _09146_ (.B1(_02680_),
    .Y(_00591_),
    .A1(_02639_),
    .A2(_02686_));
 sg13g2_nand2_1 _09147_ (.Y(_02687_),
    .A(\cpu.registers[1][8] ),
    .B(net3955));
 sg13g2_nand2_1 _09148_ (.Y(_02688_),
    .A(\cpu.registers[5][8] ),
    .B(net3951));
 sg13g2_a22oi_1 _09149_ (.Y(_02689_),
    .B1(net3953),
    .B2(\cpu.registers[3][8] ),
    .A2(net4095),
    .A1(\cpu.registers[4][8] ));
 sg13g2_o21ai_1 _09150_ (.B1(_02687_),
    .Y(_02690_),
    .A1(_00038_),
    .A2(net3947));
 sg13g2_a221oi_1 _09151_ (.B2(\cpu.registers[6][8] ),
    .C1(_02690_),
    .B1(net3949),
    .A1(\cpu.registers[2][8] ),
    .Y(_02691_),
    .A2(net3957));
 sg13g2_nand3_1 _09152_ (.B(_02689_),
    .C(_02691_),
    .A(_02688_),
    .Y(_02692_));
 sg13g2_a22oi_1 _09153_ (.Y(_02693_),
    .B1(_02640_),
    .B2(_02692_),
    .A2(net3748),
    .A1(net788));
 sg13g2_inv_1 _09154_ (.Y(_00592_),
    .A(_02693_));
 sg13g2_nor2_1 _09155_ (.A(_00039_),
    .B(net3947),
    .Y(_02694_));
 sg13g2_a221oi_1 _09156_ (.B2(\cpu.registers[1][9] ),
    .C1(_02694_),
    .B1(net3955),
    .A1(\cpu.registers[2][9] ),
    .Y(_02695_),
    .A2(net3957));
 sg13g2_a22oi_1 _09157_ (.Y(_02696_),
    .B1(net3951),
    .B2(\cpu.registers[5][9] ),
    .A2(net4095),
    .A1(\cpu.registers[4][9] ));
 sg13g2_a22oi_1 _09158_ (.Y(_02697_),
    .B1(net3949),
    .B2(\cpu.registers[6][9] ),
    .A2(net3953),
    .A1(\cpu.registers[3][9] ));
 sg13g2_nand3_1 _09159_ (.B(_02696_),
    .C(_02697_),
    .A(_02695_),
    .Y(_02698_));
 sg13g2_a22oi_1 _09160_ (.Y(_02699_),
    .B1(_02640_),
    .B2(_02698_),
    .A2(net3749),
    .A1(net756));
 sg13g2_inv_1 _09161_ (.Y(_00593_),
    .A(_02699_));
 sg13g2_nor2_1 _09162_ (.A(_00040_),
    .B(net3947),
    .Y(_02700_));
 sg13g2_a221oi_1 _09163_ (.B2(\cpu.registers[5][10] ),
    .C1(_02700_),
    .B1(net3951),
    .A1(\cpu.registers[4][10] ),
    .Y(_02701_),
    .A2(net4095));
 sg13g2_a22oi_1 _09164_ (.Y(_02702_),
    .B1(net3953),
    .B2(\cpu.registers[3][10] ),
    .A2(net3955),
    .A1(\cpu.registers[1][10] ));
 sg13g2_a22oi_1 _09165_ (.Y(_02703_),
    .B1(net3949),
    .B2(\cpu.registers[6][10] ),
    .A2(net3957),
    .A1(\cpu.registers[2][10] ));
 sg13g2_nand3_1 _09166_ (.B(_02702_),
    .C(_02703_),
    .A(_02701_),
    .Y(_02704_));
 sg13g2_a22oi_1 _09167_ (.Y(_02705_),
    .B1(_02640_),
    .B2(_02704_),
    .A2(net3748),
    .A1(net605));
 sg13g2_inv_1 _09168_ (.Y(_00594_),
    .A(_02705_));
 sg13g2_nand2_1 _09169_ (.Y(_02706_),
    .A(net565),
    .B(net3748));
 sg13g2_a22oi_1 _09170_ (.Y(_02707_),
    .B1(net3953),
    .B2(\cpu.registers[3][11] ),
    .A2(net3957),
    .A1(\cpu.registers[2][11] ));
 sg13g2_o21ai_1 _09171_ (.B1(_02707_),
    .Y(_02708_),
    .A1(_00041_),
    .A2(net3947));
 sg13g2_a22oi_1 _09172_ (.Y(_02709_),
    .B1(net3951),
    .B2(\cpu.registers[5][11] ),
    .A2(net3955),
    .A1(\cpu.registers[1][11] ));
 sg13g2_a22oi_1 _09173_ (.Y(_02710_),
    .B1(net3949),
    .B2(\cpu.registers[6][11] ),
    .A2(net4095),
    .A1(\cpu.registers[4][11] ));
 sg13g2_nand2_1 _09174_ (.Y(_02711_),
    .A(_02709_),
    .B(_02710_));
 sg13g2_nor2_2 _09175_ (.A(_02708_),
    .B(_02711_),
    .Y(_02712_));
 sg13g2_inv_1 _09176_ (.Y(_02713_),
    .A(_02712_));
 sg13g2_o21ai_1 _09177_ (.B1(_02706_),
    .Y(_00595_),
    .A1(_02641_),
    .A2(_02712_));
 sg13g2_a22oi_1 _09178_ (.Y(_02714_),
    .B1(net3949),
    .B2(\cpu.registers[6][12] ),
    .A2(net4095),
    .A1(\cpu.registers[4][12] ));
 sg13g2_nand2_1 _09179_ (.Y(_02715_),
    .A(\cpu.registers[1][12] ),
    .B(net3955));
 sg13g2_a22oi_1 _09180_ (.Y(_02716_),
    .B1(net3953),
    .B2(\cpu.registers[3][12] ),
    .A2(net3957),
    .A1(\cpu.registers[2][12] ));
 sg13g2_a22oi_1 _09181_ (.Y(_02717_),
    .B1(_02619_),
    .B2(_00989_),
    .A2(net3951),
    .A1(\cpu.registers[5][12] ));
 sg13g2_nand4_1 _09182_ (.B(_02715_),
    .C(_02716_),
    .A(_02714_),
    .Y(_02718_),
    .D(_02717_));
 sg13g2_a22oi_1 _09183_ (.Y(_02719_),
    .B1(_02640_),
    .B2(_02718_),
    .A2(net3748),
    .A1(net429));
 sg13g2_inv_1 _09184_ (.Y(_00596_),
    .A(_02719_));
 sg13g2_nor2_1 _09185_ (.A(_00046_),
    .B(net3947),
    .Y(_02720_));
 sg13g2_a221oi_1 _09186_ (.B2(\cpu.registers[5][13] ),
    .C1(_02720_),
    .B1(net3951),
    .A1(\cpu.registers[4][13] ),
    .Y(_02721_),
    .A2(net4095));
 sg13g2_a22oi_1 _09187_ (.Y(_02722_),
    .B1(net3949),
    .B2(\cpu.registers[6][13] ),
    .A2(net3957),
    .A1(\cpu.registers[2][13] ));
 sg13g2_a22oi_1 _09188_ (.Y(_02723_),
    .B1(net3953),
    .B2(\cpu.registers[3][13] ),
    .A2(net3955),
    .A1(\cpu.registers[1][13] ));
 sg13g2_nand3_1 _09189_ (.B(_02722_),
    .C(_02723_),
    .A(_02721_),
    .Y(_02724_));
 sg13g2_a22oi_1 _09190_ (.Y(_02725_),
    .B1(_02640_),
    .B2(_02724_),
    .A2(net3748),
    .A1(net634));
 sg13g2_inv_1 _09191_ (.Y(_00597_),
    .A(_02725_));
 sg13g2_nand2_1 _09192_ (.Y(_02726_),
    .A(net135),
    .B(net3748));
 sg13g2_nor2_1 _09193_ (.A(_00047_),
    .B(net3947),
    .Y(_02727_));
 sg13g2_a221oi_1 _09194_ (.B2(\cpu.registers[1][14] ),
    .C1(_02727_),
    .B1(net3955),
    .A1(\cpu.registers[4][14] ),
    .Y(_02728_),
    .A2(net4095));
 sg13g2_a22oi_1 _09195_ (.Y(_02729_),
    .B1(net3949),
    .B2(\cpu.registers[6][14] ),
    .A2(net3951),
    .A1(\cpu.registers[5][14] ));
 sg13g2_a22oi_1 _09196_ (.Y(_02730_),
    .B1(net3953),
    .B2(\cpu.registers[3][14] ),
    .A2(net3957),
    .A1(\cpu.registers[2][14] ));
 sg13g2_and3_2 _09197_ (.X(_02731_),
    .A(_02728_),
    .B(_02729_),
    .C(_02730_));
 sg13g2_inv_1 _09198_ (.Y(_02732_),
    .A(_02731_));
 sg13g2_o21ai_1 _09199_ (.B1(_02726_),
    .Y(_00598_),
    .A1(_02641_),
    .A2(_02731_));
 sg13g2_nand2_1 _09200_ (.Y(_02733_),
    .A(net451),
    .B(net3748));
 sg13g2_nor2_1 _09201_ (.A(_00048_),
    .B(net3947),
    .Y(_02734_));
 sg13g2_a221oi_1 _09202_ (.B2(\cpu.registers[6][15] ),
    .C1(_02734_),
    .B1(net3949),
    .A1(\cpu.registers[1][15] ),
    .Y(_02735_),
    .A2(net3955));
 sg13g2_a22oi_1 _09203_ (.Y(_02736_),
    .B1(net3953),
    .B2(\cpu.registers[3][15] ),
    .A2(net3957),
    .A1(\cpu.registers[2][15] ));
 sg13g2_a22oi_1 _09204_ (.Y(_02737_),
    .B1(net3951),
    .B2(\cpu.registers[5][15] ),
    .A2(net4095),
    .A1(\cpu.registers[4][15] ));
 sg13g2_and3_2 _09205_ (.X(_02738_),
    .A(_02735_),
    .B(_02736_),
    .C(_02737_));
 sg13g2_inv_1 _09206_ (.Y(_02739_),
    .A(_02738_));
 sg13g2_o21ai_1 _09207_ (.B1(_02733_),
    .Y(_00599_),
    .A1(_02641_),
    .A2(_02738_));
 sg13g2_nor3_2 _09208_ (.A(_00018_),
    .B(_01257_),
    .C(net4039),
    .Y(_02740_));
 sg13g2_inv_1 _09209_ (.Y(_02741_),
    .A(_02740_));
 sg13g2_nor2_1 _09210_ (.A(_00018_),
    .B(_01233_),
    .Y(_02742_));
 sg13g2_a22oi_1 _09211_ (.Y(_02743_),
    .B1(_02740_),
    .B2(net3803),
    .A2(_02626_),
    .A1(net4143));
 sg13g2_o21ai_1 _09212_ (.B1(_02627_),
    .Y(_02744_),
    .A1(net3799),
    .A2(_02741_));
 sg13g2_nand2_1 _09213_ (.Y(_02745_),
    .A(net4465),
    .B(net3745));
 sg13g2_o21ai_1 _09214_ (.B1(net4307),
    .Y(_02746_),
    .A1(_00049_),
    .A2(net4036));
 sg13g2_a221oi_1 _09215_ (.B2(_02161_),
    .C1(_02746_),
    .B1(net3752),
    .A1(\cpu.current_address[0] ),
    .Y(_02747_),
    .A2(net3799));
 sg13g2_o21ai_1 _09216_ (.B1(net3747),
    .Y(_02748_),
    .A1(net4309),
    .A2(net824));
 sg13g2_o21ai_1 _09217_ (.B1(_02745_),
    .Y(_00600_),
    .A1(_02747_),
    .A2(_02748_));
 sg13g2_nand2_1 _09218_ (.Y(_02749_),
    .A(net4463),
    .B(net3745));
 sg13g2_o21ai_1 _09219_ (.B1(net4310),
    .Y(_02750_),
    .A1(_00050_),
    .A2(net4037));
 sg13g2_a221oi_1 _09220_ (.B2(_02168_),
    .C1(_02750_),
    .B1(net3751),
    .A1(net819),
    .Y(_02751_),
    .A2(net3798));
 sg13g2_o21ai_1 _09221_ (.B1(net3747),
    .Y(_02752_),
    .A1(net4309),
    .A2(\cpu.request_address[1] ));
 sg13g2_o21ai_1 _09222_ (.B1(_02749_),
    .Y(_00601_),
    .A1(_02751_),
    .A2(_02752_));
 sg13g2_nand2_1 _09223_ (.Y(_02753_),
    .A(net4461),
    .B(net3745));
 sg13g2_o21ai_1 _09224_ (.B1(net4309),
    .Y(_02754_),
    .A1(_00051_),
    .A2(net4036));
 sg13g2_a221oi_1 _09225_ (.B2(_02176_),
    .C1(_02754_),
    .B1(net3752),
    .A1(net466),
    .Y(_02755_),
    .A2(net3799));
 sg13g2_o21ai_1 _09226_ (.B1(net3747),
    .Y(_02756_),
    .A1(net4309),
    .A2(net875));
 sg13g2_o21ai_1 _09227_ (.B1(_02753_),
    .Y(_00602_),
    .A1(_02755_),
    .A2(_02756_));
 sg13g2_nand2_1 _09228_ (.Y(_02757_),
    .A(net4460),
    .B(net3745));
 sg13g2_o21ai_1 _09229_ (.B1(net4310),
    .Y(_02758_),
    .A1(_00052_),
    .A2(net4036));
 sg13g2_a221oi_1 _09230_ (.B2(_02184_),
    .C1(_02758_),
    .B1(net3751),
    .A1(net145),
    .Y(_02759_),
    .A2(net3800));
 sg13g2_o21ai_1 _09231_ (.B1(net3747),
    .Y(_02760_),
    .A1(net4310),
    .A2(\cpu.request_address[3] ));
 sg13g2_o21ai_1 _09232_ (.B1(_02757_),
    .Y(_00603_),
    .A1(_02759_),
    .A2(_02760_));
 sg13g2_nand2_1 _09233_ (.Y(_02761_),
    .A(net4458),
    .B(net3745));
 sg13g2_o21ai_1 _09234_ (.B1(net4310),
    .Y(_02762_),
    .A1(_00053_),
    .A2(net4036));
 sg13g2_a221oi_1 _09235_ (.B2(_02192_),
    .C1(_02762_),
    .B1(net3751),
    .A1(net136),
    .Y(_02763_),
    .A2(net3800));
 sg13g2_o21ai_1 _09236_ (.B1(net3747),
    .Y(_02764_),
    .A1(net4310),
    .A2(\cpu.request_address[4] ));
 sg13g2_o21ai_1 _09237_ (.B1(_02761_),
    .Y(_00604_),
    .A1(_02763_),
    .A2(_02764_));
 sg13g2_nand2_1 _09238_ (.Y(_02765_),
    .A(net4455),
    .B(net3745));
 sg13g2_o21ai_1 _09239_ (.B1(net4309),
    .Y(_02766_),
    .A1(_00054_),
    .A2(net4037));
 sg13g2_a221oi_1 _09240_ (.B2(_02199_),
    .C1(_02766_),
    .B1(net3751),
    .A1(net158),
    .Y(_02767_),
    .A2(net3798));
 sg13g2_o21ai_1 _09241_ (.B1(net3747),
    .Y(_02768_),
    .A1(net4311),
    .A2(\cpu.request_address[5] ));
 sg13g2_o21ai_1 _09242_ (.B1(_02765_),
    .Y(_00605_),
    .A1(_02767_),
    .A2(_02768_));
 sg13g2_nand2_1 _09243_ (.Y(_02769_),
    .A(net427),
    .B(net3745));
 sg13g2_o21ai_1 _09244_ (.B1(net4310),
    .Y(_02770_),
    .A1(_00055_),
    .A2(net4036));
 sg13g2_a221oi_1 _09245_ (.B2(_02207_),
    .C1(_02770_),
    .B1(net3751),
    .A1(net142),
    .Y(_02771_),
    .A2(net3798));
 sg13g2_o21ai_1 _09246_ (.B1(net3747),
    .Y(_02772_),
    .A1(net4310),
    .A2(\cpu.request_address[6] ));
 sg13g2_o21ai_1 _09247_ (.B1(_02769_),
    .Y(_00606_),
    .A1(_02771_),
    .A2(_02772_));
 sg13g2_nand2_1 _09248_ (.Y(_02773_),
    .A(net4453),
    .B(net3745));
 sg13g2_o21ai_1 _09249_ (.B1(net4309),
    .Y(_02774_),
    .A1(_00056_),
    .A2(net4036));
 sg13g2_a221oi_1 _09250_ (.B2(_02215_),
    .C1(_02774_),
    .B1(net3751),
    .A1(net541),
    .Y(_02775_),
    .A2(net3798));
 sg13g2_o21ai_1 _09251_ (.B1(net3747),
    .Y(_02776_),
    .A1(net4311),
    .A2(\cpu.request_address[7] ));
 sg13g2_o21ai_1 _09252_ (.B1(_02773_),
    .Y(_00607_),
    .A1(_02775_),
    .A2(_02776_));
 sg13g2_nand2_1 _09253_ (.Y(_02777_),
    .A(net868),
    .B(net3744));
 sg13g2_o21ai_1 _09254_ (.B1(net4304),
    .Y(_02778_),
    .A1(_00057_),
    .A2(net4035));
 sg13g2_a221oi_1 _09255_ (.B2(_02223_),
    .C1(_02778_),
    .B1(net3750),
    .A1(net235),
    .Y(_02779_),
    .A2(net3796));
 sg13g2_o21ai_1 _09256_ (.B1(net3746),
    .Y(_02780_),
    .A1(net4305),
    .A2(net855));
 sg13g2_o21ai_1 _09257_ (.B1(_02777_),
    .Y(_00608_),
    .A1(_02779_),
    .A2(_02780_));
 sg13g2_nand2_1 _09258_ (.Y(_02781_),
    .A(net833),
    .B(net3744));
 sg13g2_o21ai_1 _09259_ (.B1(net4308),
    .Y(_02782_),
    .A1(_00058_),
    .A2(net4035));
 sg13g2_a221oi_1 _09260_ (.B2(_02230_),
    .C1(_02782_),
    .B1(net3750),
    .A1(net130),
    .Y(_02783_),
    .A2(net3797));
 sg13g2_o21ai_1 _09261_ (.B1(net3746),
    .Y(_02784_),
    .A1(net4305),
    .A2(net743));
 sg13g2_o21ai_1 _09262_ (.B1(_02781_),
    .Y(_00609_),
    .A1(_02783_),
    .A2(_02784_));
 sg13g2_nand2_1 _09263_ (.Y(_02785_),
    .A(net867),
    .B(net3744));
 sg13g2_o21ai_1 _09264_ (.B1(net4304),
    .Y(_02786_),
    .A1(_00059_),
    .A2(net4035));
 sg13g2_a221oi_1 _09265_ (.B2(_02237_),
    .C1(_02786_),
    .B1(net3750),
    .A1(net355),
    .Y(_02787_),
    .A2(net3796));
 sg13g2_o21ai_1 _09266_ (.B1(net3746),
    .Y(_02788_),
    .A1(net4304),
    .A2(net717));
 sg13g2_o21ai_1 _09267_ (.B1(_02785_),
    .Y(_00610_),
    .A1(_02787_),
    .A2(_02788_));
 sg13g2_nand2_1 _09268_ (.Y(_02789_),
    .A(net815),
    .B(net3744));
 sg13g2_o21ai_1 _09269_ (.B1(net4305),
    .Y(_02790_),
    .A1(_00060_),
    .A2(net4035));
 sg13g2_a221oi_1 _09270_ (.B2(_02244_),
    .C1(_02790_),
    .B1(net3750),
    .A1(net319),
    .Y(_02791_),
    .A2(net3797));
 sg13g2_o21ai_1 _09271_ (.B1(net3746),
    .Y(_02792_),
    .A1(net4305),
    .A2(net584));
 sg13g2_o21ai_1 _09272_ (.B1(_02789_),
    .Y(_00611_),
    .A1(_02791_),
    .A2(_02792_));
 sg13g2_nand2_1 _09273_ (.Y(_02793_),
    .A(net744),
    .B(net3744));
 sg13g2_o21ai_1 _09274_ (.B1(net4305),
    .Y(_02794_),
    .A1(_00061_),
    .A2(net4035));
 sg13g2_a221oi_1 _09275_ (.B2(_02251_),
    .C1(_02794_),
    .B1(net3750),
    .A1(net317),
    .Y(_02795_),
    .A2(net3797));
 sg13g2_o21ai_1 _09276_ (.B1(net3746),
    .Y(_02796_),
    .A1(net4305),
    .A2(net611));
 sg13g2_o21ai_1 _09277_ (.B1(_02793_),
    .Y(_00612_),
    .A1(_02795_),
    .A2(_02796_));
 sg13g2_nand2_1 _09278_ (.Y(_02797_),
    .A(net853),
    .B(net3744));
 sg13g2_nor2_1 _09279_ (.A(_00046_),
    .B(net3981),
    .Y(_02798_));
 sg13g2_a221oi_1 _09280_ (.B2(\cpu.registers[2][13] ),
    .C1(_02798_),
    .B1(net3969),
    .A1(\cpu.registers[4][13] ),
    .Y(_02799_),
    .A2(net3971));
 sg13g2_a22oi_1 _09281_ (.Y(_02800_),
    .B1(net3975),
    .B2(\cpu.registers[6][13] ),
    .A2(net3977),
    .A1(\cpu.registers[5][13] ));
 sg13g2_a22oi_1 _09282_ (.Y(_02801_),
    .B1(net3973),
    .B2(\cpu.registers[3][13] ),
    .A2(net3979),
    .A1(\cpu.registers[1][13] ));
 sg13g2_and3_1 _09283_ (.X(_02802_),
    .A(_02799_),
    .B(_02800_),
    .C(_02801_));
 sg13g2_inv_1 _09284_ (.Y(_02803_),
    .A(_02802_));
 sg13g2_o21ai_1 _09285_ (.B1(net4304),
    .Y(_02804_),
    .A1(_00062_),
    .A2(net4035));
 sg13g2_a221oi_1 _09286_ (.B2(_02803_),
    .C1(_02804_),
    .B1(net3750),
    .A1(net324),
    .Y(_02805_),
    .A2(net3796));
 sg13g2_o21ai_1 _09287_ (.B1(net3746),
    .Y(_02806_),
    .A1(net4304),
    .A2(net763));
 sg13g2_o21ai_1 _09288_ (.B1(_02797_),
    .Y(_00613_),
    .A1(_02805_),
    .A2(_02806_));
 sg13g2_nand2_1 _09289_ (.Y(_02807_),
    .A(net663),
    .B(net3744));
 sg13g2_or2_1 _09290_ (.X(_02808_),
    .B(net3981),
    .A(_00047_));
 sg13g2_a22oi_1 _09291_ (.Y(_02809_),
    .B1(net3977),
    .B2(\cpu.registers[5][14] ),
    .A2(net3979),
    .A1(\cpu.registers[1][14] ));
 sg13g2_a22oi_1 _09292_ (.Y(_02810_),
    .B1(net3969),
    .B2(\cpu.registers[2][14] ),
    .A2(net3973),
    .A1(\cpu.registers[3][14] ));
 sg13g2_a22oi_1 _09293_ (.Y(_02811_),
    .B1(net3971),
    .B2(\cpu.registers[4][14] ),
    .A2(net3975),
    .A1(\cpu.registers[6][14] ));
 sg13g2_nand4_1 _09294_ (.B(_02809_),
    .C(_02810_),
    .A(_02808_),
    .Y(_02812_),
    .D(_02811_));
 sg13g2_o21ai_1 _09295_ (.B1(net4304),
    .Y(_02813_),
    .A1(_00063_),
    .A2(net4035));
 sg13g2_a221oi_1 _09296_ (.B2(_02812_),
    .C1(_02813_),
    .B1(net3750),
    .A1(\cpu.current_address[14] ),
    .Y(_02814_),
    .A2(net3796));
 sg13g2_o21ai_1 _09297_ (.B1(net3746),
    .Y(_02815_),
    .A1(net4305),
    .A2(\cpu.request_address[14] ));
 sg13g2_o21ai_1 _09298_ (.B1(_02807_),
    .Y(_00614_),
    .A1(_02814_),
    .A2(_02815_));
 sg13g2_nand2_1 _09299_ (.Y(_02816_),
    .A(net803),
    .B(net3744));
 sg13g2_nor2_1 _09300_ (.A(_00048_),
    .B(net3981),
    .Y(_02817_));
 sg13g2_a221oi_1 _09301_ (.B2(\cpu.registers[2][15] ),
    .C1(_02817_),
    .B1(net3969),
    .A1(\cpu.registers[6][15] ),
    .Y(_02818_),
    .A2(net3975));
 sg13g2_a22oi_1 _09302_ (.Y(_02819_),
    .B1(net3971),
    .B2(\cpu.registers[4][15] ),
    .A2(net3979),
    .A1(\cpu.registers[1][15] ));
 sg13g2_a22oi_1 _09303_ (.Y(_02820_),
    .B1(net3973),
    .B2(\cpu.registers[3][15] ),
    .A2(net3977),
    .A1(\cpu.registers[5][15] ));
 sg13g2_nand3_1 _09304_ (.B(_02819_),
    .C(_02820_),
    .A(_02818_),
    .Y(_02821_));
 sg13g2_o21ai_1 _09305_ (.B1(net4304),
    .Y(_02822_),
    .A1(_00064_),
    .A2(net4035));
 sg13g2_a221oi_1 _09306_ (.B2(_02821_),
    .C1(_02822_),
    .B1(net3750),
    .A1(net470),
    .Y(_02823_),
    .A2(net3796));
 sg13g2_o21ai_1 _09307_ (.B1(net3746),
    .Y(_02824_),
    .A1(net4304),
    .A2(net357));
 sg13g2_o21ai_1 _09308_ (.B1(_02816_),
    .Y(_00615_),
    .A1(_02823_),
    .A2(_02824_));
 sg13g2_nor2_1 _09309_ (.A(net4307),
    .B(\cpu.execution_stage[1] ),
    .Y(_02825_));
 sg13g2_nor2_2 _09310_ (.A(_02740_),
    .B(_02825_),
    .Y(_02826_));
 sg13g2_nand2_1 _09311_ (.Y(_02827_),
    .A(net789),
    .B(net4037));
 sg13g2_nor2_1 _09312_ (.A(_00017_),
    .B(_02827_),
    .Y(_02828_));
 sg13g2_mux2_1 _09313_ (.A0(\cpu.ALU.mode[0] ),
    .A1(net790),
    .S(_02826_),
    .X(_00616_));
 sg13g2_o21ai_1 _09314_ (.B1(_00894_),
    .Y(_02829_),
    .A1(net4449),
    .A2(net4038));
 sg13g2_a21oi_1 _09315_ (.A1(net4239),
    .A2(net4038),
    .Y(_02830_),
    .B1(_02829_));
 sg13g2_mux2_1 _09316_ (.A0(net792),
    .A1(_02830_),
    .S(_02826_),
    .X(_00617_));
 sg13g2_nor2_1 _09317_ (.A(_00026_),
    .B(_02827_),
    .Y(_02831_));
 sg13g2_mux2_1 _09318_ (.A0(net68),
    .A1(_02831_),
    .S(_02826_),
    .X(_00618_));
 sg13g2_mux2_1 _09319_ (.A0(net203),
    .A1(net73),
    .S(net4023),
    .X(_00619_));
 sg13g2_mux2_1 _09320_ (.A0(net268),
    .A1(net75),
    .S(net4022),
    .X(_00620_));
 sg13g2_mux2_1 _09321_ (.A0(net238),
    .A1(net52),
    .S(net4023),
    .X(_00621_));
 sg13g2_mux2_1 _09322_ (.A0(net208),
    .A1(net67),
    .S(net4023),
    .X(_00622_));
 sg13g2_nor2_1 _09323_ (.A(net54),
    .B(net4141),
    .Y(_02832_));
 sg13g2_a21oi_1 _09324_ (.A1(net4238),
    .A2(net4140),
    .Y(_00623_),
    .B1(_02832_));
 sg13g2_mux2_1 _09325_ (.A0(net121),
    .A1(net65),
    .S(net4023),
    .X(_00624_));
 sg13g2_mux2_1 _09326_ (.A0(net351),
    .A1(net79),
    .S(net4022),
    .X(_00625_));
 sg13g2_mux2_1 _09327_ (.A0(net4445),
    .A1(net91),
    .S(net4022),
    .X(_00626_));
 sg13g2_mux2_1 _09328_ (.A0(net4440),
    .A1(net61),
    .S(net4022),
    .X(_00627_));
 sg13g2_nor2_1 _09329_ (.A(net53),
    .B(net4141),
    .Y(_02833_));
 sg13g2_a21oi_2 _09330_ (.B1(_02833_),
    .Y(_00628_),
    .A2(net4141),
    .A1(net4201));
 sg13g2_mux2_1 _09331_ (.A0(net4433),
    .A1(net71),
    .S(net4022),
    .X(_00629_));
 sg13g2_mux2_1 _09332_ (.A0(net4431),
    .A1(net64),
    .S(net4022),
    .X(_00630_));
 sg13g2_mux2_1 _09333_ (.A0(net4418),
    .A1(net120),
    .S(net4022),
    .X(_00631_));
 sg13g2_mux2_1 _09334_ (.A0(net4396),
    .A1(net78),
    .S(net4022),
    .X(_00632_));
 sg13g2_nor2_1 _09335_ (.A(net241),
    .B(net4140),
    .Y(_02834_));
 sg13g2_a21oi_1 _09336_ (.A1(net4216),
    .A2(net4140),
    .Y(_00633_),
    .B1(_02834_));
 sg13g2_nor2_1 _09337_ (.A(net92),
    .B(net4140),
    .Y(_02835_));
 sg13g2_a21oi_1 _09338_ (.A1(net4208),
    .A2(net4140),
    .Y(_00634_),
    .B1(_02835_));
 sg13g2_mux2_1 _09339_ (.A0(net677),
    .A1(\cpu.request_address[0] ),
    .S(net4024),
    .X(_00635_));
 sg13g2_mux2_1 _09340_ (.A0(net819),
    .A1(\cpu.request_address[1] ),
    .S(net4024),
    .X(_00636_));
 sg13g2_nand2_1 _09341_ (.Y(_02836_),
    .A(net466),
    .B(net4143));
 sg13g2_o21ai_1 _09342_ (.B1(_02836_),
    .Y(_00637_),
    .A1(_01146_),
    .A2(net4143));
 sg13g2_nand2_1 _09343_ (.Y(_02837_),
    .A(net145),
    .B(net4143));
 sg13g2_o21ai_1 _09344_ (.B1(_02837_),
    .Y(_00638_),
    .A1(_01147_),
    .A2(net4142));
 sg13g2_nand2_1 _09345_ (.Y(_02838_),
    .A(net136),
    .B(net4143));
 sg13g2_o21ai_1 _09346_ (.B1(_02838_),
    .Y(_00639_),
    .A1(_01148_),
    .A2(net4142));
 sg13g2_nand2_1 _09347_ (.Y(_02839_),
    .A(net158),
    .B(net4142));
 sg13g2_o21ai_1 _09348_ (.B1(_02839_),
    .Y(_00640_),
    .A1(_01149_),
    .A2(net4142));
 sg13g2_nand2_1 _09349_ (.Y(_02840_),
    .A(net142),
    .B(net4142));
 sg13g2_o21ai_1 _09350_ (.B1(_02840_),
    .Y(_00641_),
    .A1(_01150_),
    .A2(net4142));
 sg13g2_nor2_1 _09351_ (.A(\cpu.request_address[7] ),
    .B(net4142),
    .Y(_02841_));
 sg13g2_a21oi_1 _09352_ (.A1(_01151_),
    .A2(net4142),
    .Y(_00642_),
    .B1(_02841_));
 sg13g2_nor2_1 _09353_ (.A(\cpu.request_address[8] ),
    .B(net4138),
    .Y(_02842_));
 sg13g2_a21oi_1 _09354_ (.A1(_01153_),
    .A2(net4138),
    .Y(_00643_),
    .B1(_02842_));
 sg13g2_nand2_1 _09355_ (.Y(_02843_),
    .A(net130),
    .B(net4140));
 sg13g2_o21ai_1 _09356_ (.B1(_02843_),
    .Y(_00644_),
    .A1(_01154_),
    .A2(net4140));
 sg13g2_nor2_1 _09357_ (.A(\cpu.request_address[10] ),
    .B(net4138),
    .Y(_02844_));
 sg13g2_a21oi_1 _09358_ (.A1(_01155_),
    .A2(net4138),
    .Y(_00645_),
    .B1(_02844_));
 sg13g2_nor2_1 _09359_ (.A(\cpu.request_address[11] ),
    .B(net4139),
    .Y(_02845_));
 sg13g2_a21oi_1 _09360_ (.A1(_01157_),
    .A2(net4139),
    .Y(_00646_),
    .B1(_02845_));
 sg13g2_nor2_1 _09361_ (.A(\cpu.request_address[12] ),
    .B(net4139),
    .Y(_02846_));
 sg13g2_a21oi_1 _09362_ (.A1(_01159_),
    .A2(net4139),
    .Y(_00647_),
    .B1(_02846_));
 sg13g2_nor2_1 _09363_ (.A(\cpu.request_address[13] ),
    .B(net4139),
    .Y(_02847_));
 sg13g2_a21oi_1 _09364_ (.A1(_01161_),
    .A2(net4139),
    .Y(_00648_),
    .B1(_02847_));
 sg13g2_nand2_1 _09365_ (.Y(_02848_),
    .A(net140),
    .B(net4138));
 sg13g2_o21ai_1 _09366_ (.B1(_02848_),
    .Y(_00649_),
    .A1(_01163_),
    .A2(net4138));
 sg13g2_nor2_1 _09367_ (.A(net357),
    .B(net4138),
    .Y(_02849_));
 sg13g2_a21oi_1 _09368_ (.A1(_01164_),
    .A2(net4138),
    .Y(_00650_),
    .B1(_02849_));
 sg13g2_nand2b_1 _09369_ (.Y(_02850_),
    .B(net4427),
    .A_N(\cpu.keccak_alu.registers[144] ));
 sg13g2_o21ai_1 _09370_ (.B1(_02850_),
    .Y(_02851_),
    .A1(net4427),
    .A2(net4575));
 sg13g2_a22oi_1 _09371_ (.Y(_02852_),
    .B1(net4107),
    .B2(net4497),
    .A2(net4120),
    .A1(\cpu.keccak_alu.registers[176] ));
 sg13g2_o21ai_1 _09372_ (.B1(_02852_),
    .Y(_02853_),
    .A1(net4400),
    .A2(_02851_));
 sg13g2_nand2b_1 _09373_ (.Y(_02854_),
    .B(net4428),
    .A_N(\cpu.keccak_alu.registers[80] ));
 sg13g2_o21ai_1 _09374_ (.B1(_02854_),
    .Y(_02855_),
    .A1(net4428),
    .A2(\cpu.keccak_alu.registers[64] ));
 sg13g2_a22oi_1 _09375_ (.Y(_02856_),
    .B1(net4107),
    .B2(\cpu.keccak_alu.registers[96] ),
    .A2(net4120),
    .A1(\cpu.keccak_alu.registers[112] ));
 sg13g2_o21ai_1 _09376_ (.B1(_02856_),
    .Y(_02857_),
    .A1(net4400),
    .A2(_02855_));
 sg13g2_a22oi_1 _09377_ (.Y(_02858_),
    .B1(_02857_),
    .B2(_02146_),
    .A2(_02853_),
    .A1(_02151_));
 sg13g2_a21oi_1 _09378_ (.A1(net4427),
    .A2(_00998_),
    .Y(_02859_),
    .B1(net4400));
 sg13g2_o21ai_1 _09379_ (.B1(_02859_),
    .Y(_02860_),
    .A1(net4427),
    .A2(\cpu.keccak_alu.registers[256] ));
 sg13g2_a22oi_1 _09380_ (.Y(_02861_),
    .B1(net4107),
    .B2(\cpu.keccak_alu.registers[288] ),
    .A2(net4120),
    .A1(\cpu.keccak_alu.registers[304] ));
 sg13g2_nand3_1 _09381_ (.B(_02860_),
    .C(_02861_),
    .A(net4438),
    .Y(_02862_));
 sg13g2_a21oi_1 _09382_ (.A1(net4427),
    .A2(_00996_),
    .Y(_02863_),
    .B1(net4400));
 sg13g2_o21ai_1 _09383_ (.B1(_02863_),
    .Y(_02864_),
    .A1(net4427),
    .A2(\cpu.keccak_alu.registers[0] ));
 sg13g2_a221oi_1 _09384_ (.B2(\cpu.keccak_alu.registers[32] ),
    .C1(net4438),
    .B1(net4107),
    .A1(\cpu.keccak_alu.registers[48] ),
    .Y(_02865_),
    .A2(net4120));
 sg13g2_a21oi_1 _09385_ (.A1(_02864_),
    .A2(_02865_),
    .Y(_02866_),
    .B1(net4124));
 sg13g2_nand2b_1 _09386_ (.Y(_02867_),
    .B(net4427),
    .A_N(\cpu.keccak_alu.registers[208] ));
 sg13g2_o21ai_1 _09387_ (.B1(_02867_),
    .Y(_02868_),
    .A1(net4427),
    .A2(\cpu.keccak_alu.registers[192] ));
 sg13g2_a22oi_1 _09388_ (.Y(_02869_),
    .B1(net4107),
    .B2(\cpu.keccak_alu.registers[224] ),
    .A2(net4120),
    .A1(\cpu.keccak_alu.registers[240] ));
 sg13g2_o21ai_1 _09389_ (.B1(_02869_),
    .Y(_02870_),
    .A1(net4400),
    .A2(_02868_));
 sg13g2_a22oi_1 _09390_ (.Y(_02871_),
    .B1(_02870_),
    .B2(net3974),
    .A2(_02866_),
    .A1(_02862_));
 sg13g2_o21ai_1 _09391_ (.B1(_02871_),
    .Y(_02872_),
    .A1(net4438),
    .A2(_02858_));
 sg13g2_a21oi_2 _09392_ (.B1(net4070),
    .Y(_02873_),
    .A2(_02872_),
    .A1(_02259_));
 sg13g2_nor2_1 _09393_ (.A(net4074),
    .B(_02621_),
    .Y(_02874_));
 sg13g2_a21oi_1 _09394_ (.A1(net4307),
    .A2(_01251_),
    .Y(_02875_),
    .B1(_02825_));
 sg13g2_nand2b_2 _09395_ (.Y(_02876_),
    .B(_02875_),
    .A_N(_02742_));
 sg13g2_nor4_2 _09396_ (.A(\cpu.execution_stage[1] ),
    .B(_02873_),
    .C(_02874_),
    .Y(_02877_),
    .D(net3743));
 sg13g2_a21o_1 _09397_ (.A2(net3743),
    .A1(net694),
    .B1(_02877_),
    .X(_00651_));
 sg13g2_nand2_1 _09398_ (.Y(_02878_),
    .A(net393),
    .B(_02876_));
 sg13g2_nand3b_1 _09399_ (.B(_02875_),
    .C(_00045_),
    .Y(_02879_),
    .A_N(_02742_));
 sg13g2_nand2b_1 _09400_ (.Y(_02880_),
    .B(net4426),
    .A_N(\cpu.keccak_alu.registers[17] ));
 sg13g2_o21ai_1 _09401_ (.B1(_02880_),
    .Y(_02881_),
    .A1(net4426),
    .A2(\cpu.keccak_alu.registers[1] ));
 sg13g2_a221oi_1 _09402_ (.B2(\cpu.keccak_alu.registers[33] ),
    .C1(net4437),
    .B1(net4108),
    .A1(\cpu.keccak_alu.registers[49] ),
    .Y(_02882_),
    .A2(net4121));
 sg13g2_o21ai_1 _09403_ (.B1(_02882_),
    .Y(_02883_),
    .A1(net4399),
    .A2(_02881_));
 sg13g2_nand2b_1 _09404_ (.Y(_02884_),
    .B(net4426),
    .A_N(\cpu.keccak_alu.registers[209] ));
 sg13g2_o21ai_1 _09405_ (.B1(_02884_),
    .Y(_02885_),
    .A1(net4426),
    .A2(\cpu.keccak_alu.registers[193] ));
 sg13g2_a22oi_1 _09406_ (.Y(_02886_),
    .B1(net4108),
    .B2(\cpu.keccak_alu.registers[225] ),
    .A2(net4121),
    .A1(\cpu.keccak_alu.registers[241] ));
 sg13g2_o21ai_1 _09407_ (.B1(_02886_),
    .Y(_02887_),
    .A1(net4399),
    .A2(_02885_));
 sg13g2_nand2b_1 _09408_ (.Y(_02888_),
    .B(net4426),
    .A_N(\cpu.keccak_alu.registers[81] ));
 sg13g2_o21ai_1 _09409_ (.B1(_02888_),
    .Y(_02889_),
    .A1(net4426),
    .A2(\cpu.keccak_alu.registers[65] ));
 sg13g2_a22oi_1 _09410_ (.Y(_02890_),
    .B1(net4108),
    .B2(\cpu.keccak_alu.registers[97] ),
    .A2(net4121),
    .A1(\cpu.keccak_alu.registers[113] ));
 sg13g2_o21ai_1 _09411_ (.B1(_02890_),
    .Y(_02891_),
    .A1(net4401),
    .A2(_02889_));
 sg13g2_mux2_1 _09412_ (.A0(_01003_),
    .A1(_01004_),
    .S(net4426),
    .X(_02892_));
 sg13g2_a22oi_1 _09413_ (.Y(_02893_),
    .B1(net4108),
    .B2(\cpu.keccak_alu.registers[161] ),
    .A2(net4121),
    .A1(\cpu.keccak_alu.registers[177] ));
 sg13g2_o21ai_1 _09414_ (.B1(_02893_),
    .Y(_02894_),
    .A1(net4399),
    .A2(_02892_));
 sg13g2_a22oi_1 _09415_ (.Y(_02895_),
    .B1(_02891_),
    .B2(net4131),
    .A2(_02887_),
    .A1(_02142_));
 sg13g2_a22oi_1 _09416_ (.Y(_02896_),
    .B1(_02894_),
    .B2(_02151_),
    .A2(_02883_),
    .A1(net4127));
 sg13g2_mux2_1 _09417_ (.A0(_01005_),
    .A1(_01006_),
    .S(net4423),
    .X(_02897_));
 sg13g2_a22oi_1 _09418_ (.Y(_02898_),
    .B1(net4108),
    .B2(\cpu.keccak_alu.registers[289] ),
    .A2(net4121),
    .A1(\cpu.keccak_alu.registers[305] ));
 sg13g2_o21ai_1 _09419_ (.B1(_02898_),
    .Y(_02899_),
    .A1(net4399),
    .A2(_02897_));
 sg13g2_nand2_1 _09420_ (.Y(_02900_),
    .A(net4126),
    .B(_02899_));
 sg13g2_nand2_1 _09421_ (.Y(_02901_),
    .A(net4074),
    .B(_02259_));
 sg13g2_a221oi_1 _09422_ (.B2(net4438),
    .C1(net3847),
    .B1(_02900_),
    .A1(_02895_),
    .Y(_02902_),
    .A2(_02896_));
 sg13g2_a21oi_2 _09423_ (.B1(_02902_),
    .Y(_02903_),
    .A2(_02638_),
    .A1(net4072));
 sg13g2_o21ai_1 _09424_ (.B1(_02878_),
    .Y(_00652_),
    .A1(net3741),
    .A2(_02903_));
 sg13g2_nand2_1 _09425_ (.Y(_02904_),
    .A(net111),
    .B(net3743));
 sg13g2_a21oi_1 _09426_ (.A1(net4423),
    .A2(_01009_),
    .Y(_02905_),
    .B1(net4399));
 sg13g2_o21ai_1 _09427_ (.B1(_02905_),
    .Y(_02906_),
    .A1(net4423),
    .A2(\cpu.keccak_alu.registers[2] ));
 sg13g2_a22oi_1 _09428_ (.Y(_02907_),
    .B1(net4106),
    .B2(\cpu.keccak_alu.registers[34] ),
    .A2(net4119),
    .A1(\cpu.keccak_alu.registers[50] ));
 sg13g2_nand3_1 _09429_ (.B(_02906_),
    .C(_02907_),
    .A(_00906_),
    .Y(_02908_));
 sg13g2_nand2b_1 _09430_ (.Y(_02909_),
    .B(net4423),
    .A_N(\cpu.keccak_alu.registers[82] ));
 sg13g2_o21ai_1 _09431_ (.B1(_02909_),
    .Y(_02910_),
    .A1(net4423),
    .A2(\cpu.keccak_alu.registers[66] ));
 sg13g2_a22oi_1 _09432_ (.Y(_02911_),
    .B1(net4107),
    .B2(\cpu.keccak_alu.registers[98] ),
    .A2(net4120),
    .A1(\cpu.keccak_alu.registers[114] ));
 sg13g2_o21ai_1 _09433_ (.B1(_02911_),
    .Y(_02912_),
    .A1(net4399),
    .A2(_02910_));
 sg13g2_nand2b_1 _09434_ (.Y(_02913_),
    .B(net4423),
    .A_N(\cpu.keccak_alu.registers[210] ));
 sg13g2_o21ai_1 _09435_ (.B1(_02913_),
    .Y(_02914_),
    .A1(net4423),
    .A2(\cpu.keccak_alu.registers[194] ));
 sg13g2_a22oi_1 _09436_ (.Y(_02915_),
    .B1(net4106),
    .B2(\cpu.keccak_alu.registers[226] ),
    .A2(net4119),
    .A1(\cpu.keccak_alu.registers[242] ));
 sg13g2_o21ai_1 _09437_ (.B1(_02915_),
    .Y(_02916_),
    .A1(net4399),
    .A2(_02914_));
 sg13g2_mux2_1 _09438_ (.A0(net4188),
    .A1(_01012_),
    .S(net4423),
    .X(_02917_));
 sg13g2_a22oi_1 _09439_ (.Y(_02918_),
    .B1(net4106),
    .B2(\cpu.keccak_alu.registers[162] ),
    .A2(net4119),
    .A1(\cpu.keccak_alu.registers[178] ));
 sg13g2_o21ai_1 _09440_ (.B1(_02918_),
    .Y(_02919_),
    .A1(net4399),
    .A2(_02917_));
 sg13g2_a22oi_1 _09441_ (.Y(_02920_),
    .B1(_02916_),
    .B2(_02142_),
    .A2(_02912_),
    .A1(net4131));
 sg13g2_a22oi_1 _09442_ (.Y(_02921_),
    .B1(_02919_),
    .B2(_02151_),
    .A2(_02908_),
    .A1(net4127));
 sg13g2_mux2_1 _09443_ (.A0(_01013_),
    .A1(_01014_),
    .S(net4424),
    .X(_02922_));
 sg13g2_a22oi_1 _09444_ (.Y(_02923_),
    .B1(net4106),
    .B2(\cpu.keccak_alu.registers[290] ),
    .A2(net4119),
    .A1(\cpu.keccak_alu.registers[306] ));
 sg13g2_o21ai_1 _09445_ (.B1(_02923_),
    .Y(_02924_),
    .A1(net4400),
    .A2(_02922_));
 sg13g2_nand2_1 _09446_ (.Y(_02925_),
    .A(net4126),
    .B(_02924_));
 sg13g2_a221oi_1 _09447_ (.B2(net4438),
    .C1(net3847),
    .B1(_02925_),
    .A1(_02920_),
    .Y(_02926_),
    .A2(_02921_));
 sg13g2_a21oi_2 _09448_ (.B1(_02926_),
    .Y(_02927_),
    .A2(_02649_),
    .A1(net4071));
 sg13g2_o21ai_1 _09449_ (.B1(_02904_),
    .Y(_00653_),
    .A1(net3741),
    .A2(_02927_));
 sg13g2_nand2_1 _09450_ (.Y(_02928_),
    .A(net468),
    .B(net3743));
 sg13g2_nand2b_1 _09451_ (.Y(_02929_),
    .B(net4424),
    .A_N(\cpu.keccak_alu.registers[19] ));
 sg13g2_o21ai_1 _09452_ (.B1(_02929_),
    .Y(_02930_),
    .A1(net4424),
    .A2(\cpu.keccak_alu.registers[3] ));
 sg13g2_a221oi_1 _09453_ (.B2(\cpu.keccak_alu.registers[35] ),
    .C1(net4438),
    .B1(net4108),
    .A1(\cpu.keccak_alu.registers[51] ),
    .Y(_02931_),
    .A2(net4121));
 sg13g2_o21ai_1 _09454_ (.B1(_02931_),
    .Y(_02932_),
    .A1(net4401),
    .A2(_02930_));
 sg13g2_nand2_1 _09455_ (.Y(_02933_),
    .A(net4424),
    .B(_01018_));
 sg13g2_o21ai_1 _09456_ (.B1(_02933_),
    .Y(_02934_),
    .A1(net4425),
    .A2(\cpu.keccak_alu.registers[67] ));
 sg13g2_a22oi_1 _09457_ (.Y(_02935_),
    .B1(net4106),
    .B2(\cpu.keccak_alu.registers[99] ),
    .A2(net4119),
    .A1(\cpu.keccak_alu.registers[115] ));
 sg13g2_o21ai_1 _09458_ (.B1(_02935_),
    .Y(_02936_),
    .A1(net4401),
    .A2(_02934_));
 sg13g2_nand2b_1 _09459_ (.Y(_02937_),
    .B(net4424),
    .A_N(\cpu.keccak_alu.registers[211] ));
 sg13g2_o21ai_1 _09460_ (.B1(_02937_),
    .Y(_02938_),
    .A1(net4428),
    .A2(\cpu.keccak_alu.registers[195] ));
 sg13g2_a22oi_1 _09461_ (.Y(_02939_),
    .B1(net4106),
    .B2(\cpu.keccak_alu.registers[227] ),
    .A2(net4119),
    .A1(\cpu.keccak_alu.registers[243] ));
 sg13g2_o21ai_1 _09462_ (.B1(_02939_),
    .Y(_02940_),
    .A1(net4400),
    .A2(_02938_));
 sg13g2_nand2b_1 _09463_ (.Y(_02941_),
    .B(net4425),
    .A_N(\cpu.keccak_alu.registers[147] ));
 sg13g2_o21ai_1 _09464_ (.B1(_02941_),
    .Y(_02942_),
    .A1(net4425),
    .A2(net4530));
 sg13g2_a22oi_1 _09465_ (.Y(_02943_),
    .B1(net4106),
    .B2(net4495),
    .A2(net4119),
    .A1(\cpu.keccak_alu.registers[179] ));
 sg13g2_o21ai_1 _09466_ (.B1(_02943_),
    .Y(_02944_),
    .A1(net4401),
    .A2(_02942_));
 sg13g2_a22oi_1 _09467_ (.Y(_02945_),
    .B1(_02944_),
    .B2(net4129),
    .A2(_02940_),
    .A1(net4133));
 sg13g2_a22oi_1 _09468_ (.Y(_02946_),
    .B1(_02936_),
    .B2(net4131),
    .A2(_02932_),
    .A1(net4127));
 sg13g2_mux2_1 _09469_ (.A0(_01022_),
    .A1(_01023_),
    .S(net4424),
    .X(_02947_));
 sg13g2_a22oi_1 _09470_ (.Y(_02948_),
    .B1(net4106),
    .B2(\cpu.keccak_alu.registers[291] ),
    .A2(net4119),
    .A1(\cpu.keccak_alu.registers[307] ));
 sg13g2_o21ai_1 _09471_ (.B1(_02948_),
    .Y(_02949_),
    .A1(net4400),
    .A2(_02947_));
 sg13g2_nand2_1 _09472_ (.Y(_02950_),
    .A(net4126),
    .B(_02949_));
 sg13g2_a221oi_1 _09473_ (.B2(net4437),
    .C1(net3847),
    .B1(_02950_),
    .A1(_02945_),
    .Y(_02951_),
    .A2(_02946_));
 sg13g2_a21oi_2 _09474_ (.B1(_02951_),
    .Y(_02952_),
    .A2(_02656_),
    .A1(net4072));
 sg13g2_o21ai_1 _09475_ (.B1(_02928_),
    .Y(_00654_),
    .A1(net3741),
    .A2(_02952_));
 sg13g2_nand2_1 _09476_ (.Y(_02953_),
    .A(net97),
    .B(net3742));
 sg13g2_nand2b_1 _09477_ (.Y(_02954_),
    .B(net4421),
    .A_N(\cpu.keccak_alu.registers[20] ));
 sg13g2_o21ai_1 _09478_ (.B1(_02954_),
    .Y(_02955_),
    .A1(net4421),
    .A2(\cpu.keccak_alu.registers[4] ));
 sg13g2_a221oi_1 _09479_ (.B2(\cpu.keccak_alu.registers[36] ),
    .C1(net4437),
    .B1(net4104),
    .A1(\cpu.keccak_alu.registers[52] ),
    .Y(_02956_),
    .A2(net4117));
 sg13g2_o21ai_1 _09480_ (.B1(_02956_),
    .Y(_02957_),
    .A1(net4398),
    .A2(_02955_));
 sg13g2_nand2_1 _09481_ (.Y(_02958_),
    .A(net4419),
    .B(_01027_));
 sg13g2_o21ai_1 _09482_ (.B1(_02958_),
    .Y(_02959_),
    .A1(net4422),
    .A2(\cpu.keccak_alu.registers[68] ));
 sg13g2_a22oi_1 _09483_ (.Y(_02960_),
    .B1(net4107),
    .B2(\cpu.keccak_alu.registers[100] ),
    .A2(net4120),
    .A1(\cpu.keccak_alu.registers[116] ));
 sg13g2_o21ai_1 _09484_ (.B1(_02960_),
    .Y(_02961_),
    .A1(net4398),
    .A2(_02959_));
 sg13g2_nand2b_1 _09485_ (.Y(_02962_),
    .B(net4421),
    .A_N(\cpu.keccak_alu.registers[212] ));
 sg13g2_o21ai_1 _09486_ (.B1(_02962_),
    .Y(_02963_),
    .A1(net4421),
    .A2(\cpu.keccak_alu.registers[196] ));
 sg13g2_a22oi_1 _09487_ (.Y(_02964_),
    .B1(net4104),
    .B2(\cpu.keccak_alu.registers[228] ),
    .A2(net4117),
    .A1(\cpu.keccak_alu.registers[244] ));
 sg13g2_o21ai_1 _09488_ (.B1(_02964_),
    .Y(_02965_),
    .A1(net4397),
    .A2(_02963_));
 sg13g2_a22oi_1 _09489_ (.Y(_02966_),
    .B1(_02965_),
    .B2(net4133),
    .A2(_02961_),
    .A1(net4131));
 sg13g2_nand2b_1 _09490_ (.Y(_02967_),
    .B(net4421),
    .A_N(\cpu.keccak_alu.registers[148] ));
 sg13g2_o21ai_1 _09491_ (.B1(_02967_),
    .Y(_02968_),
    .A1(net4422),
    .A2(net4521));
 sg13g2_a22oi_1 _09492_ (.Y(_02969_),
    .B1(net4104),
    .B2(\cpu.keccak_alu.registers[164] ),
    .A2(net4117),
    .A1(\cpu.keccak_alu.registers[180] ));
 sg13g2_o21ai_1 _09493_ (.B1(_02969_),
    .Y(_02970_),
    .A1(net4397),
    .A2(_02968_));
 sg13g2_a22oi_1 _09494_ (.Y(_02971_),
    .B1(_02970_),
    .B2(net4129),
    .A2(_02957_),
    .A1(net4126));
 sg13g2_mux2_1 _09495_ (.A0(_01030_),
    .A1(_01031_),
    .S(net4421),
    .X(_02972_));
 sg13g2_a22oi_1 _09496_ (.Y(_02973_),
    .B1(net4104),
    .B2(\cpu.keccak_alu.registers[292] ),
    .A2(net4117),
    .A1(\cpu.keccak_alu.registers[308] ));
 sg13g2_o21ai_1 _09497_ (.B1(_02973_),
    .Y(_02974_),
    .A1(net4397),
    .A2(_02972_));
 sg13g2_nand2_1 _09498_ (.Y(_02975_),
    .A(net4126),
    .B(_02974_));
 sg13g2_a221oi_1 _09499_ (.B2(net4437),
    .C1(net3847),
    .B1(_02975_),
    .A1(_02966_),
    .Y(_02976_),
    .A2(_02971_));
 sg13g2_a21oi_2 _09500_ (.B1(_02976_),
    .Y(_02977_),
    .A2(_02663_),
    .A1(net4073));
 sg13g2_o21ai_1 _09501_ (.B1(_02953_),
    .Y(_00655_),
    .A1(net3740),
    .A2(_02977_));
 sg13g2_nand2_1 _09502_ (.Y(_02978_),
    .A(net72),
    .B(net3742));
 sg13g2_nand2b_1 _09503_ (.Y(_02979_),
    .B(net4420),
    .A_N(\cpu.keccak_alu.registers[21] ));
 sg13g2_o21ai_1 _09504_ (.B1(_02979_),
    .Y(_02980_),
    .A1(net4420),
    .A2(\cpu.keccak_alu.registers[5] ));
 sg13g2_a221oi_1 _09505_ (.B2(\cpu.keccak_alu.registers[37] ),
    .C1(net4437),
    .B1(net4105),
    .A1(\cpu.keccak_alu.registers[53] ),
    .Y(_02981_),
    .A2(net4118));
 sg13g2_o21ai_1 _09506_ (.B1(_02981_),
    .Y(_02982_),
    .A1(net4398),
    .A2(_02980_));
 sg13g2_nand2b_1 _09507_ (.Y(_02983_),
    .B(net4420),
    .A_N(\cpu.keccak_alu.registers[85] ));
 sg13g2_o21ai_1 _09508_ (.B1(_02983_),
    .Y(_02984_),
    .A1(net4420),
    .A2(\cpu.keccak_alu.registers[69] ));
 sg13g2_a22oi_1 _09509_ (.Y(_02985_),
    .B1(net4105),
    .B2(\cpu.keccak_alu.registers[101] ),
    .A2(net4118),
    .A1(\cpu.keccak_alu.registers[117] ));
 sg13g2_o21ai_1 _09510_ (.B1(_02985_),
    .Y(_02986_),
    .A1(net4398),
    .A2(_02984_));
 sg13g2_nand2b_1 _09511_ (.Y(_02987_),
    .B(net4420),
    .A_N(\cpu.keccak_alu.registers[213] ));
 sg13g2_o21ai_1 _09512_ (.B1(_02987_),
    .Y(_02988_),
    .A1(net4420),
    .A2(\cpu.keccak_alu.registers[197] ));
 sg13g2_a22oi_1 _09513_ (.Y(_02989_),
    .B1(net4102),
    .B2(\cpu.keccak_alu.registers[229] ),
    .A2(net4115),
    .A1(\cpu.keccak_alu.registers[245] ));
 sg13g2_o21ai_1 _09514_ (.B1(_02989_),
    .Y(_02990_),
    .A1(net4398),
    .A2(_02988_));
 sg13g2_mux2_1 _09515_ (.A0(net4161),
    .A1(_01037_),
    .S(net4420),
    .X(_02991_));
 sg13g2_a22oi_1 _09516_ (.Y(_02992_),
    .B1(net4105),
    .B2(\cpu.keccak_alu.registers[165] ),
    .A2(net4118),
    .A1(net4486));
 sg13g2_o21ai_1 _09517_ (.B1(_02992_),
    .Y(_02993_),
    .A1(net4398),
    .A2(_02991_));
 sg13g2_a22oi_1 _09518_ (.Y(_02994_),
    .B1(_02990_),
    .B2(net4133),
    .A2(_02986_),
    .A1(net4131));
 sg13g2_a22oi_1 _09519_ (.Y(_02995_),
    .B1(_02993_),
    .B2(net4129),
    .A2(_02982_),
    .A1(net4126));
 sg13g2_a21oi_1 _09520_ (.A1(net4421),
    .A2(_01039_),
    .Y(_02996_),
    .B1(net4398));
 sg13g2_o21ai_1 _09521_ (.B1(_02996_),
    .Y(_02997_),
    .A1(net4421),
    .A2(\cpu.keccak_alu.registers[261] ));
 sg13g2_a22oi_1 _09522_ (.Y(_02998_),
    .B1(net4105),
    .B2(\cpu.keccak_alu.registers[293] ),
    .A2(net4118),
    .A1(\cpu.keccak_alu.registers[309] ));
 sg13g2_a21o_1 _09523_ (.A2(_02998_),
    .A1(_02997_),
    .B1(net4124),
    .X(_02999_));
 sg13g2_a221oi_1 _09524_ (.B2(net4437),
    .C1(net3847),
    .B1(_02999_),
    .A1(_02994_),
    .Y(_03000_),
    .A2(_02995_));
 sg13g2_a21oi_2 _09525_ (.B1(_03000_),
    .Y(_03001_),
    .A2(_02670_),
    .A1(net4073));
 sg13g2_o21ai_1 _09526_ (.B1(_02978_),
    .Y(_00656_),
    .A1(net3740),
    .A2(_03001_));
 sg13g2_nand2_1 _09527_ (.Y(_03002_),
    .A(net186),
    .B(net3742));
 sg13g2_a21oi_1 _09528_ (.A1(net4419),
    .A2(_01042_),
    .Y(_03003_),
    .B1(net4397));
 sg13g2_o21ai_1 _09529_ (.B1(_03003_),
    .Y(_03004_),
    .A1(net4419),
    .A2(\cpu.keccak_alu.registers[6] ));
 sg13g2_a22oi_1 _09530_ (.Y(_03005_),
    .B1(net4104),
    .B2(\cpu.keccak_alu.registers[38] ),
    .A2(net4117),
    .A1(\cpu.keccak_alu.registers[54] ));
 sg13g2_nand3_1 _09531_ (.B(_03004_),
    .C(_03005_),
    .A(net4201),
    .Y(_03006_));
 sg13g2_nand2b_1 _09532_ (.Y(_03007_),
    .B(net4419),
    .A_N(\cpu.keccak_alu.registers[86] ));
 sg13g2_o21ai_1 _09533_ (.B1(_03007_),
    .Y(_03008_),
    .A1(net4419),
    .A2(\cpu.keccak_alu.registers[70] ));
 sg13g2_a22oi_1 _09534_ (.Y(_03009_),
    .B1(net4104),
    .B2(\cpu.keccak_alu.registers[102] ),
    .A2(net4117),
    .A1(\cpu.keccak_alu.registers[118] ));
 sg13g2_o21ai_1 _09535_ (.B1(_03009_),
    .Y(_03010_),
    .A1(net4397),
    .A2(_03008_));
 sg13g2_nand2b_1 _09536_ (.Y(_03011_),
    .B(net4419),
    .A_N(\cpu.keccak_alu.registers[214] ));
 sg13g2_o21ai_1 _09537_ (.B1(_03011_),
    .Y(_03012_),
    .A1(net4419),
    .A2(\cpu.keccak_alu.registers[198] ));
 sg13g2_a22oi_1 _09538_ (.Y(_03013_),
    .B1(net4105),
    .B2(\cpu.keccak_alu.registers[230] ),
    .A2(net4118),
    .A1(\cpu.keccak_alu.registers[246] ));
 sg13g2_o21ai_1 _09539_ (.B1(_03013_),
    .Y(_03014_),
    .A1(net4397),
    .A2(_03012_));
 sg13g2_a22oi_1 _09540_ (.Y(_03015_),
    .B1(_03014_),
    .B2(net4133),
    .A2(_03010_),
    .A1(net4131));
 sg13g2_mux2_1 _09541_ (.A0(net4158),
    .A1(_01047_),
    .S(net4420),
    .X(_03016_));
 sg13g2_a22oi_1 _09542_ (.Y(_03017_),
    .B1(net4104),
    .B2(\cpu.keccak_alu.registers[166] ),
    .A2(net4117),
    .A1(net4485));
 sg13g2_o21ai_1 _09543_ (.B1(_03017_),
    .Y(_03018_),
    .A1(net4397),
    .A2(_03016_));
 sg13g2_a22oi_1 _09544_ (.Y(_03019_),
    .B1(_03018_),
    .B2(net4129),
    .A2(_03006_),
    .A1(net4126));
 sg13g2_mux2_1 _09545_ (.A0(_01048_),
    .A1(_01049_),
    .S(net4419),
    .X(_03020_));
 sg13g2_a22oi_1 _09546_ (.Y(_03021_),
    .B1(net4104),
    .B2(\cpu.keccak_alu.registers[294] ),
    .A2(net4117),
    .A1(\cpu.keccak_alu.registers[310] ));
 sg13g2_o21ai_1 _09547_ (.B1(_03021_),
    .Y(_03022_),
    .A1(net4397),
    .A2(_03020_));
 sg13g2_nand2_1 _09548_ (.Y(_03023_),
    .A(net4126),
    .B(_03022_));
 sg13g2_a221oi_1 _09549_ (.B2(net4437),
    .C1(net3847),
    .B1(_03023_),
    .A1(_03015_),
    .Y(_03024_),
    .A2(_03019_));
 sg13g2_a21oi_2 _09550_ (.B1(_03024_),
    .Y(_03025_),
    .A2(_02678_),
    .A1(net4072));
 sg13g2_o21ai_1 _09551_ (.B1(_03002_),
    .Y(_00657_),
    .A1(net3740),
    .A2(_03025_));
 sg13g2_nand2_1 _09552_ (.Y(_03026_),
    .A(net306),
    .B(_02876_));
 sg13g2_nand2b_1 _09553_ (.Y(_03027_),
    .B(net4415),
    .A_N(\cpu.keccak_alu.registers[23] ));
 sg13g2_o21ai_1 _09554_ (.B1(_03027_),
    .Y(_03028_),
    .A1(net4415),
    .A2(\cpu.keccak_alu.registers[7] ));
 sg13g2_a221oi_1 _09555_ (.B2(\cpu.keccak_alu.registers[39] ),
    .C1(net4436),
    .B1(net4103),
    .A1(\cpu.keccak_alu.registers[55] ),
    .Y(_03029_),
    .A2(net4115));
 sg13g2_o21ai_1 _09556_ (.B1(_03029_),
    .Y(_03030_),
    .A1(net4394),
    .A2(_03028_));
 sg13g2_nand2b_1 _09557_ (.Y(_03031_),
    .B(net4415),
    .A_N(\cpu.keccak_alu.registers[215] ));
 sg13g2_o21ai_1 _09558_ (.B1(_03031_),
    .Y(_03032_),
    .A1(net4415),
    .A2(\cpu.keccak_alu.registers[199] ));
 sg13g2_a22oi_1 _09559_ (.Y(_03033_),
    .B1(net4103),
    .B2(\cpu.keccak_alu.registers[231] ),
    .A2(net4115),
    .A1(\cpu.keccak_alu.registers[247] ));
 sg13g2_o21ai_1 _09560_ (.B1(_03033_),
    .Y(_03034_),
    .A1(net4394),
    .A2(_03032_));
 sg13g2_nand2_1 _09561_ (.Y(_03035_),
    .A(net4417),
    .B(_01052_));
 sg13g2_o21ai_1 _09562_ (.B1(_03035_),
    .Y(_03036_),
    .A1(net4417),
    .A2(\cpu.keccak_alu.registers[71] ));
 sg13g2_a22oi_1 _09563_ (.Y(_03037_),
    .B1(net4103),
    .B2(\cpu.keccak_alu.registers[103] ),
    .A2(net4115),
    .A1(\cpu.keccak_alu.registers[119] ));
 sg13g2_o21ai_1 _09564_ (.B1(_03037_),
    .Y(_03038_),
    .A1(net4393),
    .A2(_03036_));
 sg13g2_nand2b_1 _09565_ (.Y(_03039_),
    .B(net4415),
    .A_N(\cpu.keccak_alu.registers[151] ));
 sg13g2_o21ai_1 _09566_ (.B1(_03039_),
    .Y(_03040_),
    .A1(net4415),
    .A2(net4512));
 sg13g2_a22oi_1 _09567_ (.Y(_03041_),
    .B1(net4103),
    .B2(\cpu.keccak_alu.registers[167] ),
    .A2(net4122),
    .A1(\cpu.keccak_alu.registers[183] ));
 sg13g2_o21ai_1 _09568_ (.B1(_03041_),
    .Y(_03042_),
    .A1(net4394),
    .A2(_03040_));
 sg13g2_a22oi_1 _09569_ (.Y(_03043_),
    .B1(_03038_),
    .B2(net4130),
    .A2(_03034_),
    .A1(net4132));
 sg13g2_a22oi_1 _09570_ (.Y(_03044_),
    .B1(_03042_),
    .B2(net4128),
    .A2(_03030_),
    .A1(net4125));
 sg13g2_a21oi_1 _09571_ (.A1(net4415),
    .A2(_01058_),
    .Y(_03045_),
    .B1(net4395));
 sg13g2_o21ai_1 _09572_ (.B1(_03045_),
    .Y(_03046_),
    .A1(net4415),
    .A2(\cpu.keccak_alu.registers[263] ));
 sg13g2_a22oi_1 _09573_ (.Y(_03047_),
    .B1(net4103),
    .B2(\cpu.keccak_alu.registers[295] ),
    .A2(net4115),
    .A1(\cpu.keccak_alu.registers[311] ));
 sg13g2_a21o_1 _09574_ (.A2(_03047_),
    .A1(_03046_),
    .B1(net4124),
    .X(_03048_));
 sg13g2_a221oi_1 _09575_ (.B2(net4436),
    .C1(net3846),
    .B1(_03048_),
    .A1(_03043_),
    .Y(_03049_),
    .A2(_03044_));
 sg13g2_a21oi_2 _09576_ (.B1(_03049_),
    .Y(_03050_),
    .A2(_02685_),
    .A1(net4070));
 sg13g2_o21ai_1 _09577_ (.B1(_03026_),
    .Y(_00658_),
    .A1(net3741),
    .A2(_03050_));
 sg13g2_nand2_1 _09578_ (.Y(_03051_),
    .A(net216),
    .B(net3743));
 sg13g2_nand2b_1 _09579_ (.Y(_03052_),
    .B(net4413),
    .A_N(\cpu.keccak_alu.registers[24] ));
 sg13g2_o21ai_1 _09580_ (.B1(_03052_),
    .Y(_03053_),
    .A1(net4413),
    .A2(\cpu.keccak_alu.registers[8] ));
 sg13g2_a221oi_1 _09581_ (.B2(\cpu.keccak_alu.registers[40] ),
    .C1(net4436),
    .B1(net4099),
    .A1(\cpu.keccak_alu.registers[56] ),
    .Y(_03054_),
    .A2(net4112));
 sg13g2_o21ai_1 _09582_ (.B1(_03054_),
    .Y(_03055_),
    .A1(net4393),
    .A2(_03053_));
 sg13g2_nand2b_1 _09583_ (.Y(_03056_),
    .B(net4413),
    .A_N(\cpu.keccak_alu.registers[216] ));
 sg13g2_o21ai_1 _09584_ (.B1(_03056_),
    .Y(_03057_),
    .A1(net4413),
    .A2(\cpu.keccak_alu.registers[200] ));
 sg13g2_a22oi_1 _09585_ (.Y(_03058_),
    .B1(net4099),
    .B2(\cpu.keccak_alu.registers[232] ),
    .A2(net4112),
    .A1(\cpu.keccak_alu.registers[248] ));
 sg13g2_o21ai_1 _09586_ (.B1(_03058_),
    .Y(_03059_),
    .A1(net4393),
    .A2(_03057_));
 sg13g2_mux2_1 _09587_ (.A0(_01062_),
    .A1(_01063_),
    .S(net4413),
    .X(_03060_));
 sg13g2_a22oi_1 _09588_ (.Y(_03061_),
    .B1(net4102),
    .B2(\cpu.keccak_alu.registers[104] ),
    .A2(net4116),
    .A1(\cpu.keccak_alu.registers[120] ));
 sg13g2_o21ai_1 _09589_ (.B1(_03061_),
    .Y(_03062_),
    .A1(net4393),
    .A2(_03060_));
 sg13g2_a22oi_1 _09590_ (.Y(_03063_),
    .B1(_03062_),
    .B2(net4130),
    .A2(_03059_),
    .A1(net4133));
 sg13g2_nand2b_1 _09591_ (.Y(_03064_),
    .B(net4413),
    .A_N(\cpu.keccak_alu.registers[152] ));
 sg13g2_o21ai_1 _09592_ (.B1(_03064_),
    .Y(_03065_),
    .A1(net4413),
    .A2(net4511));
 sg13g2_a22oi_1 _09593_ (.Y(_03066_),
    .B1(net4102),
    .B2(\cpu.keccak_alu.registers[168] ),
    .A2(net4116),
    .A1(\cpu.keccak_alu.registers[184] ));
 sg13g2_o21ai_1 _09594_ (.B1(_03066_),
    .Y(_03067_),
    .A1(net4393),
    .A2(_03065_));
 sg13g2_a22oi_1 _09595_ (.Y(_03068_),
    .B1(_03067_),
    .B2(net4129),
    .A2(_03055_),
    .A1(net4127));
 sg13g2_a21oi_1 _09596_ (.A1(net4413),
    .A2(_01067_),
    .Y(_03069_),
    .B1(net4393));
 sg13g2_o21ai_1 _09597_ (.B1(_03069_),
    .Y(_03070_),
    .A1(net4414),
    .A2(\cpu.keccak_alu.registers[264] ));
 sg13g2_a22oi_1 _09598_ (.Y(_03071_),
    .B1(net4099),
    .B2(\cpu.keccak_alu.registers[296] ),
    .A2(net4112),
    .A1(\cpu.keccak_alu.registers[312] ));
 sg13g2_a21o_1 _09599_ (.A2(_03071_),
    .A1(_03070_),
    .B1(net4124),
    .X(_03072_));
 sg13g2_a221oi_1 _09600_ (.B2(net4434),
    .C1(net3846),
    .B1(_03072_),
    .A1(_03063_),
    .Y(_03073_),
    .A2(_03068_));
 sg13g2_a21oi_2 _09601_ (.B1(_03073_),
    .Y(_03074_),
    .A2(_02692_),
    .A1(net4069));
 sg13g2_o21ai_1 _09602_ (.B1(_03051_),
    .Y(_00659_),
    .A1(net3741),
    .A2(_03074_));
 sg13g2_a21oi_1 _09603_ (.A1(net4403),
    .A2(_01070_),
    .Y(_03075_),
    .B1(net4388));
 sg13g2_o21ai_1 _09604_ (.B1(_03075_),
    .Y(_03076_),
    .A1(net4403),
    .A2(\cpu.keccak_alu.registers[9] ));
 sg13g2_a221oi_1 _09605_ (.B2(\cpu.keccak_alu.registers[41] ),
    .C1(net4434),
    .B1(net4097),
    .A1(\cpu.keccak_alu.registers[57] ),
    .Y(_03077_),
    .A2(net4110));
 sg13g2_a21oi_1 _09606_ (.A1(_03076_),
    .A2(_03077_),
    .Y(_03078_),
    .B1(net4123));
 sg13g2_nand2b_1 _09607_ (.Y(_03079_),
    .B(net4403),
    .A_N(net4500));
 sg13g2_o21ai_1 _09608_ (.B1(_03079_),
    .Y(_03080_),
    .A1(net4406),
    .A2(net4509));
 sg13g2_a22oi_1 _09609_ (.Y(_03081_),
    .B1(net4097),
    .B2(\cpu.keccak_alu.registers[169] ),
    .A2(net4110),
    .A1(\cpu.keccak_alu.registers[185] ));
 sg13g2_o21ai_1 _09610_ (.B1(_03081_),
    .Y(_03082_),
    .A1(net4388),
    .A2(_03080_));
 sg13g2_mux2_1 _09611_ (.A0(_01072_),
    .A1(_01073_),
    .S(net4403),
    .X(_03083_));
 sg13g2_a22oi_1 _09612_ (.Y(_03084_),
    .B1(net4097),
    .B2(\cpu.keccak_alu.registers[105] ),
    .A2(net4110),
    .A1(\cpu.keccak_alu.registers[121] ));
 sg13g2_o21ai_1 _09613_ (.B1(_03084_),
    .Y(_03085_),
    .A1(net4388),
    .A2(_03083_));
 sg13g2_nand2_1 _09614_ (.Y(_03086_),
    .A(net4130),
    .B(_03085_));
 sg13g2_nand2b_1 _09615_ (.Y(_03087_),
    .B(net4403),
    .A_N(\cpu.keccak_alu.registers[217] ));
 sg13g2_o21ai_1 _09616_ (.B1(_03087_),
    .Y(_03088_),
    .A1(net4403),
    .A2(\cpu.keccak_alu.registers[201] ));
 sg13g2_a22oi_1 _09617_ (.Y(_03089_),
    .B1(net4097),
    .B2(\cpu.keccak_alu.registers[233] ),
    .A2(net4110),
    .A1(\cpu.keccak_alu.registers[249] ));
 sg13g2_o21ai_1 _09618_ (.B1(_03089_),
    .Y(_03090_),
    .A1(net4389),
    .A2(_03088_));
 sg13g2_a221oi_1 _09619_ (.B2(net4132),
    .C1(_03078_),
    .B1(_03090_),
    .A1(net4128),
    .Y(_03091_),
    .A2(_03082_));
 sg13g2_a21oi_1 _09620_ (.A1(net4404),
    .A2(_01075_),
    .Y(_03092_),
    .B1(net4388));
 sg13g2_o21ai_1 _09621_ (.B1(_03092_),
    .Y(_03093_),
    .A1(net4403),
    .A2(\cpu.keccak_alu.registers[265] ));
 sg13g2_a22oi_1 _09622_ (.Y(_03094_),
    .B1(net4097),
    .B2(\cpu.keccak_alu.registers[297] ),
    .A2(net4110),
    .A1(\cpu.keccak_alu.registers[313] ));
 sg13g2_a21o_1 _09623_ (.A2(_03094_),
    .A1(_03093_),
    .B1(net4123),
    .X(_03095_));
 sg13g2_a221oi_1 _09624_ (.B2(net4434),
    .C1(net3846),
    .B1(_03095_),
    .A1(_03086_),
    .Y(_03096_),
    .A2(_03091_));
 sg13g2_a21oi_1 _09625_ (.A1(net4068),
    .A2(_02698_),
    .Y(_03097_),
    .B1(_03096_));
 sg13g2_nand2_1 _09626_ (.Y(_03098_),
    .A(net110),
    .B(net3742));
 sg13g2_o21ai_1 _09627_ (.B1(_03098_),
    .Y(_00660_),
    .A1(net3740),
    .A2(_03097_));
 sg13g2_nand2_1 _09628_ (.Y(_03099_),
    .A(net74),
    .B(net3742));
 sg13g2_nand2b_1 _09629_ (.Y(_03100_),
    .B(net4404),
    .A_N(\cpu.keccak_alu.registers[26] ));
 sg13g2_o21ai_1 _09630_ (.B1(_03100_),
    .Y(_03101_),
    .A1(net4404),
    .A2(\cpu.keccak_alu.registers[10] ));
 sg13g2_a221oi_1 _09631_ (.B2(\cpu.keccak_alu.registers[42] ),
    .C1(net4434),
    .B1(net4098),
    .A1(\cpu.keccak_alu.registers[58] ),
    .Y(_03102_),
    .A2(net4111));
 sg13g2_o21ai_1 _09632_ (.B1(_03102_),
    .Y(_03103_),
    .A1(net4388),
    .A2(_03101_));
 sg13g2_mux2_1 _09633_ (.A0(_01078_),
    .A1(_01079_),
    .S(net4406),
    .X(_03104_));
 sg13g2_a22oi_1 _09634_ (.Y(_03105_),
    .B1(net4097),
    .B2(\cpu.keccak_alu.registers[106] ),
    .A2(net4110),
    .A1(\cpu.keccak_alu.registers[122] ));
 sg13g2_o21ai_1 _09635_ (.B1(_03105_),
    .Y(_03106_),
    .A1(net4388),
    .A2(_03104_));
 sg13g2_nand2b_1 _09636_ (.Y(_03107_),
    .B(net4404),
    .A_N(\cpu.keccak_alu.registers[218] ));
 sg13g2_o21ai_1 _09637_ (.B1(_03107_),
    .Y(_03108_),
    .A1(net4403),
    .A2(\cpu.keccak_alu.registers[202] ));
 sg13g2_a22oi_1 _09638_ (.Y(_03109_),
    .B1(net4097),
    .B2(\cpu.keccak_alu.registers[234] ),
    .A2(net4110),
    .A1(\cpu.keccak_alu.registers[250] ));
 sg13g2_o21ai_1 _09639_ (.B1(_03109_),
    .Y(_03110_),
    .A1(net4389),
    .A2(_03108_));
 sg13g2_nand2b_1 _09640_ (.Y(_03111_),
    .B(net4407),
    .A_N(\cpu.keccak_alu.registers[154] ));
 sg13g2_o21ai_1 _09641_ (.B1(_03111_),
    .Y(_03112_),
    .A1(net4407),
    .A2(\cpu.keccak_alu.registers[138] ));
 sg13g2_a22oi_1 _09642_ (.Y(_03113_),
    .B1(net4097),
    .B2(net4492),
    .A2(net4110),
    .A1(\cpu.keccak_alu.registers[186] ));
 sg13g2_o21ai_1 _09643_ (.B1(_03113_),
    .Y(_03114_),
    .A1(net4388),
    .A2(_03112_));
 sg13g2_a22oi_1 _09644_ (.Y(_03115_),
    .B1(_03114_),
    .B2(net4128),
    .A2(_03110_),
    .A1(net4132));
 sg13g2_a22oi_1 _09645_ (.Y(_03116_),
    .B1(_03106_),
    .B2(net4130),
    .A2(_03103_),
    .A1(net4125));
 sg13g2_a21oi_1 _09646_ (.A1(net4405),
    .A2(_01082_),
    .Y(_03117_),
    .B1(net4389));
 sg13g2_o21ai_1 _09647_ (.B1(_03117_),
    .Y(_03118_),
    .A1(net4404),
    .A2(\cpu.keccak_alu.registers[266] ));
 sg13g2_a22oi_1 _09648_ (.Y(_03119_),
    .B1(net4098),
    .B2(\cpu.keccak_alu.registers[298] ),
    .A2(net4111),
    .A1(\cpu.keccak_alu.registers[314] ));
 sg13g2_a21o_1 _09649_ (.A2(_03119_),
    .A1(_03118_),
    .B1(net4123),
    .X(_03120_));
 sg13g2_a221oi_1 _09650_ (.B2(net4434),
    .C1(net3846),
    .B1(_03120_),
    .A1(_03115_),
    .Y(_03121_),
    .A2(_03116_));
 sg13g2_a21oi_1 _09651_ (.A1(net4068),
    .A2(_02704_),
    .Y(_03122_),
    .B1(_03121_));
 sg13g2_o21ai_1 _09652_ (.B1(_03099_),
    .Y(_00661_),
    .A1(net3740),
    .A2(_03122_));
 sg13g2_nand2_1 _09653_ (.Y(_03123_),
    .A(net87),
    .B(net3743));
 sg13g2_a21oi_1 _09654_ (.A1(net4409),
    .A2(_01085_),
    .Y(_03124_),
    .B1(net4390));
 sg13g2_o21ai_1 _09655_ (.B1(_03124_),
    .Y(_03125_),
    .A1(net4409),
    .A2(\cpu.keccak_alu.registers[11] ));
 sg13g2_a22oi_1 _09656_ (.Y(_03126_),
    .B1(net4099),
    .B2(\cpu.keccak_alu.registers[43] ),
    .A2(net4112),
    .A1(\cpu.keccak_alu.registers[59] ));
 sg13g2_nand3_1 _09657_ (.B(_03125_),
    .C(_03126_),
    .A(net4201),
    .Y(_03127_));
 sg13g2_nand2b_1 _09658_ (.Y(_03128_),
    .B(net4409),
    .A_N(\cpu.keccak_alu.registers[219] ));
 sg13g2_o21ai_1 _09659_ (.B1(_03128_),
    .Y(_03129_),
    .A1(net4409),
    .A2(\cpu.keccak_alu.registers[203] ));
 sg13g2_a22oi_1 _09660_ (.Y(_03130_),
    .B1(net4101),
    .B2(\cpu.keccak_alu.registers[235] ),
    .A2(net4114),
    .A1(\cpu.keccak_alu.registers[251] ));
 sg13g2_o21ai_1 _09661_ (.B1(_03130_),
    .Y(_03131_),
    .A1(net4390),
    .A2(_03129_));
 sg13g2_nand2b_1 _09662_ (.Y(_03132_),
    .B(net4410),
    .A_N(\cpu.keccak_alu.registers[91] ));
 sg13g2_o21ai_1 _09663_ (.B1(_03132_),
    .Y(_03133_),
    .A1(net4409),
    .A2(\cpu.keccak_alu.registers[75] ));
 sg13g2_a22oi_1 _09664_ (.Y(_03134_),
    .B1(net4099),
    .B2(\cpu.keccak_alu.registers[107] ),
    .A2(net4112),
    .A1(\cpu.keccak_alu.registers[123] ));
 sg13g2_o21ai_1 _09665_ (.B1(_03134_),
    .Y(_03135_),
    .A1(net4390),
    .A2(_03133_));
 sg13g2_nand2b_1 _09666_ (.Y(_03136_),
    .B(net4410),
    .A_N(\cpu.keccak_alu.registers[155] ));
 sg13g2_o21ai_1 _09667_ (.B1(_03136_),
    .Y(_03137_),
    .A1(net4410),
    .A2(\cpu.keccak_alu.registers[139] ));
 sg13g2_a22oi_1 _09668_ (.Y(_03138_),
    .B1(net4099),
    .B2(net4490),
    .A2(net4112),
    .A1(net4484));
 sg13g2_o21ai_1 _09669_ (.B1(_03138_),
    .Y(_03139_),
    .A1(net4390),
    .A2(_03137_));
 sg13g2_a22oi_1 _09670_ (.Y(_03140_),
    .B1(_03139_),
    .B2(net4128),
    .A2(_03135_),
    .A1(net4130));
 sg13g2_a22oi_1 _09671_ (.Y(_03141_),
    .B1(_03131_),
    .B2(net4132),
    .A2(_03127_),
    .A1(net4125));
 sg13g2_a21oi_1 _09672_ (.A1(net4407),
    .A2(_01091_),
    .Y(_03142_),
    .B1(net4388));
 sg13g2_o21ai_1 _09673_ (.B1(_03142_),
    .Y(_03143_),
    .A1(net4409),
    .A2(\cpu.keccak_alu.registers[267] ));
 sg13g2_a22oi_1 _09674_ (.Y(_03144_),
    .B1(net4099),
    .B2(\cpu.keccak_alu.registers[299] ),
    .A2(net4112),
    .A1(\cpu.keccak_alu.registers[315] ));
 sg13g2_a21o_1 _09675_ (.A2(_03144_),
    .A1(_03143_),
    .B1(net4123),
    .X(_03145_));
 sg13g2_a221oi_1 _09676_ (.B2(net4434),
    .C1(net3846),
    .B1(_03145_),
    .A1(_03140_),
    .Y(_03146_),
    .A2(_03141_));
 sg13g2_a21oi_2 _09677_ (.B1(_03146_),
    .Y(_03147_),
    .A2(_02713_),
    .A1(net4068));
 sg13g2_o21ai_1 _09678_ (.B1(_03123_),
    .Y(_00662_),
    .A1(net3741),
    .A2(_03147_));
 sg13g2_nand2_1 _09679_ (.Y(_03148_),
    .A(net70),
    .B(net3742));
 sg13g2_a21oi_1 _09680_ (.A1(net4416),
    .A2(_01094_),
    .Y(_03149_),
    .B1(net4394));
 sg13g2_o21ai_1 _09681_ (.B1(_03149_),
    .Y(_03150_),
    .A1(net4416),
    .A2(\cpu.keccak_alu.registers[12] ));
 sg13g2_a22oi_1 _09682_ (.Y(_03151_),
    .B1(net4102),
    .B2(\cpu.keccak_alu.registers[44] ),
    .A2(net4116),
    .A1(\cpu.keccak_alu.registers[60] ));
 sg13g2_nand3_1 _09683_ (.B(_03150_),
    .C(_03151_),
    .A(net4201),
    .Y(_03152_));
 sg13g2_nand2b_1 _09684_ (.Y(_03153_),
    .B(net4414),
    .A_N(\cpu.keccak_alu.registers[220] ));
 sg13g2_o21ai_1 _09685_ (.B1(_03153_),
    .Y(_03154_),
    .A1(net4416),
    .A2(\cpu.keccak_alu.registers[204] ));
 sg13g2_a22oi_1 _09686_ (.Y(_03155_),
    .B1(net4102),
    .B2(\cpu.keccak_alu.registers[236] ),
    .A2(net4116),
    .A1(\cpu.keccak_alu.registers[252] ));
 sg13g2_o21ai_1 _09687_ (.B1(_03155_),
    .Y(_03156_),
    .A1(net4394),
    .A2(_03154_));
 sg13g2_nand2b_1 _09688_ (.Y(_03157_),
    .B(net4416),
    .A_N(\cpu.keccak_alu.registers[92] ));
 sg13g2_o21ai_1 _09689_ (.B1(_03157_),
    .Y(_03158_),
    .A1(net4416),
    .A2(\cpu.keccak_alu.registers[76] ));
 sg13g2_a22oi_1 _09690_ (.Y(_03159_),
    .B1(net4102),
    .B2(\cpu.keccak_alu.registers[108] ),
    .A2(net4116),
    .A1(\cpu.keccak_alu.registers[124] ));
 sg13g2_o21ai_1 _09691_ (.B1(_03159_),
    .Y(_03160_),
    .A1(net4393),
    .A2(_03158_));
 sg13g2_a22oi_1 _09692_ (.Y(_03161_),
    .B1(_03160_),
    .B2(net4131),
    .A2(_03156_),
    .A1(net4133));
 sg13g2_nand2_1 _09693_ (.Y(_03162_),
    .A(net4414),
    .B(_01097_));
 sg13g2_o21ai_1 _09694_ (.B1(_03162_),
    .Y(_03163_),
    .A1(net4414),
    .A2(net4507));
 sg13g2_a22oi_1 _09695_ (.Y(_03164_),
    .B1(net4102),
    .B2(net4489),
    .A2(net4116),
    .A1(\cpu.keccak_alu.registers[188] ));
 sg13g2_o21ai_1 _09696_ (.B1(_03164_),
    .Y(_03165_),
    .A1(net4393),
    .A2(_03163_));
 sg13g2_a22oi_1 _09697_ (.Y(_03166_),
    .B1(_03165_),
    .B2(net4129),
    .A2(_03152_),
    .A1(net4127));
 sg13g2_a21oi_1 _09698_ (.A1(net4416),
    .A2(_01100_),
    .Y(_03167_),
    .B1(net4394));
 sg13g2_o21ai_1 _09699_ (.B1(_03167_),
    .Y(_03168_),
    .A1(net4416),
    .A2(\cpu.keccak_alu.registers[268] ));
 sg13g2_a22oi_1 _09700_ (.Y(_03169_),
    .B1(net4102),
    .B2(\cpu.keccak_alu.registers[300] ),
    .A2(net4116),
    .A1(\cpu.keccak_alu.registers[316] ));
 sg13g2_a21o_1 _09701_ (.A2(_03169_),
    .A1(_03168_),
    .B1(net4124),
    .X(_03170_));
 sg13g2_a221oi_1 _09702_ (.B2(net4436),
    .C1(net3847),
    .B1(_03170_),
    .A1(_03161_),
    .Y(_03171_),
    .A2(_03166_));
 sg13g2_a21oi_2 _09703_ (.B1(_03171_),
    .Y(_03172_),
    .A2(_02718_),
    .A1(net4070));
 sg13g2_o21ai_1 _09704_ (.B1(_03148_),
    .Y(_00663_),
    .A1(net3740),
    .A2(_03172_));
 sg13g2_nand2_1 _09705_ (.Y(_03173_),
    .A(net105),
    .B(net3742));
 sg13g2_nand2b_1 _09706_ (.Y(_03174_),
    .B(net4408),
    .A_N(\cpu.keccak_alu.registers[29] ));
 sg13g2_o21ai_1 _09707_ (.B1(_03174_),
    .Y(_03175_),
    .A1(net4408),
    .A2(\cpu.keccak_alu.registers[13] ));
 sg13g2_a221oi_1 _09708_ (.B2(\cpu.keccak_alu.registers[45] ),
    .C1(net4435),
    .B1(net4100),
    .A1(\cpu.keccak_alu.registers[61] ),
    .Y(_03176_),
    .A2(net4113));
 sg13g2_o21ai_1 _09709_ (.B1(_03176_),
    .Y(_03177_),
    .A1(net4391),
    .A2(_03175_));
 sg13g2_mux2_1 _09710_ (.A0(_01103_),
    .A1(_01104_),
    .S(net4408),
    .X(_03178_));
 sg13g2_a22oi_1 _09711_ (.Y(_03179_),
    .B1(net4100),
    .B2(\cpu.keccak_alu.registers[109] ),
    .A2(net4113),
    .A1(\cpu.keccak_alu.registers[125] ));
 sg13g2_o21ai_1 _09712_ (.B1(_03179_),
    .Y(_03180_),
    .A1(net4391),
    .A2(_03178_));
 sg13g2_nand2b_1 _09713_ (.Y(_03181_),
    .B(net4408),
    .A_N(\cpu.keccak_alu.registers[221] ));
 sg13g2_o21ai_1 _09714_ (.B1(_03181_),
    .Y(_03182_),
    .A1(net4408),
    .A2(\cpu.keccak_alu.registers[205] ));
 sg13g2_a22oi_1 _09715_ (.Y(_03183_),
    .B1(net4100),
    .B2(\cpu.keccak_alu.registers[237] ),
    .A2(net4113),
    .A1(\cpu.keccak_alu.registers[253] ));
 sg13g2_o21ai_1 _09716_ (.B1(_03183_),
    .Y(_03184_),
    .A1(net4391),
    .A2(_03182_));
 sg13g2_nand2b_1 _09717_ (.Y(_03185_),
    .B(net4411),
    .A_N(net4498));
 sg13g2_o21ai_1 _09718_ (.B1(_03185_),
    .Y(_03186_),
    .A1(net4408),
    .A2(net4506));
 sg13g2_a22oi_1 _09719_ (.Y(_03187_),
    .B1(net4100),
    .B2(net4488),
    .A2(net4113),
    .A1(net4482));
 sg13g2_o21ai_1 _09720_ (.B1(_03187_),
    .Y(_03188_),
    .A1(net4391),
    .A2(_03186_));
 sg13g2_a22oi_1 _09721_ (.Y(_03189_),
    .B1(_03184_),
    .B2(net4132),
    .A2(_03180_),
    .A1(net4130));
 sg13g2_a22oi_1 _09722_ (.Y(_03190_),
    .B1(_03188_),
    .B2(net4128),
    .A2(_03177_),
    .A1(net4125));
 sg13g2_a21oi_1 _09723_ (.A1(net4408),
    .A2(_01108_),
    .Y(_03191_),
    .B1(net4391));
 sg13g2_o21ai_1 _09724_ (.B1(_03191_),
    .Y(_03192_),
    .A1(net4408),
    .A2(\cpu.keccak_alu.registers[269] ));
 sg13g2_a22oi_1 _09725_ (.Y(_03193_),
    .B1(net4100),
    .B2(\cpu.keccak_alu.registers[301] ),
    .A2(net4113),
    .A1(\cpu.keccak_alu.registers[317] ));
 sg13g2_a21o_1 _09726_ (.A2(_03193_),
    .A1(_03192_),
    .B1(net4123),
    .X(_03194_));
 sg13g2_a221oi_1 _09727_ (.B2(net4435),
    .C1(net3846),
    .B1(_03194_),
    .A1(_03189_),
    .Y(_03195_),
    .A2(_03190_));
 sg13g2_a21oi_1 _09728_ (.A1(net4069),
    .A2(_02724_),
    .Y(_03196_),
    .B1(_03195_));
 sg13g2_o21ai_1 _09729_ (.B1(_03173_),
    .Y(_00664_),
    .A1(net3740),
    .A2(_03196_));
 sg13g2_nand2_1 _09730_ (.Y(_03197_),
    .A(net107),
    .B(net3742));
 sg13g2_nand2b_1 _09731_ (.Y(_03198_),
    .B(net4404),
    .A_N(\cpu.keccak_alu.registers[30] ));
 sg13g2_o21ai_1 _09732_ (.B1(_03198_),
    .Y(_03199_),
    .A1(net4404),
    .A2(\cpu.keccak_alu.registers[14] ));
 sg13g2_a221oi_1 _09733_ (.B2(\cpu.keccak_alu.registers[46] ),
    .C1(net4434),
    .B1(net4098),
    .A1(\cpu.keccak_alu.registers[62] ),
    .Y(_03200_),
    .A2(net4111));
 sg13g2_o21ai_1 _09734_ (.B1(_03200_),
    .Y(_03201_),
    .A1(net4389),
    .A2(_03199_));
 sg13g2_nand2b_1 _09735_ (.Y(_03202_),
    .B(net4405),
    .A_N(\cpu.keccak_alu.registers[222] ));
 sg13g2_o21ai_1 _09736_ (.B1(_03202_),
    .Y(_03203_),
    .A1(net4405),
    .A2(\cpu.keccak_alu.registers[206] ));
 sg13g2_a22oi_1 _09737_ (.Y(_03204_),
    .B1(net4098),
    .B2(\cpu.keccak_alu.registers[238] ),
    .A2(net4111),
    .A1(\cpu.keccak_alu.registers[254] ));
 sg13g2_o21ai_1 _09738_ (.B1(_03204_),
    .Y(_03205_),
    .A1(net4389),
    .A2(_03203_));
 sg13g2_mux2_1 _09739_ (.A0(_01118_),
    .A1(_01119_),
    .S(net4406),
    .X(_03206_));
 sg13g2_a22oi_1 _09740_ (.Y(_03207_),
    .B1(net4098),
    .B2(\cpu.keccak_alu.registers[110] ),
    .A2(net4111),
    .A1(\cpu.keccak_alu.registers[126] ));
 sg13g2_o21ai_1 _09741_ (.B1(_03207_),
    .Y(_03208_),
    .A1(net4389),
    .A2(_03206_));
 sg13g2_nand2_1 _09742_ (.Y(_03209_),
    .A(net4409),
    .B(_01121_));
 sg13g2_o21ai_1 _09743_ (.B1(_03209_),
    .Y(_03210_),
    .A1(net4409),
    .A2(net4505));
 sg13g2_a22oi_1 _09744_ (.Y(_03211_),
    .B1(net4098),
    .B2(\cpu.keccak_alu.registers[174] ),
    .A2(net4111),
    .A1(\cpu.keccak_alu.registers[190] ));
 sg13g2_o21ai_1 _09745_ (.B1(_03211_),
    .Y(_03212_),
    .A1(net4390),
    .A2(_03210_));
 sg13g2_a22oi_1 _09746_ (.Y(_03213_),
    .B1(_03212_),
    .B2(net4128),
    .A2(_03208_),
    .A1(net4130));
 sg13g2_a22oi_1 _09747_ (.Y(_03214_),
    .B1(_03205_),
    .B2(net4132),
    .A2(_03201_),
    .A1(net4125));
 sg13g2_a21oi_1 _09748_ (.A1(net4404),
    .A2(_01123_),
    .Y(_03215_),
    .B1(net4389));
 sg13g2_o21ai_1 _09749_ (.B1(_03215_),
    .Y(_03216_),
    .A1(net4405),
    .A2(\cpu.keccak_alu.registers[270] ));
 sg13g2_a22oi_1 _09750_ (.Y(_03217_),
    .B1(net4098),
    .B2(\cpu.keccak_alu.registers[302] ),
    .A2(net4111),
    .A1(\cpu.keccak_alu.registers[318] ));
 sg13g2_a21o_1 _09751_ (.A2(_03217_),
    .A1(_03216_),
    .B1(net4123),
    .X(_03218_));
 sg13g2_a221oi_1 _09752_ (.B2(net4434),
    .C1(net3846),
    .B1(_03218_),
    .A1(_03213_),
    .Y(_03219_),
    .A2(_03214_));
 sg13g2_a21oi_1 _09753_ (.A1(net4069),
    .A2(_02732_),
    .Y(_03220_),
    .B1(_03219_));
 sg13g2_o21ai_1 _09754_ (.B1(_03197_),
    .Y(_00665_),
    .A1(net3740),
    .A2(_03220_));
 sg13g2_nand2_1 _09755_ (.Y(_03221_),
    .A(net76),
    .B(net3743));
 sg13g2_nand2b_1 _09756_ (.Y(_03222_),
    .B(net4410),
    .A_N(\cpu.keccak_alu.registers[31] ));
 sg13g2_o21ai_1 _09757_ (.B1(_03222_),
    .Y(_03223_),
    .A1(net4411),
    .A2(\cpu.keccak_alu.registers[15] ));
 sg13g2_a221oi_1 _09758_ (.B2(\cpu.keccak_alu.registers[47] ),
    .C1(net4435),
    .B1(net4101),
    .A1(\cpu.keccak_alu.registers[63] ),
    .Y(_03224_),
    .A2(net4113));
 sg13g2_o21ai_1 _09759_ (.B1(_03224_),
    .Y(_03225_),
    .A1(net4392),
    .A2(_03223_));
 sg13g2_nand2b_1 _09760_ (.Y(_03226_),
    .B(net4410),
    .A_N(\cpu.keccak_alu.registers[223] ));
 sg13g2_o21ai_1 _09761_ (.B1(_03226_),
    .Y(_03227_),
    .A1(net4412),
    .A2(\cpu.keccak_alu.registers[207] ));
 sg13g2_a22oi_1 _09762_ (.Y(_03228_),
    .B1(net4100),
    .B2(\cpu.keccak_alu.registers[239] ),
    .A2(net4113),
    .A1(\cpu.keccak_alu.registers[255] ));
 sg13g2_o21ai_1 _09763_ (.B1(_03228_),
    .Y(_03229_),
    .A1(net4392),
    .A2(_03227_));
 sg13g2_nand2b_1 _09764_ (.Y(_03230_),
    .B(net4411),
    .A_N(\cpu.keccak_alu.registers[95] ));
 sg13g2_o21ai_1 _09765_ (.B1(_03230_),
    .Y(_03231_),
    .A1(net4411),
    .A2(\cpu.keccak_alu.registers[79] ));
 sg13g2_a22oi_1 _09766_ (.Y(_03232_),
    .B1(net4100),
    .B2(\cpu.keccak_alu.registers[111] ),
    .A2(net4114),
    .A1(\cpu.keccak_alu.registers[127] ));
 sg13g2_o21ai_1 _09767_ (.B1(_03232_),
    .Y(_03233_),
    .A1(net4392),
    .A2(_03231_));
 sg13g2_a22oi_1 _09768_ (.Y(_03234_),
    .B1(_03233_),
    .B2(net4130),
    .A2(_03229_),
    .A1(net4132));
 sg13g2_nand2b_1 _09769_ (.Y(_03235_),
    .B(net4410),
    .A_N(\cpu.keccak_alu.registers[159] ));
 sg13g2_o21ai_1 _09770_ (.B1(_03235_),
    .Y(_03236_),
    .A1(net4410),
    .A2(net4504));
 sg13g2_a22oi_1 _09771_ (.Y(_03237_),
    .B1(net4100),
    .B2(\cpu.keccak_alu.registers[175] ),
    .A2(net4113),
    .A1(\cpu.keccak_alu.registers[191] ));
 sg13g2_o21ai_1 _09772_ (.B1(_03237_),
    .Y(_03238_),
    .A1(net4392),
    .A2(_03236_));
 sg13g2_a22oi_1 _09773_ (.Y(_03239_),
    .B1(_03238_),
    .B2(net4128),
    .A2(_03225_),
    .A1(net4125));
 sg13g2_a21oi_1 _09774_ (.A1(net4412),
    .A2(\cpu.keccak_alu.registers[287] ),
    .Y(_03240_),
    .B1(net4395));
 sg13g2_o21ai_1 _09775_ (.B1(_03240_),
    .Y(_03241_),
    .A1(net4412),
    .A2(_01135_));
 sg13g2_a221oi_1 _09776_ (.B2(_01137_),
    .C1(net4123),
    .B1(net4101),
    .A1(_01138_),
    .Y(_03242_),
    .A2(net4114));
 sg13g2_nand2_1 _09777_ (.Y(_03243_),
    .A(_03241_),
    .B(_03242_));
 sg13g2_a221oi_1 _09778_ (.B2(net4435),
    .C1(net3846),
    .B1(_03243_),
    .A1(_03234_),
    .Y(_03244_),
    .A2(_03239_));
 sg13g2_a21oi_2 _09779_ (.B1(_03244_),
    .Y(_03245_),
    .A2(_02739_),
    .A1(net4069));
 sg13g2_o21ai_1 _09780_ (.B1(_03221_),
    .Y(_00666_),
    .A1(net3741),
    .A2(_03245_));
 sg13g2_nand2_1 _09781_ (.Y(_03246_),
    .A(net4316),
    .B(net4078));
 sg13g2_a221oi_1 _09782_ (.B2(_00894_),
    .C1(_02742_),
    .B1(_01371_),
    .A1(net4316),
    .Y(_03247_),
    .A2(net4078));
 sg13g2_o21ai_1 _09783_ (.B1(_00017_),
    .Y(_03248_),
    .A1(net4325),
    .A2(net4450));
 sg13g2_nor2_1 _09784_ (.A(net4312),
    .B(net4078),
    .Y(_03249_));
 sg13g2_o21ai_1 _09785_ (.B1(_00896_),
    .Y(_03250_),
    .A1(_00020_),
    .A2(net4051));
 sg13g2_a22oi_1 _09786_ (.Y(_03251_),
    .B1(_03248_),
    .B2(_03249_),
    .A2(_01276_),
    .A1(net4306));
 sg13g2_nand3_1 _09787_ (.B(_03250_),
    .C(_03251_),
    .A(_03247_),
    .Y(_03252_));
 sg13g2_nor2_1 _09788_ (.A(net4301),
    .B(net809),
    .Y(_03253_));
 sg13g2_mux2_1 _09789_ (.A0(_03253_),
    .A1(net211),
    .S(_03252_),
    .X(_00667_));
 sg13g2_and3_1 _09790_ (.X(_03254_),
    .A(net4312),
    .B(_00888_),
    .C(net4233));
 sg13g2_nand3_1 _09791_ (.B(_00888_),
    .C(net4233),
    .A(net4312),
    .Y(_03255_));
 sg13g2_nor2b_1 _09792_ (.A(net4326),
    .B_N(_00149_),
    .Y(_03256_));
 sg13g2_a21oi_1 _09793_ (.A1(net4326),
    .A2(_01357_),
    .Y(_03257_),
    .B1(_03256_));
 sg13g2_a21oi_1 _09794_ (.A1(net4330),
    .A2(net4365),
    .Y(_03258_),
    .B1(_03256_));
 sg13g2_a22oi_1 _09795_ (.Y(_03259_),
    .B1(_03258_),
    .B2(_01227_),
    .A2(net4051),
    .A1(_01170_));
 sg13g2_o21ai_1 _09796_ (.B1(net3799),
    .Y(_03260_),
    .A1(net4450),
    .A2(_03259_));
 sg13g2_nor2_1 _09797_ (.A(net4335),
    .B(_00149_),
    .Y(_03261_));
 sg13g2_a21oi_1 _09798_ (.A1(net4335),
    .A2(_01356_),
    .Y(_03262_),
    .B1(_03261_));
 sg13g2_a221oi_1 _09799_ (.B2(_01251_),
    .C1(_03260_),
    .B1(_03257_),
    .A1(_01248_),
    .Y(_03263_),
    .A2(_01356_));
 sg13g2_o21ai_1 _09800_ (.B1(_03263_),
    .Y(_03264_),
    .A1(net3860),
    .A2(_03262_));
 sg13g2_a21oi_1 _09801_ (.A1(net4067),
    .A2(_03258_),
    .Y(_03265_),
    .B1(net3799));
 sg13g2_o21ai_1 _09802_ (.B1(_03265_),
    .Y(_03266_),
    .A1(net4067),
    .A2(_02160_));
 sg13g2_nand3_1 _09803_ (.B(_03264_),
    .C(_03266_),
    .A(net4317),
    .Y(_03267_));
 sg13g2_o21ai_1 _09804_ (.B1(_02625_),
    .Y(_03268_),
    .A1(_01225_),
    .A2(_03246_));
 sg13g2_nor3_1 _09805_ (.A(net4312),
    .B(\cpu.jump_con ),
    .C(_01239_),
    .Y(_03269_));
 sg13g2_a221oi_1 _09806_ (.B2(net4243),
    .C1(_03269_),
    .B1(_01425_),
    .A1(_00888_),
    .Y(_03270_),
    .A2(_01371_));
 sg13g2_o21ai_1 _09807_ (.B1(_03270_),
    .Y(_03271_),
    .A1(_00018_),
    .A2(_01289_));
 sg13g2_a21o_2 _09808_ (.A2(_03268_),
    .A1(net4071),
    .B1(_03271_),
    .X(_03272_));
 sg13g2_or2_1 _09809_ (.X(_03273_),
    .B(net3998),
    .A(_00147_));
 sg13g2_a22oi_1 _09810_ (.Y(_03274_),
    .B1(net3984),
    .B2(\cpu.registers[5][0] ),
    .A2(net3989),
    .A1(\cpu.registers[2][0] ));
 sg13g2_a21oi_1 _09811_ (.A1(\cpu.registers[7][0] ),
    .A2(_02133_),
    .Y(_03275_),
    .B1(net4070));
 sg13g2_o21ai_1 _09812_ (.B1(_03273_),
    .Y(_03276_),
    .A1(_00146_),
    .A2(net4065));
 sg13g2_a221oi_1 _09813_ (.B2(\cpu.registers[3][0] ),
    .C1(_03276_),
    .B1(net3995),
    .A1(\cpu.registers[1][0] ),
    .Y(_03277_),
    .A2(_01363_));
 sg13g2_nand3_1 _09814_ (.B(_03275_),
    .C(_03277_),
    .A(_03274_),
    .Y(_03278_));
 sg13g2_o21ai_1 _09815_ (.B1(net3944),
    .Y(_03279_),
    .A1(net3806),
    .A2(_03262_));
 sg13g2_a221oi_1 _09816_ (.B2(_01292_),
    .C1(_03279_),
    .B1(_03257_),
    .A1(net4303),
    .Y(_03280_),
    .A2(_01356_));
 sg13g2_o21ai_1 _09817_ (.B1(_03278_),
    .Y(_03281_),
    .A1(net4074),
    .A2(_02161_));
 sg13g2_a221oi_1 _09818_ (.B2(_03254_),
    .C1(net3644),
    .B1(_03281_),
    .A1(_03267_),
    .Y(_03282_),
    .A2(_03280_));
 sg13g2_a21o_1 _09819_ (.A2(net3644),
    .A1(net824),
    .B1(_03282_),
    .X(_00668_));
 sg13g2_nor2_1 _09820_ (.A(net4067),
    .B(_02167_),
    .Y(_03283_));
 sg13g2_nor2b_1 _09821_ (.A(net4329),
    .B_N(_00153_),
    .Y(_03284_));
 sg13g2_a21o_1 _09822_ (.A2(net4362),
    .A1(net4329),
    .B1(_03284_),
    .X(_03285_));
 sg13g2_o21ai_1 _09823_ (.B1(net3803),
    .Y(_03286_),
    .A1(net4065),
    .A2(_03285_));
 sg13g2_o21ai_1 _09824_ (.B1(net4319),
    .Y(_03287_),
    .A1(_03283_),
    .A2(_03286_));
 sg13g2_nor2b_1 _09825_ (.A(net4323),
    .B_N(_00210_),
    .Y(_03288_));
 sg13g2_a21o_1 _09826_ (.A2(net4271),
    .A1(net4324),
    .B1(_03288_),
    .X(_03289_));
 sg13g2_o21ai_1 _09827_ (.B1(net3801),
    .Y(_03290_),
    .A1(net4062),
    .A2(_03289_));
 sg13g2_a21oi_1 _09828_ (.A1(net4060),
    .A2(_02821_),
    .Y(_03291_),
    .B1(_03290_));
 sg13g2_nand4_1 _09829_ (.B(net4216),
    .C(net4207),
    .A(net4316),
    .Y(_03292_),
    .D(net4074));
 sg13g2_and2_2 _09830_ (.A(_01293_),
    .B(_03292_),
    .X(_03293_));
 sg13g2_nand2_2 _09831_ (.Y(_03294_),
    .A(_01293_),
    .B(_03292_));
 sg13g2_a21oi_1 _09832_ (.A1(net4329),
    .A2(_01394_),
    .Y(_03295_),
    .B1(_03284_));
 sg13g2_nor3_1 _09833_ (.A(\cpu.current_instruction[4] ),
    .B(net4078),
    .C(_03285_),
    .Y(_03296_));
 sg13g2_o21ai_1 _09834_ (.B1(net3799),
    .Y(_03297_),
    .A1(net4362),
    .A2(_01247_));
 sg13g2_nor2_1 _09835_ (.A(_03296_),
    .B(_03297_),
    .Y(_03298_));
 sg13g2_o21ai_1 _09836_ (.B1(net3944),
    .Y(_03299_),
    .A1(_03287_),
    .A2(_03298_));
 sg13g2_or2_2 _09837_ (.X(_03300_),
    .B(_03287_),
    .A(net3860));
 sg13g2_nor2_1 _09838_ (.A(net4204),
    .B(_01395_),
    .Y(_03301_));
 sg13g2_a221oi_1 _09839_ (.B2(_03300_),
    .C1(_03301_),
    .B1(net3806),
    .A1(net4204),
    .Y(_03302_),
    .A2(_00153_));
 sg13g2_o21ai_1 _09840_ (.B1(_00888_),
    .Y(_03303_),
    .A1(_01249_),
    .A2(_03287_));
 sg13g2_a21oi_1 _09841_ (.A1(_03294_),
    .A2(_03295_),
    .Y(_03304_),
    .B1(_03302_));
 sg13g2_a21oi_1 _09842_ (.A1(_01395_),
    .A2(_03303_),
    .Y(_03305_),
    .B1(_03299_));
 sg13g2_nand2b_1 _09843_ (.Y(_03306_),
    .B(_02133_),
    .A_N(_00031_));
 sg13g2_or2_1 _09844_ (.X(_03307_),
    .B(net3998),
    .A(_00151_));
 sg13g2_a22oi_1 _09845_ (.Y(_03308_),
    .B1(net3990),
    .B2(\cpu.registers[2][1] ),
    .A2(_01363_),
    .A1(_01181_));
 sg13g2_o21ai_1 _09846_ (.B1(_03307_),
    .Y(_03309_),
    .A1(_00150_),
    .A2(net4063));
 sg13g2_a221oi_1 _09847_ (.B2(\cpu.registers[5][1] ),
    .C1(_03309_),
    .B1(net3985),
    .A1(\cpu.registers[3][1] ),
    .Y(_03310_),
    .A2(net3995));
 sg13g2_nand4_1 _09848_ (.B(_03306_),
    .C(_03308_),
    .A(net4075),
    .Y(_03311_),
    .D(_03310_));
 sg13g2_o21ai_1 _09849_ (.B1(_03311_),
    .Y(_03312_),
    .A1(net4075),
    .A2(_02168_));
 sg13g2_a221oi_1 _09850_ (.B2(_03254_),
    .C1(net3642),
    .B1(_03312_),
    .A1(_03304_),
    .Y(_03313_),
    .A2(_03305_));
 sg13g2_a21o_1 _09851_ (.A2(net3642),
    .A1(net863),
    .B1(_03313_),
    .X(_00669_));
 sg13g2_nand2_1 _09852_ (.Y(_03314_),
    .A(net4303),
    .B(_01475_));
 sg13g2_nor2b_1 _09853_ (.A(net4329),
    .B_N(_00157_),
    .Y(_03315_));
 sg13g2_o21ai_1 _09854_ (.B1(_03294_),
    .Y(_03316_),
    .A1(net4242),
    .A2(_01475_));
 sg13g2_nor2_1 _09855_ (.A(net4067),
    .B(_02175_),
    .Y(_03317_));
 sg13g2_a21o_1 _09856_ (.A2(net4354),
    .A1(net4329),
    .B1(_03315_),
    .X(_03318_));
 sg13g2_o21ai_1 _09857_ (.B1(net3804),
    .Y(_03319_),
    .A1(net4064),
    .A2(_03318_));
 sg13g2_o21ai_1 _09858_ (.B1(net4319),
    .Y(_03320_),
    .A1(_03317_),
    .A2(_03319_));
 sg13g2_a21oi_1 _09859_ (.A1(net4240),
    .A2(net4354),
    .Y(_03321_),
    .B1(net3866));
 sg13g2_or2_1 _09860_ (.X(_03322_),
    .B(_03318_),
    .A(net4079));
 sg13g2_o21ai_1 _09861_ (.B1(_03322_),
    .Y(_03323_),
    .A1(net4354),
    .A2(net3866));
 sg13g2_a221oi_1 _09862_ (.B2(net4241),
    .C1(net3803),
    .B1(_03323_),
    .A1(_01475_),
    .Y(_03324_),
    .A2(_03321_));
 sg13g2_a21o_1 _09863_ (.A2(_03322_),
    .A1(net3860),
    .B1(_03320_),
    .X(_03325_));
 sg13g2_a22oi_1 _09864_ (.Y(_03326_),
    .B1(net3806),
    .B2(_03325_),
    .A2(_00157_),
    .A1(net4204));
 sg13g2_o21ai_1 _09865_ (.B1(_03326_),
    .Y(_03327_),
    .A1(net4204),
    .A2(_01475_));
 sg13g2_o21ai_1 _09866_ (.B1(_03314_),
    .Y(_03328_),
    .A1(_03320_),
    .A2(_03324_));
 sg13g2_o21ai_1 _09867_ (.B1(_03327_),
    .Y(_03329_),
    .A1(_03315_),
    .A2(_03316_));
 sg13g2_o21ai_1 _09868_ (.B1(net3944),
    .Y(_03330_),
    .A1(_03328_),
    .A2(_03329_));
 sg13g2_nor2_1 _09869_ (.A(_00156_),
    .B(net4148),
    .Y(_03331_));
 sg13g2_nand2_1 _09870_ (.Y(_03332_),
    .A(\cpu.registers[3][2] ),
    .B(net3995));
 sg13g2_o21ai_1 _09871_ (.B1(net4074),
    .Y(_03333_),
    .A1(_00155_),
    .A2(net3998));
 sg13g2_nor2_1 _09872_ (.A(_00032_),
    .B(net3987),
    .Y(_03334_));
 sg13g2_o21ai_1 _09873_ (.B1(_03332_),
    .Y(_03335_),
    .A1(_00154_),
    .A2(net4065));
 sg13g2_a221oi_1 _09874_ (.B2(\cpu.registers[5][2] ),
    .C1(_03335_),
    .B1(net3984),
    .A1(\cpu.registers[2][2] ),
    .Y(_03336_),
    .A2(net3989));
 sg13g2_nor3_1 _09875_ (.A(_03331_),
    .B(_03333_),
    .C(_03334_),
    .Y(_03337_));
 sg13g2_a22oi_1 _09876_ (.Y(_03338_),
    .B1(_03336_),
    .B2(_03337_),
    .A2(_02175_),
    .A1(net4070));
 sg13g2_a21oi_1 _09877_ (.A1(net3946),
    .A2(_03338_),
    .Y(_03339_),
    .B1(net3644));
 sg13g2_a22oi_1 _09878_ (.Y(_00670_),
    .B1(_03330_),
    .B2(_03339_),
    .A2(net3644),
    .A1(_01146_));
 sg13g2_nor2_1 _09879_ (.A(net4327),
    .B(_00161_),
    .Y(_03340_));
 sg13g2_a21oi_1 _09880_ (.A1(net4327),
    .A2(_01171_),
    .Y(_03341_),
    .B1(_03340_));
 sg13g2_nor2_1 _09881_ (.A(net4065),
    .B(_03341_),
    .Y(_03342_));
 sg13g2_a21oi_1 _09882_ (.A1(net4064),
    .A2(_02184_),
    .Y(_03343_),
    .B1(_03342_));
 sg13g2_a21oi_1 _09883_ (.A1(net3803),
    .A2(_03343_),
    .Y(_03344_),
    .B1(net4261));
 sg13g2_nor2_1 _09884_ (.A(net4079),
    .B(_03341_),
    .Y(_03345_));
 sg13g2_nand2b_1 _09885_ (.Y(_03346_),
    .B(_01254_),
    .A_N(_03345_));
 sg13g2_a21oi_1 _09886_ (.A1(_03344_),
    .A2(_03346_),
    .Y(_03347_),
    .B1(_01290_));
 sg13g2_a21oi_1 _09887_ (.A1(net4240),
    .A2(net4352),
    .Y(_03348_),
    .B1(net3867));
 sg13g2_a221oi_1 _09888_ (.B2(_03348_),
    .C1(net4303),
    .B1(_03344_),
    .A1(net4327),
    .Y(_03349_),
    .A2(_03294_));
 sg13g2_o21ai_1 _09889_ (.B1(_03349_),
    .Y(_03350_),
    .A1(net4205),
    .A2(_03347_));
 sg13g2_nor3_1 _09890_ (.A(net4335),
    .B(net891),
    .C(_03347_),
    .Y(_03351_));
 sg13g2_nor3_1 _09891_ (.A(net4327),
    .B(_00161_),
    .C(_03293_),
    .Y(_03352_));
 sg13g2_a21oi_1 _09892_ (.A1(_01171_),
    .A2(net4055),
    .Y(_03353_),
    .B1(_03345_));
 sg13g2_o21ai_1 _09893_ (.B1(net3800),
    .Y(_03354_),
    .A1(net4452),
    .A2(_03353_));
 sg13g2_a221oi_1 _09894_ (.B2(_03344_),
    .C1(_03352_),
    .B1(_03354_),
    .A1(_01509_),
    .Y(_03355_),
    .A2(_03350_));
 sg13g2_inv_1 _09895_ (.Y(_03356_),
    .A(_03355_));
 sg13g2_o21ai_1 _09896_ (.B1(net3944),
    .Y(_03357_),
    .A1(_03351_),
    .A2(_03356_));
 sg13g2_nand2_1 _09897_ (.Y(_03358_),
    .A(\cpu.registers[2][3] ),
    .B(net3989));
 sg13g2_nand2_1 _09898_ (.Y(_03359_),
    .A(\cpu.registers[5][3] ),
    .B(net3984));
 sg13g2_a22oi_1 _09899_ (.Y(_03360_),
    .B1(net3995),
    .B2(\cpu.registers[3][3] ),
    .A2(_01363_),
    .A1(_01182_));
 sg13g2_o21ai_1 _09900_ (.B1(_03359_),
    .Y(_03361_),
    .A1(_00159_),
    .A2(net3999));
 sg13g2_o21ai_1 _09901_ (.B1(_03358_),
    .Y(_03362_),
    .A1(_00158_),
    .A2(net4063));
 sg13g2_o21ai_1 _09902_ (.B1(net4075),
    .Y(_03363_),
    .A1(_00033_),
    .A2(net3987));
 sg13g2_nor3_1 _09903_ (.A(_03361_),
    .B(_03362_),
    .C(_03363_),
    .Y(_03364_));
 sg13g2_a22oi_1 _09904_ (.Y(_03365_),
    .B1(_03360_),
    .B2(_03364_),
    .A2(_02183_),
    .A1(net4072));
 sg13g2_a21oi_1 _09905_ (.A1(net3946),
    .A2(_03365_),
    .Y(_03366_),
    .B1(net3643));
 sg13g2_a22oi_1 _09906_ (.Y(_00671_),
    .B1(_03357_),
    .B2(_03366_),
    .A2(net3642),
    .A1(_01147_));
 sg13g2_nor2b_1 _09907_ (.A(net4327),
    .B_N(_00165_),
    .Y(_03367_));
 sg13g2_a21oi_1 _09908_ (.A1(net4327),
    .A2(_01551_),
    .Y(_03368_),
    .B1(_03367_));
 sg13g2_a21o_1 _09909_ (.A2(net4348),
    .A1(net4327),
    .B1(_03367_),
    .X(_03369_));
 sg13g2_nor2_1 _09910_ (.A(net4063),
    .B(_03369_),
    .Y(_03370_));
 sg13g2_a21oi_1 _09911_ (.A1(net4065),
    .A2(_02192_),
    .Y(_03371_),
    .B1(_03370_));
 sg13g2_a21oi_1 _09912_ (.A1(net3803),
    .A2(_03371_),
    .Y(_03372_),
    .B1(net4261));
 sg13g2_nor2_1 _09913_ (.A(net4079),
    .B(_03369_),
    .Y(_03373_));
 sg13g2_nand2b_1 _09914_ (.Y(_03374_),
    .B(net3860),
    .A_N(_03373_));
 sg13g2_nand2_1 _09915_ (.Y(_03375_),
    .A(_03372_),
    .B(_03374_));
 sg13g2_nor2b_1 _09916_ (.A(net4335),
    .B_N(_00165_),
    .Y(_03376_));
 sg13g2_a221oi_1 _09917_ (.B2(net3806),
    .C1(_03376_),
    .B1(_03375_),
    .A1(net4335),
    .Y(_03377_),
    .A2(_01551_));
 sg13g2_a21oi_1 _09918_ (.A1(net4240),
    .A2(net4348),
    .Y(_03378_),
    .B1(net3868));
 sg13g2_a21oi_1 _09919_ (.A1(_03372_),
    .A2(_03378_),
    .Y(_03379_),
    .B1(net4303));
 sg13g2_a21oi_1 _09920_ (.A1(net4156),
    .A2(net4055),
    .Y(_03380_),
    .B1(_03373_));
 sg13g2_o21ai_1 _09921_ (.B1(net3798),
    .Y(_03381_),
    .A1(net4452),
    .A2(_03380_));
 sg13g2_a221oi_1 _09922_ (.B2(_03381_),
    .C1(_03377_),
    .B1(_03372_),
    .A1(_03294_),
    .Y(_03382_),
    .A2(_03368_));
 sg13g2_o21ai_1 _09923_ (.B1(_03382_),
    .Y(_03383_),
    .A1(_01551_),
    .A2(_03379_));
 sg13g2_nand2_1 _09924_ (.Y(_03384_),
    .A(net3944),
    .B(_03383_));
 sg13g2_nand2_1 _09925_ (.Y(_03385_),
    .A(\cpu.registers[2][4] ),
    .B(net3989));
 sg13g2_nor2_1 _09926_ (.A(_00034_),
    .B(net3987),
    .Y(_03386_));
 sg13g2_nor2_1 _09927_ (.A(_00163_),
    .B(net3998),
    .Y(_03387_));
 sg13g2_a22oi_1 _09928_ (.Y(_03388_),
    .B1(net3984),
    .B2(\cpu.registers[5][4] ),
    .A2(net3995),
    .A1(\cpu.registers[3][4] ));
 sg13g2_o21ai_1 _09929_ (.B1(_03385_),
    .Y(_03389_),
    .A1(_00164_),
    .A2(net4148));
 sg13g2_o21ai_1 _09930_ (.B1(net4074),
    .Y(_03390_),
    .A1(_00162_),
    .A2(net4063));
 sg13g2_nor4_1 _09931_ (.A(_03386_),
    .B(_03387_),
    .C(_03389_),
    .D(_03390_),
    .Y(_03391_));
 sg13g2_a22oi_1 _09932_ (.Y(_03392_),
    .B1(_03388_),
    .B2(_03391_),
    .A2(_02191_),
    .A1(net4072));
 sg13g2_a21oi_1 _09933_ (.A1(net3946),
    .A2(_03392_),
    .Y(_03393_),
    .B1(net3643));
 sg13g2_a22oi_1 _09934_ (.Y(_00672_),
    .B1(_03384_),
    .B2(_03393_),
    .A2(net3642),
    .A1(_01148_));
 sg13g2_nor2b_1 _09935_ (.A(net4328),
    .B_N(_00169_),
    .Y(_03394_));
 sg13g2_a21o_1 _09936_ (.A2(net4345),
    .A1(net4328),
    .B1(_03394_),
    .X(_03395_));
 sg13g2_nor2_1 _09937_ (.A(net4064),
    .B(_03395_),
    .Y(_03396_));
 sg13g2_a21oi_1 _09938_ (.A1(net4064),
    .A2(_02199_),
    .Y(_03397_),
    .B1(_03396_));
 sg13g2_a21oi_1 _09939_ (.A1(net3803),
    .A2(_03397_),
    .Y(_03398_),
    .B1(net4261));
 sg13g2_nor2_1 _09940_ (.A(net4079),
    .B(_03395_),
    .Y(_03399_));
 sg13g2_nand2b_1 _09941_ (.Y(_03400_),
    .B(net3860),
    .A_N(_03399_));
 sg13g2_nand2_1 _09942_ (.Y(_03401_),
    .A(_03398_),
    .B(_03400_));
 sg13g2_a22oi_1 _09943_ (.Y(_03402_),
    .B1(net3805),
    .B2(_03401_),
    .A2(_00169_),
    .A1(net4204));
 sg13g2_a21oi_1 _09944_ (.A1(net4240),
    .A2(net4345),
    .Y(_03403_),
    .B1(net3867));
 sg13g2_a21oi_1 _09945_ (.A1(_03398_),
    .A2(_03403_),
    .Y(_03404_),
    .B1(net4303));
 sg13g2_o21ai_1 _09946_ (.B1(_03404_),
    .Y(_03405_),
    .A1(_03293_),
    .A2(_03394_));
 sg13g2_nor2_1 _09947_ (.A(_03402_),
    .B(_03405_),
    .Y(_03406_));
 sg13g2_a21oi_1 _09948_ (.A1(_01173_),
    .A2(net4055),
    .Y(_03407_),
    .B1(_03399_));
 sg13g2_o21ai_1 _09949_ (.B1(net3798),
    .Y(_03408_),
    .A1(net4452),
    .A2(_03407_));
 sg13g2_nor3_1 _09950_ (.A(net4328),
    .B(_00169_),
    .C(_03293_),
    .Y(_03409_));
 sg13g2_a221oi_1 _09951_ (.B2(_03398_),
    .C1(_03409_),
    .B1(_03408_),
    .A1(net4204),
    .Y(_03410_),
    .A2(_03402_));
 sg13g2_o21ai_1 _09952_ (.B1(_03410_),
    .Y(_03411_),
    .A1(_01595_),
    .A2(_03406_));
 sg13g2_nand2_1 _09953_ (.Y(_03412_),
    .A(net3944),
    .B(_03411_));
 sg13g2_nand2_1 _09954_ (.Y(_03413_),
    .A(\cpu.registers[3][5] ),
    .B(_01924_));
 sg13g2_o21ai_1 _09955_ (.B1(_03413_),
    .Y(_03414_),
    .A1(_00166_),
    .A2(net4063));
 sg13g2_a221oi_1 _09956_ (.B2(\cpu.registers[5][5] ),
    .C1(_03414_),
    .B1(net3984),
    .A1(\cpu.registers[2][5] ),
    .Y(_03415_),
    .A2(net3989));
 sg13g2_o21ai_1 _09957_ (.B1(net4075),
    .Y(_03416_),
    .A1(_00168_),
    .A2(net4148));
 sg13g2_nor2_1 _09958_ (.A(_00167_),
    .B(net3998),
    .Y(_03417_));
 sg13g2_nor2_1 _09959_ (.A(_00035_),
    .B(net3987),
    .Y(_03418_));
 sg13g2_nor3_1 _09960_ (.A(_03416_),
    .B(_03417_),
    .C(_03418_),
    .Y(_03419_));
 sg13g2_a22oi_1 _09961_ (.Y(_03420_),
    .B1(_03415_),
    .B2(_03419_),
    .A2(_02198_),
    .A1(net4072));
 sg13g2_a21oi_1 _09962_ (.A1(net3946),
    .A2(_03420_),
    .Y(_03421_),
    .B1(net3643));
 sg13g2_a22oi_1 _09963_ (.Y(_00673_),
    .B1(_03412_),
    .B2(_03421_),
    .A2(net3642),
    .A1(_01149_));
 sg13g2_nand2_1 _09964_ (.Y(_03422_),
    .A(net4242),
    .B(_00173_));
 sg13g2_o21ai_1 _09965_ (.B1(_03422_),
    .Y(_03423_),
    .A1(net4243),
    .A2(net4155));
 sg13g2_nor2_1 _09966_ (.A(net4063),
    .B(_03423_),
    .Y(_03424_));
 sg13g2_a21oi_1 _09967_ (.A1(net4063),
    .A2(_02207_),
    .Y(_03425_),
    .B1(_03424_));
 sg13g2_a21oi_1 _09968_ (.A1(net3803),
    .A2(_03425_),
    .Y(_03426_),
    .B1(net4261));
 sg13g2_nor2_1 _09969_ (.A(net4078),
    .B(_03423_),
    .Y(_03427_));
 sg13g2_o21ai_1 _09970_ (.B1(net3860),
    .Y(_03428_),
    .A1(net4078),
    .A2(_03423_));
 sg13g2_a21oi_1 _09971_ (.A1(_03426_),
    .A2(_03428_),
    .Y(_03429_),
    .B1(_01290_));
 sg13g2_a21o_1 _09972_ (.A2(_00173_),
    .A1(net4205),
    .B1(_03429_),
    .X(_03430_));
 sg13g2_a21oi_1 _09973_ (.A1(net4240),
    .A2(net4341),
    .Y(_03431_),
    .B1(net3867));
 sg13g2_a221oi_1 _09974_ (.B2(_03431_),
    .C1(net4303),
    .B1(_03426_),
    .A1(_03294_),
    .Y(_03432_),
    .A2(_03422_));
 sg13g2_a21oi_1 _09975_ (.A1(_03430_),
    .A2(_03432_),
    .Y(_03433_),
    .B1(_01648_));
 sg13g2_a21oi_1 _09976_ (.A1(net4155),
    .A2(net4055),
    .Y(_03434_),
    .B1(_03427_));
 sg13g2_o21ai_1 _09977_ (.B1(net3798),
    .Y(_03435_),
    .A1(net4452),
    .A2(_03434_));
 sg13g2_nor3_1 _09978_ (.A(net4328),
    .B(_00173_),
    .C(net3795),
    .Y(_03436_));
 sg13g2_a21oi_1 _09979_ (.A1(_03426_),
    .A2(_03435_),
    .Y(_03437_),
    .B1(_03436_));
 sg13g2_o21ai_1 _09980_ (.B1(_03437_),
    .Y(_03438_),
    .A1(net4335),
    .A2(_03430_));
 sg13g2_o21ai_1 _09981_ (.B1(net3943),
    .Y(_03439_),
    .A1(_03433_),
    .A2(_03438_));
 sg13g2_nor2_1 _09982_ (.A(_00172_),
    .B(net4148),
    .Y(_03440_));
 sg13g2_o21ai_1 _09983_ (.B1(net4075),
    .Y(_03441_),
    .A1(_00171_),
    .A2(net3998));
 sg13g2_nand2_1 _09984_ (.Y(_03442_),
    .A(\cpu.registers[2][6] ),
    .B(net3989));
 sg13g2_nor2_1 _09985_ (.A(_00036_),
    .B(net3986),
    .Y(_03443_));
 sg13g2_o21ai_1 _09986_ (.B1(_03442_),
    .Y(_03444_),
    .A1(_00170_),
    .A2(net4063));
 sg13g2_a221oi_1 _09987_ (.B2(\cpu.registers[5][6] ),
    .C1(_03444_),
    .B1(net3984),
    .A1(\cpu.registers[3][6] ),
    .Y(_03445_),
    .A2(net3995));
 sg13g2_nor3_1 _09988_ (.A(_03440_),
    .B(_03441_),
    .C(_03443_),
    .Y(_03446_));
 sg13g2_a22oi_1 _09989_ (.Y(_03447_),
    .B1(_03445_),
    .B2(_03446_),
    .A2(_02206_),
    .A1(net4072));
 sg13g2_a21oi_1 _09990_ (.A1(net3946),
    .A2(_03447_),
    .Y(_03448_),
    .B1(net3643));
 sg13g2_a22oi_1 _09991_ (.Y(_00674_),
    .B1(_03439_),
    .B2(_03448_),
    .A2(net3642),
    .A1(_01150_));
 sg13g2_nor2b_1 _09992_ (.A(net4329),
    .B_N(_00177_),
    .Y(_03449_));
 sg13g2_a21o_1 _09993_ (.A2(net4338),
    .A1(net4329),
    .B1(_03449_),
    .X(_03450_));
 sg13g2_nor2_1 _09994_ (.A(net4064),
    .B(_03450_),
    .Y(_03451_));
 sg13g2_a21oi_1 _09995_ (.A1(net4064),
    .A2(_02215_),
    .Y(_03452_),
    .B1(_03451_));
 sg13g2_a21oi_1 _09996_ (.A1(net3803),
    .A2(_03452_),
    .Y(_03453_),
    .B1(net4262));
 sg13g2_nor2_1 _09997_ (.A(net4079),
    .B(_03450_),
    .Y(_03454_));
 sg13g2_nand2b_1 _09998_ (.Y(_03455_),
    .B(net3860),
    .A_N(_03454_));
 sg13g2_nand2_1 _09999_ (.Y(_03456_),
    .A(_03453_),
    .B(_03455_));
 sg13g2_a22oi_1 _10000_ (.Y(_03457_),
    .B1(net3805),
    .B2(_03456_),
    .A2(_00177_),
    .A1(net4204));
 sg13g2_a21oi_1 _10001_ (.A1(net4240),
    .A2(net4338),
    .Y(_03458_),
    .B1(net3865));
 sg13g2_a21oi_1 _10002_ (.A1(_03453_),
    .A2(_03458_),
    .Y(_03459_),
    .B1(net4302));
 sg13g2_o21ai_1 _10003_ (.B1(_03459_),
    .Y(_03460_),
    .A1(net3795),
    .A2(_03449_));
 sg13g2_nor2_1 _10004_ (.A(_03457_),
    .B(_03460_),
    .Y(_03461_));
 sg13g2_a21oi_1 _10005_ (.A1(_01175_),
    .A2(net4053),
    .Y(_03462_),
    .B1(_03454_));
 sg13g2_o21ai_1 _10006_ (.B1(net3799),
    .Y(_03463_),
    .A1(net4452),
    .A2(_03462_));
 sg13g2_nor3_1 _10007_ (.A(net4329),
    .B(_00177_),
    .C(net3795),
    .Y(_03464_));
 sg13g2_a221oi_1 _10008_ (.B2(_03453_),
    .C1(_03464_),
    .B1(_03463_),
    .A1(net4204),
    .Y(_03465_),
    .A2(_03457_));
 sg13g2_o21ai_1 _10009_ (.B1(_03465_),
    .Y(_03466_),
    .A1(_01706_),
    .A2(_03461_));
 sg13g2_nand2_1 _10010_ (.Y(_03467_),
    .A(net3944),
    .B(_03466_));
 sg13g2_nor2_1 _10011_ (.A(_00175_),
    .B(net3998),
    .Y(_03468_));
 sg13g2_nor2_1 _10012_ (.A(_00174_),
    .B(net4064),
    .Y(_03469_));
 sg13g2_nand2_1 _10013_ (.Y(_03470_),
    .A(\cpu.registers[2][7] ),
    .B(net3989));
 sg13g2_a22oi_1 _10014_ (.Y(_03471_),
    .B1(net3984),
    .B2(\cpu.registers[5][7] ),
    .A2(net3995),
    .A1(\cpu.registers[3][7] ));
 sg13g2_o21ai_1 _10015_ (.B1(_03470_),
    .Y(_03472_),
    .A1(_00176_),
    .A2(net4148));
 sg13g2_o21ai_1 _10016_ (.B1(net4075),
    .Y(_03473_),
    .A1(_00037_),
    .A2(net3986));
 sg13g2_nor4_1 _10017_ (.A(_03468_),
    .B(_03469_),
    .C(_03472_),
    .D(_03473_),
    .Y(_03474_));
 sg13g2_a22oi_1 _10018_ (.Y(_03475_),
    .B1(_03471_),
    .B2(_03474_),
    .A2(_02214_),
    .A1(net4072));
 sg13g2_a21oi_1 _10019_ (.A1(net3946),
    .A2(_03475_),
    .Y(_03476_),
    .B1(net3642));
 sg13g2_a22oi_1 _10020_ (.Y(_00675_),
    .B1(_03467_),
    .B2(_03476_),
    .A2(net3642),
    .A1(_01152_));
 sg13g2_nand2b_1 _10021_ (.Y(_03477_),
    .B(net3640),
    .A_N(net855));
 sg13g2_nor2b_1 _10022_ (.A(net4322),
    .B_N(_00181_),
    .Y(_03478_));
 sg13g2_or2_1 _10023_ (.X(_03479_),
    .B(_03478_),
    .A(net3795));
 sg13g2_nand2_1 _10024_ (.Y(_03480_),
    .A(net4202),
    .B(_00181_));
 sg13g2_a21o_1 _10025_ (.A2(net4297),
    .A1(net4322),
    .B1(_03478_),
    .X(_03481_));
 sg13g2_nor2_1 _10026_ (.A(net4060),
    .B(_03481_),
    .Y(_03482_));
 sg13g2_o21ai_1 _10027_ (.B1(net3801),
    .Y(_03483_),
    .A1(net4067),
    .A2(_02222_));
 sg13g2_o21ai_1 _10028_ (.B1(net4314),
    .Y(_03484_),
    .A1(_03482_),
    .A2(_03483_));
 sg13g2_or2_1 _10029_ (.X(_03485_),
    .B(_03481_),
    .A(net4077));
 sg13g2_a21oi_1 _10030_ (.A1(net3861),
    .A2(_03485_),
    .Y(_03486_),
    .B1(_03484_));
 sg13g2_o21ai_1 _10031_ (.B1(_03480_),
    .Y(_03487_),
    .A1(_01290_),
    .A2(_03486_));
 sg13g2_nand2_1 _10032_ (.Y(_03488_),
    .A(net4237),
    .B(net4297));
 sg13g2_nand3_1 _10033_ (.B(net4050),
    .C(_03488_),
    .A(net4314),
    .Y(_03489_));
 sg13g2_nand4_1 _10034_ (.B(_03479_),
    .C(_03487_),
    .A(_00888_),
    .Y(_03490_),
    .D(_03489_));
 sg13g2_o21ai_1 _10035_ (.B1(_03485_),
    .Y(_03491_),
    .A1(net4297),
    .A2(net3863));
 sg13g2_a21oi_1 _10036_ (.A1(net4237),
    .A2(_03491_),
    .Y(_03492_),
    .B1(net3801));
 sg13g2_nor2_1 _10037_ (.A(_03484_),
    .B(_03492_),
    .Y(_03493_));
 sg13g2_nor2_1 _10038_ (.A(net4323),
    .B(_03479_),
    .Y(_03494_));
 sg13g2_nor2_1 _10039_ (.A(_03493_),
    .B(_03494_),
    .Y(_03495_));
 sg13g2_o21ai_1 _10040_ (.B1(_03495_),
    .Y(_03496_),
    .A1(net4334),
    .A2(_03487_));
 sg13g2_a21oi_1 _10041_ (.A1(_01755_),
    .A2(_03490_),
    .Y(_03497_),
    .B1(_03496_));
 sg13g2_nor2_1 _10042_ (.A(_00961_),
    .B(_01925_),
    .Y(_03498_));
 sg13g2_or2_1 _10043_ (.X(_03499_),
    .B(net3997),
    .A(_00179_));
 sg13g2_nand2_1 _10044_ (.Y(_03500_),
    .A(\cpu.registers[2][8] ),
    .B(net3988));
 sg13g2_a22oi_1 _10045_ (.Y(_03501_),
    .B1(net3983),
    .B2(\cpu.registers[5][8] ),
    .A2(_01363_),
    .A1(_01183_));
 sg13g2_o21ai_1 _10046_ (.B1(_03500_),
    .Y(_03502_),
    .A1(_00178_),
    .A2(net4060));
 sg13g2_o21ai_1 _10047_ (.B1(_03499_),
    .Y(_03503_),
    .A1(_00038_),
    .A2(net3986));
 sg13g2_nor4_1 _10048_ (.A(net4068),
    .B(_03498_),
    .C(_03502_),
    .D(_03503_),
    .Y(_03504_));
 sg13g2_a22oi_1 _10049_ (.Y(_03505_),
    .B1(_03501_),
    .B2(_03504_),
    .A2(_02222_),
    .A1(net4068));
 sg13g2_a21oi_1 _10050_ (.A1(net3945),
    .A2(_03505_),
    .Y(_03506_),
    .B1(net3640));
 sg13g2_o21ai_1 _10051_ (.B1(_03506_),
    .Y(_03507_),
    .A1(net3945),
    .A2(_03497_));
 sg13g2_and2_1 _10052_ (.A(_03477_),
    .B(_03507_),
    .X(_00676_));
 sg13g2_nand2_1 _10053_ (.Y(_03508_),
    .A(net4242),
    .B(_00185_));
 sg13g2_o21ai_1 _10054_ (.B1(_03508_),
    .Y(_03509_),
    .A1(net4242),
    .A2(net4154));
 sg13g2_nor2_1 _10055_ (.A(net4062),
    .B(_03509_),
    .Y(_03510_));
 sg13g2_a21oi_1 _10056_ (.A1(net4062),
    .A2(_02230_),
    .Y(_03511_),
    .B1(_03510_));
 sg13g2_a21oi_1 _10057_ (.A1(net3802),
    .A2(_03511_),
    .Y(_03512_),
    .B1(net4256));
 sg13g2_or2_1 _10058_ (.X(_03513_),
    .B(_03509_),
    .A(net4077));
 sg13g2_nand2_1 _10059_ (.Y(_03514_),
    .A(net3861),
    .B(_03513_));
 sg13g2_nand2_1 _10060_ (.Y(_03515_),
    .A(_03512_),
    .B(_03514_));
 sg13g2_a22oi_1 _10061_ (.Y(_03516_),
    .B1(net3805),
    .B2(_03515_),
    .A2(_00185_),
    .A1(net4202));
 sg13g2_a21oi_1 _10062_ (.A1(net4238),
    .A2(net4293),
    .Y(_03517_),
    .B1(net3863));
 sg13g2_a21oi_1 _10063_ (.A1(_03512_),
    .A2(_03517_),
    .Y(_03518_),
    .B1(net4302));
 sg13g2_o21ai_1 _10064_ (.B1(_03513_),
    .Y(_03519_),
    .A1(net4293),
    .A2(net3863));
 sg13g2_a21oi_1 _10065_ (.A1(net4237),
    .A2(_03519_),
    .Y(_03520_),
    .B1(net3802));
 sg13g2_nand2b_1 _10066_ (.Y(_03521_),
    .B(_03512_),
    .A_N(_03520_));
 sg13g2_a21oi_1 _10067_ (.A1(net4323),
    .A2(_01779_),
    .Y(_03522_),
    .B1(net3795));
 sg13g2_nand2_1 _10068_ (.Y(_03523_),
    .A(net4334),
    .B(_01779_));
 sg13g2_nor2_1 _10069_ (.A(_01779_),
    .B(_03518_),
    .Y(_03524_));
 sg13g2_a221oi_1 _10070_ (.B2(_03516_),
    .C1(_03524_),
    .B1(_03523_),
    .A1(_03508_),
    .Y(_03525_),
    .A2(_03522_));
 sg13g2_a21oi_1 _10071_ (.A1(_03521_),
    .A2(_03525_),
    .Y(_03526_),
    .B1(net3945));
 sg13g2_nand2_1 _10072_ (.Y(_03527_),
    .A(\cpu.registers[5][9] ),
    .B(net3985));
 sg13g2_nor2_1 _10073_ (.A(_00039_),
    .B(net3986),
    .Y(_03528_));
 sg13g2_nor2_1 _10074_ (.A(_00184_),
    .B(net4149),
    .Y(_03529_));
 sg13g2_a22oi_1 _10075_ (.Y(_03530_),
    .B1(net3990),
    .B2(\cpu.registers[2][9] ),
    .A2(net3996),
    .A1(\cpu.registers[3][9] ));
 sg13g2_o21ai_1 _10076_ (.B1(_03527_),
    .Y(_03531_),
    .A1(_00183_),
    .A2(net3997));
 sg13g2_o21ai_1 _10077_ (.B1(net4076),
    .Y(_03532_),
    .A1(_00182_),
    .A2(net4062));
 sg13g2_nor4_1 _10078_ (.A(_03528_),
    .B(_03529_),
    .C(_03531_),
    .D(_03532_),
    .Y(_03533_));
 sg13g2_a221oi_1 _10079_ (.B2(_03533_),
    .C1(net3943),
    .B1(_03530_),
    .A1(net4069),
    .Y(_03534_),
    .A2(_02229_));
 sg13g2_nor3_1 _10080_ (.A(net3641),
    .B(_03526_),
    .C(_03534_),
    .Y(_03535_));
 sg13g2_a21oi_1 _10081_ (.A1(_01154_),
    .A2(net3641),
    .Y(_00677_),
    .B1(_03535_));
 sg13g2_nor2_1 _10082_ (.A(net4322),
    .B(_01186_),
    .Y(_03536_));
 sg13g2_a21o_1 _10083_ (.A2(net4289),
    .A1(net4322),
    .B1(_03536_),
    .X(_03537_));
 sg13g2_nor2_1 _10084_ (.A(net4061),
    .B(_03537_),
    .Y(_03538_));
 sg13g2_a21oi_1 _10085_ (.A1(net4060),
    .A2(_02237_),
    .Y(_03539_),
    .B1(_03538_));
 sg13g2_a21oi_1 _10086_ (.A1(net3801),
    .A2(_03539_),
    .Y(_03540_),
    .B1(net4253));
 sg13g2_nor2_1 _10087_ (.A(net4077),
    .B(_03537_),
    .Y(_03541_));
 sg13g2_nand2b_1 _10088_ (.Y(_03542_),
    .B(net3861),
    .A_N(_03541_));
 sg13g2_nand2_1 _10089_ (.Y(_03543_),
    .A(_03540_),
    .B(_03542_));
 sg13g2_a21oi_1 _10090_ (.A1(net4237),
    .A2(net4289),
    .Y(_03544_),
    .B1(net3862));
 sg13g2_a21oi_1 _10091_ (.A1(_03540_),
    .A2(_03544_),
    .Y(_03545_),
    .B1(net4302));
 sg13g2_a21oi_1 _10092_ (.A1(net4153),
    .A2(net4045),
    .Y(_03546_),
    .B1(_03541_));
 sg13g2_o21ai_1 _10093_ (.B1(net3796),
    .Y(_03547_),
    .A1(net4451),
    .A2(_03546_));
 sg13g2_a21oi_1 _10094_ (.A1(net4322),
    .A2(_01802_),
    .Y(_03548_),
    .B1(_03536_));
 sg13g2_a22oi_1 _10095_ (.Y(_03549_),
    .B1(_03543_),
    .B2(net3805),
    .A2(_01802_),
    .A1(net4334));
 sg13g2_o21ai_1 _10096_ (.B1(_03549_),
    .Y(_03550_),
    .A1(net4334),
    .A2(_01186_));
 sg13g2_nor2_1 _10097_ (.A(_01802_),
    .B(_03545_),
    .Y(_03551_));
 sg13g2_a221oi_1 _10098_ (.B2(_03294_),
    .C1(_03551_),
    .B1(_03548_),
    .A1(_03540_),
    .Y(_03552_),
    .A2(_03547_));
 sg13g2_a21o_1 _10099_ (.A2(_03552_),
    .A1(_03550_),
    .B1(net3945),
    .X(_03553_));
 sg13g2_nand2b_1 _10100_ (.Y(_03554_),
    .B(net4067),
    .A_N(_00186_));
 sg13g2_o21ai_1 _10101_ (.B1(_03554_),
    .Y(_03555_),
    .A1(_00188_),
    .A2(net4149));
 sg13g2_a221oi_1 _10102_ (.B2(\cpu.registers[5][10] ),
    .C1(_03555_),
    .B1(net3983),
    .A1(\cpu.registers[3][10] ),
    .Y(_03556_),
    .A2(net3996));
 sg13g2_o21ai_1 _10103_ (.B1(net4076),
    .Y(_03557_),
    .A1(_00187_),
    .A2(net3997));
 sg13g2_a221oi_1 _10104_ (.B2(_00973_),
    .C1(_03557_),
    .B1(_02133_),
    .A1(\cpu.registers[2][10] ),
    .Y(_03558_),
    .A2(net3988));
 sg13g2_a22oi_1 _10105_ (.Y(_03559_),
    .B1(_03556_),
    .B2(_03558_),
    .A2(_02236_),
    .A1(net4068));
 sg13g2_a21oi_1 _10106_ (.A1(net3945),
    .A2(_03559_),
    .Y(_03560_),
    .B1(net3640));
 sg13g2_a22oi_1 _10107_ (.Y(_00678_),
    .B1(_03553_),
    .B2(_03560_),
    .A2(net3640),
    .A1(_01156_));
 sg13g2_o21ai_1 _10108_ (.B1(_03294_),
    .Y(_03561_),
    .A1(net4323),
    .A2(_01189_));
 sg13g2_nor2_1 _10109_ (.A(net4067),
    .B(_02243_),
    .Y(_03562_));
 sg13g2_nand2_1 _10110_ (.Y(_03563_),
    .A(net4323),
    .B(net4284));
 sg13g2_o21ai_1 _10111_ (.B1(_03563_),
    .Y(_03564_),
    .A1(net4323),
    .A2(_01189_));
 sg13g2_o21ai_1 _10112_ (.B1(net3802),
    .Y(_03565_),
    .A1(net4062),
    .A2(_03564_));
 sg13g2_o21ai_1 _10113_ (.B1(net4314),
    .Y(_03566_),
    .A1(_03562_),
    .A2(_03565_));
 sg13g2_inv_1 _10114_ (.Y(_03567_),
    .A(_03566_));
 sg13g2_nor2_1 _10115_ (.A(net4284),
    .B(net3863),
    .Y(_03568_));
 sg13g2_a21oi_1 _10116_ (.A1(net4237),
    .A2(net4284),
    .Y(_03569_),
    .B1(net3863));
 sg13g2_nor2_1 _10117_ (.A(net4077),
    .B(_03564_),
    .Y(_03570_));
 sg13g2_nor2b_1 _10118_ (.A(_03570_),
    .B_N(net3861),
    .Y(_03571_));
 sg13g2_o21ai_1 _10119_ (.B1(net3805),
    .Y(_03572_),
    .A1(_03566_),
    .A2(_03571_));
 sg13g2_nand2_1 _10120_ (.Y(_03573_),
    .A(net4202),
    .B(_00193_));
 sg13g2_a221oi_1 _10121_ (.B2(_03573_),
    .C1(net4302),
    .B1(_03572_),
    .A1(_03567_),
    .Y(_03574_),
    .A2(_03569_));
 sg13g2_a21oi_1 _10122_ (.A1(_03561_),
    .A2(_03574_),
    .Y(_03575_),
    .B1(_01825_));
 sg13g2_and3_1 _10123_ (.X(_03576_),
    .A(net4203),
    .B(_01189_),
    .C(_03572_));
 sg13g2_o21ai_1 _10124_ (.B1(net4237),
    .Y(_03577_),
    .A1(_03568_),
    .A2(_03570_));
 sg13g2_a21oi_1 _10125_ (.A1(net3796),
    .A2(_03577_),
    .Y(_03578_),
    .B1(_03566_));
 sg13g2_nor2_1 _10126_ (.A(net4323),
    .B(_03561_),
    .Y(_03579_));
 sg13g2_or4_1 _10127_ (.A(_03575_),
    .B(_03576_),
    .C(_03578_),
    .D(_03579_),
    .X(_03580_));
 sg13g2_nand2_1 _10128_ (.Y(_03581_),
    .A(net4069),
    .B(_02243_));
 sg13g2_nand2_1 _10129_ (.Y(_03582_),
    .A(\cpu.registers[2][11] ),
    .B(net3988));
 sg13g2_o21ai_1 _10130_ (.B1(_03582_),
    .Y(_03583_),
    .A1(_00191_),
    .A2(net3997));
 sg13g2_a221oi_1 _10131_ (.B2(_00981_),
    .C1(_03583_),
    .B1(_02133_),
    .A1(_01187_),
    .Y(_03584_),
    .A2(_01363_));
 sg13g2_o21ai_1 _10132_ (.B1(net4076),
    .Y(_03585_),
    .A1(_00190_),
    .A2(net4062));
 sg13g2_a221oi_1 _10133_ (.B2(\cpu.registers[5][11] ),
    .C1(_03585_),
    .B1(net3983),
    .A1(\cpu.registers[3][11] ),
    .Y(_03586_),
    .A2(net3996));
 sg13g2_a21oi_1 _10134_ (.A1(_03584_),
    .A2(_03586_),
    .Y(_03587_),
    .B1(net3943));
 sg13g2_a221oi_1 _10135_ (.B2(_03587_),
    .C1(net3641),
    .B1(_03581_),
    .A1(net3943),
    .Y(_03588_),
    .A2(_03580_));
 sg13g2_a21oi_1 _10136_ (.A1(_01158_),
    .A2(net3641),
    .Y(_00679_),
    .B1(_03588_));
 sg13g2_nor2_1 _10137_ (.A(net4067),
    .B(_02250_),
    .Y(_03589_));
 sg13g2_nor2b_1 _10138_ (.A(net4323),
    .B_N(_00197_),
    .Y(_03590_));
 sg13g2_a21o_1 _10139_ (.A2(net4280),
    .A1(net4325),
    .B1(_03590_),
    .X(_03591_));
 sg13g2_o21ai_1 _10140_ (.B1(net3802),
    .Y(_03592_),
    .A1(net4062),
    .A2(_03591_));
 sg13g2_o21ai_1 _10141_ (.B1(net4318),
    .Y(_03593_),
    .A1(_03589_),
    .A2(_03592_));
 sg13g2_o21ai_1 _10142_ (.B1(net3861),
    .Y(_03594_),
    .A1(net4077),
    .A2(_03591_));
 sg13g2_nand2b_1 _10143_ (.Y(_03595_),
    .B(_03594_),
    .A_N(_03593_));
 sg13g2_a22oi_1 _10144_ (.Y(_03596_),
    .B1(net3805),
    .B2(_03595_),
    .A2(_00197_),
    .A1(net4203));
 sg13g2_nor2_1 _10145_ (.A(net3795),
    .B(_03590_),
    .Y(_03597_));
 sg13g2_nand2b_1 _10146_ (.Y(_03598_),
    .B(net4049),
    .A_N(net4280));
 sg13g2_a21oi_1 _10147_ (.A1(_01249_),
    .A2(_03598_),
    .Y(_03599_),
    .B1(_03593_));
 sg13g2_or3_1 _10148_ (.A(net4302),
    .B(_03597_),
    .C(_03599_),
    .X(_03600_));
 sg13g2_o21ai_1 _10149_ (.B1(_01851_),
    .Y(_03601_),
    .A1(_03596_),
    .A2(_03600_));
 sg13g2_o21ai_1 _10150_ (.B1(_03598_),
    .Y(_03602_),
    .A1(net4077),
    .A2(_03591_));
 sg13g2_a21oi_1 _10151_ (.A1(net4238),
    .A2(_03602_),
    .Y(_03603_),
    .B1(net3801));
 sg13g2_nor2_1 _10152_ (.A(_03593_),
    .B(_03603_),
    .Y(_03604_));
 sg13g2_a221oi_1 _10153_ (.B2(net4242),
    .C1(_03604_),
    .B1(_03597_),
    .A1(net4203),
    .Y(_03605_),
    .A2(_03596_));
 sg13g2_a21oi_1 _10154_ (.A1(_03601_),
    .A2(_03605_),
    .Y(_03606_),
    .B1(net3946));
 sg13g2_nand2_1 _10155_ (.Y(_03607_),
    .A(\cpu.registers[2][12] ),
    .B(net3988));
 sg13g2_o21ai_1 _10156_ (.B1(_03607_),
    .Y(_03608_),
    .A1(_00195_),
    .A2(net3997));
 sg13g2_a221oi_1 _10157_ (.B2(_00989_),
    .C1(_03608_),
    .B1(_02133_),
    .A1(_01190_),
    .Y(_03609_),
    .A2(_01363_));
 sg13g2_o21ai_1 _10158_ (.B1(net4076),
    .Y(_03610_),
    .A1(_00194_),
    .A2(net4062));
 sg13g2_a221oi_1 _10159_ (.B2(\cpu.registers[5][12] ),
    .C1(_03610_),
    .B1(net3983),
    .A1(\cpu.registers[3][12] ),
    .Y(_03611_),
    .A2(net3996));
 sg13g2_a221oi_1 _10160_ (.B2(_03611_),
    .C1(net3943),
    .B1(_03609_),
    .A1(net4069),
    .Y(_03612_),
    .A2(_02250_));
 sg13g2_nor3_1 _10161_ (.A(_03272_),
    .B(_03606_),
    .C(_03612_),
    .Y(_03613_));
 sg13g2_a21oi_1 _10162_ (.A1(_01160_),
    .A2(net3641),
    .Y(_00680_),
    .B1(_03613_));
 sg13g2_nor2b_1 _10163_ (.A(net4324),
    .B_N(_00202_),
    .Y(_03614_));
 sg13g2_a21o_1 _10164_ (.A2(_00143_),
    .A1(net4322),
    .B1(_03614_),
    .X(_03615_));
 sg13g2_nor2_1 _10165_ (.A(net4060),
    .B(_03615_),
    .Y(_03616_));
 sg13g2_a21oi_1 _10166_ (.A1(net4060),
    .A2(_02803_),
    .Y(_03617_),
    .B1(_03616_));
 sg13g2_a21oi_1 _10167_ (.A1(net3801),
    .A2(_03617_),
    .Y(_03618_),
    .B1(net4253));
 sg13g2_nor2_1 _10168_ (.A(net4077),
    .B(_03615_),
    .Y(_03619_));
 sg13g2_nand2b_1 _10169_ (.Y(_03620_),
    .B(net3861),
    .A_N(_03619_));
 sg13g2_a21oi_1 _10170_ (.A1(_03618_),
    .A2(_03620_),
    .Y(_03621_),
    .B1(_01290_));
 sg13g2_a21oi_1 _10171_ (.A1(net4238),
    .A2(_00143_),
    .Y(_03622_),
    .B1(net3862));
 sg13g2_a21oi_1 _10172_ (.A1(_03618_),
    .A2(_03622_),
    .Y(_03623_),
    .B1(net4302));
 sg13g2_a21oi_1 _10173_ (.A1(net4152),
    .A2(net4045),
    .Y(_03624_),
    .B1(_03619_));
 sg13g2_o21ai_1 _10174_ (.B1(net3796),
    .Y(_03625_),
    .A1(net4451),
    .A2(_03624_));
 sg13g2_nand2_1 _10175_ (.Y(_03626_),
    .A(_03618_),
    .B(_03625_));
 sg13g2_a21oi_1 _10176_ (.A1(net4324),
    .A2(_01870_),
    .Y(_03627_),
    .B1(_03614_));
 sg13g2_a21o_1 _10177_ (.A2(_01870_),
    .A1(net4334),
    .B1(_03621_),
    .X(_03628_));
 sg13g2_a21oi_1 _10178_ (.A1(net4202),
    .A2(_00202_),
    .Y(_03629_),
    .B1(_03628_));
 sg13g2_o21ai_1 _10179_ (.B1(_03626_),
    .Y(_03630_),
    .A1(_01870_),
    .A2(_03623_));
 sg13g2_a21o_1 _10180_ (.A2(_03627_),
    .A1(_03294_),
    .B1(_03630_),
    .X(_03631_));
 sg13g2_o21ai_1 _10181_ (.B1(net3943),
    .Y(_03632_),
    .A1(_03629_),
    .A2(_03631_));
 sg13g2_nor2_1 _10182_ (.A(_00046_),
    .B(net3986),
    .Y(_03633_));
 sg13g2_nor2_1 _10183_ (.A(_00200_),
    .B(net4149),
    .Y(_03634_));
 sg13g2_nand2_1 _10184_ (.Y(_03635_),
    .A(\cpu.registers[2][13] ),
    .B(net3988));
 sg13g2_o21ai_1 _10185_ (.B1(_03635_),
    .Y(_03636_),
    .A1(_00199_),
    .A2(net3997));
 sg13g2_nor3_1 _10186_ (.A(_03633_),
    .B(_03634_),
    .C(_03636_),
    .Y(_03637_));
 sg13g2_o21ai_1 _10187_ (.B1(net4076),
    .Y(_03638_),
    .A1(_00198_),
    .A2(net4061));
 sg13g2_a221oi_1 _10188_ (.B2(\cpu.registers[5][13] ),
    .C1(_03638_),
    .B1(net3983),
    .A1(\cpu.registers[3][13] ),
    .Y(_03639_),
    .A2(net3996));
 sg13g2_a22oi_1 _10189_ (.Y(_03640_),
    .B1(_03637_),
    .B2(_03639_),
    .A2(_02802_),
    .A1(net4068));
 sg13g2_a21oi_1 _10190_ (.A1(net3945),
    .A2(_03640_),
    .Y(_03641_),
    .B1(net3641));
 sg13g2_a22oi_1 _10191_ (.Y(_00681_),
    .B1(_03632_),
    .B2(_03641_),
    .A2(net3641),
    .A1(_01162_));
 sg13g2_nand2_1 _10192_ (.Y(_03642_),
    .A(net4242),
    .B(_00206_));
 sg13g2_o21ai_1 _10193_ (.B1(_03642_),
    .Y(_03643_),
    .A1(net4242),
    .A2(net4151));
 sg13g2_o21ai_1 _10194_ (.B1(net3801),
    .Y(_03644_),
    .A1(net4060),
    .A2(_03643_));
 sg13g2_a21oi_1 _10195_ (.A1(net4060),
    .A2(_02812_),
    .Y(_03645_),
    .B1(_03644_));
 sg13g2_nor2_1 _10196_ (.A(net4253),
    .B(_03645_),
    .Y(_03646_));
 sg13g2_or2_1 _10197_ (.X(_03647_),
    .B(_03643_),
    .A(net4077));
 sg13g2_nand2_1 _10198_ (.Y(_03648_),
    .A(net3861),
    .B(_03647_));
 sg13g2_nand2_1 _10199_ (.Y(_03649_),
    .A(_03646_),
    .B(_03648_));
 sg13g2_a22oi_1 _10200_ (.Y(_03650_),
    .B1(net3805),
    .B2(_03649_),
    .A2(_00206_),
    .A1(net4202));
 sg13g2_a21oi_1 _10201_ (.A1(net4237),
    .A2(net4274),
    .Y(_03651_),
    .B1(net3863));
 sg13g2_a21oi_1 _10202_ (.A1(_03646_),
    .A2(_03651_),
    .Y(_03652_),
    .B1(net4302));
 sg13g2_o21ai_1 _10203_ (.B1(_03647_),
    .Y(_03653_),
    .A1(net4274),
    .A2(net3862));
 sg13g2_a21oi_1 _10204_ (.A1(net4237),
    .A2(_03653_),
    .Y(_03654_),
    .B1(net3801));
 sg13g2_nand2b_1 _10205_ (.Y(_03655_),
    .B(_03646_),
    .A_N(_03654_));
 sg13g2_a21oi_1 _10206_ (.A1(net4322),
    .A2(_01891_),
    .Y(_03656_),
    .B1(net3795));
 sg13g2_nand2_1 _10207_ (.Y(_03657_),
    .A(net4334),
    .B(_01891_));
 sg13g2_o21ai_1 _10208_ (.B1(_03655_),
    .Y(_03658_),
    .A1(_01891_),
    .A2(_03652_));
 sg13g2_a221oi_1 _10209_ (.B2(_03650_),
    .C1(_03658_),
    .B1(_03657_),
    .A1(_03642_),
    .Y(_03659_),
    .A2(_03656_));
 sg13g2_or2_1 _10210_ (.X(_03660_),
    .B(_03659_),
    .A(net3945));
 sg13g2_nor2_1 _10211_ (.A(net4076),
    .B(_02812_),
    .Y(_03661_));
 sg13g2_nor2_1 _10212_ (.A(_00205_),
    .B(net4149),
    .Y(_03662_));
 sg13g2_nand2_1 _10213_ (.Y(_03663_),
    .A(\cpu.registers[5][14] ),
    .B(net3983));
 sg13g2_o21ai_1 _10214_ (.B1(net4076),
    .Y(_03664_),
    .A1(_00047_),
    .A2(net3986));
 sg13g2_nor2_1 _10215_ (.A(_00203_),
    .B(net4061),
    .Y(_03665_));
 sg13g2_o21ai_1 _10216_ (.B1(_03663_),
    .Y(_03666_),
    .A1(_00204_),
    .A2(net3997));
 sg13g2_a221oi_1 _10217_ (.B2(\cpu.registers[2][14] ),
    .C1(_03666_),
    .B1(net3988),
    .A1(\cpu.registers[3][14] ),
    .Y(_03667_),
    .A2(net3996));
 sg13g2_nor3_1 _10218_ (.A(_03662_),
    .B(_03664_),
    .C(_03665_),
    .Y(_03668_));
 sg13g2_a21oi_1 _10219_ (.A1(_03667_),
    .A2(_03668_),
    .Y(_03669_),
    .B1(_03661_));
 sg13g2_a21oi_1 _10220_ (.A1(net3945),
    .A2(_03669_),
    .Y(_03670_),
    .B1(net3640));
 sg13g2_a22oi_1 _10221_ (.Y(_00682_),
    .B1(_03660_),
    .B2(_03670_),
    .A2(net3640),
    .A1(_01163_));
 sg13g2_a22oi_1 _10222_ (.Y(_03671_),
    .B1(net3805),
    .B2(_03300_),
    .A2(_00210_),
    .A1(net4202));
 sg13g2_nor2_1 _10223_ (.A(_03288_),
    .B(net3795),
    .Y(_03672_));
 sg13g2_nor3_1 _10224_ (.A(_03303_),
    .B(_03671_),
    .C(_03672_),
    .Y(_03673_));
 sg13g2_nor3_1 _10225_ (.A(net4451),
    .B(net4080),
    .C(_03289_),
    .Y(_03674_));
 sg13g2_o21ai_1 _10226_ (.B1(net3797),
    .Y(_03675_),
    .A1(net4271),
    .A2(_01247_));
 sg13g2_nor2_1 _10227_ (.A(_03674_),
    .B(_03675_),
    .Y(_03676_));
 sg13g2_nor3_1 _10228_ (.A(net4253),
    .B(_03291_),
    .C(_03676_),
    .Y(_03677_));
 sg13g2_a221oi_1 _10229_ (.B2(net4242),
    .C1(_03677_),
    .B1(_03672_),
    .A1(net4202),
    .Y(_03678_),
    .A2(_03671_));
 sg13g2_o21ai_1 _10230_ (.B1(_03678_),
    .Y(_03679_),
    .A1(_01911_),
    .A2(_03673_));
 sg13g2_nand2b_1 _10231_ (.Y(_03680_),
    .B(net4068),
    .A_N(_02821_));
 sg13g2_nor2_1 _10232_ (.A(_00209_),
    .B(net4149),
    .Y(_03681_));
 sg13g2_nand2_1 _10233_ (.Y(_03682_),
    .A(\cpu.registers[5][15] ),
    .B(net3983));
 sg13g2_o21ai_1 _10234_ (.B1(net4076),
    .Y(_03683_),
    .A1(_00048_),
    .A2(net3986));
 sg13g2_nor2_1 _10235_ (.A(_00207_),
    .B(net4061),
    .Y(_03684_));
 sg13g2_o21ai_1 _10236_ (.B1(_03682_),
    .Y(_03685_),
    .A1(_00208_),
    .A2(net3997));
 sg13g2_a221oi_1 _10237_ (.B2(\cpu.registers[2][15] ),
    .C1(_03685_),
    .B1(net3988),
    .A1(\cpu.registers[3][15] ),
    .Y(_03686_),
    .A2(net3996));
 sg13g2_nor3_1 _10238_ (.A(_03681_),
    .B(_03683_),
    .C(_03684_),
    .Y(_03687_));
 sg13g2_a21oi_1 _10239_ (.A1(_03686_),
    .A2(_03687_),
    .Y(_03688_),
    .B1(net3943));
 sg13g2_a221oi_1 _10240_ (.B2(_03688_),
    .C1(net3640),
    .B1(_03680_),
    .A1(net3943),
    .Y(_03689_),
    .A2(_03679_));
 sg13g2_a21oi_1 _10241_ (.A1(_01165_),
    .A2(net3640),
    .Y(_00683_),
    .B1(_03689_));
 sg13g2_and2_1 _10242_ (.A(_01301_),
    .B(_01307_),
    .X(_03690_));
 sg13g2_nor2b_2 _10243_ (.A(\memory_controller.state[4] ),
    .B_N(_03690_),
    .Y(_03691_));
 sg13g2_nand2b_2 _10244_ (.Y(_03692_),
    .B(_03690_),
    .A_N(net4332));
 sg13g2_nand2_1 _10245_ (.Y(_03693_),
    .A(net182),
    .B(_03691_));
 sg13g2_nand2b_1 _10246_ (.Y(_00684_),
    .B(_03693_),
    .A_N(net192));
 sg13g2_nand2_1 _10247_ (.Y(_03694_),
    .A(net4391),
    .B(net4012));
 sg13g2_nand2_1 _10248_ (.Y(_03695_),
    .A(_00227_),
    .B(net3843));
 sg13g2_o21ai_1 _10249_ (.B1(_03695_),
    .Y(_03696_),
    .A1(_01170_),
    .A2(net3843));
 sg13g2_nand2_1 _10250_ (.Y(_03697_),
    .A(_01420_),
    .B(net3842));
 sg13g2_nand2_1 _10251_ (.Y(_03698_),
    .A(net4445),
    .B(_01336_));
 sg13g2_a22oi_1 _10252_ (.Y(_03699_),
    .B1(_03698_),
    .B2(_01927_),
    .A2(_02138_),
    .A1(_01926_));
 sg13g2_nand4_1 _10253_ (.B(_01432_),
    .C(_03697_),
    .A(_01423_),
    .Y(_03700_),
    .D(_03699_));
 sg13g2_o21ai_1 _10254_ (.B1(_01443_),
    .Y(_03701_),
    .A1(_01410_),
    .A2(_03696_));
 sg13g2_mux2_1 _10255_ (.A0(_03701_),
    .A1(net746),
    .S(net3601),
    .X(_00685_));
 sg13g2_mux2_1 _10256_ (.A0(net4361),
    .A1(_00228_),
    .S(net3844),
    .X(_03702_));
 sg13g2_nor2_1 _10257_ (.A(_01451_),
    .B(_03702_),
    .Y(_03703_));
 sg13g2_nor3_1 _10258_ (.A(_01448_),
    .B(net3601),
    .C(_03703_),
    .Y(_03704_));
 sg13g2_a21oi_1 _10259_ (.A1(_00910_),
    .A2(net3601),
    .Y(_00686_),
    .B1(_03704_));
 sg13g2_mux2_1 _10260_ (.A0(net4353),
    .A1(_00229_),
    .S(net3843),
    .X(_03705_));
 sg13g2_nor2_1 _10261_ (.A(_01477_),
    .B(_03705_),
    .Y(_03706_));
 sg13g2_nor3_1 _10262_ (.A(_01481_),
    .B(net3601),
    .C(_03706_),
    .Y(_03707_));
 sg13g2_a21oi_1 _10263_ (.A1(_00915_),
    .A2(net3601),
    .Y(_00687_),
    .B1(_03707_));
 sg13g2_nand2b_1 _10264_ (.Y(_03708_),
    .B(net3844),
    .A_N(_00230_));
 sg13g2_o21ai_1 _10265_ (.B1(_03708_),
    .Y(_03709_),
    .A1(net4351),
    .A2(net3843));
 sg13g2_o21ai_1 _10266_ (.B1(_01511_),
    .Y(_03710_),
    .A1(net3868),
    .A2(_03709_));
 sg13g2_a21oi_1 _10267_ (.A1(net4300),
    .A2(_03709_),
    .Y(_03711_),
    .B1(_01516_));
 sg13g2_nor2b_1 _10268_ (.A(net3600),
    .B_N(_03711_),
    .Y(_03712_));
 sg13g2_a22oi_1 _10269_ (.Y(_00688_),
    .B1(_03710_),
    .B2(_03712_),
    .A2(net3600),
    .A1(_00923_));
 sg13g2_nand2_1 _10270_ (.Y(_03713_),
    .A(_00231_),
    .B(net3843));
 sg13g2_o21ai_1 _10271_ (.B1(_03713_),
    .Y(_03714_),
    .A1(net4156),
    .A2(net3844));
 sg13g2_a21o_1 _10272_ (.A2(_03714_),
    .A1(net4057),
    .B1(_01552_),
    .X(_03715_));
 sg13g2_nor2_1 _10273_ (.A(net4235),
    .B(_03714_),
    .Y(_03716_));
 sg13g2_nor3_1 _10274_ (.A(_01556_),
    .B(net3600),
    .C(_03716_),
    .Y(_03717_));
 sg13g2_a22oi_1 _10275_ (.Y(_00689_),
    .B1(_03715_),
    .B2(_03717_),
    .A2(net3600),
    .A1(_00930_));
 sg13g2_mux2_1 _10276_ (.A0(net4345),
    .A1(_00232_),
    .S(net3844),
    .X(_03718_));
 sg13g2_a21oi_1 _10277_ (.A1(net4054),
    .A2(_03718_),
    .Y(_03719_),
    .B1(net4260));
 sg13g2_nor2_1 _10278_ (.A(net4234),
    .B(_03718_),
    .Y(_03720_));
 sg13g2_a21oi_1 _10279_ (.A1(_01596_),
    .A2(_03719_),
    .Y(_03721_),
    .B1(_03720_));
 sg13g2_nor2_1 _10280_ (.A(_01601_),
    .B(net3600),
    .Y(_03722_));
 sg13g2_a22oi_1 _10281_ (.Y(_00690_),
    .B1(_03721_),
    .B2(_03722_),
    .A2(net3600),
    .A1(_00937_));
 sg13g2_nand2_1 _10282_ (.Y(_03723_),
    .A(_00233_),
    .B(net3843));
 sg13g2_o21ai_1 _10283_ (.B1(_03723_),
    .Y(_03724_),
    .A1(net4155),
    .A2(net3843));
 sg13g2_a21oi_1 _10284_ (.A1(net4056),
    .A2(_03724_),
    .Y(_03725_),
    .B1(net4262));
 sg13g2_nand2_1 _10285_ (.Y(_03726_),
    .A(_01649_),
    .B(_03725_));
 sg13g2_o21ai_1 _10286_ (.B1(_01654_),
    .Y(_03727_),
    .A1(net4235),
    .A2(_03724_));
 sg13g2_nor2_1 _10287_ (.A(net3600),
    .B(_03727_),
    .Y(_03728_));
 sg13g2_a22oi_1 _10288_ (.Y(_00691_),
    .B1(_03726_),
    .B2(_03728_),
    .A2(net3600),
    .A1(_00944_));
 sg13g2_mux2_1 _10289_ (.A0(net4338),
    .A1(_00234_),
    .S(net3843),
    .X(_03729_));
 sg13g2_a21oi_1 _10290_ (.A1(net4052),
    .A2(_03729_),
    .Y(_03730_),
    .B1(net4259));
 sg13g2_nand2_1 _10291_ (.Y(_03731_),
    .A(_01707_),
    .B(_03730_));
 sg13g2_nor2_1 _10292_ (.A(net4232),
    .B(_03729_),
    .Y(_03732_));
 sg13g2_nor3_1 _10293_ (.A(_01713_),
    .B(net3601),
    .C(_03732_),
    .Y(_03733_));
 sg13g2_a22oi_1 _10294_ (.Y(_00692_),
    .B1(_03731_),
    .B2(_03733_),
    .A2(net3601),
    .A1(_00952_));
 sg13g2_mux2_1 _10295_ (.A0(net4297),
    .A1(_00235_),
    .S(net3841),
    .X(_03734_));
 sg13g2_a21oi_1 _10296_ (.A1(net4044),
    .A2(_03734_),
    .Y(_03735_),
    .B1(net4251));
 sg13g2_nor2_1 _10297_ (.A(net4225),
    .B(_03734_),
    .Y(_03736_));
 sg13g2_a21oi_1 _10298_ (.A1(_01756_),
    .A2(_03735_),
    .Y(_03737_),
    .B1(_03736_));
 sg13g2_nor2_1 _10299_ (.A(_01761_),
    .B(net3599),
    .Y(_03738_));
 sg13g2_a22oi_1 _10300_ (.Y(_00693_),
    .B1(_03737_),
    .B2(_03738_),
    .A2(net3599),
    .A1(_00959_));
 sg13g2_nand2_1 _10301_ (.Y(_03739_),
    .A(_00236_),
    .B(net3842));
 sg13g2_o21ai_1 _10302_ (.B1(_03739_),
    .Y(_03740_),
    .A1(net4154),
    .A2(net3842));
 sg13g2_a21oi_1 _10303_ (.A1(net4047),
    .A2(_03740_),
    .Y(_03741_),
    .B1(net4256));
 sg13g2_nand2_1 _10304_ (.Y(_03742_),
    .A(_01780_),
    .B(_03741_));
 sg13g2_nor2_1 _10305_ (.A(net4228),
    .B(_03740_),
    .Y(_03743_));
 sg13g2_nor3_1 _10306_ (.A(_01786_),
    .B(net3599),
    .C(_03743_),
    .Y(_03744_));
 sg13g2_a22oi_1 _10307_ (.Y(_00694_),
    .B1(_03742_),
    .B2(_03744_),
    .A2(net3599),
    .A1(_00967_));
 sg13g2_nand2_1 _10308_ (.Y(_03745_),
    .A(_00237_),
    .B(net3841));
 sg13g2_o21ai_1 _10309_ (.B1(_03745_),
    .Y(_03746_),
    .A1(net4153),
    .A2(net3841));
 sg13g2_a21oi_1 _10310_ (.A1(net4043),
    .A2(_03746_),
    .Y(_03747_),
    .B1(net4246));
 sg13g2_nor2_1 _10311_ (.A(net4224),
    .B(_03746_),
    .Y(_03748_));
 sg13g2_a21oi_1 _10312_ (.A1(_01803_),
    .A2(_03747_),
    .Y(_03749_),
    .B1(_03748_));
 sg13g2_nor2_1 _10313_ (.A(_01809_),
    .B(net3598),
    .Y(_03750_));
 sg13g2_a22oi_1 _10314_ (.Y(_00695_),
    .B1(_03749_),
    .B2(_03750_),
    .A2(net3598),
    .A1(_00975_));
 sg13g2_mux2_1 _10315_ (.A0(net4284),
    .A1(_00238_),
    .S(net3842),
    .X(_03751_));
 sg13g2_a21oi_1 _10316_ (.A1(net4046),
    .A2(_03751_),
    .Y(_03752_),
    .B1(net4252));
 sg13g2_nand2_1 _10317_ (.Y(_03753_),
    .A(_01826_),
    .B(_03752_));
 sg13g2_nor2_1 _10318_ (.A(net4229),
    .B(_03751_),
    .Y(_03754_));
 sg13g2_nor3_1 _10319_ (.A(_01831_),
    .B(_03700_),
    .C(_03754_),
    .Y(_03755_));
 sg13g2_a22oi_1 _10320_ (.Y(_00696_),
    .B1(_03753_),
    .B2(_03755_),
    .A2(net3599),
    .A1(_00983_));
 sg13g2_mux2_1 _10321_ (.A0(net4280),
    .A1(_00239_),
    .S(net3842),
    .X(_03756_));
 sg13g2_a21oi_1 _10322_ (.A1(net4047),
    .A2(_03756_),
    .Y(_03757_),
    .B1(net4255));
 sg13g2_nor2_1 _10323_ (.A(net4227),
    .B(_03756_),
    .Y(_03758_));
 sg13g2_a21oi_1 _10324_ (.A1(_01852_),
    .A2(_03757_),
    .Y(_03759_),
    .B1(_03758_));
 sg13g2_nor2_1 _10325_ (.A(_01857_),
    .B(net3599),
    .Y(_03760_));
 sg13g2_a22oi_1 _10326_ (.Y(_00697_),
    .B1(_03759_),
    .B2(_03760_),
    .A2(net3599),
    .A1(_00991_));
 sg13g2_nand2_1 _10327_ (.Y(_03761_),
    .A(_00240_),
    .B(net3841));
 sg13g2_o21ai_1 _10328_ (.B1(_03761_),
    .Y(_03762_),
    .A1(net4152),
    .A2(net3841));
 sg13g2_a21oi_1 _10329_ (.A1(net4041),
    .A2(_03762_),
    .Y(_03763_),
    .B1(net4247));
 sg13g2_nand2_1 _10330_ (.Y(_03764_),
    .A(_01871_),
    .B(_03763_));
 sg13g2_nor2_1 _10331_ (.A(net4222),
    .B(_03762_),
    .Y(_03765_));
 sg13g2_nor3_1 _10332_ (.A(_01877_),
    .B(net3598),
    .C(_03765_),
    .Y(_03766_));
 sg13g2_a22oi_1 _10333_ (.Y(_00698_),
    .B1(_03764_),
    .B2(_03766_),
    .A2(net3598),
    .A1(_01113_));
 sg13g2_nand2_1 _10334_ (.Y(_03767_),
    .A(_00241_),
    .B(net3841));
 sg13g2_o21ai_1 _10335_ (.B1(_03767_),
    .Y(_03768_),
    .A1(net4151),
    .A2(net3841));
 sg13g2_a21oi_1 _10336_ (.A1(net4040),
    .A2(_03768_),
    .Y(_03769_),
    .B1(net4246));
 sg13g2_nand2_1 _10337_ (.Y(_03770_),
    .A(_01892_),
    .B(_03769_));
 sg13g2_nor2_1 _10338_ (.A(net4221),
    .B(_03768_),
    .Y(_03771_));
 sg13g2_nor3_1 _10339_ (.A(_01898_),
    .B(net3598),
    .C(_03771_),
    .Y(_03772_));
 sg13g2_a22oi_1 _10340_ (.Y(_00699_),
    .B1(_03770_),
    .B2(_03772_),
    .A2(net3598),
    .A1(_01128_));
 sg13g2_mux2_1 _10341_ (.A0(net4268),
    .A1(_00242_),
    .S(net3841),
    .X(_03773_));
 sg13g2_a21oi_1 _10342_ (.A1(net4041),
    .A2(_03773_),
    .Y(_03774_),
    .B1(net4248));
 sg13g2_nand2_1 _10343_ (.Y(_03775_),
    .A(_01912_),
    .B(_03774_));
 sg13g2_nor2_1 _10344_ (.A(net4222),
    .B(_03773_),
    .Y(_03776_));
 sg13g2_nor3_1 _10345_ (.A(_01917_),
    .B(net3598),
    .C(_03776_),
    .Y(_03777_));
 sg13g2_a22oi_1 _10346_ (.Y(_00700_),
    .B1(_03775_),
    .B2(_03777_),
    .A2(net3598),
    .A1(_01141_));
 sg13g2_nor3_1 _10347_ (.A(net4215),
    .B(net4207),
    .C(net4396),
    .Y(_03778_));
 sg13g2_mux2_1 _10348_ (.A0(_00146_),
    .A1(net4365),
    .S(net3940),
    .X(_03779_));
 sg13g2_nand2b_1 _10349_ (.Y(_03780_),
    .B(_01420_),
    .A_N(net3940));
 sg13g2_nand2_1 _10350_ (.Y(_03781_),
    .A(net4445),
    .B(_01433_));
 sg13g2_a22oi_1 _10351_ (.Y(_03782_),
    .B1(_01927_),
    .B2(_03781_),
    .A2(_01436_),
    .A1(net4066));
 sg13g2_nand4_1 _10352_ (.B(_01432_),
    .C(_03780_),
    .A(_01423_),
    .Y(_03783_),
    .D(_03782_));
 sg13g2_o21ai_1 _10353_ (.B1(_01443_),
    .Y(_03784_),
    .A1(_01410_),
    .A2(_03779_));
 sg13g2_mux2_1 _10354_ (.A0(_03784_),
    .A1(net308),
    .S(net3597),
    .X(_00701_));
 sg13g2_mux2_1 _10355_ (.A0(_00150_),
    .A1(net4362),
    .S(net3941),
    .X(_03785_));
 sg13g2_nor2_1 _10356_ (.A(_01451_),
    .B(_03785_),
    .Y(_03786_));
 sg13g2_nor3_1 _10357_ (.A(_01448_),
    .B(net3595),
    .C(_03786_),
    .Y(_03787_));
 sg13g2_a21oi_1 _10358_ (.A1(_00909_),
    .A2(net3596),
    .Y(_00702_),
    .B1(_03787_));
 sg13g2_nor2b_1 _10359_ (.A(net3940),
    .B_N(_00154_),
    .Y(_03788_));
 sg13g2_a221oi_1 _10360_ (.B2(net4353),
    .C1(_03788_),
    .B1(net3940),
    .A1(net4231),
    .Y(_03789_),
    .A2(_01476_));
 sg13g2_nor3_1 _10361_ (.A(_01481_),
    .B(net3597),
    .C(_03789_),
    .Y(_03790_));
 sg13g2_a21oi_1 _10362_ (.A1(_00914_),
    .A2(net3597),
    .Y(_00703_),
    .B1(_03790_));
 sg13g2_mux2_1 _10363_ (.A0(_00158_),
    .A1(net4351),
    .S(net3941),
    .X(_03791_));
 sg13g2_a21oi_1 _10364_ (.A1(net4057),
    .A2(_03791_),
    .Y(_03792_),
    .B1(_01512_));
 sg13g2_nor2_1 _10365_ (.A(net4236),
    .B(_03791_),
    .Y(_03793_));
 sg13g2_nor4_1 _10366_ (.A(_01516_),
    .B(net3596),
    .C(_03792_),
    .D(_03793_),
    .Y(_03794_));
 sg13g2_a21oi_1 _10367_ (.A1(_00922_),
    .A2(net3595),
    .Y(_00704_),
    .B1(_03794_));
 sg13g2_nor2_1 _10368_ (.A(_00162_),
    .B(net3940),
    .Y(_03795_));
 sg13g2_a21oi_1 _10369_ (.A1(net4156),
    .A2(net3940),
    .Y(_03796_),
    .B1(_03795_));
 sg13g2_a21oi_1 _10370_ (.A1(net4056),
    .A2(_03796_),
    .Y(_03797_),
    .B1(_01552_));
 sg13g2_nor2_1 _10371_ (.A(net4235),
    .B(_03796_),
    .Y(_03798_));
 sg13g2_nor4_1 _10372_ (.A(_01556_),
    .B(net3595),
    .C(_03797_),
    .D(_03798_),
    .Y(_03799_));
 sg13g2_a21oi_1 _10373_ (.A1(_00929_),
    .A2(net3595),
    .Y(_00705_),
    .B1(_03799_));
 sg13g2_mux2_1 _10374_ (.A0(_00166_),
    .A1(net4345),
    .S(net3940),
    .X(_03800_));
 sg13g2_a21oi_1 _10375_ (.A1(net4054),
    .A2(_03800_),
    .Y(_03801_),
    .B1(net4260));
 sg13g2_nand2_1 _10376_ (.Y(_03802_),
    .A(_01596_),
    .B(_03801_));
 sg13g2_nor2_1 _10377_ (.A(net4234),
    .B(_03800_),
    .Y(_03803_));
 sg13g2_nor3_1 _10378_ (.A(_01601_),
    .B(net3595),
    .C(_03803_),
    .Y(_03804_));
 sg13g2_a22oi_1 _10379_ (.Y(_00706_),
    .B1(_03802_),
    .B2(_03804_),
    .A2(net3595),
    .A1(_00936_));
 sg13g2_nor2_1 _10380_ (.A(_00170_),
    .B(net3940),
    .Y(_03805_));
 sg13g2_a21oi_1 _10381_ (.A1(net4155),
    .A2(net3941),
    .Y(_03806_),
    .B1(_03805_));
 sg13g2_inv_1 _10382_ (.Y(_03807_),
    .A(_03806_));
 sg13g2_a21oi_1 _10383_ (.A1(net4056),
    .A2(_03806_),
    .Y(_03808_),
    .B1(net4262));
 sg13g2_a221oi_1 _10384_ (.B2(_01649_),
    .C1(net3595),
    .B1(_03808_),
    .A1(net4299),
    .Y(_03809_),
    .A2(_03807_));
 sg13g2_a22oi_1 _10385_ (.Y(_00707_),
    .B1(_03809_),
    .B2(_01654_),
    .A2(net3595),
    .A1(_00943_));
 sg13g2_mux2_1 _10386_ (.A0(_00174_),
    .A1(net4338),
    .S(net3941),
    .X(_03810_));
 sg13g2_a21oi_1 _10387_ (.A1(net4052),
    .A2(_03810_),
    .Y(_03811_),
    .B1(net4259));
 sg13g2_nand2_1 _10388_ (.Y(_03812_),
    .A(_01707_),
    .B(_03811_));
 sg13g2_nor2_1 _10389_ (.A(net4231),
    .B(_03810_),
    .Y(_03813_));
 sg13g2_nor3_1 _10390_ (.A(_01713_),
    .B(net3596),
    .C(_03813_),
    .Y(_03814_));
 sg13g2_a22oi_1 _10391_ (.Y(_00708_),
    .B1(_03812_),
    .B2(_03814_),
    .A2(net3596),
    .A1(_00951_));
 sg13g2_mux2_1 _10392_ (.A0(_00178_),
    .A1(net4297),
    .S(net3938),
    .X(_03815_));
 sg13g2_a21oi_1 _10393_ (.A1(net4044),
    .A2(_03815_),
    .Y(_03816_),
    .B1(net4251));
 sg13g2_nand2_1 _10394_ (.Y(_03817_),
    .A(_01756_),
    .B(_03816_));
 sg13g2_nor2_1 _10395_ (.A(net4225),
    .B(_03815_),
    .Y(_03818_));
 sg13g2_nor3_1 _10396_ (.A(_01761_),
    .B(net3594),
    .C(_03818_),
    .Y(_03819_));
 sg13g2_a22oi_1 _10397_ (.Y(_00709_),
    .B1(_03817_),
    .B2(_03819_),
    .A2(net3594),
    .A1(_00958_));
 sg13g2_nor2_1 _10398_ (.A(_00182_),
    .B(net3939),
    .Y(_03820_));
 sg13g2_a21oi_1 _10399_ (.A1(net4154),
    .A2(net3939),
    .Y(_03821_),
    .B1(_03820_));
 sg13g2_a21oi_1 _10400_ (.A1(net4048),
    .A2(_03821_),
    .Y(_03822_),
    .B1(net4255));
 sg13g2_nand2_1 _10401_ (.Y(_03823_),
    .A(_01780_),
    .B(_03822_));
 sg13g2_nor2_1 _10402_ (.A(net4228),
    .B(_03821_),
    .Y(_03824_));
 sg13g2_nor3_1 _10403_ (.A(_01786_),
    .B(net3594),
    .C(_03824_),
    .Y(_03825_));
 sg13g2_a22oi_1 _10404_ (.Y(_00710_),
    .B1(_03823_),
    .B2(_03825_),
    .A2(net3594),
    .A1(_00966_));
 sg13g2_nor2_1 _10405_ (.A(_00186_),
    .B(net3938),
    .Y(_03826_));
 sg13g2_a21oi_1 _10406_ (.A1(net4153),
    .A2(net3938),
    .Y(_03827_),
    .B1(_03826_));
 sg13g2_a21oi_1 _10407_ (.A1(net4040),
    .A2(_03827_),
    .Y(_03828_),
    .B1(net4246));
 sg13g2_nand2_1 _10408_ (.Y(_03829_),
    .A(_01803_),
    .B(_03828_));
 sg13g2_nor2_1 _10409_ (.A(net4221),
    .B(_03827_),
    .Y(_03830_));
 sg13g2_nor3_1 _10410_ (.A(_01809_),
    .B(net3593),
    .C(_03830_),
    .Y(_03831_));
 sg13g2_a22oi_1 _10411_ (.Y(_00711_),
    .B1(_03829_),
    .B2(_03831_),
    .A2(net3593),
    .A1(_00974_));
 sg13g2_mux2_1 _10412_ (.A0(_00190_),
    .A1(net4284),
    .S(net3939),
    .X(_03832_));
 sg13g2_a21oi_1 _10413_ (.A1(net4046),
    .A2(_03832_),
    .Y(_03833_),
    .B1(net4252));
 sg13g2_nand2_1 _10414_ (.Y(_03834_),
    .A(_01826_),
    .B(_03833_));
 sg13g2_nor2_1 _10415_ (.A(net4229),
    .B(_03832_),
    .Y(_03835_));
 sg13g2_nor3_1 _10416_ (.A(_01831_),
    .B(_03783_),
    .C(_03835_),
    .Y(_03836_));
 sg13g2_a22oi_1 _10417_ (.Y(_00712_),
    .B1(_03834_),
    .B2(_03836_),
    .A2(net3594),
    .A1(_00982_));
 sg13g2_mux2_1 _10418_ (.A0(_00194_),
    .A1(net4280),
    .S(net3939),
    .X(_03837_));
 sg13g2_a21oi_1 _10419_ (.A1(net4046),
    .A2(_03837_),
    .Y(_03838_),
    .B1(net4255));
 sg13g2_nand2_1 _10420_ (.Y(_03839_),
    .A(_01852_),
    .B(_03838_));
 sg13g2_nor2_1 _10421_ (.A(net4229),
    .B(_03837_),
    .Y(_03840_));
 sg13g2_nor3_1 _10422_ (.A(_01857_),
    .B(net3594),
    .C(_03840_),
    .Y(_03841_));
 sg13g2_a22oi_1 _10423_ (.Y(_00713_),
    .B1(_03839_),
    .B2(_03841_),
    .A2(net3594),
    .A1(_00990_));
 sg13g2_nor2_1 _10424_ (.A(_00198_),
    .B(net3938),
    .Y(_03842_));
 sg13g2_a21oi_1 _10425_ (.A1(net4152),
    .A2(net3938),
    .Y(_03843_),
    .B1(_03842_));
 sg13g2_a21oi_1 _10426_ (.A1(net4041),
    .A2(_03843_),
    .Y(_03844_),
    .B1(net4247));
 sg13g2_nand2_1 _10427_ (.Y(_03845_),
    .A(_01871_),
    .B(_03844_));
 sg13g2_nor2_1 _10428_ (.A(net4222),
    .B(_03843_),
    .Y(_03846_));
 sg13g2_nor3_1 _10429_ (.A(_01877_),
    .B(net3593),
    .C(_03846_),
    .Y(_03847_));
 sg13g2_a22oi_1 _10430_ (.Y(_00714_),
    .B1(_03845_),
    .B2(_03847_),
    .A2(net3593),
    .A1(_01112_));
 sg13g2_nor2_1 _10431_ (.A(_00203_),
    .B(net3938),
    .Y(_03848_));
 sg13g2_a21oi_1 _10432_ (.A1(net4151),
    .A2(net3938),
    .Y(_03849_),
    .B1(_03848_));
 sg13g2_a21oi_1 _10433_ (.A1(net4040),
    .A2(_03849_),
    .Y(_03850_),
    .B1(net4246));
 sg13g2_nand2_1 _10434_ (.Y(_03851_),
    .A(_01892_),
    .B(_03850_));
 sg13g2_nor2_1 _10435_ (.A(net4221),
    .B(_03849_),
    .Y(_03852_));
 sg13g2_nor3_1 _10436_ (.A(_01898_),
    .B(net3593),
    .C(_03852_),
    .Y(_03853_));
 sg13g2_a22oi_1 _10437_ (.Y(_00715_),
    .B1(_03851_),
    .B2(_03853_),
    .A2(net3593),
    .A1(_01127_));
 sg13g2_mux2_1 _10438_ (.A0(_00207_),
    .A1(net4268),
    .S(net3938),
    .X(_03854_));
 sg13g2_a21oi_1 _10439_ (.A1(net4041),
    .A2(_03854_),
    .Y(_03855_),
    .B1(net4248));
 sg13g2_nand2_1 _10440_ (.Y(_03856_),
    .A(_01912_),
    .B(_03855_));
 sg13g2_nor2_1 _10441_ (.A(net4222),
    .B(_03854_),
    .Y(_03857_));
 sg13g2_nor3_1 _10442_ (.A(_01917_),
    .B(net3593),
    .C(_03857_),
    .Y(_03858_));
 sg13g2_a22oi_1 _10443_ (.Y(_00716_),
    .B1(_03856_),
    .B2(_03858_),
    .A2(net3593),
    .A1(_01140_));
 sg13g2_o21ai_1 _10444_ (.B1(_02253_),
    .Y(_03859_),
    .A1(_00022_),
    .A2(_01250_));
 sg13g2_nand2_1 _10445_ (.Y(_03860_),
    .A(net4316),
    .B(net4070));
 sg13g2_o21ai_1 _10446_ (.B1(net4307),
    .Y(_03861_),
    .A1(_01256_),
    .A2(_01263_));
 sg13g2_and4_2 _10447_ (.A(_01370_),
    .B(_03859_),
    .C(_03860_),
    .D(_03861_),
    .X(_03862_));
 sg13g2_nand4_1 _10448_ (.B(_03859_),
    .C(_03860_),
    .A(_01370_),
    .Y(_03863_),
    .D(_03861_));
 sg13g2_nor2b_1 _10449_ (.A(\cpu.keccak_alu.registers[64] ),
    .B_N(net4572),
    .Y(_03864_));
 sg13g2_nor2_2 _10450_ (.A(net4532),
    .B(net4530),
    .Y(_03865_));
 sg13g2_nand2_1 _10451_ (.Y(_03866_),
    .A(net4184),
    .B(net4179));
 sg13g2_nor2_1 _10452_ (.A(net4570),
    .B(net4546),
    .Y(_03867_));
 sg13g2_nor4_2 _10453_ (.A(net4561),
    .B(net4538),
    .C(net4531),
    .Y(_03868_),
    .D(net4525));
 sg13g2_nor2_1 _10454_ (.A(net4523),
    .B(net4519),
    .Y(_03869_));
 sg13g2_nand2_1 _10455_ (.Y(_03870_),
    .A(net4165),
    .B(net4162));
 sg13g2_nor2_1 _10456_ (.A(net4518),
    .B(net4514),
    .Y(_03871_));
 sg13g2_nand2_2 _10457_ (.Y(_03872_),
    .A(net4162),
    .B(net4158));
 sg13g2_nand3_1 _10458_ (.B(net4157),
    .C(_03868_),
    .A(net4164),
    .Y(_03873_));
 sg13g2_nand2_1 _10459_ (.Y(_03874_),
    .A(net3931),
    .B(_03873_));
 sg13g2_a22oi_1 _10460_ (.Y(_03875_),
    .B1(net3931),
    .B2(_03873_),
    .A2(net4091),
    .A1(_03868_));
 sg13g2_xnor2_1 _10461_ (.Y(_03876_),
    .A(net4521),
    .B(_03868_));
 sg13g2_xnor2_1 _10462_ (.Y(_03877_),
    .A(net4165),
    .B(_03868_));
 sg13g2_nand2_1 _10463_ (.Y(_03878_),
    .A(_00069_),
    .B(net4093));
 sg13g2_nand2_2 _10464_ (.Y(_03879_),
    .A(net4528),
    .B(_03878_));
 sg13g2_nand3_1 _10465_ (.B(_00069_),
    .C(net4093),
    .A(net4174),
    .Y(_03880_));
 sg13g2_and2_1 _10466_ (.A(_03879_),
    .B(_03880_),
    .X(_03881_));
 sg13g2_nand2_1 _10467_ (.Y(_03882_),
    .A(_03879_),
    .B(_03880_));
 sg13g2_xor2_1 _10468_ (.B(net4094),
    .A(_00069_),
    .X(_03883_));
 sg13g2_xnor2_1 _10469_ (.Y(_03884_),
    .A(_00069_),
    .B(net4094));
 sg13g2_and2_1 _10470_ (.A(net4570),
    .B(net4546),
    .X(_03885_));
 sg13g2_nand2_1 _10471_ (.Y(_03886_),
    .A(net4570),
    .B(net4546));
 sg13g2_nor2_2 _10472_ (.A(net4093),
    .B(_03885_),
    .Y(_03887_));
 sg13g2_nand2b_1 _10473_ (.Y(_03888_),
    .B(_03886_),
    .A_N(net4093));
 sg13g2_nor2_1 _10474_ (.A(net4487),
    .B(net4486),
    .Y(_03889_));
 sg13g2_nor3_1 _10475_ (.A(net4487),
    .B(net4486),
    .C(net4485),
    .Y(_03890_));
 sg13g2_nor4_2 _10476_ (.A(net4487),
    .B(net4486),
    .C(net4485),
    .Y(_03891_),
    .D(\cpu.keccak_alu.registers[183] ));
 sg13g2_nor2_1 _10477_ (.A(\cpu.keccak_alu.registers[172] ),
    .B(\cpu.keccak_alu.registers[173] ),
    .Y(_03892_));
 sg13g2_nor2_1 _10478_ (.A(\cpu.keccak_alu.registers[168] ),
    .B(\cpu.keccak_alu.registers[169] ),
    .Y(_03893_));
 sg13g2_nor2_1 _10479_ (.A(\cpu.keccak_alu.registers[170] ),
    .B(net4491),
    .Y(_03894_));
 sg13g2_nor4_2 _10480_ (.A(\cpu.keccak_alu.registers[168] ),
    .B(\cpu.keccak_alu.registers[169] ),
    .C(net4492),
    .Y(_03895_),
    .D(net4491));
 sg13g2_a21oi_2 _10481_ (.B1(net4157),
    .Y(_03896_),
    .A2(net4091),
    .A1(_03868_));
 sg13g2_a21o_2 _10482_ (.A2(net4091),
    .A1(_03868_),
    .B1(net4157),
    .X(_03897_));
 sg13g2_nor2_1 _10483_ (.A(net4512),
    .B(_03896_),
    .Y(_03898_));
 sg13g2_nor3_1 _10484_ (.A(net4510),
    .B(\cpu.keccak_alu.registers[137] ),
    .C(\cpu.keccak_alu.registers[139] ),
    .Y(_03899_));
 sg13g2_nor4_2 _10485_ (.A(net4510),
    .B(\cpu.keccak_alu.registers[137] ),
    .C(\cpu.keccak_alu.registers[138] ),
    .Y(_03900_),
    .D(\cpu.keccak_alu.registers[139] ));
 sg13g2_nor2_1 _10486_ (.A(net4508),
    .B(\cpu.keccak_alu.registers[141] ),
    .Y(_03901_));
 sg13g2_and2_1 _10487_ (.A(_03900_),
    .B(_03901_),
    .X(_03902_));
 sg13g2_nand3_1 _10488_ (.B(_03897_),
    .C(_03902_),
    .A(_01055_),
    .Y(_03903_));
 sg13g2_nor2_2 _10489_ (.A(\cpu.keccak_alu.registers[146] ),
    .B(\cpu.keccak_alu.registers[147] ),
    .Y(_03904_));
 sg13g2_nor2_1 _10490_ (.A(\cpu.keccak_alu.registers[148] ),
    .B(\cpu.keccak_alu.registers[149] ),
    .Y(_03905_));
 sg13g2_nor4_2 _10491_ (.A(\cpu.keccak_alu.registers[148] ),
    .B(\cpu.keccak_alu.registers[149] ),
    .C(\cpu.keccak_alu.registers[150] ),
    .Y(_03906_),
    .D(net4502));
 sg13g2_nor2_2 _10492_ (.A(\cpu.keccak_alu.registers[142] ),
    .B(net4504),
    .Y(_03907_));
 sg13g2_nor2_1 _10493_ (.A(net4503),
    .B(\cpu.keccak_alu.registers[145] ),
    .Y(_03908_));
 sg13g2_nor4_2 _10494_ (.A(net4503),
    .B(\cpu.keccak_alu.registers[145] ),
    .C(net4505),
    .Y(_03909_),
    .D(net4504));
 sg13g2_and4_2 _10495_ (.A(_01055_),
    .B(_03897_),
    .C(_03902_),
    .D(_03907_),
    .X(_03910_));
 sg13g2_nand4_1 _10496_ (.B(_03897_),
    .C(_03902_),
    .A(_01055_),
    .Y(_03911_),
    .D(_03907_));
 sg13g2_and4_2 _10497_ (.A(_01055_),
    .B(_03897_),
    .C(_03902_),
    .D(_03909_),
    .X(_03912_));
 sg13g2_and3_2 _10498_ (.X(_03913_),
    .A(_03904_),
    .B(_03906_),
    .C(_03908_));
 sg13g2_nand3_1 _10499_ (.B(_03906_),
    .C(_03908_),
    .A(_03904_),
    .Y(_03914_));
 sg13g2_nor2_2 _10500_ (.A(_03911_),
    .B(_03914_),
    .Y(_03915_));
 sg13g2_nor4_2 _10501_ (.A(net4501),
    .B(\cpu.keccak_alu.registers[153] ),
    .C(\cpu.keccak_alu.registers[154] ),
    .Y(_03916_),
    .D(net4499));
 sg13g2_inv_1 _10502_ (.Y(_03917_),
    .A(_03916_));
 sg13g2_or2_1 _10503_ (.X(_03918_),
    .B(\cpu.keccak_alu.registers[157] ),
    .A(\cpu.keccak_alu.registers[156] ));
 sg13g2_nor4_2 _10504_ (.A(\cpu.keccak_alu.registers[156] ),
    .B(\cpu.keccak_alu.registers[157] ),
    .C(\cpu.keccak_alu.registers[158] ),
    .Y(_03919_),
    .D(\cpu.keccak_alu.registers[159] ));
 sg13g2_nor2_1 _10505_ (.A(net4497),
    .B(net4496),
    .Y(_03920_));
 sg13g2_nor3_1 _10506_ (.A(net4497),
    .B(net4496),
    .C(\cpu.keccak_alu.registers[166] ),
    .Y(_03921_));
 sg13g2_nor2_1 _10507_ (.A(net4494),
    .B(net4493),
    .Y(_03922_));
 sg13g2_nor4_1 _10508_ (.A(\cpu.keccak_alu.registers[162] ),
    .B(net4495),
    .C(net4494),
    .D(net4493),
    .Y(_03923_));
 sg13g2_nand4_1 _10509_ (.B(_03919_),
    .C(_03921_),
    .A(_03916_),
    .Y(_03924_),
    .D(_03923_));
 sg13g2_nor2_2 _10510_ (.A(\cpu.keccak_alu.registers[167] ),
    .B(_03924_),
    .Y(_03925_));
 sg13g2_nor3_2 _10511_ (.A(_03911_),
    .B(_03914_),
    .C(_03917_),
    .Y(_03926_));
 sg13g2_nand3_1 _10512_ (.B(_03913_),
    .C(_03916_),
    .A(_03910_),
    .Y(_03927_));
 sg13g2_nor4_2 _10513_ (.A(_03911_),
    .B(_03914_),
    .C(_03917_),
    .Y(_03928_),
    .D(_03918_));
 sg13g2_and3_1 _10514_ (.X(_03929_),
    .A(_03913_),
    .B(_03916_),
    .C(_03919_));
 sg13g2_and2_1 _10515_ (.A(_03910_),
    .B(_03929_),
    .X(_03930_));
 sg13g2_nand2_2 _10516_ (.Y(_03931_),
    .A(_03910_),
    .B(_03929_));
 sg13g2_nor4_2 _10517_ (.A(net4497),
    .B(net4496),
    .C(\cpu.keccak_alu.registers[162] ),
    .Y(_03932_),
    .D(net4495));
 sg13g2_nor4_1 _10518_ (.A(net4494),
    .B(net4493),
    .C(\cpu.keccak_alu.registers[166] ),
    .D(\cpu.keccak_alu.registers[167] ),
    .Y(_03933_));
 sg13g2_nand3_1 _10519_ (.B(_03913_),
    .C(_03925_),
    .A(_03910_),
    .Y(_03934_));
 sg13g2_nand4_1 _10520_ (.B(_03910_),
    .C(_03913_),
    .A(_03893_),
    .Y(_03935_),
    .D(_03925_));
 sg13g2_nor3_2 _10521_ (.A(net4492),
    .B(net4491),
    .C(_03935_),
    .Y(_03936_));
 sg13g2_nand3_1 _10522_ (.B(_03915_),
    .C(_03925_),
    .A(_03895_),
    .Y(_03937_));
 sg13g2_nand4_1 _10523_ (.B(_03895_),
    .C(_03932_),
    .A(_03892_),
    .Y(_03938_),
    .D(_03933_));
 sg13g2_nor3_1 _10524_ (.A(\cpu.keccak_alu.registers[174] ),
    .B(\cpu.keccak_alu.registers[175] ),
    .C(_03938_),
    .Y(_03939_));
 sg13g2_inv_1 _10525_ (.Y(_03940_),
    .A(net3835));
 sg13g2_nor4_2 _10526_ (.A(\cpu.keccak_alu.registers[176] ),
    .B(\cpu.keccak_alu.registers[177] ),
    .C(\cpu.keccak_alu.registers[178] ),
    .Y(_03941_),
    .D(\cpu.keccak_alu.registers[179] ));
 sg13g2_and3_1 _10527_ (.X(_03942_),
    .A(net3780),
    .B(_03939_),
    .C(_03941_));
 sg13g2_nand3_1 _10528_ (.B(net3835),
    .C(_03941_),
    .A(net3780),
    .Y(_03943_));
 sg13g2_and2_1 _10529_ (.A(_03891_),
    .B(_03941_),
    .X(_03944_));
 sg13g2_nor2_2 _10530_ (.A(\cpu.keccak_alu.registers[186] ),
    .B(\cpu.keccak_alu.registers[187] ),
    .Y(_03945_));
 sg13g2_nor2_1 _10531_ (.A(\cpu.keccak_alu.registers[184] ),
    .B(\cpu.keccak_alu.registers[185] ),
    .Y(_03946_));
 sg13g2_nor4_2 _10532_ (.A(\cpu.keccak_alu.registers[184] ),
    .B(\cpu.keccak_alu.registers[185] ),
    .C(\cpu.keccak_alu.registers[186] ),
    .Y(_03947_),
    .D(net4484));
 sg13g2_nand4_1 _10533_ (.B(net3835),
    .C(_03944_),
    .A(net3780),
    .Y(_03948_),
    .D(_03946_));
 sg13g2_nand4_1 _10534_ (.B(net3835),
    .C(_03944_),
    .A(net3780),
    .Y(_03949_),
    .D(_03947_));
 sg13g2_nand2b_1 _10535_ (.Y(_03950_),
    .B(_03949_),
    .A_N(net4483));
 sg13g2_nand4_1 _10536_ (.B(_03930_),
    .C(net3835),
    .A(_03889_),
    .Y(_03951_),
    .D(_03941_));
 sg13g2_nand4_1 _10537_ (.B(_03930_),
    .C(net3835),
    .A(_03890_),
    .Y(_03952_),
    .D(_03941_));
 sg13g2_xor2_1 _10538_ (.B(_03951_),
    .A(net4485),
    .X(_03953_));
 sg13g2_xnor2_1 _10539_ (.Y(_03954_),
    .A(net4485),
    .B(_03951_));
 sg13g2_a22oi_1 _10540_ (.Y(_03955_),
    .B1(_03952_),
    .B2(\cpu.keccak_alu.registers[183] ),
    .A2(_03942_),
    .A1(_03891_));
 sg13g2_inv_1 _10541_ (.Y(_03956_),
    .A(_03955_));
 sg13g2_nand4_1 _10542_ (.B(\cpu.keccak_alu.registers[185] ),
    .C(\cpu.keccak_alu.registers[186] ),
    .A(\cpu.keccak_alu.registers[184] ),
    .Y(_03957_),
    .D(net4484));
 sg13g2_a21o_1 _10543_ (.A2(_03942_),
    .A1(_03891_),
    .B1(_03957_),
    .X(_03958_));
 sg13g2_nand2_1 _10544_ (.Y(_03959_),
    .A(_03949_),
    .B(_03958_));
 sg13g2_nand4_1 _10545_ (.B(_03954_),
    .C(_03956_),
    .A(_03950_),
    .Y(_03960_),
    .D(_03959_));
 sg13g2_nor4_2 _10546_ (.A(\cpu.keccak_alu.registers[176] ),
    .B(\cpu.keccak_alu.registers[177] ),
    .C(_03931_),
    .Y(_03961_),
    .D(_03940_));
 sg13g2_nand2_1 _10547_ (.Y(_03962_),
    .A(\cpu.keccak_alu.registers[178] ),
    .B(\cpu.keccak_alu.registers[179] ));
 sg13g2_or2_1 _10548_ (.X(_03963_),
    .B(_03962_),
    .A(_03961_));
 sg13g2_o21ai_1 _10549_ (.B1(_03943_),
    .Y(_03964_),
    .A1(_03961_),
    .A2(_03962_));
 sg13g2_nand4_1 _10550_ (.B(_03930_),
    .C(net3835),
    .A(net4487),
    .Y(_03965_),
    .D(_03941_));
 sg13g2_xnor2_1 _10551_ (.Y(_03966_),
    .A(_01029_),
    .B(_03942_));
 sg13g2_and2_1 _10552_ (.A(\cpu.keccak_alu.registers[174] ),
    .B(\cpu.keccak_alu.registers[175] ),
    .X(_03967_));
 sg13g2_o21ai_1 _10553_ (.B1(_03967_),
    .Y(_03968_),
    .A1(_03931_),
    .A2(_03938_));
 sg13g2_o21ai_1 _10554_ (.B1(_03968_),
    .Y(_03969_),
    .A1(_03931_),
    .A2(_03940_));
 sg13g2_nand3_1 _10555_ (.B(_03920_),
    .C(_03929_),
    .A(_03910_),
    .Y(_03970_));
 sg13g2_nand3b_1 _10556_ (.B(net3780),
    .C(_03932_),
    .Y(_03971_),
    .A_N(net4494));
 sg13g2_nand4_1 _10557_ (.B(net4495),
    .C(net4494),
    .A(\cpu.keccak_alu.registers[162] ),
    .Y(_03972_),
    .D(_03970_));
 sg13g2_and2_1 _10558_ (.A(_03971_),
    .B(_03972_),
    .X(_03973_));
 sg13g2_nand2_2 _10559_ (.Y(_03974_),
    .A(_03904_),
    .B(_03912_));
 sg13g2_and3_1 _10560_ (.X(_03975_),
    .A(\cpu.keccak_alu.registers[148] ),
    .B(\cpu.keccak_alu.registers[149] ),
    .C(net4502));
 sg13g2_a21oi_1 _10561_ (.A1(_03904_),
    .A2(_03912_),
    .Y(_03976_),
    .B1(_03975_));
 sg13g2_and2_1 _10562_ (.A(\cpu.keccak_alu.registers[168] ),
    .B(\cpu.keccak_alu.registers[169] ),
    .X(_03977_));
 sg13g2_mux2_1 _10563_ (.A0(_03893_),
    .A1(_03977_),
    .S(_03934_),
    .X(_03978_));
 sg13g2_inv_1 _10564_ (.Y(_03979_),
    .A(_03978_));
 sg13g2_nand2b_1 _10565_ (.Y(_03980_),
    .B(\cpu.keccak_alu.registers[150] ),
    .A_N(net4502));
 sg13g2_a21oi_1 _10566_ (.A1(_03905_),
    .A2(_03980_),
    .Y(_03981_),
    .B1(_03974_));
 sg13g2_nor4_1 _10567_ (.A(_03973_),
    .B(_03976_),
    .C(_03979_),
    .D(_03981_),
    .Y(_03982_));
 sg13g2_nand4_1 _10568_ (.B(_03966_),
    .C(_03969_),
    .A(_03964_),
    .Y(_03983_),
    .D(_03982_));
 sg13g2_nor2_2 _10569_ (.A(\cpu.keccak_alu.registers[190] ),
    .B(\cpu.keccak_alu.registers[191] ),
    .Y(_03984_));
 sg13g2_inv_1 _10570_ (.Y(_03985_),
    .A(_03984_));
 sg13g2_a21oi_1 _10571_ (.A1(_01106_),
    .A2(_03985_),
    .Y(_03986_),
    .B1(\cpu.keccak_alu.registers[188] ));
 sg13g2_nor2_1 _10572_ (.A(_03949_),
    .B(_03986_),
    .Y(_03987_));
 sg13g2_nand2_1 _10573_ (.Y(_03988_),
    .A(\cpu.keccak_alu.registers[158] ),
    .B(\cpu.keccak_alu.registers[159] ));
 sg13g2_nor2_1 _10574_ (.A(_03928_),
    .B(_03988_),
    .Y(_03989_));
 sg13g2_o21ai_1 _10575_ (.B1(_03931_),
    .Y(_03990_),
    .A1(_03928_),
    .A2(_03988_));
 sg13g2_inv_1 _10576_ (.Y(_03991_),
    .A(_03990_));
 sg13g2_and2_1 _10577_ (.A(net4492),
    .B(net4491),
    .X(_03992_));
 sg13g2_mux2_2 _10578_ (.A0(_03894_),
    .A1(_03992_),
    .S(_03935_),
    .X(_03993_));
 sg13g2_a21o_1 _10579_ (.A2(_03974_),
    .A1(\cpu.keccak_alu.registers[150] ),
    .B1(_03915_),
    .X(_03994_));
 sg13g2_nand3_1 _10580_ (.B(_03993_),
    .C(_03994_),
    .A(_03990_),
    .Y(_03995_));
 sg13g2_nand2_1 _10581_ (.Y(_03996_),
    .A(net4489),
    .B(_03936_));
 sg13g2_xnor2_1 _10582_ (.Y(_03997_),
    .A(net4489),
    .B(_03936_));
 sg13g2_nand2_1 _10583_ (.Y(_03998_),
    .A(net4497),
    .B(net4496));
 sg13g2_o21ai_1 _10584_ (.B1(_03970_),
    .Y(_03999_),
    .A1(net3780),
    .A2(_03998_));
 sg13g2_or4_1 _10585_ (.A(net4501),
    .B(net4500),
    .C(_03911_),
    .D(_03914_),
    .X(_04000_));
 sg13g2_and2_1 _10586_ (.A(\cpu.keccak_alu.registers[154] ),
    .B(\cpu.keccak_alu.registers[155] ),
    .X(_04001_));
 sg13g2_a21oi_1 _10587_ (.A1(_04000_),
    .A2(_04001_),
    .Y(_04002_),
    .B1(_03926_));
 sg13g2_a21o_1 _10588_ (.A2(_04001_),
    .A1(_04000_),
    .B1(_03926_),
    .X(_04003_));
 sg13g2_nand2_1 _10589_ (.Y(_04004_),
    .A(_03999_),
    .B(_04003_));
 sg13g2_nand3_1 _10590_ (.B(net4504),
    .C(_03903_),
    .A(net4505),
    .Y(_04005_));
 sg13g2_a21o_1 _10591_ (.A2(_03916_),
    .A1(\cpu.keccak_alu.registers[156] ),
    .B1(net4501),
    .X(_04006_));
 sg13g2_a21oi_1 _10592_ (.A1(_03910_),
    .A2(_03913_),
    .Y(_04007_),
    .B1(\cpu.keccak_alu.registers[152] ));
 sg13g2_a221oi_1 _10593_ (.B2(_03915_),
    .C1(_04007_),
    .B1(_04006_),
    .A1(_03911_),
    .Y(_04008_),
    .A2(_04005_));
 sg13g2_nand2b_1 _10594_ (.Y(_04009_),
    .B(net4507),
    .A_N(\cpu.keccak_alu.registers[138] ));
 sg13g2_nand4_1 _10595_ (.B(_03898_),
    .C(_03899_),
    .A(_00065_),
    .Y(_04010_),
    .D(_04009_));
 sg13g2_nor2b_1 _10596_ (.A(_00065_),
    .B_N(\cpu.keccak_alu.registers[139] ),
    .Y(_04011_));
 sg13g2_nand2_1 _10597_ (.Y(_04012_),
    .A(net4512),
    .B(\cpu.keccak_alu.registers[137] ));
 sg13g2_nand3_1 _10598_ (.B(net4509),
    .C(_04011_),
    .A(net4512),
    .Y(_04013_));
 sg13g2_o21ai_1 _10599_ (.B1(net4511),
    .Y(_04014_),
    .A1(_03897_),
    .A2(_04013_));
 sg13g2_or2_1 _10600_ (.X(_04015_),
    .B(_03902_),
    .A(net4508));
 sg13g2_xor2_1 _10601_ (.B(net4482),
    .A(net4484),
    .X(_04016_));
 sg13g2_or2_1 _10602_ (.X(_04017_),
    .B(net4482),
    .A(net4483));
 sg13g2_nand2_2 _10603_ (.Y(_04018_),
    .A(\cpu.keccak_alu.registers[190] ),
    .B(\cpu.keccak_alu.registers[191] ));
 sg13g2_a221oi_1 _10604_ (.B2(_04018_),
    .C1(_04016_),
    .B1(_04017_),
    .A1(net4503),
    .Y(_04019_),
    .A2(_03907_));
 sg13g2_nand2b_1 _10605_ (.Y(_04020_),
    .B(net4500),
    .A_N(net4502));
 sg13g2_nand2b_1 _10606_ (.Y(_04021_),
    .B(net4498),
    .A_N(net4499));
 sg13g2_nand2b_1 _10607_ (.Y(_04022_),
    .B(net4502),
    .A_N(net4500));
 sg13g2_nand2b_1 _10608_ (.Y(_04023_),
    .B(net4495),
    .A_N(net4493));
 sg13g2_nand4_1 _10609_ (.B(_04021_),
    .C(_04022_),
    .A(_04020_),
    .Y(_04024_),
    .D(_04023_));
 sg13g2_xnor2_1 _10610_ (.Y(_04025_),
    .A(\cpu.keccak_alu.registers[179] ),
    .B(net4486));
 sg13g2_nand2b_1 _10611_ (.Y(_04026_),
    .B(net4499),
    .A_N(net4498));
 sg13g2_nand2b_1 _10612_ (.Y(_04027_),
    .B(net4508),
    .A_N(net4506));
 sg13g2_nand3_1 _10613_ (.B(_04026_),
    .C(_04027_),
    .A(_04025_),
    .Y(_04028_));
 sg13g2_a21oi_1 _10614_ (.A1(net4503),
    .A2(\cpu.keccak_alu.registers[145] ),
    .Y(_04029_),
    .B1(_03909_));
 sg13g2_nand2b_1 _10615_ (.Y(_04030_),
    .B(net4490),
    .A_N(\cpu.keccak_alu.registers[173] ));
 sg13g2_nand2b_1 _10616_ (.Y(_04031_),
    .B(net4493),
    .A_N(net4495));
 sg13g2_nand2b_1 _10617_ (.Y(_04032_),
    .B(net4488),
    .A_N(net4490));
 sg13g2_nand3_1 _10618_ (.B(_04031_),
    .C(_04032_),
    .A(_04030_),
    .Y(_04033_));
 sg13g2_nor4_1 _10619_ (.A(_04024_),
    .B(_04028_),
    .C(_04029_),
    .D(_04033_),
    .Y(_04034_));
 sg13g2_nand4_1 _10620_ (.B(_04015_),
    .C(_04019_),
    .A(_04014_),
    .Y(_04035_),
    .D(_04034_));
 sg13g2_a221oi_1 _10621_ (.B2(_01064_),
    .C1(_04035_),
    .B1(_04010_),
    .A1(_01097_),
    .Y(_04036_),
    .A2(_03927_));
 sg13g2_nand3b_1 _10622_ (.B(\cpu.keccak_alu.registers[147] ),
    .C(\cpu.keccak_alu.registers[146] ),
    .Y(_04037_),
    .A_N(_03912_));
 sg13g2_nand2_1 _10623_ (.Y(_04038_),
    .A(_03974_),
    .B(_04037_));
 sg13g2_nor3_2 _10624_ (.A(_03911_),
    .B(_03914_),
    .C(_03924_),
    .Y(_04039_));
 sg13g2_o21ai_1 _10625_ (.B1(_03934_),
    .Y(_04040_),
    .A1(_01056_),
    .A2(_04039_));
 sg13g2_nand4_1 _10626_ (.B(_04036_),
    .C(_04038_),
    .A(_04008_),
    .Y(_04041_),
    .D(_04040_));
 sg13g2_or4_1 _10627_ (.A(_03995_),
    .B(_03997_),
    .C(_04004_),
    .D(_04041_),
    .X(_04042_));
 sg13g2_nand3_1 _10628_ (.B(net3780),
    .C(_03932_),
    .A(_03922_),
    .Y(_04043_));
 sg13g2_a21oi_2 _10629_ (.B1(_04039_),
    .Y(_04044_),
    .A2(_04043_),
    .A1(\cpu.keccak_alu.registers[166] ));
 sg13g2_nand2_1 _10630_ (.Y(_04045_),
    .A(\cpu.keccak_alu.registers[176] ),
    .B(\cpu.keccak_alu.registers[177] ));
 sg13g2_a21oi_1 _10631_ (.A1(net3780),
    .A2(net3835),
    .Y(_04046_),
    .B1(_04045_));
 sg13g2_nor2_1 _10632_ (.A(_03961_),
    .B(_04046_),
    .Y(_04047_));
 sg13g2_or2_1 _10633_ (.X(_04048_),
    .B(_04046_),
    .A(_03961_));
 sg13g2_or4_2 _10634_ (.A(_03987_),
    .B(_04042_),
    .C(_04044_),
    .D(_04047_),
    .X(_04049_));
 sg13g2_nor2b_2 _10635_ (.A(net4551),
    .B_N(_00108_),
    .Y(_04050_));
 sg13g2_and2_1 _10636_ (.A(net4550),
    .B(_00109_),
    .X(_04051_));
 sg13g2_nor2_1 _10637_ (.A(_04050_),
    .B(_04051_),
    .Y(_04052_));
 sg13g2_nor2b_2 _10638_ (.A(net4551),
    .B_N(_00106_),
    .Y(_04053_));
 sg13g2_and2_1 _10639_ (.A(net4551),
    .B(_00107_),
    .X(_04054_));
 sg13g2_nor2_1 _10640_ (.A(_04053_),
    .B(_04054_),
    .Y(_04055_));
 sg13g2_nor2_1 _10641_ (.A(_03949_),
    .B(_04017_),
    .Y(_04056_));
 sg13g2_nand2_1 _10642_ (.Y(_04057_),
    .A(_03984_),
    .B(_04056_));
 sg13g2_o21ai_1 _10643_ (.B1(_04057_),
    .Y(_04058_),
    .A1(_04018_),
    .A2(_04056_));
 sg13g2_mux2_2 _10644_ (.A0(_04018_),
    .A1(_03985_),
    .S(_04056_),
    .X(_04059_));
 sg13g2_xnor2_1 _10645_ (.Y(_04060_),
    .A(net4483),
    .B(_03949_));
 sg13g2_nand2b_1 _10646_ (.Y(_04061_),
    .B(_03961_),
    .A_N(\cpu.keccak_alu.registers[178] ));
 sg13g2_a22oi_1 _10647_ (.Y(_04062_),
    .B1(_03963_),
    .B2(_04061_),
    .A2(_03958_),
    .A1(_03948_));
 sg13g2_or2_1 _10648_ (.X(_04063_),
    .B(_04061_),
    .A(_01021_));
 sg13g2_and4_2 _10649_ (.A(_03956_),
    .B(_04060_),
    .C(_04062_),
    .D(_04063_),
    .X(_04064_));
 sg13g2_nand4_1 _10650_ (.B(_04060_),
    .C(_04062_),
    .A(_03956_),
    .Y(_04065_),
    .D(_04063_));
 sg13g2_o21ai_1 _10651_ (.B1(net4504),
    .Y(_04066_),
    .A1(net4505),
    .A2(_03903_));
 sg13g2_a22oi_1 _10652_ (.Y(_04067_),
    .B1(_04066_),
    .B2(_03911_),
    .A2(_04037_),
    .A1(_03974_));
 sg13g2_or4_1 _10653_ (.A(net4512),
    .B(net4511),
    .C(net4509),
    .D(_03896_),
    .X(_04068_));
 sg13g2_and4_1 _10654_ (.A(_01055_),
    .B(_00065_),
    .C(_03897_),
    .D(_03899_),
    .X(_04069_));
 sg13g2_a21oi_1 _10655_ (.A1(_04011_),
    .A2(_04068_),
    .Y(_04070_),
    .B1(_04069_));
 sg13g2_xor2_1 _10656_ (.B(_03903_),
    .A(net4505),
    .X(_04071_));
 sg13g2_o21ai_1 _10657_ (.B1(net4510),
    .Y(_04072_),
    .A1(_03897_),
    .A2(_04012_));
 sg13g2_xnor2_1 _10658_ (.Y(_04073_),
    .A(net4495),
    .B(net4493));
 sg13g2_xnor2_1 _10659_ (.Y(_04074_),
    .A(net4499),
    .B(net4498));
 sg13g2_xnor2_1 _10660_ (.Y(_04075_),
    .A(net4508),
    .B(net4506));
 sg13g2_nand3_1 _10661_ (.B(_04074_),
    .C(_04075_),
    .A(_04073_),
    .Y(_04076_));
 sg13g2_a21oi_1 _10662_ (.A1(net4503),
    .A2(_03907_),
    .Y(_04077_),
    .B1(_04076_));
 sg13g2_a21oi_1 _10663_ (.A1(net4508),
    .A2(_03900_),
    .Y(_04078_),
    .B1(net4509));
 sg13g2_a21oi_1 _10664_ (.A1(_03898_),
    .A2(_04078_),
    .Y(_04079_),
    .B1(net4510));
 sg13g2_nand3b_1 _10665_ (.B(_04020_),
    .C(_04022_),
    .Y(_04080_),
    .A_N(_04016_));
 sg13g2_xnor2_1 _10666_ (.Y(_04081_),
    .A(net4490),
    .B(net4488));
 sg13g2_nand2_1 _10667_ (.Y(_04082_),
    .A(_04025_),
    .B(_04081_));
 sg13g2_nor2_1 _10668_ (.A(net4507),
    .B(_03900_),
    .Y(_04083_));
 sg13g2_nor4_1 _10669_ (.A(_04029_),
    .B(_04080_),
    .C(_04082_),
    .D(_04083_),
    .Y(_04084_));
 sg13g2_nand3_1 _10670_ (.B(_04077_),
    .C(_04084_),
    .A(_04072_),
    .Y(_04085_));
 sg13g2_nor4_1 _10671_ (.A(_04070_),
    .B(_04071_),
    .C(_04079_),
    .D(_04085_),
    .Y(_04086_));
 sg13g2_xnor2_1 _10672_ (.Y(_04087_),
    .A(\cpu.keccak_alu.registers[156] ),
    .B(_03926_));
 sg13g2_xnor2_1 _10673_ (.Y(_04088_),
    .A(net4501),
    .B(_03915_));
 sg13g2_xor2_1 _10674_ (.B(_03915_),
    .A(net4501),
    .X(_04089_));
 sg13g2_and3_1 _10675_ (.X(_04090_),
    .A(_03904_),
    .B(_03905_),
    .C(_03912_));
 sg13g2_nand3_1 _10676_ (.B(_03905_),
    .C(_03912_),
    .A(_03904_),
    .Y(_04091_));
 sg13g2_a22oi_1 _10677_ (.Y(_04092_),
    .B1(_03980_),
    .B2(_04090_),
    .A2(_03975_),
    .A1(_03974_));
 sg13g2_nor3_1 _10678_ (.A(_04087_),
    .B(_04088_),
    .C(_04092_),
    .Y(_04093_));
 sg13g2_and4_1 _10679_ (.A(_03969_),
    .B(_04067_),
    .C(_04086_),
    .D(_04093_),
    .X(_04094_));
 sg13g2_a21oi_1 _10680_ (.A1(\cpu.keccak_alu.registers[150] ),
    .A2(_04091_),
    .Y(_04095_),
    .B1(_03915_));
 sg13g2_a21oi_1 _10681_ (.A1(_01098_),
    .A2(_03937_),
    .Y(_04096_),
    .B1(_04095_));
 sg13g2_and4_1 _10682_ (.A(_03996_),
    .B(_03999_),
    .C(_04040_),
    .D(_04096_),
    .X(_04097_));
 sg13g2_nand3_1 _10683_ (.B(\cpu.keccak_alu.registers[159] ),
    .C(_03928_),
    .A(_01121_),
    .Y(_04098_));
 sg13g2_o21ai_1 _10684_ (.B1(_04098_),
    .Y(_04099_),
    .A1(_03945_),
    .A2(_03948_));
 sg13g2_a21oi_1 _10685_ (.A1(_01121_),
    .A2(_03928_),
    .Y(_04100_),
    .B1(_03989_));
 sg13g2_nor3_1 _10686_ (.A(_04044_),
    .B(_04099_),
    .C(_04100_),
    .Y(_04101_));
 sg13g2_a22oi_1 _10687_ (.Y(_04102_),
    .B1(_03971_),
    .B2(_03972_),
    .A2(_03943_),
    .A1(_01029_));
 sg13g2_and4_1 _10688_ (.A(_03965_),
    .B(_03978_),
    .C(_03993_),
    .D(_04003_),
    .X(_04103_));
 sg13g2_and4_1 _10689_ (.A(_03954_),
    .B(_04048_),
    .C(_04102_),
    .D(_04103_),
    .X(_04104_));
 sg13g2_and4_2 _10690_ (.A(_04094_),
    .B(_04097_),
    .C(_04101_),
    .D(_04104_),
    .X(_04105_));
 sg13g2_nand4_1 _10691_ (.B(_04097_),
    .C(_04101_),
    .A(_04094_),
    .Y(_04106_),
    .D(_04104_));
 sg13g2_and4_1 _10692_ (.A(_04052_),
    .B(net3588),
    .C(net3583),
    .D(net3574),
    .X(_04107_));
 sg13g2_nand4_1 _10693_ (.B(net3588),
    .C(net3583),
    .A(_04052_),
    .Y(_04108_),
    .D(net3574));
 sg13g2_and4_1 _10694_ (.A(_04055_),
    .B(net3588),
    .C(net3583),
    .D(net3574),
    .X(_04109_));
 sg13g2_nand4_1 _10695_ (.B(net3588),
    .C(net3583),
    .A(_04055_),
    .Y(_04110_),
    .D(net3574));
 sg13g2_mux2_1 _10696_ (.A0(_04108_),
    .A1(_04110_),
    .S(net3878),
    .X(_04111_));
 sg13g2_mux2_1 _10697_ (.A0(_04107_),
    .A1(_04109_),
    .S(net3877),
    .X(_04112_));
 sg13g2_nor2b_1 _10698_ (.A(net4552),
    .B_N(_00112_),
    .Y(_04113_));
 sg13g2_and2_1 _10699_ (.A(net4553),
    .B(_00113_),
    .X(_04114_));
 sg13g2_nor2_1 _10700_ (.A(_04113_),
    .B(_04114_),
    .Y(_04115_));
 sg13g2_nor2b_1 _10701_ (.A(net4550),
    .B_N(_00110_),
    .Y(_04116_));
 sg13g2_and2_1 _10702_ (.A(net4553),
    .B(_00111_),
    .X(_04117_));
 sg13g2_nor2_1 _10703_ (.A(_04116_),
    .B(_04117_),
    .Y(_04118_));
 sg13g2_nor2b_1 _10704_ (.A(_03955_),
    .B_N(_04060_),
    .Y(_04119_));
 sg13g2_nor3_1 _10705_ (.A(_03997_),
    .B(_04044_),
    .C(_04047_),
    .Y(_04120_));
 sg13g2_nor4_1 _10706_ (.A(_04070_),
    .B(_04071_),
    .C(_04079_),
    .D(_04085_),
    .Y(_04121_));
 sg13g2_nand4_1 _10707_ (.B(_04067_),
    .C(_04089_),
    .A(_03999_),
    .Y(_04122_),
    .D(_04121_));
 sg13g2_nor4_2 _10708_ (.A(_03973_),
    .B(_03979_),
    .C(_03991_),
    .Y(_04123_),
    .D(_04122_));
 sg13g2_and4_2 _10709_ (.A(_03959_),
    .B(_04119_),
    .C(_04120_),
    .D(_04123_),
    .X(_04124_));
 sg13g2_nand4_1 _10710_ (.B(_04119_),
    .C(_04120_),
    .A(_03959_),
    .Y(_04125_),
    .D(_04123_));
 sg13g2_nand2_1 _10711_ (.Y(_04126_),
    .A(_03966_),
    .B(_03993_));
 sg13g2_nor4_1 _10712_ (.A(_04002_),
    .B(_04087_),
    .C(_04092_),
    .D(_04095_),
    .Y(_04127_));
 sg13g2_nand4_1 _10713_ (.B(_03969_),
    .C(_04040_),
    .A(_03964_),
    .Y(_04128_),
    .D(_04127_));
 sg13g2_nor4_2 _10714_ (.A(_03953_),
    .B(net3636),
    .C(_04126_),
    .Y(_04129_),
    .D(_04128_));
 sg13g2_or4_1 _10715_ (.A(_03953_),
    .B(net3636),
    .C(_04126_),
    .D(_04128_),
    .X(_04130_));
 sg13g2_nor2_1 _10716_ (.A(net3563),
    .B(net3552),
    .Y(_04131_));
 sg13g2_nand2_1 _10717_ (.Y(_04132_),
    .A(net3568),
    .B(net3557));
 sg13g2_nor4_1 _10718_ (.A(_04116_),
    .B(_04117_),
    .C(net3559),
    .D(net3548),
    .Y(_04133_));
 sg13g2_and4_2 _10719_ (.A(_04058_),
    .B(_04064_),
    .C(_04105_),
    .D(_04115_),
    .X(_04134_));
 sg13g2_and4_1 _10720_ (.A(net3588),
    .B(net3583),
    .C(net3574),
    .D(_04118_),
    .X(_04135_));
 sg13g2_mux2_2 _10721_ (.A0(_04134_),
    .A1(_04135_),
    .S(net3878),
    .X(_04136_));
 sg13g2_nor2b_1 _10722_ (.A(net4556),
    .B_N(_00100_),
    .Y(_04137_));
 sg13g2_and2_1 _10723_ (.A(net4557),
    .B(_00101_),
    .X(_04138_));
 sg13g2_nor2b_2 _10724_ (.A(net4556),
    .B_N(_00098_),
    .Y(_04139_));
 sg13g2_and2_1 _10725_ (.A(net4556),
    .B(_00099_),
    .X(_04140_));
 sg13g2_nor4_2 _10726_ (.A(net3560),
    .B(net3549),
    .C(_04139_),
    .Y(_04141_),
    .D(_04140_));
 sg13g2_or4_1 _10727_ (.A(net3560),
    .B(net3549),
    .C(_04139_),
    .D(_04140_),
    .X(_04142_));
 sg13g2_nor4_1 _10728_ (.A(net3560),
    .B(net3549),
    .C(_04137_),
    .D(_04138_),
    .Y(_04143_));
 sg13g2_or4_1 _10729_ (.A(net3560),
    .B(net3549),
    .C(_04137_),
    .D(_04138_),
    .X(_04144_));
 sg13g2_mux2_2 _10730_ (.A0(_04141_),
    .A1(_04143_),
    .S(net3887),
    .X(_04145_));
 sg13g2_mux2_1 _10731_ (.A0(_04142_),
    .A1(_04144_),
    .S(net3887),
    .X(_04146_));
 sg13g2_nor2b_2 _10732_ (.A(net4557),
    .B_N(_00104_),
    .Y(_04147_));
 sg13g2_and2_1 _10733_ (.A(net4554),
    .B(_00105_),
    .X(_04148_));
 sg13g2_nor2_2 _10734_ (.A(_04147_),
    .B(_04148_),
    .Y(_04149_));
 sg13g2_nor2b_2 _10735_ (.A(net4563),
    .B_N(_00102_),
    .Y(_04150_));
 sg13g2_and2_1 _10736_ (.A(net4554),
    .B(_00103_),
    .X(_04151_));
 sg13g2_nor2_2 _10737_ (.A(_04150_),
    .B(_04151_),
    .Y(_04152_));
 sg13g2_and4_1 _10738_ (.A(net3590),
    .B(net3585),
    .C(net3576),
    .D(_04149_),
    .X(_04153_));
 sg13g2_nand4_1 _10739_ (.B(net3586),
    .C(net3577),
    .A(net3591),
    .Y(_04154_),
    .D(_04149_));
 sg13g2_and4_1 _10740_ (.A(net3590),
    .B(net3585),
    .C(net3576),
    .D(_04152_),
    .X(_04155_));
 sg13g2_nand4_1 _10741_ (.B(net3586),
    .C(net3577),
    .A(net3591),
    .Y(_04156_),
    .D(_04152_));
 sg13g2_mux2_1 _10742_ (.A0(_04154_),
    .A1(_04156_),
    .S(net3879),
    .X(_04157_));
 sg13g2_mux2_1 _10743_ (.A0(_04153_),
    .A1(_04155_),
    .S(net3879),
    .X(_04158_));
 sg13g2_mux4_1 _10744_ (.S0(net3906),
    .A0(_04112_),
    .A1(_04136_),
    .A2(_04145_),
    .A3(_04158_),
    .S1(net3781),
    .X(_04159_));
 sg13g2_nor2b_2 _10745_ (.A(net4548),
    .B_N(_00124_),
    .Y(_04160_));
 sg13g2_and2_1 _10746_ (.A(net4548),
    .B(_00125_),
    .X(_04161_));
 sg13g2_or2_1 _10747_ (.X(_04162_),
    .B(_04161_),
    .A(_04160_));
 sg13g2_nor2b_1 _10748_ (.A(net4550),
    .B_N(_00122_),
    .Y(_04163_));
 sg13g2_nand2_1 _10749_ (.Y(_04164_),
    .A(net4549),
    .B(_00123_));
 sg13g2_nand2b_1 _10750_ (.Y(_04165_),
    .B(_04164_),
    .A_N(_04163_));
 sg13g2_nor4_1 _10751_ (.A(_03960_),
    .B(_03983_),
    .C(_04049_),
    .D(_04165_),
    .Y(_04166_));
 sg13g2_nor4_2 _10752_ (.A(net3636),
    .B(net3582),
    .C(net3573),
    .Y(_04167_),
    .D(_04162_));
 sg13g2_or4_1 _10753_ (.A(net3636),
    .B(net3582),
    .C(net3573),
    .D(_04162_),
    .X(_04168_));
 sg13g2_nor4_1 _10754_ (.A(net3636),
    .B(net3582),
    .C(net3573),
    .D(_04165_),
    .Y(_04169_));
 sg13g2_or4_1 _10755_ (.A(net3636),
    .B(net3582),
    .C(net3573),
    .D(_04165_),
    .X(_04170_));
 sg13g2_mux2_1 _10756_ (.A0(_04167_),
    .A1(_04169_),
    .S(net3877),
    .X(_04171_));
 sg13g2_nor2b_1 _10757_ (.A(net4548),
    .B_N(_00126_),
    .Y(_04172_));
 sg13g2_and2_1 _10758_ (.A(net4549),
    .B(_00127_),
    .X(_04173_));
 sg13g2_nor2_1 _10759_ (.A(_04172_),
    .B(_04173_),
    .Y(_04174_));
 sg13g2_nor2b_1 _10760_ (.A(net4549),
    .B_N(_00128_),
    .Y(_04175_));
 sg13g2_and2_1 _10761_ (.A(net4549),
    .B(net4576),
    .X(_04176_));
 sg13g2_or2_1 _10762_ (.X(_04177_),
    .B(_04176_),
    .A(_04175_));
 sg13g2_nor4_1 _10763_ (.A(net3559),
    .B(net3548),
    .C(_04172_),
    .D(_04173_),
    .Y(_04178_));
 sg13g2_nor4_2 _10764_ (.A(net3559),
    .B(net3548),
    .C(_04175_),
    .Y(_04179_),
    .D(_04176_));
 sg13g2_nor4_2 _10765_ (.A(net3636),
    .B(net3582),
    .C(net3573),
    .Y(_04180_),
    .D(_04177_));
 sg13g2_and4_1 _10766_ (.A(net3588),
    .B(net3583),
    .C(net3574),
    .D(_04174_),
    .X(_04181_));
 sg13g2_nand4_1 _10767_ (.B(net3584),
    .C(net3575),
    .A(net3589),
    .Y(_04182_),
    .D(_04174_));
 sg13g2_mux2_2 _10768_ (.A0(_04180_),
    .A1(_04181_),
    .S(net3877),
    .X(_04183_));
 sg13g2_mux4_1 _10769_ (.S0(net3877),
    .A0(_04167_),
    .A1(_04169_),
    .A2(_04180_),
    .A3(_04181_),
    .S1(net3905),
    .X(_04184_));
 sg13g2_nor2_1 _10770_ (.A(net4552),
    .B(_01168_),
    .Y(_04185_));
 sg13g2_and2_1 _10771_ (.A(net4552),
    .B(_00117_),
    .X(_04186_));
 sg13g2_nor2_1 _10772_ (.A(_04185_),
    .B(_04186_),
    .Y(_04187_));
 sg13g2_nor2b_1 _10773_ (.A(net4554),
    .B_N(_00114_),
    .Y(_04188_));
 sg13g2_nand2_1 _10774_ (.Y(_04189_),
    .A(net4554),
    .B(_00115_));
 sg13g2_nand2b_2 _10775_ (.Y(_04190_),
    .B(_04189_),
    .A_N(_04188_));
 sg13g2_nor4_2 _10776_ (.A(_03960_),
    .B(_03983_),
    .C(_04049_),
    .Y(_04191_),
    .D(_04190_));
 sg13g2_nor4_1 _10777_ (.A(net3559),
    .B(net3548),
    .C(_04185_),
    .D(_04186_),
    .Y(_04192_));
 sg13g2_and4_1 _10778_ (.A(net3588),
    .B(net3583),
    .C(net3574),
    .D(_04187_),
    .X(_04193_));
 sg13g2_nor4_1 _10779_ (.A(net3636),
    .B(net3582),
    .C(net3573),
    .D(_04190_),
    .Y(_04194_));
 sg13g2_mux2_2 _10780_ (.A0(_04193_),
    .A1(_04194_),
    .S(net3878),
    .X(_04195_));
 sg13g2_nor2b_1 _10781_ (.A(net4553),
    .B_N(_00120_),
    .Y(_04196_));
 sg13g2_a21oi_2 _10782_ (.B1(_04196_),
    .Y(_04197_),
    .A2(_00121_),
    .A1(net4553));
 sg13g2_nor2b_2 _10783_ (.A(net4554),
    .B_N(_00118_),
    .Y(_04198_));
 sg13g2_and2_1 _10784_ (.A(net4552),
    .B(_00119_),
    .X(_04199_));
 sg13g2_nor2_1 _10785_ (.A(_04198_),
    .B(_04199_),
    .Y(_04200_));
 sg13g2_and4_1 _10786_ (.A(net3589),
    .B(net3584),
    .C(net3575),
    .D(_04197_),
    .X(_04201_));
 sg13g2_nand4_1 _10787_ (.B(net3584),
    .C(net3575),
    .A(net3589),
    .Y(_04202_),
    .D(_04197_));
 sg13g2_and4_1 _10788_ (.A(net3588),
    .B(net3583),
    .C(net3574),
    .D(_04200_),
    .X(_04203_));
 sg13g2_nand4_1 _10789_ (.B(net3584),
    .C(net3575),
    .A(net3589),
    .Y(_04204_),
    .D(_04200_));
 sg13g2_mux2_1 _10790_ (.A0(_04201_),
    .A1(_04203_),
    .S(net3877),
    .X(_04205_));
 sg13g2_mux4_1 _10791_ (.S0(net3905),
    .A0(_04171_),
    .A1(_04183_),
    .A2(_04195_),
    .A3(_04205_),
    .S1(net3781),
    .X(_04206_));
 sg13g2_mux2_1 _10792_ (.A0(_04159_),
    .A1(_04206_),
    .S(net3925),
    .X(_04207_));
 sg13g2_nand2_1 _10793_ (.Y(_04208_),
    .A(net3838),
    .B(_04207_));
 sg13g2_nor2b_1 _10794_ (.A(net4556),
    .B_N(_00092_),
    .Y(_04209_));
 sg13g2_and2_1 _10795_ (.A(net4557),
    .B(_00093_),
    .X(_04210_));
 sg13g2_nor2_1 _10796_ (.A(_04209_),
    .B(_04210_),
    .Y(_04211_));
 sg13g2_nor2b_1 _10797_ (.A(net4557),
    .B_N(_00090_),
    .Y(_04212_));
 sg13g2_and2_1 _10798_ (.A(net4556),
    .B(_00091_),
    .X(_04213_));
 sg13g2_nor2_1 _10799_ (.A(_04212_),
    .B(_04213_),
    .Y(_04214_));
 sg13g2_and4_1 _10800_ (.A(net3591),
    .B(net3586),
    .C(net3577),
    .D(_04211_),
    .X(_04215_));
 sg13g2_nand4_1 _10801_ (.B(net3586),
    .C(net3578),
    .A(net3592),
    .Y(_04216_),
    .D(_04211_));
 sg13g2_and4_1 _10802_ (.A(net3591),
    .B(net3586),
    .C(net3577),
    .D(_04214_),
    .X(_04217_));
 sg13g2_nand4_1 _10803_ (.B(net3587),
    .C(net3578),
    .A(net3591),
    .Y(_04218_),
    .D(_04214_));
 sg13g2_mux2_1 _10804_ (.A0(_04215_),
    .A1(_04217_),
    .S(net3881),
    .X(_04219_));
 sg13g2_mux2_1 _10805_ (.A0(_04216_),
    .A1(_04218_),
    .S(net3881),
    .X(_04220_));
 sg13g2_nor2b_2 _10806_ (.A(net4556),
    .B_N(_00096_),
    .Y(_04221_));
 sg13g2_and2_1 _10807_ (.A(net4556),
    .B(_00097_),
    .X(_04222_));
 sg13g2_nor2_1 _10808_ (.A(_04221_),
    .B(_04222_),
    .Y(_04223_));
 sg13g2_nor2b_2 _10809_ (.A(net4557),
    .B_N(_00094_),
    .Y(_04224_));
 sg13g2_and2_1 _10810_ (.A(net4557),
    .B(_00095_),
    .X(_04225_));
 sg13g2_nor2_1 _10811_ (.A(_04224_),
    .B(_04225_),
    .Y(_04226_));
 sg13g2_nand4_1 _10812_ (.B(net3587),
    .C(net3577),
    .A(net3592),
    .Y(_04227_),
    .D(_04223_));
 sg13g2_and4_1 _10813_ (.A(net3591),
    .B(net3586),
    .C(net3577),
    .D(_04226_),
    .X(_04228_));
 sg13g2_nand4_1 _10814_ (.B(net3587),
    .C(net3578),
    .A(net3592),
    .Y(_04229_),
    .D(_04226_));
 sg13g2_mux2_1 _10815_ (.A0(_04227_),
    .A1(_04229_),
    .S(net3881),
    .X(_04230_));
 sg13g2_nor2b_2 _10816_ (.A(net4559),
    .B_N(_00086_),
    .Y(_04231_));
 sg13g2_and2_1 _10817_ (.A(net4560),
    .B(_00087_),
    .X(_04232_));
 sg13g2_nor2_1 _10818_ (.A(_04231_),
    .B(_04232_),
    .Y(_04233_));
 sg13g2_nand4_1 _10819_ (.B(net3586),
    .C(net3577),
    .A(net3591),
    .Y(_04234_),
    .D(_04233_));
 sg13g2_nor2b_2 _10820_ (.A(net4560),
    .B_N(_00088_),
    .Y(_04235_));
 sg13g2_and2_1 _10821_ (.A(net4556),
    .B(_00089_),
    .X(_04236_));
 sg13g2_or2_1 _10822_ (.X(_04237_),
    .B(_04236_),
    .A(_04235_));
 sg13g2_nor4_1 _10823_ (.A(_03960_),
    .B(_03983_),
    .C(_04049_),
    .D(_04237_),
    .Y(_04238_));
 sg13g2_or4_1 _10824_ (.A(_04059_),
    .B(net3582),
    .C(net3573),
    .D(_04237_),
    .X(_04239_));
 sg13g2_nor2b_2 _10825_ (.A(net4568),
    .B_N(_00082_),
    .Y(_04240_));
 sg13g2_and2_2 _10826_ (.A(net4569),
    .B(_00083_),
    .X(_04241_));
 sg13g2_nor2b_2 _10827_ (.A(net4569),
    .B_N(_00084_),
    .Y(_04242_));
 sg13g2_and2_2 _10828_ (.A(net4571),
    .B(_00085_),
    .X(_04243_));
 sg13g2_nor2_1 _10829_ (.A(_04242_),
    .B(_04243_),
    .Y(_04244_));
 sg13g2_nand4_1 _10830_ (.B(net3586),
    .C(net3577),
    .A(net3591),
    .Y(_04245_),
    .D(_04244_));
 sg13g2_nor4_2 _10831_ (.A(net3560),
    .B(net3549),
    .C(_04242_),
    .Y(_04246_),
    .D(_04243_));
 sg13g2_nor4_2 _10832_ (.A(net3564),
    .B(net3553),
    .C(_04240_),
    .Y(_04247_),
    .D(_04241_));
 sg13g2_mux2_1 _10833_ (.A0(_04246_),
    .A1(_04247_),
    .S(net3880),
    .X(_04248_));
 sg13g2_nor4_1 _10834_ (.A(net3561),
    .B(net3550),
    .C(_04235_),
    .D(_04236_),
    .Y(_04249_));
 sg13g2_nor4_2 _10835_ (.A(net3561),
    .B(net3550),
    .C(_04231_),
    .Y(_04250_),
    .D(_04232_));
 sg13g2_mux2_1 _10836_ (.A0(_04249_),
    .A1(_04250_),
    .S(net3880),
    .X(_04251_));
 sg13g2_mux4_1 _10837_ (.S0(net3881),
    .A0(_04246_),
    .A1(_04247_),
    .A2(_04249_),
    .A3(_04250_),
    .S1(net3907),
    .X(_04252_));
 sg13g2_nor4_1 _10838_ (.A(net3560),
    .B(net3549),
    .C(_04224_),
    .D(_04225_),
    .Y(_04253_));
 sg13g2_nor4_2 _10839_ (.A(net3560),
    .B(net3549),
    .C(_04221_),
    .Y(_04254_),
    .D(_04222_));
 sg13g2_or4_1 _10840_ (.A(net3560),
    .B(net3549),
    .C(_04221_),
    .D(_04222_),
    .X(_04255_));
 sg13g2_mux2_2 _10841_ (.A0(_04253_),
    .A1(_04254_),
    .S(net3887),
    .X(_04256_));
 sg13g2_mux4_1 _10842_ (.S0(net3783),
    .A0(_04219_),
    .A1(_04248_),
    .A2(_04256_),
    .A3(_04251_),
    .S1(net3907),
    .X(_04257_));
 sg13g2_nor2_1 _10843_ (.A(_03874_),
    .B(_03896_),
    .Y(_04258_));
 sg13g2_nand3_1 _10844_ (.B(_03873_),
    .C(_03897_),
    .A(net3931),
    .Y(_04259_));
 sg13g2_nand2_1 _10845_ (.Y(_04260_),
    .A(net4559),
    .B(_00073_));
 sg13g2_o21ai_1 _10846_ (.B1(_04260_),
    .Y(_04261_),
    .A1(net4559),
    .A2(_01167_));
 sg13g2_nand2_1 _10847_ (.Y(_04262_),
    .A(net4565),
    .B(_00071_));
 sg13g2_nand2b_1 _10848_ (.Y(_04263_),
    .B(_00070_),
    .A_N(net4566));
 sg13g2_nand2_1 _10849_ (.Y(_04264_),
    .A(_04262_),
    .B(_04263_));
 sg13g2_mux2_1 _10850_ (.A0(_04261_),
    .A1(_04264_),
    .S(net3880),
    .X(_04265_));
 sg13g2_nand2_1 _10851_ (.Y(_04266_),
    .A(net4572),
    .B(_00068_));
 sg13g2_nor2_1 _10852_ (.A(net4570),
    .B(_01166_),
    .Y(_04267_));
 sg13g2_a21oi_2 _10853_ (.B1(_04267_),
    .Y(_04268_),
    .A2(_00068_),
    .A1(net4569));
 sg13g2_o21ai_1 _10854_ (.B1(net3904),
    .Y(_04269_),
    .A1(_00066_),
    .A2(_03886_));
 sg13g2_a221oi_1 _10855_ (.B2(_04268_),
    .C1(_04269_),
    .B1(net3893),
    .A1(\cpu.keccak_alu.registers[64] ),
    .Y(_04270_),
    .A2(net4093));
 sg13g2_a221oi_1 _10856_ (.B2(_04265_),
    .C1(_04270_),
    .B1(net3909),
    .A1(_03879_),
    .Y(_04271_),
    .A2(_03880_));
 sg13g2_a21oi_1 _10857_ (.A1(_04131_),
    .A2(_04271_),
    .Y(_04272_),
    .B1(net3925));
 sg13g2_nand2_1 _10858_ (.Y(_04273_),
    .A(net4559),
    .B(_00081_));
 sg13g2_nand2b_1 _10859_ (.Y(_04274_),
    .B(_00080_),
    .A_N(net4558));
 sg13g2_nand2_1 _10860_ (.Y(_04275_),
    .A(_04273_),
    .B(_04274_));
 sg13g2_nand2_1 _10861_ (.Y(_04276_),
    .A(net3888),
    .B(_04275_));
 sg13g2_nand2_1 _10862_ (.Y(_04277_),
    .A(net4558),
    .B(_00079_));
 sg13g2_nand2b_1 _10863_ (.Y(_04278_),
    .B(_00078_),
    .A_N(net4558));
 sg13g2_and2_1 _10864_ (.A(_04277_),
    .B(_04278_),
    .X(_04279_));
 sg13g2_o21ai_1 _10865_ (.B1(_04276_),
    .Y(_04280_),
    .A1(net3888),
    .A2(_04279_));
 sg13g2_nand2_1 _10866_ (.Y(_04281_),
    .A(net4558),
    .B(_00075_));
 sg13g2_nor2b_1 _10867_ (.A(net4560),
    .B_N(_00074_),
    .Y(_04282_));
 sg13g2_a21oi_1 _10868_ (.A1(net4558),
    .A2(_00075_),
    .Y(_04283_),
    .B1(_04282_));
 sg13g2_and2_1 _10869_ (.A(net3882),
    .B(_04283_),
    .X(_04284_));
 sg13g2_nand2_1 _10870_ (.Y(_04285_),
    .A(net4558),
    .B(_00077_));
 sg13g2_nand2b_1 _10871_ (.Y(_04286_),
    .B(_00076_),
    .A_N(net4559));
 sg13g2_and2_1 _10872_ (.A(_04285_),
    .B(_04286_),
    .X(_04287_));
 sg13g2_a21oi_1 _10873_ (.A1(net3887),
    .A2(_04287_),
    .Y(_04288_),
    .B1(_04284_));
 sg13g2_o21ai_1 _10874_ (.B1(net3900),
    .Y(_04289_),
    .A1(net3541),
    .A2(_04288_));
 sg13g2_nor2_1 _10875_ (.A(net3541),
    .B(_04280_),
    .Y(_04290_));
 sg13g2_o21ai_1 _10876_ (.B1(net3907),
    .Y(_04291_),
    .A1(net3541),
    .A2(_04280_));
 sg13g2_nand3_1 _10877_ (.B(_04289_),
    .C(_04291_),
    .A(net3790),
    .Y(_04292_));
 sg13g2_a21oi_1 _10878_ (.A1(_04272_),
    .A2(_04292_),
    .Y(_04293_),
    .B1(net3833));
 sg13g2_o21ai_1 _10879_ (.B1(_04293_),
    .Y(_04294_),
    .A1(net3916),
    .A2(_04257_));
 sg13g2_nand4_1 _10880_ (.B(_03900_),
    .C(_03906_),
    .A(_03891_),
    .Y(_04295_),
    .D(_03909_));
 sg13g2_nand3_1 _10881_ (.B(_03941_),
    .C(_03947_),
    .A(_03895_),
    .Y(_04296_));
 sg13g2_nor4_1 _10882_ (.A(net4483),
    .B(net4482),
    .C(\cpu.keccak_alu.registers[174] ),
    .D(\cpu.keccak_alu.registers[175] ),
    .Y(_04297_));
 sg13g2_nor4_1 _10883_ (.A(net4512),
    .B(\cpu.keccak_alu.registers[167] ),
    .C(net4489),
    .D(net4488),
    .Y(_04298_));
 sg13g2_nor4_1 _10884_ (.A(\cpu.keccak_alu.registers[146] ),
    .B(\cpu.keccak_alu.registers[147] ),
    .C(net4507),
    .D(net4506),
    .Y(_04299_));
 sg13g2_nand4_1 _10885_ (.B(_04297_),
    .C(_04298_),
    .A(_03984_),
    .Y(_04300_),
    .D(_04299_));
 sg13g2_nor4_2 _10886_ (.A(_03924_),
    .B(_04295_),
    .C(_04296_),
    .Y(_04301_),
    .D(_04300_));
 sg13g2_or4_1 _10887_ (.A(_03924_),
    .B(_04295_),
    .C(_04296_),
    .D(_04300_),
    .X(_04302_));
 sg13g2_and3_2 _10888_ (.X(_04303_),
    .A(\cpu.keccak_alu.registers[64] ),
    .B(net4094),
    .C(net3831));
 sg13g2_nand2_1 _10889_ (.Y(_04304_),
    .A(_03865_),
    .B(_04303_));
 sg13g2_nand4_1 _10890_ (.B(_03865_),
    .C(net4089),
    .A(net4167),
    .Y(_04305_),
    .D(_04303_));
 sg13g2_nor4_1 _10891_ (.A(net3559),
    .B(net3548),
    .C(_04198_),
    .D(_04199_),
    .Y(_04306_));
 sg13g2_nor4_1 _10892_ (.A(net3559),
    .B(net3548),
    .C(_04160_),
    .D(_04161_),
    .Y(_04307_));
 sg13g2_nor4_2 _10893_ (.A(net3562),
    .B(net3551),
    .C(_04150_),
    .Y(_04308_),
    .D(_04151_));
 sg13g2_nor4_2 _10894_ (.A(net3562),
    .B(net3551),
    .C(_04147_),
    .Y(_04309_),
    .D(_04148_));
 sg13g2_mux2_1 _10895_ (.A0(_04308_),
    .A1(_04309_),
    .S(net3889),
    .X(_04310_));
 sg13g2_nor4_1 _10896_ (.A(_04053_),
    .B(_04054_),
    .C(net3559),
    .D(net3548),
    .Y(_04311_));
 sg13g2_nor4_1 _10897_ (.A(_04050_),
    .B(_04051_),
    .C(net3559),
    .D(net3548),
    .Y(_04312_));
 sg13g2_mux2_1 _10898_ (.A0(_04311_),
    .A1(_04312_),
    .S(net3886),
    .X(_04313_));
 sg13g2_nand4_1 _10899_ (.B(_04208_),
    .C(_04294_),
    .A(net4018),
    .Y(_04314_),
    .D(_04305_));
 sg13g2_o21ai_1 _10900_ (.B1(_04314_),
    .Y(_04315_),
    .A1(net4019),
    .A2(_03864_));
 sg13g2_xor2_1 _10901_ (.B(_04315_),
    .A(\cpu.keccak_alu.registers[0] ),
    .X(_04316_));
 sg13g2_o21ai_1 _10902_ (.B1(net4210),
    .Y(_04317_),
    .A1(net4574),
    .A2(\cpu.keccak_alu.registers[192] ));
 sg13g2_a21oi_1 _10903_ (.A1(net4574),
    .A2(\cpu.keccak_alu.registers[192] ),
    .Y(_04318_),
    .B1(_04317_));
 sg13g2_xor2_1 _10904_ (.B(\cpu.keccak_alu.registers[64] ),
    .A(\cpu.keccak_alu.registers[0] ),
    .X(_04319_));
 sg13g2_o21ai_1 _10905_ (.B1(net4385),
    .Y(_04320_),
    .A1(_04318_),
    .A2(_04319_));
 sg13g2_a21o_1 _10906_ (.A2(_04319_),
    .A1(_04318_),
    .B1(_04320_),
    .X(_04321_));
 sg13g2_o21ai_1 _10907_ (.B1(_04321_),
    .Y(_04322_),
    .A1(net4385),
    .A2(_04316_));
 sg13g2_nor3_1 _10908_ (.A(net4070),
    .B(_01250_),
    .C(_01288_),
    .Y(_04323_));
 sg13g2_or3_2 _10909_ (.A(net4070),
    .B(_01250_),
    .C(_01288_),
    .X(_04324_));
 sg13g2_nor2b_2 _10910_ (.A(net3755),
    .B_N(net3754),
    .Y(_04325_));
 sg13g2_nand3_1 _10911_ (.B(_02279_),
    .C(net3754),
    .A(_02256_),
    .Y(_04326_));
 sg13g2_a22oi_1 _10912_ (.Y(_04327_),
    .B1(_04326_),
    .B2(net267),
    .A2(_02482_),
    .A1(_02459_));
 sg13g2_o21ai_1 _10913_ (.B1(net3739),
    .Y(_04328_),
    .A1(net3814),
    .A2(_04327_));
 sg13g2_a21oi_1 _10914_ (.A1(net4265),
    .A2(_04322_),
    .Y(_04329_),
    .B1(_04328_));
 sg13g2_a21oi_1 _10915_ (.A1(_00997_),
    .A2(net3733),
    .Y(_00717_),
    .B1(_04329_));
 sg13g2_nand2b_1 _10916_ (.Y(_04330_),
    .B(_00066_),
    .A_N(net4572));
 sg13g2_nand3b_1 _10917_ (.B(net3832),
    .C(_04330_),
    .Y(_04331_),
    .A_N(_03864_));
 sg13g2_nor2_1 _10918_ (.A(net4545),
    .B(_04331_),
    .Y(_04332_));
 sg13g2_nand2_1 _10919_ (.Y(_04333_),
    .A(_03865_),
    .B(_04332_));
 sg13g2_nor3_1 _10920_ (.A(net4523),
    .B(net3933),
    .C(_04333_),
    .Y(_04334_));
 sg13g2_nor2_1 _10921_ (.A(net4565),
    .B(_00101_),
    .Y(_04335_));
 sg13g2_nand2b_1 _10922_ (.Y(_04336_),
    .B(net4563),
    .A_N(_00102_));
 sg13g2_nor2b_2 _10923_ (.A(_04335_),
    .B_N(_04336_),
    .Y(_04337_));
 sg13g2_nor4_1 _10924_ (.A(net3638),
    .B(net3580),
    .C(net3571),
    .D(_04337_),
    .Y(_04338_));
 sg13g2_nor2_1 _10925_ (.A(net4565),
    .B(_00099_),
    .Y(_04339_));
 sg13g2_nand2b_1 _10926_ (.Y(_04340_),
    .B(net4565),
    .A_N(_00100_));
 sg13g2_nor2b_2 _10927_ (.A(_04339_),
    .B_N(_04340_),
    .Y(_04341_));
 sg13g2_nor4_1 _10928_ (.A(net3638),
    .B(net3580),
    .C(net3571),
    .D(_04341_),
    .Y(_04342_));
 sg13g2_mux2_1 _10929_ (.A0(_04338_),
    .A1(_04342_),
    .S(net3884),
    .X(_04343_));
 sg13g2_nor2_2 _10930_ (.A(net4554),
    .B(_00105_),
    .Y(_04344_));
 sg13g2_nand2b_1 _10931_ (.Y(_04345_),
    .B(net4551),
    .A_N(_00106_));
 sg13g2_nor2b_2 _10932_ (.A(_04344_),
    .B_N(_04345_),
    .Y(_04346_));
 sg13g2_nor4_2 _10933_ (.A(net3638),
    .B(net3580),
    .C(net3571),
    .Y(_04347_),
    .D(_04346_));
 sg13g2_nor2_1 _10934_ (.A(net4563),
    .B(_00103_),
    .Y(_04348_));
 sg13g2_nand2b_1 _10935_ (.Y(_04349_),
    .B(net4563),
    .A_N(_00104_));
 sg13g2_nor2b_2 _10936_ (.A(_04348_),
    .B_N(_04349_),
    .Y(_04350_));
 sg13g2_nor4_1 _10937_ (.A(net3638),
    .B(net3580),
    .C(net3571),
    .D(_04350_),
    .Y(_04351_));
 sg13g2_mux2_1 _10938_ (.A0(_04347_),
    .A1(_04351_),
    .S(net3885),
    .X(_04352_));
 sg13g2_mux2_1 _10939_ (.A0(_04343_),
    .A1(_04352_),
    .S(net3911),
    .X(_04353_));
 sg13g2_nor2_1 _10940_ (.A(net4550),
    .B(_00109_),
    .Y(_04354_));
 sg13g2_nor2b_1 _10941_ (.A(_00110_),
    .B_N(net4550),
    .Y(_04355_));
 sg13g2_nor2_2 _10942_ (.A(_04354_),
    .B(_04355_),
    .Y(_04356_));
 sg13g2_nor2_1 _10943_ (.A(net4551),
    .B(_00107_),
    .Y(_04357_));
 sg13g2_nor2b_1 _10944_ (.A(_00108_),
    .B_N(net4550),
    .Y(_04358_));
 sg13g2_nor2_2 _10945_ (.A(_04357_),
    .B(_04358_),
    .Y(_04359_));
 sg13g2_nor3_2 _10946_ (.A(net3564),
    .B(net3553),
    .C(_04359_),
    .Y(_04360_));
 sg13g2_nor3_2 _10947_ (.A(net3563),
    .B(net3552),
    .C(_04356_),
    .Y(_04361_));
 sg13g2_nor4_1 _10948_ (.A(net3638),
    .B(net3580),
    .C(net3571),
    .D(_04359_),
    .Y(_04362_));
 sg13g2_mux2_2 _10949_ (.A0(_04360_),
    .A1(_04361_),
    .S(net3892),
    .X(_04363_));
 sg13g2_nor2_2 _10950_ (.A(net4552),
    .B(_00113_),
    .Y(_04364_));
 sg13g2_nor2b_1 _10951_ (.A(_00114_),
    .B_N(net4567),
    .Y(_04365_));
 sg13g2_nor2_2 _10952_ (.A(_04364_),
    .B(_04365_),
    .Y(_04366_));
 sg13g2_nor4_2 _10953_ (.A(net3637),
    .B(net3579),
    .C(net3570),
    .Y(_04367_),
    .D(_04366_));
 sg13g2_nor2_1 _10954_ (.A(net4552),
    .B(_00111_),
    .Y(_04368_));
 sg13g2_nor2b_1 _10955_ (.A(_00112_),
    .B_N(net4552),
    .Y(_04369_));
 sg13g2_nor2_2 _10956_ (.A(_04368_),
    .B(_04369_),
    .Y(_04370_));
 sg13g2_nor4_1 _10957_ (.A(net3637),
    .B(net3579),
    .C(net3570),
    .D(_04370_),
    .Y(_04371_));
 sg13g2_mux2_2 _10958_ (.A0(_04367_),
    .A1(_04371_),
    .S(net3883),
    .X(_04372_));
 sg13g2_mux2_1 _10959_ (.A0(_04363_),
    .A1(_04372_),
    .S(net3911),
    .X(_04373_));
 sg13g2_mux4_1 _10960_ (.S0(net3911),
    .A0(_04343_),
    .A1(_04352_),
    .A2(_04363_),
    .A3(_04372_),
    .S1(net3792),
    .X(_04374_));
 sg13g2_mux2_2 _10961_ (.A0(_00125_),
    .A1(_00126_),
    .S(net4548),
    .X(_04375_));
 sg13g2_nor4_2 _10962_ (.A(_03960_),
    .B(_03983_),
    .C(_04049_),
    .Y(_04376_),
    .D(_04375_));
 sg13g2_or4_1 _10963_ (.A(net3639),
    .B(net3581),
    .C(net3572),
    .D(_04375_),
    .X(_04377_));
 sg13g2_nor2_2 _10964_ (.A(net4549),
    .B(_00123_),
    .Y(_04378_));
 sg13g2_nand2b_1 _10965_ (.Y(_04379_),
    .B(net4548),
    .A_N(_00124_));
 sg13g2_nor2b_2 _10966_ (.A(_04378_),
    .B_N(_04379_),
    .Y(_04380_));
 sg13g2_nor4_1 _10967_ (.A(net3639),
    .B(net3579),
    .C(net3570),
    .D(_04380_),
    .Y(_04381_));
 sg13g2_or4_1 _10968_ (.A(net3637),
    .B(net3581),
    .C(net3572),
    .D(_04380_),
    .X(_04382_));
 sg13g2_mux2_1 _10969_ (.A0(_04377_),
    .A1(_04382_),
    .S(net3885),
    .X(_04383_));
 sg13g2_mux2_1 _10970_ (.A0(_04376_),
    .A1(_04381_),
    .S(net3883),
    .X(_04384_));
 sg13g2_nor2b_1 _10971_ (.A(net4548),
    .B_N(_00127_),
    .Y(_04385_));
 sg13g2_a21o_2 _10972_ (.A2(_00128_),
    .A1(net4549),
    .B1(_04385_),
    .X(_04386_));
 sg13g2_nor4_2 _10973_ (.A(_03960_),
    .B(_03983_),
    .C(_04049_),
    .Y(_04387_),
    .D(_04386_));
 sg13g2_nor2_2 _10974_ (.A(net4564),
    .B(net4198),
    .Y(_04388_));
 sg13g2_nor4_2 _10975_ (.A(_00129_),
    .B(_03960_),
    .C(_03983_),
    .Y(_04389_),
    .D(_04049_));
 sg13g2_nor4_1 _10976_ (.A(net3637),
    .B(net3579),
    .C(net3572),
    .D(_04386_),
    .Y(_04390_));
 sg13g2_nor4_1 _10977_ (.A(net4576),
    .B(net3639),
    .C(net3581),
    .D(net3570),
    .Y(_04391_));
 sg13g2_a22oi_1 _10978_ (.Y(_04392_),
    .B1(_04391_),
    .B2(_04388_),
    .A2(_04390_),
    .A1(net3883));
 sg13g2_a221oi_1 _10979_ (.B2(_04388_),
    .C1(net3903),
    .B1(_04391_),
    .A1(net3883),
    .Y(_04393_),
    .A2(_04390_));
 sg13g2_a21oi_1 _10980_ (.A1(net3903),
    .A2(_04383_),
    .Y(_04394_),
    .B1(_04393_));
 sg13g2_nor2_1 _10981_ (.A(net4566),
    .B(_00117_),
    .Y(_04395_));
 sg13g2_nor2b_1 _10982_ (.A(_00118_),
    .B_N(net4566),
    .Y(_04396_));
 sg13g2_nor2_1 _10983_ (.A(_04395_),
    .B(_04396_),
    .Y(_04397_));
 sg13g2_nor2_1 _10984_ (.A(net4566),
    .B(_00115_),
    .Y(_04398_));
 sg13g2_a21oi_2 _10985_ (.B1(_04398_),
    .Y(_04399_),
    .A2(_01168_),
    .A1(net4566));
 sg13g2_nor3_2 _10986_ (.A(net3563),
    .B(net3552),
    .C(_04399_),
    .Y(_04400_));
 sg13g2_nor3_2 _10987_ (.A(net3563),
    .B(net3552),
    .C(_04397_),
    .Y(_04401_));
 sg13g2_nor4_1 _10988_ (.A(net3637),
    .B(net3579),
    .C(net3570),
    .D(_04399_),
    .Y(_04402_));
 sg13g2_mux2_1 _10989_ (.A0(_04400_),
    .A1(_04401_),
    .S(net3890),
    .X(_04403_));
 sg13g2_nor2_2 _10990_ (.A(net4552),
    .B(_00121_),
    .Y(_04404_));
 sg13g2_nor2b_1 _10991_ (.A(_00122_),
    .B_N(net4550),
    .Y(_04405_));
 sg13g2_nor2_2 _10992_ (.A(_04404_),
    .B(_04405_),
    .Y(_04406_));
 sg13g2_nor4_1 _10993_ (.A(net3637),
    .B(net3579),
    .C(net3570),
    .D(_04406_),
    .Y(_04407_));
 sg13g2_nor2_2 _10994_ (.A(net4554),
    .B(_00119_),
    .Y(_04408_));
 sg13g2_nor2b_1 _10995_ (.A(_00120_),
    .B_N(net4561),
    .Y(_04409_));
 sg13g2_nor2_1 _10996_ (.A(_04408_),
    .B(_04409_),
    .Y(_04410_));
 sg13g2_nor3_2 _10997_ (.A(net3563),
    .B(net3552),
    .C(_04410_),
    .Y(_04411_));
 sg13g2_nor3_2 _10998_ (.A(net3563),
    .B(net3552),
    .C(_04406_),
    .Y(_04412_));
 sg13g2_mux2_1 _10999_ (.A0(_04411_),
    .A1(_04412_),
    .S(net3891),
    .X(_04413_));
 sg13g2_mux2_1 _11000_ (.A0(_04403_),
    .A1(_04413_),
    .S(net3908),
    .X(_04414_));
 sg13g2_mux4_1 _11001_ (.S0(net3792),
    .A0(_04353_),
    .A1(_04373_),
    .A2(_04414_),
    .A3(_04394_),
    .S1(net3928),
    .X(_04415_));
 sg13g2_nor2_1 _11002_ (.A(net4564),
    .B(_00093_),
    .Y(_04416_));
 sg13g2_nand2b_1 _11003_ (.Y(_04417_),
    .B(net4564),
    .A_N(_00094_));
 sg13g2_nor2b_2 _11004_ (.A(_04416_),
    .B_N(_04417_),
    .Y(_04418_));
 sg13g2_nor4_1 _11005_ (.A(net3639),
    .B(net3580),
    .C(net3571),
    .D(_04418_),
    .Y(_04419_));
 sg13g2_nand2b_1 _11006_ (.Y(_04420_),
    .B(net4562),
    .A_N(_00092_));
 sg13g2_o21ai_1 _11007_ (.B1(_04420_),
    .Y(_04421_),
    .A1(net4564),
    .A2(_00091_));
 sg13g2_and3_1 _11008_ (.X(_04422_),
    .A(net3569),
    .B(net3558),
    .C(_04421_));
 sg13g2_nand3_1 _11009_ (.B(net3558),
    .C(_04421_),
    .A(net3569),
    .Y(_04423_));
 sg13g2_nor3_2 _11010_ (.A(net3566),
    .B(net3555),
    .C(_04418_),
    .Y(_04424_));
 sg13g2_nand3b_1 _11011_ (.B(net3558),
    .C(net3569),
    .Y(_04425_),
    .A_N(_04418_));
 sg13g2_mux2_1 _11012_ (.A0(_04422_),
    .A1(_04424_),
    .S(net3895),
    .X(_04426_));
 sg13g2_nor2_1 _11013_ (.A(net4564),
    .B(_00097_),
    .Y(_04427_));
 sg13g2_nand2b_1 _11014_ (.Y(_04428_),
    .B(net4564),
    .A_N(_00098_));
 sg13g2_nor2b_1 _11015_ (.A(_04427_),
    .B_N(_04428_),
    .Y(_04429_));
 sg13g2_nor2_1 _11016_ (.A(net4565),
    .B(_00095_),
    .Y(_04430_));
 sg13g2_nand2b_1 _11017_ (.Y(_04431_),
    .B(net4564),
    .A_N(_00096_));
 sg13g2_nor2b_2 _11018_ (.A(_04430_),
    .B_N(_04431_),
    .Y(_04432_));
 sg13g2_nor4_1 _11019_ (.A(net3638),
    .B(net3580),
    .C(net3571),
    .D(_04432_),
    .Y(_04433_));
 sg13g2_or2_1 _11020_ (.X(_04434_),
    .B(_00085_),
    .A(net4569));
 sg13g2_nand2b_2 _11021_ (.Y(_04435_),
    .B(net4562),
    .A_N(_00086_));
 sg13g2_nand2_1 _11022_ (.Y(_04436_),
    .A(_04434_),
    .B(_04435_));
 sg13g2_nor2_1 _11023_ (.A(net4569),
    .B(_00083_),
    .Y(_04437_));
 sg13g2_nand2b_1 _11024_ (.Y(_04438_),
    .B(net4569),
    .A_N(_00084_));
 sg13g2_nor2b_2 _11025_ (.A(_04437_),
    .B_N(_04438_),
    .Y(_04439_));
 sg13g2_nor3_1 _11026_ (.A(net3565),
    .B(net3554),
    .C(_04439_),
    .Y(_04440_));
 sg13g2_nand3b_1 _11027_ (.B(net3556),
    .C(net3567),
    .Y(_04441_),
    .A_N(_04439_));
 sg13g2_and3_1 _11028_ (.X(_04442_),
    .A(net3567),
    .B(net3556),
    .C(_04436_));
 sg13g2_nand3_1 _11029_ (.B(net3556),
    .C(_04436_),
    .A(net3567),
    .Y(_04443_));
 sg13g2_nor4_1 _11030_ (.A(net3638),
    .B(net3581),
    .C(net3572),
    .D(_04439_),
    .Y(_04444_));
 sg13g2_or2_1 _11031_ (.X(_04445_),
    .B(_00089_),
    .A(net4562));
 sg13g2_nand2b_1 _11032_ (.Y(_04446_),
    .B(net4562),
    .A_N(_00090_));
 sg13g2_nand2_2 _11033_ (.Y(_04447_),
    .A(_04445_),
    .B(_04446_));
 sg13g2_nand2b_1 _11034_ (.Y(_04448_),
    .B(net4559),
    .A_N(_00088_));
 sg13g2_o21ai_1 _11035_ (.B1(_04448_),
    .Y(_04449_),
    .A1(net4562),
    .A2(_00087_));
 sg13g2_and3_1 _11036_ (.X(_04450_),
    .A(net3567),
    .B(net3556),
    .C(_04449_));
 sg13g2_nand3_1 _11037_ (.B(net3556),
    .C(_04449_),
    .A(net3567),
    .Y(_04451_));
 sg13g2_and3_2 _11038_ (.X(_04452_),
    .A(net3567),
    .B(net3556),
    .C(_04447_));
 sg13g2_nand3_1 _11039_ (.B(net3556),
    .C(_04447_),
    .A(net3567),
    .Y(_04453_));
 sg13g2_mux2_1 _11040_ (.A0(_04450_),
    .A1(_04452_),
    .S(net3895),
    .X(_04454_));
 sg13g2_mux4_1 _11041_ (.S0(net3894),
    .A0(_04441_),
    .A1(_04443_),
    .A2(_04451_),
    .A3(_04453_),
    .S1(net3910),
    .X(_04455_));
 sg13g2_nor3_1 _11042_ (.A(net3566),
    .B(net3555),
    .C(_04432_),
    .Y(_04456_));
 sg13g2_nand3b_1 _11043_ (.B(net3558),
    .C(net3569),
    .Y(_04457_),
    .A_N(_04432_));
 sg13g2_nor3_1 _11044_ (.A(net3565),
    .B(net3554),
    .C(_04429_),
    .Y(_04458_));
 sg13g2_nand3b_1 _11045_ (.B(net3558),
    .C(net3569),
    .Y(_04459_),
    .A_N(_04429_));
 sg13g2_mux2_1 _11046_ (.A0(_04456_),
    .A1(_04458_),
    .S(net3895),
    .X(_04460_));
 sg13g2_mux4_1 _11047_ (.S0(net3894),
    .A0(_04423_),
    .A1(_04425_),
    .A2(_04457_),
    .A3(_04459_),
    .S1(net3910),
    .X(_04461_));
 sg13g2_mux2_1 _11048_ (.A0(_04455_),
    .A1(_04461_),
    .S(net3792),
    .X(_04462_));
 sg13g2_mux2_1 _11049_ (.A0(_00077_),
    .A1(_00078_),
    .S(net4568),
    .X(_04463_));
 sg13g2_nand2b_1 _11050_ (.Y(_04464_),
    .B(net4568),
    .A_N(_00076_));
 sg13g2_or2_1 _11051_ (.X(_04465_),
    .B(_00075_),
    .A(net4568));
 sg13g2_nand2_1 _11052_ (.Y(_04466_),
    .A(_04464_),
    .B(_04465_));
 sg13g2_nor4_2 _11053_ (.A(net3639),
    .B(net3580),
    .C(net3572),
    .Y(_04467_),
    .D(_04463_));
 sg13g2_nand2b_1 _11054_ (.Y(_04468_),
    .B(net4571),
    .A_N(_00082_));
 sg13g2_mux2_1 _11055_ (.A0(_00081_),
    .A1(_00082_),
    .S(net4568),
    .X(_04469_));
 sg13g2_nor4_2 _11056_ (.A(net3638),
    .B(net3581),
    .C(net3571),
    .Y(_04470_),
    .D(_04469_));
 sg13g2_nand2b_2 _11057_ (.Y(_04471_),
    .B(net4558),
    .A_N(_00080_));
 sg13g2_o21ai_1 _11058_ (.B1(_04471_),
    .Y(_04472_),
    .A1(net4558),
    .A2(_00079_));
 sg13g2_nor3_1 _11059_ (.A(net3565),
    .B(net3554),
    .C(_04469_),
    .Y(_04473_));
 sg13g2_and4_2 _11060_ (.A(net3592),
    .B(net3587),
    .C(net3578),
    .D(_04472_),
    .X(_04474_));
 sg13g2_and3_1 _11061_ (.X(_04475_),
    .A(net3568),
    .B(net3556),
    .C(_04466_));
 sg13g2_nor3_1 _11062_ (.A(net3565),
    .B(net3554),
    .C(_04463_),
    .Y(_04476_));
 sg13g2_mux2_1 _11063_ (.A0(_04475_),
    .A1(_04476_),
    .S(net3893),
    .X(_04477_));
 sg13g2_mux4_1 _11064_ (.S0(net3884),
    .A0(_04470_),
    .A1(_04474_),
    .A2(_04476_),
    .A3(_04475_),
    .S1(net3902),
    .X(_04478_));
 sg13g2_a21oi_1 _11065_ (.A1(net3794),
    .A2(_04478_),
    .Y(_04479_),
    .B1(net3929));
 sg13g2_o21ai_1 _11066_ (.B1(net4093),
    .Y(_04480_),
    .A1(_00066_),
    .A2(net3542));
 sg13g2_nand2b_1 _11067_ (.Y(_04481_),
    .B(net4572),
    .A_N(_00070_));
 sg13g2_nor2_1 _11068_ (.A(net4572),
    .B(_00068_),
    .Y(_04482_));
 sg13g2_o21ai_1 _11069_ (.B1(_04481_),
    .Y(_04483_),
    .A1(net4569),
    .A2(_00068_));
 sg13g2_nand3_1 _11070_ (.B(net3557),
    .C(_04483_),
    .A(net3568),
    .Y(_04484_));
 sg13g2_nand3_1 _11071_ (.B(net3568),
    .C(net3557),
    .A(_01166_),
    .Y(_04485_));
 sg13g2_a22oi_1 _11072_ (.Y(_04486_),
    .B1(_04485_),
    .B2(_03885_),
    .A2(_04484_),
    .A1(net3893));
 sg13g2_a21oi_1 _11073_ (.A1(_04480_),
    .A2(_04486_),
    .Y(_04487_),
    .B1(net3910));
 sg13g2_nand2b_1 _11074_ (.Y(_04488_),
    .B(net4568),
    .A_N(_00074_));
 sg13g2_o21ai_1 _11075_ (.B1(_04488_),
    .Y(_04489_),
    .A1(net4571),
    .A2(_00073_));
 sg13g2_nand2_1 _11076_ (.Y(_04490_),
    .A(net4573),
    .B(_01167_));
 sg13g2_or2_1 _11077_ (.X(_04491_),
    .B(_00071_),
    .A(net4571));
 sg13g2_and2_1 _11078_ (.A(_04490_),
    .B(_04491_),
    .X(_04492_));
 sg13g2_nor3_1 _11079_ (.A(net3565),
    .B(net3554),
    .C(_04492_),
    .Y(_04493_));
 sg13g2_and3_1 _11080_ (.X(_04494_),
    .A(net3567),
    .B(net3557),
    .C(_04489_));
 sg13g2_mux2_1 _11081_ (.A0(_04493_),
    .A1(_04494_),
    .S(net3893),
    .X(_04495_));
 sg13g2_o21ai_1 _11082_ (.B1(net3787),
    .Y(_04496_),
    .A1(net3904),
    .A2(_04495_));
 sg13g2_o21ai_1 _11083_ (.B1(_04479_),
    .Y(_04497_),
    .A1(_04487_),
    .A2(_04496_));
 sg13g2_a21oi_1 _11084_ (.A1(net3928),
    .A2(_04462_),
    .Y(_04498_),
    .B1(net3834));
 sg13g2_a22oi_1 _11085_ (.Y(_04499_),
    .B1(_04497_),
    .B2(_04498_),
    .A2(_04415_),
    .A1(net3839));
 sg13g2_nor3_1 _11086_ (.A(net3564),
    .B(net3553),
    .C(_04386_),
    .Y(_04500_));
 sg13g2_or4_1 _11087_ (.A(net3892),
    .B(net3564),
    .C(net3553),
    .D(_04386_),
    .X(_04501_));
 sg13g2_nand4_1 _11088_ (.B(_04124_),
    .C(_04129_),
    .A(_01169_),
    .Y(_04502_),
    .D(_04388_));
 sg13g2_nand2_1 _11089_ (.Y(_04503_),
    .A(_04501_),
    .B(_04502_));
 sg13g2_nor3_2 _11090_ (.A(net3564),
    .B(net3553),
    .C(_04380_),
    .Y(_04504_));
 sg13g2_nor3_2 _11091_ (.A(net3564),
    .B(net3553),
    .C(_04375_),
    .Y(_04505_));
 sg13g2_mux2_1 _11092_ (.A0(_04504_),
    .A1(_04505_),
    .S(net3892),
    .X(_04506_));
 sg13g2_mux4_1 _11093_ (.S0(net3908),
    .A0(_04403_),
    .A1(_04413_),
    .A2(_04506_),
    .A3(_04503_),
    .S1(net3793),
    .X(_04507_));
 sg13g2_nor3_2 _11094_ (.A(net3563),
    .B(net3552),
    .C(_04370_),
    .Y(_04508_));
 sg13g2_nor3_1 _11095_ (.A(net3563),
    .B(net3552),
    .C(_04366_),
    .Y(_04509_));
 sg13g2_nor3_2 _11096_ (.A(net3565),
    .B(net3554),
    .C(_04350_),
    .Y(_04510_));
 sg13g2_nor3_2 _11097_ (.A(net3565),
    .B(net3554),
    .C(_04346_),
    .Y(_04511_));
 sg13g2_mux2_1 _11098_ (.A0(_04510_),
    .A1(_04511_),
    .S(net3896),
    .X(_04512_));
 sg13g2_nor3_1 _11099_ (.A(net3566),
    .B(net3555),
    .C(_04341_),
    .Y(_04513_));
 sg13g2_nor3_1 _11100_ (.A(net3565),
    .B(net3554),
    .C(_04337_),
    .Y(_04514_));
 sg13g2_mux2_1 _11101_ (.A0(_04513_),
    .A1(_04514_),
    .S(net3896),
    .X(_04515_));
 sg13g2_o21ai_1 _11102_ (.B1(net4006),
    .Y(_04516_),
    .A1(\cpu.keccak_alu.registers[65] ),
    .A2(net4200));
 sg13g2_xnor2_1 _11103_ (.Y(_04517_),
    .A(_04334_),
    .B(_04499_));
 sg13g2_o21ai_1 _11104_ (.B1(_04516_),
    .Y(_04518_),
    .A1(net4006),
    .A2(_04517_));
 sg13g2_o21ai_1 _11105_ (.B1(net4218),
    .Y(_04519_),
    .A1(_01001_),
    .A2(_04518_));
 sg13g2_a21oi_1 _11106_ (.A1(_01001_),
    .A2(_04518_),
    .Y(_04520_),
    .B1(_04519_));
 sg13g2_a21oi_1 _11107_ (.A1(net4546),
    .A2(\cpu.keccak_alu.registers[193] ),
    .Y(_04521_),
    .B1(net4370));
 sg13g2_o21ai_1 _11108_ (.B1(_04521_),
    .Y(_04522_),
    .A1(net4546),
    .A2(\cpu.keccak_alu.registers[193] ));
 sg13g2_xnor2_1 _11109_ (.Y(_04523_),
    .A(\cpu.keccak_alu.registers[1] ),
    .B(\cpu.keccak_alu.registers[65] ));
 sg13g2_o21ai_1 _11110_ (.B1(net4386),
    .Y(_04524_),
    .A1(_04522_),
    .A2(_04523_));
 sg13g2_a21oi_1 _11111_ (.A1(_04522_),
    .A2(_04523_),
    .Y(_04525_),
    .B1(_04524_));
 sg13g2_o21ai_1 _11112_ (.B1(net4264),
    .Y(_04526_),
    .A1(_04520_),
    .A2(_04525_));
 sg13g2_a22oi_1 _11113_ (.Y(_04527_),
    .B1(_04326_),
    .B2(net389),
    .A2(_02482_),
    .A1(_02461_));
 sg13g2_nor2_1 _11114_ (.A(net3813),
    .B(_04527_),
    .Y(_04528_));
 sg13g2_nor2_1 _11115_ (.A(net3734),
    .B(_04528_),
    .Y(_04529_));
 sg13g2_a22oi_1 _11116_ (.Y(_00718_),
    .B1(_04526_),
    .B2(_04529_),
    .A2(net3735),
    .A1(_01005_));
 sg13g2_nor3_1 _11117_ (.A(\cpu.keccak_alu.registers[66] ),
    .B(net4189),
    .C(net4019),
    .Y(_04530_));
 sg13g2_a21oi_2 _11118_ (.B1(_04267_),
    .Y(_04531_),
    .A2(_00066_),
    .A1(net4569));
 sg13g2_a22oi_1 _11119_ (.Y(_04532_),
    .B1(_04531_),
    .B2(net4194),
    .A2(_04388_),
    .A1(\cpu.keccak_alu.registers[64] ));
 sg13g2_nand2b_1 _11120_ (.Y(_04533_),
    .B(net3831),
    .A_N(_04532_));
 sg13g2_or2_1 _11121_ (.X(_04534_),
    .B(_04533_),
    .A(_03866_));
 sg13g2_nor3_1 _11122_ (.A(net4521),
    .B(net3932),
    .C(_04534_),
    .Y(_04535_));
 sg13g2_mux2_1 _11123_ (.A0(_04143_),
    .A1(_04308_),
    .S(net3889),
    .X(_04536_));
 sg13g2_mux2_1 _11124_ (.A0(_04109_),
    .A1(_04153_),
    .S(net3879),
    .X(_04537_));
 sg13g2_mux2_1 _11125_ (.A0(_04107_),
    .A1(_04135_),
    .S(net3886),
    .X(_04538_));
 sg13g2_mux2_1 _11126_ (.A0(_04134_),
    .A1(_04191_),
    .S(net3886),
    .X(_04539_));
 sg13g2_mux4_1 _11127_ (.S0(net3906),
    .A0(_04536_),
    .A1(_04537_),
    .A2(_04538_),
    .A3(_04539_),
    .S1(net3788),
    .X(_04540_));
 sg13g2_mux2_1 _11128_ (.A0(_04168_),
    .A1(_04182_),
    .S(net3886),
    .X(_04541_));
 sg13g2_mux2_1 _11129_ (.A0(_04167_),
    .A1(_04181_),
    .S(net3886),
    .X(_04542_));
 sg13g2_and2_1 _11130_ (.A(net3877),
    .B(_04180_),
    .X(_04543_));
 sg13g2_a21oi_1 _11131_ (.A1(net3878),
    .A2(_04180_),
    .Y(_04544_),
    .B1(net3898));
 sg13g2_mux2_1 _11132_ (.A0(_04193_),
    .A1(_04203_),
    .S(net3886),
    .X(_04545_));
 sg13g2_mux2_1 _11133_ (.A0(_04166_),
    .A1(_04201_),
    .S(net3877),
    .X(_04546_));
 sg13g2_mux4_1 _11134_ (.S0(net3905),
    .A0(_04542_),
    .A1(_04543_),
    .A2(_04545_),
    .A3(_04546_),
    .S1(net3781),
    .X(_04547_));
 sg13g2_mux2_2 _11135_ (.A0(_04540_),
    .A1(_04547_),
    .S(net3923),
    .X(_04548_));
 sg13g2_mux2_1 _11136_ (.A0(_04217_),
    .A1(_04238_),
    .S(net3881),
    .X(_04549_));
 sg13g2_mux2_1 _11137_ (.A0(_04218_),
    .A1(_04239_),
    .S(net3880),
    .X(_04550_));
 sg13g2_mux2_1 _11138_ (.A0(_04234_),
    .A1(_04245_),
    .S(net3880),
    .X(_04551_));
 sg13g2_mux2_1 _11139_ (.A0(_04216_),
    .A1(_04229_),
    .S(net3887),
    .X(_04552_));
 sg13g2_mux2_1 _11140_ (.A0(_04215_),
    .A1(_04228_),
    .S(net3887),
    .X(_04553_));
 sg13g2_mux2_1 _11141_ (.A0(_04141_),
    .A1(_04254_),
    .S(net3881),
    .X(_04554_));
 sg13g2_mux2_1 _11142_ (.A0(_04142_),
    .A1(_04255_),
    .S(net3881),
    .X(_04555_));
 sg13g2_mux4_1 _11143_ (.S0(net3899),
    .A0(_04550_),
    .A1(_04551_),
    .A2(_04555_),
    .A3(_04552_),
    .S1(net3790),
    .X(_04556_));
 sg13g2_a21oi_1 _11144_ (.A1(net3891),
    .A2(_04264_),
    .Y(_04557_),
    .B1(net3909));
 sg13g2_o21ai_1 _11145_ (.B1(_04557_),
    .Y(_04558_),
    .A1(net3891),
    .A2(_04268_));
 sg13g2_nand2_1 _11146_ (.Y(_04559_),
    .A(net3880),
    .B(_04261_));
 sg13g2_o21ai_1 _11147_ (.B1(_04559_),
    .Y(_04560_),
    .A1(net3880),
    .A2(_04283_));
 sg13g2_or4_1 _11148_ (.A(net3899),
    .B(net3564),
    .C(net3553),
    .D(_04560_),
    .X(_04561_));
 sg13g2_o21ai_1 _11149_ (.B1(_04561_),
    .Y(_04562_),
    .A1(net3541),
    .A2(_04558_));
 sg13g2_a21oi_1 _11150_ (.A1(net3783),
    .A2(_04562_),
    .Y(_04563_),
    .B1(net3925));
 sg13g2_and2_1 _11151_ (.A(net3882),
    .B(_04287_),
    .X(_04564_));
 sg13g2_a21oi_1 _11152_ (.A1(net3888),
    .A2(_04279_),
    .Y(_04565_),
    .B1(_04564_));
 sg13g2_nand2b_1 _11153_ (.Y(_04566_),
    .B(_04131_),
    .A_N(_04565_));
 sg13g2_nor3_1 _11154_ (.A(net3561),
    .B(net3550),
    .C(_04275_),
    .Y(_04567_));
 sg13g2_nor4_1 _11155_ (.A(net3888),
    .B(net3561),
    .C(net3550),
    .D(_04275_),
    .Y(_04568_));
 sg13g2_a21oi_1 _11156_ (.A1(net3888),
    .A2(_04247_),
    .Y(_04569_),
    .B1(_04568_));
 sg13g2_mux2_1 _11157_ (.A0(_04566_),
    .A1(_04569_),
    .S(net3907),
    .X(_04570_));
 sg13g2_nor4_1 _11158_ (.A(net3637),
    .B(net3579),
    .C(net3570),
    .D(_04560_),
    .Y(_04571_));
 sg13g2_nor4_1 _11159_ (.A(net3637),
    .B(net3579),
    .C(net3570),
    .D(_04565_),
    .Y(_04572_));
 sg13g2_o21ai_1 _11160_ (.B1(_04563_),
    .Y(_04573_),
    .A1(net3783),
    .A2(_04570_));
 sg13g2_mux2_1 _11161_ (.A0(_04192_),
    .A1(_04306_),
    .S(net3886),
    .X(_04574_));
 sg13g2_and2_1 _11162_ (.A(net3879),
    .B(_04179_),
    .X(_04575_));
 sg13g2_mux2_1 _11163_ (.A0(_04178_),
    .A1(_04307_),
    .S(net3878),
    .X(_04576_));
 sg13g2_mux4_1 _11164_ (.S0(net3897),
    .A0(_04546_),
    .A1(_04574_),
    .A2(_04575_),
    .A3(_04576_),
    .S1(net3789),
    .X(_04577_));
 sg13g2_a21oi_1 _11165_ (.A1(net3925),
    .A2(_04556_),
    .Y(_04578_),
    .B1(net3833));
 sg13g2_a22oi_1 _11166_ (.Y(_04579_),
    .B1(_04573_),
    .B2(_04578_),
    .A2(_04548_),
    .A1(net3838));
 sg13g2_xnor2_1 _11167_ (.Y(_04580_),
    .A(_04535_),
    .B(_04579_));
 sg13g2_a21oi_1 _11168_ (.A1(net4019),
    .A2(_04580_),
    .Y(_04581_),
    .B1(_04530_));
 sg13g2_xor2_1 _11169_ (.B(_04581_),
    .A(\cpu.keccak_alu.registers[2] ),
    .X(_04582_));
 sg13g2_o21ai_1 _11170_ (.B1(net4209),
    .Y(_04583_),
    .A1(net4533),
    .A2(\cpu.keccak_alu.registers[194] ));
 sg13g2_a21oi_1 _11171_ (.A1(net4532),
    .A2(\cpu.keccak_alu.registers[194] ),
    .Y(_04584_),
    .B1(_04583_));
 sg13g2_xor2_1 _11172_ (.B(\cpu.keccak_alu.registers[66] ),
    .A(\cpu.keccak_alu.registers[2] ),
    .X(_04585_));
 sg13g2_a21oi_1 _11173_ (.A1(_04584_),
    .A2(_04585_),
    .Y(_04586_),
    .B1(net4218));
 sg13g2_o21ai_1 _11174_ (.B1(_04586_),
    .Y(_04587_),
    .A1(_04584_),
    .A2(_04585_));
 sg13g2_o21ai_1 _11175_ (.B1(_04587_),
    .Y(_04588_),
    .A1(net4384),
    .A2(_04582_));
 sg13g2_a22oi_1 _11176_ (.Y(_04589_),
    .B1(_04326_),
    .B2(net282),
    .A2(net3754),
    .A1(_02463_));
 sg13g2_o21ai_1 _11177_ (.B1(net3739),
    .Y(_04590_),
    .A1(net3813),
    .A2(_04589_));
 sg13g2_a21oi_1 _11178_ (.A1(net4264),
    .A2(_04588_),
    .Y(_04591_),
    .B1(_04590_));
 sg13g2_a21oi_1 _11179_ (.A1(_01013_),
    .A2(net3734),
    .Y(_00719_),
    .B1(_04591_));
 sg13g2_a21oi_1 _11180_ (.A1(net4572),
    .A2(_01166_),
    .Y(_04592_),
    .B1(_04482_));
 sg13g2_nor2_1 _11181_ (.A(net3826),
    .B(_04592_),
    .Y(_04593_));
 sg13g2_nor2_1 _11182_ (.A(net4200),
    .B(_04331_),
    .Y(_04594_));
 sg13g2_a21oi_1 _11183_ (.A1(net4200),
    .A2(_04593_),
    .Y(_04595_),
    .B1(_04594_));
 sg13g2_nand2b_1 _11184_ (.Y(_04596_),
    .B(_03865_),
    .A_N(_04595_));
 sg13g2_nor3_1 _11185_ (.A(net4523),
    .B(net3933),
    .C(_04596_),
    .Y(_04597_));
 sg13g2_mux2_1 _11186_ (.A0(_04510_),
    .A1(_04514_),
    .S(net3884),
    .X(_04598_));
 sg13g2_mux2_1 _11187_ (.A0(_04347_),
    .A1(_04362_),
    .S(net3892),
    .X(_04599_));
 sg13g2_mux2_2 _11188_ (.A0(_04361_),
    .A1(_04508_),
    .S(net3890),
    .X(_04600_));
 sg13g2_mux2_1 _11189_ (.A0(_04367_),
    .A1(_04402_),
    .S(net3890),
    .X(_04601_));
 sg13g2_mux4_1 _11190_ (.S0(net3911),
    .A0(_04598_),
    .A1(_04599_),
    .A2(_04600_),
    .A3(_04601_),
    .S1(net3792),
    .X(_04602_));
 sg13g2_nand2b_1 _11191_ (.Y(_04603_),
    .B(net3922),
    .A_N(_04602_));
 sg13g2_mux2_1 _11192_ (.A0(_04401_),
    .A1(_04411_),
    .S(net3890),
    .X(_04604_));
 sg13g2_mux2_1 _11193_ (.A0(_04381_),
    .A1(_04407_),
    .S(net3883),
    .X(_04605_));
 sg13g2_mux2_1 _11194_ (.A0(_04376_),
    .A1(_04387_),
    .S(net3890),
    .X(_04606_));
 sg13g2_nor3_1 _11195_ (.A(net4567),
    .B(net4541),
    .C(_00069_),
    .Y(_04607_));
 sg13g2_and2_1 _11196_ (.A(_04389_),
    .B(_04607_),
    .X(_04608_));
 sg13g2_a21o_1 _11197_ (.A2(_04606_),
    .A1(net3903),
    .B1(_04608_),
    .X(_04609_));
 sg13g2_mux4_1 _11198_ (.S0(net3890),
    .A0(_04401_),
    .A1(_04411_),
    .A2(_04412_),
    .A3(_04504_),
    .S1(net3908),
    .X(_04610_));
 sg13g2_nor2_1 _11199_ (.A(net3792),
    .B(_04610_),
    .Y(_04611_));
 sg13g2_mux2_1 _11200_ (.A0(_04500_),
    .A1(_04505_),
    .S(net3883),
    .X(_04612_));
 sg13g2_nor3_1 _11201_ (.A(_00069_),
    .B(net4576),
    .C(net3542),
    .Y(_04613_));
 sg13g2_a22oi_1 _11202_ (.Y(_04614_),
    .B1(_04613_),
    .B2(net4093),
    .A2(_04612_),
    .A1(net3903));
 sg13g2_a221oi_1 _11203_ (.B2(net4093),
    .C1(net3785),
    .B1(_04613_),
    .A1(net3903),
    .Y(_04615_),
    .A2(_04612_));
 sg13g2_o21ai_1 _11204_ (.B1(net3928),
    .Y(_04616_),
    .A1(_04611_),
    .A2(_04615_));
 sg13g2_and3_1 _11205_ (.X(_04617_),
    .A(_03875_),
    .B(_04603_),
    .C(_04616_));
 sg13g2_mux2_1 _11206_ (.A0(_04419_),
    .A1(_04433_),
    .S(net3895),
    .X(_04618_));
 sg13g2_mux2_1 _11207_ (.A0(_04458_),
    .A1(_04513_),
    .S(net3896),
    .X(_04619_));
 sg13g2_mux2_1 _11208_ (.A0(_04442_),
    .A1(_04450_),
    .S(net3895),
    .X(_04620_));
 sg13g2_mux2_1 _11209_ (.A0(_04422_),
    .A1(_04452_),
    .S(net3885),
    .X(_04621_));
 sg13g2_mux4_1 _11210_ (.S0(net3910),
    .A0(_04618_),
    .A1(_04619_),
    .A2(_04620_),
    .A3(_04621_),
    .S1(net3786),
    .X(_04622_));
 sg13g2_nor2_1 _11211_ (.A(net3922),
    .B(_04622_),
    .Y(_04623_));
 sg13g2_mux2_1 _11212_ (.A0(_04467_),
    .A1(_04474_),
    .S(net3893),
    .X(_04624_));
 sg13g2_mux2_1 _11213_ (.A0(_04444_),
    .A1(_04470_),
    .S(net3884),
    .X(_04625_));
 sg13g2_mux2_1 _11214_ (.A0(_04624_),
    .A1(_04625_),
    .S(net3911),
    .X(_04626_));
 sg13g2_nor2_1 _11215_ (.A(net3894),
    .B(_04494_),
    .Y(_04627_));
 sg13g2_nor2_1 _11216_ (.A(net3884),
    .B(_04475_),
    .Y(_04628_));
 sg13g2_o21ai_1 _11217_ (.B1(net3910),
    .Y(_04629_),
    .A1(_04627_),
    .A2(_04628_));
 sg13g2_a21oi_1 _11218_ (.A1(net3893),
    .A2(_04493_),
    .Y(_04630_),
    .B1(net3910));
 sg13g2_nand2b_1 _11219_ (.Y(_04631_),
    .B(net3884),
    .A_N(_04484_));
 sg13g2_a21oi_1 _11220_ (.A1(_04630_),
    .A2(_04631_),
    .Y(_04632_),
    .B1(net3791));
 sg13g2_a221oi_1 _11221_ (.B2(_04632_),
    .C1(net3929),
    .B1(_04629_),
    .A1(net3791),
    .Y(_04633_),
    .A2(_04626_));
 sg13g2_nor3_2 _11222_ (.A(net3834),
    .B(_04623_),
    .C(_04633_),
    .Y(_04634_));
 sg13g2_o21ai_1 _11223_ (.B1(_04597_),
    .Y(_04635_),
    .A1(_04617_),
    .A2(_04634_));
 sg13g2_or3_1 _11224_ (.A(_04597_),
    .B(_04617_),
    .C(_04634_),
    .X(_04636_));
 sg13g2_and2_1 _11225_ (.A(net4019),
    .B(_04636_),
    .X(_04637_));
 sg13g2_nor2_1 _11226_ (.A(\cpu.keccak_alu.registers[67] ),
    .B(net4177),
    .Y(_04638_));
 sg13g2_nor2_1 _11227_ (.A(net4020),
    .B(_04638_),
    .Y(_04639_));
 sg13g2_a21oi_1 _11228_ (.A1(_04635_),
    .A2(_04636_),
    .Y(_04640_),
    .B1(net4005));
 sg13g2_a221oi_1 _11229_ (.B2(net4007),
    .C1(\cpu.keccak_alu.registers[3] ),
    .B1(_04638_),
    .A1(_04635_),
    .Y(_04641_),
    .A2(_04637_));
 sg13g2_nor3_1 _11230_ (.A(_01017_),
    .B(_04639_),
    .C(_04640_),
    .Y(_04642_));
 sg13g2_or3_1 _11231_ (.A(net4386),
    .B(_04641_),
    .C(_04642_),
    .X(_04643_));
 sg13g2_o21ai_1 _11232_ (.B1(net4210),
    .Y(_04644_),
    .A1(net4530),
    .A2(\cpu.keccak_alu.registers[195] ));
 sg13g2_a21oi_1 _11233_ (.A1(net4530),
    .A2(\cpu.keccak_alu.registers[195] ),
    .Y(_04645_),
    .B1(_04644_));
 sg13g2_xor2_1 _11234_ (.B(\cpu.keccak_alu.registers[67] ),
    .A(\cpu.keccak_alu.registers[3] ),
    .X(_04646_));
 sg13g2_a21oi_1 _11235_ (.A1(_04645_),
    .A2(_04646_),
    .Y(_04647_),
    .B1(net4219));
 sg13g2_o21ai_1 _11236_ (.B1(_04647_),
    .Y(_04648_),
    .A1(_04645_),
    .A2(_04646_));
 sg13g2_a21o_1 _11237_ (.A2(_04648_),
    .A1(_04643_),
    .B1(net4321),
    .X(_04649_));
 sg13g2_a22oi_1 _11238_ (.Y(_04650_),
    .B1(_04326_),
    .B2(net453),
    .A2(net3754),
    .A1(_02465_));
 sg13g2_nor2_1 _11239_ (.A(net3813),
    .B(_04650_),
    .Y(_04651_));
 sg13g2_nor2_1 _11240_ (.A(net3734),
    .B(_04651_),
    .Y(_04652_));
 sg13g2_a22oi_1 _11241_ (.Y(_00720_),
    .B1(_04649_),
    .B2(_04652_),
    .A2(net3734),
    .A1(_01022_));
 sg13g2_o21ai_1 _11242_ (.B1(net4211),
    .Y(_04653_),
    .A1(net4522),
    .A2(\cpu.keccak_alu.registers[196] ));
 sg13g2_a21oi_1 _11243_ (.A1(net4522),
    .A2(\cpu.keccak_alu.registers[196] ),
    .Y(_04654_),
    .B1(_04653_));
 sg13g2_xor2_1 _11244_ (.B(\cpu.keccak_alu.registers[68] ),
    .A(\cpu.keccak_alu.registers[4] ),
    .X(_04655_));
 sg13g2_o21ai_1 _11245_ (.B1(net4382),
    .Y(_04656_),
    .A1(_04654_),
    .A2(_04655_));
 sg13g2_a21oi_1 _11246_ (.A1(_04654_),
    .A2(_04655_),
    .Y(_04657_),
    .B1(_04656_));
 sg13g2_nand3b_1 _11247_ (.B(net4522),
    .C(net4004),
    .Y(_04658_),
    .A_N(\cpu.keccak_alu.registers[68] ));
 sg13g2_nand2_1 _11248_ (.Y(_04659_),
    .A(_04263_),
    .B(_04266_));
 sg13g2_nor2_1 _11249_ (.A(net4538),
    .B(_04659_),
    .Y(_04660_));
 sg13g2_a21oi_1 _11250_ (.A1(net4538),
    .A2(_04531_),
    .Y(_04661_),
    .B1(_04660_));
 sg13g2_nor3_1 _11251_ (.A(net4534),
    .B(net3824),
    .C(_04661_),
    .Y(_04662_));
 sg13g2_a21oi_2 _11252_ (.B1(_04662_),
    .Y(_04663_),
    .A2(_04303_),
    .A1(net4531));
 sg13g2_or3_1 _11253_ (.A(net4527),
    .B(net4521),
    .C(_04663_),
    .X(_04664_));
 sg13g2_or2_1 _11254_ (.X(_04665_),
    .B(_04664_),
    .A(net3931));
 sg13g2_mux2_1 _11255_ (.A0(_04171_),
    .A1(_04205_),
    .S(net3897),
    .X(_04666_));
 sg13g2_mux4_1 _11256_ (.S0(net3877),
    .A0(_04168_),
    .A1(_04170_),
    .A2(_04202_),
    .A3(_04204_),
    .S1(net3897),
    .X(_04667_));
 sg13g2_nand2_1 _11257_ (.Y(_04668_),
    .A(net3782),
    .B(_04667_));
 sg13g2_and2_1 _11258_ (.A(net3897),
    .B(_04183_),
    .X(_04669_));
 sg13g2_a21o_1 _11259_ (.A2(_04183_),
    .A1(net3898),
    .B1(net3781),
    .X(_04670_));
 sg13g2_mux2_1 _11260_ (.A0(_04112_),
    .A1(_04158_),
    .S(net3897),
    .X(_04671_));
 sg13g2_mux2_1 _11261_ (.A0(_04136_),
    .A1(_04195_),
    .S(net3905),
    .X(_04672_));
 sg13g2_mux4_1 _11262_ (.S0(net3897),
    .A0(_04112_),
    .A1(_04158_),
    .A2(_04195_),
    .A3(_04136_),
    .S1(net3788),
    .X(_04673_));
 sg13g2_mux4_1 _11263_ (.S0(net3788),
    .A0(_04666_),
    .A1(_04669_),
    .A2(_04671_),
    .A3(_04672_),
    .S1(net3913),
    .X(_04674_));
 sg13g2_nand2_1 _11264_ (.Y(_04675_),
    .A(net3838),
    .B(_04674_));
 sg13g2_mux4_1 _11265_ (.S0(net3880),
    .A0(_04216_),
    .A1(_04218_),
    .A2(_04239_),
    .A3(_04234_),
    .S1(net3900),
    .X(_04676_));
 sg13g2_mux4_1 _11266_ (.S0(net3783),
    .A0(_04145_),
    .A1(_04219_),
    .A2(_04256_),
    .A3(_04251_),
    .S1(net3899),
    .X(_04677_));
 sg13g2_nor2_1 _11267_ (.A(net3916),
    .B(_04677_),
    .Y(_04678_));
 sg13g2_mux2_1 _11268_ (.A0(_04248_),
    .A1(_04290_),
    .S(net3900),
    .X(_04679_));
 sg13g2_o21ai_1 _11269_ (.B1(net3899),
    .Y(_04680_),
    .A1(net3541),
    .A2(_04265_));
 sg13g2_o21ai_1 _11270_ (.B1(net3907),
    .Y(_04681_),
    .A1(net3541),
    .A2(_04288_));
 sg13g2_and2_1 _11271_ (.A(net3784),
    .B(_04681_),
    .X(_04682_));
 sg13g2_a221oi_1 _11272_ (.B2(_04682_),
    .C1(net3925),
    .B1(_04680_),
    .A1(net3790),
    .Y(_04683_),
    .A2(_04679_));
 sg13g2_or3_1 _11273_ (.A(net3833),
    .B(_04678_),
    .C(_04683_),
    .X(_04684_));
 sg13g2_nand3_1 _11274_ (.B(_04675_),
    .C(_04684_),
    .A(_04665_),
    .Y(_04685_));
 sg13g2_or4_1 _11275_ (.A(net4518),
    .B(net4515),
    .C(_04664_),
    .D(_04675_),
    .X(_04686_));
 sg13g2_nand3_1 _11276_ (.B(_04685_),
    .C(_04686_),
    .A(net4018),
    .Y(_04687_));
 sg13g2_a21oi_1 _11277_ (.A1(_04658_),
    .A2(_04687_),
    .Y(_04688_),
    .B1(_01026_));
 sg13g2_and3_1 _11278_ (.X(_04689_),
    .A(_01026_),
    .B(_04658_),
    .C(_04687_));
 sg13g2_nor3_1 _11279_ (.A(net4382),
    .B(_04688_),
    .C(_04689_),
    .Y(_04690_));
 sg13g2_o21ai_1 _11280_ (.B1(net4265),
    .Y(_04691_),
    .A1(_04657_),
    .A2(_04690_));
 sg13g2_a22oi_1 _11281_ (.Y(_04692_),
    .B1(_04326_),
    .B2(net484),
    .A2(net3754),
    .A1(_02467_));
 sg13g2_nor2_1 _11282_ (.A(net3814),
    .B(_04692_),
    .Y(_04693_));
 sg13g2_nor2_1 _11283_ (.A(net3732),
    .B(_04693_),
    .Y(_04694_));
 sg13g2_a22oi_1 _11284_ (.Y(_00721_),
    .B1(_04691_),
    .B2(_04694_),
    .A2(net3732),
    .A1(_01030_));
 sg13g2_o21ai_1 _11285_ (.B1(net4211),
    .Y(_04695_),
    .A1(net4517),
    .A2(\cpu.keccak_alu.registers[197] ));
 sg13g2_a21oi_1 _11286_ (.A1(net4517),
    .A2(\cpu.keccak_alu.registers[197] ),
    .Y(_04696_),
    .B1(_04695_));
 sg13g2_xor2_1 _11287_ (.B(\cpu.keccak_alu.registers[69] ),
    .A(\cpu.keccak_alu.registers[5] ),
    .X(_04697_));
 sg13g2_a21oi_1 _11288_ (.A1(_04696_),
    .A2(_04697_),
    .Y(_04698_),
    .B1(net4220));
 sg13g2_o21ai_1 _11289_ (.B1(_04698_),
    .Y(_04699_),
    .A1(_04696_),
    .A2(_04697_));
 sg13g2_o21ai_1 _11290_ (.B1(net4532),
    .Y(_04700_),
    .A1(net4547),
    .A2(_04331_));
 sg13g2_a21oi_1 _11291_ (.A1(_04481_),
    .A2(_04491_),
    .Y(_04701_),
    .B1(net3826));
 sg13g2_mux2_1 _11292_ (.A0(_04593_),
    .A1(_04701_),
    .S(net4200),
    .X(_04702_));
 sg13g2_o21ai_1 _11293_ (.B1(_04700_),
    .Y(_04703_),
    .A1(net4532),
    .A2(_04702_));
 sg13g2_nand2b_1 _11294_ (.Y(_04704_),
    .B(net4175),
    .A_N(_04703_));
 sg13g2_nor2_1 _11295_ (.A(net4524),
    .B(_04704_),
    .Y(_04705_));
 sg13g2_nand2_1 _11296_ (.Y(_04706_),
    .A(net4089),
    .B(_04705_));
 sg13g2_mux4_1 _11297_ (.S0(net3893),
    .A0(_04440_),
    .A1(_04442_),
    .A2(_04474_),
    .A3(_04470_),
    .S1(net3902),
    .X(_04707_));
 sg13g2_a21o_1 _11298_ (.A2(_04707_),
    .A1(net3791),
    .B1(net3929),
    .X(_04708_));
 sg13g2_mux2_1 _11299_ (.A0(_04477_),
    .A1(_04495_),
    .S(net3904),
    .X(_04709_));
 sg13g2_a21oi_2 _11300_ (.B1(_04708_),
    .Y(_04710_),
    .A2(_04709_),
    .A1(net3787));
 sg13g2_mux4_1 _11301_ (.S0(net3895),
    .A0(_04422_),
    .A1(_04424_),
    .A2(_04450_),
    .A3(_04452_),
    .S1(net3902),
    .X(_04711_));
 sg13g2_mux4_1 _11302_ (.S0(net3902),
    .A0(_04426_),
    .A1(_04454_),
    .A2(_04515_),
    .A3(_04460_),
    .S1(net3791),
    .X(_04712_));
 sg13g2_o21ai_1 _11303_ (.B1(net3777),
    .Y(_04713_),
    .A1(net3918),
    .A2(_04712_));
 sg13g2_a21oi_2 _11304_ (.B1(net3908),
    .Y(_04714_),
    .A2(_04502_),
    .A1(_04501_));
 sg13g2_mux4_1 _11305_ (.S0(net3890),
    .A0(_04411_),
    .A1(_04412_),
    .A2(_04504_),
    .A3(_04505_),
    .S1(net3908),
    .X(_04715_));
 sg13g2_mux2_1 _11306_ (.A0(_04714_),
    .A1(_04715_),
    .S(net3785),
    .X(_04716_));
 sg13g2_mux4_1 _11307_ (.S0(net3892),
    .A0(_04360_),
    .A1(_04361_),
    .A2(_04510_),
    .A3(_04511_),
    .S1(net3903),
    .X(_04717_));
 sg13g2_mux4_1 _11308_ (.S0(net3890),
    .A0(_04400_),
    .A1(_04401_),
    .A2(_04508_),
    .A3(_04509_),
    .S1(net3903),
    .X(_04718_));
 sg13g2_mux2_1 _11309_ (.A0(_04717_),
    .A1(_04718_),
    .S(net3793),
    .X(_04719_));
 sg13g2_mux4_1 _11310_ (.S0(net3785),
    .A0(_04714_),
    .A1(_04715_),
    .A2(_04718_),
    .A3(_04717_),
    .S1(net3919),
    .X(_04720_));
 sg13g2_nand2_1 _11311_ (.Y(_04721_),
    .A(net3840),
    .B(_04720_));
 sg13g2_o21ai_1 _11312_ (.B1(_04721_),
    .Y(_04722_),
    .A1(_04710_),
    .A2(_04713_));
 sg13g2_o21ai_1 _11313_ (.B1(net4004),
    .Y(_04723_),
    .A1(\cpu.keccak_alu.registers[69] ),
    .A2(net4162));
 sg13g2_xnor2_1 _11314_ (.Y(_04724_),
    .A(_04706_),
    .B(_04722_));
 sg13g2_o21ai_1 _11315_ (.B1(_04723_),
    .Y(_04725_),
    .A1(net4008),
    .A2(_04724_));
 sg13g2_xor2_1 _11316_ (.B(_04725_),
    .A(\cpu.keccak_alu.registers[5] ),
    .X(_04726_));
 sg13g2_o21ai_1 _11317_ (.B1(_04699_),
    .Y(_04727_),
    .A1(net4383),
    .A2(_04726_));
 sg13g2_nor2_1 _11318_ (.A(net181),
    .B(net3698),
    .Y(_04728_));
 sg13g2_a21oi_1 _11319_ (.A1(net4344),
    .A2(net3698),
    .Y(_04729_),
    .B1(_04728_));
 sg13g2_a221oi_1 _11320_ (.B2(net3819),
    .C1(net3731),
    .B1(_04729_),
    .A1(net4263),
    .Y(_04730_),
    .A2(_04727_));
 sg13g2_a21oi_1 _11321_ (.A1(_01038_),
    .A2(net3731),
    .Y(_00722_),
    .B1(_04730_));
 sg13g2_o21ai_1 _11322_ (.B1(_04262_),
    .Y(_04731_),
    .A1(net4562),
    .A2(_01167_));
 sg13g2_mux2_1 _11323_ (.A0(_04659_),
    .A1(_04731_),
    .S(net4196),
    .X(_04732_));
 sg13g2_nor2_1 _11324_ (.A(net3824),
    .B(_04732_),
    .Y(_04733_));
 sg13g2_nor2_1 _11325_ (.A(net4182),
    .B(_04533_),
    .Y(_04734_));
 sg13g2_a21oi_1 _11326_ (.A1(net4183),
    .A2(_04733_),
    .Y(_04735_),
    .B1(_04734_));
 sg13g2_or2_1 _11327_ (.X(_04736_),
    .B(_04735_),
    .A(net4525));
 sg13g2_nand2b_1 _11328_ (.Y(_04737_),
    .B(net4166),
    .A_N(_04736_));
 sg13g2_nor2_1 _11329_ (.A(net3932),
    .B(_04737_),
    .Y(_04738_));
 sg13g2_mux4_1 _11330_ (.S0(net3887),
    .A0(_04215_),
    .A1(_04228_),
    .A2(_04238_),
    .A3(_04217_),
    .S1(net3899),
    .X(_04739_));
 sg13g2_mux4_1 _11331_ (.S0(net3782),
    .A0(_04536_),
    .A1(_04553_),
    .A2(_04554_),
    .A3(_04549_),
    .S1(net3899),
    .X(_04740_));
 sg13g2_mux2_1 _11332_ (.A0(_04571_),
    .A1(_04572_),
    .S(net3907),
    .X(_04741_));
 sg13g2_mux4_1 _11333_ (.S0(net3887),
    .A0(_04246_),
    .A1(_04250_),
    .A2(_04567_),
    .A3(_04247_),
    .S1(net3900),
    .X(_04742_));
 sg13g2_mux2_1 _11334_ (.A0(_04741_),
    .A1(_04742_),
    .S(net3790),
    .X(_04743_));
 sg13g2_nor2_1 _11335_ (.A(net3925),
    .B(_04743_),
    .Y(_04744_));
 sg13g2_o21ai_1 _11336_ (.B1(net3773),
    .Y(_04745_),
    .A1(net3914),
    .A2(_04740_));
 sg13g2_mux4_1 _11337_ (.S0(net3898),
    .A0(_04133_),
    .A1(_04311_),
    .A2(_04312_),
    .A3(_04309_),
    .S1(net3879),
    .X(_04746_));
 sg13g2_mux4_1 _11338_ (.S0(net3886),
    .A0(_04134_),
    .A1(_04191_),
    .A2(_04192_),
    .A3(_04306_),
    .S1(net3906),
    .X(_04747_));
 sg13g2_mux2_1 _11339_ (.A0(_04746_),
    .A1(_04747_),
    .S(net3789),
    .X(_04748_));
 sg13g2_and3_1 _11340_ (.X(_04749_),
    .A(net3898),
    .B(net3878),
    .C(_04179_));
 sg13g2_mux4_1 _11341_ (.S0(net3906),
    .A0(_04166_),
    .A1(_04178_),
    .A2(_04201_),
    .A3(_04307_),
    .S1(net3878),
    .X(_04750_));
 sg13g2_mux2_1 _11342_ (.A0(_04749_),
    .A1(_04750_),
    .S(net3782),
    .X(_04751_));
 sg13g2_mux4_1 _11343_ (.S0(net3789),
    .A0(_04746_),
    .A1(_04747_),
    .A2(_04750_),
    .A3(_04749_),
    .S1(net3923),
    .X(_04752_));
 sg13g2_nand2_1 _11344_ (.Y(_04753_),
    .A(net3837),
    .B(_04752_));
 sg13g2_o21ai_1 _11345_ (.B1(_04753_),
    .Y(_04754_),
    .A1(_04744_),
    .A2(_04745_));
 sg13g2_a21oi_1 _11346_ (.A1(_01043_),
    .A2(net4514),
    .Y(_04755_),
    .B1(net4016));
 sg13g2_xnor2_1 _11347_ (.Y(_04756_),
    .A(_04738_),
    .B(_04754_));
 sg13g2_a21oi_1 _11348_ (.A1(net4016),
    .A2(_04756_),
    .Y(_04757_),
    .B1(_04755_));
 sg13g2_xnor2_1 _11349_ (.Y(_04758_),
    .A(\cpu.keccak_alu.registers[6] ),
    .B(_04757_));
 sg13g2_o21ai_1 _11350_ (.B1(net4211),
    .Y(_04759_),
    .A1(net4513),
    .A2(\cpu.keccak_alu.registers[198] ));
 sg13g2_a21oi_1 _11351_ (.A1(net4515),
    .A2(\cpu.keccak_alu.registers[198] ),
    .Y(_04760_),
    .B1(_04759_));
 sg13g2_xor2_1 _11352_ (.B(\cpu.keccak_alu.registers[70] ),
    .A(\cpu.keccak_alu.registers[6] ),
    .X(_04761_));
 sg13g2_a21oi_1 _11353_ (.A1(_04760_),
    .A2(_04761_),
    .Y(_04762_),
    .B1(net4220));
 sg13g2_o21ai_1 _11354_ (.B1(_04762_),
    .Y(_04763_),
    .A1(_04760_),
    .A2(_04761_));
 sg13g2_o21ai_1 _11355_ (.B1(_04763_),
    .Y(_04764_),
    .A1(net4383),
    .A2(_04758_));
 sg13g2_a22oi_1 _11356_ (.Y(_04765_),
    .B1(_04326_),
    .B2(net251),
    .A2(net3754),
    .A1(_02470_));
 sg13g2_o21ai_1 _11357_ (.B1(net3739),
    .Y(_04766_),
    .A1(net3814),
    .A2(_04765_));
 sg13g2_a21oi_1 _11358_ (.A1(net4263),
    .A2(_04764_),
    .Y(_04767_),
    .B1(_04766_));
 sg13g2_a21oi_1 _11359_ (.A1(_01048_),
    .A2(net3732),
    .Y(_00723_),
    .B1(_04767_));
 sg13g2_nor3_1 _11360_ (.A(\cpu.keccak_alu.registers[71] ),
    .B(_01055_),
    .C(net4015),
    .Y(_04768_));
 sg13g2_o21ai_1 _11361_ (.B1(_04490_),
    .Y(_04769_),
    .A1(net4568),
    .A2(_00073_));
 sg13g2_nand2_1 _11362_ (.Y(_04770_),
    .A(net3832),
    .B(_04769_));
 sg13g2_nand2_1 _11363_ (.Y(_04771_),
    .A(net4545),
    .B(_04701_));
 sg13g2_o21ai_1 _11364_ (.B1(_04771_),
    .Y(_04772_),
    .A1(net4545),
    .A2(_04770_));
 sg13g2_nor2_1 _11365_ (.A(net4532),
    .B(_04772_),
    .Y(_04773_));
 sg13g2_a21oi_1 _11366_ (.A1(net4532),
    .A2(_04595_),
    .Y(_04774_),
    .B1(_04773_));
 sg13g2_inv_1 _11367_ (.Y(_04775_),
    .A(_04774_));
 sg13g2_nor3_1 _11368_ (.A(net4529),
    .B(net4524),
    .C(_04775_),
    .Y(_04776_));
 sg13g2_nand2_1 _11369_ (.Y(_04777_),
    .A(net4089),
    .B(_04776_));
 sg13g2_mux4_1 _11370_ (.S0(net3893),
    .A0(_04467_),
    .A1(_04474_),
    .A2(_04494_),
    .A3(_04475_),
    .S1(net3902),
    .X(_04778_));
 sg13g2_nand2_1 _11371_ (.Y(_04779_),
    .A(net3786),
    .B(_04778_));
 sg13g2_mux4_1 _11372_ (.S0(net3912),
    .A0(_04440_),
    .A1(_04450_),
    .A2(_04473_),
    .A3(_04442_),
    .S1(net3884),
    .X(_04780_));
 sg13g2_a21oi_1 _11373_ (.A1(net3791),
    .A2(_04780_),
    .Y(_04781_),
    .B1(net3929));
 sg13g2_mux4_1 _11374_ (.S0(net3786),
    .A0(_04598_),
    .A1(_04618_),
    .A2(_04619_),
    .A3(_04621_),
    .S1(net3902),
    .X(_04782_));
 sg13g2_mux4_1 _11375_ (.S0(net3884),
    .A0(_04422_),
    .A1(_04452_),
    .A2(_04456_),
    .A3(_04424_),
    .S1(net3910),
    .X(_04783_));
 sg13g2_or2_1 _11376_ (.X(_04784_),
    .B(_04782_),
    .A(net3921));
 sg13g2_a21oi_1 _11377_ (.A1(_04779_),
    .A2(_04781_),
    .Y(_04785_),
    .B1(net3834));
 sg13g2_mux4_1 _11378_ (.S0(net3909),
    .A0(_04400_),
    .A1(_04411_),
    .A2(_04509_),
    .A3(_04401_),
    .S1(net3883),
    .X(_04786_));
 sg13g2_mux4_1 _11379_ (.S0(net3908),
    .A0(_04360_),
    .A1(_04508_),
    .A2(_04511_),
    .A3(_04361_),
    .S1(net3883),
    .X(_04787_));
 sg13g2_mux2_1 _11380_ (.A0(_04786_),
    .A1(_04787_),
    .S(net3787),
    .X(_04788_));
 sg13g2_mux4_1 _11381_ (.S0(net3892),
    .A0(_04412_),
    .A1(_04504_),
    .A2(_04505_),
    .A3(_04500_),
    .S1(net3908),
    .X(_04789_));
 sg13g2_nor4_1 _11382_ (.A(net4174),
    .B(net4576),
    .C(_03878_),
    .D(net3542),
    .Y(_04790_));
 sg13g2_a21o_1 _11383_ (.A2(_04789_),
    .A1(net3785),
    .B1(_04790_),
    .X(_04791_));
 sg13g2_mux2_1 _11384_ (.A0(_04788_),
    .A1(_04791_),
    .S(net3926),
    .X(_04792_));
 sg13g2_a22oi_1 _11385_ (.Y(_04793_),
    .B1(_04792_),
    .B2(net3839),
    .A2(_04785_),
    .A1(_04784_));
 sg13g2_xor2_1 _11386_ (.B(_04793_),
    .A(_04777_),
    .X(_04794_));
 sg13g2_a21oi_1 _11387_ (.A1(net4015),
    .A2(_04794_),
    .Y(_04795_),
    .B1(_04768_));
 sg13g2_xor2_1 _11388_ (.B(_04795_),
    .A(\cpu.keccak_alu.registers[7] ),
    .X(_04796_));
 sg13g2_o21ai_1 _11389_ (.B1(net4207),
    .Y(_04797_),
    .A1(net4512),
    .A2(\cpu.keccak_alu.registers[199] ));
 sg13g2_a21oi_1 _11390_ (.A1(net4512),
    .A2(\cpu.keccak_alu.registers[199] ),
    .Y(_04798_),
    .B1(_04797_));
 sg13g2_xor2_1 _11391_ (.B(\cpu.keccak_alu.registers[71] ),
    .A(\cpu.keccak_alu.registers[7] ),
    .X(_04799_));
 sg13g2_o21ai_1 _11392_ (.B1(net4378),
    .Y(_04800_),
    .A1(_04798_),
    .A2(_04799_));
 sg13g2_a21o_1 _11393_ (.A2(_04799_),
    .A1(_04798_),
    .B1(_04800_),
    .X(_04801_));
 sg13g2_o21ai_1 _11394_ (.B1(_04801_),
    .Y(_04802_),
    .A1(net4378),
    .A2(_04796_));
 sg13g2_nor2_1 _11395_ (.A(net156),
    .B(net3698),
    .Y(_04803_));
 sg13g2_a21oi_1 _11396_ (.A1(net4337),
    .A2(net3698),
    .Y(_04804_),
    .B1(_04803_));
 sg13g2_a221oi_1 _11397_ (.B2(net3818),
    .C1(net3728),
    .B1(_04804_),
    .A1(net4258),
    .Y(_04805_),
    .A2(_04802_));
 sg13g2_a21oi_1 _11398_ (.A1(_01057_),
    .A2(net3728),
    .Y(_00724_),
    .B1(_04805_));
 sg13g2_a21oi_1 _11399_ (.A1(net4510),
    .A2(\cpu.keccak_alu.registers[200] ),
    .Y(_04806_),
    .B1(net4369));
 sg13g2_o21ai_1 _11400_ (.B1(_04806_),
    .Y(_04807_),
    .A1(net4510),
    .A2(\cpu.keccak_alu.registers[200] ));
 sg13g2_xor2_1 _11401_ (.B(\cpu.keccak_alu.registers[72] ),
    .A(\cpu.keccak_alu.registers[8] ),
    .X(_04808_));
 sg13g2_xnor2_1 _11402_ (.Y(_04809_),
    .A(_04807_),
    .B(_04808_));
 sg13g2_nor2_2 _11403_ (.A(net4532),
    .B(net4177),
    .Y(_04810_));
 sg13g2_nand2_1 _11404_ (.Y(_04811_),
    .A(_04303_),
    .B(_04810_));
 sg13g2_a21o_1 _11405_ (.A2(_00073_),
    .A1(net4560),
    .B1(_04282_),
    .X(_04812_));
 sg13g2_mux2_1 _11406_ (.A0(_04731_),
    .A1(_04812_),
    .S(net4194),
    .X(_04813_));
 sg13g2_nor2_1 _11407_ (.A(net3823),
    .B(_04813_),
    .Y(_04814_));
 sg13g2_nor3_1 _11408_ (.A(net4184),
    .B(net3824),
    .C(_04661_),
    .Y(_04815_));
 sg13g2_a21oi_1 _11409_ (.A1(net4184),
    .A2(_04814_),
    .Y(_04816_),
    .B1(_04815_));
 sg13g2_o21ai_1 _11410_ (.B1(_04811_),
    .Y(_04817_),
    .A1(net4527),
    .A2(_04816_));
 sg13g2_nand3_1 _11411_ (.B(net4090),
    .C(_04817_),
    .A(net4164),
    .Y(_04818_));
 sg13g2_mux4_1 _11412_ (.S0(net3905),
    .A0(_04112_),
    .A1(_04136_),
    .A2(_04195_),
    .A3(_04205_),
    .S1(net3788),
    .X(_04819_));
 sg13g2_and2_1 _11413_ (.A(net3782),
    .B(_04184_),
    .X(_04820_));
 sg13g2_mux2_1 _11414_ (.A0(_04819_),
    .A1(_04820_),
    .S(net3923),
    .X(_04821_));
 sg13g2_mux4_1 _11415_ (.S0(net3907),
    .A0(_04146_),
    .A1(_04157_),
    .A2(_04220_),
    .A3(_04230_),
    .S1(net3782),
    .X(_04822_));
 sg13g2_nand3_1 _11416_ (.B(_04289_),
    .C(_04291_),
    .A(net3784),
    .Y(_04823_));
 sg13g2_a21oi_1 _11417_ (.A1(net3790),
    .A2(_04252_),
    .Y(_04824_),
    .B1(net3925));
 sg13g2_a221oi_1 _11418_ (.B2(_04824_),
    .C1(net3833),
    .B1(_04823_),
    .A1(net3924),
    .Y(_04825_),
    .A2(_04822_));
 sg13g2_a21oi_1 _11419_ (.A1(net3836),
    .A2(_04821_),
    .Y(_04826_),
    .B1(_04825_));
 sg13g2_xnor2_1 _11420_ (.Y(_04827_),
    .A(_04818_),
    .B(_04826_));
 sg13g2_a21oi_1 _11421_ (.A1(_01062_),
    .A2(net4510),
    .Y(_04828_),
    .B1(net4014));
 sg13g2_a21oi_1 _11422_ (.A1(net4014),
    .A2(_04827_),
    .Y(_04829_),
    .B1(_04828_));
 sg13g2_or2_1 _11423_ (.X(_04830_),
    .B(_04829_),
    .A(\cpu.keccak_alu.registers[8] ));
 sg13g2_a21oi_1 _11424_ (.A1(\cpu.keccak_alu.registers[8] ),
    .A2(_04829_),
    .Y(_04831_),
    .B1(net4379));
 sg13g2_a22oi_1 _11425_ (.Y(_04832_),
    .B1(_04830_),
    .B2(_04831_),
    .A2(_04809_),
    .A1(net4379));
 sg13g2_or2_1 _11426_ (.X(_04833_),
    .B(_04832_),
    .A(net4315));
 sg13g2_o21ai_1 _11427_ (.B1(net3820),
    .Y(_04834_),
    .A1(net454),
    .A2(_04325_));
 sg13g2_a21oi_1 _11428_ (.A1(net4295),
    .A2(_04325_),
    .Y(_04835_),
    .B1(_04834_));
 sg13g2_nor2_1 _11429_ (.A(net3726),
    .B(_04835_),
    .Y(_04836_));
 sg13g2_a22oi_1 _11430_ (.Y(_00725_),
    .B1(_04833_),
    .B2(_04836_),
    .A2(net3726),
    .A1(_01066_));
 sg13g2_a21oi_1 _11431_ (.A1(net4509),
    .A2(\cpu.keccak_alu.registers[201] ),
    .Y(_04837_),
    .B1(net4366));
 sg13g2_o21ai_1 _11432_ (.B1(_04837_),
    .Y(_04838_),
    .A1(net4509),
    .A2(\cpu.keccak_alu.registers[201] ));
 sg13g2_xor2_1 _11433_ (.B(\cpu.keccak_alu.registers[73] ),
    .A(\cpu.keccak_alu.registers[9] ),
    .X(_04839_));
 sg13g2_xnor2_1 _11434_ (.Y(_04840_),
    .A(_04838_),
    .B(_04839_));
 sg13g2_a21oi_1 _11435_ (.A1(_04465_),
    .A2(_04488_),
    .Y(_04841_),
    .B1(net3826));
 sg13g2_nor2_1 _11436_ (.A(net4544),
    .B(_04841_),
    .Y(_04842_));
 sg13g2_a21oi_1 _11437_ (.A1(net4545),
    .A2(_04770_),
    .Y(_04843_),
    .B1(_04842_));
 sg13g2_mux2_1 _11438_ (.A0(_04702_),
    .A1(_04843_),
    .S(net4188),
    .X(_04844_));
 sg13g2_a22oi_1 _11439_ (.Y(_04845_),
    .B1(_04844_),
    .B2(net4177),
    .A2(_04810_),
    .A1(_04332_));
 sg13g2_nor2_1 _11440_ (.A(net4523),
    .B(_04845_),
    .Y(_04846_));
 sg13g2_nand2_1 _11441_ (.Y(_04847_),
    .A(net4089),
    .B(_04846_));
 sg13g2_mux4_1 _11442_ (.S0(net3911),
    .A0(_04426_),
    .A1(_04460_),
    .A2(_04515_),
    .A3(_04512_),
    .S1(net3792),
    .X(_04848_));
 sg13g2_nand2b_1 _11443_ (.Y(_04849_),
    .B(net3928),
    .A_N(_04848_));
 sg13g2_nand2b_1 _11444_ (.Y(_04850_),
    .B(net3791),
    .A_N(_04455_));
 sg13g2_a21oi_1 _11445_ (.A1(net3786),
    .A2(_04478_),
    .Y(_04851_),
    .B1(net3928));
 sg13g2_a21oi_1 _11446_ (.A1(_04850_),
    .A2(_04851_),
    .Y(_04852_),
    .B1(net3834));
 sg13g2_mux4_1 _11447_ (.S0(net3908),
    .A0(_04363_),
    .A1(_04372_),
    .A2(_04403_),
    .A3(_04413_),
    .S1(net3793),
    .X(_04853_));
 sg13g2_a221oi_1 _11448_ (.B2(_04383_),
    .C1(_04393_),
    .B1(net3903),
    .A1(_03879_),
    .Y(_04854_),
    .A2(_03880_));
 sg13g2_mux2_1 _11449_ (.A0(_04853_),
    .A1(_04854_),
    .S(net3926),
    .X(_04855_));
 sg13g2_a22oi_1 _11450_ (.Y(_04856_),
    .B1(_04855_),
    .B2(net3839),
    .A2(_04852_),
    .A1(_04849_));
 sg13g2_a21oi_1 _11451_ (.A1(_01072_),
    .A2(net4509),
    .Y(_04857_),
    .B1(net4009));
 sg13g2_xnor2_1 _11452_ (.Y(_04858_),
    .A(_04847_),
    .B(_04856_));
 sg13g2_a21oi_1 _11453_ (.A1(net4009),
    .A2(_04858_),
    .Y(_04859_),
    .B1(_04857_));
 sg13g2_or2_1 _11454_ (.X(_04860_),
    .B(_04859_),
    .A(\cpu.keccak_alu.registers[9] ));
 sg13g2_a21oi_1 _11455_ (.A1(\cpu.keccak_alu.registers[9] ),
    .A2(_04859_),
    .Y(_04861_),
    .B1(net4371));
 sg13g2_a22oi_1 _11456_ (.Y(_04862_),
    .B1(_04860_),
    .B2(_04861_),
    .A2(_04840_),
    .A1(net4371));
 sg13g2_or2_1 _11457_ (.X(_04863_),
    .B(_04862_),
    .A(net4313));
 sg13g2_o21ai_1 _11458_ (.B1(net3815),
    .Y(_04864_),
    .A1(net310),
    .A2(net3697));
 sg13g2_a21oi_1 _11459_ (.A1(net4290),
    .A2(net3697),
    .Y(_04865_),
    .B1(_04864_));
 sg13g2_nor2_1 _11460_ (.A(net3719),
    .B(_04865_),
    .Y(_04866_));
 sg13g2_a22oi_1 _11461_ (.Y(_00726_),
    .B1(_04863_),
    .B2(_04866_),
    .A2(net3719),
    .A1(_01074_));
 sg13g2_a21oi_1 _11462_ (.A1(\cpu.keccak_alu.registers[138] ),
    .A2(\cpu.keccak_alu.registers[202] ),
    .Y(_04867_),
    .B1(net4366));
 sg13g2_o21ai_1 _11463_ (.B1(_04867_),
    .Y(_04868_),
    .A1(\cpu.keccak_alu.registers[138] ),
    .A2(\cpu.keccak_alu.registers[202] ));
 sg13g2_xnor2_1 _11464_ (.Y(_04869_),
    .A(\cpu.keccak_alu.registers[10] ),
    .B(\cpu.keccak_alu.registers[74] ));
 sg13g2_o21ai_1 _11465_ (.B1(net4371),
    .Y(_04870_),
    .A1(_04868_),
    .A2(_04869_));
 sg13g2_a21oi_1 _11466_ (.A1(_04868_),
    .A2(_04869_),
    .Y(_04871_),
    .B1(_04870_));
 sg13g2_nand2b_1 _11467_ (.Y(_04872_),
    .B(_04810_),
    .A_N(_04533_));
 sg13g2_nand2_1 _11468_ (.Y(_04873_),
    .A(_04281_),
    .B(_04286_));
 sg13g2_mux2_1 _11469_ (.A0(_04812_),
    .A1(_04873_),
    .S(net4194),
    .X(_04874_));
 sg13g2_nor2_1 _11470_ (.A(net3824),
    .B(_04874_),
    .Y(_04875_));
 sg13g2_nor3_1 _11471_ (.A(net4534),
    .B(net3824),
    .C(_04874_),
    .Y(_04876_));
 sg13g2_a21oi_1 _11472_ (.A1(net4534),
    .A2(_04733_),
    .Y(_04877_),
    .B1(_04876_));
 sg13g2_o21ai_1 _11473_ (.B1(_04872_),
    .Y(_04878_),
    .A1(net4525),
    .A2(_04877_));
 sg13g2_nand2_1 _11474_ (.Y(_04879_),
    .A(net4164),
    .B(_04878_));
 sg13g2_nor2_1 _11475_ (.A(net3931),
    .B(_04879_),
    .Y(_04880_));
 sg13g2_mux4_1 _11476_ (.S0(net3905),
    .A0(_04538_),
    .A1(_04539_),
    .A2(_04545_),
    .A3(_04546_),
    .S1(net3788),
    .X(_04881_));
 sg13g2_a221oi_1 _11477_ (.B2(_04541_),
    .C1(_04544_),
    .B1(net3897),
    .A1(_03879_),
    .Y(_04882_),
    .A2(_03880_));
 sg13g2_mux2_1 _11478_ (.A0(_04881_),
    .A1(_04882_),
    .S(net3924),
    .X(_04883_));
 sg13g2_mux4_1 _11479_ (.S0(net3906),
    .A0(_04536_),
    .A1(_04537_),
    .A2(_04553_),
    .A3(_04554_),
    .S1(net3781),
    .X(_04884_));
 sg13g2_or2_1 _11480_ (.X(_04885_),
    .B(_04884_),
    .A(net3915));
 sg13g2_mux4_1 _11481_ (.S0(net3899),
    .A0(_04550_),
    .A1(_04551_),
    .A2(_04569_),
    .A3(_04566_),
    .S1(net3783),
    .X(_04886_));
 sg13g2_a21oi_1 _11482_ (.A1(net3913),
    .A2(_04886_),
    .Y(_04887_),
    .B1(net3833));
 sg13g2_a22oi_1 _11483_ (.Y(_04888_),
    .B1(_04885_),
    .B2(_04887_),
    .A2(_04883_),
    .A1(net3837));
 sg13g2_a21oi_1 _11484_ (.A1(_01078_),
    .A2(\cpu.keccak_alu.registers[138] ),
    .Y(_04889_),
    .B1(net4009));
 sg13g2_xor2_1 _11485_ (.B(_04888_),
    .A(_04880_),
    .X(_04890_));
 sg13g2_a21oi_1 _11486_ (.A1(net4009),
    .A2(_04890_),
    .Y(_04891_),
    .B1(_04889_));
 sg13g2_o21ai_1 _11487_ (.B1(net4213),
    .Y(_04892_),
    .A1(\cpu.keccak_alu.registers[10] ),
    .A2(_04891_));
 sg13g2_a21oi_1 _11488_ (.A1(\cpu.keccak_alu.registers[10] ),
    .A2(_04891_),
    .Y(_04893_),
    .B1(_04892_));
 sg13g2_o21ai_1 _11489_ (.B1(net4244),
    .Y(_04894_),
    .A1(_04871_),
    .A2(_04893_));
 sg13g2_o21ai_1 _11490_ (.B1(net3815),
    .Y(_04895_),
    .A1(net338),
    .A2(net3697));
 sg13g2_a21oi_1 _11491_ (.A1(net4286),
    .A2(net3697),
    .Y(_04896_),
    .B1(_04895_));
 sg13g2_nor2_1 _11492_ (.A(net3719),
    .B(_04896_),
    .Y(_04897_));
 sg13g2_a22oi_1 _11493_ (.Y(_00727_),
    .B1(_04894_),
    .B2(_04897_),
    .A2(net3719),
    .A1(_01081_));
 sg13g2_o21ai_1 _11494_ (.B1(_04464_),
    .Y(_04898_),
    .A1(net4568),
    .A2(_00077_));
 sg13g2_nand2_1 _11495_ (.Y(_04899_),
    .A(net3832),
    .B(_04898_));
 sg13g2_nand2_1 _11496_ (.Y(_04900_),
    .A(net4544),
    .B(_04841_));
 sg13g2_o21ai_1 _11497_ (.B1(_04900_),
    .Y(_04901_),
    .A1(net4544),
    .A2(_04899_));
 sg13g2_mux2_1 _11498_ (.A0(_04772_),
    .A1(_04901_),
    .S(net4188),
    .X(_04902_));
 sg13g2_inv_1 _11499_ (.Y(_04903_),
    .A(_04902_));
 sg13g2_nand2b_1 _11500_ (.Y(_04904_),
    .B(_04810_),
    .A_N(_04595_));
 sg13g2_o21ai_1 _11501_ (.B1(_04904_),
    .Y(_04905_),
    .A1(net4528),
    .A2(_04903_));
 sg13g2_nand3_1 _11502_ (.B(net4089),
    .C(_04905_),
    .A(net4168),
    .Y(_04906_));
 sg13g2_mux4_1 _11503_ (.S0(net3911),
    .A0(_04598_),
    .A1(_04599_),
    .A2(_04618_),
    .A3(_04619_),
    .S1(net3786),
    .X(_04907_));
 sg13g2_nor2_1 _11504_ (.A(net3921),
    .B(_04907_),
    .Y(_04908_));
 sg13g2_mux4_1 _11505_ (.S0(net3910),
    .A0(_04620_),
    .A1(_04621_),
    .A2(_04624_),
    .A3(_04625_),
    .S1(net3786),
    .X(_04909_));
 sg13g2_o21ai_1 _11506_ (.B1(net3777),
    .Y(_04910_),
    .A1(net3928),
    .A2(_04909_));
 sg13g2_or2_1 _11507_ (.X(_04911_),
    .B(_04910_),
    .A(_04908_));
 sg13g2_mux4_1 _11508_ (.S0(net3909),
    .A0(_04600_),
    .A1(_04601_),
    .A2(_04604_),
    .A3(_04605_),
    .S1(net3793),
    .X(_04912_));
 sg13g2_nand2b_1 _11509_ (.Y(_04913_),
    .B(net3920),
    .A_N(_04912_));
 sg13g2_a21o_1 _11510_ (.A2(_04609_),
    .A1(net3785),
    .B1(net3920),
    .X(_04914_));
 sg13g2_nand3_1 _11511_ (.B(_04913_),
    .C(_04914_),
    .A(net3840),
    .Y(_04915_));
 sg13g2_and3_1 _11512_ (.X(_04916_),
    .A(_04906_),
    .B(_04911_),
    .C(_04915_));
 sg13g2_a21oi_1 _11513_ (.A1(_04911_),
    .A2(_04915_),
    .Y(_04917_),
    .B1(_04906_));
 sg13g2_o21ai_1 _11514_ (.B1(net4000),
    .Y(_04918_),
    .A1(\cpu.keccak_alu.registers[75] ),
    .A2(_01088_));
 sg13g2_o21ai_1 _11515_ (.B1(net4019),
    .Y(_04919_),
    .A1(_04916_),
    .A2(_04917_));
 sg13g2_a21oi_1 _11516_ (.A1(_04918_),
    .A2(_04919_),
    .Y(_04920_),
    .B1(\cpu.keccak_alu.registers[11] ));
 sg13g2_and3_1 _11517_ (.X(_04921_),
    .A(\cpu.keccak_alu.registers[11] ),
    .B(_04918_),
    .C(_04919_));
 sg13g2_nor3_1 _11518_ (.A(net4374),
    .B(_04920_),
    .C(_04921_),
    .Y(_04922_));
 sg13g2_a21oi_1 _11519_ (.A1(\cpu.keccak_alu.registers[139] ),
    .A2(\cpu.keccak_alu.registers[203] ),
    .Y(_04923_),
    .B1(net4367));
 sg13g2_o21ai_1 _11520_ (.B1(_04923_),
    .Y(_04924_),
    .A1(\cpu.keccak_alu.registers[139] ),
    .A2(\cpu.keccak_alu.registers[203] ));
 sg13g2_xnor2_1 _11521_ (.Y(_04925_),
    .A(\cpu.keccak_alu.registers[11] ),
    .B(\cpu.keccak_alu.registers[75] ));
 sg13g2_o21ai_1 _11522_ (.B1(net4374),
    .Y(_04926_),
    .A1(_04924_),
    .A2(_04925_));
 sg13g2_a21oi_1 _11523_ (.A1(_04924_),
    .A2(_04925_),
    .Y(_04927_),
    .B1(_04926_));
 sg13g2_o21ai_1 _11524_ (.B1(net4244),
    .Y(_04928_),
    .A1(_04922_),
    .A2(_04927_));
 sg13g2_o21ai_1 _11525_ (.B1(net3817),
    .Y(_04929_),
    .A1(net283),
    .A2(net3697));
 sg13g2_a21oi_1 _11526_ (.A1(net4282),
    .A2(net3698),
    .Y(_04930_),
    .B1(_04929_));
 sg13g2_nor2_1 _11527_ (.A(net3723),
    .B(_04930_),
    .Y(_04931_));
 sg13g2_a22oi_1 _11528_ (.Y(_00728_),
    .B1(_04928_),
    .B2(_04931_),
    .A2(net3723),
    .A1(_01090_));
 sg13g2_nand3_1 _11529_ (.B(_04278_),
    .C(_04285_),
    .A(net4194),
    .Y(_04932_));
 sg13g2_nand3_1 _11530_ (.B(_04281_),
    .C(_04286_),
    .A(net4538),
    .Y(_04933_));
 sg13g2_a21oi_1 _11531_ (.A1(_04932_),
    .A2(_04933_),
    .Y(_04934_),
    .B1(net3823));
 sg13g2_mux2_1 _11532_ (.A0(_04814_),
    .A1(_04934_),
    .S(net4183),
    .X(_04935_));
 sg13g2_nor2_1 _11533_ (.A(net4525),
    .B(_04935_),
    .Y(_04936_));
 sg13g2_a21oi_1 _11534_ (.A1(net4525),
    .A2(_04663_),
    .Y(_04937_),
    .B1(_04936_));
 sg13g2_nand2_1 _11535_ (.Y(_04938_),
    .A(net4164),
    .B(_04937_));
 sg13g2_nor2_1 _11536_ (.A(net3931),
    .B(_04938_),
    .Y(_04939_));
 sg13g2_mux4_1 _11537_ (.S0(net3905),
    .A0(_04136_),
    .A1(_04195_),
    .A2(_04205_),
    .A3(_04171_),
    .S1(net3788),
    .X(_04940_));
 sg13g2_and3_1 _11538_ (.X(_04941_),
    .A(net3781),
    .B(net3901),
    .C(_04183_));
 sg13g2_nand3_1 _11539_ (.B(net3898),
    .C(_04183_),
    .A(net3782),
    .Y(_04942_));
 sg13g2_mux2_1 _11540_ (.A0(_04940_),
    .A1(_04941_),
    .S(net3923),
    .X(_04943_));
 sg13g2_o21ai_1 _11541_ (.B1(net3916),
    .Y(_04944_),
    .A1(net3783),
    .A2(_04676_));
 sg13g2_a21o_1 _11542_ (.A2(_04679_),
    .A1(net3783),
    .B1(_04944_),
    .X(_04945_));
 sg13g2_mux4_1 _11543_ (.S0(net3782),
    .A0(_04111_),
    .A1(_04146_),
    .A2(_04157_),
    .A3(_04230_),
    .S1(net3899),
    .X(_04946_));
 sg13g2_mux4_1 _11544_ (.S0(net3898),
    .A0(_04145_),
    .A1(_04256_),
    .A2(_04313_),
    .A3(_04310_),
    .S1(net3789),
    .X(_04947_));
 sg13g2_a21oi_1 _11545_ (.A1(net3924),
    .A2(_04946_),
    .Y(_04948_),
    .B1(net3833));
 sg13g2_a22oi_1 _11546_ (.Y(_04949_),
    .B1(_04945_),
    .B2(_04948_),
    .A2(_04943_),
    .A1(net3836));
 sg13g2_a21oi_1 _11547_ (.A1(_01095_),
    .A2(net4507),
    .Y(_04950_),
    .B1(net4014));
 sg13g2_xor2_1 _11548_ (.B(_04949_),
    .A(_04939_),
    .X(_04951_));
 sg13g2_a21oi_1 _11549_ (.A1(net4015),
    .A2(_04951_),
    .Y(_04952_),
    .B1(_04950_));
 sg13g2_a21oi_1 _11550_ (.A1(\cpu.keccak_alu.registers[12] ),
    .A2(_04952_),
    .Y(_04953_),
    .B1(net4377));
 sg13g2_o21ai_1 _11551_ (.B1(_04953_),
    .Y(_04954_),
    .A1(\cpu.keccak_alu.registers[12] ),
    .A2(_04952_));
 sg13g2_o21ai_1 _11552_ (.B1(net4208),
    .Y(_04955_),
    .A1(net4507),
    .A2(\cpu.keccak_alu.registers[204] ));
 sg13g2_a21oi_1 _11553_ (.A1(net4507),
    .A2(\cpu.keccak_alu.registers[204] ),
    .Y(_04956_),
    .B1(_04955_));
 sg13g2_xor2_1 _11554_ (.B(\cpu.keccak_alu.registers[76] ),
    .A(\cpu.keccak_alu.registers[12] ),
    .X(_04957_));
 sg13g2_a21oi_1 _11555_ (.A1(_04956_),
    .A2(_04957_),
    .Y(_04958_),
    .B1(net4216));
 sg13g2_o21ai_1 _11556_ (.B1(_04958_),
    .Y(_04959_),
    .A1(_04956_),
    .A2(_04957_));
 sg13g2_a21o_1 _11557_ (.A2(_04959_),
    .A1(_04954_),
    .B1(net4318),
    .X(_04960_));
 sg13g2_o21ai_1 _11558_ (.B1(net3818),
    .Y(_04961_),
    .A1(\cpu.keccak_alu.registers[268] ),
    .A2(_04325_));
 sg13g2_a21oi_1 _11559_ (.A1(net4278),
    .A2(net3698),
    .Y(_04962_),
    .B1(_04961_));
 sg13g2_nor2_1 _11560_ (.A(net3726),
    .B(_04962_),
    .Y(_04963_));
 sg13g2_a22oi_1 _11561_ (.Y(_00729_),
    .B1(_04960_),
    .B2(_04963_),
    .A2(net3727),
    .A1(_01099_));
 sg13g2_a21oi_1 _11562_ (.A1(net4506),
    .A2(\cpu.keccak_alu.registers[205] ),
    .Y(_04964_),
    .B1(net4366));
 sg13g2_o21ai_1 _11563_ (.B1(_04964_),
    .Y(_04965_),
    .A1(net4506),
    .A2(\cpu.keccak_alu.registers[205] ));
 sg13g2_xnor2_1 _11564_ (.Y(_04966_),
    .A(\cpu.keccak_alu.registers[13] ),
    .B(\cpu.keccak_alu.registers[77] ));
 sg13g2_o21ai_1 _11565_ (.B1(net4373),
    .Y(_04967_),
    .A1(_04965_),
    .A2(_04966_));
 sg13g2_a21oi_1 _11566_ (.A1(_04965_),
    .A2(_04966_),
    .Y(_04968_),
    .B1(_04967_));
 sg13g2_a21oi_1 _11567_ (.A1(_01103_),
    .A2(net4506),
    .Y(_04969_),
    .B1(net4012));
 sg13g2_mux2_1 _11568_ (.A0(_00079_),
    .A1(_00078_),
    .S(net4573),
    .X(_04970_));
 sg13g2_nor2_1 _11569_ (.A(net3826),
    .B(_04970_),
    .Y(_04971_));
 sg13g2_nor2_1 _11570_ (.A(net4544),
    .B(_04971_),
    .Y(_04972_));
 sg13g2_a21oi_1 _11571_ (.A1(net4544),
    .A2(_04899_),
    .Y(_04973_),
    .B1(_04972_));
 sg13g2_mux2_1 _11572_ (.A0(_04843_),
    .A1(_04973_),
    .S(net4188),
    .X(_04974_));
 sg13g2_nand2_1 _11573_ (.Y(_04975_),
    .A(net4177),
    .B(_04974_));
 sg13g2_o21ai_1 _11574_ (.B1(_04975_),
    .Y(_04976_),
    .A1(net4175),
    .A2(_04703_));
 sg13g2_nand2_1 _11575_ (.Y(_04977_),
    .A(net4168),
    .B(_04976_));
 sg13g2_nor2_1 _11576_ (.A(net3933),
    .B(_04977_),
    .Y(_04978_));
 sg13g2_mux4_1 _11577_ (.S0(net3902),
    .A0(_04363_),
    .A1(_04512_),
    .A2(_04515_),
    .A3(_04460_),
    .S1(net3786),
    .X(_04979_));
 sg13g2_nand2b_1 _11578_ (.Y(_04980_),
    .B(net3926),
    .A_N(_04979_));
 sg13g2_nand2_1 _11579_ (.Y(_04981_),
    .A(net3791),
    .B(_04711_));
 sg13g2_a21oi_1 _11580_ (.A1(net3786),
    .A2(_04707_),
    .Y(_04982_),
    .B1(net3929));
 sg13g2_a21oi_2 _11581_ (.B1(net3834),
    .Y(_04983_),
    .A2(_04982_),
    .A1(_04981_));
 sg13g2_mux4_1 _11582_ (.S0(net3909),
    .A0(_04372_),
    .A1(_04403_),
    .A2(_04413_),
    .A3(_04384_),
    .S1(net3793),
    .X(_04984_));
 sg13g2_nor3_1 _11583_ (.A(net3793),
    .B(net3909),
    .C(_04392_),
    .Y(_04985_));
 sg13g2_mux2_1 _11584_ (.A0(_04984_),
    .A1(_04985_),
    .S(net3926),
    .X(_04986_));
 sg13g2_a22oi_1 _11585_ (.Y(_04987_),
    .B1(_04986_),
    .B2(net3839),
    .A2(_04983_),
    .A1(_04980_));
 sg13g2_xor2_1 _11586_ (.B(_04987_),
    .A(_04978_),
    .X(_04988_));
 sg13g2_a21oi_1 _11587_ (.A1(net4012),
    .A2(_04988_),
    .Y(_04989_),
    .B1(_04969_));
 sg13g2_o21ai_1 _11588_ (.B1(net4213),
    .Y(_04990_),
    .A1(\cpu.keccak_alu.registers[13] ),
    .A2(_04989_));
 sg13g2_a21oi_1 _11589_ (.A1(net953),
    .A2(_04989_),
    .Y(_04991_),
    .B1(_04990_));
 sg13g2_o21ai_1 _11590_ (.B1(net4244),
    .Y(_04992_),
    .A1(_04968_),
    .A2(_04991_));
 sg13g2_o21ai_1 _11591_ (.B1(net3816),
    .Y(_04993_),
    .A1(net386),
    .A2(net3698));
 sg13g2_a21oi_1 _11592_ (.A1(net4275),
    .A2(net3697),
    .Y(_04994_),
    .B1(_04993_));
 sg13g2_nor2_1 _11593_ (.A(net3725),
    .B(_04994_),
    .Y(_04995_));
 sg13g2_a22oi_1 _11594_ (.Y(_00730_),
    .B1(_04992_),
    .B2(_04995_),
    .A2(net3722),
    .A1(_01107_));
 sg13g2_a21oi_1 _11595_ (.A1(net4505),
    .A2(\cpu.keccak_alu.registers[206] ),
    .Y(_04996_),
    .B1(net4366));
 sg13g2_o21ai_1 _11596_ (.B1(_04996_),
    .Y(_04997_),
    .A1(net4505),
    .A2(\cpu.keccak_alu.registers[206] ));
 sg13g2_xor2_1 _11597_ (.B(\cpu.keccak_alu.registers[78] ),
    .A(\cpu.keccak_alu.registers[14] ),
    .X(_04998_));
 sg13g2_xnor2_1 _11598_ (.Y(_04999_),
    .A(_04997_),
    .B(_04998_));
 sg13g2_nand3_1 _11599_ (.B(_04274_),
    .C(_04277_),
    .A(net4194),
    .Y(_05000_));
 sg13g2_nand3_1 _11600_ (.B(_04278_),
    .C(_04285_),
    .A(net4539),
    .Y(_05001_));
 sg13g2_a21oi_1 _11601_ (.A1(_05000_),
    .A2(_05001_),
    .Y(_05002_),
    .B1(net3823));
 sg13g2_mux2_1 _11602_ (.A0(_04875_),
    .A1(_05002_),
    .S(net4182),
    .X(_05003_));
 sg13g2_nor2_1 _11603_ (.A(net4526),
    .B(_05003_),
    .Y(_05004_));
 sg13g2_a21oi_1 _11604_ (.A1(net4526),
    .A2(_04735_),
    .Y(_05005_),
    .B1(_05004_));
 sg13g2_and2_1 _11605_ (.A(net4165),
    .B(_05005_),
    .X(_05006_));
 sg13g2_nand2_1 _11606_ (.Y(_05007_),
    .A(net4090),
    .B(_05006_));
 sg13g2_mux4_1 _11607_ (.S0(net3905),
    .A0(_04539_),
    .A1(_04545_),
    .A2(_04546_),
    .A3(_04542_),
    .S1(net3788),
    .X(_05008_));
 sg13g2_and3_1 _11608_ (.X(_05009_),
    .A(net3781),
    .B(net3897),
    .C(_04543_));
 sg13g2_mux2_1 _11609_ (.A0(_05008_),
    .A1(_05009_),
    .S(net3923),
    .X(_05010_));
 sg13g2_mux4_1 _11610_ (.S0(net3788),
    .A0(_04536_),
    .A1(_04538_),
    .A2(_04554_),
    .A3(_04537_),
    .S1(net3898),
    .X(_05011_));
 sg13g2_or2_1 _11611_ (.X(_05012_),
    .B(_05011_),
    .A(net3913));
 sg13g2_nand2_1 _11612_ (.Y(_05013_),
    .A(net3783),
    .B(_04742_));
 sg13g2_a21oi_1 _11613_ (.A1(net3790),
    .A2(_04739_),
    .Y(_05014_),
    .B1(net3924));
 sg13g2_a21oi_1 _11614_ (.A1(_05013_),
    .A2(_05014_),
    .Y(_05015_),
    .B1(net3833));
 sg13g2_a22oi_1 _11615_ (.Y(_05016_),
    .B1(_05012_),
    .B2(_05015_),
    .A2(_05010_),
    .A1(net3836));
 sg13g2_a21oi_1 _11616_ (.A1(_01118_),
    .A2(net4505),
    .Y(_05017_),
    .B1(net4009));
 sg13g2_xnor2_1 _11617_ (.Y(_05018_),
    .A(_05007_),
    .B(_05016_));
 sg13g2_a21oi_1 _11618_ (.A1(net4009),
    .A2(_05018_),
    .Y(_05019_),
    .B1(_05017_));
 sg13g2_or2_1 _11619_ (.X(_05020_),
    .B(_05019_),
    .A(\cpu.keccak_alu.registers[14] ));
 sg13g2_a21oi_1 _11620_ (.A1(\cpu.keccak_alu.registers[14] ),
    .A2(_05019_),
    .Y(_05021_),
    .B1(net4371));
 sg13g2_a22oi_1 _11621_ (.Y(_05022_),
    .B1(_05020_),
    .B2(_05021_),
    .A2(_04999_),
    .A1(net4371));
 sg13g2_or2_1 _11622_ (.X(_05023_),
    .B(_05022_),
    .A(net4313));
 sg13g2_o21ai_1 _11623_ (.B1(net3815),
    .Y(_05024_),
    .A1(net277),
    .A2(net3697));
 sg13g2_a21oi_1 _11624_ (.A1(net4273),
    .A2(net3697),
    .Y(_05025_),
    .B1(_05024_));
 sg13g2_nor2_1 _11625_ (.A(net3719),
    .B(_05025_),
    .Y(_05026_));
 sg13g2_a22oi_1 _11626_ (.Y(_00731_),
    .B1(_05023_),
    .B2(_05026_),
    .A2(net3719),
    .A1(_01122_));
 sg13g2_o21ai_1 _11627_ (.B1(_04471_),
    .Y(_05027_),
    .A1(net4567),
    .A2(_00081_));
 sg13g2_nand2_1 _11628_ (.Y(_05028_),
    .A(net3832),
    .B(_05027_));
 sg13g2_nand2_1 _11629_ (.Y(_05029_),
    .A(net4544),
    .B(_04971_));
 sg13g2_o21ai_1 _11630_ (.B1(_05029_),
    .Y(_05030_),
    .A1(net4543),
    .A2(_05028_));
 sg13g2_mux2_1 _11631_ (.A0(_04901_),
    .A1(_05030_),
    .S(net4188),
    .X(_05031_));
 sg13g2_nand2_1 _11632_ (.Y(_05032_),
    .A(net4178),
    .B(_05031_));
 sg13g2_o21ai_1 _11633_ (.B1(_05032_),
    .Y(_05033_),
    .A1(net4178),
    .A2(_04775_));
 sg13g2_nand3_1 _11634_ (.B(net4090),
    .C(_05033_),
    .A(net4170),
    .Y(_05034_));
 sg13g2_nand2_1 _11635_ (.Y(_05035_),
    .A(net3791),
    .B(_04783_));
 sg13g2_a21oi_1 _11636_ (.A1(net3787),
    .A2(_04780_),
    .Y(_05036_),
    .B1(net3929));
 sg13g2_mux4_1 _11637_ (.S0(net3792),
    .A0(_04598_),
    .A1(_04600_),
    .A2(_04619_),
    .A3(_04599_),
    .S1(net3902),
    .X(_05037_));
 sg13g2_or2_1 _11638_ (.X(_05038_),
    .B(_05037_),
    .A(net3921));
 sg13g2_nor4_1 _11639_ (.A(net4576),
    .B(net3918),
    .C(_03880_),
    .D(net3541),
    .Y(_05039_));
 sg13g2_mux2_1 _11640_ (.A0(_04786_),
    .A1(_04789_),
    .S(net3793),
    .X(_05040_));
 sg13g2_a21o_1 _11641_ (.A2(_05040_),
    .A1(net3918),
    .B1(_05039_),
    .X(_05041_));
 sg13g2_a21oi_1 _11642_ (.A1(_05035_),
    .A2(_05036_),
    .Y(_05042_),
    .B1(net3834));
 sg13g2_a22oi_1 _11643_ (.Y(_05043_),
    .B1(_05042_),
    .B2(_05038_),
    .A2(_05041_),
    .A1(net3839));
 sg13g2_a21oi_1 _11644_ (.A1(_01133_),
    .A2(\cpu.keccak_alu.registers[143] ),
    .Y(_05044_),
    .B1(net4013));
 sg13g2_xnor2_1 _11645_ (.Y(_05045_),
    .A(_05034_),
    .B(_05043_));
 sg13g2_a21oi_1 _11646_ (.A1(net4021),
    .A2(_05045_),
    .Y(_05046_),
    .B1(_05044_));
 sg13g2_or2_1 _11647_ (.X(_05047_),
    .B(_05046_),
    .A(\cpu.keccak_alu.registers[15] ));
 sg13g2_a21oi_1 _11648_ (.A1(\cpu.keccak_alu.registers[15] ),
    .A2(_05046_),
    .Y(_05048_),
    .B1(net4380));
 sg13g2_a21oi_1 _11649_ (.A1(net4504),
    .A2(\cpu.keccak_alu.registers[207] ),
    .Y(_05049_),
    .B1(net4368));
 sg13g2_o21ai_1 _11650_ (.B1(_05049_),
    .Y(_05050_),
    .A1(net4504),
    .A2(\cpu.keccak_alu.registers[207] ));
 sg13g2_xor2_1 _11651_ (.B(\cpu.keccak_alu.registers[79] ),
    .A(\cpu.keccak_alu.registers[15] ),
    .X(_05051_));
 sg13g2_xnor2_1 _11652_ (.Y(_05052_),
    .A(_05050_),
    .B(_05051_));
 sg13g2_a22oi_1 _11653_ (.Y(_05053_),
    .B1(_05052_),
    .B2(net4376),
    .A2(_05048_),
    .A1(_05047_));
 sg13g2_or2_1 _11654_ (.X(_05054_),
    .B(_05053_),
    .A(net4315));
 sg13g2_a22oi_1 _11655_ (.Y(_05055_),
    .B1(_04326_),
    .B2(net606),
    .A2(net3754),
    .A1(_02480_));
 sg13g2_nor2_1 _11656_ (.A(net3811),
    .B(_05055_),
    .Y(_05056_));
 sg13g2_nor2_1 _11657_ (.A(net3729),
    .B(_05056_),
    .Y(_05057_));
 sg13g2_a22oi_1 _11658_ (.Y(_00732_),
    .B1(_05054_),
    .B2(_05057_),
    .A2(net3726),
    .A1(_01135_));
 sg13g2_and2_1 _11659_ (.A(net3917),
    .B(_04206_),
    .X(_05058_));
 sg13g2_nor2b_1 _11660_ (.A(_04240_),
    .B_N(_04273_),
    .Y(_05059_));
 sg13g2_nand2_1 _11661_ (.Y(_05060_),
    .A(net4194),
    .B(_05059_));
 sg13g2_nand3_1 _11662_ (.B(_04274_),
    .C(_04277_),
    .A(net4538),
    .Y(_05061_));
 sg13g2_a21oi_1 _11663_ (.A1(_05060_),
    .A2(_05061_),
    .Y(_05062_),
    .B1(net3823));
 sg13g2_mux2_1 _11664_ (.A0(_04934_),
    .A1(_05062_),
    .S(net4183),
    .X(_05063_));
 sg13g2_nor2_1 _11665_ (.A(net4525),
    .B(_05063_),
    .Y(_05064_));
 sg13g2_a21oi_1 _11666_ (.A1(net4527),
    .A2(_04816_),
    .Y(_05065_),
    .B1(_05064_));
 sg13g2_nor2_1 _11667_ (.A(net4167),
    .B(_04304_),
    .Y(_05066_));
 sg13g2_a21oi_1 _11668_ (.A1(net4167),
    .A2(_05065_),
    .Y(_05067_),
    .B1(_05066_));
 sg13g2_nor2_1 _11669_ (.A(net3932),
    .B(_05067_),
    .Y(_05068_));
 sg13g2_mux2_1 _11670_ (.A0(_04159_),
    .A1(_04257_),
    .S(net3916),
    .X(_05069_));
 sg13g2_a221oi_1 _11671_ (.B2(net3775),
    .C1(_05068_),
    .B1(_05069_),
    .A1(net3838),
    .Y(_05070_),
    .A2(_05058_));
 sg13g2_nand3b_1 _11672_ (.B(\cpu.keccak_alu.registers[144] ),
    .C(net4005),
    .Y(_05071_),
    .A_N(\cpu.keccak_alu.registers[80] ));
 sg13g2_o21ai_1 _11673_ (.B1(_05071_),
    .Y(_05072_),
    .A1(net4005),
    .A2(_05070_));
 sg13g2_a21oi_1 _11674_ (.A1(\cpu.keccak_alu.registers[16] ),
    .A2(_05072_),
    .Y(_05073_),
    .B1(net4386));
 sg13g2_o21ai_1 _11675_ (.B1(_05073_),
    .Y(_05074_),
    .A1(\cpu.keccak_alu.registers[16] ),
    .A2(_05072_));
 sg13g2_o21ai_1 _11676_ (.B1(net4210),
    .Y(_05075_),
    .A1(net4503),
    .A2(\cpu.keccak_alu.registers[208] ));
 sg13g2_a21oi_1 _11677_ (.A1(net4503),
    .A2(\cpu.keccak_alu.registers[208] ),
    .Y(_05076_),
    .B1(_05075_));
 sg13g2_xor2_1 _11678_ (.B(\cpu.keccak_alu.registers[80] ),
    .A(\cpu.keccak_alu.registers[16] ),
    .X(_05077_));
 sg13g2_a21oi_1 _11679_ (.A1(_05076_),
    .A2(_05077_),
    .Y(_05078_),
    .B1(net4219));
 sg13g2_o21ai_1 _11680_ (.B1(_05078_),
    .Y(_05079_),
    .A1(_05076_),
    .A2(_05077_));
 sg13g2_a21oi_1 _11681_ (.A1(_05074_),
    .A2(_05079_),
    .Y(_05080_),
    .B1(net4321));
 sg13g2_a21oi_2 _11682_ (.B1(_02286_),
    .Y(_05081_),
    .A2(_02258_),
    .A1(net4432));
 sg13g2_and2_2 _11683_ (.A(_02289_),
    .B(net3770),
    .X(_05082_));
 sg13g2_nand2_2 _11684_ (.Y(_05083_),
    .A(_02289_),
    .B(net3771));
 sg13g2_nor2_2 _11685_ (.A(_02285_),
    .B(_05083_),
    .Y(_05084_));
 sg13g2_nand2_1 _11686_ (.Y(_05085_),
    .A(_02284_),
    .B(_05082_));
 sg13g2_o21ai_1 _11687_ (.B1(net3820),
    .Y(_05086_),
    .A1(net254),
    .A2(_05084_));
 sg13g2_a21oi_1 _11688_ (.A1(net4364),
    .A2(_05084_),
    .Y(_05087_),
    .B1(_05086_));
 sg13g2_nor3_1 _11689_ (.A(net3733),
    .B(_05080_),
    .C(_05087_),
    .Y(_05088_));
 sg13g2_a21oi_1 _11690_ (.A1(_00998_),
    .A2(net3733),
    .Y(_00733_),
    .B1(_05088_));
 sg13g2_o21ai_1 _11691_ (.B1(net4209),
    .Y(_05089_),
    .A1(\cpu.keccak_alu.registers[145] ),
    .A2(\cpu.keccak_alu.registers[209] ));
 sg13g2_a21oi_1 _11692_ (.A1(\cpu.keccak_alu.registers[145] ),
    .A2(\cpu.keccak_alu.registers[209] ),
    .Y(_05090_),
    .B1(_05089_));
 sg13g2_xor2_1 _11693_ (.B(\cpu.keccak_alu.registers[81] ),
    .A(\cpu.keccak_alu.registers[17] ),
    .X(_05091_));
 sg13g2_a21oi_1 _11694_ (.A1(_05090_),
    .A2(_05091_),
    .Y(_05092_),
    .B1(net4218));
 sg13g2_o21ai_1 _11695_ (.B1(_05092_),
    .Y(_05093_),
    .A1(_05090_),
    .A2(_05091_));
 sg13g2_nand2b_1 _11696_ (.Y(_05094_),
    .B(_04468_),
    .A_N(_04437_));
 sg13g2_nand3_1 _11697_ (.B(net3832),
    .C(_05094_),
    .A(net4200),
    .Y(_05095_));
 sg13g2_o21ai_1 _11698_ (.B1(_05095_),
    .Y(_05096_),
    .A1(net4200),
    .A2(_05028_));
 sg13g2_mux2_1 _11699_ (.A0(_04973_),
    .A1(_05096_),
    .S(net4188),
    .X(_05097_));
 sg13g2_mux2_1 _11700_ (.A0(_04844_),
    .A1(_05097_),
    .S(net4177),
    .X(_05098_));
 sg13g2_nor2_1 _11701_ (.A(net4169),
    .B(_04333_),
    .Y(_05099_));
 sg13g2_a21oi_1 _11702_ (.A1(net4169),
    .A2(_05098_),
    .Y(_05100_),
    .B1(_05099_));
 sg13g2_nor2_1 _11703_ (.A(net3933),
    .B(_05100_),
    .Y(_05101_));
 sg13g2_nor2_1 _11704_ (.A(net3921),
    .B(_04374_),
    .Y(_05102_));
 sg13g2_o21ai_1 _11705_ (.B1(net4006),
    .Y(_05103_),
    .A1(\cpu.keccak_alu.registers[81] ),
    .A2(_01004_));
 sg13g2_a21o_1 _11706_ (.A2(_04462_),
    .A1(net3921),
    .B1(net3834),
    .X(_05104_));
 sg13g2_nand3_1 _11707_ (.B(net3921),
    .C(_04507_),
    .A(net3839),
    .Y(_05105_));
 sg13g2_o21ai_1 _11708_ (.B1(_05105_),
    .Y(_05106_),
    .A1(_05102_),
    .A2(_05104_));
 sg13g2_xor2_1 _11709_ (.B(_05106_),
    .A(_05101_),
    .X(_05107_));
 sg13g2_o21ai_1 _11710_ (.B1(_05103_),
    .Y(_05108_),
    .A1(net4006),
    .A2(_05107_));
 sg13g2_xor2_1 _11711_ (.B(_05108_),
    .A(\cpu.keccak_alu.registers[17] ),
    .X(_05109_));
 sg13g2_o21ai_1 _11712_ (.B1(_05093_),
    .Y(_05110_),
    .A1(net4384),
    .A2(_05109_));
 sg13g2_a22oi_1 _11713_ (.Y(_05111_),
    .B1(net3696),
    .B2(net94),
    .A2(_05082_),
    .A1(_02294_));
 sg13g2_o21ai_1 _11714_ (.B1(net3739),
    .Y(_05112_),
    .A1(net3813),
    .A2(_05111_));
 sg13g2_a21oi_1 _11715_ (.A1(net4264),
    .A2(_05110_),
    .Y(_05113_),
    .B1(_05112_));
 sg13g2_a21oi_1 _11716_ (.A1(_01006_),
    .A2(net3735),
    .Y(_00734_),
    .B1(_05113_));
 sg13g2_o21ai_1 _11717_ (.B1(net4209),
    .Y(_05114_),
    .A1(\cpu.keccak_alu.registers[146] ),
    .A2(\cpu.keccak_alu.registers[210] ));
 sg13g2_a21oi_1 _11718_ (.A1(\cpu.keccak_alu.registers[146] ),
    .A2(\cpu.keccak_alu.registers[210] ),
    .Y(_05115_),
    .B1(_05114_));
 sg13g2_xor2_1 _11719_ (.B(\cpu.keccak_alu.registers[82] ),
    .A(\cpu.keccak_alu.registers[18] ),
    .X(_05116_));
 sg13g2_o21ai_1 _11720_ (.B1(net4384),
    .Y(_05117_),
    .A1(_05115_),
    .A2(_05116_));
 sg13g2_a21oi_1 _11721_ (.A1(_05115_),
    .A2(_05116_),
    .Y(_05118_),
    .B1(_05117_));
 sg13g2_nor3_1 _11722_ (.A(net4539),
    .B(_04241_),
    .C(_04242_),
    .Y(_05119_));
 sg13g2_a21oi_1 _11723_ (.A1(net4539),
    .A2(_05059_),
    .Y(_05120_),
    .B1(_05119_));
 sg13g2_nor2_1 _11724_ (.A(net3823),
    .B(_05120_),
    .Y(_05121_));
 sg13g2_mux2_1 _11725_ (.A0(_05002_),
    .A1(_05121_),
    .S(net4183),
    .X(_05122_));
 sg13g2_nand2_1 _11726_ (.Y(_05123_),
    .A(net4172),
    .B(_05122_));
 sg13g2_o21ai_1 _11727_ (.B1(_05123_),
    .Y(_05124_),
    .A1(net4172),
    .A2(_04877_));
 sg13g2_nor2_1 _11728_ (.A(net4521),
    .B(_05124_),
    .Y(_05125_));
 sg13g2_a21oi_1 _11729_ (.A1(net4521),
    .A2(_04534_),
    .Y(_05126_),
    .B1(_05125_));
 sg13g2_nand2_1 _11730_ (.Y(_05127_),
    .A(net4090),
    .B(_05126_));
 sg13g2_and2_1 _11731_ (.A(net3916),
    .B(_04556_),
    .X(_05128_));
 sg13g2_o21ai_1 _11732_ (.B1(net3774),
    .Y(_05129_),
    .A1(net3916),
    .A2(_04540_));
 sg13g2_nand3_1 _11733_ (.B(net3916),
    .C(_04577_),
    .A(net3838),
    .Y(_05130_));
 sg13g2_o21ai_1 _11734_ (.B1(_05130_),
    .Y(_05131_),
    .A1(_05128_),
    .A2(_05129_));
 sg13g2_o21ai_1 _11735_ (.B1(net4006),
    .Y(_05132_),
    .A1(\cpu.keccak_alu.registers[82] ),
    .A2(_01012_));
 sg13g2_xnor2_1 _11736_ (.Y(_05133_),
    .A(_05127_),
    .B(_05131_));
 sg13g2_o21ai_1 _11737_ (.B1(_05132_),
    .Y(_05134_),
    .A1(net4006),
    .A2(_05133_));
 sg13g2_o21ai_1 _11738_ (.B1(net4218),
    .Y(_05135_),
    .A1(_01009_),
    .A2(_05134_));
 sg13g2_a21oi_1 _11739_ (.A1(_01009_),
    .A2(_05134_),
    .Y(_05136_),
    .B1(_05135_));
 sg13g2_o21ai_1 _11740_ (.B1(net4264),
    .Y(_05137_),
    .A1(_05118_),
    .A2(_05136_));
 sg13g2_nand2_1 _11741_ (.Y(_05138_),
    .A(_01014_),
    .B(net3696));
 sg13g2_a21oi_1 _11742_ (.A1(net4355),
    .A2(_05084_),
    .Y(_05139_),
    .B1(_04324_));
 sg13g2_a21oi_1 _11743_ (.A1(_05138_),
    .A2(_05139_),
    .Y(_05140_),
    .B1(net3733));
 sg13g2_a22oi_1 _11744_ (.Y(_00735_),
    .B1(_05137_),
    .B2(_05140_),
    .A2(net3734),
    .A1(_01014_));
 sg13g2_o21ai_1 _11745_ (.B1(net4209),
    .Y(_05141_),
    .A1(\cpu.keccak_alu.registers[147] ),
    .A2(\cpu.keccak_alu.registers[211] ));
 sg13g2_a21oi_1 _11746_ (.A1(\cpu.keccak_alu.registers[147] ),
    .A2(\cpu.keccak_alu.registers[211] ),
    .Y(_05142_),
    .B1(_05141_));
 sg13g2_xor2_1 _11747_ (.B(\cpu.keccak_alu.registers[83] ),
    .A(\cpu.keccak_alu.registers[19] ),
    .X(_05143_));
 sg13g2_a21oi_1 _11748_ (.A1(_05142_),
    .A2(_05143_),
    .Y(_05144_),
    .B1(net4218));
 sg13g2_o21ai_1 _11749_ (.B1(_05144_),
    .Y(_05145_),
    .A1(_05142_),
    .A2(_05143_));
 sg13g2_a21oi_1 _11750_ (.A1(_04434_),
    .A2(_04438_),
    .Y(_05146_),
    .B1(net3826));
 sg13g2_a21oi_1 _11751_ (.A1(net3832),
    .A2(_05094_),
    .Y(_05147_),
    .B1(net4200));
 sg13g2_nor2_1 _11752_ (.A(net4544),
    .B(_05146_),
    .Y(_05148_));
 sg13g2_nor2_1 _11753_ (.A(_05147_),
    .B(_05148_),
    .Y(_05149_));
 sg13g2_mux2_1 _11754_ (.A0(_05030_),
    .A1(_05149_),
    .S(net4188),
    .X(_05150_));
 sg13g2_nand2_1 _11755_ (.Y(_05151_),
    .A(net4177),
    .B(_05150_));
 sg13g2_o21ai_1 _11756_ (.B1(_05151_),
    .Y(_05152_),
    .A1(net4177),
    .A2(_04903_));
 sg13g2_nor2_1 _11757_ (.A(net4169),
    .B(_04596_),
    .Y(_05153_));
 sg13g2_a21oi_1 _11758_ (.A1(net4169),
    .A2(_05152_),
    .Y(_05154_),
    .B1(_05153_));
 sg13g2_nor2_1 _11759_ (.A(net3933),
    .B(_05154_),
    .Y(_05155_));
 sg13g2_nor3_1 _11760_ (.A(net3928),
    .B(_04611_),
    .C(_04615_),
    .Y(_05156_));
 sg13g2_mux2_1 _11761_ (.A0(_04602_),
    .A1(_04622_),
    .S(net3922),
    .X(_05157_));
 sg13g2_a22oi_1 _11762_ (.Y(_05158_),
    .B1(_05157_),
    .B2(net3778),
    .A2(_05156_),
    .A1(net3839));
 sg13g2_a21oi_1 _11763_ (.A1(_01018_),
    .A2(\cpu.keccak_alu.registers[147] ),
    .Y(_05159_),
    .B1(net4020));
 sg13g2_xor2_1 _11764_ (.B(_05158_),
    .A(_05155_),
    .X(_05160_));
 sg13g2_a21oi_1 _11765_ (.A1(net4019),
    .A2(_05160_),
    .Y(_05161_),
    .B1(_05159_));
 sg13g2_xnor2_1 _11766_ (.Y(_05162_),
    .A(\cpu.keccak_alu.registers[19] ),
    .B(_05161_));
 sg13g2_o21ai_1 _11767_ (.B1(_05145_),
    .Y(_05163_),
    .A1(net4384),
    .A2(_05162_));
 sg13g2_a22oi_1 _11768_ (.Y(_05164_),
    .B1(net3696),
    .B2(net116),
    .A2(_05082_),
    .A1(_02297_));
 sg13g2_o21ai_1 _11769_ (.B1(net3739),
    .Y(_05165_),
    .A1(net3813),
    .A2(_05164_));
 sg13g2_a21oi_1 _11770_ (.A1(net4264),
    .A2(_05163_),
    .Y(_05166_),
    .B1(_05165_));
 sg13g2_a21oi_1 _11771_ (.A1(_01023_),
    .A2(net3734),
    .Y(_00736_),
    .B1(_05166_));
 sg13g2_o21ai_1 _11772_ (.B1(net4211),
    .Y(_05167_),
    .A1(\cpu.keccak_alu.registers[148] ),
    .A2(\cpu.keccak_alu.registers[212] ));
 sg13g2_a21oi_1 _11773_ (.A1(\cpu.keccak_alu.registers[148] ),
    .A2(\cpu.keccak_alu.registers[212] ),
    .Y(_05168_),
    .B1(_05167_));
 sg13g2_xor2_1 _11774_ (.B(\cpu.keccak_alu.registers[84] ),
    .A(\cpu.keccak_alu.registers[20] ),
    .X(_05169_));
 sg13g2_a21oi_1 _11775_ (.A1(_05168_),
    .A2(_05169_),
    .Y(_05170_),
    .B1(net4220));
 sg13g2_o21ai_1 _11776_ (.B1(_05170_),
    .Y(_05171_),
    .A1(_05168_),
    .A2(_05169_));
 sg13g2_nor3_1 _11777_ (.A(net4539),
    .B(_04231_),
    .C(_04243_),
    .Y(_05172_));
 sg13g2_nor3_1 _11778_ (.A(net4194),
    .B(_04241_),
    .C(_04242_),
    .Y(_05173_));
 sg13g2_nor2_1 _11779_ (.A(_05172_),
    .B(_05173_),
    .Y(_05174_));
 sg13g2_nor2_1 _11780_ (.A(net3823),
    .B(_05174_),
    .Y(_05175_));
 sg13g2_mux2_1 _11781_ (.A0(_05062_),
    .A1(_05175_),
    .S(net4182),
    .X(_05176_));
 sg13g2_mux2_1 _11782_ (.A0(_04935_),
    .A1(_05176_),
    .S(net4171),
    .X(_05177_));
 sg13g2_nor3_1 _11783_ (.A(net4525),
    .B(net4167),
    .C(_04663_),
    .Y(_05178_));
 sg13g2_a21oi_1 _11784_ (.A1(net4167),
    .A2(_05177_),
    .Y(_05179_),
    .B1(_05178_));
 sg13g2_nor2_1 _11785_ (.A(net3932),
    .B(_05179_),
    .Y(_05180_));
 sg13g2_nand4_1 _11786_ (.B(net3914),
    .C(_04668_),
    .A(net3837),
    .Y(_05181_),
    .D(_04670_));
 sg13g2_nor2_1 _11787_ (.A(net3914),
    .B(_04673_),
    .Y(_05182_));
 sg13g2_o21ai_1 _11788_ (.B1(net3774),
    .Y(_05183_),
    .A1(net3924),
    .A2(_04677_));
 sg13g2_o21ai_1 _11789_ (.B1(_05181_),
    .Y(_05184_),
    .A1(_05182_),
    .A2(_05183_));
 sg13g2_a21oi_1 _11790_ (.A1(_01027_),
    .A2(\cpu.keccak_alu.registers[148] ),
    .Y(_05185_),
    .B1(net4016));
 sg13g2_xnor2_1 _11791_ (.Y(_05186_),
    .A(_05180_),
    .B(_05184_));
 sg13g2_a21oi_1 _11792_ (.A1(net4017),
    .A2(_05186_),
    .Y(_05187_),
    .B1(_05185_));
 sg13g2_xnor2_1 _11793_ (.Y(_05188_),
    .A(\cpu.keccak_alu.registers[20] ),
    .B(_05187_));
 sg13g2_o21ai_1 _11794_ (.B1(_05171_),
    .Y(_05189_),
    .A1(net4382),
    .A2(_05188_));
 sg13g2_nand2_1 _11795_ (.Y(_05190_),
    .A(net101),
    .B(net3696));
 sg13g2_o21ai_1 _11796_ (.B1(_05190_),
    .Y(_05191_),
    .A1(_02302_),
    .A2(_05083_));
 sg13g2_a221oi_1 _11797_ (.B2(net3819),
    .C1(net3732),
    .B1(_05191_),
    .A1(net4263),
    .Y(_05192_),
    .A2(_05189_));
 sg13g2_a21oi_1 _11798_ (.A1(_01031_),
    .A2(net3732),
    .Y(_00737_),
    .B1(_05192_));
 sg13g2_o21ai_1 _11799_ (.B1(_04435_),
    .Y(_05193_),
    .A1(net4562),
    .A2(_00087_));
 sg13g2_nand2_1 _11800_ (.Y(_05194_),
    .A(net3828),
    .B(_05193_));
 sg13g2_nand2_1 _11801_ (.Y(_05195_),
    .A(net4544),
    .B(_05146_));
 sg13g2_o21ai_1 _11802_ (.B1(_05195_),
    .Y(_05196_),
    .A1(net4543),
    .A2(_05194_));
 sg13g2_mux2_1 _11803_ (.A0(_05096_),
    .A1(_05196_),
    .S(net4188),
    .X(_05197_));
 sg13g2_mux2_1 _11804_ (.A0(_04974_),
    .A1(_05197_),
    .S(net4175),
    .X(_05198_));
 sg13g2_nand2_1 _11805_ (.Y(_05199_),
    .A(net4168),
    .B(_05198_));
 sg13g2_o21ai_1 _11806_ (.B1(_05199_),
    .Y(_05200_),
    .A1(net4168),
    .A2(_04704_));
 sg13g2_nand2_1 _11807_ (.Y(_05201_),
    .A(net4089),
    .B(_05200_));
 sg13g2_nand3_1 _11808_ (.B(net3918),
    .C(_04716_),
    .A(net3840),
    .Y(_05202_));
 sg13g2_nor2_1 _11809_ (.A(net3926),
    .B(_04712_),
    .Y(_05203_));
 sg13g2_o21ai_1 _11810_ (.B1(net3776),
    .Y(_05204_),
    .A1(net3919),
    .A2(_04719_));
 sg13g2_o21ai_1 _11811_ (.B1(_05202_),
    .Y(_05205_),
    .A1(_05203_),
    .A2(_05204_));
 sg13g2_o21ai_1 _11812_ (.B1(net4003),
    .Y(_05206_),
    .A1(\cpu.keccak_alu.registers[85] ),
    .A2(_01037_));
 sg13g2_xnor2_1 _11813_ (.Y(_05207_),
    .A(_05201_),
    .B(_05205_));
 sg13g2_o21ai_1 _11814_ (.B1(_05206_),
    .Y(_05208_),
    .A1(net4004),
    .A2(_05207_));
 sg13g2_xor2_1 _11815_ (.B(_05208_),
    .A(\cpu.keccak_alu.registers[21] ),
    .X(_05209_));
 sg13g2_o21ai_1 _11816_ (.B1(net4211),
    .Y(_05210_),
    .A1(\cpu.keccak_alu.registers[149] ),
    .A2(\cpu.keccak_alu.registers[213] ));
 sg13g2_a21oi_1 _11817_ (.A1(\cpu.keccak_alu.registers[149] ),
    .A2(\cpu.keccak_alu.registers[213] ),
    .Y(_05211_),
    .B1(_05210_));
 sg13g2_xor2_1 _11818_ (.B(\cpu.keccak_alu.registers[85] ),
    .A(\cpu.keccak_alu.registers[21] ),
    .X(_05212_));
 sg13g2_o21ai_1 _11819_ (.B1(net4383),
    .Y(_05213_),
    .A1(_05211_),
    .A2(_05212_));
 sg13g2_a21o_1 _11820_ (.A2(_05212_),
    .A1(_05211_),
    .B1(_05213_),
    .X(_05214_));
 sg13g2_o21ai_1 _11821_ (.B1(_05214_),
    .Y(_05215_),
    .A1(net4383),
    .A2(_05209_));
 sg13g2_a22oi_1 _11822_ (.Y(_05216_),
    .B1(net3696),
    .B2(net221),
    .A2(_05081_),
    .A1(_02303_));
 sg13g2_o21ai_1 _11823_ (.B1(net3738),
    .Y(_05217_),
    .A1(net3812),
    .A2(_05216_));
 sg13g2_a21oi_1 _11824_ (.A1(net4263),
    .A2(_05215_),
    .Y(_05218_),
    .B1(_05217_));
 sg13g2_a21oi_1 _11825_ (.A1(_01039_),
    .A2(net3730),
    .Y(_00738_),
    .B1(_05218_));
 sg13g2_a21oi_1 _11826_ (.A1(\cpu.keccak_alu.registers[150] ),
    .A2(\cpu.keccak_alu.registers[214] ),
    .Y(_05219_),
    .B1(net4370));
 sg13g2_o21ai_1 _11827_ (.B1(_05219_),
    .Y(_05220_),
    .A1(\cpu.keccak_alu.registers[150] ),
    .A2(\cpu.keccak_alu.registers[214] ));
 sg13g2_xor2_1 _11828_ (.B(\cpu.keccak_alu.registers[86] ),
    .A(\cpu.keccak_alu.registers[22] ),
    .X(_05221_));
 sg13g2_xnor2_1 _11829_ (.Y(_05222_),
    .A(_05220_),
    .B(_05221_));
 sg13g2_nor3_1 _11830_ (.A(\cpu.keccak_alu.registers[86] ),
    .B(_01047_),
    .C(net4016),
    .Y(_05223_));
 sg13g2_nor3_1 _11831_ (.A(net4538),
    .B(_04232_),
    .C(_04235_),
    .Y(_05224_));
 sg13g2_nor3_1 _11832_ (.A(net4194),
    .B(_04231_),
    .C(_04243_),
    .Y(_05225_));
 sg13g2_nor2_1 _11833_ (.A(_05224_),
    .B(_05225_),
    .Y(_05226_));
 sg13g2_nor2_1 _11834_ (.A(net3823),
    .B(_05226_),
    .Y(_05227_));
 sg13g2_mux2_1 _11835_ (.A0(_05121_),
    .A1(_05227_),
    .S(net4182),
    .X(_05228_));
 sg13g2_mux2_1 _11836_ (.A0(_05003_),
    .A1(_05228_),
    .S(net4172),
    .X(_05229_));
 sg13g2_nand2_1 _11837_ (.Y(_05230_),
    .A(net4166),
    .B(_05229_));
 sg13g2_o21ai_1 _11838_ (.B1(_05230_),
    .Y(_05231_),
    .A1(net4166),
    .A2(_04736_));
 sg13g2_nand2_1 _11839_ (.Y(_05232_),
    .A(net4090),
    .B(_05231_));
 sg13g2_nor2_1 _11840_ (.A(net3913),
    .B(_04748_),
    .Y(_05233_));
 sg13g2_o21ai_1 _11841_ (.B1(net3773),
    .Y(_05234_),
    .A1(net3924),
    .A2(_04740_));
 sg13g2_nand3_1 _11842_ (.B(net3915),
    .C(_04751_),
    .A(net3836),
    .Y(_05235_));
 sg13g2_o21ai_1 _11843_ (.B1(_05235_),
    .Y(_05236_),
    .A1(_05233_),
    .A2(_05234_));
 sg13g2_xnor2_1 _11844_ (.Y(_05237_),
    .A(_05232_),
    .B(_05236_));
 sg13g2_a21oi_1 _11845_ (.A1(net4016),
    .A2(_05237_),
    .Y(_05238_),
    .B1(_05223_));
 sg13g2_nand2b_1 _11846_ (.Y(_05239_),
    .B(\cpu.keccak_alu.registers[22] ),
    .A_N(_05238_));
 sg13g2_a21oi_1 _11847_ (.A1(_01042_),
    .A2(_05238_),
    .Y(_05240_),
    .B1(net4383));
 sg13g2_a22oi_1 _11848_ (.Y(_05241_),
    .B1(_05239_),
    .B2(_05240_),
    .A2(_05222_),
    .A1(net4383));
 sg13g2_or2_1 _11849_ (.X(_05242_),
    .B(_05241_),
    .A(net4320));
 sg13g2_a22oi_1 _11850_ (.Y(_05243_),
    .B1(net3696),
    .B2(net444),
    .A2(net3771),
    .A1(_02305_));
 sg13g2_nor2_1 _11851_ (.A(net3814),
    .B(_05243_),
    .Y(_05244_));
 sg13g2_nor2_1 _11852_ (.A(net3731),
    .B(_05244_),
    .Y(_05245_));
 sg13g2_a22oi_1 _11853_ (.Y(_00739_),
    .B1(_05242_),
    .B2(_05245_),
    .A2(net3730),
    .A1(_01049_));
 sg13g2_a21oi_1 _11854_ (.A1(net4502),
    .A2(\cpu.keccak_alu.registers[215] ),
    .Y(_05246_),
    .B1(net4369));
 sg13g2_o21ai_1 _11855_ (.B1(_05246_),
    .Y(_05247_),
    .A1(\cpu.keccak_alu.registers[151] ),
    .A2(\cpu.keccak_alu.registers[215] ));
 sg13g2_xor2_1 _11856_ (.B(\cpu.keccak_alu.registers[87] ),
    .A(\cpu.keccak_alu.registers[23] ),
    .X(_05248_));
 sg13g2_xnor2_1 _11857_ (.Y(_05249_),
    .A(_05247_),
    .B(_05248_));
 sg13g2_a21oi_2 _11858_ (.B1(net3825),
    .Y(_05250_),
    .A2(_04448_),
    .A1(_04445_));
 sg13g2_nor2_1 _11859_ (.A(net4541),
    .B(_05250_),
    .Y(_05251_));
 sg13g2_a21oi_1 _11860_ (.A1(net4542),
    .A2(_05194_),
    .Y(_05252_),
    .B1(_05251_));
 sg13g2_mux2_1 _11861_ (.A0(_05149_),
    .A1(_05252_),
    .S(net4187),
    .X(_05253_));
 sg13g2_and2_1 _11862_ (.A(net4176),
    .B(_05253_),
    .X(_05254_));
 sg13g2_a21oi_1 _11863_ (.A1(net4529),
    .A2(_05031_),
    .Y(_05255_),
    .B1(_05254_));
 sg13g2_a21oi_1 _11864_ (.A1(net4178),
    .A2(_04774_),
    .Y(_05256_),
    .B1(net4170));
 sg13g2_a21o_1 _11865_ (.A2(_05255_),
    .A1(net4170),
    .B1(_05256_),
    .X(_05257_));
 sg13g2_nor2_1 _11866_ (.A(net3933),
    .B(_05257_),
    .Y(_05258_));
 sg13g2_nor2_1 _11867_ (.A(net3919),
    .B(_04788_),
    .Y(_05259_));
 sg13g2_o21ai_1 _11868_ (.B1(net3777),
    .Y(_05260_),
    .A1(net3927),
    .A2(_04782_));
 sg13g2_nand3_1 _11869_ (.B(net3919),
    .C(_04791_),
    .A(net3840),
    .Y(_05261_));
 sg13g2_o21ai_1 _11870_ (.B1(_05261_),
    .Y(_05262_),
    .A1(_05259_),
    .A2(_05260_));
 sg13g2_a21oi_1 _11871_ (.A1(_01052_),
    .A2(net4502),
    .Y(_05263_),
    .B1(net4015));
 sg13g2_xnor2_1 _11872_ (.Y(_05264_),
    .A(_05258_),
    .B(_05262_));
 sg13g2_a21oi_1 _11873_ (.A1(net4015),
    .A2(_05264_),
    .Y(_05265_),
    .B1(_05263_));
 sg13g2_or2_1 _11874_ (.X(_05266_),
    .B(_05265_),
    .A(\cpu.keccak_alu.registers[23] ));
 sg13g2_a21oi_1 _11875_ (.A1(\cpu.keccak_alu.registers[23] ),
    .A2(_05265_),
    .Y(_05267_),
    .B1(net4378));
 sg13g2_a22oi_1 _11876_ (.Y(_05268_),
    .B1(_05266_),
    .B2(_05267_),
    .A2(_05249_),
    .A1(net4378));
 sg13g2_or2_1 _11877_ (.X(_05269_),
    .B(_05268_),
    .A(net4315));
 sg13g2_a22oi_1 _11878_ (.Y(_05270_),
    .B1(net3695),
    .B2(net556),
    .A2(net3771),
    .A1(_02307_));
 sg13g2_nor2_1 _11879_ (.A(net3812),
    .B(_05270_),
    .Y(_05271_));
 sg13g2_nor2_1 _11880_ (.A(net3728),
    .B(_05271_),
    .Y(_05272_));
 sg13g2_a22oi_1 _11881_ (.Y(_00740_),
    .B1(_05269_),
    .B2(_05272_),
    .A2(net3728),
    .A1(_01058_));
 sg13g2_o21ai_1 _11882_ (.B1(net4206),
    .Y(_05273_),
    .A1(net4501),
    .A2(\cpu.keccak_alu.registers[216] ));
 sg13g2_a21oi_1 _11883_ (.A1(net4501),
    .A2(\cpu.keccak_alu.registers[216] ),
    .Y(_05274_),
    .B1(_05273_));
 sg13g2_xor2_1 _11884_ (.B(\cpu.keccak_alu.registers[88] ),
    .A(\cpu.keccak_alu.registers[24] ),
    .X(_05275_));
 sg13g2_a21oi_1 _11885_ (.A1(_05274_),
    .A2(_05275_),
    .Y(_05276_),
    .B1(net4214));
 sg13g2_o21ai_1 _11886_ (.B1(_05276_),
    .Y(_05277_),
    .A1(_05274_),
    .A2(_05275_));
 sg13g2_nor3_1 _11887_ (.A(net4538),
    .B(_04212_),
    .C(_04236_),
    .Y(_05278_));
 sg13g2_nor3_1 _11888_ (.A(net4195),
    .B(_04232_),
    .C(_04235_),
    .Y(_05279_));
 sg13g2_nor2_1 _11889_ (.A(_05278_),
    .B(_05279_),
    .Y(_05280_));
 sg13g2_nor2_1 _11890_ (.A(net3823),
    .B(_05280_),
    .Y(_05281_));
 sg13g2_mux2_1 _11891_ (.A0(_05175_),
    .A1(_05281_),
    .S(net4182),
    .X(_05282_));
 sg13g2_mux2_1 _11892_ (.A0(_05063_),
    .A1(_05282_),
    .S(net4171),
    .X(_05283_));
 sg13g2_mux2_1 _11893_ (.A0(_04817_),
    .A1(_05283_),
    .S(net4164),
    .X(_05284_));
 sg13g2_inv_1 _11894_ (.Y(_05285_),
    .A(_05284_));
 sg13g2_nor2_1 _11895_ (.A(net3931),
    .B(_05285_),
    .Y(_05286_));
 sg13g2_nand3_1 _11896_ (.B(net3917),
    .C(_04820_),
    .A(net3836),
    .Y(_05287_));
 sg13g2_and2_1 _11897_ (.A(net3914),
    .B(_04822_),
    .X(_05288_));
 sg13g2_o21ai_1 _11898_ (.B1(net3772),
    .Y(_05289_),
    .A1(net3913),
    .A2(_04819_));
 sg13g2_o21ai_1 _11899_ (.B1(_05287_),
    .Y(_05290_),
    .A1(_05288_),
    .A2(_05289_));
 sg13g2_a21oi_1 _11900_ (.A1(_01063_),
    .A2(\cpu.keccak_alu.registers[152] ),
    .Y(_05291_),
    .B1(net4014));
 sg13g2_or4_1 _11901_ (.A(net4517),
    .B(net4513),
    .C(_05285_),
    .D(_05287_),
    .X(_05292_));
 sg13g2_o21ai_1 _11902_ (.B1(_05292_),
    .Y(_05293_),
    .A1(_05286_),
    .A2(_05290_));
 sg13g2_a21oi_1 _11903_ (.A1(net4014),
    .A2(_05293_),
    .Y(_05294_),
    .B1(_05291_));
 sg13g2_xnor2_1 _11904_ (.Y(_05295_),
    .A(\cpu.keccak_alu.registers[24] ),
    .B(_05294_));
 sg13g2_o21ai_1 _11905_ (.B1(_05277_),
    .Y(_05296_),
    .A1(net4379),
    .A2(_05295_));
 sg13g2_a22oi_1 _11906_ (.Y(_05297_),
    .B1(net3695),
    .B2(net346),
    .A2(net3771),
    .A1(_02309_));
 sg13g2_o21ai_1 _11907_ (.B1(net3738),
    .Y(_05298_),
    .A1(net3812),
    .A2(_05297_));
 sg13g2_a21oi_1 _11908_ (.A1(net4258),
    .A2(_05296_),
    .Y(_05299_),
    .B1(_05298_));
 sg13g2_a21oi_1 _11909_ (.A1(_01067_),
    .A2(net3726),
    .Y(_00741_),
    .B1(_05299_));
 sg13g2_o21ai_1 _11910_ (.B1(_04446_),
    .Y(_05300_),
    .A1(net4564),
    .A2(_00091_));
 sg13g2_nand2_1 _11911_ (.Y(_05301_),
    .A(net3828),
    .B(_05300_));
 sg13g2_nand2_1 _11912_ (.Y(_05302_),
    .A(net4541),
    .B(_05250_));
 sg13g2_o21ai_1 _11913_ (.B1(_05302_),
    .Y(_05303_),
    .A1(net4541),
    .A2(_05301_));
 sg13g2_mux2_1 _11914_ (.A0(_05196_),
    .A1(_05303_),
    .S(net4187),
    .X(_05304_));
 sg13g2_mux2_1 _11915_ (.A0(_05097_),
    .A1(_05304_),
    .S(net4177),
    .X(_05305_));
 sg13g2_nor2_1 _11916_ (.A(net4169),
    .B(_04845_),
    .Y(_05306_));
 sg13g2_a21oi_1 _11917_ (.A1(net4169),
    .A2(_05305_),
    .Y(_05307_),
    .B1(_05306_));
 sg13g2_nor2_1 _11918_ (.A(_03872_),
    .B(_05307_),
    .Y(_05308_));
 sg13g2_and2_1 _11919_ (.A(net3921),
    .B(_04854_),
    .X(_05309_));
 sg13g2_mux2_1 _11920_ (.A0(_04848_),
    .A1(_04853_),
    .S(net3926),
    .X(_05310_));
 sg13g2_a22oi_1 _11921_ (.Y(_05311_),
    .B1(_05310_),
    .B2(net3777),
    .A2(_05309_),
    .A1(net3839));
 sg13g2_a21oi_1 _11922_ (.A1(_01073_),
    .A2(net4500),
    .Y(_05312_),
    .B1(net4009));
 sg13g2_xor2_1 _11923_ (.B(_05311_),
    .A(_05308_),
    .X(_05313_));
 sg13g2_a21oi_1 _11924_ (.A1(net4009),
    .A2(_05313_),
    .Y(_05314_),
    .B1(_05312_));
 sg13g2_or2_1 _11925_ (.X(_05315_),
    .B(_05314_),
    .A(\cpu.keccak_alu.registers[25] ));
 sg13g2_a21oi_1 _11926_ (.A1(\cpu.keccak_alu.registers[25] ),
    .A2(_05314_),
    .Y(_05316_),
    .B1(net4371));
 sg13g2_a21oi_1 _11927_ (.A1(net4500),
    .A2(\cpu.keccak_alu.registers[217] ),
    .Y(_05317_),
    .B1(net4366));
 sg13g2_o21ai_1 _11928_ (.B1(_05317_),
    .Y(_05318_),
    .A1(net4500),
    .A2(\cpu.keccak_alu.registers[217] ));
 sg13g2_xor2_1 _11929_ (.B(\cpu.keccak_alu.registers[89] ),
    .A(\cpu.keccak_alu.registers[25] ),
    .X(_05319_));
 sg13g2_xnor2_1 _11930_ (.Y(_05320_),
    .A(_05318_),
    .B(_05319_));
 sg13g2_a22oi_1 _11931_ (.Y(_05321_),
    .B1(_05320_),
    .B2(net4371),
    .A2(_05316_),
    .A1(_05315_));
 sg13g2_or2_1 _11932_ (.X(_05322_),
    .B(_05321_),
    .A(net4313));
 sg13g2_nand2_1 _11933_ (.Y(_05323_),
    .A(net562),
    .B(net3695));
 sg13g2_o21ai_1 _11934_ (.B1(_05323_),
    .Y(_05324_),
    .A1(_02312_),
    .A2(net3718));
 sg13g2_a21oi_1 _11935_ (.A1(net3815),
    .A2(_05324_),
    .Y(_05325_),
    .B1(net3720));
 sg13g2_a22oi_1 _11936_ (.Y(_00742_),
    .B1(_05322_),
    .B2(_05325_),
    .A2(net3719),
    .A1(_01075_));
 sg13g2_nor3_1 _11937_ (.A(net4538),
    .B(_04209_),
    .C(_04213_),
    .Y(_05326_));
 sg13g2_nor3_1 _11938_ (.A(net4195),
    .B(_04212_),
    .C(_04236_),
    .Y(_05327_));
 sg13g2_nor2_1 _11939_ (.A(_05326_),
    .B(_05327_),
    .Y(_05328_));
 sg13g2_nor2_1 _11940_ (.A(net3822),
    .B(_05328_),
    .Y(_05329_));
 sg13g2_mux2_1 _11941_ (.A0(_05227_),
    .A1(_05329_),
    .S(net4182),
    .X(_05330_));
 sg13g2_mux2_1 _11942_ (.A0(_05122_),
    .A1(_05330_),
    .S(net4171),
    .X(_05331_));
 sg13g2_mux2_1 _11943_ (.A0(_04878_),
    .A1(_05331_),
    .S(net4164),
    .X(_05332_));
 sg13g2_inv_1 _11944_ (.Y(_05333_),
    .A(_05332_));
 sg13g2_nor2_1 _11945_ (.A(net3931),
    .B(_05333_),
    .Y(_05334_));
 sg13g2_nand3_1 _11946_ (.B(net3917),
    .C(_04882_),
    .A(net3836),
    .Y(_05335_));
 sg13g2_nor2_1 _11947_ (.A(net3924),
    .B(_04884_),
    .Y(_05336_));
 sg13g2_o21ai_1 _11948_ (.B1(net3772),
    .Y(_05337_),
    .A1(net3915),
    .A2(_04881_));
 sg13g2_o21ai_1 _11949_ (.B1(_05335_),
    .Y(_05338_),
    .A1(_05336_),
    .A2(_05337_));
 sg13g2_a21oi_1 _11950_ (.A1(_01079_),
    .A2(\cpu.keccak_alu.registers[154] ),
    .Y(_05339_),
    .B1(net4010));
 sg13g2_or4_1 _11951_ (.A(net4517),
    .B(net4513),
    .C(_05333_),
    .D(_05335_),
    .X(_05340_));
 sg13g2_o21ai_1 _11952_ (.B1(_05340_),
    .Y(_05341_),
    .A1(_05334_),
    .A2(_05338_));
 sg13g2_a21oi_1 _11953_ (.A1(net4010),
    .A2(_05341_),
    .Y(_05342_),
    .B1(_05339_));
 sg13g2_o21ai_1 _11954_ (.B1(net4213),
    .Y(_05343_),
    .A1(\cpu.keccak_alu.registers[26] ),
    .A2(_05342_));
 sg13g2_a21oi_1 _11955_ (.A1(\cpu.keccak_alu.registers[26] ),
    .A2(_05342_),
    .Y(_05344_),
    .B1(_05343_));
 sg13g2_a21oi_1 _11956_ (.A1(\cpu.keccak_alu.registers[154] ),
    .A2(\cpu.keccak_alu.registers[218] ),
    .Y(_05345_),
    .B1(net4366));
 sg13g2_o21ai_1 _11957_ (.B1(_05345_),
    .Y(_05346_),
    .A1(\cpu.keccak_alu.registers[154] ),
    .A2(\cpu.keccak_alu.registers[218] ));
 sg13g2_xnor2_1 _11958_ (.Y(_05347_),
    .A(\cpu.keccak_alu.registers[26] ),
    .B(\cpu.keccak_alu.registers[90] ));
 sg13g2_o21ai_1 _11959_ (.B1(net4371),
    .Y(_05348_),
    .A1(_05346_),
    .A2(_05347_));
 sg13g2_a21oi_1 _11960_ (.A1(_05346_),
    .A2(_05347_),
    .Y(_05349_),
    .B1(_05348_));
 sg13g2_o21ai_1 _11961_ (.B1(net4244),
    .Y(_05350_),
    .A1(_05344_),
    .A2(_05349_));
 sg13g2_nand2_1 _11962_ (.Y(_05351_),
    .A(net697),
    .B(net3695));
 sg13g2_o21ai_1 _11963_ (.B1(_05351_),
    .Y(_05352_),
    .A1(_02314_),
    .A2(net3718));
 sg13g2_a21oi_1 _11964_ (.A1(net3815),
    .A2(_05352_),
    .Y(_05353_),
    .B1(net3720));
 sg13g2_a22oi_1 _11965_ (.Y(_00743_),
    .B1(_05350_),
    .B2(_05353_),
    .A2(net3720),
    .A1(_01082_));
 sg13g2_nor2b_1 _11966_ (.A(\cpu.keccak_alu.registers[91] ),
    .B_N(net4499),
    .Y(_05354_));
 sg13g2_nand2b_1 _11967_ (.Y(_05355_),
    .B(_04420_),
    .A_N(_04416_));
 sg13g2_nand3_1 _11968_ (.B(net3828),
    .C(_05355_),
    .A(net4199),
    .Y(_05356_));
 sg13g2_o21ai_1 _11969_ (.B1(_05356_),
    .Y(_05357_),
    .A1(net4199),
    .A2(_05301_));
 sg13g2_mux2_1 _11970_ (.A0(_05252_),
    .A1(_05357_),
    .S(net4187),
    .X(_05358_));
 sg13g2_mux2_1 _11971_ (.A0(_05150_),
    .A1(_05358_),
    .S(net4174),
    .X(_05359_));
 sg13g2_mux2_1 _11972_ (.A0(_04905_),
    .A1(_05359_),
    .S(net4168),
    .X(_05360_));
 sg13g2_inv_1 _11973_ (.Y(_05361_),
    .A(_05360_));
 sg13g2_nor2_2 _11974_ (.A(_03872_),
    .B(_05361_),
    .Y(_05362_));
 sg13g2_nand4_1 _11975_ (.B(net3920),
    .C(net3785),
    .A(net3840),
    .Y(_05363_),
    .D(_04609_));
 sg13g2_nor2_1 _11976_ (.A(net3928),
    .B(_04907_),
    .Y(_05364_));
 sg13g2_o21ai_1 _11977_ (.B1(net3776),
    .Y(_05365_),
    .A1(net3920),
    .A2(_04912_));
 sg13g2_o21ai_1 _11978_ (.B1(_05363_),
    .Y(_05366_),
    .A1(_05364_),
    .A2(_05365_));
 sg13g2_or2_1 _11979_ (.X(_05367_),
    .B(_05366_),
    .A(_05362_));
 sg13g2_a21oi_1 _11980_ (.A1(_05362_),
    .A2(_05366_),
    .Y(_05368_),
    .B1(net4001));
 sg13g2_a22oi_1 _11981_ (.Y(_05369_),
    .B1(_05367_),
    .B2(_05368_),
    .A2(_05354_),
    .A1(net4000));
 sg13g2_nand2b_1 _11982_ (.Y(_05370_),
    .B(\cpu.keccak_alu.registers[27] ),
    .A_N(_05369_));
 sg13g2_a21oi_1 _11983_ (.A1(_01085_),
    .A2(_05369_),
    .Y(_05371_),
    .B1(net4374));
 sg13g2_a21oi_1 _11984_ (.A1(net4499),
    .A2(\cpu.keccak_alu.registers[219] ),
    .Y(_05372_),
    .B1(net4367));
 sg13g2_o21ai_1 _11985_ (.B1(_05372_),
    .Y(_05373_),
    .A1(net4499),
    .A2(\cpu.keccak_alu.registers[219] ));
 sg13g2_xor2_1 _11986_ (.B(\cpu.keccak_alu.registers[91] ),
    .A(\cpu.keccak_alu.registers[27] ),
    .X(_05374_));
 sg13g2_xnor2_1 _11987_ (.Y(_05375_),
    .A(_05373_),
    .B(_05374_));
 sg13g2_a22oi_1 _11988_ (.Y(_05376_),
    .B1(_05375_),
    .B2(net4374),
    .A2(_05371_),
    .A1(_05370_));
 sg13g2_or2_1 _11989_ (.X(_05377_),
    .B(_05376_),
    .A(net4313));
 sg13g2_nand2_1 _11990_ (.Y(_05378_),
    .A(net499),
    .B(net3695));
 sg13g2_o21ai_1 _11991_ (.B1(_05378_),
    .Y(_05379_),
    .A1(_02316_),
    .A2(net3718));
 sg13g2_a21oi_1 _11992_ (.A1(net3815),
    .A2(_05379_),
    .Y(_05380_),
    .B1(net3721));
 sg13g2_a22oi_1 _11993_ (.Y(_00744_),
    .B1(_05377_),
    .B2(_05380_),
    .A2(net3721),
    .A1(_01091_));
 sg13g2_nor3_1 _11994_ (.A(net4537),
    .B(_04210_),
    .C(_04224_),
    .Y(_05381_));
 sg13g2_nor3_1 _11995_ (.A(net4195),
    .B(_04209_),
    .C(_04213_),
    .Y(_05382_));
 sg13g2_nor2_1 _11996_ (.A(_05381_),
    .B(_05382_),
    .Y(_05383_));
 sg13g2_nor2_1 _11997_ (.A(net3822),
    .B(_05383_),
    .Y(_05384_));
 sg13g2_mux2_1 _11998_ (.A0(_05281_),
    .A1(_05384_),
    .S(net4182),
    .X(_05385_));
 sg13g2_mux2_1 _11999_ (.A0(_05176_),
    .A1(_05385_),
    .S(net4171),
    .X(_05386_));
 sg13g2_mux2_1 _12000_ (.A0(_04937_),
    .A1(_05386_),
    .S(net4164),
    .X(_05387_));
 sg13g2_nand2_1 _12001_ (.Y(_05388_),
    .A(net4090),
    .B(_05387_));
 sg13g2_nor2_1 _12002_ (.A(net3923),
    .B(_04942_),
    .Y(_05389_));
 sg13g2_mux2_1 _12003_ (.A0(_04940_),
    .A1(_04947_),
    .S(net3913),
    .X(_05390_));
 sg13g2_a22oi_1 _12004_ (.Y(_05391_),
    .B1(_05390_),
    .B2(net3772),
    .A2(_05389_),
    .A1(net3836));
 sg13g2_o21ai_1 _12005_ (.B1(net4003),
    .Y(_05392_),
    .A1(\cpu.keccak_alu.registers[92] ),
    .A2(_01097_));
 sg13g2_xor2_1 _12006_ (.B(_05391_),
    .A(_05388_),
    .X(_05393_));
 sg13g2_o21ai_1 _12007_ (.B1(_05392_),
    .Y(_05394_),
    .A1(net4003),
    .A2(_05393_));
 sg13g2_nand2b_1 _12008_ (.Y(_05395_),
    .B(\cpu.keccak_alu.registers[28] ),
    .A_N(_05394_));
 sg13g2_a21oi_1 _12009_ (.A1(_01094_),
    .A2(_05394_),
    .Y(_05396_),
    .B1(net4377));
 sg13g2_a21oi_1 _12010_ (.A1(\cpu.keccak_alu.registers[156] ),
    .A2(\cpu.keccak_alu.registers[220] ),
    .Y(_05397_),
    .B1(net4369));
 sg13g2_o21ai_1 _12011_ (.B1(_05397_),
    .Y(_05398_),
    .A1(\cpu.keccak_alu.registers[156] ),
    .A2(\cpu.keccak_alu.registers[220] ));
 sg13g2_xor2_1 _12012_ (.B(\cpu.keccak_alu.registers[92] ),
    .A(\cpu.keccak_alu.registers[28] ),
    .X(_05399_));
 sg13g2_xnor2_1 _12013_ (.Y(_05400_),
    .A(_05398_),
    .B(_05399_));
 sg13g2_a22oi_1 _12014_ (.Y(_05401_),
    .B1(_05400_),
    .B2(net4377),
    .A2(_05396_),
    .A1(_05395_));
 sg13g2_or2_1 _12015_ (.X(_05402_),
    .B(_05401_),
    .A(net4318));
 sg13g2_nand2_1 _12016_ (.Y(_05403_),
    .A(net546),
    .B(net3696));
 sg13g2_o21ai_1 _12017_ (.B1(_05403_),
    .Y(_05404_),
    .A1(_02317_),
    .A2(net3718));
 sg13g2_a21oi_1 _12018_ (.A1(net3818),
    .A2(_05404_),
    .Y(_05405_),
    .B1(net3727));
 sg13g2_a22oi_1 _12019_ (.Y(_00745_),
    .B1(_05402_),
    .B2(_05405_),
    .A2(net3727),
    .A1(_01100_));
 sg13g2_o21ai_1 _12020_ (.B1(net4206),
    .Y(_05406_),
    .A1(net4498),
    .A2(\cpu.keccak_alu.registers[221] ));
 sg13g2_a21oi_1 _12021_ (.A1(net4498),
    .A2(\cpu.keccak_alu.registers[221] ),
    .Y(_05407_),
    .B1(_05406_));
 sg13g2_xor2_1 _12022_ (.B(\cpu.keccak_alu.registers[93] ),
    .A(\cpu.keccak_alu.registers[29] ),
    .X(_05408_));
 sg13g2_a21oi_1 _12023_ (.A1(_05407_),
    .A2(_05408_),
    .Y(_05409_),
    .B1(net4213));
 sg13g2_o21ai_1 _12024_ (.B1(_05409_),
    .Y(_05410_),
    .A1(_05407_),
    .A2(_05408_));
 sg13g2_o21ai_1 _12025_ (.B1(_04417_),
    .Y(_05411_),
    .A1(net4565),
    .A2(_00095_));
 sg13g2_nand3_1 _12026_ (.B(net3830),
    .C(_05411_),
    .A(net4199),
    .Y(_05412_));
 sg13g2_nand3_1 _12027_ (.B(net3830),
    .C(_05355_),
    .A(net4541),
    .Y(_05413_));
 sg13g2_nand2_1 _12028_ (.Y(_05414_),
    .A(_05412_),
    .B(_05413_));
 sg13g2_mux2_1 _12029_ (.A0(_05303_),
    .A1(_05414_),
    .S(net4187),
    .X(_05415_));
 sg13g2_mux2_1 _12030_ (.A0(_05197_),
    .A1(_05415_),
    .S(net4175),
    .X(_05416_));
 sg13g2_mux2_1 _12031_ (.A0(_04976_),
    .A1(_05416_),
    .S(net4168),
    .X(_05417_));
 sg13g2_nand2_1 _12032_ (.Y(_05418_),
    .A(net4089),
    .B(_05417_));
 sg13g2_nor2_1 _12033_ (.A(net3926),
    .B(_04979_),
    .Y(_05419_));
 sg13g2_o21ai_1 _12034_ (.B1(net3776),
    .Y(_05420_),
    .A1(net3919),
    .A2(_04984_));
 sg13g2_nand4_1 _12035_ (.B(net3918),
    .C(net3785),
    .A(net3840),
    .Y(_05421_),
    .D(_04714_));
 sg13g2_o21ai_1 _12036_ (.B1(_05421_),
    .Y(_05422_),
    .A1(_05419_),
    .A2(_05420_));
 sg13g2_a21oi_1 _12037_ (.A1(_01104_),
    .A2(net4498),
    .Y(_05423_),
    .B1(net4012));
 sg13g2_xor2_1 _12038_ (.B(_05422_),
    .A(_05418_),
    .X(_05424_));
 sg13g2_a21oi_1 _12039_ (.A1(net4012),
    .A2(_05424_),
    .Y(_05425_),
    .B1(_05423_));
 sg13g2_xnor2_1 _12040_ (.Y(_05426_),
    .A(\cpu.keccak_alu.registers[29] ),
    .B(_05425_));
 sg13g2_o21ai_1 _12041_ (.B1(_05410_),
    .Y(_05427_),
    .A1(net4373),
    .A2(_05426_));
 sg13g2_nand2_1 _12042_ (.Y(_05428_),
    .A(net165),
    .B(net3695));
 sg13g2_o21ai_1 _12043_ (.B1(_05428_),
    .Y(_05429_),
    .A1(_02320_),
    .A2(net3718));
 sg13g2_a221oi_1 _12044_ (.B2(net3816),
    .C1(net3722),
    .B1(_05429_),
    .A1(net4244),
    .Y(_05430_),
    .A2(_05427_));
 sg13g2_a21oi_1 _12045_ (.A1(_01108_),
    .A2(net3722),
    .Y(_00746_),
    .B1(_05430_));
 sg13g2_nor3_1 _12046_ (.A(net4536),
    .B(_04221_),
    .C(_04225_),
    .Y(_05431_));
 sg13g2_nor3_1 _12047_ (.A(net4195),
    .B(_04210_),
    .C(_04224_),
    .Y(_05432_));
 sg13g2_nor2_1 _12048_ (.A(_05431_),
    .B(_05432_),
    .Y(_05433_));
 sg13g2_nor2_1 _12049_ (.A(net3822),
    .B(_05433_),
    .Y(_05434_));
 sg13g2_mux2_1 _12050_ (.A0(_05329_),
    .A1(_05434_),
    .S(net4181),
    .X(_05435_));
 sg13g2_mux2_1 _12051_ (.A0(_05228_),
    .A1(_05435_),
    .S(net4172),
    .X(_05436_));
 sg13g2_mux2_1 _12052_ (.A0(_05005_),
    .A1(_05436_),
    .S(net4165),
    .X(_05437_));
 sg13g2_nand2_1 _12053_ (.Y(_05438_),
    .A(net4090),
    .B(_05437_));
 sg13g2_nor2_1 _12054_ (.A(net3923),
    .B(_05011_),
    .Y(_05439_));
 sg13g2_and3_1 _12055_ (.X(_05440_),
    .A(net3913),
    .B(net3781),
    .C(_04749_));
 sg13g2_nand2_1 _12056_ (.Y(_05441_),
    .A(net3836),
    .B(_05440_));
 sg13g2_o21ai_1 _12057_ (.B1(net3772),
    .Y(_05442_),
    .A1(net3913),
    .A2(_05008_));
 sg13g2_o21ai_1 _12058_ (.B1(_05441_),
    .Y(_05443_),
    .A1(_05439_),
    .A2(_05442_));
 sg13g2_a21oi_1 _12059_ (.A1(_01119_),
    .A2(\cpu.keccak_alu.registers[158] ),
    .Y(_05444_),
    .B1(net4010));
 sg13g2_xor2_1 _12060_ (.B(_05443_),
    .A(_05438_),
    .X(_05445_));
 sg13g2_a21oi_1 _12061_ (.A1(net4010),
    .A2(_05445_),
    .Y(_05446_),
    .B1(_05444_));
 sg13g2_o21ai_1 _12062_ (.B1(net4213),
    .Y(_05447_),
    .A1(\cpu.keccak_alu.registers[30] ),
    .A2(_05446_));
 sg13g2_a21oi_1 _12063_ (.A1(net952),
    .A2(_05446_),
    .Y(_05448_),
    .B1(_05447_));
 sg13g2_o21ai_1 _12064_ (.B1(net4206),
    .Y(_05449_),
    .A1(\cpu.keccak_alu.registers[158] ),
    .A2(\cpu.keccak_alu.registers[222] ));
 sg13g2_a21oi_1 _12065_ (.A1(\cpu.keccak_alu.registers[158] ),
    .A2(\cpu.keccak_alu.registers[222] ),
    .Y(_05450_),
    .B1(_05449_));
 sg13g2_xor2_1 _12066_ (.B(\cpu.keccak_alu.registers[94] ),
    .A(\cpu.keccak_alu.registers[30] ),
    .X(_05451_));
 sg13g2_o21ai_1 _12067_ (.B1(net4373),
    .Y(_05452_),
    .A1(_05450_),
    .A2(_05451_));
 sg13g2_a21oi_1 _12068_ (.A1(_05450_),
    .A2(_05451_),
    .Y(_05453_),
    .B1(_05452_));
 sg13g2_o21ai_1 _12069_ (.B1(net4244),
    .Y(_05454_),
    .A1(_05448_),
    .A2(_05453_));
 sg13g2_nand2_1 _12070_ (.Y(_05455_),
    .A(net511),
    .B(net3695));
 sg13g2_o21ai_1 _12071_ (.B1(_05455_),
    .Y(_05456_),
    .A1(_02321_),
    .A2(net3718));
 sg13g2_a21oi_1 _12072_ (.A1(net3815),
    .A2(_05456_),
    .Y(_05457_),
    .B1(net3719));
 sg13g2_a22oi_1 _12073_ (.Y(_00747_),
    .B1(_05454_),
    .B2(_05457_),
    .A2(net3720),
    .A1(_01123_));
 sg13g2_nand3b_1 _12074_ (.B(\cpu.keccak_alu.registers[159] ),
    .C(net4002),
    .Y(_05458_),
    .A_N(\cpu.keccak_alu.registers[95] ));
 sg13g2_nand2b_1 _12075_ (.Y(_05459_),
    .B(_04431_),
    .A_N(_04427_));
 sg13g2_nand3_1 _12076_ (.B(net3830),
    .C(_05459_),
    .A(net4199),
    .Y(_05460_));
 sg13g2_nand3_1 _12077_ (.B(net3830),
    .C(_05411_),
    .A(net4541),
    .Y(_05461_));
 sg13g2_nand2_1 _12078_ (.Y(_05462_),
    .A(_05460_),
    .B(_05461_));
 sg13g2_mux2_1 _12079_ (.A0(_05357_),
    .A1(_05462_),
    .S(net4187),
    .X(_05463_));
 sg13g2_mux2_1 _12080_ (.A0(_05253_),
    .A1(_05463_),
    .S(net4176),
    .X(_05464_));
 sg13g2_mux2_1 _12081_ (.A0(_05033_),
    .A1(_05464_),
    .S(net4170),
    .X(_05465_));
 sg13g2_nand2_1 _12082_ (.Y(_05466_),
    .A(net4089),
    .B(_05465_));
 sg13g2_nor2_1 _12083_ (.A(net3918),
    .B(_05040_),
    .Y(_05467_));
 sg13g2_o21ai_1 _12084_ (.B1(net3777),
    .Y(_05468_),
    .A1(net3927),
    .A2(_05037_));
 sg13g2_nor4_2 _12085_ (.A(net4576),
    .B(net3926),
    .C(_03880_),
    .Y(_05469_),
    .D(net3541));
 sg13g2_nand2_1 _12086_ (.Y(_05470_),
    .A(net3840),
    .B(_05469_));
 sg13g2_o21ai_1 _12087_ (.B1(_05470_),
    .Y(_05471_),
    .A1(_05467_),
    .A2(_05468_));
 sg13g2_xor2_1 _12088_ (.B(_05471_),
    .A(_05466_),
    .X(_05472_));
 sg13g2_o21ai_1 _12089_ (.B1(_05458_),
    .Y(_05473_),
    .A1(net4002),
    .A2(_05472_));
 sg13g2_xnor2_1 _12090_ (.Y(_05474_),
    .A(\cpu.keccak_alu.registers[31] ),
    .B(_05473_));
 sg13g2_o21ai_1 _12091_ (.B1(net4207),
    .Y(_05475_),
    .A1(\cpu.keccak_alu.registers[159] ),
    .A2(\cpu.keccak_alu.registers[223] ));
 sg13g2_a21oi_1 _12092_ (.A1(\cpu.keccak_alu.registers[159] ),
    .A2(\cpu.keccak_alu.registers[223] ),
    .Y(_05476_),
    .B1(_05475_));
 sg13g2_xor2_1 _12093_ (.B(\cpu.keccak_alu.registers[95] ),
    .A(\cpu.keccak_alu.registers[31] ),
    .X(_05477_));
 sg13g2_a21oi_1 _12094_ (.A1(_05476_),
    .A2(_05477_),
    .Y(_05478_),
    .B1(net4213));
 sg13g2_o21ai_1 _12095_ (.B1(_05478_),
    .Y(_05479_),
    .A1(_05476_),
    .A2(_05477_));
 sg13g2_o21ai_1 _12096_ (.B1(_05479_),
    .Y(_05480_),
    .A1(net4375),
    .A2(_05474_));
 sg13g2_nand2_1 _12097_ (.Y(_05481_),
    .A(net196),
    .B(net3695));
 sg13g2_o21ai_1 _12098_ (.B1(_05481_),
    .Y(_05482_),
    .A1(_02324_),
    .A2(net3718));
 sg13g2_a221oi_1 _12099_ (.B2(net3818),
    .C1(net3724),
    .B1(_05482_),
    .A1(net4258),
    .Y(_05483_),
    .A2(_05480_));
 sg13g2_a21oi_1 _12100_ (.A1(_01136_),
    .A2(net3724),
    .Y(_00748_),
    .B1(_05483_));
 sg13g2_a21oi_1 _12101_ (.A1(net4497),
    .A2(\cpu.keccak_alu.registers[224] ),
    .Y(_05484_),
    .B1(\cpu.current_instruction[15] ));
 sg13g2_o21ai_1 _12102_ (.B1(_05484_),
    .Y(_05485_),
    .A1(net4497),
    .A2(\cpu.keccak_alu.registers[224] ));
 sg13g2_xnor2_1 _12103_ (.Y(_05486_),
    .A(\cpu.keccak_alu.registers[32] ),
    .B(\cpu.keccak_alu.registers[96] ));
 sg13g2_xnor2_1 _12104_ (.Y(_05487_),
    .A(_05485_),
    .B(_05486_));
 sg13g2_nor2_1 _12105_ (.A(net4167),
    .B(_05065_),
    .Y(_05488_));
 sg13g2_nor3_1 _12106_ (.A(net4536),
    .B(_04139_),
    .C(_04222_),
    .Y(_05489_));
 sg13g2_nor3_1 _12107_ (.A(net4195),
    .B(_04221_),
    .C(_04225_),
    .Y(_05490_));
 sg13g2_nor2_1 _12108_ (.A(_05489_),
    .B(_05490_),
    .Y(_05491_));
 sg13g2_nor2_1 _12109_ (.A(net3821),
    .B(_05491_),
    .Y(_05492_));
 sg13g2_mux2_1 _12110_ (.A0(_05384_),
    .A1(_05492_),
    .S(net4182),
    .X(_05493_));
 sg13g2_mux2_1 _12111_ (.A0(_05282_),
    .A1(_05493_),
    .S(net4171),
    .X(_05494_));
 sg13g2_o21ai_1 _12112_ (.B1(net4518),
    .Y(_05495_),
    .A1(net4521),
    .A2(_04304_));
 sg13g2_o21ai_1 _12113_ (.B1(_05495_),
    .Y(_05496_),
    .A1(net3937),
    .A2(_05494_));
 sg13g2_nor2_1 _12114_ (.A(_05488_),
    .B(_05496_),
    .Y(_05497_));
 sg13g2_a22oi_1 _12115_ (.Y(_05498_),
    .B1(_05497_),
    .B2(net4158),
    .A2(net3774),
    .A1(_04207_));
 sg13g2_nand3b_1 _12116_ (.B(\cpu.keccak_alu.registers[160] ),
    .C(net4005),
    .Y(_05499_),
    .A_N(\cpu.keccak_alu.registers[96] ));
 sg13g2_o21ai_1 _12117_ (.B1(_05499_),
    .Y(_05500_),
    .A1(net4005),
    .A2(_05498_));
 sg13g2_a21oi_1 _12118_ (.A1(\cpu.keccak_alu.registers[32] ),
    .A2(_05500_),
    .Y(_05501_),
    .B1(net4385));
 sg13g2_o21ai_1 _12119_ (.B1(_05501_),
    .Y(_05502_),
    .A1(\cpu.keccak_alu.registers[32] ),
    .A2(_05500_));
 sg13g2_o21ai_1 _12120_ (.B1(_05502_),
    .Y(_05503_),
    .A1(net4219),
    .A2(_05487_));
 sg13g2_nor3_1 _12121_ (.A(net4447),
    .B(net3760),
    .C(_05083_),
    .Y(_05504_));
 sg13g2_nand2_1 _12122_ (.Y(_05505_),
    .A(_02328_),
    .B(_05082_));
 sg13g2_a22oi_1 _12123_ (.Y(_05506_),
    .B1(_05505_),
    .B2(net153),
    .A2(_05082_),
    .A1(_02330_));
 sg13g2_o21ai_1 _12124_ (.B1(net3739),
    .Y(_05507_),
    .A1(net3813),
    .A2(_05506_));
 sg13g2_a21oi_1 _12125_ (.A1(net4265),
    .A2(_05503_),
    .Y(_05508_),
    .B1(_05507_));
 sg13g2_a21oi_1 _12126_ (.A1(_00999_),
    .A2(net3736),
    .Y(_00749_),
    .B1(_05508_));
 sg13g2_o21ai_1 _12127_ (.B1(net4209),
    .Y(_05509_),
    .A1(net4496),
    .A2(\cpu.keccak_alu.registers[225] ));
 sg13g2_a21oi_1 _12128_ (.A1(net4496),
    .A2(\cpu.keccak_alu.registers[225] ),
    .Y(_05510_),
    .B1(_05509_));
 sg13g2_xor2_1 _12129_ (.B(\cpu.keccak_alu.registers[97] ),
    .A(\cpu.keccak_alu.registers[33] ),
    .X(_05511_));
 sg13g2_a21oi_1 _12130_ (.A1(_05510_),
    .A2(_05511_),
    .Y(_05512_),
    .B1(net4218));
 sg13g2_o21ai_1 _12131_ (.B1(_05512_),
    .Y(_05513_),
    .A1(_05510_),
    .A2(_05511_));
 sg13g2_a21oi_1 _12132_ (.A1(_01002_),
    .A2(net4496),
    .Y(_05514_),
    .B1(net4019));
 sg13g2_nand2b_1 _12133_ (.Y(_05515_),
    .B(_04428_),
    .A_N(_04339_));
 sg13g2_nand3_1 _12134_ (.B(net3828),
    .C(_05515_),
    .A(net4198),
    .Y(_05516_));
 sg13g2_nand3_1 _12135_ (.B(net3828),
    .C(_05459_),
    .A(net4541),
    .Y(_05517_));
 sg13g2_nand2_1 _12136_ (.Y(_05518_),
    .A(_05516_),
    .B(_05517_));
 sg13g2_mux2_1 _12137_ (.A0(_05414_),
    .A1(_05518_),
    .S(net4189),
    .X(_05519_));
 sg13g2_mux2_1 _12138_ (.A0(_05304_),
    .A1(_05519_),
    .S(net4174),
    .X(_05520_));
 sg13g2_o21ai_1 _12139_ (.B1(net4519),
    .Y(_05521_),
    .A1(net4523),
    .A2(_04333_));
 sg13g2_o21ai_1 _12140_ (.B1(_05521_),
    .Y(_05522_),
    .A1(net3935),
    .A2(_05520_));
 sg13g2_o21ai_1 _12141_ (.B1(net4159),
    .Y(_05523_),
    .A1(net4169),
    .A2(_05098_));
 sg13g2_or2_1 _12142_ (.X(_05524_),
    .B(_05523_),
    .A(_05522_));
 sg13g2_nand2_1 _12143_ (.Y(_05525_),
    .A(net3778),
    .B(_04415_));
 sg13g2_xnor2_1 _12144_ (.Y(_05526_),
    .A(_05524_),
    .B(_05525_));
 sg13g2_a21oi_1 _12145_ (.A1(net4019),
    .A2(_05526_),
    .Y(_05527_),
    .B1(_05514_));
 sg13g2_xnor2_1 _12146_ (.Y(_05528_),
    .A(\cpu.keccak_alu.registers[33] ),
    .B(_05527_));
 sg13g2_o21ai_1 _12147_ (.B1(_05513_),
    .Y(_05529_),
    .A1(net4384),
    .A2(_05528_));
 sg13g2_nand2_1 _12148_ (.Y(_05530_),
    .A(net4359),
    .B(_05504_));
 sg13g2_a21oi_1 _12149_ (.A1(_01007_),
    .A2(net3635),
    .Y(_05531_),
    .B1(net3814));
 sg13g2_a221oi_1 _12150_ (.B2(_05531_),
    .C1(net3735),
    .B1(_05530_),
    .A1(net4264),
    .Y(_05532_),
    .A2(_05529_));
 sg13g2_a21oi_1 _12151_ (.A1(_01007_),
    .A2(net3735),
    .Y(_00750_),
    .B1(_05532_));
 sg13g2_o21ai_1 _12152_ (.B1(net4209),
    .Y(_05533_),
    .A1(\cpu.keccak_alu.registers[162] ),
    .A2(\cpu.keccak_alu.registers[226] ));
 sg13g2_a21oi_1 _12153_ (.A1(\cpu.keccak_alu.registers[162] ),
    .A2(\cpu.keccak_alu.registers[226] ),
    .Y(_05534_),
    .B1(_05533_));
 sg13g2_xor2_1 _12154_ (.B(\cpu.keccak_alu.registers[98] ),
    .A(\cpu.keccak_alu.registers[34] ),
    .X(_05535_));
 sg13g2_a21oi_1 _12155_ (.A1(_05534_),
    .A2(_05535_),
    .Y(_05536_),
    .B1(net4218));
 sg13g2_o21ai_1 _12156_ (.B1(_05536_),
    .Y(_05537_),
    .A1(_05534_),
    .A2(_05535_));
 sg13g2_nand2b_1 _12157_ (.Y(_05538_),
    .B(\cpu.keccak_alu.registers[162] ),
    .A_N(\cpu.keccak_alu.registers[98] ));
 sg13g2_nor3_1 _12158_ (.A(net4536),
    .B(_04137_),
    .C(_04140_),
    .Y(_05539_));
 sg13g2_nor3_1 _12159_ (.A(net4195),
    .B(_04139_),
    .C(_04222_),
    .Y(_05540_));
 sg13g2_nor2_1 _12160_ (.A(_05539_),
    .B(_05540_),
    .Y(_05541_));
 sg13g2_nor2_1 _12161_ (.A(net3821),
    .B(_05541_),
    .Y(_05542_));
 sg13g2_mux2_1 _12162_ (.A0(_05434_),
    .A1(_05542_),
    .S(net4181),
    .X(_05543_));
 sg13g2_mux2_1 _12163_ (.A0(_05330_),
    .A1(_05543_),
    .S(net4173),
    .X(_05544_));
 sg13g2_o21ai_1 _12164_ (.B1(net4518),
    .Y(_05545_),
    .A1(net4521),
    .A2(_04534_));
 sg13g2_o21ai_1 _12165_ (.B1(_05545_),
    .Y(_05546_),
    .A1(net3937),
    .A2(_05544_));
 sg13g2_o21ai_1 _12166_ (.B1(net4158),
    .Y(_05547_),
    .A1(net4167),
    .A2(_05124_));
 sg13g2_nor2_1 _12167_ (.A(_05546_),
    .B(_05547_),
    .Y(_05548_));
 sg13g2_nand3_1 _12168_ (.B(_04548_),
    .C(_05548_),
    .A(net3774),
    .Y(_05549_));
 sg13g2_a21o_1 _12169_ (.A2(_04548_),
    .A1(net3774),
    .B1(_05548_),
    .X(_05550_));
 sg13g2_a21oi_2 _12170_ (.B1(net4004),
    .Y(_05551_),
    .A2(_05550_),
    .A1(_05549_));
 sg13g2_a21oi_1 _12171_ (.A1(net4005),
    .A2(_05538_),
    .Y(_05552_),
    .B1(_05551_));
 sg13g2_xnor2_1 _12172_ (.Y(_05553_),
    .A(\cpu.keccak_alu.registers[34] ),
    .B(_05552_));
 sg13g2_o21ai_1 _12173_ (.B1(_05537_),
    .Y(_05554_),
    .A1(net4384),
    .A2(_05553_));
 sg13g2_nand2_1 _12174_ (.Y(_05555_),
    .A(net4355),
    .B(_05504_));
 sg13g2_a21oi_1 _12175_ (.A1(_01015_),
    .A2(net3635),
    .Y(_05556_),
    .B1(net3813));
 sg13g2_a221oi_1 _12176_ (.B2(_05556_),
    .C1(net3736),
    .B1(_05555_),
    .A1(net4264),
    .Y(_05557_),
    .A2(_05554_));
 sg13g2_a21oi_1 _12177_ (.A1(_01015_),
    .A2(net3736),
    .Y(_00751_),
    .B1(_05557_));
 sg13g2_o21ai_1 _12178_ (.B1(net4210),
    .Y(_05558_),
    .A1(\cpu.keccak_alu.registers[163] ),
    .A2(\cpu.keccak_alu.registers[227] ));
 sg13g2_a21oi_1 _12179_ (.A1(\cpu.keccak_alu.registers[163] ),
    .A2(\cpu.keccak_alu.registers[227] ),
    .Y(_05559_),
    .B1(_05558_));
 sg13g2_xor2_1 _12180_ (.B(\cpu.keccak_alu.registers[99] ),
    .A(\cpu.keccak_alu.registers[35] ),
    .X(_05560_));
 sg13g2_o21ai_1 _12181_ (.B1(net4385),
    .Y(_05561_),
    .A1(_05559_),
    .A2(_05560_));
 sg13g2_a21o_1 _12182_ (.A2(_05560_),
    .A1(_05559_),
    .B1(_05561_),
    .X(_05562_));
 sg13g2_o21ai_1 _12183_ (.B1(net4005),
    .Y(_05563_),
    .A1(\cpu.keccak_alu.registers[99] ),
    .A2(_01020_));
 sg13g2_nand2b_1 _12184_ (.Y(_05564_),
    .B(_04340_),
    .A_N(_04335_));
 sg13g2_nand3_1 _12185_ (.B(net3828),
    .C(_05564_),
    .A(net4198),
    .Y(_05565_));
 sg13g2_nand3_1 _12186_ (.B(net3828),
    .C(_05515_),
    .A(net4541),
    .Y(_05566_));
 sg13g2_nand2_1 _12187_ (.Y(_05567_),
    .A(_05565_),
    .B(_05566_));
 sg13g2_mux2_1 _12188_ (.A0(_05462_),
    .A1(_05567_),
    .S(net4187),
    .X(_05568_));
 sg13g2_mux2_1 _12189_ (.A0(_05358_),
    .A1(_05568_),
    .S(net4174),
    .X(_05569_));
 sg13g2_o21ai_1 _12190_ (.B1(net4519),
    .Y(_05570_),
    .A1(net4523),
    .A2(_04596_));
 sg13g2_o21ai_1 _12191_ (.B1(_05570_),
    .Y(_05571_),
    .A1(net3935),
    .A2(_05569_));
 sg13g2_o21ai_1 _12192_ (.B1(net4159),
    .Y(_05572_),
    .A1(net4169),
    .A2(_05152_));
 sg13g2_or2_1 _12193_ (.X(_05573_),
    .B(_05572_),
    .A(_05571_));
 sg13g2_nand3_1 _12194_ (.B(_04603_),
    .C(_04616_),
    .A(net3778),
    .Y(_05574_));
 sg13g2_xor2_1 _12195_ (.B(_05574_),
    .A(_05573_),
    .X(_05575_));
 sg13g2_o21ai_1 _12196_ (.B1(_05563_),
    .Y(_05576_),
    .A1(net4007),
    .A2(_05575_));
 sg13g2_xor2_1 _12197_ (.B(_05576_),
    .A(\cpu.keccak_alu.registers[35] ),
    .X(_05577_));
 sg13g2_o21ai_1 _12198_ (.B1(_05562_),
    .Y(_05578_),
    .A1(net4385),
    .A2(_05577_));
 sg13g2_a22oi_1 _12199_ (.Y(_05579_),
    .B1(net3635),
    .B2(net108),
    .A2(_05082_),
    .A1(_02334_));
 sg13g2_o21ai_1 _12200_ (.B1(net3739),
    .Y(_05580_),
    .A1(net3813),
    .A2(_05579_));
 sg13g2_a21oi_1 _12201_ (.A1(net4265),
    .A2(_05578_),
    .Y(_05581_),
    .B1(_05580_));
 sg13g2_a21oi_1 _12202_ (.A1(_01024_),
    .A2(net3736),
    .Y(_00752_),
    .B1(_05581_));
 sg13g2_a21oi_1 _12203_ (.A1(net4494),
    .A2(\cpu.keccak_alu.registers[228] ),
    .Y(_05582_),
    .B1(net4370));
 sg13g2_o21ai_1 _12204_ (.B1(_05582_),
    .Y(_05583_),
    .A1(net4494),
    .A2(\cpu.keccak_alu.registers[228] ));
 sg13g2_xor2_1 _12205_ (.B(\cpu.keccak_alu.registers[100] ),
    .A(\cpu.keccak_alu.registers[36] ),
    .X(_05584_));
 sg13g2_xnor2_1 _12206_ (.Y(_05585_),
    .A(_05583_),
    .B(_05584_));
 sg13g2_nand3b_1 _12207_ (.B(\cpu.keccak_alu.registers[164] ),
    .C(net4004),
    .Y(_05586_),
    .A_N(\cpu.keccak_alu.registers[100] ));
 sg13g2_and2_1 _12208_ (.A(net4518),
    .B(_04664_),
    .X(_05587_));
 sg13g2_nand2_1 _12209_ (.Y(_05588_),
    .A(net4524),
    .B(net4163));
 sg13g2_nor2_1 _12210_ (.A(_05177_),
    .B(net3873),
    .Y(_05589_));
 sg13g2_nor3_1 _12211_ (.A(net4536),
    .B(_04138_),
    .C(_04150_),
    .Y(_05590_));
 sg13g2_nor3_1 _12212_ (.A(net4195),
    .B(_04137_),
    .C(_04140_),
    .Y(_05591_));
 sg13g2_nor2_1 _12213_ (.A(_05590_),
    .B(_05591_),
    .Y(_05592_));
 sg13g2_nor2_1 _12214_ (.A(net3821),
    .B(_05592_),
    .Y(_05593_));
 sg13g2_mux2_1 _12215_ (.A0(_05492_),
    .A1(_05593_),
    .S(net4181),
    .X(_05594_));
 sg13g2_mux2_1 _12216_ (.A0(_05385_),
    .A1(_05594_),
    .S(net4173),
    .X(_05595_));
 sg13g2_nor2_1 _12217_ (.A(net3934),
    .B(_05595_),
    .Y(_05596_));
 sg13g2_nor4_1 _12218_ (.A(net4513),
    .B(_05587_),
    .C(_05589_),
    .D(_05596_),
    .Y(_05597_));
 sg13g2_nand3_1 _12219_ (.B(_04674_),
    .C(_05597_),
    .A(net3774),
    .Y(_05598_));
 sg13g2_a21oi_1 _12220_ (.A1(net3774),
    .A2(_04674_),
    .Y(_05599_),
    .B1(_05597_));
 sg13g2_nand2_1 _12221_ (.Y(_05600_),
    .A(net4016),
    .B(_05598_));
 sg13g2_o21ai_1 _12222_ (.B1(_05586_),
    .Y(_05601_),
    .A1(_05599_),
    .A2(_05600_));
 sg13g2_or2_1 _12223_ (.X(_05602_),
    .B(_05601_),
    .A(\cpu.keccak_alu.registers[36] ));
 sg13g2_a21oi_1 _12224_ (.A1(\cpu.keccak_alu.registers[36] ),
    .A2(_05601_),
    .Y(_05603_),
    .B1(net4387));
 sg13g2_a22oi_1 _12225_ (.Y(_05604_),
    .B1(_05602_),
    .B2(_05603_),
    .A2(_05585_),
    .A1(net4387));
 sg13g2_or2_1 _12226_ (.X(_05605_),
    .B(_05604_),
    .A(net4319));
 sg13g2_a22oi_1 _12227_ (.Y(_05606_),
    .B1(net3635),
    .B2(net390),
    .A2(net3771),
    .A1(_02336_));
 sg13g2_nor2_1 _12228_ (.A(net3814),
    .B(_05606_),
    .Y(_05607_));
 sg13g2_nor2_1 _12229_ (.A(net3732),
    .B(_05607_),
    .Y(_05608_));
 sg13g2_a22oi_1 _12230_ (.Y(_00753_),
    .B1(_05605_),
    .B2(_05608_),
    .A2(net3732),
    .A1(_01032_));
 sg13g2_a21oi_1 _12231_ (.A1(\cpu.keccak_alu.registers[165] ),
    .A2(\cpu.keccak_alu.registers[229] ),
    .Y(_05609_),
    .B1(net4369));
 sg13g2_o21ai_1 _12232_ (.B1(_05609_),
    .Y(_05610_),
    .A1(\cpu.keccak_alu.registers[165] ),
    .A2(\cpu.keccak_alu.registers[229] ));
 sg13g2_xnor2_1 _12233_ (.Y(_05611_),
    .A(\cpu.keccak_alu.registers[37] ),
    .B(\cpu.keccak_alu.registers[101] ));
 sg13g2_a21oi_1 _12234_ (.A1(_05610_),
    .A2(_05611_),
    .Y(_05612_),
    .B1(net4216));
 sg13g2_o21ai_1 _12235_ (.B1(_05612_),
    .Y(_05613_),
    .A1(_05610_),
    .A2(_05611_));
 sg13g2_a21oi_1 _12236_ (.A1(_01034_),
    .A2(net4493),
    .Y(_05614_),
    .B1(net4017));
 sg13g2_o21ai_1 _12237_ (.B1(_04336_),
    .Y(_05615_),
    .A1(net4562),
    .A2(_00103_));
 sg13g2_nand3_1 _12238_ (.B(net3829),
    .C(_05615_),
    .A(net4197),
    .Y(_05616_));
 sg13g2_nand3_1 _12239_ (.B(net3828),
    .C(_05564_),
    .A(net4542),
    .Y(_05617_));
 sg13g2_nand2_1 _12240_ (.Y(_05618_),
    .A(_05616_),
    .B(_05617_));
 sg13g2_mux2_1 _12241_ (.A0(_05518_),
    .A1(_05618_),
    .S(net4189),
    .X(_05619_));
 sg13g2_mux2_1 _12242_ (.A0(_05415_),
    .A1(_05619_),
    .S(net4175),
    .X(_05620_));
 sg13g2_nor2_1 _12243_ (.A(net3935),
    .B(_05620_),
    .Y(_05621_));
 sg13g2_nor2_1 _12244_ (.A(_05198_),
    .B(net3875),
    .Y(_05622_));
 sg13g2_o21ai_1 _12245_ (.B1(net4159),
    .Y(_05623_),
    .A1(net4163),
    .A2(_04705_));
 sg13g2_nor3_1 _12246_ (.A(_05621_),
    .B(_05622_),
    .C(_05623_),
    .Y(_05624_));
 sg13g2_nand2_1 _12247_ (.Y(_05625_),
    .A(net3776),
    .B(_04720_));
 sg13g2_xor2_1 _12248_ (.B(_05625_),
    .A(_05624_),
    .X(_05626_));
 sg13g2_a21oi_2 _12249_ (.B1(_05614_),
    .Y(_05627_),
    .A2(_05626_),
    .A1(net4017));
 sg13g2_xnor2_1 _12250_ (.Y(_05628_),
    .A(\cpu.keccak_alu.registers[37] ),
    .B(_05627_));
 sg13g2_o21ai_1 _12251_ (.B1(_05613_),
    .Y(_05629_),
    .A1(net4382),
    .A2(_05628_));
 sg13g2_a22oi_1 _12252_ (.Y(_05630_),
    .B1(net3635),
    .B2(net218),
    .A2(net3771),
    .A1(_02338_));
 sg13g2_o21ai_1 _12253_ (.B1(net3738),
    .Y(_05631_),
    .A1(net3812),
    .A2(_05630_));
 sg13g2_a21oi_1 _12254_ (.A1(net4263),
    .A2(_05629_),
    .Y(_05632_),
    .B1(_05631_));
 sg13g2_a21oi_1 _12255_ (.A1(_01040_),
    .A2(net3730),
    .Y(_00754_),
    .B1(_05632_));
 sg13g2_o21ai_1 _12256_ (.B1(net4211),
    .Y(_05633_),
    .A1(\cpu.keccak_alu.registers[166] ),
    .A2(\cpu.keccak_alu.registers[230] ));
 sg13g2_a21oi_1 _12257_ (.A1(\cpu.keccak_alu.registers[166] ),
    .A2(\cpu.keccak_alu.registers[230] ),
    .Y(_05634_),
    .B1(_05633_));
 sg13g2_xor2_1 _12258_ (.B(\cpu.keccak_alu.registers[102] ),
    .A(\cpu.keccak_alu.registers[38] ),
    .X(_05635_));
 sg13g2_a21oi_1 _12259_ (.A1(_05634_),
    .A2(_05635_),
    .Y(_05636_),
    .B1(net4220));
 sg13g2_o21ai_1 _12260_ (.B1(_05636_),
    .Y(_05637_),
    .A1(_05634_),
    .A2(_05635_));
 sg13g2_a21oi_1 _12261_ (.A1(net4518),
    .A2(_04737_),
    .Y(_05638_),
    .B1(net4514));
 sg13g2_nor2_1 _12262_ (.A(_05229_),
    .B(net3872),
    .Y(_05639_));
 sg13g2_nor3_1 _12263_ (.A(net4536),
    .B(_04147_),
    .C(_04151_),
    .Y(_05640_));
 sg13g2_nor3_1 _12264_ (.A(net4193),
    .B(_04138_),
    .C(_04150_),
    .Y(_05641_));
 sg13g2_nor2_1 _12265_ (.A(_05640_),
    .B(_05641_),
    .Y(_05642_));
 sg13g2_nor2_1 _12266_ (.A(net3822),
    .B(_05642_),
    .Y(_05643_));
 sg13g2_mux2_1 _12267_ (.A0(_05542_),
    .A1(_05643_),
    .S(net4181),
    .X(_05644_));
 sg13g2_mux2_1 _12268_ (.A0(_05435_),
    .A1(_05644_),
    .S(net4172),
    .X(_05645_));
 sg13g2_o21ai_1 _12269_ (.B1(_05638_),
    .Y(_05646_),
    .A1(net3934),
    .A2(_05645_));
 sg13g2_or2_1 _12270_ (.X(_05647_),
    .B(_05646_),
    .A(_05639_));
 sg13g2_nand2_1 _12271_ (.Y(_05648_),
    .A(net3773),
    .B(_04752_));
 sg13g2_a21oi_1 _12272_ (.A1(_01044_),
    .A2(\cpu.keccak_alu.registers[166] ),
    .Y(_05649_),
    .B1(net4016));
 sg13g2_xnor2_1 _12273_ (.Y(_05650_),
    .A(_05647_),
    .B(_05648_));
 sg13g2_a21oi_1 _12274_ (.A1(net4016),
    .A2(_05650_),
    .Y(_05651_),
    .B1(_05649_));
 sg13g2_xnor2_1 _12275_ (.Y(_05652_),
    .A(\cpu.keccak_alu.registers[38] ),
    .B(_05651_));
 sg13g2_o21ai_1 _12276_ (.B1(_05637_),
    .Y(_05653_),
    .A1(net4382),
    .A2(_05652_));
 sg13g2_a22oi_1 _12277_ (.Y(_05654_),
    .B1(net3635),
    .B2(net167),
    .A2(_05082_),
    .A1(_02340_));
 sg13g2_o21ai_1 _12278_ (.B1(net3739),
    .Y(_05655_),
    .A1(net3814),
    .A2(_05654_));
 sg13g2_a21oi_1 _12279_ (.A1(net4263),
    .A2(_05653_),
    .Y(_05656_),
    .B1(_05655_));
 sg13g2_a21oi_1 _12280_ (.A1(_01050_),
    .A2(net3730),
    .Y(_00755_),
    .B1(_05656_));
 sg13g2_a21oi_1 _12281_ (.A1(_01053_),
    .A2(\cpu.keccak_alu.registers[167] ),
    .Y(_05657_),
    .B1(net4015));
 sg13g2_a21oi_1 _12282_ (.A1(net4523),
    .A2(_05255_),
    .Y(_05658_),
    .B1(net4519));
 sg13g2_nand2b_1 _12283_ (.Y(_05659_),
    .B(_04349_),
    .A_N(_04344_));
 sg13g2_nand3_1 _12284_ (.B(net3829),
    .C(_05659_),
    .A(net4197),
    .Y(_05660_));
 sg13g2_nand3_1 _12285_ (.B(net3829),
    .C(_05615_),
    .A(net4542),
    .Y(_05661_));
 sg13g2_nand2_1 _12286_ (.Y(_05662_),
    .A(_05660_),
    .B(_05661_));
 sg13g2_mux2_1 _12287_ (.A0(_05567_),
    .A1(_05662_),
    .S(net4185),
    .X(_05663_));
 sg13g2_mux2_1 _12288_ (.A0(_05463_),
    .A1(_05663_),
    .S(net4174),
    .X(_05664_));
 sg13g2_nor2_1 _12289_ (.A(net3935),
    .B(_05664_),
    .Y(_05665_));
 sg13g2_nor2_1 _12290_ (.A(net4515),
    .B(_05665_),
    .Y(_05666_));
 sg13g2_o21ai_1 _12291_ (.B1(_05666_),
    .Y(_05667_),
    .A1(_04776_),
    .A2(_05658_));
 sg13g2_nand2_1 _12292_ (.Y(_05668_),
    .A(net3777),
    .B(_04792_));
 sg13g2_xnor2_1 _12293_ (.Y(_05669_),
    .A(_05667_),
    .B(_05668_));
 sg13g2_a21oi_1 _12294_ (.A1(net4015),
    .A2(_05669_),
    .Y(_05670_),
    .B1(_05657_));
 sg13g2_or2_1 _12295_ (.X(_05671_),
    .B(_05670_),
    .A(\cpu.keccak_alu.registers[39] ));
 sg13g2_a21oi_1 _12296_ (.A1(\cpu.keccak_alu.registers[39] ),
    .A2(_05670_),
    .Y(_05672_),
    .B1(net4377));
 sg13g2_a21oi_1 _12297_ (.A1(\cpu.keccak_alu.registers[167] ),
    .A2(\cpu.keccak_alu.registers[231] ),
    .Y(_05673_),
    .B1(net4369));
 sg13g2_o21ai_1 _12298_ (.B1(_05673_),
    .Y(_05674_),
    .A1(\cpu.keccak_alu.registers[167] ),
    .A2(\cpu.keccak_alu.registers[231] ));
 sg13g2_xor2_1 _12299_ (.B(\cpu.keccak_alu.registers[103] ),
    .A(\cpu.keccak_alu.registers[39] ),
    .X(_05675_));
 sg13g2_xnor2_1 _12300_ (.Y(_05676_),
    .A(_05674_),
    .B(_05675_));
 sg13g2_a22oi_1 _12301_ (.Y(_05677_),
    .B1(_05676_),
    .B2(net4377),
    .A2(_05672_),
    .A1(_05671_));
 sg13g2_or2_1 _12302_ (.X(_05678_),
    .B(_05677_),
    .A(net4315));
 sg13g2_a22oi_1 _12303_ (.Y(_05679_),
    .B1(net3635),
    .B2(net276),
    .A2(net3771),
    .A1(_02342_));
 sg13g2_nor2_1 _12304_ (.A(net3812),
    .B(_05679_),
    .Y(_05680_));
 sg13g2_nor2_1 _12305_ (.A(net3727),
    .B(_05680_),
    .Y(_05681_));
 sg13g2_a22oi_1 _12306_ (.Y(_00756_),
    .B1(_05678_),
    .B2(_05681_),
    .A2(net3727),
    .A1(_01059_));
 sg13g2_a21oi_1 _12307_ (.A1(\cpu.keccak_alu.registers[168] ),
    .A2(\cpu.keccak_alu.registers[232] ),
    .Y(_05682_),
    .B1(net4369));
 sg13g2_o21ai_1 _12308_ (.B1(_05682_),
    .Y(_05683_),
    .A1(\cpu.keccak_alu.registers[168] ),
    .A2(\cpu.keccak_alu.registers[232] ));
 sg13g2_xnor2_1 _12309_ (.Y(_05684_),
    .A(\cpu.keccak_alu.registers[40] ),
    .B(\cpu.keccak_alu.registers[104] ));
 sg13g2_a21oi_1 _12310_ (.A1(_05683_),
    .A2(_05684_),
    .Y(_05685_),
    .B1(net4216));
 sg13g2_o21ai_1 _12311_ (.B1(_05685_),
    .Y(_05686_),
    .A1(_05683_),
    .A2(_05684_));
 sg13g2_nand3b_1 _12312_ (.B(\cpu.keccak_alu.registers[168] ),
    .C(net4001),
    .Y(_05687_),
    .A_N(\cpu.keccak_alu.registers[104] ));
 sg13g2_a21oi_1 _12313_ (.A1(net4164),
    .A2(_04817_),
    .Y(_05688_),
    .B1(net4161));
 sg13g2_o21ai_1 _12314_ (.B1(net4157),
    .Y(_05689_),
    .A1(_05283_),
    .A2(net3871));
 sg13g2_nor3_1 _12315_ (.A(net4193),
    .B(_04147_),
    .C(_04151_),
    .Y(_05690_));
 sg13g2_nor3_1 _12316_ (.A(net4535),
    .B(_04053_),
    .C(_04148_),
    .Y(_05691_));
 sg13g2_nor2_1 _12317_ (.A(_05690_),
    .B(_05691_),
    .Y(_05692_));
 sg13g2_nor2_1 _12318_ (.A(net3821),
    .B(_05692_),
    .Y(_05693_));
 sg13g2_mux2_1 _12319_ (.A0(_05593_),
    .A1(_05693_),
    .S(net4181),
    .X(_05694_));
 sg13g2_mux2_1 _12320_ (.A0(_05493_),
    .A1(_05694_),
    .S(net4171),
    .X(_05695_));
 sg13g2_nor2_1 _12321_ (.A(net3934),
    .B(_05695_),
    .Y(_05696_));
 sg13g2_nor3_1 _12322_ (.A(_05688_),
    .B(_05689_),
    .C(_05696_),
    .Y(_05697_));
 sg13g2_nand2_1 _12323_ (.Y(_05698_),
    .A(net3772),
    .B(_04821_));
 sg13g2_xor2_1 _12324_ (.B(_05698_),
    .A(_05697_),
    .X(_05699_));
 sg13g2_o21ai_1 _12325_ (.B1(_05687_),
    .Y(_05700_),
    .A1(net4001),
    .A2(_05699_));
 sg13g2_xnor2_1 _12326_ (.Y(_05701_),
    .A(\cpu.keccak_alu.registers[40] ),
    .B(_05700_));
 sg13g2_o21ai_1 _12327_ (.B1(_05686_),
    .Y(_05702_),
    .A1(net4379),
    .A2(_05701_));
 sg13g2_a22oi_1 _12328_ (.Y(_05703_),
    .B1(net3634),
    .B2(net125),
    .A2(net3770),
    .A1(_02344_));
 sg13g2_o21ai_1 _12329_ (.B1(net3738),
    .Y(_05704_),
    .A1(net3811),
    .A2(_05703_));
 sg13g2_a21oi_1 _12330_ (.A1(net4258),
    .A2(_05702_),
    .Y(_05705_),
    .B1(_05704_));
 sg13g2_a21oi_1 _12331_ (.A1(_01068_),
    .A2(net3723),
    .Y(_00757_),
    .B1(_05705_));
 sg13g2_o21ai_1 _12332_ (.B1(net4206),
    .Y(_05706_),
    .A1(\cpu.keccak_alu.registers[169] ),
    .A2(\cpu.keccak_alu.registers[233] ));
 sg13g2_a21oi_1 _12333_ (.A1(\cpu.keccak_alu.registers[169] ),
    .A2(\cpu.keccak_alu.registers[233] ),
    .Y(_05707_),
    .B1(_05706_));
 sg13g2_xor2_1 _12334_ (.B(\cpu.keccak_alu.registers[105] ),
    .A(\cpu.keccak_alu.registers[41] ),
    .X(_05708_));
 sg13g2_o21ai_1 _12335_ (.B1(net4372),
    .Y(_05709_),
    .A1(_05707_),
    .A2(_05708_));
 sg13g2_a21o_1 _12336_ (.A2(_05708_),
    .A1(_05707_),
    .B1(_05709_),
    .X(_05710_));
 sg13g2_nand3b_1 _12337_ (.B(\cpu.keccak_alu.registers[169] ),
    .C(net4000),
    .Y(_05711_),
    .A_N(\cpu.keccak_alu.registers[105] ));
 sg13g2_nor2_1 _12338_ (.A(_05305_),
    .B(net3874),
    .Y(_05712_));
 sg13g2_o21ai_1 _12339_ (.B1(_04345_),
    .Y(_05713_),
    .A1(net4554),
    .A2(_00107_));
 sg13g2_nand3_1 _12340_ (.B(net3829),
    .C(_05713_),
    .A(net4197),
    .Y(_05714_));
 sg13g2_nand3_1 _12341_ (.B(net3829),
    .C(_05659_),
    .A(net4542),
    .Y(_05715_));
 sg13g2_nand2_1 _12342_ (.Y(_05716_),
    .A(_05714_),
    .B(_05715_));
 sg13g2_mux2_1 _12343_ (.A0(_05618_),
    .A1(_05716_),
    .S(net4185),
    .X(_05717_));
 sg13g2_mux2_1 _12344_ (.A0(_05519_),
    .A1(_05717_),
    .S(net4174),
    .X(_05718_));
 sg13g2_o21ai_1 _12345_ (.B1(net4159),
    .Y(_05719_),
    .A1(net3935),
    .A2(_05718_));
 sg13g2_nor2_1 _12346_ (.A(_05712_),
    .B(_05719_),
    .Y(_05720_));
 sg13g2_o21ai_1 _12347_ (.B1(_05720_),
    .Y(_05721_),
    .A1(net4163),
    .A2(_04846_));
 sg13g2_nand2_1 _12348_ (.Y(_05722_),
    .A(net3777),
    .B(_04855_));
 sg13g2_xnor2_1 _12349_ (.Y(_05723_),
    .A(_05721_),
    .B(_05722_));
 sg13g2_o21ai_1 _12350_ (.B1(_05711_),
    .Y(_05724_),
    .A1(net4000),
    .A2(_05723_));
 sg13g2_xnor2_1 _12351_ (.Y(_05725_),
    .A(\cpu.keccak_alu.registers[41] ),
    .B(_05724_));
 sg13g2_o21ai_1 _12352_ (.B1(_05710_),
    .Y(_05726_),
    .A1(net4372),
    .A2(_05725_));
 sg13g2_a22oi_1 _12353_ (.Y(_05727_),
    .B1(net3634),
    .B2(net209),
    .A2(net3770),
    .A1(_02346_));
 sg13g2_o21ai_1 _12354_ (.B1(net3738),
    .Y(_05728_),
    .A1(net3811),
    .A2(_05727_));
 sg13g2_a21oi_1 _12355_ (.A1(net4245),
    .A2(_05726_),
    .Y(_05729_),
    .B1(_05728_));
 sg13g2_a21oi_1 _12356_ (.A1(_01076_),
    .A2(net3723),
    .Y(_00758_),
    .B1(_05729_));
 sg13g2_o21ai_1 _12357_ (.B1(net4206),
    .Y(_05730_),
    .A1(net4492),
    .A2(\cpu.keccak_alu.registers[234] ));
 sg13g2_a21oi_1 _12358_ (.A1(net4492),
    .A2(\cpu.keccak_alu.registers[234] ),
    .Y(_05731_),
    .B1(_05730_));
 sg13g2_xor2_1 _12359_ (.B(\cpu.keccak_alu.registers[106] ),
    .A(\cpu.keccak_alu.registers[42] ),
    .X(_05732_));
 sg13g2_a21oi_1 _12360_ (.A1(_05731_),
    .A2(_05732_),
    .Y(_05733_),
    .B1(net4213));
 sg13g2_o21ai_1 _12361_ (.B1(_05733_),
    .Y(_05734_),
    .A1(_05731_),
    .A2(_05732_));
 sg13g2_nor3_1 _12362_ (.A(net4191),
    .B(_04053_),
    .C(_04148_),
    .Y(_05735_));
 sg13g2_nor3_1 _12363_ (.A(net4536),
    .B(_04050_),
    .C(_04054_),
    .Y(_05736_));
 sg13g2_nor2_1 _12364_ (.A(_05735_),
    .B(_05736_),
    .Y(_05737_));
 sg13g2_nor2_1 _12365_ (.A(net3821),
    .B(_05737_),
    .Y(_05738_));
 sg13g2_mux2_1 _12366_ (.A0(_05643_),
    .A1(_05738_),
    .S(net4180),
    .X(_05739_));
 sg13g2_mux2_1 _12367_ (.A0(_05543_),
    .A1(_05739_),
    .S(net4172),
    .X(_05740_));
 sg13g2_nor2_1 _12368_ (.A(net3934),
    .B(_05740_),
    .Y(_05741_));
 sg13g2_nor2_1 _12369_ (.A(net4513),
    .B(_05741_),
    .Y(_05742_));
 sg13g2_o21ai_1 _12370_ (.B1(_05742_),
    .Y(_05743_),
    .A1(_05331_),
    .A2(net3871));
 sg13g2_a21oi_1 _12371_ (.A1(net4517),
    .A2(_04879_),
    .Y(_05744_),
    .B1(_05743_));
 sg13g2_nand2_1 _12372_ (.Y(_05745_),
    .A(net3773),
    .B(_04883_));
 sg13g2_a21oi_1 _12373_ (.A1(_01080_),
    .A2(net4492),
    .Y(_05746_),
    .B1(net4010));
 sg13g2_xor2_1 _12374_ (.B(_05745_),
    .A(_05744_),
    .X(_05747_));
 sg13g2_a21oi_1 _12375_ (.A1(net4010),
    .A2(_05747_),
    .Y(_05748_),
    .B1(_05746_));
 sg13g2_xnor2_1 _12376_ (.Y(_05749_),
    .A(\cpu.keccak_alu.registers[42] ),
    .B(_05748_));
 sg13g2_o21ai_1 _12377_ (.B1(_05734_),
    .Y(_05750_),
    .A1(net4372),
    .A2(_05749_));
 sg13g2_a22oi_1 _12378_ (.Y(_05751_),
    .B1(net3634),
    .B2(net129),
    .A2(net3770),
    .A1(_02348_));
 sg13g2_o21ai_1 _12379_ (.B1(net3738),
    .Y(_05752_),
    .A1(net3811),
    .A2(_05751_));
 sg13g2_a21oi_1 _12380_ (.A1(net4245),
    .A2(_05750_),
    .Y(_05753_),
    .B1(_05752_));
 sg13g2_a21oi_1 _12381_ (.A1(_01083_),
    .A2(net3721),
    .Y(_00759_),
    .B1(_05753_));
 sg13g2_o21ai_1 _12382_ (.B1(net4206),
    .Y(_05754_),
    .A1(net4490),
    .A2(\cpu.keccak_alu.registers[235] ));
 sg13g2_a21oi_1 _12383_ (.A1(net4490),
    .A2(\cpu.keccak_alu.registers[235] ),
    .Y(_05755_),
    .B1(_05754_));
 sg13g2_xor2_1 _12384_ (.B(\cpu.keccak_alu.registers[107] ),
    .A(\cpu.keccak_alu.registers[43] ),
    .X(_05756_));
 sg13g2_a21oi_1 _12385_ (.A1(_05755_),
    .A2(_05756_),
    .Y(_05757_),
    .B1(net4214));
 sg13g2_o21ai_1 _12386_ (.B1(_05757_),
    .Y(_05758_),
    .A1(_05755_),
    .A2(_05756_));
 sg13g2_a21oi_1 _12387_ (.A1(net4168),
    .A2(_04905_),
    .Y(_05759_),
    .B1(net4163));
 sg13g2_nor2_1 _12388_ (.A(_05359_),
    .B(net3874),
    .Y(_05760_));
 sg13g2_o21ai_1 _12389_ (.B1(net3827),
    .Y(_05761_),
    .A1(_04354_),
    .A2(_04358_));
 sg13g2_nand3_1 _12390_ (.B(net3829),
    .C(_05713_),
    .A(net4542),
    .Y(_05762_));
 sg13g2_o21ai_1 _12391_ (.B1(_05762_),
    .Y(_05763_),
    .A1(net4542),
    .A2(_05761_));
 sg13g2_mux2_1 _12392_ (.A0(_05662_),
    .A1(_05763_),
    .S(net4185),
    .X(_05764_));
 sg13g2_mux2_1 _12393_ (.A0(_05568_),
    .A1(_05764_),
    .S(net4174),
    .X(_05765_));
 sg13g2_o21ai_1 _12394_ (.B1(net4159),
    .Y(_05766_),
    .A1(net3935),
    .A2(_05765_));
 sg13g2_nor3_2 _12395_ (.A(_05759_),
    .B(_05760_),
    .C(_05766_),
    .Y(_05767_));
 sg13g2_nand3_1 _12396_ (.B(_04913_),
    .C(_04914_),
    .A(net3779),
    .Y(_05768_));
 sg13g2_a21oi_1 _12397_ (.A1(_01087_),
    .A2(net4490),
    .Y(_05769_),
    .B1(net4011));
 sg13g2_xor2_1 _12398_ (.B(_05768_),
    .A(_05767_),
    .X(_05770_));
 sg13g2_a21oi_1 _12399_ (.A1(net4011),
    .A2(_05770_),
    .Y(_05771_),
    .B1(_05769_));
 sg13g2_xnor2_1 _12400_ (.Y(_05772_),
    .A(\cpu.keccak_alu.registers[43] ),
    .B(_05771_));
 sg13g2_o21ai_1 _12401_ (.B1(_05758_),
    .Y(_05773_),
    .A1(net4374),
    .A2(_05772_));
 sg13g2_a22oi_1 _12402_ (.Y(_05774_),
    .B1(net3634),
    .B2(net144),
    .A2(net3770),
    .A1(_02350_));
 sg13g2_o21ai_1 _12403_ (.B1(net3738),
    .Y(_05775_),
    .A1(net3811),
    .A2(_05774_));
 sg13g2_a21oi_1 _12404_ (.A1(net4244),
    .A2(_05773_),
    .Y(_05776_),
    .B1(_05775_));
 sg13g2_a21oi_1 _12405_ (.A1(_01092_),
    .A2(net3723),
    .Y(_00760_),
    .B1(_05776_));
 sg13g2_nand3b_1 _12406_ (.B(net4489),
    .C(net4003),
    .Y(_05777_),
    .A_N(\cpu.keccak_alu.registers[108] ));
 sg13g2_nand2_2 _12407_ (.Y(_05778_),
    .A(net4172),
    .B(net3827));
 sg13g2_or2_1 _12408_ (.X(_05779_),
    .B(_04116_),
    .A(_04051_));
 sg13g2_nor2_1 _12409_ (.A(net4536),
    .B(_05779_),
    .Y(_05780_));
 sg13g2_nor3_1 _12410_ (.A(net4191),
    .B(_04050_),
    .C(_04054_),
    .Y(_05781_));
 sg13g2_nor2_1 _12411_ (.A(_05780_),
    .B(_05781_),
    .Y(_05782_));
 sg13g2_nor3_1 _12412_ (.A(net4531),
    .B(net3821),
    .C(_05782_),
    .Y(_05783_));
 sg13g2_a21o_1 _12413_ (.A2(_05693_),
    .A1(net4531),
    .B1(_05783_),
    .X(_05784_));
 sg13g2_mux2_1 _12414_ (.A0(_05594_),
    .A1(_05784_),
    .S(net4171),
    .X(_05785_));
 sg13g2_o21ai_1 _12415_ (.B1(net4157),
    .Y(_05786_),
    .A1(net3934),
    .A2(_05785_));
 sg13g2_a21oi_1 _12416_ (.A1(net4517),
    .A2(_04938_),
    .Y(_05787_),
    .B1(_05786_));
 sg13g2_o21ai_1 _12417_ (.B1(_05787_),
    .Y(_05788_),
    .A1(_05386_),
    .A2(net3871));
 sg13g2_nand2_1 _12418_ (.Y(_05789_),
    .A(net3772),
    .B(_04943_));
 sg13g2_xnor2_1 _12419_ (.Y(_05790_),
    .A(_05788_),
    .B(_05789_));
 sg13g2_o21ai_1 _12420_ (.B1(_05777_),
    .Y(_05791_),
    .A1(net4003),
    .A2(_05790_));
 sg13g2_or2_1 _12421_ (.X(_05792_),
    .B(_05791_),
    .A(\cpu.keccak_alu.registers[44] ));
 sg13g2_a21oi_1 _12422_ (.A1(\cpu.keccak_alu.registers[44] ),
    .A2(_05791_),
    .Y(_05793_),
    .B1(net4377));
 sg13g2_a21oi_1 _12423_ (.A1(net4489),
    .A2(\cpu.keccak_alu.registers[236] ),
    .Y(_05794_),
    .B1(net4369));
 sg13g2_o21ai_1 _12424_ (.B1(_05794_),
    .Y(_05795_),
    .A1(net4489),
    .A2(\cpu.keccak_alu.registers[236] ));
 sg13g2_xor2_1 _12425_ (.B(\cpu.keccak_alu.registers[108] ),
    .A(\cpu.keccak_alu.registers[44] ),
    .X(_05796_));
 sg13g2_xnor2_1 _12426_ (.Y(_05797_),
    .A(_05795_),
    .B(_05796_));
 sg13g2_a22oi_1 _12427_ (.Y(_05798_),
    .B1(_05797_),
    .B2(net4377),
    .A2(_05793_),
    .A1(_05792_));
 sg13g2_or2_1 _12428_ (.X(_05799_),
    .B(_05798_),
    .A(net4315));
 sg13g2_a22oi_1 _12429_ (.Y(_05800_),
    .B1(net3634),
    .B2(\cpu.keccak_alu.registers[300] ),
    .A2(_05082_),
    .A1(_02352_));
 sg13g2_nor2_1 _12430_ (.A(net3812),
    .B(_05800_),
    .Y(_05801_));
 sg13g2_nor2_1 _12431_ (.A(net3727),
    .B(_05801_),
    .Y(_05802_));
 sg13g2_a22oi_1 _12432_ (.Y(_00761_),
    .B1(_05799_),
    .B2(_05802_),
    .A2(net3727),
    .A1(_01101_));
 sg13g2_nor2b_1 _12433_ (.A(\cpu.keccak_alu.registers[109] ),
    .B_N(net4488),
    .Y(_05803_));
 sg13g2_nor2_1 _12434_ (.A(_05416_),
    .B(net3875),
    .Y(_05804_));
 sg13g2_nor2_1 _12435_ (.A(net4515),
    .B(_05804_),
    .Y(_05805_));
 sg13g2_o21ai_1 _12436_ (.B1(net3827),
    .Y(_05806_),
    .A1(_04355_),
    .A2(_04368_));
 sg13g2_nand2b_1 _12437_ (.Y(_05807_),
    .B(net4197),
    .A_N(_05806_));
 sg13g2_o21ai_1 _12438_ (.B1(_05807_),
    .Y(_05808_),
    .A1(net4197),
    .A2(_05761_));
 sg13g2_mux2_1 _12439_ (.A0(_05716_),
    .A1(_05808_),
    .S(net4185),
    .X(_05809_));
 sg13g2_mux2_1 _12440_ (.A0(_05619_),
    .A1(_05809_),
    .S(net4175),
    .X(_05810_));
 sg13g2_o21ai_1 _12441_ (.B1(_05805_),
    .Y(_05811_),
    .A1(net3935),
    .A2(_05810_));
 sg13g2_a21oi_1 _12442_ (.A1(net4520),
    .A2(_04977_),
    .Y(_05812_),
    .B1(_05811_));
 sg13g2_nand2_1 _12443_ (.Y(_05813_),
    .A(net3778),
    .B(_04986_));
 sg13g2_xnor2_1 _12444_ (.Y(_05814_),
    .A(_05812_),
    .B(_05813_));
 sg13g2_mux2_1 _12445_ (.A0(_05803_),
    .A1(_05814_),
    .S(net4012),
    .X(_05815_));
 sg13g2_o21ai_1 _12446_ (.B1(net4215),
    .Y(_05816_),
    .A1(\cpu.keccak_alu.registers[45] ),
    .A2(_05815_));
 sg13g2_a21oi_1 _12447_ (.A1(\cpu.keccak_alu.registers[45] ),
    .A2(_05815_),
    .Y(_05817_),
    .B1(_05816_));
 sg13g2_a21oi_1 _12448_ (.A1(net4488),
    .A2(\cpu.keccak_alu.registers[237] ),
    .Y(_05818_),
    .B1(net4367));
 sg13g2_o21ai_1 _12449_ (.B1(_05818_),
    .Y(_05819_),
    .A1(net4488),
    .A2(\cpu.keccak_alu.registers[237] ));
 sg13g2_xnor2_1 _12450_ (.Y(_05820_),
    .A(\cpu.keccak_alu.registers[45] ),
    .B(\cpu.keccak_alu.registers[109] ));
 sg13g2_o21ai_1 _12451_ (.B1(net4376),
    .Y(_05821_),
    .A1(_05819_),
    .A2(_05820_));
 sg13g2_a21oi_1 _12452_ (.A1(_05819_),
    .A2(_05820_),
    .Y(_05822_),
    .B1(_05821_));
 sg13g2_o21ai_1 _12453_ (.B1(net4245),
    .Y(_05823_),
    .A1(_05817_),
    .A2(_05822_));
 sg13g2_a22oi_1 _12454_ (.Y(_05824_),
    .B1(net3634),
    .B2(net269),
    .A2(net3770),
    .A1(_02354_));
 sg13g2_nor2_1 _12455_ (.A(net3811),
    .B(_05824_),
    .Y(_05825_));
 sg13g2_nor2_1 _12456_ (.A(net3722),
    .B(_05825_),
    .Y(_05826_));
 sg13g2_a22oi_1 _12457_ (.Y(_00762_),
    .B1(_05823_),
    .B2(_05826_),
    .A2(net3722),
    .A1(_01109_));
 sg13g2_nor2_1 _12458_ (.A(net4161),
    .B(_05006_),
    .Y(_05827_));
 sg13g2_nor2_1 _12459_ (.A(_05436_),
    .B(net3871),
    .Y(_05828_));
 sg13g2_nor2_1 _12460_ (.A(_04113_),
    .B(_04117_),
    .Y(_05829_));
 sg13g2_nor2_1 _12461_ (.A(net4192),
    .B(_05779_),
    .Y(_05830_));
 sg13g2_a21oi_1 _12462_ (.A1(net4192),
    .A2(_05829_),
    .Y(_05831_),
    .B1(_05830_));
 sg13g2_nor3_1 _12463_ (.A(net4531),
    .B(net3821),
    .C(_05831_),
    .Y(_05832_));
 sg13g2_a21o_1 _12464_ (.A2(_05738_),
    .A1(net4531),
    .B1(_05832_),
    .X(_05833_));
 sg13g2_mux2_1 _12465_ (.A0(_05644_),
    .A1(_05833_),
    .S(net4172),
    .X(_05834_));
 sg13g2_o21ai_1 _12466_ (.B1(net4157),
    .Y(_05835_),
    .A1(net3934),
    .A2(_05834_));
 sg13g2_nor3_1 _12467_ (.A(_05827_),
    .B(_05828_),
    .C(_05835_),
    .Y(_05836_));
 sg13g2_nand2_1 _12468_ (.Y(_05837_),
    .A(net3775),
    .B(_05010_));
 sg13g2_a21oi_1 _12469_ (.A1(_01120_),
    .A2(\cpu.keccak_alu.registers[174] ),
    .Y(_05838_),
    .B1(net4011));
 sg13g2_xor2_1 _12470_ (.B(_05837_),
    .A(_05836_),
    .X(_05839_));
 sg13g2_a21oi_1 _12471_ (.A1(net4011),
    .A2(_05839_),
    .Y(_05840_),
    .B1(_05838_));
 sg13g2_xnor2_1 _12472_ (.Y(_05841_),
    .A(\cpu.keccak_alu.registers[46] ),
    .B(_05840_));
 sg13g2_o21ai_1 _12473_ (.B1(net4206),
    .Y(_05842_),
    .A1(\cpu.keccak_alu.registers[174] ),
    .A2(\cpu.keccak_alu.registers[238] ));
 sg13g2_a21oi_1 _12474_ (.A1(\cpu.keccak_alu.registers[174] ),
    .A2(\cpu.keccak_alu.registers[238] ),
    .Y(_05843_),
    .B1(_05842_));
 sg13g2_xor2_1 _12475_ (.B(\cpu.keccak_alu.registers[110] ),
    .A(\cpu.keccak_alu.registers[46] ),
    .X(_05844_));
 sg13g2_a21oi_1 _12476_ (.A1(_05843_),
    .A2(_05844_),
    .Y(_05845_),
    .B1(net4214));
 sg13g2_o21ai_1 _12477_ (.B1(_05845_),
    .Y(_05846_),
    .A1(_05843_),
    .A2(_05844_));
 sg13g2_o21ai_1 _12478_ (.B1(_05846_),
    .Y(_05847_),
    .A1(net4375),
    .A2(_05841_));
 sg13g2_a22oi_1 _12479_ (.Y(_05848_),
    .B1(net3634),
    .B2(net138),
    .A2(net3770),
    .A1(_02356_));
 sg13g2_o21ai_1 _12480_ (.B1(net3738),
    .Y(_05849_),
    .A1(net3811),
    .A2(_05848_));
 sg13g2_a21oi_1 _12481_ (.A1(net4244),
    .A2(_05847_),
    .Y(_05850_),
    .B1(_05849_));
 sg13g2_a21oi_1 _12482_ (.A1(_01124_),
    .A2(net3723),
    .Y(_00763_),
    .B1(_05850_));
 sg13g2_a21oi_1 _12483_ (.A1(_01134_),
    .A2(\cpu.keccak_alu.registers[175] ),
    .Y(_05851_),
    .B1(net4013));
 sg13g2_a21oi_1 _12484_ (.A1(net4168),
    .A2(_05033_),
    .Y(_05852_),
    .B1(net4163));
 sg13g2_nor2_1 _12485_ (.A(_05464_),
    .B(net3874),
    .Y(_05853_));
 sg13g2_o21ai_1 _12486_ (.B1(net3827),
    .Y(_05854_),
    .A1(_04364_),
    .A2(_04369_));
 sg13g2_nand2b_1 _12487_ (.Y(_05855_),
    .B(net4198),
    .A_N(_05854_));
 sg13g2_o21ai_1 _12488_ (.B1(_05855_),
    .Y(_05856_),
    .A1(net4198),
    .A2(_05806_));
 sg13g2_mux2_1 _12489_ (.A0(_05763_),
    .A1(_05856_),
    .S(net4185),
    .X(_05857_));
 sg13g2_mux2_1 _12490_ (.A0(_05663_),
    .A1(_05857_),
    .S(net4175),
    .X(_05858_));
 sg13g2_o21ai_1 _12491_ (.B1(net4160),
    .Y(_05859_),
    .A1(net3935),
    .A2(_05858_));
 sg13g2_nor3_1 _12492_ (.A(_05852_),
    .B(_05853_),
    .C(_05859_),
    .Y(_05860_));
 sg13g2_nand2_1 _12493_ (.Y(_05861_),
    .A(net3778),
    .B(_05041_));
 sg13g2_xor2_1 _12494_ (.B(_05861_),
    .A(_05860_),
    .X(_05862_));
 sg13g2_a21oi_2 _12495_ (.B1(_05851_),
    .Y(_05863_),
    .A2(_05862_),
    .A1(net4013));
 sg13g2_or2_1 _12496_ (.X(_05864_),
    .B(_05863_),
    .A(\cpu.keccak_alu.registers[47] ));
 sg13g2_a21oi_1 _12497_ (.A1(\cpu.keccak_alu.registers[47] ),
    .A2(_05863_),
    .Y(_05865_),
    .B1(net4381));
 sg13g2_a21oi_1 _12498_ (.A1(\cpu.keccak_alu.registers[175] ),
    .A2(\cpu.keccak_alu.registers[239] ),
    .Y(_05866_),
    .B1(net4368));
 sg13g2_o21ai_1 _12499_ (.B1(_05866_),
    .Y(_05867_),
    .A1(\cpu.keccak_alu.registers[175] ),
    .A2(\cpu.keccak_alu.registers[239] ));
 sg13g2_xor2_1 _12500_ (.B(\cpu.keccak_alu.registers[111] ),
    .A(\cpu.keccak_alu.registers[47] ),
    .X(_05868_));
 sg13g2_xnor2_1 _12501_ (.Y(_05869_),
    .A(_05867_),
    .B(_05868_));
 sg13g2_a22oi_1 _12502_ (.Y(_05870_),
    .B1(_05869_),
    .B2(net4376),
    .A2(_05865_),
    .A1(_05864_));
 sg13g2_or2_1 _12503_ (.X(_05871_),
    .B(_05870_),
    .A(net4314));
 sg13g2_a22oi_1 _12504_ (.Y(_05872_),
    .B1(net3634),
    .B2(net296),
    .A2(net3770),
    .A1(_02358_));
 sg13g2_nor2_1 _12505_ (.A(net3811),
    .B(_05872_),
    .Y(_05873_));
 sg13g2_nor2_1 _12506_ (.A(net3724),
    .B(_05873_),
    .Y(_05874_));
 sg13g2_a22oi_1 _12507_ (.Y(_00764_),
    .B1(_05871_),
    .B2(_05874_),
    .A2(net3724),
    .A1(_01137_));
 sg13g2_nand3_1 _12508_ (.B(_04206_),
    .C(net3775),
    .A(net3917),
    .Y(_05875_));
 sg13g2_nand2_1 _12509_ (.Y(_05876_),
    .A(net4525),
    .B(_05694_));
 sg13g2_nor2_1 _12510_ (.A(_04114_),
    .B(_04188_),
    .Y(_05877_));
 sg13g2_nor3_1 _12511_ (.A(net4537),
    .B(_04114_),
    .C(_04188_),
    .Y(_05878_));
 sg13g2_a21oi_1 _12512_ (.A1(net4537),
    .A2(_05829_),
    .Y(_05879_),
    .B1(_05878_));
 sg13g2_mux2_1 _12513_ (.A0(_05782_),
    .A1(_05879_),
    .S(net4180),
    .X(_05880_));
 sg13g2_nor2_2 _12514_ (.A(net3821),
    .B(_05880_),
    .Y(_05881_));
 sg13g2_a21oi_1 _12515_ (.A1(net4171),
    .A2(_05881_),
    .Y(_05882_),
    .B1(net3934));
 sg13g2_nor2_1 _12516_ (.A(_05494_),
    .B(net3873),
    .Y(_05883_));
 sg13g2_a221oi_1 _12517_ (.B2(_05882_),
    .C1(_05883_),
    .B1(_05876_),
    .A1(net4518),
    .Y(_05884_),
    .A2(_05067_));
 sg13g2_a21oi_1 _12518_ (.A1(net4158),
    .A2(_05884_),
    .Y(_05885_),
    .B1(net4004));
 sg13g2_nand2b_1 _12519_ (.Y(_05886_),
    .B(\cpu.keccak_alu.registers[176] ),
    .A_N(\cpu.keccak_alu.registers[112] ));
 sg13g2_a22oi_1 _12520_ (.Y(_05887_),
    .B1(_05886_),
    .B2(net4004),
    .A2(_05885_),
    .A1(_05875_));
 sg13g2_a21oi_1 _12521_ (.A1(\cpu.keccak_alu.registers[48] ),
    .A2(_05887_),
    .Y(_05888_),
    .B1(net4385));
 sg13g2_o21ai_1 _12522_ (.B1(_05888_),
    .Y(_05889_),
    .A1(\cpu.keccak_alu.registers[48] ),
    .A2(_05887_));
 sg13g2_a21oi_1 _12523_ (.A1(\cpu.keccak_alu.registers[176] ),
    .A2(\cpu.keccak_alu.registers[240] ),
    .Y(_05890_),
    .B1(net4370));
 sg13g2_o21ai_1 _12524_ (.B1(_05890_),
    .Y(_05891_),
    .A1(\cpu.keccak_alu.registers[176] ),
    .A2(\cpu.keccak_alu.registers[240] ));
 sg13g2_xnor2_1 _12525_ (.Y(_05892_),
    .A(\cpu.keccak_alu.registers[48] ),
    .B(\cpu.keccak_alu.registers[112] ));
 sg13g2_xnor2_1 _12526_ (.Y(_05893_),
    .A(_05891_),
    .B(_05892_));
 sg13g2_o21ai_1 _12527_ (.B1(_05889_),
    .Y(_05894_),
    .A1(net4219),
    .A2(_05893_));
 sg13g2_nor3_2 _12528_ (.A(net3962),
    .B(_02360_),
    .C(net3718),
    .Y(_05895_));
 sg13g2_nor2_1 _12529_ (.A(net172),
    .B(net3633),
    .Y(_05896_));
 sg13g2_a21oi_1 _12530_ (.A1(net4363),
    .A2(net3633),
    .Y(_05897_),
    .B1(_05896_));
 sg13g2_a221oi_1 _12531_ (.B2(net3819),
    .C1(net3736),
    .B1(_05897_),
    .A1(net4265),
    .Y(_05898_),
    .A2(_05894_));
 sg13g2_a21oi_1 _12532_ (.A1(_01000_),
    .A2(net3736),
    .Y(_00765_),
    .B1(_05898_));
 sg13g2_nand3b_1 _12533_ (.B(\cpu.keccak_alu.registers[177] ),
    .C(net4006),
    .Y(_05899_),
    .A_N(\cpu.keccak_alu.registers[113] ));
 sg13g2_or2_1 _12534_ (.X(_05900_),
    .B(_05808_),
    .A(net4185));
 sg13g2_o21ai_1 _12535_ (.B1(net3831),
    .Y(_05901_),
    .A1(_04365_),
    .A2(_04398_));
 sg13g2_nand2b_1 _12536_ (.Y(_05902_),
    .B(net4197),
    .A_N(_05901_));
 sg13g2_o21ai_1 _12537_ (.B1(_05902_),
    .Y(_05903_),
    .A1(net4197),
    .A2(_05854_));
 sg13g2_o21ai_1 _12538_ (.B1(_05900_),
    .Y(_05904_),
    .A1(net4533),
    .A2(_05903_));
 sg13g2_nor2_1 _12539_ (.A(net4528),
    .B(_05904_),
    .Y(_05905_));
 sg13g2_a21oi_1 _12540_ (.A1(net4528),
    .A2(_05717_),
    .Y(_05906_),
    .B1(_05905_));
 sg13g2_o21ai_1 _12541_ (.B1(net4159),
    .Y(_05907_),
    .A1(_05520_),
    .A2(net3875));
 sg13g2_a221oi_1 _12542_ (.B2(net4092),
    .C1(_05907_),
    .B1(_05906_),
    .A1(net4519),
    .Y(_05908_),
    .A2(_05100_));
 sg13g2_nand3_1 _12543_ (.B(net3778),
    .C(_04507_),
    .A(net3921),
    .Y(_05909_));
 sg13g2_xor2_1 _12544_ (.B(_05909_),
    .A(_05908_),
    .X(_05910_));
 sg13g2_o21ai_1 _12545_ (.B1(_05899_),
    .Y(_05911_),
    .A1(net4006),
    .A2(_05910_));
 sg13g2_a21oi_1 _12546_ (.A1(\cpu.keccak_alu.registers[49] ),
    .A2(_05911_),
    .Y(_05912_),
    .B1(net4384));
 sg13g2_o21ai_1 _12547_ (.B1(_05912_),
    .Y(_05913_),
    .A1(\cpu.keccak_alu.registers[49] ),
    .A2(_05911_));
 sg13g2_o21ai_1 _12548_ (.B1(net4209),
    .Y(_05914_),
    .A1(\cpu.keccak_alu.registers[177] ),
    .A2(\cpu.keccak_alu.registers[241] ));
 sg13g2_a21oi_1 _12549_ (.A1(\cpu.keccak_alu.registers[177] ),
    .A2(\cpu.keccak_alu.registers[241] ),
    .Y(_05915_),
    .B1(_05914_));
 sg13g2_xor2_1 _12550_ (.B(\cpu.keccak_alu.registers[113] ),
    .A(\cpu.keccak_alu.registers[49] ),
    .X(_05916_));
 sg13g2_a21oi_1 _12551_ (.A1(_05915_),
    .A2(_05916_),
    .Y(_05917_),
    .B1(net4219));
 sg13g2_o21ai_1 _12552_ (.B1(_05917_),
    .Y(_05918_),
    .A1(_05915_),
    .A2(_05916_));
 sg13g2_a21oi_1 _12553_ (.A1(_05913_),
    .A2(_05918_),
    .Y(_05919_),
    .B1(net4321));
 sg13g2_o21ai_1 _12554_ (.B1(net3819),
    .Y(_05920_),
    .A1(net171),
    .A2(net3633));
 sg13g2_a21oi_1 _12555_ (.A1(net4358),
    .A2(net3633),
    .Y(_05921_),
    .B1(_05920_));
 sg13g2_nor3_1 _12556_ (.A(net3735),
    .B(_05919_),
    .C(_05921_),
    .Y(_05922_));
 sg13g2_a21oi_1 _12557_ (.A1(_01008_),
    .A2(net3735),
    .Y(_00766_),
    .B1(_05922_));
 sg13g2_a21oi_1 _12558_ (.A1(_01010_),
    .A2(\cpu.keccak_alu.registers[178] ),
    .Y(_05923_),
    .B1(net4020));
 sg13g2_nor2_1 _12559_ (.A(_05544_),
    .B(net3873),
    .Y(_05924_));
 sg13g2_o21ai_1 _12560_ (.B1(_04189_),
    .Y(_05925_),
    .A1(net4555),
    .A2(_01168_));
 sg13g2_nor2_1 _12561_ (.A(net4537),
    .B(_05925_),
    .Y(_05926_));
 sg13g2_a21oi_1 _12562_ (.A1(net4537),
    .A2(_05877_),
    .Y(_05927_),
    .B1(_05926_));
 sg13g2_mux2_1 _12563_ (.A0(_05831_),
    .A1(_05927_),
    .S(net4180),
    .X(_05928_));
 sg13g2_o21ai_1 _12564_ (.B1(net4092),
    .Y(_05929_),
    .A1(_05778_),
    .A2(_05928_));
 sg13g2_a21oi_1 _12565_ (.A1(net4526),
    .A2(_05739_),
    .Y(_05930_),
    .B1(_05929_));
 sg13g2_nor3_1 _12566_ (.A(net4514),
    .B(_05924_),
    .C(_05930_),
    .Y(_05931_));
 sg13g2_o21ai_1 _12567_ (.B1(_05931_),
    .Y(_05932_),
    .A1(net4162),
    .A2(_05126_));
 sg13g2_nand3_1 _12568_ (.B(net3774),
    .C(_04577_),
    .A(net3916),
    .Y(_05933_));
 sg13g2_xnor2_1 _12569_ (.Y(_05934_),
    .A(_05932_),
    .B(_05933_));
 sg13g2_a21oi_1 _12570_ (.A1(net4020),
    .A2(_05934_),
    .Y(_05935_),
    .B1(_05923_));
 sg13g2_a21oi_1 _12571_ (.A1(\cpu.keccak_alu.registers[50] ),
    .A2(_05935_),
    .Y(_05936_),
    .B1(net4384));
 sg13g2_o21ai_1 _12572_ (.B1(_05936_),
    .Y(_05937_),
    .A1(\cpu.keccak_alu.registers[50] ),
    .A2(_05935_));
 sg13g2_o21ai_1 _12573_ (.B1(net4209),
    .Y(_05938_),
    .A1(\cpu.keccak_alu.registers[178] ),
    .A2(\cpu.keccak_alu.registers[242] ));
 sg13g2_a21oi_1 _12574_ (.A1(\cpu.keccak_alu.registers[178] ),
    .A2(\cpu.keccak_alu.registers[242] ),
    .Y(_05939_),
    .B1(_05938_));
 sg13g2_xor2_1 _12575_ (.B(\cpu.keccak_alu.registers[114] ),
    .A(\cpu.keccak_alu.registers[50] ),
    .X(_05940_));
 sg13g2_a21oi_1 _12576_ (.A1(_05939_),
    .A2(_05940_),
    .Y(_05941_),
    .B1(net4218));
 sg13g2_o21ai_1 _12577_ (.B1(_05941_),
    .Y(_05942_),
    .A1(_05939_),
    .A2(_05940_));
 sg13g2_a21oi_1 _12578_ (.A1(_05937_),
    .A2(_05942_),
    .Y(_05943_),
    .B1(net4321));
 sg13g2_o21ai_1 _12579_ (.B1(net3819),
    .Y(_05944_),
    .A1(net132),
    .A2(net3633));
 sg13g2_a21oi_1 _12580_ (.A1(net4355),
    .A2(net3633),
    .Y(_05945_),
    .B1(_05944_));
 sg13g2_nor3_1 _12581_ (.A(net3733),
    .B(_05943_),
    .C(_05945_),
    .Y(_05946_));
 sg13g2_a21oi_1 _12582_ (.A1(_01016_),
    .A2(net3733),
    .Y(_00767_),
    .B1(_05946_));
 sg13g2_o21ai_1 _12583_ (.B1(net4005),
    .Y(_05947_),
    .A1(\cpu.keccak_alu.registers[115] ),
    .A2(_01021_));
 sg13g2_a21oi_1 _12584_ (.A1(net4567),
    .A2(_01168_),
    .Y(_05948_),
    .B1(_04395_));
 sg13g2_nor2_1 _12585_ (.A(net3825),
    .B(_05948_),
    .Y(_05949_));
 sg13g2_nor2_1 _12586_ (.A(net4540),
    .B(_05949_),
    .Y(_05950_));
 sg13g2_a21oi_1 _12587_ (.A1(net4540),
    .A2(_05901_),
    .Y(_05951_),
    .B1(_05950_));
 sg13g2_mux2_1 _12588_ (.A0(_05856_),
    .A1(_05951_),
    .S(net4186),
    .X(_05952_));
 sg13g2_inv_1 _12589_ (.Y(_05953_),
    .A(_05952_));
 sg13g2_nand2_1 _12590_ (.Y(_05954_),
    .A(net4176),
    .B(_05952_));
 sg13g2_a21oi_1 _12591_ (.A1(net4529),
    .A2(_05764_),
    .Y(_05955_),
    .B1(net3936));
 sg13g2_o21ai_1 _12592_ (.B1(net4159),
    .Y(_05956_),
    .A1(_05569_),
    .A2(net3874));
 sg13g2_a221oi_1 _12593_ (.B2(_05955_),
    .C1(_05956_),
    .B1(_05954_),
    .A1(net4519),
    .Y(_05957_),
    .A2(_05154_));
 sg13g2_nand2_1 _12594_ (.Y(_05958_),
    .A(net3778),
    .B(_05156_));
 sg13g2_xnor2_1 _12595_ (.Y(_05959_),
    .A(_05957_),
    .B(_05958_));
 sg13g2_o21ai_1 _12596_ (.B1(_05947_),
    .Y(_05960_),
    .A1(net4007),
    .A2(_05959_));
 sg13g2_xor2_1 _12597_ (.B(_05960_),
    .A(\cpu.keccak_alu.registers[51] ),
    .X(_05961_));
 sg13g2_o21ai_1 _12598_ (.B1(net4210),
    .Y(_05962_),
    .A1(\cpu.keccak_alu.registers[179] ),
    .A2(\cpu.keccak_alu.registers[243] ));
 sg13g2_a21oi_1 _12599_ (.A1(\cpu.keccak_alu.registers[179] ),
    .A2(\cpu.keccak_alu.registers[243] ),
    .Y(_05963_),
    .B1(_05962_));
 sg13g2_xor2_1 _12600_ (.B(\cpu.keccak_alu.registers[115] ),
    .A(\cpu.keccak_alu.registers[51] ),
    .X(_05964_));
 sg13g2_a21oi_1 _12601_ (.A1(_05963_),
    .A2(_05964_),
    .Y(_05965_),
    .B1(net4219));
 sg13g2_o21ai_1 _12602_ (.B1(_05965_),
    .Y(_05966_),
    .A1(_05963_),
    .A2(_05964_));
 sg13g2_o21ai_1 _12603_ (.B1(_05966_),
    .Y(_05967_),
    .A1(net4385),
    .A2(_05961_));
 sg13g2_nor2_1 _12604_ (.A(net180),
    .B(net3632),
    .Y(_05968_));
 sg13g2_a21oi_1 _12605_ (.A1(net4350),
    .A2(net3632),
    .Y(_05969_),
    .B1(_05968_));
 sg13g2_a221oi_1 _12606_ (.B2(net3819),
    .C1(net3733),
    .B1(_05969_),
    .A1(net4264),
    .Y(_05970_),
    .A2(_05967_));
 sg13g2_a21oi_1 _12607_ (.A1(_01025_),
    .A2(net3733),
    .Y(_00768_),
    .B1(_05970_));
 sg13g2_nand2b_1 _12608_ (.Y(_05971_),
    .B(\cpu.keccak_alu.registers[180] ),
    .A_N(\cpu.keccak_alu.registers[116] ));
 sg13g2_nand2_1 _12609_ (.Y(_05972_),
    .A(net4526),
    .B(_04301_));
 sg13g2_nor2_1 _12610_ (.A(net4191),
    .B(_05925_),
    .Y(_05973_));
 sg13g2_nor2_1 _12611_ (.A(_04186_),
    .B(_04198_),
    .Y(_05974_));
 sg13g2_a21oi_1 _12612_ (.A1(net4191),
    .A2(_05974_),
    .Y(_05975_),
    .B1(_05973_));
 sg13g2_mux2_1 _12613_ (.A0(_05879_),
    .A1(_05975_),
    .S(net4180),
    .X(_05976_));
 sg13g2_or2_1 _12614_ (.X(_05977_),
    .B(_05976_),
    .A(_05778_));
 sg13g2_a21oi_1 _12615_ (.A1(net4526),
    .A2(_05784_),
    .Y(_05978_),
    .B1(net3934));
 sg13g2_o21ai_1 _12616_ (.B1(net4157),
    .Y(_05979_),
    .A1(net3872),
    .A2(_05595_));
 sg13g2_a221oi_1 _12617_ (.B2(_05978_),
    .C1(_05979_),
    .B1(_05977_),
    .A1(\cpu.keccak_alu.registers[133] ),
    .Y(_05980_),
    .A2(_05179_));
 sg13g2_nand4_1 _12618_ (.B(net3773),
    .C(_04668_),
    .A(net3914),
    .Y(_05981_),
    .D(_04670_));
 sg13g2_xnor2_1 _12619_ (.Y(_05982_),
    .A(_05980_),
    .B(_05981_));
 sg13g2_nor2_1 _12620_ (.A(net4008),
    .B(_05982_),
    .Y(_05983_));
 sg13g2_a21oi_1 _12621_ (.A1(net4004),
    .A2(_05971_),
    .Y(_05984_),
    .B1(_05983_));
 sg13g2_a21oi_1 _12622_ (.A1(\cpu.keccak_alu.registers[52] ),
    .A2(_05984_),
    .Y(_05985_),
    .B1(net4382));
 sg13g2_o21ai_1 _12623_ (.B1(_05985_),
    .Y(_05986_),
    .A1(\cpu.keccak_alu.registers[52] ),
    .A2(_05984_));
 sg13g2_o21ai_1 _12624_ (.B1(net4211),
    .Y(_05987_),
    .A1(net4487),
    .A2(\cpu.keccak_alu.registers[244] ));
 sg13g2_a21oi_1 _12625_ (.A1(net4487),
    .A2(\cpu.keccak_alu.registers[244] ),
    .Y(_05988_),
    .B1(_05987_));
 sg13g2_xor2_1 _12626_ (.B(\cpu.keccak_alu.registers[116] ),
    .A(\cpu.keccak_alu.registers[52] ),
    .X(_05989_));
 sg13g2_a21oi_1 _12627_ (.A1(_05988_),
    .A2(_05989_),
    .Y(_05990_),
    .B1(net4220));
 sg13g2_o21ai_1 _12628_ (.B1(_05990_),
    .Y(_05991_),
    .A1(_05988_),
    .A2(_05989_));
 sg13g2_a21o_1 _12629_ (.A2(_05991_),
    .A1(_05986_),
    .B1(net4319),
    .X(_05992_));
 sg13g2_o21ai_1 _12630_ (.B1(net3820),
    .Y(_05993_),
    .A1(net332),
    .A2(net3632));
 sg13g2_a21oi_1 _12631_ (.A1(net4347),
    .A2(net3632),
    .Y(_05994_),
    .B1(_05993_));
 sg13g2_nor2_1 _12632_ (.A(net3732),
    .B(_05994_),
    .Y(_05995_));
 sg13g2_a22oi_1 _12633_ (.Y(_00769_),
    .B1(_05992_),
    .B2(_05995_),
    .A2(net3737),
    .A1(_01033_));
 sg13g2_a21oi_1 _12634_ (.A1(_01035_),
    .A2(net4486),
    .Y(_05996_),
    .B1(net4017));
 sg13g2_nor2_1 _12635_ (.A(net4163),
    .B(_05200_),
    .Y(_05997_));
 sg13g2_nor2_1 _12636_ (.A(net4185),
    .B(_05903_),
    .Y(_05998_));
 sg13g2_o21ai_1 _12637_ (.B1(net3831),
    .Y(_05999_),
    .A1(_04396_),
    .A2(_04408_));
 sg13g2_nor2_1 _12638_ (.A(net4540),
    .B(_05999_),
    .Y(_06000_));
 sg13g2_a21oi_1 _12639_ (.A1(net4540),
    .A2(_05949_),
    .Y(_06001_),
    .B1(_06000_));
 sg13g2_a21oi_1 _12640_ (.A1(net4186),
    .A2(_06001_),
    .Y(_06002_),
    .B1(_05998_));
 sg13g2_inv_1 _12641_ (.Y(_06003_),
    .A(_06002_));
 sg13g2_a21oi_1 _12642_ (.A1(net4528),
    .A2(_05809_),
    .Y(_06004_),
    .B1(net3936));
 sg13g2_o21ai_1 _12643_ (.B1(_06004_),
    .Y(_06005_),
    .A1(net4528),
    .A2(_06003_));
 sg13g2_o21ai_1 _12644_ (.B1(_06005_),
    .Y(_06006_),
    .A1(net3874),
    .A2(_05620_));
 sg13g2_nor3_1 _12645_ (.A(net4515),
    .B(_05997_),
    .C(_06006_),
    .Y(_06007_));
 sg13g2_nand3_1 _12646_ (.B(net3776),
    .C(_04716_),
    .A(net3918),
    .Y(_06008_));
 sg13g2_xor2_1 _12647_ (.B(_06008_),
    .A(_06007_),
    .X(_06009_));
 sg13g2_a21oi_2 _12648_ (.B1(_05996_),
    .Y(_06010_),
    .A2(_06009_),
    .A1(net4017));
 sg13g2_a21oi_1 _12649_ (.A1(\cpu.keccak_alu.registers[53] ),
    .A2(_06010_),
    .Y(_06011_),
    .B1(net4382));
 sg13g2_o21ai_1 _12650_ (.B1(_06011_),
    .Y(_06012_),
    .A1(\cpu.keccak_alu.registers[53] ),
    .A2(_06010_));
 sg13g2_a21oi_1 _12651_ (.A1(net4486),
    .A2(\cpu.keccak_alu.registers[245] ),
    .Y(_06013_),
    .B1(net4370));
 sg13g2_o21ai_1 _12652_ (.B1(_06013_),
    .Y(_06014_),
    .A1(net4486),
    .A2(\cpu.keccak_alu.registers[245] ));
 sg13g2_xnor2_1 _12653_ (.Y(_06015_),
    .A(\cpu.keccak_alu.registers[53] ),
    .B(\cpu.keccak_alu.registers[117] ));
 sg13g2_a21oi_1 _12654_ (.A1(_06014_),
    .A2(_06015_),
    .Y(_06016_),
    .B1(net4216));
 sg13g2_o21ai_1 _12655_ (.B1(_06016_),
    .Y(_06017_),
    .A1(_06014_),
    .A2(_06015_));
 sg13g2_a21oi_1 _12656_ (.A1(_06012_),
    .A2(_06017_),
    .Y(_06018_),
    .B1(net4320));
 sg13g2_o21ai_1 _12657_ (.B1(net3819),
    .Y(_06019_),
    .A1(net164),
    .A2(net3632));
 sg13g2_a21oi_1 _12658_ (.A1(net4343),
    .A2(net3632),
    .Y(_06020_),
    .B1(_06019_));
 sg13g2_nor3_1 _12659_ (.A(net3730),
    .B(_06018_),
    .C(_06020_),
    .Y(_06021_));
 sg13g2_a21oi_1 _12660_ (.A1(_01041_),
    .A2(net3730),
    .Y(_00770_),
    .B1(_06021_));
 sg13g2_a21oi_1 _12661_ (.A1(net4485),
    .A2(\cpu.keccak_alu.registers[246] ),
    .Y(_06022_),
    .B1(net4370));
 sg13g2_o21ai_1 _12662_ (.B1(_06022_),
    .Y(_06023_),
    .A1(net4485),
    .A2(\cpu.keccak_alu.registers[246] ));
 sg13g2_xnor2_1 _12663_ (.Y(_06024_),
    .A(\cpu.keccak_alu.registers[54] ),
    .B(\cpu.keccak_alu.registers[118] ));
 sg13g2_xnor2_1 _12664_ (.Y(_06025_),
    .A(_06023_),
    .B(_06024_));
 sg13g2_a21oi_1 _12665_ (.A1(_01045_),
    .A2(\cpu.keccak_alu.registers[182] ),
    .Y(_06026_),
    .B1(net4017));
 sg13g2_nor2_1 _12666_ (.A(net3871),
    .B(_05645_),
    .Y(_06027_));
 sg13g2_nor3_1 _12667_ (.A(net4537),
    .B(_04196_),
    .C(_04199_),
    .Y(_06028_));
 sg13g2_a21oi_1 _12668_ (.A1(net4537),
    .A2(_05974_),
    .Y(_06029_),
    .B1(_06028_));
 sg13g2_mux2_1 _12669_ (.A0(_05927_),
    .A1(_06029_),
    .S(net4180),
    .X(_06030_));
 sg13g2_o21ai_1 _12670_ (.B1(net4091),
    .Y(_06031_),
    .A1(_05778_),
    .A2(_06030_));
 sg13g2_a21oi_1 _12671_ (.A1(net4526),
    .A2(_05833_),
    .Y(_06032_),
    .B1(_06031_));
 sg13g2_nor3_1 _12672_ (.A(net4514),
    .B(_06027_),
    .C(_06032_),
    .Y(_06033_));
 sg13g2_o21ai_1 _12673_ (.B1(_06033_),
    .Y(_06034_),
    .A1(net4161),
    .A2(_05231_));
 sg13g2_nand3_1 _12674_ (.B(net3772),
    .C(_04751_),
    .A(net3915),
    .Y(_06035_));
 sg13g2_xnor2_1 _12675_ (.Y(_06036_),
    .A(_06034_),
    .B(_06035_));
 sg13g2_a21oi_1 _12676_ (.A1(net4017),
    .A2(_06036_),
    .Y(_06037_),
    .B1(_06026_));
 sg13g2_a21oi_1 _12677_ (.A1(\cpu.keccak_alu.registers[54] ),
    .A2(_06037_),
    .Y(_06038_),
    .B1(net4383));
 sg13g2_o21ai_1 _12678_ (.B1(_06038_),
    .Y(_06039_),
    .A1(\cpu.keccak_alu.registers[54] ),
    .A2(_06037_));
 sg13g2_o21ai_1 _12679_ (.B1(_06039_),
    .Y(_06040_),
    .A1(net4220),
    .A2(_06025_));
 sg13g2_nor2_1 _12680_ (.A(net195),
    .B(net3632),
    .Y(_06041_));
 sg13g2_a21oi_1 _12681_ (.A1(net4339),
    .A2(net3632),
    .Y(_06042_),
    .B1(_06041_));
 sg13g2_a221oi_1 _12682_ (.B2(net3819),
    .C1(net3730),
    .B1(_06042_),
    .A1(net4259),
    .Y(_06043_),
    .A2(_06040_));
 sg13g2_a21oi_1 _12683_ (.A1(_01051_),
    .A2(net3730),
    .Y(_00771_),
    .B1(_06043_));
 sg13g2_a21oi_1 _12684_ (.A1(_01054_),
    .A2(\cpu.keccak_alu.registers[183] ),
    .Y(_06044_),
    .B1(net4014));
 sg13g2_nor2_1 _12685_ (.A(net4186),
    .B(_05951_),
    .Y(_06045_));
 sg13g2_o21ai_1 _12686_ (.B1(net3831),
    .Y(_06046_),
    .A1(_04404_),
    .A2(_04409_));
 sg13g2_mux2_1 _12687_ (.A0(_05999_),
    .A1(_06046_),
    .S(net4197),
    .X(_06047_));
 sg13g2_a21oi_1 _12688_ (.A1(net4186),
    .A2(_06047_),
    .Y(_06048_),
    .B1(_06045_));
 sg13g2_nand2_1 _12689_ (.Y(_06049_),
    .A(net4175),
    .B(_06048_));
 sg13g2_a21oi_1 _12690_ (.A1(net4528),
    .A2(_05857_),
    .Y(_06050_),
    .B1(net3936));
 sg13g2_o21ai_1 _12691_ (.B1(net4159),
    .Y(_06051_),
    .A1(net3874),
    .A2(_05664_));
 sg13g2_a221oi_1 _12692_ (.B2(_06050_),
    .C1(_06051_),
    .B1(_06049_),
    .A1(net4519),
    .Y(_06052_),
    .A2(_05257_));
 sg13g2_nand3_1 _12693_ (.B(net3776),
    .C(_04791_),
    .A(net3922),
    .Y(_06053_));
 sg13g2_xor2_1 _12694_ (.B(_06053_),
    .A(_06052_),
    .X(_06054_));
 sg13g2_a21oi_2 _12695_ (.B1(_06044_),
    .Y(_06055_),
    .A2(_06054_),
    .A1(net4018));
 sg13g2_a21oi_1 _12696_ (.A1(\cpu.keccak_alu.registers[55] ),
    .A2(_06055_),
    .Y(_06056_),
    .B1(net4378));
 sg13g2_o21ai_1 _12697_ (.B1(_06056_),
    .Y(_06057_),
    .A1(\cpu.keccak_alu.registers[55] ),
    .A2(_06055_));
 sg13g2_o21ai_1 _12698_ (.B1(net4207),
    .Y(_06058_),
    .A1(\cpu.keccak_alu.registers[183] ),
    .A2(\cpu.keccak_alu.registers[247] ));
 sg13g2_a21oi_1 _12699_ (.A1(\cpu.keccak_alu.registers[183] ),
    .A2(\cpu.keccak_alu.registers[247] ),
    .Y(_06059_),
    .B1(_06058_));
 sg13g2_xor2_1 _12700_ (.B(\cpu.keccak_alu.registers[119] ),
    .A(\cpu.keccak_alu.registers[55] ),
    .X(_06060_));
 sg13g2_a21oi_1 _12701_ (.A1(_06059_),
    .A2(_06060_),
    .Y(_06061_),
    .B1(net4216));
 sg13g2_o21ai_1 _12702_ (.B1(_06061_),
    .Y(_06062_),
    .A1(_06059_),
    .A2(_06060_));
 sg13g2_a21oi_1 _12703_ (.A1(_06057_),
    .A2(_06062_),
    .Y(_06063_),
    .B1(net4315));
 sg13g2_o21ai_1 _12704_ (.B1(net3818),
    .Y(_06064_),
    .A1(net173),
    .A2(net3631));
 sg13g2_a21oi_1 _12705_ (.A1(net4336),
    .A2(net3631),
    .Y(_06065_),
    .B1(_06064_));
 sg13g2_nor3_1 _12706_ (.A(net3728),
    .B(_06063_),
    .C(_06065_),
    .Y(_06066_));
 sg13g2_a21oi_1 _12707_ (.A1(_01060_),
    .A2(net3728),
    .Y(_00772_),
    .B1(_06066_));
 sg13g2_a21oi_1 _12708_ (.A1(\cpu.keccak_alu.registers[184] ),
    .A2(\cpu.keccak_alu.registers[248] ),
    .Y(_06067_),
    .B1(net4369));
 sg13g2_o21ai_1 _12709_ (.B1(_06067_),
    .Y(_06068_),
    .A1(\cpu.keccak_alu.registers[184] ),
    .A2(\cpu.keccak_alu.registers[248] ));
 sg13g2_xor2_1 _12710_ (.B(\cpu.keccak_alu.registers[120] ),
    .A(\cpu.keccak_alu.registers[56] ),
    .X(_06069_));
 sg13g2_xnor2_1 _12711_ (.Y(_06070_),
    .A(_06068_),
    .B(_06069_));
 sg13g2_a21oi_1 _12712_ (.A1(net4553),
    .A2(_00121_),
    .Y(_06071_),
    .B1(_04163_));
 sg13g2_nor3_1 _12713_ (.A(net4192),
    .B(_04196_),
    .C(_04199_),
    .Y(_06072_));
 sg13g2_a21oi_1 _12714_ (.A1(net4192),
    .A2(_06071_),
    .Y(_06073_),
    .B1(_06072_));
 sg13g2_mux2_1 _12715_ (.A0(_05975_),
    .A1(_06073_),
    .S(net4180),
    .X(_06074_));
 sg13g2_o21ai_1 _12716_ (.B1(net4091),
    .Y(_06075_),
    .A1(_05778_),
    .A2(_06074_));
 sg13g2_a21oi_1 _12717_ (.A1(net4526),
    .A2(_05881_),
    .Y(_06076_),
    .B1(_06075_));
 sg13g2_nor2_1 _12718_ (.A(net4513),
    .B(_06076_),
    .Y(_06077_));
 sg13g2_o21ai_1 _12719_ (.B1(_06077_),
    .Y(_06078_),
    .A1(net3871),
    .A2(_05695_));
 sg13g2_a21oi_1 _12720_ (.A1(net4517),
    .A2(_05285_),
    .Y(_06079_),
    .B1(_06078_));
 sg13g2_nand3_1 _12721_ (.B(net3773),
    .C(_04820_),
    .A(net3915),
    .Y(_06080_));
 sg13g2_o21ai_1 _12722_ (.B1(net4001),
    .Y(_06081_),
    .A1(\cpu.keccak_alu.registers[120] ),
    .A2(_01065_));
 sg13g2_xnor2_1 _12723_ (.Y(_06082_),
    .A(_06079_),
    .B(_06080_));
 sg13g2_o21ai_1 _12724_ (.B1(_06081_),
    .Y(_06083_),
    .A1(net4001),
    .A2(_06082_));
 sg13g2_nand2b_1 _12725_ (.Y(_06084_),
    .B(\cpu.keccak_alu.registers[56] ),
    .A_N(_06083_));
 sg13g2_a21oi_1 _12726_ (.A1(_01061_),
    .A2(_06083_),
    .Y(_06085_),
    .B1(net4379));
 sg13g2_a22oi_1 _12727_ (.Y(_06086_),
    .B1(_06084_),
    .B2(_06085_),
    .A2(_06070_),
    .A1(net4379));
 sg13g2_nor2_1 _12728_ (.A(net4315),
    .B(_06086_),
    .Y(_06087_));
 sg13g2_o21ai_1 _12729_ (.B1(net3818),
    .Y(_06088_),
    .A1(net157),
    .A2(net3630));
 sg13g2_a21oi_1 _12730_ (.A1(net4295),
    .A2(net3629),
    .Y(_06089_),
    .B1(_06088_));
 sg13g2_nor3_1 _12731_ (.A(net3726),
    .B(_06087_),
    .C(_06089_),
    .Y(_06090_));
 sg13g2_a21oi_1 _12732_ (.A1(_01069_),
    .A2(net3726),
    .Y(_00773_),
    .B1(_06090_));
 sg13g2_nand2b_1 _12733_ (.Y(_06091_),
    .B(\cpu.keccak_alu.registers[185] ),
    .A_N(\cpu.keccak_alu.registers[121] ));
 sg13g2_nand2_1 _12734_ (.Y(_06092_),
    .A(net4528),
    .B(_05904_));
 sg13g2_nor2_2 _12735_ (.A(net4185),
    .B(net4527),
    .Y(_06093_));
 sg13g2_o21ai_1 _12736_ (.B1(net3827),
    .Y(_06094_),
    .A1(_04378_),
    .A2(_04405_));
 sg13g2_mux2_1 _12737_ (.A0(_06046_),
    .A1(_06094_),
    .S(net4196),
    .X(_06095_));
 sg13g2_a22oi_1 _12738_ (.Y(_06096_),
    .B1(_06095_),
    .B2(_03865_),
    .A2(_06093_),
    .A1(_06001_));
 sg13g2_a21oi_1 _12739_ (.A1(_06092_),
    .A2(_06096_),
    .Y(_06097_),
    .B1(net3936));
 sg13g2_nor2_1 _12740_ (.A(net4515),
    .B(_06097_),
    .Y(_06098_));
 sg13g2_o21ai_1 _12741_ (.B1(_06098_),
    .Y(_06099_),
    .A1(net3875),
    .A2(_05718_));
 sg13g2_a21oi_1 _12742_ (.A1(net4519),
    .A2(_05307_),
    .Y(_06100_),
    .B1(_06099_));
 sg13g2_nand2_1 _12743_ (.Y(_06101_),
    .A(net3777),
    .B(_05309_));
 sg13g2_xor2_1 _12744_ (.B(_06101_),
    .A(_06100_),
    .X(_06102_));
 sg13g2_mux2_1 _12745_ (.A0(_06091_),
    .A1(_06102_),
    .S(net4010),
    .X(_06103_));
 sg13g2_a21oi_1 _12746_ (.A1(_01071_),
    .A2(_06103_),
    .Y(_06104_),
    .B1(net4372));
 sg13g2_o21ai_1 _12747_ (.B1(_06104_),
    .Y(_06105_),
    .A1(_01071_),
    .A2(_06103_));
 sg13g2_a21oi_1 _12748_ (.A1(\cpu.keccak_alu.registers[185] ),
    .A2(\cpu.keccak_alu.registers[249] ),
    .Y(_06106_),
    .B1(net4366));
 sg13g2_o21ai_1 _12749_ (.B1(_06106_),
    .Y(_06107_),
    .A1(\cpu.keccak_alu.registers[185] ),
    .A2(\cpu.keccak_alu.registers[249] ));
 sg13g2_xnor2_1 _12750_ (.Y(_06108_),
    .A(\cpu.keccak_alu.registers[57] ),
    .B(\cpu.keccak_alu.registers[121] ));
 sg13g2_o21ai_1 _12751_ (.B1(net4372),
    .Y(_06109_),
    .A1(_06107_),
    .A2(_06108_));
 sg13g2_a21o_1 _12752_ (.A2(_06108_),
    .A1(_06107_),
    .B1(_06109_),
    .X(_06110_));
 sg13g2_a21o_1 _12753_ (.A2(_06110_),
    .A1(_06105_),
    .B1(net4313),
    .X(_06111_));
 sg13g2_o21ai_1 _12754_ (.B1(net3815),
    .Y(_06112_),
    .A1(net237),
    .A2(net3629));
 sg13g2_a21oi_1 _12755_ (.A1(net4290),
    .A2(net3629),
    .Y(_06113_),
    .B1(_06112_));
 sg13g2_nor2_1 _12756_ (.A(net3721),
    .B(_06113_),
    .Y(_06114_));
 sg13g2_a22oi_1 _12757_ (.Y(_00774_),
    .B1(_06111_),
    .B2(_06114_),
    .A2(net3721),
    .A1(_01077_));
 sg13g2_nand3b_1 _12758_ (.B(\cpu.keccak_alu.registers[186] ),
    .C(net4000),
    .Y(_06115_),
    .A_N(\cpu.keccak_alu.registers[122] ));
 sg13g2_nor2b_2 _12759_ (.A(_04160_),
    .B_N(_04164_),
    .Y(_06116_));
 sg13g2_and2_1 _12760_ (.A(net4192),
    .B(_06116_),
    .X(_06117_));
 sg13g2_a21oi_1 _12761_ (.A1(net4535),
    .A2(_06071_),
    .Y(_06118_),
    .B1(_06117_));
 sg13g2_mux2_1 _12762_ (.A0(_06029_),
    .A1(_06118_),
    .S(net4180),
    .X(_06119_));
 sg13g2_nor2_1 _12763_ (.A(_05778_),
    .B(_06119_),
    .Y(_06120_));
 sg13g2_o21ai_1 _12764_ (.B1(net4091),
    .Y(_06121_),
    .A1(_05928_),
    .A2(_05972_));
 sg13g2_o21ai_1 _12765_ (.B1(net4157),
    .Y(_06122_),
    .A1(_06120_),
    .A2(_06121_));
 sg13g2_nor2_1 _12766_ (.A(net3872),
    .B(_05740_),
    .Y(_06123_));
 sg13g2_nor2_1 _12767_ (.A(_06122_),
    .B(_06123_),
    .Y(_06124_));
 sg13g2_o21ai_1 _12768_ (.B1(_06124_),
    .Y(_06125_),
    .A1(net4161),
    .A2(_05332_));
 sg13g2_nand3_1 _12769_ (.B(net3773),
    .C(_04882_),
    .A(net3915),
    .Y(_06126_));
 sg13g2_xnor2_1 _12770_ (.Y(_06127_),
    .A(_06125_),
    .B(_06126_));
 sg13g2_o21ai_1 _12771_ (.B1(_06115_),
    .Y(_06128_),
    .A1(net4000),
    .A2(_06127_));
 sg13g2_a21oi_1 _12772_ (.A1(\cpu.keccak_alu.registers[58] ),
    .A2(_06128_),
    .Y(_06129_),
    .B1(net4372));
 sg13g2_o21ai_1 _12773_ (.B1(_06129_),
    .Y(_06130_),
    .A1(\cpu.keccak_alu.registers[58] ),
    .A2(_06128_));
 sg13g2_a21oi_1 _12774_ (.A1(\cpu.keccak_alu.registers[186] ),
    .A2(\cpu.keccak_alu.registers[250] ),
    .Y(_06131_),
    .B1(net4366));
 sg13g2_o21ai_1 _12775_ (.B1(_06131_),
    .Y(_06132_),
    .A1(\cpu.keccak_alu.registers[186] ),
    .A2(\cpu.keccak_alu.registers[250] ));
 sg13g2_xnor2_1 _12776_ (.Y(_06133_),
    .A(\cpu.keccak_alu.registers[58] ),
    .B(\cpu.keccak_alu.registers[122] ));
 sg13g2_o21ai_1 _12777_ (.B1(net4372),
    .Y(_06134_),
    .A1(_06132_),
    .A2(_06133_));
 sg13g2_a21o_1 _12778_ (.A2(_06133_),
    .A1(_06132_),
    .B1(_06134_),
    .X(_06135_));
 sg13g2_a21oi_1 _12779_ (.A1(_06130_),
    .A2(_06135_),
    .Y(_06136_),
    .B1(net4313));
 sg13g2_o21ai_1 _12780_ (.B1(net3816),
    .Y(_06137_),
    .A1(net128),
    .A2(net3629));
 sg13g2_a21oi_1 _12781_ (.A1(net4286),
    .A2(net3629),
    .Y(_06138_),
    .B1(_06137_));
 sg13g2_nor3_1 _12782_ (.A(net3721),
    .B(_06136_),
    .C(_06138_),
    .Y(_06139_));
 sg13g2_a21oi_1 _12783_ (.A1(_01084_),
    .A2(net3722),
    .Y(_00775_),
    .B1(_06139_));
 sg13g2_o21ai_1 _12784_ (.B1(_04379_),
    .Y(_06140_),
    .A1(net4548),
    .A2(_00125_));
 sg13g2_and2_1 _12785_ (.A(net3827),
    .B(_06140_),
    .X(_06141_));
 sg13g2_nor2_1 _12786_ (.A(net4535),
    .B(_06141_),
    .Y(_06142_));
 sg13g2_a21oi_2 _12787_ (.B1(_06142_),
    .Y(_06143_),
    .A2(_06094_),
    .A1(net4535));
 sg13g2_inv_1 _12788_ (.Y(_06144_),
    .A(_06143_));
 sg13g2_a22oi_1 _12789_ (.Y(_06145_),
    .B1(_06047_),
    .B2(_06093_),
    .A2(_05953_),
    .A1(net4527));
 sg13g2_o21ai_1 _12790_ (.B1(_06145_),
    .Y(_06146_),
    .A1(_03866_),
    .A2(_06143_));
 sg13g2_o21ai_1 _12791_ (.B1(net4160),
    .Y(_06147_),
    .A1(net3876),
    .A2(_05765_));
 sg13g2_a221oi_1 _12792_ (.B2(net4092),
    .C1(_06147_),
    .B1(_06146_),
    .A1(net4520),
    .Y(_06148_),
    .A2(_05361_));
 sg13g2_nor4_2 _12793_ (.A(net3927),
    .B(net3793),
    .C(net3834),
    .Y(_06149_),
    .D(_04614_));
 sg13g2_o21ai_1 _12794_ (.B1(net4001),
    .Y(_06150_),
    .A1(\cpu.keccak_alu.registers[123] ),
    .A2(_01089_));
 sg13g2_xor2_1 _12795_ (.B(_06149_),
    .A(_06148_),
    .X(_06151_));
 sg13g2_o21ai_1 _12796_ (.B1(_06150_),
    .Y(_06152_),
    .A1(net4001),
    .A2(_06151_));
 sg13g2_nand2b_1 _12797_ (.Y(_06153_),
    .B(\cpu.keccak_alu.registers[59] ),
    .A_N(_06152_));
 sg13g2_a21oi_1 _12798_ (.A1(_01086_),
    .A2(_06152_),
    .Y(_06154_),
    .B1(net4374));
 sg13g2_a21oi_1 _12799_ (.A1(net4484),
    .A2(\cpu.keccak_alu.registers[251] ),
    .Y(_06155_),
    .B1(net4367));
 sg13g2_o21ai_1 _12800_ (.B1(_06155_),
    .Y(_06156_),
    .A1(net4484),
    .A2(\cpu.keccak_alu.registers[251] ));
 sg13g2_xor2_1 _12801_ (.B(\cpu.keccak_alu.registers[123] ),
    .A(\cpu.keccak_alu.registers[59] ),
    .X(_06157_));
 sg13g2_xnor2_1 _12802_ (.Y(_06158_),
    .A(_06156_),
    .B(_06157_));
 sg13g2_a22oi_1 _12803_ (.Y(_06159_),
    .B1(_06158_),
    .B2(net4374),
    .A2(_06154_),
    .A1(_06153_));
 sg13g2_nor2_1 _12804_ (.A(net4314),
    .B(_06159_),
    .Y(_06160_));
 sg13g2_o21ai_1 _12805_ (.B1(net3817),
    .Y(_06161_),
    .A1(net152),
    .A2(net3629));
 sg13g2_a21oi_1 _12806_ (.A1(net4282),
    .A2(net3630),
    .Y(_06162_),
    .B1(_06161_));
 sg13g2_nor3_1 _12807_ (.A(net3724),
    .B(_06160_),
    .C(_06162_),
    .Y(_06163_));
 sg13g2_a21oi_1 _12808_ (.A1(_01093_),
    .A2(net3724),
    .Y(_00776_),
    .B1(_06163_));
 sg13g2_a21oi_1 _12809_ (.A1(_01096_),
    .A2(net4483),
    .Y(_06164_),
    .B1(net4014));
 sg13g2_nor2_1 _12810_ (.A(_04161_),
    .B(_04172_),
    .Y(_06165_));
 sg13g2_nand2_1 _12811_ (.Y(_06166_),
    .A(net4191),
    .B(_06165_));
 sg13g2_a21oi_1 _12812_ (.A1(net4535),
    .A2(_06116_),
    .Y(_06167_),
    .B1(net4531));
 sg13g2_a221oi_1 _12813_ (.B2(_06167_),
    .C1(_05778_),
    .B1(_06166_),
    .A1(net4531),
    .Y(_06168_),
    .A2(_06073_));
 sg13g2_o21ai_1 _12814_ (.B1(net4091),
    .Y(_06169_),
    .A1(_05972_),
    .A2(_05976_));
 sg13g2_nor2_1 _12815_ (.A(_06168_),
    .B(_06169_),
    .Y(_06170_));
 sg13g2_nor2_1 _12816_ (.A(net3871),
    .B(_05785_),
    .Y(_06171_));
 sg13g2_nor3_1 _12817_ (.A(net4513),
    .B(_06170_),
    .C(_06171_),
    .Y(_06172_));
 sg13g2_o21ai_1 _12818_ (.B1(_06172_),
    .Y(_06173_),
    .A1(net4161),
    .A2(_05387_));
 sg13g2_nor3_1 _12819_ (.A(net3923),
    .B(net3833),
    .C(_04942_),
    .Y(_06174_));
 sg13g2_xor2_1 _12820_ (.B(_06174_),
    .A(_06173_),
    .X(_06175_));
 sg13g2_a21oi_1 _12821_ (.A1(net4014),
    .A2(_06175_),
    .Y(_06176_),
    .B1(_06164_));
 sg13g2_a21oi_1 _12822_ (.A1(\cpu.keccak_alu.registers[60] ),
    .A2(_06176_),
    .Y(_06177_),
    .B1(net4377));
 sg13g2_o21ai_1 _12823_ (.B1(_06177_),
    .Y(_06178_),
    .A1(\cpu.keccak_alu.registers[60] ),
    .A2(_06176_));
 sg13g2_o21ai_1 _12824_ (.B1(net4207),
    .Y(_06179_),
    .A1(net4483),
    .A2(\cpu.keccak_alu.registers[252] ));
 sg13g2_a21oi_1 _12825_ (.A1(net4483),
    .A2(\cpu.keccak_alu.registers[252] ),
    .Y(_06180_),
    .B1(_06179_));
 sg13g2_xor2_1 _12826_ (.B(\cpu.keccak_alu.registers[124] ),
    .A(\cpu.keccak_alu.registers[60] ),
    .X(_06181_));
 sg13g2_a21oi_1 _12827_ (.A1(_06180_),
    .A2(_06181_),
    .Y(_06182_),
    .B1(net4216));
 sg13g2_o21ai_1 _12828_ (.B1(_06182_),
    .Y(_06183_),
    .A1(_06180_),
    .A2(_06181_));
 sg13g2_a21oi_1 _12829_ (.A1(_06178_),
    .A2(_06183_),
    .Y(_06184_),
    .B1(net4315));
 sg13g2_o21ai_1 _12830_ (.B1(net3818),
    .Y(_06185_),
    .A1(net189),
    .A2(net3631));
 sg13g2_a21oi_1 _12831_ (.A1(net4277),
    .A2(net3631),
    .Y(_06186_),
    .B1(_06185_));
 sg13g2_nor3_1 _12832_ (.A(net3727),
    .B(_06184_),
    .C(_06186_),
    .Y(_06187_));
 sg13g2_a21oi_1 _12833_ (.A1(_01102_),
    .A2(net3726),
    .Y(_00777_),
    .B1(_06187_));
 sg13g2_o21ai_1 _12834_ (.B1(net4160),
    .Y(_06188_),
    .A1(net3874),
    .A2(_05810_));
 sg13g2_a21o_1 _12835_ (.A2(_00126_),
    .A1(net4548),
    .B1(_04385_),
    .X(_06189_));
 sg13g2_nor2_1 _12836_ (.A(net4535),
    .B(_06189_),
    .Y(_06190_));
 sg13g2_a22oi_1 _12837_ (.Y(_06191_),
    .B1(_06190_),
    .B2(net3827),
    .A2(_06141_),
    .A1(net4535));
 sg13g2_a22oi_1 _12838_ (.Y(_06192_),
    .B1(_06191_),
    .B2(_03865_),
    .A2(_06095_),
    .A1(_06093_));
 sg13g2_o21ai_1 _12839_ (.B1(_06192_),
    .Y(_06193_),
    .A1(net4179),
    .A2(_06002_));
 sg13g2_a21oi_1 _12840_ (.A1(net4092),
    .A2(_06193_),
    .Y(_06194_),
    .B1(_06188_));
 sg13g2_o21ai_1 _12841_ (.B1(_06194_),
    .Y(_06195_),
    .A1(net4163),
    .A2(_05417_));
 sg13g2_nand4_1 _12842_ (.B(net3785),
    .C(net3776),
    .A(net3918),
    .Y(_06196_),
    .D(_04714_));
 sg13g2_xnor2_1 _12843_ (.Y(_06197_),
    .A(_06195_),
    .B(_06196_));
 sg13g2_a21oi_1 _12844_ (.A1(_01105_),
    .A2(net4482),
    .Y(_06198_),
    .B1(net4012));
 sg13g2_a21oi_1 _12845_ (.A1(net4012),
    .A2(_06197_),
    .Y(_06199_),
    .B1(_06198_));
 sg13g2_a21oi_1 _12846_ (.A1(\cpu.keccak_alu.registers[61] ),
    .A2(_06199_),
    .Y(_06200_),
    .B1(net4376));
 sg13g2_o21ai_1 _12847_ (.B1(_06200_),
    .Y(_06201_),
    .A1(\cpu.keccak_alu.registers[61] ),
    .A2(_06199_));
 sg13g2_a21oi_1 _12848_ (.A1(net4482),
    .A2(\cpu.keccak_alu.registers[253] ),
    .Y(_06202_),
    .B1(net4367));
 sg13g2_o21ai_1 _12849_ (.B1(_06202_),
    .Y(_06203_),
    .A1(net4482),
    .A2(\cpu.keccak_alu.registers[253] ));
 sg13g2_xnor2_1 _12850_ (.Y(_06204_),
    .A(\cpu.keccak_alu.registers[61] ),
    .B(\cpu.keccak_alu.registers[125] ));
 sg13g2_a21oi_1 _12851_ (.A1(_06203_),
    .A2(_06204_),
    .Y(_06205_),
    .B1(net4215));
 sg13g2_o21ai_1 _12852_ (.B1(_06205_),
    .Y(_06206_),
    .A1(_06203_),
    .A2(_06204_));
 sg13g2_a21oi_1 _12853_ (.A1(_06201_),
    .A2(_06206_),
    .Y(_06207_),
    .B1(net4313));
 sg13g2_o21ai_1 _12854_ (.B1(net3816),
    .Y(_06208_),
    .A1(net122),
    .A2(net3630));
 sg13g2_a21oi_1 _12855_ (.A1(net4276),
    .A2(net3630),
    .Y(_06209_),
    .B1(_06208_));
 sg13g2_nor3_1 _12856_ (.A(net3725),
    .B(_06207_),
    .C(_06209_),
    .Y(_06210_));
 sg13g2_a21oi_1 _12857_ (.A1(_01110_),
    .A2(net3722),
    .Y(_00778_),
    .B1(_06210_));
 sg13g2_o21ai_1 _12858_ (.B1(net4206),
    .Y(_06211_),
    .A1(\cpu.keccak_alu.registers[190] ),
    .A2(\cpu.keccak_alu.registers[254] ));
 sg13g2_a21oi_1 _12859_ (.A1(\cpu.keccak_alu.registers[190] ),
    .A2(\cpu.keccak_alu.registers[254] ),
    .Y(_06212_),
    .B1(_06211_));
 sg13g2_xor2_1 _12860_ (.B(\cpu.keccak_alu.registers[126] ),
    .A(\cpu.keccak_alu.registers[62] ),
    .X(_06213_));
 sg13g2_a21oi_1 _12861_ (.A1(_06212_),
    .A2(_06213_),
    .Y(_06214_),
    .B1(net4214));
 sg13g2_o21ai_1 _12862_ (.B1(_06214_),
    .Y(_06215_),
    .A1(_06212_),
    .A2(_06213_));
 sg13g2_nand3b_1 _12863_ (.B(\cpu.keccak_alu.registers[190] ),
    .C(net4000),
    .Y(_06216_),
    .A_N(\cpu.keccak_alu.registers[126] ));
 sg13g2_nor2_1 _12864_ (.A(_05972_),
    .B(_06030_),
    .Y(_06217_));
 sg13g2_o21ai_1 _12865_ (.B1(net4191),
    .Y(_06218_),
    .A1(_04173_),
    .A2(_04175_));
 sg13g2_o21ai_1 _12866_ (.B1(_06218_),
    .Y(_06219_),
    .A1(net4191),
    .A2(_06165_));
 sg13g2_mux2_1 _12867_ (.A0(_06118_),
    .A1(_06219_),
    .S(net4180),
    .X(_06220_));
 sg13g2_o21ai_1 _12868_ (.B1(net4091),
    .Y(_06221_),
    .A1(_05778_),
    .A2(_06220_));
 sg13g2_nor2_1 _12869_ (.A(_06217_),
    .B(_06221_),
    .Y(_06222_));
 sg13g2_nor2_1 _12870_ (.A(net3871),
    .B(_05834_),
    .Y(_06223_));
 sg13g2_nor3_1 _12871_ (.A(net4513),
    .B(_06222_),
    .C(_06223_),
    .Y(_06224_));
 sg13g2_o21ai_1 _12872_ (.B1(_06224_),
    .Y(_06225_),
    .A1(net4161),
    .A2(_05437_));
 sg13g2_nand2_1 _12873_ (.Y(_06226_),
    .A(net3772),
    .B(_05440_));
 sg13g2_xnor2_1 _12874_ (.Y(_06227_),
    .A(_06225_),
    .B(_06226_));
 sg13g2_o21ai_1 _12875_ (.B1(_06216_),
    .Y(_06228_),
    .A1(net4000),
    .A2(_06227_));
 sg13g2_xnor2_1 _12876_ (.Y(_06229_),
    .A(\cpu.keccak_alu.registers[62] ),
    .B(_06228_));
 sg13g2_o21ai_1 _12877_ (.B1(_06215_),
    .Y(_06230_),
    .A1(net4374),
    .A2(_06229_));
 sg13g2_nor2_1 _12878_ (.A(net166),
    .B(net3629),
    .Y(_06231_));
 sg13g2_a21oi_1 _12879_ (.A1(net4272),
    .A2(net3629),
    .Y(_06232_),
    .B1(_06231_));
 sg13g2_a221oi_1 _12880_ (.B2(net3817),
    .C1(net3723),
    .B1(_06232_),
    .A1(net4245),
    .Y(_06233_),
    .A2(_06230_));
 sg13g2_a21oi_1 _12881_ (.A1(_01125_),
    .A2(net3723),
    .Y(_00779_),
    .B1(_06233_));
 sg13g2_nor2b_1 _12882_ (.A(net3874),
    .B_N(_05858_),
    .Y(_06234_));
 sg13g2_nand2b_1 _12883_ (.Y(_06235_),
    .B(net4527),
    .A_N(_06048_));
 sg13g2_nand3_1 _12884_ (.B(net4191),
    .C(_00128_),
    .A(net4551),
    .Y(_06236_));
 sg13g2_a22oi_1 _12885_ (.Y(_06237_),
    .B1(_06189_),
    .B2(net4535),
    .A2(net4094),
    .A1(net4576));
 sg13g2_nand3_1 _12886_ (.B(_06236_),
    .C(_06237_),
    .A(net3827),
    .Y(_06238_));
 sg13g2_a221oi_1 _12887_ (.B2(_03865_),
    .C1(net3936),
    .B1(_06238_),
    .A1(_06093_),
    .Y(_06239_),
    .A2(_06144_));
 sg13g2_a221oi_1 _12888_ (.B2(_06239_),
    .C1(_06234_),
    .B1(_06235_),
    .A1(net4520),
    .Y(_06240_),
    .A2(_05465_));
 sg13g2_nor2_1 _12889_ (.A(net4516),
    .B(_06240_),
    .Y(_06241_));
 sg13g2_nand2_2 _12890_ (.Y(_06242_),
    .A(net3776),
    .B(_05469_));
 sg13g2_xor2_1 _12891_ (.B(_06242_),
    .A(_06241_),
    .X(_06243_));
 sg13g2_nand3b_1 _12892_ (.B(\cpu.keccak_alu.registers[191] ),
    .C(net4002),
    .Y(_06244_),
    .A_N(\cpu.keccak_alu.registers[127] ));
 sg13g2_o21ai_1 _12893_ (.B1(_06244_),
    .Y(_06245_),
    .A1(net4002),
    .A2(_06243_));
 sg13g2_xor2_1 _12894_ (.B(_06245_),
    .A(net949),
    .X(_06246_));
 sg13g2_o21ai_1 _12895_ (.B1(net4207),
    .Y(_06247_),
    .A1(\cpu.keccak_alu.registers[191] ),
    .A2(\cpu.keccak_alu.registers[255] ));
 sg13g2_a21oi_1 _12896_ (.A1(\cpu.keccak_alu.registers[191] ),
    .A2(\cpu.keccak_alu.registers[255] ),
    .Y(_06248_),
    .B1(_06247_));
 sg13g2_xnor2_1 _12897_ (.Y(_06249_),
    .A(\cpu.keccak_alu.registers[63] ),
    .B(\cpu.keccak_alu.registers[127] ));
 sg13g2_o21ai_1 _12898_ (.B1(net4376),
    .Y(_06250_),
    .A1(_06248_),
    .A2(_06249_));
 sg13g2_a21oi_1 _12899_ (.A1(_06248_),
    .A2(_06249_),
    .Y(_06251_),
    .B1(_06250_));
 sg13g2_nor2_1 _12900_ (.A(net4313),
    .B(_06251_),
    .Y(_06252_));
 sg13g2_o21ai_1 _12901_ (.B1(_06252_),
    .Y(_06253_),
    .A1(net4376),
    .A2(_06246_));
 sg13g2_o21ai_1 _12902_ (.B1(net3817),
    .Y(_06254_),
    .A1(net431),
    .A2(net3630));
 sg13g2_a21oi_1 _12903_ (.A1(net4269),
    .A2(net3630),
    .Y(_06255_),
    .B1(_06254_));
 sg13g2_nor2_1 _12904_ (.A(net3725),
    .B(_06255_),
    .Y(_06256_));
 sg13g2_a22oi_1 _12905_ (.Y(_00780_),
    .B1(_06253_),
    .B2(_06256_),
    .A2(net3724),
    .A1(_01138_));
 sg13g2_and3_2 _12906_ (.X(_06257_),
    .A(net4332),
    .B(_01301_),
    .C(_01318_));
 sg13g2_nand3_1 _12907_ (.B(_01301_),
    .C(_01318_),
    .A(net4332),
    .Y(_06258_));
 sg13g2_nor2_2 _12908_ (.A(_01302_),
    .B(_01306_),
    .Y(_06259_));
 sg13g2_and2_1 _12909_ (.A(_01301_),
    .B(_01310_),
    .X(_06260_));
 sg13g2_nand2_1 _12910_ (.Y(_06261_),
    .A(net4331),
    .B(_06260_));
 sg13g2_nand2b_1 _12911_ (.Y(_06262_),
    .B(_06261_),
    .A_N(_06259_));
 sg13g2_nor2_1 _12912_ (.A(_06257_),
    .B(net3769),
    .Y(_06263_));
 sg13g2_nor3_1 _12913_ (.A(net780),
    .B(_06257_),
    .C(net3769),
    .Y(_06264_));
 sg13g2_nor2_1 _12914_ (.A(_01302_),
    .B(_01313_),
    .Y(_06265_));
 sg13g2_or2_1 _12915_ (.X(_06266_),
    .B(_01313_),
    .A(_01302_));
 sg13g2_nor3_2 _12916_ (.A(\memory_controller.state[1] ),
    .B(net4333),
    .C(_01315_),
    .Y(_06267_));
 sg13g2_nand3_1 _12917_ (.B(_01305_),
    .C(_01307_),
    .A(\memory_controller.state[4] ),
    .Y(_06268_));
 sg13g2_nor2_2 _12918_ (.A(_01299_),
    .B(_01311_),
    .Y(_06269_));
 sg13g2_o21ai_1 _12919_ (.B1(_06268_),
    .Y(_06270_),
    .A1(_01299_),
    .A2(_01311_));
 sg13g2_nor4_1 _12920_ (.A(_03691_),
    .B(_06264_),
    .C(_06265_),
    .D(_06270_),
    .Y(_00781_));
 sg13g2_nand4_1 _12921_ (.B(\memory_controller.state[2] ),
    .C(net4331),
    .A(\memory_controller.state[3] ),
    .Y(_06271_),
    .D(_01307_));
 sg13g2_nand3_1 _12922_ (.B(_01301_),
    .C(_01318_),
    .A(net4331),
    .Y(_06272_));
 sg13g2_nand2_2 _12923_ (.Y(_06273_),
    .A(_06271_),
    .B(_06272_));
 sg13g2_nor2_2 _12924_ (.A(_01302_),
    .B(_01312_),
    .Y(_06274_));
 sg13g2_nor2_2 _12925_ (.A(_01299_),
    .B(_01319_),
    .Y(_06275_));
 sg13g2_nor4_1 _12926_ (.A(net893),
    .B(net3809),
    .C(_06274_),
    .D(net3808),
    .Y(_06276_));
 sg13g2_nand3_1 _12927_ (.B(_01305_),
    .C(_01310_),
    .A(net314),
    .Y(_06277_));
 sg13g2_nand2_2 _12928_ (.Y(_06278_),
    .A(_03692_),
    .B(_06277_));
 sg13g2_nor4_1 _12929_ (.A(_06257_),
    .B(_06270_),
    .C(_06276_),
    .D(_06278_),
    .Y(_00782_));
 sg13g2_nor2_1 _12930_ (.A(net4334),
    .B(_01317_),
    .Y(_06279_));
 sg13g2_nor2_1 _12931_ (.A(_01316_),
    .B(_06278_),
    .Y(_06280_));
 sg13g2_o21ai_1 _12932_ (.B1(net381),
    .Y(_06281_),
    .A1(_06279_),
    .A2(_06280_));
 sg13g2_nand3_1 _12933_ (.B(_06268_),
    .C(_06281_),
    .A(_06261_),
    .Y(_00783_));
 sg13g2_or3_1 _12934_ (.A(_06257_),
    .B(net3769),
    .C(_06270_),
    .X(_06282_));
 sg13g2_nor4_1 _12935_ (.A(_03691_),
    .B(net3809),
    .C(_06274_),
    .D(_06275_),
    .Y(_06283_));
 sg13g2_a21o_1 _12936_ (.A2(_06283_),
    .A1(net134),
    .B1(_06282_),
    .X(_00784_));
 sg13g2_nor2_1 _12937_ (.A(\memory_controller.state[0] ),
    .B(net1),
    .Y(_06284_));
 sg13g2_nor3_2 _12938_ (.A(_00891_),
    .B(_01313_),
    .C(_06284_),
    .Y(_06285_));
 sg13g2_nor2_2 _12939_ (.A(_03691_),
    .B(net3870),
    .Y(_06286_));
 sg13g2_a22oi_1 _12940_ (.Y(_06287_),
    .B1(_06286_),
    .B2(net73),
    .A2(net3870),
    .A1(net4));
 sg13g2_inv_1 _12941_ (.Y(_00785_),
    .A(_06287_));
 sg13g2_a22oi_1 _12942_ (.Y(_06288_),
    .B1(_06286_),
    .B2(net75),
    .A2(net3870),
    .A1(net5));
 sg13g2_inv_1 _12943_ (.Y(_00786_),
    .A(_06288_));
 sg13g2_a22oi_1 _12944_ (.Y(_06289_),
    .B1(_06286_),
    .B2(net52),
    .A2(net3870),
    .A1(net6));
 sg13g2_inv_1 _12945_ (.Y(_00787_),
    .A(_06289_));
 sg13g2_a22oi_1 _12946_ (.Y(_06290_),
    .B1(_06286_),
    .B2(net67),
    .A2(net3870),
    .A1(net7));
 sg13g2_inv_1 _12947_ (.Y(_00788_),
    .A(_06290_));
 sg13g2_a22oi_1 _12948_ (.Y(_06291_),
    .B1(_06286_),
    .B2(net54),
    .A2(net3870),
    .A1(net8));
 sg13g2_inv_1 _12949_ (.Y(_00789_),
    .A(_06291_));
 sg13g2_a22oi_1 _12950_ (.Y(_06292_),
    .B1(_06286_),
    .B2(net65),
    .A2(_06285_),
    .A1(net9));
 sg13g2_inv_1 _12951_ (.Y(_00790_),
    .A(net66));
 sg13g2_a22oi_1 _12952_ (.Y(_06293_),
    .B1(_06286_),
    .B2(net79),
    .A2(net3870),
    .A1(net10));
 sg13g2_inv_1 _12953_ (.Y(_00791_),
    .A(_06293_));
 sg13g2_a22oi_1 _12954_ (.Y(_06294_),
    .B1(_06286_),
    .B2(net91),
    .A2(net3870),
    .A1(net11));
 sg13g2_inv_1 _12955_ (.Y(_00792_),
    .A(_06294_));
 sg13g2_o21ai_1 _12956_ (.B1(_06277_),
    .Y(_00793_),
    .A1(net4202),
    .A2(_03691_));
 sg13g2_nor2_1 _12957_ (.A(net4331),
    .B(_01303_),
    .Y(_06295_));
 sg13g2_a21o_1 _12958_ (.A2(_03692_),
    .A1(net4322),
    .B1(_06295_),
    .X(_00794_));
 sg13g2_nand2_1 _12959_ (.Y(_06296_),
    .A(net890),
    .B(_06266_));
 sg13g2_o21ai_1 _12960_ (.B1(_06263_),
    .Y(_00795_),
    .A1(_06278_),
    .A2(_06296_));
 sg13g2_o21ai_1 _12961_ (.B1(_03692_),
    .Y(_06297_),
    .A1(net516),
    .A2(_06259_));
 sg13g2_nor2_1 _12962_ (.A(_06295_),
    .B(_06297_),
    .Y(_00796_));
 sg13g2_nor2b_2 _12963_ (.A(_06282_),
    .B_N(_06283_),
    .Y(_06298_));
 sg13g2_a22oi_1 _12964_ (.Y(_06299_),
    .B1(_06275_),
    .B2(net216),
    .A2(net3810),
    .A1(net339));
 sg13g2_and2_2 _12965_ (.A(\memory_controller.uart_memory_address[10] ),
    .B(_06274_),
    .X(_06300_));
 sg13g2_a21oi_1 _12966_ (.A1(net694),
    .A2(_06269_),
    .Y(_06301_),
    .B1(_06300_));
 sg13g2_a22oi_1 _12967_ (.Y(_06302_),
    .B1(net3809),
    .B2(\cpu.request_address[8] ),
    .A2(net3769),
    .A1(\cpu.request_address[0] ));
 sg13g2_nand2_1 _12968_ (.Y(_06303_),
    .A(net793),
    .B(_06298_));
 sg13g2_nand4_1 _12969_ (.B(_06301_),
    .C(_06302_),
    .A(_06299_),
    .Y(_00797_),
    .D(_06303_));
 sg13g2_a22oi_1 _12970_ (.Y(_06304_),
    .B1(net3808),
    .B2(net110),
    .A2(net3810),
    .A1(net139));
 sg13g2_a21oi_1 _12971_ (.A1(net393),
    .A2(_06269_),
    .Y(_06305_),
    .B1(_06300_));
 sg13g2_a22oi_1 _12972_ (.Y(_06306_),
    .B1(_06273_),
    .B2(\cpu.request_address[9] ),
    .A2(_06262_),
    .A1(\cpu.request_address[1] ));
 sg13g2_nand2_1 _12973_ (.Y(_06307_),
    .A(net720),
    .B(_06298_));
 sg13g2_nand4_1 _12974_ (.B(_06305_),
    .C(_06306_),
    .A(_06304_),
    .Y(_00798_),
    .D(_06307_));
 sg13g2_a22oi_1 _12975_ (.Y(_06308_),
    .B1(net3808),
    .B2(net74),
    .A2(_06269_),
    .A1(net111));
 sg13g2_a21oi_1 _12976_ (.A1(net197),
    .A2(net3810),
    .Y(_06309_),
    .B1(_06300_));
 sg13g2_a22oi_1 _12977_ (.Y(_06310_),
    .B1(net3809),
    .B2(net717),
    .A2(net3769),
    .A1(\cpu.request_address[2] ));
 sg13g2_nand2_1 _12978_ (.Y(_06311_),
    .A(net782),
    .B(_06298_));
 sg13g2_nand4_1 _12979_ (.B(_06309_),
    .C(_06310_),
    .A(_06308_),
    .Y(_00799_),
    .D(_06311_));
 sg13g2_a21oi_1 _12980_ (.A1(net87),
    .A2(_06275_),
    .Y(_06312_),
    .B1(_06300_));
 sg13g2_a22oi_1 _12981_ (.Y(_06313_),
    .B1(_06269_),
    .B2(net468),
    .A2(net3810),
    .A1(net190));
 sg13g2_a22oi_1 _12982_ (.Y(_06314_),
    .B1(_06273_),
    .B2(net584),
    .A2(_06262_),
    .A1(\cpu.request_address[3] ));
 sg13g2_nand2_1 _12983_ (.Y(_06315_),
    .A(net749),
    .B(_06298_));
 sg13g2_nand4_1 _12984_ (.B(_06313_),
    .C(_06314_),
    .A(_06312_),
    .Y(_00800_),
    .D(_06315_));
 sg13g2_a22oi_1 _12985_ (.Y(_06316_),
    .B1(net3808),
    .B2(net70),
    .A2(_06269_),
    .A1(net97));
 sg13g2_a21oi_1 _12986_ (.A1(net374),
    .A2(net3810),
    .Y(_06317_),
    .B1(_06300_));
 sg13g2_a22oi_1 _12987_ (.Y(_06318_),
    .B1(net3809),
    .B2(net611),
    .A2(_06262_),
    .A1(\cpu.request_address[4] ));
 sg13g2_nand2_1 _12988_ (.Y(_06319_),
    .A(net736),
    .B(_06298_));
 sg13g2_nand4_1 _12989_ (.B(_06317_),
    .C(_06318_),
    .A(_06316_),
    .Y(_00801_),
    .D(_06319_));
 sg13g2_and2_1 _12990_ (.A(\cpu.data_out[5] ),
    .B(_06269_),
    .X(_06320_));
 sg13g2_a21oi_1 _12991_ (.A1(\cpu.request_address[5] ),
    .A2(net3769),
    .Y(_06321_),
    .B1(_06300_));
 sg13g2_a221oi_1 _12992_ (.B2(net105),
    .C1(_06320_),
    .B1(net3808),
    .A1(\data_received[5] ),
    .Y(_06322_),
    .A2(net3810));
 sg13g2_a22oi_1 _12993_ (.Y(_06323_),
    .B1(net3809),
    .B2(\cpu.request_address[13] ),
    .A2(_06257_),
    .A1(\memory_controller.uart_memory_address[10] ));
 sg13g2_nand3_1 _12994_ (.B(_06322_),
    .C(_06323_),
    .A(_06321_),
    .Y(_06324_));
 sg13g2_mux2_1 _12995_ (.A0(_06324_),
    .A1(net777),
    .S(_06298_),
    .X(_00802_));
 sg13g2_a22oi_1 _12996_ (.Y(_06325_),
    .B1(_06269_),
    .B2(net186),
    .A2(net3810),
    .A1(net151));
 sg13g2_a21oi_1 _12997_ (.A1(net107),
    .A2(net3808),
    .Y(_06326_),
    .B1(_06300_));
 sg13g2_a22oi_1 _12998_ (.Y(_06327_),
    .B1(net3809),
    .B2(net805),
    .A2(net3769),
    .A1(\cpu.request_address[6] ));
 sg13g2_nand2_1 _12999_ (.Y(_06328_),
    .A(net810),
    .B(_06298_));
 sg13g2_nand4_1 _13000_ (.B(_06326_),
    .C(_06327_),
    .A(_06325_),
    .Y(_00803_),
    .D(_06328_));
 sg13g2_a22oi_1 _13001_ (.Y(_06329_),
    .B1(net3808),
    .B2(net76),
    .A2(net3810),
    .A1(net722));
 sg13g2_a22oi_1 _13002_ (.Y(_06330_),
    .B1(_06269_),
    .B2(net306),
    .A2(_06257_),
    .A1(net192));
 sg13g2_a22oi_1 _13003_ (.Y(_06331_),
    .B1(net3809),
    .B2(net357),
    .A2(net3769),
    .A1(\cpu.request_address[7] ));
 sg13g2_nand2_1 _13004_ (.Y(_06332_),
    .A(uio_out[7]),
    .B(_06298_));
 sg13g2_nand4_1 _13005_ (.B(_06330_),
    .C(_06331_),
    .A(_06329_),
    .Y(_00804_),
    .D(_06332_));
 sg13g2_mux2_1 _13006_ (.A0(\cpu.rx_speed[0] ),
    .A1(net258),
    .S(net4150),
    .X(_00805_));
 sg13g2_mux2_1 _13007_ (.A0(\cpu.rx_speed[1] ),
    .A1(net252),
    .S(net4150),
    .X(_00806_));
 sg13g2_mux2_1 _13008_ (.A0(\cpu.rx_speed[2] ),
    .A1(net245),
    .S(net4150),
    .X(_00807_));
 sg13g2_mux2_1 _13009_ (.A0(\cpu.rx_speed[3] ),
    .A1(net233),
    .S(net4150),
    .X(_00808_));
 sg13g2_mux2_1 _13010_ (.A0(\cpu.rx_speed[4] ),
    .A1(net214),
    .S(_01281_),
    .X(_00809_));
 sg13g2_mux2_1 _13011_ (.A0(net242),
    .A1(net305),
    .S(net4150),
    .X(_00810_));
 sg13g2_mux2_1 _13012_ (.A0(\cpu.rx_speed[6] ),
    .A1(net344),
    .S(net4150),
    .X(_00811_));
 sg13g2_mux2_1 _13013_ (.A0(\cpu.rx_speed[7] ),
    .A1(net212),
    .S(net4150),
    .X(_00812_));
 sg13g2_a221oi_1 _13014_ (.B2(_01337_),
    .C1(_02099_),
    .B1(_01927_),
    .A1(_01250_),
    .Y(_06333_),
    .A2(_01417_));
 sg13g2_nand2_1 _13015_ (.Y(_06334_),
    .A(_01431_),
    .B(_06333_));
 sg13g2_mux2_1 _13016_ (.A0(net4345),
    .A1(_00168_),
    .S(net3853),
    .X(_06335_));
 sg13g2_a21oi_1 _13017_ (.A1(net4054),
    .A2(_06335_),
    .Y(_06336_),
    .B1(net4260));
 sg13g2_nand2_1 _13018_ (.Y(_06337_),
    .A(_01596_),
    .B(_06336_));
 sg13g2_nor2_1 _13019_ (.A(net4234),
    .B(_06335_),
    .Y(_06338_));
 sg13g2_nor3_1 _13020_ (.A(_01601_),
    .B(net3540),
    .C(_06338_),
    .Y(_06339_));
 sg13g2_a22oi_1 _13021_ (.Y(_00813_),
    .B1(_06337_),
    .B2(_06339_),
    .A2(net3540),
    .A1(_00941_));
 sg13g2_nor2_1 _13022_ (.A(_00172_),
    .B(net3854),
    .Y(_06340_));
 sg13g2_a21oi_1 _13023_ (.A1(net4155),
    .A2(net3854),
    .Y(_06341_),
    .B1(_06340_));
 sg13g2_inv_1 _13024_ (.Y(_06342_),
    .A(_06341_));
 sg13g2_a21oi_1 _13025_ (.A1(net4056),
    .A2(_06341_),
    .Y(_06343_),
    .B1(net4262));
 sg13g2_a221oi_1 _13026_ (.B2(_01649_),
    .C1(net3540),
    .B1(_06343_),
    .A1(net4299),
    .Y(_06344_),
    .A2(_06342_));
 sg13g2_a22oi_1 _13027_ (.Y(_00814_),
    .B1(_06344_),
    .B2(_01654_),
    .A2(net3540),
    .A1(_00948_));
 sg13g2_mux2_1 _13028_ (.A0(net4338),
    .A1(_00176_),
    .S(net3853),
    .X(_06345_));
 sg13g2_a21oi_1 _13029_ (.A1(net4052),
    .A2(_06345_),
    .Y(_06346_),
    .B1(net4259));
 sg13g2_nand2_1 _13030_ (.Y(_06347_),
    .A(_01707_),
    .B(_06346_));
 sg13g2_nor2_1 _13031_ (.A(net4231),
    .B(_06345_),
    .Y(_06348_));
 sg13g2_nor3_1 _13032_ (.A(_01713_),
    .B(net3540),
    .C(_06348_),
    .Y(_06349_));
 sg13g2_a22oi_1 _13033_ (.Y(_00815_),
    .B1(_06347_),
    .B2(_06349_),
    .A2(net3540),
    .A1(_00956_));
 sg13g2_nor2_1 _13034_ (.A(net4297),
    .B(net3852),
    .Y(_06350_));
 sg13g2_a21oi_1 _13035_ (.A1(_01183_),
    .A2(net3852),
    .Y(_06351_),
    .B1(_06350_));
 sg13g2_a21oi_1 _13036_ (.A1(net4044),
    .A2(_06351_),
    .Y(_06352_),
    .B1(net4251));
 sg13g2_nand2_1 _13037_ (.Y(_06353_),
    .A(_01756_),
    .B(_06352_));
 sg13g2_nor2_1 _13038_ (.A(net4225),
    .B(_06351_),
    .Y(_06354_));
 sg13g2_nor3_1 _13039_ (.A(_01761_),
    .B(net3539),
    .C(_06354_),
    .Y(_06355_));
 sg13g2_a22oi_1 _13040_ (.Y(_00816_),
    .B1(_06353_),
    .B2(_06355_),
    .A2(net3539),
    .A1(_00963_));
 sg13g2_nand2_1 _13041_ (.Y(_06356_),
    .A(_00184_),
    .B(net3852));
 sg13g2_o21ai_1 _13042_ (.B1(_06356_),
    .Y(_06357_),
    .A1(net4154),
    .A2(net3852));
 sg13g2_a21oi_1 _13043_ (.A1(net4047),
    .A2(_06357_),
    .Y(_06358_),
    .B1(net4255));
 sg13g2_nand2_1 _13044_ (.Y(_06359_),
    .A(_01780_),
    .B(_06358_));
 sg13g2_nor2_1 _13045_ (.A(net4228),
    .B(_06357_),
    .Y(_06360_));
 sg13g2_nor3_1 _13046_ (.A(_01786_),
    .B(net3539),
    .C(_06360_),
    .Y(_06361_));
 sg13g2_a22oi_1 _13047_ (.Y(_00817_),
    .B1(_06359_),
    .B2(_06361_),
    .A2(net3539),
    .A1(_00971_));
 sg13g2_nor2_1 _13048_ (.A(_00188_),
    .B(net3855),
    .Y(_06362_));
 sg13g2_a21oi_1 _13049_ (.A1(net4153),
    .A2(net3855),
    .Y(_06363_),
    .B1(_06362_));
 sg13g2_a21oi_1 _13050_ (.A1(net4040),
    .A2(_06363_),
    .Y(_06364_),
    .B1(net4246));
 sg13g2_nand2_1 _13051_ (.Y(_06365_),
    .A(_01803_),
    .B(_06364_));
 sg13g2_nor2_1 _13052_ (.A(net4224),
    .B(_06363_),
    .Y(_06366_));
 sg13g2_nor3_1 _13053_ (.A(_01809_),
    .B(net3538),
    .C(_06366_),
    .Y(_06367_));
 sg13g2_a22oi_1 _13054_ (.Y(_00818_),
    .B1(_06365_),
    .B2(_06367_),
    .A2(net3538),
    .A1(_00979_));
 sg13g2_mux2_1 _13055_ (.A0(net4284),
    .A1(_00192_),
    .S(net3852),
    .X(_06368_));
 sg13g2_a21oi_1 _13056_ (.A1(net4046),
    .A2(_06368_),
    .Y(_06369_),
    .B1(net4252));
 sg13g2_nand2_1 _13057_ (.Y(_06370_),
    .A(_01826_),
    .B(_06369_));
 sg13g2_nor2_1 _13058_ (.A(net4229),
    .B(_06368_),
    .Y(_06371_));
 sg13g2_nor3_1 _13059_ (.A(_01831_),
    .B(net3540),
    .C(_06371_),
    .Y(_06372_));
 sg13g2_a22oi_1 _13060_ (.Y(_00819_),
    .B1(_06370_),
    .B2(_06372_),
    .A2(net3539),
    .A1(_00987_));
 sg13g2_mux2_1 _13061_ (.A0(net4280),
    .A1(_00196_),
    .S(net3852),
    .X(_06373_));
 sg13g2_a21oi_1 _13062_ (.A1(net4047),
    .A2(_06373_),
    .Y(_06374_),
    .B1(net4256));
 sg13g2_nand2_1 _13063_ (.Y(_06375_),
    .A(_01852_),
    .B(_06374_));
 sg13g2_nor2_1 _13064_ (.A(net4227),
    .B(_06373_),
    .Y(_06376_));
 sg13g2_nor3_1 _13065_ (.A(_01857_),
    .B(net3539),
    .C(_06376_),
    .Y(_06377_));
 sg13g2_a22oi_1 _13066_ (.Y(_00820_),
    .B1(_06375_),
    .B2(_06377_),
    .A2(net3539),
    .A1(_00995_));
 sg13g2_nor2_1 _13067_ (.A(_00200_),
    .B(net3855),
    .Y(_06378_));
 sg13g2_a21oi_1 _13068_ (.A1(net4152),
    .A2(net3855),
    .Y(_06379_),
    .B1(_06378_));
 sg13g2_a21oi_1 _13069_ (.A1(net4042),
    .A2(_06379_),
    .Y(_06380_),
    .B1(net4247));
 sg13g2_nand2_1 _13070_ (.Y(_06381_),
    .A(_01871_),
    .B(_06380_));
 sg13g2_nor2_1 _13071_ (.A(net4223),
    .B(_06379_),
    .Y(_06382_));
 sg13g2_nor3_1 _13072_ (.A(_01877_),
    .B(net3538),
    .C(_06382_),
    .Y(_06383_));
 sg13g2_a22oi_1 _13073_ (.Y(_00821_),
    .B1(_06381_),
    .B2(_06383_),
    .A2(net3538),
    .A1(_01117_));
 sg13g2_nor2_1 _13074_ (.A(_00205_),
    .B(net3855),
    .Y(_06384_));
 sg13g2_a21oi_1 _13075_ (.A1(net4151),
    .A2(net3855),
    .Y(_06385_),
    .B1(_06384_));
 sg13g2_a21oi_1 _13076_ (.A1(net4040),
    .A2(_06385_),
    .Y(_06386_),
    .B1(net4247));
 sg13g2_nand2_1 _13077_ (.Y(_06387_),
    .A(_01892_),
    .B(_06386_));
 sg13g2_nor2_1 _13078_ (.A(net4221),
    .B(_06385_),
    .Y(_06388_));
 sg13g2_nor3_1 _13079_ (.A(_01898_),
    .B(net3538),
    .C(_06388_),
    .Y(_06389_));
 sg13g2_a22oi_1 _13080_ (.Y(_00822_),
    .B1(_06387_),
    .B2(_06389_),
    .A2(net3538),
    .A1(_01132_));
 sg13g2_mux2_1 _13081_ (.A0(net4268),
    .A1(_00209_),
    .S(net3852),
    .X(_06390_));
 sg13g2_a21oi_1 _13082_ (.A1(net4042),
    .A2(_06390_),
    .Y(_06391_),
    .B1(net4249));
 sg13g2_nand2_1 _13083_ (.Y(_06392_),
    .A(_01912_),
    .B(_06391_));
 sg13g2_nor2_1 _13084_ (.A(net4223),
    .B(_06390_),
    .Y(_06393_));
 sg13g2_nor3_1 _13085_ (.A(_01917_),
    .B(net3538),
    .C(_06393_),
    .Y(_06394_));
 sg13g2_a22oi_1 _13086_ (.Y(_00823_),
    .B1(_06392_),
    .B2(_06394_),
    .A2(net3538),
    .A1(_01145_));
 sg13g2_nor2b_2 _13087_ (.A(net946),
    .B_N(_06260_),
    .Y(_06395_));
 sg13g2_nor2_2 _13088_ (.A(_03691_),
    .B(_06395_),
    .Y(_06396_));
 sg13g2_a22oi_1 _13089_ (.Y(_06397_),
    .B1(_06396_),
    .B2(net61),
    .A2(net3807),
    .A1(net4));
 sg13g2_inv_1 _13090_ (.Y(_00824_),
    .A(_06397_));
 sg13g2_a22oi_1 _13091_ (.Y(_06398_),
    .B1(_06396_),
    .B2(net53),
    .A2(net3807),
    .A1(net5));
 sg13g2_inv_1 _13092_ (.Y(_00825_),
    .A(_06398_));
 sg13g2_a22oi_1 _13093_ (.Y(_06399_),
    .B1(_06396_),
    .B2(net71),
    .A2(net3807),
    .A1(net6));
 sg13g2_inv_1 _13094_ (.Y(_00826_),
    .A(_06399_));
 sg13g2_a22oi_1 _13095_ (.Y(_06400_),
    .B1(_06396_),
    .B2(net64),
    .A2(net3807),
    .A1(net7));
 sg13g2_inv_1 _13096_ (.Y(_00827_),
    .A(_06400_));
 sg13g2_a22oi_1 _13097_ (.Y(_06401_),
    .B1(_06396_),
    .B2(net120),
    .A2(net3807),
    .A1(net8));
 sg13g2_inv_1 _13098_ (.Y(_00828_),
    .A(_06401_));
 sg13g2_a22oi_1 _13099_ (.Y(_06402_),
    .B1(_06396_),
    .B2(net78),
    .A2(net3807),
    .A1(net9));
 sg13g2_inv_1 _13100_ (.Y(_00829_),
    .A(_06402_));
 sg13g2_a22oi_1 _13101_ (.Y(_06403_),
    .B1(_06396_),
    .B2(net241),
    .A2(net3807),
    .A1(net10));
 sg13g2_inv_1 _13102_ (.Y(_00830_),
    .A(_06403_));
 sg13g2_a22oi_1 _13103_ (.Y(_06404_),
    .B1(_06396_),
    .B2(net92),
    .A2(net3807),
    .A1(net11));
 sg13g2_inv_1 _13104_ (.Y(_00831_),
    .A(_06404_));
 sg13g2_nand2_1 _13105_ (.Y(_06405_),
    .A(\memory_controller.state[4] ),
    .B(_03690_));
 sg13g2_o21ai_1 _13106_ (.B1(_06405_),
    .Y(_06406_),
    .A1(_01313_),
    .A2(_01319_));
 sg13g2_nor3_1 _13107_ (.A(_06274_),
    .B(_06395_),
    .C(_06406_),
    .Y(_06407_));
 sg13g2_o21ai_1 _13108_ (.B1(_06258_),
    .Y(_06408_),
    .A1(_01311_),
    .A2(_01312_));
 sg13g2_nand4_1 _13109_ (.B(_01321_),
    .C(_06268_),
    .A(net4634),
    .Y(_06409_),
    .D(_06407_));
 sg13g2_nor2_1 _13110_ (.A(_06408_),
    .B(_06409_),
    .Y(_06410_));
 sg13g2_a22oi_1 _13111_ (.Y(_00832_),
    .B1(_03693_),
    .B2(_06410_),
    .A2(_01192_),
    .A1(net4580));
 sg13g2_nor3_2 _13112_ (.A(_00898_),
    .B(net211),
    .C(_03692_),
    .Y(_06411_));
 sg13g2_nand2b_1 _13113_ (.Y(_06412_),
    .B(_06411_),
    .A_N(\cpu.uart_inbound ));
 sg13g2_nor2_1 _13114_ (.A(_01313_),
    .B(_01318_),
    .Y(_06413_));
 sg13g2_nor4_2 _13115_ (.A(\memory_controller.wait_counter[3] ),
    .B(net174),
    .C(\memory_controller.wait_counter[5] ),
    .Y(_06414_),
    .D(net947));
 sg13g2_inv_1 _13116_ (.Y(_06415_),
    .A(_06414_));
 sg13g2_a21oi_1 _13117_ (.A1(_01320_),
    .A2(_06415_),
    .Y(_06416_),
    .B1(_01308_));
 sg13g2_nor3_2 _13118_ (.A(_06259_),
    .B(_06267_),
    .C(_06279_),
    .Y(_06417_));
 sg13g2_nand3_1 _13119_ (.B(_06416_),
    .C(_06417_),
    .A(net4633),
    .Y(_06418_));
 sg13g2_nor4_1 _13120_ (.A(_01322_),
    .B(net3808),
    .C(_06413_),
    .D(_06418_),
    .Y(_06419_));
 sg13g2_a22oi_1 _13121_ (.Y(_00833_),
    .B1(_06412_),
    .B2(_06419_),
    .A2(_01193_),
    .A1(net4580));
 sg13g2_a21oi_2 _13122_ (.B1(_06274_),
    .Y(_06420_),
    .A2(net175),
    .A1(_01320_));
 sg13g2_nand3_1 _13123_ (.B(net4331),
    .C(_01319_),
    .A(\memory_controller.state[2] ),
    .Y(_06421_));
 sg13g2_nand3_1 _13124_ (.B(_06272_),
    .C(_06421_),
    .A(net4633),
    .Y(_06422_));
 sg13g2_nor3_1 _13125_ (.A(_01306_),
    .B(_01319_),
    .C(_06414_),
    .Y(_06423_));
 sg13g2_nor3_1 _13126_ (.A(_06408_),
    .B(_06422_),
    .C(_06423_),
    .Y(_06424_));
 sg13g2_a22oi_1 _13127_ (.Y(_00834_),
    .B1(_06420_),
    .B2(_06424_),
    .A2(_01194_),
    .A1(net4580));
 sg13g2_and2_1 _13128_ (.A(_01314_),
    .B(_06415_),
    .X(_06425_));
 sg13g2_a22oi_1 _13129_ (.Y(_06426_),
    .B1(_06414_),
    .B2(_01322_),
    .A2(_03691_),
    .A1(\cpu.uart_inbound ));
 sg13g2_nor3_1 _13130_ (.A(_01299_),
    .B(_01307_),
    .C(_01318_),
    .Y(_06427_));
 sg13g2_o21ai_1 _13131_ (.B1(_06266_),
    .Y(_06428_),
    .A1(_00020_),
    .A2(_01317_));
 sg13g2_nor4_1 _13132_ (.A(net4580),
    .B(_01304_),
    .C(_06259_),
    .D(_06260_),
    .Y(_06429_));
 sg13g2_nor4_1 _13133_ (.A(_06411_),
    .B(_06425_),
    .C(_06427_),
    .D(_06428_),
    .Y(_06430_));
 sg13g2_nand4_1 _13134_ (.B(_06426_),
    .C(_06429_),
    .A(_06420_),
    .Y(_06431_),
    .D(_06430_));
 sg13g2_o21ai_1 _13135_ (.B1(_06431_),
    .Y(_06432_),
    .A1(net4629),
    .A2(net19));
 sg13g2_inv_1 _13136_ (.Y(_00835_),
    .A(_06432_));
 sg13g2_nand3_1 _13137_ (.B(\cpu.request_type ),
    .C(_03691_),
    .A(\cpu.request ),
    .Y(_06433_));
 sg13g2_nand2_1 _13138_ (.Y(_06434_),
    .A(_01314_),
    .B(_06414_));
 sg13g2_nand2_1 _13139_ (.Y(_06435_),
    .A(net1),
    .B(_06265_));
 sg13g2_nand4_1 _13140_ (.B(net81),
    .C(_06434_),
    .A(_06426_),
    .Y(_06436_),
    .D(_06435_));
 sg13g2_nor2_1 _13141_ (.A(_01309_),
    .B(net948),
    .Y(_06437_));
 sg13g2_nand2_1 _13142_ (.Y(_06438_),
    .A(_06417_),
    .B(_06420_));
 sg13g2_nand3_1 _13143_ (.B(net2),
    .C(_03690_),
    .A(net4332),
    .Y(_06439_));
 sg13g2_nand4_1 _13144_ (.B(_06258_),
    .C(_06271_),
    .A(net4633),
    .Y(_06440_),
    .D(_06439_));
 sg13g2_nor4_1 _13145_ (.A(_06436_),
    .B(_06437_),
    .C(_06438_),
    .D(_06440_),
    .Y(_06441_));
 sg13g2_a21oi_1 _13146_ (.A1(net4579),
    .A2(_01195_),
    .Y(_00836_),
    .B1(_06441_));
 sg13g2_nor2b_1 _13147_ (.A(\cpu.uart.send ),
    .B_N(\cpu.uart.stage[0] ),
    .Y(_06442_));
 sg13g2_a21oi_1 _13148_ (.A1(\cpu.uart.stage[1] ),
    .A2(_01219_),
    .Y(_06443_),
    .B1(_06442_));
 sg13g2_or2_1 _13149_ (.X(_06444_),
    .B(net30),
    .A(\cpu.uart.stage[1] ));
 sg13g2_nand3_1 _13150_ (.B(_06443_),
    .C(_06444_),
    .A(net588),
    .Y(_06445_));
 sg13g2_nor3_1 _13151_ (.A(_00007_),
    .B(_01219_),
    .C(_01222_),
    .Y(_06446_));
 sg13g2_o21ai_1 _13152_ (.B1(net342),
    .Y(_06447_),
    .A1(_06445_),
    .A2(_06446_));
 sg13g2_o21ai_1 _13153_ (.B1(_06447_),
    .Y(_00837_),
    .A1(_00905_),
    .A2(_06445_));
 sg13g2_nand3_1 _13154_ (.B(net4368),
    .C(net4396),
    .A(net4376),
    .Y(_06448_));
 sg13g2_inv_1 _13155_ (.Y(_06449_),
    .A(net4088));
 sg13g2_nand2_1 _13156_ (.Y(_06450_),
    .A(_00243_),
    .B(net4088));
 sg13g2_a21oi_1 _13157_ (.A1(net4365),
    .A2(_06449_),
    .Y(_06451_),
    .B1(_01410_));
 sg13g2_nand2_1 _13158_ (.Y(_06452_),
    .A(_01420_),
    .B(net4088));
 sg13g2_nand3_1 _13159_ (.B(\cpu.current_instruction[6] ),
    .C(net4445),
    .A(net4448),
    .Y(_06453_));
 sg13g2_a22oi_1 _13160_ (.Y(_06454_),
    .B1(_06453_),
    .B2(_01927_),
    .A2(net3986),
    .A1(_01926_));
 sg13g2_nand4_1 _13161_ (.B(_01432_),
    .C(_06452_),
    .A(_01423_),
    .Y(_06455_),
    .D(_06454_));
 sg13g2_a21oi_1 _13162_ (.A1(_06450_),
    .A2(_06451_),
    .Y(_06456_),
    .B1(_01442_));
 sg13g2_nand2_1 _13163_ (.Y(_06457_),
    .A(net347),
    .B(net3546));
 sg13g2_o21ai_1 _13164_ (.B1(_06457_),
    .Y(_00838_),
    .A1(net3546),
    .A2(_06456_));
 sg13g2_mux2_1 _13165_ (.A0(net4361),
    .A1(_00031_),
    .S(net4088),
    .X(_06458_));
 sg13g2_nor2_1 _13166_ (.A(_01451_),
    .B(_06458_),
    .Y(_06459_));
 sg13g2_nor3_1 _13167_ (.A(_01448_),
    .B(net3546),
    .C(_06459_),
    .Y(_06460_));
 sg13g2_a21oi_1 _13168_ (.A1(_00908_),
    .A2(net3547),
    .Y(_00839_),
    .B1(_06460_));
 sg13g2_and2_1 _13169_ (.A(_00032_),
    .B(net4088),
    .X(_06461_));
 sg13g2_a221oi_1 _13170_ (.B2(net4353),
    .C1(_06461_),
    .B1(_06449_),
    .A1(net4231),
    .Y(_06462_),
    .A2(_01476_));
 sg13g2_nor3_1 _13171_ (.A(_01481_),
    .B(net3546),
    .C(_06462_),
    .Y(_06463_));
 sg13g2_a21oi_1 _13172_ (.A1(_00913_),
    .A2(net3546),
    .Y(_00840_),
    .B1(_06463_));
 sg13g2_nor2_1 _13173_ (.A(net4351),
    .B(net4087),
    .Y(_06464_));
 sg13g2_a21oi_1 _13174_ (.A1(_00921_),
    .A2(net4087),
    .Y(_06465_),
    .B1(_06464_));
 sg13g2_a21oi_1 _13175_ (.A1(net4057),
    .A2(_06465_),
    .Y(_06466_),
    .B1(_01512_));
 sg13g2_nor2_1 _13176_ (.A(net4235),
    .B(_06465_),
    .Y(_06467_));
 sg13g2_nor4_1 _13177_ (.A(_01516_),
    .B(net3545),
    .C(_06466_),
    .D(_06467_),
    .Y(_06468_));
 sg13g2_a21oi_1 _13178_ (.A1(_00920_),
    .A2(net3545),
    .Y(_00841_),
    .B1(_06468_));
 sg13g2_nor2_1 _13179_ (.A(net4348),
    .B(net4087),
    .Y(_06469_));
 sg13g2_a21oi_1 _13180_ (.A1(_00928_),
    .A2(net4087),
    .Y(_06470_),
    .B1(_06469_));
 sg13g2_a21oi_1 _13181_ (.A1(net4057),
    .A2(_06470_),
    .Y(_06471_),
    .B1(_01552_));
 sg13g2_nand2b_1 _13182_ (.Y(_06472_),
    .B(net4299),
    .A_N(_06470_));
 sg13g2_nor3_1 _13183_ (.A(_01556_),
    .B(net3545),
    .C(_06471_),
    .Y(_06473_));
 sg13g2_a22oi_1 _13184_ (.Y(_00842_),
    .B1(_06472_),
    .B2(_06473_),
    .A2(net3545),
    .A1(_00927_));
 sg13g2_nor2_1 _13185_ (.A(net4345),
    .B(net4087),
    .Y(_06474_));
 sg13g2_a21oi_1 _13186_ (.A1(_00935_),
    .A2(net4087),
    .Y(_06475_),
    .B1(_06474_));
 sg13g2_a21oi_1 _13187_ (.A1(net4054),
    .A2(_06475_),
    .Y(_06476_),
    .B1(net4260));
 sg13g2_nand2_1 _13188_ (.Y(_06477_),
    .A(_01596_),
    .B(_06476_));
 sg13g2_nor2_1 _13189_ (.A(net4234),
    .B(_06475_),
    .Y(_06478_));
 sg13g2_nor3_1 _13190_ (.A(_01601_),
    .B(net3545),
    .C(_06478_),
    .Y(_06479_));
 sg13g2_a22oi_1 _13191_ (.Y(_00843_),
    .B1(_06477_),
    .B2(_06479_),
    .A2(net3545),
    .A1(_00934_));
 sg13g2_nand2_1 _13192_ (.Y(_06480_),
    .A(_00036_),
    .B(net4087));
 sg13g2_o21ai_1 _13193_ (.B1(_06480_),
    .Y(_06481_),
    .A1(net4155),
    .A2(net4087));
 sg13g2_inv_1 _13194_ (.Y(_06482_),
    .A(_06481_));
 sg13g2_a21oi_1 _13195_ (.A1(net4056),
    .A2(_06481_),
    .Y(_06483_),
    .B1(net4262));
 sg13g2_a221oi_1 _13196_ (.B2(_01649_),
    .C1(net3545),
    .B1(_06483_),
    .A1(net4299),
    .Y(_06484_),
    .A2(_06482_));
 sg13g2_a22oi_1 _13197_ (.Y(_00844_),
    .B1(_06484_),
    .B2(_01654_),
    .A2(net3545),
    .A1(_00942_));
 sg13g2_nor2_1 _13198_ (.A(net4338),
    .B(net4088),
    .Y(_06485_));
 sg13g2_a21oi_1 _13199_ (.A1(_00950_),
    .A2(net4088),
    .Y(_06486_),
    .B1(_06485_));
 sg13g2_a21oi_1 _13200_ (.A1(net4054),
    .A2(_06486_),
    .Y(_06487_),
    .B1(net4259));
 sg13g2_nand2_1 _13201_ (.Y(_06488_),
    .A(_01707_),
    .B(_06487_));
 sg13g2_nor2_1 _13202_ (.A(net4234),
    .B(_06486_),
    .Y(_06489_));
 sg13g2_nor3_1 _13203_ (.A(_01713_),
    .B(net3546),
    .C(_06489_),
    .Y(_06490_));
 sg13g2_a22oi_1 _13204_ (.Y(_00845_),
    .B1(_06488_),
    .B2(_06490_),
    .A2(net3546),
    .A1(_00949_));
 sg13g2_mux2_1 _13205_ (.A0(net4297),
    .A1(_00038_),
    .S(net4085),
    .X(_06491_));
 sg13g2_a21oi_1 _13206_ (.A1(net4045),
    .A2(_06491_),
    .Y(_06492_),
    .B1(net4251));
 sg13g2_nand2_1 _13207_ (.Y(_06493_),
    .A(_01756_),
    .B(_06492_));
 sg13g2_nor2_1 _13208_ (.A(net4226),
    .B(_06491_),
    .Y(_06494_));
 sg13g2_nor3_1 _13209_ (.A(_01761_),
    .B(net3544),
    .C(_06494_),
    .Y(_06495_));
 sg13g2_a22oi_1 _13210_ (.Y(_00846_),
    .B1(_06493_),
    .B2(_06495_),
    .A2(net3544),
    .A1(_00957_));
 sg13g2_nor2_1 _13211_ (.A(net4293),
    .B(net4086),
    .Y(_06496_));
 sg13g2_a21oi_1 _13212_ (.A1(_00965_),
    .A2(net4086),
    .Y(_06497_),
    .B1(_06496_));
 sg13g2_a21oi_1 _13213_ (.A1(net4048),
    .A2(_06497_),
    .Y(_06498_),
    .B1(net4255));
 sg13g2_nand2_1 _13214_ (.Y(_06499_),
    .A(_01780_),
    .B(_06498_));
 sg13g2_nor2_1 _13215_ (.A(net4227),
    .B(_06497_),
    .Y(_06500_));
 sg13g2_nor3_1 _13216_ (.A(_01786_),
    .B(net3544),
    .C(_06500_),
    .Y(_06501_));
 sg13g2_a22oi_1 _13217_ (.Y(_00847_),
    .B1(_06499_),
    .B2(_06501_),
    .A2(net3544),
    .A1(_00964_));
 sg13g2_nor2_1 _13218_ (.A(net4289),
    .B(net4085),
    .Y(_06502_));
 sg13g2_a21oi_1 _13219_ (.A1(_00973_),
    .A2(net4085),
    .Y(_06503_),
    .B1(_06502_));
 sg13g2_a21oi_1 _13220_ (.A1(net4044),
    .A2(_06503_),
    .Y(_06504_),
    .B1(net4250));
 sg13g2_nand2_1 _13221_ (.Y(_06505_),
    .A(_01803_),
    .B(_06504_));
 sg13g2_nor2_1 _13222_ (.A(net4225),
    .B(_06503_),
    .Y(_06506_));
 sg13g2_nor3_1 _13223_ (.A(_01809_),
    .B(net3543),
    .C(_06506_),
    .Y(_06507_));
 sg13g2_a22oi_1 _13224_ (.Y(_00848_),
    .B1(_06505_),
    .B2(_06507_),
    .A2(net3543),
    .A1(_00972_));
 sg13g2_nor2_1 _13225_ (.A(net4284),
    .B(net4086),
    .Y(_06508_));
 sg13g2_a21oi_1 _13226_ (.A1(_00981_),
    .A2(net4086),
    .Y(_06509_),
    .B1(_06508_));
 sg13g2_a21oi_1 _13227_ (.A1(net4046),
    .A2(_06509_),
    .Y(_06510_),
    .B1(net4252));
 sg13g2_nand2_1 _13228_ (.Y(_06511_),
    .A(_01826_),
    .B(_06510_));
 sg13g2_nor2_1 _13229_ (.A(net4229),
    .B(_06509_),
    .Y(_06512_));
 sg13g2_nor3_1 _13230_ (.A(_01831_),
    .B(net3544),
    .C(_06512_),
    .Y(_06513_));
 sg13g2_a22oi_1 _13231_ (.Y(_00849_),
    .B1(_06511_),
    .B2(_06513_),
    .A2(net3544),
    .A1(_00980_));
 sg13g2_nor2_1 _13232_ (.A(net4280),
    .B(net4086),
    .Y(_06514_));
 sg13g2_a21oi_1 _13233_ (.A1(_00989_),
    .A2(net4086),
    .Y(_06515_),
    .B1(_06514_));
 sg13g2_a21oi_1 _13234_ (.A1(net4047),
    .A2(_06515_),
    .Y(_06516_),
    .B1(net4255));
 sg13g2_nand2_1 _13235_ (.Y(_06517_),
    .A(_01852_),
    .B(_06516_));
 sg13g2_nor2_1 _13236_ (.A(net4227),
    .B(_06515_),
    .Y(_06518_));
 sg13g2_nor3_1 _13237_ (.A(_01857_),
    .B(net3547),
    .C(_06518_),
    .Y(_06519_));
 sg13g2_a22oi_1 _13238_ (.Y(_00850_),
    .B1(_06517_),
    .B2(_06519_),
    .A2(net3544),
    .A1(_00988_));
 sg13g2_nand2_1 _13239_ (.Y(_06520_),
    .A(_00046_),
    .B(net4085));
 sg13g2_o21ai_1 _13240_ (.B1(_06520_),
    .Y(_06521_),
    .A1(net4152),
    .A2(net4085));
 sg13g2_a21oi_1 _13241_ (.A1(net4041),
    .A2(_06521_),
    .Y(_06522_),
    .B1(net4247));
 sg13g2_nand2_1 _13242_ (.Y(_06523_),
    .A(_01871_),
    .B(_06522_));
 sg13g2_nor2_1 _13243_ (.A(net4222),
    .B(_06521_),
    .Y(_06524_));
 sg13g2_nor3_1 _13244_ (.A(_01877_),
    .B(net3543),
    .C(_06524_),
    .Y(_06525_));
 sg13g2_a22oi_1 _13245_ (.Y(_00851_),
    .B1(_06523_),
    .B2(_06525_),
    .A2(net3543),
    .A1(_01111_));
 sg13g2_nand2_1 _13246_ (.Y(_06526_),
    .A(_00047_),
    .B(net4085));
 sg13g2_o21ai_1 _13247_ (.B1(_06526_),
    .Y(_06527_),
    .A1(net4151),
    .A2(net4085));
 sg13g2_a21oi_1 _13248_ (.A1(net4040),
    .A2(_06527_),
    .Y(_06528_),
    .B1(net4247));
 sg13g2_nand2_1 _13249_ (.Y(_06529_),
    .A(_01892_),
    .B(_06528_));
 sg13g2_nor2_1 _13250_ (.A(net4221),
    .B(_06527_),
    .Y(_06530_));
 sg13g2_nor3_1 _13251_ (.A(_01898_),
    .B(net3543),
    .C(_06530_),
    .Y(_06531_));
 sg13g2_a22oi_1 _13252_ (.Y(_00852_),
    .B1(_06529_),
    .B2(_06531_),
    .A2(net3543),
    .A1(_01126_));
 sg13g2_mux2_1 _13253_ (.A0(net4268),
    .A1(_00048_),
    .S(net4085),
    .X(_06532_));
 sg13g2_a21oi_1 _13254_ (.A1(net4041),
    .A2(_06532_),
    .Y(_06533_),
    .B1(net4248));
 sg13g2_nand2_1 _13255_ (.Y(_06534_),
    .A(_01912_),
    .B(_06533_));
 sg13g2_nor2_1 _13256_ (.A(net4222),
    .B(_06532_),
    .Y(_06535_));
 sg13g2_nor3_1 _13257_ (.A(_01917_),
    .B(net3543),
    .C(_06535_),
    .Y(_06536_));
 sg13g2_a22oi_1 _13258_ (.Y(_00853_),
    .B1(_06534_),
    .B2(_06536_),
    .A2(net3543),
    .A1(_01139_));
 sg13g2_nor2_1 _13259_ (.A(\cpu.uart.stage[2] ),
    .B(_06444_),
    .Y(_06537_));
 sg13g2_nor3_2 _13260_ (.A(net4477),
    .B(_06442_),
    .C(_06537_),
    .Y(_06538_));
 sg13g2_a21oi_1 _13261_ (.A1(\cpu.uart.stage[2] ),
    .A2(_01219_),
    .Y(_06539_),
    .B1(_06537_));
 sg13g2_and2_1 _13262_ (.A(_06443_),
    .B(_06539_),
    .X(_06540_));
 sg13g2_nand2_1 _13263_ (.Y(_06541_),
    .A(_06443_),
    .B(_06539_));
 sg13g2_a21oi_1 _13264_ (.A1(_06538_),
    .A2(_06541_),
    .Y(_06542_),
    .B1(net391));
 sg13g2_a21oi_1 _13265_ (.A1(net391),
    .A2(_06538_),
    .Y(_00854_),
    .B1(_06542_));
 sg13g2_o21ai_1 _13266_ (.B1(_01219_),
    .Y(_06543_),
    .A1(\cpu.uart.stage[1] ),
    .A2(\cpu.uart.stage[2] ));
 sg13g2_and2_1 _13267_ (.A(_06538_),
    .B(_06543_),
    .X(_06544_));
 sg13g2_a21oi_1 _13268_ (.A1(\cpu.uart.cycle_counter[0] ),
    .A2(_06538_),
    .Y(_06545_),
    .B1(net264));
 sg13g2_and3_1 _13269_ (.X(_06546_),
    .A(net391),
    .B(net264),
    .C(_06538_));
 sg13g2_nor3_1 _13270_ (.A(net3628),
    .B(net265),
    .C(_06546_),
    .Y(_00855_));
 sg13g2_xnor2_1 _13271_ (.Y(_06547_),
    .A(net724),
    .B(_06546_));
 sg13g2_nor2_1 _13272_ (.A(net3628),
    .B(_06547_),
    .Y(_00856_));
 sg13g2_and3_1 _13273_ (.X(_06548_),
    .A(\cpu.uart.cycle_counter[2] ),
    .B(net117),
    .C(_06546_));
 sg13g2_a21oi_1 _13274_ (.A1(\cpu.uart.cycle_counter[2] ),
    .A2(_06546_),
    .Y(_06549_),
    .B1(net117));
 sg13g2_nor3_1 _13275_ (.A(net3628),
    .B(_06548_),
    .C(net118),
    .Y(_00857_));
 sg13g2_nor2_1 _13276_ (.A(net506),
    .B(_06548_),
    .Y(_06550_));
 sg13g2_and2_1 _13277_ (.A(net506),
    .B(_06548_),
    .X(_06551_));
 sg13g2_nor3_1 _13278_ (.A(net3628),
    .B(net507),
    .C(_06551_),
    .Y(_00858_));
 sg13g2_nor2_1 _13279_ (.A(net456),
    .B(_06551_),
    .Y(_06552_));
 sg13g2_and2_1 _13280_ (.A(net456),
    .B(_06551_),
    .X(_06553_));
 sg13g2_nor3_1 _13281_ (.A(net3627),
    .B(net457),
    .C(_06553_),
    .Y(_00859_));
 sg13g2_xnor2_1 _13282_ (.Y(_06554_),
    .A(net738),
    .B(_06553_));
 sg13g2_nor2_1 _13283_ (.A(net3627),
    .B(_06554_),
    .Y(_00860_));
 sg13g2_a21oi_1 _13284_ (.A1(\cpu.uart.cycle_counter[6] ),
    .A2(_06553_),
    .Y(_06555_),
    .B1(net113));
 sg13g2_and3_1 _13285_ (.X(_06556_),
    .A(\cpu.uart.cycle_counter[6] ),
    .B(net113),
    .C(_06553_));
 sg13g2_nor3_1 _13286_ (.A(net3627),
    .B(net114),
    .C(_06556_),
    .Y(_00861_));
 sg13g2_xnor2_1 _13287_ (.Y(_06557_),
    .A(net679),
    .B(_06556_));
 sg13g2_nor2_1 _13288_ (.A(net3627),
    .B(net680),
    .Y(_00862_));
 sg13g2_a21oi_1 _13289_ (.A1(\cpu.uart.cycle_counter[8] ),
    .A2(_06556_),
    .Y(_06558_),
    .B1(net278));
 sg13g2_and3_1 _13290_ (.X(_06559_),
    .A(\cpu.uart.cycle_counter[8] ),
    .B(net278),
    .C(_06556_));
 sg13g2_nor3_1 _13291_ (.A(net3627),
    .B(net279),
    .C(_06559_),
    .Y(_00863_));
 sg13g2_nor2_1 _13292_ (.A(net368),
    .B(_06559_),
    .Y(_06560_));
 sg13g2_and2_1 _13293_ (.A(net368),
    .B(_06559_),
    .X(_06561_));
 sg13g2_nor3_1 _13294_ (.A(net3627),
    .B(net369),
    .C(_06561_),
    .Y(_00864_));
 sg13g2_nor2_1 _13295_ (.A(net378),
    .B(_06561_),
    .Y(_06562_));
 sg13g2_and2_1 _13296_ (.A(net378),
    .B(_06561_),
    .X(_06563_));
 sg13g2_nor3_1 _13297_ (.A(net3627),
    .B(_06562_),
    .C(_06563_),
    .Y(_00865_));
 sg13g2_a21oi_1 _13298_ (.A1(net706),
    .A2(_06563_),
    .Y(_06564_),
    .B1(net3627));
 sg13g2_o21ai_1 _13299_ (.B1(_06564_),
    .Y(_06565_),
    .A1(net706),
    .A2(_06563_));
 sg13g2_inv_1 _13300_ (.Y(_00866_),
    .A(_06565_));
 sg13g2_nand2_1 _13301_ (.Y(_06566_),
    .A(net4476),
    .B(\cpu.rx_speed[0] ));
 sg13g2_o21ai_1 _13302_ (.B1(_06566_),
    .Y(_00867_),
    .A1(net4476),
    .A2(_00900_));
 sg13g2_mux2_1 _13303_ (.A0(_00253_),
    .A1(net28),
    .S(net4476),
    .X(_00868_));
 sg13g2_mux2_1 _13304_ (.A0(net198),
    .A1(\cpu.rx_speed[2] ),
    .S(net4476),
    .X(_00869_));
 sg13g2_mux2_1 _13305_ (.A0(_00254_),
    .A1(net26),
    .S(net4477),
    .X(_00870_));
 sg13g2_mux2_1 _13306_ (.A0(net187),
    .A1(\cpu.rx_speed[4] ),
    .S(net4476),
    .X(_00871_));
 sg13g2_mux2_1 _13307_ (.A0(_00255_),
    .A1(net37),
    .S(net4476),
    .X(_00872_));
 sg13g2_mux2_1 _13308_ (.A0(_00256_),
    .A1(net32),
    .S(net4475),
    .X(_00873_));
 sg13g2_mux2_1 _13309_ (.A0(net288),
    .A1(\cpu.rx_speed[7] ),
    .S(net4476),
    .X(_00874_));
 sg13g2_nand2_1 _13310_ (.Y(_06567_),
    .A(net4475),
    .B(\cpu.rx_speed[8] ));
 sg13g2_o21ai_1 _13311_ (.B1(_06567_),
    .Y(_00875_),
    .A1(net4476),
    .A2(_00903_));
 sg13g2_mux2_1 _13312_ (.A0(net352),
    .A1(net248),
    .S(net4475),
    .X(_00876_));
 sg13g2_mux2_1 _13313_ (.A0(net376),
    .A1(\cpu.rx_speed[10] ),
    .S(net4475),
    .X(_00877_));
 sg13g2_mux2_1 _13314_ (.A0(_00257_),
    .A1(net24),
    .S(net4475),
    .X(_00878_));
 sg13g2_mux2_1 _13315_ (.A0(_00258_),
    .A1(net39),
    .S(net4475),
    .X(_00879_));
 sg13g2_a21oi_1 _13316_ (.A1(_00027_),
    .A2(_06540_),
    .Y(_06568_),
    .B1(net34));
 sg13g2_mux4_1 _13317_ (.S0(net4267),
    .A0(\cpu.uart.data_sending[0] ),
    .A1(\cpu.uart.data_sending[1] ),
    .A2(\cpu.uart.data_sending[2] ),
    .A3(\cpu.uart.data_sending[3] ),
    .S1(\cpu.uart.bit_counter[1] ),
    .X(_06569_));
 sg13g2_mux2_1 _13318_ (.A0(\cpu.uart.data_sending[4] ),
    .A1(\cpu.uart.data_sending[5] ),
    .S(\cpu.uart.bit_counter[0] ),
    .X(_06570_));
 sg13g2_nor2b_1 _13319_ (.A(\cpu.uart.data_sending[7] ),
    .B_N(net4267),
    .Y(_06571_));
 sg13g2_o21ai_1 _13320_ (.B1(\cpu.uart.bit_counter[1] ),
    .Y(_06572_),
    .A1(net4267),
    .A2(\cpu.uart.data_sending[6] ));
 sg13g2_o21ai_1 _13321_ (.B1(\cpu.uart.bit_counter[2] ),
    .Y(_06573_),
    .A1(_06571_),
    .A2(_06572_));
 sg13g2_a21oi_1 _13322_ (.A1(_00904_),
    .A2(_06570_),
    .Y(_06574_),
    .B1(_06573_));
 sg13g2_nor2_1 _13323_ (.A(_00028_),
    .B(_06574_),
    .Y(_06575_));
 sg13g2_o21ai_1 _13324_ (.B1(_06575_),
    .Y(_06576_),
    .A1(\cpu.uart.bit_counter[2] ),
    .A2(_06569_));
 sg13g2_o21ai_1 _13325_ (.B1(_00027_),
    .Y(_06577_),
    .A1(\cpu.uart.stage[1] ),
    .A2(\cpu.uart.stage[2] ));
 sg13g2_a21oi_1 _13326_ (.A1(_00007_),
    .A2(_06576_),
    .Y(_06578_),
    .B1(_06577_));
 sg13g2_a21oi_1 _13327_ (.A1(_06540_),
    .A2(_06578_),
    .Y(_00880_),
    .B1(net35));
 sg13g2_nor2_1 _13328_ (.A(_00028_),
    .B(_01283_),
    .Y(_06579_));
 sg13g2_or3_2 _13329_ (.A(_01219_),
    .B(_06577_),
    .C(_06579_),
    .X(_06580_));
 sg13g2_nor3_1 _13330_ (.A(net817),
    .B(net4267),
    .C(_06580_),
    .Y(_06581_));
 sg13g2_a21o_1 _13331_ (.A2(_06580_),
    .A1(net4267),
    .B1(_06581_),
    .X(_00881_));
 sg13g2_nor2_1 _13332_ (.A(_00905_),
    .B(_01220_),
    .Y(_06582_));
 sg13g2_and2_1 _13333_ (.A(_01282_),
    .B(_06582_),
    .X(_06583_));
 sg13g2_mux2_1 _13334_ (.A0(_06583_),
    .A1(net844),
    .S(_06580_),
    .X(_00882_));
 sg13g2_o21ai_1 _13335_ (.B1(_00007_),
    .Y(_06584_),
    .A1(_00029_),
    .A2(_01282_));
 sg13g2_a21oi_1 _13336_ (.A1(_00029_),
    .A2(_01282_),
    .Y(_06585_),
    .B1(_06584_));
 sg13g2_mux2_1 _13337_ (.A0(_06585_),
    .A1(net580),
    .S(_06580_),
    .X(_00883_));
 sg13g2_dfrbp_1 _13338_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4640),
    .D(net419),
    .Q_N(_00147_),
    .Q(\cpu.registers[4][0] ));
 sg13g2_dfrbp_1 _13339_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4683),
    .D(net225),
    .Q_N(_00151_),
    .Q(\cpu.registers[4][1] ));
 sg13g2_dfrbp_1 _13340_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4641),
    .D(net201),
    .Q_N(_00155_),
    .Q(\cpu.registers[4][2] ));
 sg13g2_dfrbp_1 _13341_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4680),
    .D(net272),
    .Q_N(_00159_),
    .Q(\cpu.registers[4][3] ));
 sg13g2_dfrbp_1 _13342_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4681),
    .D(_00267_),
    .Q_N(_00163_),
    .Q(\cpu.registers[4][4] ));
 sg13g2_dfrbp_1 _13343_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4677),
    .D(net293),
    .Q_N(_00167_),
    .Q(\cpu.registers[4][5] ));
 sg13g2_dfrbp_1 _13344_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4679),
    .D(_00269_),
    .Q_N(_00171_),
    .Q(\cpu.registers[4][6] ));
 sg13g2_dfrbp_1 _13345_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4676),
    .D(net275),
    .Q_N(_00175_),
    .Q(\cpu.registers[4][7] ));
 sg13g2_dfrbp_1 _13346_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4624),
    .D(net403),
    .Q_N(_00179_),
    .Q(\cpu.registers[4][8] ));
 sg13g2_dfrbp_1 _13347_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4639),
    .D(net223),
    .Q_N(_00183_),
    .Q(\cpu.registers[4][9] ));
 sg13g2_dfrbp_1 _13348_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4623),
    .D(net313),
    .Q_N(_00187_),
    .Q(\cpu.registers[4][10] ));
 sg13g2_dfrbp_1 _13349_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4626),
    .D(net341),
    .Q_N(_00191_),
    .Q(\cpu.registers[4][11] ));
 sg13g2_dfrbp_1 _13350_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4637),
    .D(net295),
    .Q_N(_00195_),
    .Q(\cpu.registers[4][12] ));
 sg13g2_dfrbp_1 _13351_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4622),
    .D(net397),
    .Q_N(_00199_),
    .Q(\cpu.registers[4][13] ));
 sg13g2_dfrbp_1 _13352_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4620),
    .D(net330),
    .Q_N(_00204_),
    .Q(\cpu.registers[4][14] ));
 sg13g2_dfrbp_1 _13353_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4622),
    .D(net400),
    .Q_N(_00208_),
    .Q(\cpu.registers[4][15] ));
 sg13g2_dfrbp_1 _13354_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4640),
    .D(net620),
    .Q_N(_00211_),
    .Q(\cpu.registers[3][0] ));
 sg13g2_dfrbp_1 _13355_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4680),
    .D(net433),
    .Q_N(_00212_),
    .Q(\cpu.registers[3][1] ));
 sg13g2_dfrbp_1 _13356_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4641),
    .D(net486),
    .Q_N(_00213_),
    .Q(\cpu.registers[3][2] ));
 sg13g2_dfrbp_1 _13357_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4680),
    .D(net630),
    .Q_N(_00214_),
    .Q(\cpu.registers[3][3] ));
 sg13g2_dfrbp_1 _13358_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4680),
    .D(net361),
    .Q_N(_00215_),
    .Q(\cpu.registers[3][4] ));
 sg13g2_dfrbp_1 _13359_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4677),
    .D(net501),
    .Q_N(_00216_),
    .Q(\cpu.registers[3][5] ));
 sg13g2_dfrbp_1 _13360_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4679),
    .D(net476),
    .Q_N(_00217_),
    .Q(\cpu.registers[3][6] ));
 sg13g2_dfrbp_1 _13361_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4676),
    .D(net527),
    .Q_N(_00218_),
    .Q(\cpu.registers[3][7] ));
 sg13g2_dfrbp_1 _13362_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4624),
    .D(net798),
    .Q_N(_00219_),
    .Q(\cpu.registers[3][8] ));
 sg13g2_dfrbp_1 _13363_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4637),
    .D(net687),
    .Q_N(_00220_),
    .Q(\cpu.registers[3][9] ));
 sg13g2_dfrbp_1 _13364_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4620),
    .D(net704),
    .Q_N(_00221_),
    .Q(\cpu.registers[3][10] ));
 sg13g2_dfrbp_1 _13365_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4602),
    .D(net602),
    .Q_N(_00222_),
    .Q(\cpu.registers[3][11] ));
 sg13g2_dfrbp_1 _13366_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net4637),
    .D(net647),
    .Q_N(_00223_),
    .Q(\cpu.registers[3][12] ));
 sg13g2_dfrbp_1 _13367_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4621),
    .D(net653),
    .Q_N(_00224_),
    .Q(\cpu.registers[3][13] ));
 sg13g2_dfrbp_1 _13368_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4620),
    .D(net623),
    .Q_N(_00225_),
    .Q(\cpu.registers[3][14] ));
 sg13g2_dfrbp_1 _13369_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4627),
    .D(net712),
    .Q_N(_00226_),
    .Q(\cpu.registers[3][15] ));
 sg13g2_dfrbp_1 _13370_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4640),
    .D(net519),
    .Q_N(_00049_),
    .Q(\cpu.registers[2][0] ));
 sg13g2_dfrbp_1 _13371_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net4678),
    .D(net535),
    .Q_N(_00050_),
    .Q(\cpu.registers[2][1] ));
 sg13g2_dfrbp_1 _13372_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4642),
    .D(net322),
    .Q_N(_00051_),
    .Q(\cpu.registers[2][2] ));
 sg13g2_dfrbp_1 _13373_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4688),
    .D(net753),
    .Q_N(_00052_),
    .Q(\cpu.registers[2][3] ));
 sg13g2_dfrbp_1 _13374_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4687),
    .D(net594),
    .Q_N(_00053_),
    .Q(\cpu.registers[2][4] ));
 sg13g2_dfrbp_1 _13375_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4683),
    .D(net571),
    .Q_N(_00054_),
    .Q(\cpu.registers[2][5] ));
 sg13g2_dfrbp_1 _13376_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net4682),
    .D(net627),
    .Q_N(_00055_),
    .Q(\cpu.registers[2][6] ));
 sg13g2_dfrbp_1 _13377_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net4676),
    .D(net577),
    .Q_N(_00056_),
    .Q(\cpu.registers[2][7] ));
 sg13g2_dfrbp_1 _13378_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4624),
    .D(net531),
    .Q_N(_00057_),
    .Q(\cpu.registers[2][8] ));
 sg13g2_dfrbp_1 _13379_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4638),
    .D(net463),
    .Q_N(_00058_),
    .Q(\cpu.registers[2][9] ));
 sg13g2_dfrbp_1 _13380_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4620),
    .D(net481),
    .Q_N(_00059_),
    .Q(\cpu.registers[2][10] ));
 sg13g2_dfrbp_1 _13381_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4624),
    .D(net554),
    .Q_N(_00060_),
    .Q(\cpu.registers[2][11] ));
 sg13g2_dfrbp_1 _13382_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4638),
    .D(net545),
    .Q_N(_00061_),
    .Q(\cpu.registers[2][12] ));
 sg13g2_dfrbp_1 _13383_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4625),
    .D(net515),
    .Q_N(_00062_),
    .Q(\cpu.registers[2][13] ));
 sg13g2_dfrbp_1 _13384_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4625),
    .D(net537),
    .Q_N(_00063_),
    .Q(\cpu.registers[2][14] ));
 sg13g2_dfrbp_1 _13385_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4628),
    .D(net327),
    .Q_N(_00064_),
    .Q(\cpu.registers[2][15] ));
 sg13g2_dfrbp_1 _13386_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4642),
    .D(net492),
    .Q_N(_00156_),
    .Q(\cpu.registers[1][2] ));
 sg13g2_dfrbp_1 _13387_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4681),
    .D(_00312_),
    .Q_N(_00160_),
    .Q(\cpu.registers[1][3] ));
 sg13g2_dfrbp_1 _13388_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4681),
    .D(_00313_),
    .Q_N(_00164_),
    .Q(\cpu.registers[1][4] ));
 sg13g2_dfrbp_1 _13389_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4652),
    .D(net205),
    .Q_N(_06973_),
    .Q(\cpu.jump_con ));
 sg13g2_dfrbp_1 _13390_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4698),
    .D(_00315_),
    .Q_N(_06972_),
    .Q(\cpu.rx_speed[0] ));
 sg13g2_dfrbp_1 _13391_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4691),
    .D(_00316_),
    .Q_N(_00249_),
    .Q(\cpu.rx_speed[1] ));
 sg13g2_dfrbp_1 _13392_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4691),
    .D(_00317_),
    .Q_N(_06971_),
    .Q(\cpu.rx_speed[2] ));
 sg13g2_dfrbp_1 _13393_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4698),
    .D(_00318_),
    .Q_N(_00248_),
    .Q(\cpu.rx_speed[3] ));
 sg13g2_dfrbp_1 _13394_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4691),
    .D(_00319_),
    .Q_N(_06970_),
    .Q(\cpu.rx_speed[4] ));
 sg13g2_dfrbp_1 _13395_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4692),
    .D(_00320_),
    .Q_N(_00247_),
    .Q(\cpu.rx_speed[5] ));
 sg13g2_dfrbp_1 _13396_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4692),
    .D(_00321_),
    .Q_N(_00246_),
    .Q(\cpu.rx_speed[6] ));
 sg13g2_dfrbp_1 _13397_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4692),
    .D(net682),
    .Q_N(_06969_),
    .Q(\cpu.rx_speed[7] ));
 sg13g2_dfrbp_1 _13398_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4692),
    .D(_00323_),
    .Q_N(_06968_),
    .Q(\cpu.rx_speed[8] ));
 sg13g2_dfrbp_1 _13399_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4689),
    .D(net249),
    .Q_N(_06967_),
    .Q(\cpu.rx_speed[9] ));
 sg13g2_dfrbp_1 _13400_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4689),
    .D(_00325_),
    .Q_N(_06966_),
    .Q(\cpu.rx_speed[10] ));
 sg13g2_dfrbp_1 _13401_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4692),
    .D(_00326_),
    .Q_N(_00245_),
    .Q(\cpu.rx_speed[11] ));
 sg13g2_dfrbp_1 _13402_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4692),
    .D(_00327_),
    .Q_N(_00244_),
    .Q(\cpu.rx_speed[12] ));
 sg13g2_dfrbp_1 _13403_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4671),
    .D(_00328_),
    .Q_N(_06965_),
    .Q(\cpu.keccak_alu.registers[0] ));
 sg13g2_dfrbp_1 _13404_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4663),
    .D(_00329_),
    .Q_N(_06964_),
    .Q(\cpu.keccak_alu.registers[1] ));
 sg13g2_dfrbp_1 _13405_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4664),
    .D(_00330_),
    .Q_N(_06963_),
    .Q(\cpu.keccak_alu.registers[2] ));
 sg13g2_dfrbp_1 _13406_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net4669),
    .D(_00331_),
    .Q_N(_06962_),
    .Q(\cpu.keccak_alu.registers[3] ));
 sg13g2_dfrbp_1 _13407_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4660),
    .D(_00332_),
    .Q_N(_06961_),
    .Q(\cpu.keccak_alu.registers[4] ));
 sg13g2_dfrbp_1 _13408_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net4656),
    .D(_00333_),
    .Q_N(_06960_),
    .Q(\cpu.keccak_alu.registers[5] ));
 sg13g2_dfrbp_1 _13409_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4659),
    .D(_00334_),
    .Q_N(_06959_),
    .Q(\cpu.keccak_alu.registers[6] ));
 sg13g2_dfrbp_1 _13410_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net4615),
    .D(_00335_),
    .Q_N(_06958_),
    .Q(\cpu.keccak_alu.registers[7] ));
 sg13g2_dfrbp_1 _13411_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net4606),
    .D(_00336_),
    .Q_N(_06957_),
    .Q(\cpu.keccak_alu.registers[8] ));
 sg13g2_dfrbp_1 _13412_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net4586),
    .D(_00337_),
    .Q_N(_06956_),
    .Q(\cpu.keccak_alu.registers[9] ));
 sg13g2_dfrbp_1 _13413_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net4586),
    .D(_00338_),
    .Q_N(_06955_),
    .Q(\cpu.keccak_alu.registers[10] ));
 sg13g2_dfrbp_1 _13414_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net4592),
    .D(_00339_),
    .Q_N(_06954_),
    .Q(\cpu.keccak_alu.registers[11] ));
 sg13g2_dfrbp_1 _13415_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net4607),
    .D(_00340_),
    .Q_N(_06953_),
    .Q(\cpu.keccak_alu.registers[12] ));
 sg13g2_dfrbp_1 _13416_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4596),
    .D(_00341_),
    .Q_N(_06952_),
    .Q(\cpu.keccak_alu.registers[13] ));
 sg13g2_dfrbp_1 _13417_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net4586),
    .D(_00342_),
    .Q_N(_06951_),
    .Q(\cpu.keccak_alu.registers[14] ));
 sg13g2_dfrbp_1 _13418_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4601),
    .D(_00343_),
    .Q_N(_06950_),
    .Q(\cpu.keccak_alu.registers[15] ));
 sg13g2_dfrbp_1 _13419_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4668),
    .D(_00344_),
    .Q_N(_06949_),
    .Q(\cpu.keccak_alu.registers[16] ));
 sg13g2_dfrbp_1 _13420_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4663),
    .D(_00345_),
    .Q_N(_06948_),
    .Q(\cpu.keccak_alu.registers[17] ));
 sg13g2_dfrbp_1 _13421_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4670),
    .D(_00346_),
    .Q_N(_06947_),
    .Q(\cpu.keccak_alu.registers[18] ));
 sg13g2_dfrbp_1 _13422_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4670),
    .D(_00347_),
    .Q_N(_06946_),
    .Q(\cpu.keccak_alu.registers[19] ));
 sg13g2_dfrbp_1 _13423_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net4660),
    .D(_00348_),
    .Q_N(_06945_),
    .Q(\cpu.keccak_alu.registers[20] ));
 sg13g2_dfrbp_1 _13424_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4657),
    .D(_00349_),
    .Q_N(_06944_),
    .Q(\cpu.keccak_alu.registers[21] ));
 sg13g2_dfrbp_1 _13425_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net4655),
    .D(_00350_),
    .Q_N(_06943_),
    .Q(\cpu.keccak_alu.registers[22] ));
 sg13g2_dfrbp_1 _13426_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net4616),
    .D(_00351_),
    .Q_N(_06942_),
    .Q(\cpu.keccak_alu.registers[23] ));
 sg13g2_dfrbp_1 _13427_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net4606),
    .D(_00352_),
    .Q_N(_06941_),
    .Q(\cpu.keccak_alu.registers[24] ));
 sg13g2_dfrbp_1 _13428_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net4595),
    .D(_00353_),
    .Q_N(_06940_),
    .Q(\cpu.keccak_alu.registers[25] ));
 sg13g2_dfrbp_1 _13429_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net4595),
    .D(_00354_),
    .Q_N(_06939_),
    .Q(\cpu.keccak_alu.registers[26] ));
 sg13g2_dfrbp_1 _13430_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4598),
    .D(_00355_),
    .Q_N(_06938_),
    .Q(\cpu.keccak_alu.registers[27] ));
 sg13g2_dfrbp_1 _13431_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net4609),
    .D(_00356_),
    .Q_N(_06937_),
    .Q(\cpu.keccak_alu.registers[28] ));
 sg13g2_dfrbp_1 _13432_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4595),
    .D(_00357_),
    .Q_N(_06936_),
    .Q(\cpu.keccak_alu.registers[29] ));
 sg13g2_dfrbp_1 _13433_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4596),
    .D(_00358_),
    .Q_N(_06935_),
    .Q(\cpu.keccak_alu.registers[30] ));
 sg13g2_dfrbp_1 _13434_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4599),
    .D(_00359_),
    .Q_N(_06934_),
    .Q(\cpu.keccak_alu.registers[31] ));
 sg13g2_dfrbp_1 _13435_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4667),
    .D(_00360_),
    .Q_N(_06933_),
    .Q(\cpu.keccak_alu.registers[32] ));
 sg13g2_dfrbp_1 _13436_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4666),
    .D(_00361_),
    .Q_N(_06932_),
    .Q(\cpu.keccak_alu.registers[33] ));
 sg13g2_dfrbp_1 _13437_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4665),
    .D(_00362_),
    .Q_N(_06931_),
    .Q(\cpu.keccak_alu.registers[34] ));
 sg13g2_dfrbp_1 _13438_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4668),
    .D(_00363_),
    .Q_N(_06930_),
    .Q(\cpu.keccak_alu.registers[35] ));
 sg13g2_dfrbp_1 _13439_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4660),
    .D(_00364_),
    .Q_N(_06929_),
    .Q(\cpu.keccak_alu.registers[36] ));
 sg13g2_dfrbp_1 _13440_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net4656),
    .D(_00365_),
    .Q_N(_06928_),
    .Q(\cpu.keccak_alu.registers[37] ));
 sg13g2_dfrbp_1 _13441_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4657),
    .D(_00366_),
    .Q_N(_06927_),
    .Q(\cpu.keccak_alu.registers[38] ));
 sg13g2_dfrbp_1 _13442_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net4617),
    .D(_00367_),
    .Q_N(_06926_),
    .Q(\cpu.keccak_alu.registers[39] ));
 sg13g2_dfrbp_1 _13443_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net4606),
    .D(_00368_),
    .Q_N(_06925_),
    .Q(\cpu.keccak_alu.registers[40] ));
 sg13g2_dfrbp_1 _13444_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4593),
    .D(_00369_),
    .Q_N(_06924_),
    .Q(\cpu.keccak_alu.registers[41] ));
 sg13g2_dfrbp_1 _13445_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4598),
    .D(_00370_),
    .Q_N(_06923_),
    .Q(\cpu.keccak_alu.registers[42] ));
 sg13g2_dfrbp_1 _13446_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4593),
    .D(_00371_),
    .Q_N(_06922_),
    .Q(\cpu.keccak_alu.registers[43] ));
 sg13g2_dfrbp_1 _13447_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net4618),
    .D(_00372_),
    .Q_N(_06921_),
    .Q(\cpu.keccak_alu.registers[44] ));
 sg13g2_dfrbp_1 _13448_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4601),
    .D(_00373_),
    .Q_N(_06920_),
    .Q(\cpu.keccak_alu.registers[45] ));
 sg13g2_dfrbp_1 _13449_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4593),
    .D(_00374_),
    .Q_N(_06919_),
    .Q(\cpu.keccak_alu.registers[46] ));
 sg13g2_dfrbp_1 _13450_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4602),
    .D(_00375_),
    .Q_N(_06918_),
    .Q(\cpu.keccak_alu.registers[47] ));
 sg13g2_dfrbp_1 _13451_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4667),
    .D(_00376_),
    .Q_N(_06917_),
    .Q(\cpu.keccak_alu.registers[48] ));
 sg13g2_dfrbp_1 _13452_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4666),
    .D(_00377_),
    .Q_N(_06916_),
    .Q(\cpu.keccak_alu.registers[49] ));
 sg13g2_dfrbp_1 _13453_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4666),
    .D(_00378_),
    .Q_N(_06915_),
    .Q(\cpu.keccak_alu.registers[50] ));
 sg13g2_dfrbp_1 _13454_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4668),
    .D(_00379_),
    .Q_N(_06914_),
    .Q(\cpu.keccak_alu.registers[51] ));
 sg13g2_dfrbp_1 _13455_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4661),
    .D(_00380_),
    .Q_N(_06913_),
    .Q(\cpu.keccak_alu.registers[52] ));
 sg13g2_dfrbp_1 _13456_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net4617),
    .D(_00381_),
    .Q_N(_06912_),
    .Q(\cpu.keccak_alu.registers[53] ));
 sg13g2_dfrbp_1 _13457_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net4655),
    .D(_00382_),
    .Q_N(_06911_),
    .Q(\cpu.keccak_alu.registers[54] ));
 sg13g2_dfrbp_1 _13458_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net4615),
    .D(_00383_),
    .Q_N(_06910_),
    .Q(\cpu.keccak_alu.registers[55] ));
 sg13g2_dfrbp_1 _13459_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net4604),
    .D(_00384_),
    .Q_N(_06909_),
    .Q(\cpu.keccak_alu.registers[56] ));
 sg13g2_dfrbp_1 _13460_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net4587),
    .D(_00385_),
    .Q_N(_06908_),
    .Q(\cpu.keccak_alu.registers[57] ));
 sg13g2_dfrbp_1 _13461_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net4587),
    .D(_00386_),
    .Q_N(_06907_),
    .Q(\cpu.keccak_alu.registers[58] ));
 sg13g2_dfrbp_1 _13462_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net4604),
    .D(_00387_),
    .Q_N(_06906_),
    .Q(\cpu.keccak_alu.registers[59] ));
 sg13g2_dfrbp_1 _13463_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net4607),
    .D(_00388_),
    .Q_N(_06905_),
    .Q(\cpu.keccak_alu.registers[60] ));
 sg13g2_dfrbp_1 _13464_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4603),
    .D(_00389_),
    .Q_N(_06904_),
    .Q(\cpu.keccak_alu.registers[61] ));
 sg13g2_dfrbp_1 _13465_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net4587),
    .D(_00390_),
    .Q_N(_06903_),
    .Q(\cpu.keccak_alu.registers[62] ));
 sg13g2_dfrbp_1 _13466_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4601),
    .D(_00391_),
    .Q_N(_06902_),
    .Q(\cpu.keccak_alu.registers[63] ));
 sg13g2_dfrbp_1 _13467_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4672),
    .D(_00392_),
    .Q_N(_06901_),
    .Q(\cpu.keccak_alu.registers[64] ));
 sg13g2_dfrbp_1 _13468_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net4663),
    .D(_00393_),
    .Q_N(_00066_),
    .Q(\cpu.keccak_alu.registers[65] ));
 sg13g2_dfrbp_1 _13469_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net4664),
    .D(_00394_),
    .Q_N(_00067_),
    .Q(\cpu.keccak_alu.registers[66] ));
 sg13g2_dfrbp_1 _13470_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net4669),
    .D(_00395_),
    .Q_N(_00068_),
    .Q(\cpu.keccak_alu.registers[67] ));
 sg13g2_dfrbp_1 _13471_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4665),
    .D(_00396_),
    .Q_N(_00070_),
    .Q(\cpu.keccak_alu.registers[68] ));
 sg13g2_dfrbp_1 _13472_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net4658),
    .D(_00397_),
    .Q_N(_00071_),
    .Q(\cpu.keccak_alu.registers[69] ));
 sg13g2_dfrbp_1 _13473_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net4658),
    .D(_00398_),
    .Q_N(_00072_),
    .Q(\cpu.keccak_alu.registers[70] ));
 sg13g2_dfrbp_1 _13474_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net4609),
    .D(_00399_),
    .Q_N(_00073_),
    .Q(\cpu.keccak_alu.registers[71] ));
 sg13g2_dfrbp_1 _13475_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net4605),
    .D(_00400_),
    .Q_N(_00074_),
    .Q(\cpu.keccak_alu.registers[72] ));
 sg13g2_dfrbp_1 _13476_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net4587),
    .D(_00401_),
    .Q_N(_00075_),
    .Q(\cpu.keccak_alu.registers[73] ));
 sg13g2_dfrbp_1 _13477_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net4586),
    .D(_00402_),
    .Q_N(_00076_),
    .Q(\cpu.keccak_alu.registers[74] ));
 sg13g2_dfrbp_1 _13478_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net4604),
    .D(_00403_),
    .Q_N(_00077_),
    .Q(\cpu.keccak_alu.registers[75] ));
 sg13g2_dfrbp_1 _13479_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net4608),
    .D(_00404_),
    .Q_N(_00078_),
    .Q(\cpu.keccak_alu.registers[76] ));
 sg13g2_dfrbp_1 _13480_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net4596),
    .D(_00405_),
    .Q_N(_00079_),
    .Q(\cpu.keccak_alu.registers[77] ));
 sg13g2_dfrbp_1 _13481_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net4586),
    .D(net263),
    .Q_N(_00080_),
    .Q(\cpu.keccak_alu.registers[78] ));
 sg13g2_dfrbp_1 _13482_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net4611),
    .D(_00407_),
    .Q_N(_00081_),
    .Q(\cpu.keccak_alu.registers[79] ));
 sg13g2_dfrbp_1 _13483_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net4669),
    .D(_00408_),
    .Q_N(_00082_),
    .Q(\cpu.keccak_alu.registers[80] ));
 sg13g2_dfrbp_1 _13484_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net4663),
    .D(_00409_),
    .Q_N(_00083_),
    .Q(\cpu.keccak_alu.registers[81] ));
 sg13g2_dfrbp_1 _13485_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4664),
    .D(_00410_),
    .Q_N(_00084_),
    .Q(\cpu.keccak_alu.registers[82] ));
 sg13g2_dfrbp_1 _13486_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net4669),
    .D(_00411_),
    .Q_N(_00085_),
    .Q(\cpu.keccak_alu.registers[83] ));
 sg13g2_dfrbp_1 _13487_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net4661),
    .D(_00412_),
    .Q_N(_00086_),
    .Q(\cpu.keccak_alu.registers[84] ));
 sg13g2_dfrbp_1 _13488_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net4658),
    .D(_00413_),
    .Q_N(_00087_),
    .Q(\cpu.keccak_alu.registers[85] ));
 sg13g2_dfrbp_1 _13489_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net4658),
    .D(_00414_),
    .Q_N(_00088_),
    .Q(\cpu.keccak_alu.registers[86] ));
 sg13g2_dfrbp_1 _13490_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net4618),
    .D(_00415_),
    .Q_N(_00089_),
    .Q(\cpu.keccak_alu.registers[87] ));
 sg13g2_dfrbp_1 _13491_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net4605),
    .D(_00416_),
    .Q_N(_00090_),
    .Q(\cpu.keccak_alu.registers[88] ));
 sg13g2_dfrbp_1 _13492_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net4587),
    .D(_00417_),
    .Q_N(_00091_),
    .Q(\cpu.keccak_alu.registers[89] ));
 sg13g2_dfrbp_1 _13493_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4589),
    .D(_00418_),
    .Q_N(_00092_),
    .Q(\cpu.keccak_alu.registers[90] ));
 sg13g2_dfrbp_1 _13494_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net4591),
    .D(_00419_),
    .Q_N(_00093_),
    .Q(\cpu.keccak_alu.registers[91] ));
 sg13g2_dfrbp_1 _13495_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net4608),
    .D(_00420_),
    .Q_N(_00094_),
    .Q(\cpu.keccak_alu.registers[92] ));
 sg13g2_dfrbp_1 _13496_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4596),
    .D(_00421_),
    .Q_N(_00095_),
    .Q(\cpu.keccak_alu.registers[93] ));
 sg13g2_dfrbp_1 _13497_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4589),
    .D(_00422_),
    .Q_N(_00096_),
    .Q(\cpu.keccak_alu.registers[94] ));
 sg13g2_dfrbp_1 _13498_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net4611),
    .D(_00423_),
    .Q_N(_00097_),
    .Q(\cpu.keccak_alu.registers[95] ));
 sg13g2_dfrbp_1 _13499_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4665),
    .D(_00424_),
    .Q_N(_00098_),
    .Q(\cpu.keccak_alu.registers[96] ));
 sg13g2_dfrbp_1 _13500_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net4675),
    .D(_00425_),
    .Q_N(_00099_),
    .Q(\cpu.keccak_alu.registers[97] ));
 sg13g2_dfrbp_1 _13501_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4665),
    .D(_00426_),
    .Q_N(_00100_),
    .Q(\cpu.keccak_alu.registers[98] ));
 sg13g2_dfrbp_1 _13502_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4665),
    .D(_00427_),
    .Q_N(_00101_),
    .Q(\cpu.keccak_alu.registers[99] ));
 sg13g2_dfrbp_1 _13503_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4659),
    .D(_00428_),
    .Q_N(_00102_),
    .Q(\cpu.keccak_alu.registers[100] ));
 sg13g2_dfrbp_1 _13504_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net4654),
    .D(_00429_),
    .Q_N(_00103_),
    .Q(\cpu.keccak_alu.registers[101] ));
 sg13g2_dfrbp_1 _13505_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net4658),
    .D(_00430_),
    .Q_N(_00104_),
    .Q(\cpu.keccak_alu.registers[102] ));
 sg13g2_dfrbp_1 _13506_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net4654),
    .D(_00431_),
    .Q_N(_00105_),
    .Q(\cpu.keccak_alu.registers[103] ));
 sg13g2_dfrbp_1 _13507_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net4611),
    .D(_00432_),
    .Q_N(_00106_),
    .Q(\cpu.keccak_alu.registers[104] ));
 sg13g2_dfrbp_1 _13508_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net4593),
    .D(net489),
    .Q_N(_00107_),
    .Q(\cpu.keccak_alu.registers[105] ));
 sg13g2_dfrbp_1 _13509_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net4594),
    .D(net550),
    .Q_N(_00108_),
    .Q(\cpu.keccak_alu.registers[106] ));
 sg13g2_dfrbp_1 _13510_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net4604),
    .D(_00435_),
    .Q_N(_00109_),
    .Q(\cpu.keccak_alu.registers[107] ));
 sg13g2_dfrbp_1 _13511_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net4608),
    .D(_00436_),
    .Q_N(_00110_),
    .Q(\cpu.keccak_alu.registers[108] ));
 sg13g2_dfrbp_1 _13512_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net4598),
    .D(_00437_),
    .Q_N(_00111_),
    .Q(\cpu.keccak_alu.registers[109] ));
 sg13g2_dfrbp_1 _13513_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net4593),
    .D(_00438_),
    .Q_N(_00112_),
    .Q(\cpu.keccak_alu.registers[110] ));
 sg13g2_dfrbp_1 _13514_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4599),
    .D(_00439_),
    .Q_N(_00113_),
    .Q(\cpu.keccak_alu.registers[111] ));
 sg13g2_dfrbp_1 _13515_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4659),
    .D(_00440_),
    .Q_N(_00114_),
    .Q(\cpu.keccak_alu.registers[112] ));
 sg13g2_dfrbp_1 _13516_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4675),
    .D(_00441_),
    .Q_N(_00115_),
    .Q(\cpu.keccak_alu.registers[113] ));
 sg13g2_dfrbp_1 _13517_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4665),
    .D(_00442_),
    .Q_N(_00116_),
    .Q(\cpu.keccak_alu.registers[114] ));
 sg13g2_dfrbp_1 _13518_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4659),
    .D(_00443_),
    .Q_N(_00117_),
    .Q(\cpu.keccak_alu.registers[115] ));
 sg13g2_dfrbp_1 _13519_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4659),
    .D(_00444_),
    .Q_N(_00118_),
    .Q(\cpu.keccak_alu.registers[116] ));
 sg13g2_dfrbp_1 _13520_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net4655),
    .D(_00445_),
    .Q_N(_00119_),
    .Q(\cpu.keccak_alu.registers[117] ));
 sg13g2_dfrbp_1 _13521_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net4655),
    .D(_00446_),
    .Q_N(_00120_),
    .Q(\cpu.keccak_alu.registers[118] ));
 sg13g2_dfrbp_1 _13522_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net4609),
    .D(_00447_),
    .Q_N(_00121_),
    .Q(\cpu.keccak_alu.registers[119] ));
 sg13g2_dfrbp_1 _13523_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net4605),
    .D(_00448_),
    .Q_N(_00122_),
    .Q(\cpu.keccak_alu.registers[120] ));
 sg13g2_dfrbp_1 _13524_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net4605),
    .D(net760),
    .Q_N(_00123_),
    .Q(\cpu.keccak_alu.registers[121] ));
 sg13g2_dfrbp_1 _13525_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net4591),
    .D(net800),
    .Q_N(_00124_),
    .Q(\cpu.keccak_alu.registers[122] ));
 sg13g2_dfrbp_1 _13526_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net4604),
    .D(_00451_),
    .Q_N(_00125_),
    .Q(\cpu.keccak_alu.registers[123] ));
 sg13g2_dfrbp_1 _13527_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net4608),
    .D(_00452_),
    .Q_N(_00126_),
    .Q(\cpu.keccak_alu.registers[124] ));
 sg13g2_dfrbp_1 _13528_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4599),
    .D(net568),
    .Q_N(_00127_),
    .Q(\cpu.keccak_alu.registers[125] ));
 sg13g2_dfrbp_1 _13529_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net4591),
    .D(_00454_),
    .Q_N(_00128_),
    .Q(\cpu.keccak_alu.registers[126] ));
 sg13g2_dfrbp_1 _13530_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4599),
    .D(_00455_),
    .Q_N(_00129_),
    .Q(\cpu.keccak_alu.registers[127] ));
 sg13g2_dfrbp_1 _13531_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4672),
    .D(_00456_),
    .Q_N(_06900_),
    .Q(\cpu.keccak_alu.registers[128] ));
 sg13g2_dfrbp_1 _13532_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net4670),
    .D(_00457_),
    .Q_N(_06899_),
    .Q(\cpu.keccak_alu.registers[129] ));
 sg13g2_dfrbp_1 _13533_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net4663),
    .D(_00458_),
    .Q_N(_00069_),
    .Q(\cpu.keccak_alu.registers[130] ));
 sg13g2_dfrbp_1 _13534_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4671),
    .D(_00459_),
    .Q_N(_06898_),
    .Q(\cpu.keccak_alu.registers[131] ));
 sg13g2_dfrbp_1 _13535_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4667),
    .D(_00460_),
    .Q_N(_06897_),
    .Q(\cpu.keccak_alu.registers[132] ));
 sg13g2_dfrbp_1 _13536_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net4654),
    .D(_00461_),
    .Q_N(_06896_),
    .Q(\cpu.keccak_alu.registers[133] ));
 sg13g2_dfrbp_1 _13537_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net4665),
    .D(_00462_),
    .Q_N(_06895_),
    .Q(\cpu.keccak_alu.registers[134] ));
 sg13g2_dfrbp_1 _13538_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net4615),
    .D(_00463_),
    .Q_N(_06894_),
    .Q(\cpu.keccak_alu.registers[135] ));
 sg13g2_dfrbp_1 _13539_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net4606),
    .D(_00464_),
    .Q_N(_06893_),
    .Q(\cpu.keccak_alu.registers[136] ));
 sg13g2_dfrbp_1 _13540_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net4591),
    .D(net928),
    .Q_N(_06892_),
    .Q(\cpu.keccak_alu.registers[137] ));
 sg13g2_dfrbp_1 _13541_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net4606),
    .D(_00466_),
    .Q_N(_00065_),
    .Q(\cpu.keccak_alu.registers[138] ));
 sg13g2_dfrbp_1 _13542_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net4591),
    .D(_00467_),
    .Q_N(_06891_),
    .Q(\cpu.keccak_alu.registers[139] ));
 sg13g2_dfrbp_1 _13543_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net4605),
    .D(net830),
    .Q_N(_06890_),
    .Q(\cpu.keccak_alu.registers[140] ));
 sg13g2_dfrbp_1 _13544_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4600),
    .D(net903),
    .Q_N(_06889_),
    .Q(\cpu.keccak_alu.registers[141] ));
 sg13g2_dfrbp_1 _13545_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net4591),
    .D(_00470_),
    .Q_N(_06888_),
    .Q(\cpu.keccak_alu.registers[142] ));
 sg13g2_dfrbp_1 _13546_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4614),
    .D(_00471_),
    .Q_N(_06887_),
    .Q(\cpu.keccak_alu.registers[143] ));
 sg13g2_dfrbp_1 _13547_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4654),
    .D(_00472_),
    .Q_N(_06886_),
    .Q(\cpu.keccak_alu.registers[144] ));
 sg13g2_dfrbp_1 _13548_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net4612),
    .D(net925),
    .Q_N(_06885_),
    .Q(\cpu.keccak_alu.registers[145] ));
 sg13g2_dfrbp_1 _13549_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net4655),
    .D(_00474_),
    .Q_N(_06884_),
    .Q(\cpu.keccak_alu.registers[146] ));
 sg13g2_dfrbp_1 _13550_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net4613),
    .D(_00475_),
    .Q_N(_06883_),
    .Q(\cpu.keccak_alu.registers[147] ));
 sg13g2_dfrbp_1 _13551_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4617),
    .D(_00476_),
    .Q_N(_06882_),
    .Q(\cpu.keccak_alu.registers[148] ));
 sg13g2_dfrbp_1 _13552_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net4654),
    .D(_00477_),
    .Q_N(_06881_),
    .Q(\cpu.keccak_alu.registers[149] ));
 sg13g2_dfrbp_1 _13553_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net4655),
    .D(_00478_),
    .Q_N(_06880_),
    .Q(\cpu.keccak_alu.registers[150] ));
 sg13g2_dfrbp_1 _13554_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4612),
    .D(_00479_),
    .Q_N(_06879_),
    .Q(\cpu.keccak_alu.registers[151] ));
 sg13g2_dfrbp_1 _13555_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4611),
    .D(_00480_),
    .Q_N(_06878_),
    .Q(\cpu.keccak_alu.registers[152] ));
 sg13g2_dfrbp_1 _13556_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net4595),
    .D(_00481_),
    .Q_N(_06877_),
    .Q(\cpu.keccak_alu.registers[153] ));
 sg13g2_dfrbp_1 _13557_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4595),
    .D(_00482_),
    .Q_N(_06876_),
    .Q(\cpu.keccak_alu.registers[154] ));
 sg13g2_dfrbp_1 _13558_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net4598),
    .D(_00483_),
    .Q_N(_06875_),
    .Q(\cpu.keccak_alu.registers[155] ));
 sg13g2_dfrbp_1 _13559_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net4612),
    .D(_00484_),
    .Q_N(_06874_),
    .Q(\cpu.keccak_alu.registers[156] ));
 sg13g2_dfrbp_1 _13560_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net4595),
    .D(_00485_),
    .Q_N(_06873_),
    .Q(\cpu.keccak_alu.registers[157] ));
 sg13g2_dfrbp_1 _13561_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net4595),
    .D(_00486_),
    .Q_N(_06872_),
    .Q(\cpu.keccak_alu.registers[158] ));
 sg13g2_dfrbp_1 _13562_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4611),
    .D(_00487_),
    .Q_N(_06871_),
    .Q(\cpu.keccak_alu.registers[159] ));
 sg13g2_dfrbp_1 _13563_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4616),
    .D(net643),
    .Q_N(_06870_),
    .Q(\cpu.keccak_alu.registers[160] ));
 sg13g2_dfrbp_1 _13564_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net4612),
    .D(net938),
    .Q_N(_06869_),
    .Q(\cpu.keccak_alu.registers[161] ));
 sg13g2_dfrbp_1 _13565_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net4612),
    .D(_00490_),
    .Q_N(_06868_),
    .Q(\cpu.keccak_alu.registers[162] ));
 sg13g2_dfrbp_1 _13566_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net4613),
    .D(_00491_),
    .Q_N(_06867_),
    .Q(\cpu.keccak_alu.registers[163] ));
 sg13g2_dfrbp_1 _13567_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net4616),
    .D(_00492_),
    .Q_N(_06866_),
    .Q(\cpu.keccak_alu.registers[164] ));
 sg13g2_dfrbp_1 _13568_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4613),
    .D(net923),
    .Q_N(_06865_),
    .Q(\cpu.keccak_alu.registers[165] ));
 sg13g2_dfrbp_1 _13569_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net4616),
    .D(_00494_),
    .Q_N(_06864_),
    .Q(\cpu.keccak_alu.registers[166] ));
 sg13g2_dfrbp_1 _13570_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net4615),
    .D(_00495_),
    .Q_N(_06863_),
    .Q(\cpu.keccak_alu.registers[167] ));
 sg13g2_dfrbp_1 _13571_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4611),
    .D(_00496_),
    .Q_N(_06862_),
    .Q(\cpu.keccak_alu.registers[168] ));
 sg13g2_dfrbp_1 _13572_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4598),
    .D(_00497_),
    .Q_N(_06861_),
    .Q(\cpu.keccak_alu.registers[169] ));
 sg13g2_dfrbp_1 _13573_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4598),
    .D(_00498_),
    .Q_N(_06860_),
    .Q(\cpu.keccak_alu.registers[170] ));
 sg13g2_dfrbp_1 _13574_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4599),
    .D(_00499_),
    .Q_N(_06859_),
    .Q(\cpu.keccak_alu.registers[171] ));
 sg13g2_dfrbp_1 _13575_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net4615),
    .D(_00500_),
    .Q_N(_06858_),
    .Q(\cpu.keccak_alu.registers[172] ));
 sg13g2_dfrbp_1 _13576_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4598),
    .D(_00501_),
    .Q_N(_06857_),
    .Q(\cpu.keccak_alu.registers[173] ));
 sg13g2_dfrbp_1 _13577_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4599),
    .D(_00502_),
    .Q_N(_06856_),
    .Q(\cpu.keccak_alu.registers[174] ));
 sg13g2_dfrbp_1 _13578_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net4613),
    .D(_00503_),
    .Q_N(_06855_),
    .Q(\cpu.keccak_alu.registers[175] ));
 sg13g2_dfrbp_1 _13579_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4667),
    .D(_00504_),
    .Q_N(_06854_),
    .Q(\cpu.keccak_alu.registers[176] ));
 sg13g2_dfrbp_1 _13580_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4666),
    .D(_00505_),
    .Q_N(_06853_),
    .Q(\cpu.keccak_alu.registers[177] ));
 sg13g2_dfrbp_1 _13581_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4665),
    .D(_00506_),
    .Q_N(_06852_),
    .Q(\cpu.keccak_alu.registers[178] ));
 sg13g2_dfrbp_1 _13582_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4668),
    .D(_00507_),
    .Q_N(_06851_),
    .Q(\cpu.keccak_alu.registers[179] ));
 sg13g2_dfrbp_1 _13583_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net4616),
    .D(net852),
    .Q_N(_06850_),
    .Q(\cpu.keccak_alu.registers[180] ));
 sg13g2_dfrbp_1 _13584_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4617),
    .D(net124),
    .Q_N(_06849_),
    .Q(\cpu.keccak_alu.registers[181] ));
 sg13g2_dfrbp_1 _13585_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net4654),
    .D(net847),
    .Q_N(_06848_),
    .Q(\cpu.keccak_alu.registers[182] ));
 sg13g2_dfrbp_1 _13586_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net4654),
    .D(_00511_),
    .Q_N(_06847_),
    .Q(\cpu.keccak_alu.registers[183] ));
 sg13g2_dfrbp_1 _13587_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net4605),
    .D(_00512_),
    .Q_N(_06846_),
    .Q(\cpu.keccak_alu.registers[184] ));
 sg13g2_dfrbp_1 _13588_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net4592),
    .D(_00513_),
    .Q_N(_06845_),
    .Q(\cpu.keccak_alu.registers[185] ));
 sg13g2_dfrbp_1 _13589_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net4592),
    .D(_00514_),
    .Q_N(_06844_),
    .Q(\cpu.keccak_alu.registers[186] ));
 sg13g2_dfrbp_1 _13590_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net4604),
    .D(_00515_),
    .Q_N(_06843_),
    .Q(\cpu.keccak_alu.registers[187] ));
 sg13g2_dfrbp_1 _13591_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net4607),
    .D(_00516_),
    .Q_N(_06842_),
    .Q(\cpu.keccak_alu.registers[188] ));
 sg13g2_dfrbp_1 _13592_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4600),
    .D(_00517_),
    .Q_N(_06841_),
    .Q(\cpu.keccak_alu.registers[189] ));
 sg13g2_dfrbp_1 _13593_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net4592),
    .D(_00518_),
    .Q_N(_06840_),
    .Q(\cpu.keccak_alu.registers[190] ));
 sg13g2_dfrbp_1 _13594_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4601),
    .D(net886),
    .Q_N(_06839_),
    .Q(\cpu.keccak_alu.registers[191] ));
 sg13g2_dfrbp_1 _13595_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4671),
    .D(net413),
    .Q_N(_06838_),
    .Q(\cpu.keccak_alu.registers[192] ));
 sg13g2_dfrbp_1 _13596_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net4663),
    .D(_00521_),
    .Q_N(_06837_),
    .Q(\cpu.keccak_alu.registers[193] ));
 sg13g2_dfrbp_1 _13597_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4664),
    .D(_00522_),
    .Q_N(_06836_),
    .Q(\cpu.keccak_alu.registers[194] ));
 sg13g2_dfrbp_1 _13598_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4671),
    .D(_00523_),
    .Q_N(_06835_),
    .Q(\cpu.keccak_alu.registers[195] ));
 sg13g2_dfrbp_1 _13599_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4660),
    .D(_00524_),
    .Q_N(_06834_),
    .Q(\cpu.keccak_alu.registers[196] ));
 sg13g2_dfrbp_1 _13600_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net4654),
    .D(_00525_),
    .Q_N(_06833_),
    .Q(\cpu.keccak_alu.registers[197] ));
 sg13g2_dfrbp_1 _13601_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4658),
    .D(_00526_),
    .Q_N(_06832_),
    .Q(\cpu.keccak_alu.registers[198] ));
 sg13g2_dfrbp_1 _13602_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net4615),
    .D(_00527_),
    .Q_N(_06831_),
    .Q(\cpu.keccak_alu.registers[199] ));
 sg13g2_dfrbp_1 _13603_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net4604),
    .D(_00528_),
    .Q_N(_06830_),
    .Q(\cpu.keccak_alu.registers[200] ));
 sg13g2_dfrbp_1 _13604_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net4586),
    .D(_00529_),
    .Q_N(_06829_),
    .Q(\cpu.keccak_alu.registers[201] ));
 sg13g2_dfrbp_1 _13605_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4588),
    .D(_00530_),
    .Q_N(_06828_),
    .Q(\cpu.keccak_alu.registers[202] ));
 sg13g2_dfrbp_1 _13606_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net4591),
    .D(_00531_),
    .Q_N(_06827_),
    .Q(\cpu.keccak_alu.registers[203] ));
 sg13g2_dfrbp_1 _13607_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net4607),
    .D(_00532_),
    .Q_N(_06826_),
    .Q(\cpu.keccak_alu.registers[204] ));
 sg13g2_dfrbp_1 _13608_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4597),
    .D(_00533_),
    .Q_N(_06825_),
    .Q(\cpu.keccak_alu.registers[205] ));
 sg13g2_dfrbp_1 _13609_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net4586),
    .D(_00534_),
    .Q_N(_06824_),
    .Q(\cpu.keccak_alu.registers[206] ));
 sg13g2_dfrbp_1 _13610_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net4613),
    .D(_00535_),
    .Q_N(_06823_),
    .Q(\cpu.keccak_alu.registers[207] ));
 sg13g2_dfrbp_1 _13611_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4671),
    .D(net388),
    .Q_N(_06822_),
    .Q(\cpu.keccak_alu.registers[208] ));
 sg13g2_dfrbp_1 _13612_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4663),
    .D(_00537_),
    .Q_N(_06821_),
    .Q(\cpu.keccak_alu.registers[209] ));
 sg13g2_dfrbp_1 _13613_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4670),
    .D(_00538_),
    .Q_N(_06820_),
    .Q(\cpu.keccak_alu.registers[210] ));
 sg13g2_dfrbp_1 _13614_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4671),
    .D(_00539_),
    .Q_N(_06819_),
    .Q(\cpu.keccak_alu.registers[211] ));
 sg13g2_dfrbp_1 _13615_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4660),
    .D(_00540_),
    .Q_N(_06818_),
    .Q(\cpu.keccak_alu.registers[212] ));
 sg13g2_dfrbp_1 _13616_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4612),
    .D(net779),
    .Q_N(_06817_),
    .Q(\cpu.keccak_alu.registers[213] ));
 sg13g2_dfrbp_1 _13617_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4658),
    .D(_00542_),
    .Q_N(_06816_),
    .Q(\cpu.keccak_alu.registers[214] ));
 sg13g2_dfrbp_1 _13618_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net4616),
    .D(_00543_),
    .Q_N(_06815_),
    .Q(\cpu.keccak_alu.registers[215] ));
 sg13g2_dfrbp_1 _13619_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4611),
    .D(_00544_),
    .Q_N(_06814_),
    .Q(\cpu.keccak_alu.registers[216] ));
 sg13g2_dfrbp_1 _13620_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4588),
    .D(_00545_),
    .Q_N(_06813_),
    .Q(\cpu.keccak_alu.registers[217] ));
 sg13g2_dfrbp_1 _13621_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4588),
    .D(_00546_),
    .Q_N(_06812_),
    .Q(\cpu.keccak_alu.registers[218] ));
 sg13g2_dfrbp_1 _13622_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net4592),
    .D(_00547_),
    .Q_N(_06811_),
    .Q(\cpu.keccak_alu.registers[219] ));
 sg13g2_dfrbp_1 _13623_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net4606),
    .D(net474),
    .Q_N(_06810_),
    .Q(\cpu.keccak_alu.registers[220] ));
 sg13g2_dfrbp_1 _13624_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4599),
    .D(_00549_),
    .Q_N(_06809_),
    .Q(\cpu.keccak_alu.registers[221] ));
 sg13g2_dfrbp_1 _13625_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4588),
    .D(_00550_),
    .Q_N(_06808_),
    .Q(\cpu.keccak_alu.registers[222] ));
 sg13g2_dfrbp_1 _13626_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4602),
    .D(_00551_),
    .Q_N(_06807_),
    .Q(\cpu.keccak_alu.registers[223] ));
 sg13g2_dfrbp_1 _13627_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4689),
    .D(_00552_),
    .Q_N(_06806_),
    .Q(\cpu.keccak_alu.registers[224] ));
 sg13g2_dfrbp_1 _13628_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4669),
    .D(_00553_),
    .Q_N(_06805_),
    .Q(\cpu.keccak_alu.registers[225] ));
 sg13g2_dfrbp_1 _13629_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net4666),
    .D(_00554_),
    .Q_N(_06804_),
    .Q(\cpu.keccak_alu.registers[226] ));
 sg13g2_dfrbp_1 _13630_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4667),
    .D(_00555_),
    .Q_N(_06803_),
    .Q(\cpu.keccak_alu.registers[227] ));
 sg13g2_dfrbp_1 _13631_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4679),
    .D(_00556_),
    .Q_N(_06802_),
    .Q(\cpu.keccak_alu.registers[228] ));
 sg13g2_dfrbp_1 _13632_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net4618),
    .D(_00557_),
    .Q_N(_06801_),
    .Q(\cpu.keccak_alu.registers[229] ));
 sg13g2_dfrbp_1 _13633_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4657),
    .D(_00558_),
    .Q_N(_06800_),
    .Q(\cpu.keccak_alu.registers[230] ));
 sg13g2_dfrbp_1 _13634_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net4615),
    .D(_00559_),
    .Q_N(_06799_),
    .Q(\cpu.keccak_alu.registers[231] ));
 sg13g2_dfrbp_1 _13635_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net4611),
    .D(_00560_),
    .Q_N(_06798_),
    .Q(\cpu.keccak_alu.registers[232] ));
 sg13g2_dfrbp_1 _13636_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net4592),
    .D(_00561_),
    .Q_N(_06797_),
    .Q(\cpu.keccak_alu.registers[233] ));
 sg13g2_dfrbp_1 _13637_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net4589),
    .D(_00562_),
    .Q_N(_06796_),
    .Q(\cpu.keccak_alu.registers[234] ));
 sg13g2_dfrbp_1 _13638_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net4594),
    .D(_00563_),
    .Q_N(_06795_),
    .Q(\cpu.keccak_alu.registers[235] ));
 sg13g2_dfrbp_1 _13639_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net4607),
    .D(_00564_),
    .Q_N(_06794_),
    .Q(\cpu.keccak_alu.registers[236] ));
 sg13g2_dfrbp_1 _13640_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net4598),
    .D(_00565_),
    .Q_N(_06793_),
    .Q(\cpu.keccak_alu.registers[237] ));
 sg13g2_dfrbp_1 _13641_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net4593),
    .D(net498),
    .Q_N(_06792_),
    .Q(\cpu.keccak_alu.registers[238] ));
 sg13g2_dfrbp_1 _13642_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4601),
    .D(_00567_),
    .Q_N(_06791_),
    .Q(\cpu.keccak_alu.registers[239] ));
 sg13g2_dfrbp_1 _13643_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4689),
    .D(_00568_),
    .Q_N(_06790_),
    .Q(\cpu.keccak_alu.registers[240] ));
 sg13g2_dfrbp_1 _13644_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4690),
    .D(net598),
    .Q_N(_06789_),
    .Q(\cpu.keccak_alu.registers[241] ));
 sg13g2_dfrbp_1 _13645_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4667),
    .D(_00570_),
    .Q_N(_06788_),
    .Q(\cpu.keccak_alu.registers[242] ));
 sg13g2_dfrbp_1 _13646_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4667),
    .D(_00571_),
    .Q_N(_06787_),
    .Q(\cpu.keccak_alu.registers[243] ));
 sg13g2_dfrbp_1 _13647_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4682),
    .D(_00572_),
    .Q_N(_06786_),
    .Q(\cpu.keccak_alu.registers[244] ));
 sg13g2_dfrbp_1 _13648_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4617),
    .D(_00573_),
    .Q_N(_06785_),
    .Q(\cpu.keccak_alu.registers[245] ));
 sg13g2_dfrbp_1 _13649_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4656),
    .D(_00574_),
    .Q_N(_06784_),
    .Q(\cpu.keccak_alu.registers[246] ));
 sg13g2_dfrbp_1 _13650_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net4615),
    .D(_00575_),
    .Q_N(_06783_),
    .Q(\cpu.keccak_alu.registers[247] ));
 sg13g2_dfrbp_1 _13651_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net4604),
    .D(_00576_),
    .Q_N(_06782_),
    .Q(\cpu.keccak_alu.registers[248] ));
 sg13g2_dfrbp_1 _13652_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net4587),
    .D(_00577_),
    .Q_N(_06781_),
    .Q(\cpu.keccak_alu.registers[249] ));
 sg13g2_dfrbp_1 _13653_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net4587),
    .D(_00578_),
    .Q_N(_06780_),
    .Q(\cpu.keccak_alu.registers[250] ));
 sg13g2_dfrbp_1 _13654_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net4591),
    .D(_00579_),
    .Q_N(_06779_),
    .Q(\cpu.keccak_alu.registers[251] ));
 sg13g2_dfrbp_1 _13655_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net4607),
    .D(_00580_),
    .Q_N(_06778_),
    .Q(\cpu.keccak_alu.registers[252] ));
 sg13g2_dfrbp_1 _13656_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4597),
    .D(_00581_),
    .Q_N(_06777_),
    .Q(\cpu.keccak_alu.registers[253] ));
 sg13g2_dfrbp_1 _13657_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net4592),
    .D(_00582_),
    .Q_N(_06776_),
    .Q(\cpu.keccak_alu.registers[254] ));
 sg13g2_dfrbp_1 _13658_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4601),
    .D(net436),
    .Q_N(_06974_),
    .Q(\cpu.keccak_alu.registers[255] ));
 sg13g2_dfrbp_1 _13659_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net4696),
    .D(_00009_),
    .Q_N(_00027_),
    .Q(\cpu.set_rx_speed ));
 sg13g2_dfrbp_1 _13660_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net4696),
    .D(net343),
    .Q_N(_06775_),
    .Q(\cpu.uart.send ));
 sg13g2_dfrbp_1 _13661_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4648),
    .D(net866),
    .Q_N(_06774_),
    .Q(\cpu.ALU.b[0] ));
 sg13g2_dfrbp_1 _13662_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net4684),
    .D(_00585_),
    .Q_N(_06773_),
    .Q(\cpu.ALU.b[1] ));
 sg13g2_dfrbp_1 _13663_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4686),
    .D(_00586_),
    .Q_N(_06772_),
    .Q(\cpu.ALU.b[2] ));
 sg13g2_dfrbp_1 _13664_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4688),
    .D(_00587_),
    .Q_N(_06771_),
    .Q(\cpu.ALU.b[3] ));
 sg13g2_dfrbp_1 _13665_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4687),
    .D(_00588_),
    .Q_N(_06770_),
    .Q(\cpu.ALU.b[4] ));
 sg13g2_dfrbp_1 _13666_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net4684),
    .D(_00589_),
    .Q_N(_06769_),
    .Q(\cpu.ALU.b[5] ));
 sg13g2_dfrbp_1 _13667_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4687),
    .D(_00590_),
    .Q_N(_06768_),
    .Q(\cpu.ALU.b[6] ));
 sg13g2_dfrbp_1 _13668_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4686),
    .D(_00591_),
    .Q_N(_06767_),
    .Q(\cpu.ALU.b[7] ));
 sg13g2_dfrbp_1 _13669_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net4650),
    .D(_00592_),
    .Q_N(_06766_),
    .Q(\cpu.ALU.b[8] ));
 sg13g2_dfrbp_1 _13670_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net4649),
    .D(_00593_),
    .Q_N(_06765_),
    .Q(\cpu.ALU.b[9] ));
 sg13g2_dfrbp_1 _13671_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net4650),
    .D(_00594_),
    .Q_N(_06764_),
    .Q(\cpu.ALU.b[10] ));
 sg13g2_dfrbp_1 _13672_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net4649),
    .D(_00595_),
    .Q_N(_06763_),
    .Q(\cpu.ALU.b[11] ));
 sg13g2_dfrbp_1 _13673_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net4649),
    .D(_00596_),
    .Q_N(_06762_),
    .Q(\cpu.ALU.b[12] ));
 sg13g2_dfrbp_1 _13674_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net4649),
    .D(_00597_),
    .Q_N(_06761_),
    .Q(\cpu.ALU.b[13] ));
 sg13g2_dfrbp_1 _13675_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net4649),
    .D(_00598_),
    .Q_N(_06760_),
    .Q(\cpu.ALU.b[14] ));
 sg13g2_dfrbp_1 _13676_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4648),
    .D(_00599_),
    .Q_N(_06759_),
    .Q(\cpu.ALU.b[15] ));
 sg13g2_dfrbp_1 _13677_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net4684),
    .D(net857),
    .Q_N(_06758_),
    .Q(\cpu.ALU.a[0] ));
 sg13g2_dfrbp_1 _13678_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net4685),
    .D(net850),
    .Q_N(_06757_),
    .Q(\cpu.ALU.a[1] ));
 sg13g2_dfrbp_1 _13679_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net4684),
    .D(net888),
    .Q_N(_06756_),
    .Q(\cpu.ALU.a[2] ));
 sg13g2_dfrbp_1 _13680_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4687),
    .D(net884),
    .Q_N(_06755_),
    .Q(\cpu.ALU.a[3] ));
 sg13g2_dfrbp_1 _13681_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net4688),
    .D(net843),
    .Q_N(_06754_),
    .Q(\cpu.ALU.a[4] ));
 sg13g2_dfrbp_1 _13682_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net4685),
    .D(net823),
    .Q_N(_06753_),
    .Q(\cpu.ALU.a[5] ));
 sg13g2_dfrbp_1 _13683_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net4688),
    .D(net428),
    .Q_N(_06752_),
    .Q(\cpu.ALU.a[6] ));
 sg13g2_dfrbp_1 _13684_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4684),
    .D(net839),
    .Q_N(_06751_),
    .Q(\cpu.ALU.a[7] ));
 sg13g2_dfrbp_1 _13685_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4634),
    .D(net869),
    .Q_N(_06750_),
    .Q(\cpu.ALU.a[8] ));
 sg13g2_dfrbp_1 _13686_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4646),
    .D(net834),
    .Q_N(_06749_),
    .Q(\cpu.ALU.a[9] ));
 sg13g2_dfrbp_1 _13687_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4634),
    .D(_00610_),
    .Q_N(_06748_),
    .Q(\cpu.ALU.a[10] ));
 sg13g2_dfrbp_1 _13688_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4646),
    .D(net816),
    .Q_N(_06747_),
    .Q(\cpu.ALU.a[11] ));
 sg13g2_dfrbp_1 _13689_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4643),
    .D(net745),
    .Q_N(_06746_),
    .Q(\cpu.ALU.a[12] ));
 sg13g2_dfrbp_1 _13690_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4634),
    .D(net854),
    .Q_N(_06745_),
    .Q(\cpu.ALU.a[13] ));
 sg13g2_dfrbp_1 _13691_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4634),
    .D(net664),
    .Q_N(_00201_),
    .Q(\cpu.ALU.a[14] ));
 sg13g2_dfrbp_1 _13692_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4632),
    .D(net804),
    .Q_N(_06744_),
    .Q(\cpu.ALU.a[15] ));
 sg13g2_dfrbp_1 _13693_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4649),
    .D(net791),
    .Q_N(_06743_),
    .Q(\cpu.ALU.mode[0] ));
 sg13g2_dfrbp_1 _13694_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4650),
    .D(_00617_),
    .Q_N(_06742_),
    .Q(\cpu.ALU.mode[1] ));
 sg13g2_dfrbp_1 _13695_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4649),
    .D(net69),
    .Q_N(_00148_),
    .Q(\cpu.ALU.mode[2] ));
 sg13g2_dfrbp_1 _13696_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4645),
    .D(_00619_),
    .Q_N(_06741_),
    .Q(\cpu.current_instruction[0] ));
 sg13g2_dfrbp_1 _13697_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4643),
    .D(_00620_),
    .Q_N(_06740_),
    .Q(\cpu.current_instruction[1] ));
 sg13g2_dfrbp_1 _13698_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4645),
    .D(_00621_),
    .Q_N(_06739_),
    .Q(\cpu.current_instruction[2] ));
 sg13g2_dfrbp_1 _13699_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4645),
    .D(_00622_),
    .Q_N(_06738_),
    .Q(\cpu.current_instruction[3] ));
 sg13g2_dfrbp_1 _13700_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4643),
    .D(_00623_),
    .Q_N(_00017_),
    .Q(\cpu.current_instruction[4] ));
 sg13g2_dfrbp_1 _13701_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net4647),
    .D(_00624_),
    .Q_N(_06737_),
    .Q(\cpu.current_instruction[5] ));
 sg13g2_dfrbp_1 _13702_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4648),
    .D(_00625_),
    .Q_N(_00026_),
    .Q(\cpu.current_instruction[6] ));
 sg13g2_dfrbp_1 _13703_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4638),
    .D(_00626_),
    .Q_N(_00024_),
    .Q(\cpu.current_instruction[7] ));
 sg13g2_dfrbp_1 _13704_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4643),
    .D(_00627_),
    .Q_N(_00043_),
    .Q(\cpu.current_instruction[8] ));
 sg13g2_dfrbp_1 _13705_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4640),
    .D(_00628_),
    .Q_N(_00030_),
    .Q(\cpu.current_instruction[9] ));
 sg13g2_dfrbp_1 _13706_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4645),
    .D(_00629_),
    .Q_N(_06736_),
    .Q(\cpu.current_instruction[10] ));
 sg13g2_dfrbp_1 _13707_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4645),
    .D(_00630_),
    .Q_N(_06735_),
    .Q(\cpu.current_instruction[11] ));
 sg13g2_dfrbp_1 _13708_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4639),
    .D(_00631_),
    .Q_N(_00044_),
    .Q(\cpu.current_instruction[12] ));
 sg13g2_dfrbp_1 _13709_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4646),
    .D(_00632_),
    .Q_N(_06734_),
    .Q(\cpu.current_instruction[13] ));
 sg13g2_dfrbp_1 _13710_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net4639),
    .D(_00633_),
    .Q_N(_06733_),
    .Q(\cpu.current_instruction[14] ));
 sg13g2_dfrbp_1 _13711_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net4639),
    .D(_00634_),
    .Q_N(_00025_),
    .Q(\cpu.current_instruction[15] ));
 sg13g2_dfrbp_1 _13712_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4648),
    .D(net678),
    .Q_N(_06732_),
    .Q(\cpu.current_address[0] ));
 sg13g2_dfrbp_1 _13713_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net4684),
    .D(net820),
    .Q_N(_06731_),
    .Q(\cpu.current_address[1] ));
 sg13g2_dfrbp_1 _13714_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net4642),
    .D(net467),
    .Q_N(_06730_),
    .Q(\cpu.current_address[2] ));
 sg13g2_dfrbp_1 _13715_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net4687),
    .D(net146),
    .Q_N(_06729_),
    .Q(\cpu.current_address[3] ));
 sg13g2_dfrbp_1 _13716_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net4687),
    .D(net137),
    .Q_N(_06728_),
    .Q(\cpu.current_address[4] ));
 sg13g2_dfrbp_1 _13717_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net4678),
    .D(net159),
    .Q_N(_06727_),
    .Q(\cpu.current_address[5] ));
 sg13g2_dfrbp_1 _13718_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net4687),
    .D(net143),
    .Q_N(_06726_),
    .Q(\cpu.current_address[6] ));
 sg13g2_dfrbp_1 _13719_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4678),
    .D(net542),
    .Q_N(_06725_),
    .Q(\cpu.current_address[7] ));
 sg13g2_dfrbp_1 _13720_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4626),
    .D(net236),
    .Q_N(_06724_),
    .Q(\cpu.current_address[8] ));
 sg13g2_dfrbp_1 _13721_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4638),
    .D(net131),
    .Q_N(_06723_),
    .Q(\cpu.current_address[9] ));
 sg13g2_dfrbp_1 _13722_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4625),
    .D(net356),
    .Q_N(_06722_),
    .Q(\cpu.current_address[10] ));
 sg13g2_dfrbp_1 _13723_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4625),
    .D(net320),
    .Q_N(_06721_),
    .Q(\cpu.current_address[11] ));
 sg13g2_dfrbp_1 _13724_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4638),
    .D(net318),
    .Q_N(_06720_),
    .Q(\cpu.current_address[12] ));
 sg13g2_dfrbp_1 _13725_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4631),
    .D(net325),
    .Q_N(_06719_),
    .Q(\cpu.current_address[13] ));
 sg13g2_dfrbp_1 _13726_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4625),
    .D(net141),
    .Q_N(_06718_),
    .Q(\cpu.current_address[14] ));
 sg13g2_dfrbp_1 _13727_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4631),
    .D(_00650_),
    .Q_N(_06717_),
    .Q(\cpu.current_address[15] ));
 sg13g2_dfrbp_1 _13728_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4649),
    .D(net695),
    .Q_N(_06716_),
    .Q(\cpu.data_out[0] ));
 sg13g2_dfrbp_1 _13729_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4644),
    .D(net394),
    .Q_N(_06715_),
    .Q(\cpu.data_out[1] ));
 sg13g2_dfrbp_1 _13730_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4632),
    .D(net112),
    .Q_N(_06714_),
    .Q(\cpu.data_out[2] ));
 sg13g2_dfrbp_1 _13731_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4645),
    .D(net469),
    .Q_N(_06713_),
    .Q(\cpu.data_out[3] ));
 sg13g2_dfrbp_1 _13732_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4628),
    .D(_00655_),
    .Q_N(_06712_),
    .Q(\cpu.data_out[4] ));
 sg13g2_dfrbp_1 _13733_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net4631),
    .D(_00656_),
    .Q_N(_06711_),
    .Q(\cpu.data_out[5] ));
 sg13g2_dfrbp_1 _13734_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4628),
    .D(_00657_),
    .Q_N(_06710_),
    .Q(\cpu.data_out[6] ));
 sg13g2_dfrbp_1 _13735_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4646),
    .D(net307),
    .Q_N(_06709_),
    .Q(\cpu.data_out[7] ));
 sg13g2_dfrbp_1 _13736_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4644),
    .D(net217),
    .Q_N(_06708_),
    .Q(\cpu.data_out[8] ));
 sg13g2_dfrbp_1 _13737_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4628),
    .D(_00660_),
    .Q_N(_06707_),
    .Q(\cpu.data_out[9] ));
 sg13g2_dfrbp_1 _13738_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net4628),
    .D(_00661_),
    .Q_N(_06706_),
    .Q(\cpu.data_out[10] ));
 sg13g2_dfrbp_1 _13739_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net4635),
    .D(net88),
    .Q_N(_06705_),
    .Q(\cpu.data_out[11] ));
 sg13g2_dfrbp_1 _13740_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4627),
    .D(_00663_),
    .Q_N(_06704_),
    .Q(\cpu.data_out[12] ));
 sg13g2_dfrbp_1 _13741_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4628),
    .D(_00664_),
    .Q_N(_06703_),
    .Q(\cpu.data_out[13] ));
 sg13g2_dfrbp_1 _13742_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4628),
    .D(_00665_),
    .Q_N(_06702_),
    .Q(\cpu.data_out[14] ));
 sg13g2_dfrbp_1 _13743_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net4634),
    .D(net77),
    .Q_N(_06701_),
    .Q(\cpu.data_out[15] ));
 sg13g2_dfrbp_1 _13744_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net4648),
    .D(_00667_),
    .Q_N(_06700_),
    .Q(\cpu.request_type ));
 sg13g2_dfrbp_1 _13745_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4632),
    .D(_00260_),
    .Q_N(\cpu.request ),
    .Q(_00250_));
 sg13g2_dfrbp_1 _13746_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4648),
    .D(_00668_),
    .Q_N(_00149_),
    .Q(\cpu.request_address[0] ));
 sg13g2_dfrbp_1 _13747_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4684),
    .D(net864),
    .Q_N(_00153_),
    .Q(\cpu.request_address[1] ));
 sg13g2_dfrbp_1 _13748_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4678),
    .D(_00670_),
    .Q_N(_00157_),
    .Q(\cpu.request_address[2] ));
 sg13g2_dfrbp_1 _13749_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net4685),
    .D(net892),
    .Q_N(_00161_),
    .Q(\cpu.request_address[3] ));
 sg13g2_dfrbp_1 _13750_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net4685),
    .D(_00672_),
    .Q_N(_00165_),
    .Q(\cpu.request_address[4] ));
 sg13g2_dfrbp_1 _13751_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net4678),
    .D(_00673_),
    .Q_N(_00169_),
    .Q(\cpu.request_address[5] ));
 sg13g2_dfrbp_1 _13752_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net4685),
    .D(_00674_),
    .Q_N(_00173_),
    .Q(\cpu.request_address[6] ));
 sg13g2_dfrbp_1 _13753_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4678),
    .D(_00675_),
    .Q_N(_00177_),
    .Q(\cpu.request_address[7] ));
 sg13g2_dfrbp_1 _13754_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4632),
    .D(_00676_),
    .Q_N(_00181_),
    .Q(\cpu.request_address[8] ));
 sg13g2_dfrbp_1 _13755_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4638),
    .D(_00677_),
    .Q_N(_00185_),
    .Q(\cpu.request_address[9] ));
 sg13g2_dfrbp_1 _13756_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4625),
    .D(net718),
    .Q_N(_00189_),
    .Q(\cpu.request_address[10] ));
 sg13g2_dfrbp_1 _13757_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4625),
    .D(_00679_),
    .Q_N(_00193_),
    .Q(\cpu.request_address[11] ));
 sg13g2_dfrbp_1 _13758_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4644),
    .D(_00680_),
    .Q_N(_00197_),
    .Q(\cpu.request_address[12] ));
 sg13g2_dfrbp_1 _13759_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4631),
    .D(net764),
    .Q_N(_00202_),
    .Q(\cpu.request_address[13] ));
 sg13g2_dfrbp_1 _13760_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4625),
    .D(_00682_),
    .Q_N(_00206_),
    .Q(\cpu.request_address[14] ));
 sg13g2_dfrbp_1 _13761_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net4632),
    .D(_00683_),
    .Q_N(_00210_),
    .Q(\cpu.request_address[15] ));
 sg13g2_dfrbp_1 _13762_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4635),
    .D(_00684_),
    .Q_N(_06699_),
    .Q(\memory_controller.uart_memory_address[10] ));
 sg13g2_dfrbp_1 _13763_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4640),
    .D(net747),
    .Q_N(_00227_),
    .Q(\cpu.registers[5][0] ));
 sg13g2_dfrbp_1 _13764_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4680),
    .D(net423),
    .Q_N(_00228_),
    .Q(\cpu.registers[5][1] ));
 sg13g2_dfrbp_1 _13765_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4641),
    .D(net448),
    .Q_N(_00229_),
    .Q(\cpu.registers[5][2] ));
 sg13g2_dfrbp_1 _13766_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4681),
    .D(net727),
    .Q_N(_00230_),
    .Q(\cpu.registers[5][3] ));
 sg13g2_dfrbp_1 _13767_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4680),
    .D(net596),
    .Q_N(_00231_),
    .Q(\cpu.registers[5][4] ));
 sg13g2_dfrbp_1 _13768_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4676),
    .D(net509),
    .Q_N(_00232_),
    .Q(\cpu.registers[5][5] ));
 sg13g2_dfrbp_1 _13769_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4679),
    .D(net472),
    .Q_N(_00233_),
    .Q(\cpu.registers[5][6] ));
 sg13g2_dfrbp_1 _13770_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4656),
    .D(net592),
    .Q_N(_00234_),
    .Q(\cpu.registers[5][7] ));
 sg13g2_dfrbp_1 _13771_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4601),
    .D(net731),
    .Q_N(_00235_),
    .Q(\cpu.registers[5][8] ));
 sg13g2_dfrbp_1 _13772_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4639),
    .D(net525),
    .Q_N(_00236_),
    .Q(\cpu.registers[5][9] ));
 sg13g2_dfrbp_1 _13773_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4597),
    .D(net772),
    .Q_N(_00237_),
    .Q(\cpu.registers[5][10] ));
 sg13g2_dfrbp_1 _13774_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4602),
    .D(net714),
    .Q_N(_00238_),
    .Q(\cpu.registers[5][11] ));
 sg13g2_dfrbp_1 _13775_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net4613),
    .D(net669),
    .Q_N(_00239_),
    .Q(\cpu.registers[5][12] ));
 sg13g2_dfrbp_1 _13776_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4621),
    .D(net733),
    .Q_N(_00240_),
    .Q(\cpu.registers[5][13] ));
 sg13g2_dfrbp_1 _13777_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4620),
    .D(net692),
    .Q_N(_00241_),
    .Q(\cpu.registers[5][14] ));
 sg13g2_dfrbp_1 _13778_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4621),
    .D(net657),
    .Q_N(_00242_),
    .Q(\cpu.registers[5][15] ));
 sg13g2_dfrbp_1 _13779_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4640),
    .D(net309),
    .Q_N(_00146_),
    .Q(\cpu.registers[6][0] ));
 sg13g2_dfrbp_1 _13780_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net4681),
    .D(net161),
    .Q_N(_00150_),
    .Q(\cpu.registers[6][1] ));
 sg13g2_dfrbp_1 _13781_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4640),
    .D(net163),
    .Q_N(_00154_),
    .Q(\cpu.registers[6][2] ));
 sg13g2_dfrbp_1 _13782_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4687),
    .D(net220),
    .Q_N(_00158_),
    .Q(\cpu.registers[6][3] ));
 sg13g2_dfrbp_1 _13783_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4681),
    .D(net299),
    .Q_N(_00162_),
    .Q(\cpu.registers[6][4] ));
 sg13g2_dfrbp_1 _13784_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4677),
    .D(net365),
    .Q_N(_00166_),
    .Q(\cpu.registers[6][5] ));
 sg13g2_dfrbp_1 _13785_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4679),
    .D(_00707_),
    .Q_N(_00170_),
    .Q(\cpu.registers[6][6] ));
 sg13g2_dfrbp_1 _13786_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net4676),
    .D(net373),
    .Q_N(_00174_),
    .Q(\cpu.registers[6][7] ));
 sg13g2_dfrbp_1 _13787_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4624),
    .D(net335),
    .Q_N(_00178_),
    .Q(\cpu.registers[6][8] ));
 sg13g2_dfrbp_1 _13788_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4637),
    .D(net244),
    .Q_N(_00182_),
    .Q(\cpu.registers[6][9] ));
 sg13g2_dfrbp_1 _13789_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4620),
    .D(net483),
    .Q_N(_00186_),
    .Q(\cpu.registers[6][10] ));
 sg13g2_dfrbp_1 _13790_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4624),
    .D(net367),
    .Q_N(_00190_),
    .Q(\cpu.registers[6][11] ));
 sg13g2_dfrbp_1 _13791_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4637),
    .D(net337),
    .Q_N(_00194_),
    .Q(\cpu.registers[6][12] ));
 sg13g2_dfrbp_1 _13792_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4621),
    .D(net407),
    .Q_N(_00198_),
    .Q(\cpu.registers[6][13] ));
 sg13g2_dfrbp_1 _13793_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4620),
    .D(net513),
    .Q_N(_00203_),
    .Q(\cpu.registers[6][14] ));
 sg13g2_dfrbp_1 _13794_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4621),
    .D(net440),
    .Q_N(_00207_),
    .Q(\cpu.registers[6][15] ));
 sg13g2_dfrbp_1 _13795_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4672),
    .D(_00717_),
    .Q_N(_06698_),
    .Q(\cpu.keccak_alu.registers[256] ));
 sg13g2_dfrbp_1 _13796_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net4670),
    .D(_00718_),
    .Q_N(_06697_),
    .Q(\cpu.keccak_alu.registers[257] ));
 sg13g2_dfrbp_1 _13797_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4670),
    .D(_00719_),
    .Q_N(_06696_),
    .Q(\cpu.keccak_alu.registers[258] ));
 sg13g2_dfrbp_1 _13798_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4671),
    .D(_00720_),
    .Q_N(_06695_),
    .Q(\cpu.keccak_alu.registers[259] ));
 sg13g2_dfrbp_1 _13799_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4660),
    .D(_00721_),
    .Q_N(_06694_),
    .Q(\cpu.keccak_alu.registers[260] ));
 sg13g2_dfrbp_1 _13800_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4657),
    .D(_00722_),
    .Q_N(_06693_),
    .Q(\cpu.keccak_alu.registers[261] ));
 sg13g2_dfrbp_1 _13801_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net4658),
    .D(_00723_),
    .Q_N(_06692_),
    .Q(\cpu.keccak_alu.registers[262] ));
 sg13g2_dfrbp_1 _13802_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net4616),
    .D(_00724_),
    .Q_N(_06691_),
    .Q(\cpu.keccak_alu.registers[263] ));
 sg13g2_dfrbp_1 _13803_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net4605),
    .D(_00725_),
    .Q_N(_06690_),
    .Q(\cpu.keccak_alu.registers[264] ));
 sg13g2_dfrbp_1 _13804_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net4586),
    .D(_00726_),
    .Q_N(_06689_),
    .Q(\cpu.keccak_alu.registers[265] ));
 sg13g2_dfrbp_1 _13805_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4588),
    .D(_00727_),
    .Q_N(_06688_),
    .Q(\cpu.keccak_alu.registers[266] ));
 sg13g2_dfrbp_1 _13806_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net4592),
    .D(_00728_),
    .Q_N(_06687_),
    .Q(\cpu.keccak_alu.registers[267] ));
 sg13g2_dfrbp_1 _13807_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net4607),
    .D(_00729_),
    .Q_N(_06686_),
    .Q(\cpu.keccak_alu.registers[268] ));
 sg13g2_dfrbp_1 _13808_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4597),
    .D(_00730_),
    .Q_N(_06685_),
    .Q(\cpu.keccak_alu.registers[269] ));
 sg13g2_dfrbp_1 _13809_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4588),
    .D(_00731_),
    .Q_N(_06684_),
    .Q(\cpu.keccak_alu.registers[270] ));
 sg13g2_dfrbp_1 _13810_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net4613),
    .D(_00732_),
    .Q_N(_06683_),
    .Q(\cpu.keccak_alu.registers[271] ));
 sg13g2_dfrbp_1 _13811_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4672),
    .D(_00733_),
    .Q_N(_06682_),
    .Q(\cpu.keccak_alu.registers[272] ));
 sg13g2_dfrbp_1 _13812_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4663),
    .D(_00734_),
    .Q_N(_06681_),
    .Q(\cpu.keccak_alu.registers[273] ));
 sg13g2_dfrbp_1 _13813_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net4669),
    .D(_00735_),
    .Q_N(_06680_),
    .Q(\cpu.keccak_alu.registers[274] ));
 sg13g2_dfrbp_1 _13814_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net4671),
    .D(_00736_),
    .Q_N(_06679_),
    .Q(\cpu.keccak_alu.registers[275] ));
 sg13g2_dfrbp_1 _13815_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net4660),
    .D(_00737_),
    .Q_N(_06678_),
    .Q(\cpu.keccak_alu.registers[276] ));
 sg13g2_dfrbp_1 _13816_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4656),
    .D(_00738_),
    .Q_N(_06677_),
    .Q(\cpu.keccak_alu.registers[277] ));
 sg13g2_dfrbp_1 _13817_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4657),
    .D(_00739_),
    .Q_N(_06676_),
    .Q(\cpu.keccak_alu.registers[278] ));
 sg13g2_dfrbp_1 _13818_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net4616),
    .D(_00740_),
    .Q_N(_06675_),
    .Q(\cpu.keccak_alu.registers[279] ));
 sg13g2_dfrbp_1 _13819_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net4606),
    .D(_00741_),
    .Q_N(_06674_),
    .Q(\cpu.keccak_alu.registers[280] ));
 sg13g2_dfrbp_1 _13820_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4588),
    .D(_00742_),
    .Q_N(_06673_),
    .Q(\cpu.keccak_alu.registers[281] ));
 sg13g2_dfrbp_1 _13821_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net4588),
    .D(_00743_),
    .Q_N(_06672_),
    .Q(\cpu.keccak_alu.registers[282] ));
 sg13g2_dfrbp_1 _13822_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4589),
    .D(_00744_),
    .Q_N(_06671_),
    .Q(\cpu.keccak_alu.registers[283] ));
 sg13g2_dfrbp_1 _13823_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net4609),
    .D(_00745_),
    .Q_N(_06670_),
    .Q(\cpu.keccak_alu.registers[284] ));
 sg13g2_dfrbp_1 _13824_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4597),
    .D(_00746_),
    .Q_N(_06669_),
    .Q(\cpu.keccak_alu.registers[285] ));
 sg13g2_dfrbp_1 _13825_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net4595),
    .D(_00747_),
    .Q_N(_06668_),
    .Q(\cpu.keccak_alu.registers[286] ));
 sg13g2_dfrbp_1 _13826_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net4613),
    .D(_00748_),
    .Q_N(_06667_),
    .Q(\cpu.keccak_alu.registers[287] ));
 sg13g2_dfrbp_1 _13827_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4689),
    .D(_00749_),
    .Q_N(_06666_),
    .Q(\cpu.keccak_alu.registers[288] ));
 sg13g2_dfrbp_1 _13828_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4669),
    .D(_00750_),
    .Q_N(_06665_),
    .Q(\cpu.keccak_alu.registers[289] ));
 sg13g2_dfrbp_1 _13829_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4666),
    .D(_00751_),
    .Q_N(_06664_),
    .Q(\cpu.keccak_alu.registers[290] ));
 sg13g2_dfrbp_1 _13830_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4667),
    .D(_00752_),
    .Q_N(_06663_),
    .Q(\cpu.keccak_alu.registers[291] ));
 sg13g2_dfrbp_1 _13831_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4660),
    .D(_00753_),
    .Q_N(_06662_),
    .Q(\cpu.keccak_alu.registers[292] ));
 sg13g2_dfrbp_1 _13832_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4656),
    .D(_00754_),
    .Q_N(_06661_),
    .Q(\cpu.keccak_alu.registers[293] ));
 sg13g2_dfrbp_1 _13833_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net4657),
    .D(_00755_),
    .Q_N(_06660_),
    .Q(\cpu.keccak_alu.registers[294] ));
 sg13g2_dfrbp_1 _13834_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net4617),
    .D(_00756_),
    .Q_N(_06659_),
    .Q(\cpu.keccak_alu.registers[295] ));
 sg13g2_dfrbp_1 _13835_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net4610),
    .D(_00757_),
    .Q_N(_06658_),
    .Q(\cpu.keccak_alu.registers[296] ));
 sg13g2_dfrbp_1 _13836_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4593),
    .D(_00758_),
    .Q_N(_06657_),
    .Q(\cpu.keccak_alu.registers[297] ));
 sg13g2_dfrbp_1 _13837_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4593),
    .D(_00759_),
    .Q_N(_06656_),
    .Q(\cpu.keccak_alu.registers[298] ));
 sg13g2_dfrbp_1 _13838_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4594),
    .D(_00760_),
    .Q_N(_06655_),
    .Q(\cpu.keccak_alu.registers[299] ));
 sg13g2_dfrbp_1 _13839_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net4609),
    .D(net673),
    .Q_N(_06654_),
    .Q(\cpu.keccak_alu.registers[300] ));
 sg13g2_dfrbp_1 _13840_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4601),
    .D(_00762_),
    .Q_N(_06653_),
    .Q(\cpu.keccak_alu.registers[301] ));
 sg13g2_dfrbp_1 _13841_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net4599),
    .D(_00763_),
    .Q_N(_06652_),
    .Q(\cpu.keccak_alu.registers[302] ));
 sg13g2_dfrbp_1 _13842_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net4602),
    .D(_00764_),
    .Q_N(_06651_),
    .Q(\cpu.keccak_alu.registers[303] ));
 sg13g2_dfrbp_1 _13843_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4689),
    .D(_00765_),
    .Q_N(_06650_),
    .Q(\cpu.keccak_alu.registers[304] ));
 sg13g2_dfrbp_1 _13844_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net4674),
    .D(_00766_),
    .Q_N(_06649_),
    .Q(\cpu.keccak_alu.registers[305] ));
 sg13g2_dfrbp_1 _13845_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4669),
    .D(_00767_),
    .Q_N(_06648_),
    .Q(\cpu.keccak_alu.registers[306] ));
 sg13g2_dfrbp_1 _13846_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net4672),
    .D(_00768_),
    .Q_N(_06647_),
    .Q(\cpu.keccak_alu.registers[307] ));
 sg13g2_dfrbp_1 _13847_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4679),
    .D(_00769_),
    .Q_N(_06646_),
    .Q(\cpu.keccak_alu.registers[308] ));
 sg13g2_dfrbp_1 _13848_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4656),
    .D(_00770_),
    .Q_N(_06645_),
    .Q(\cpu.keccak_alu.registers[309] ));
 sg13g2_dfrbp_1 _13849_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net4656),
    .D(_00771_),
    .Q_N(_06644_),
    .Q(\cpu.keccak_alu.registers[310] ));
 sg13g2_dfrbp_1 _13850_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net4617),
    .D(_00772_),
    .Q_N(_06643_),
    .Q(\cpu.keccak_alu.registers[311] ));
 sg13g2_dfrbp_1 _13851_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net4610),
    .D(_00773_),
    .Q_N(_06642_),
    .Q(\cpu.keccak_alu.registers[312] ));
 sg13g2_dfrbp_1 _13852_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net4587),
    .D(_00774_),
    .Q_N(_06641_),
    .Q(\cpu.keccak_alu.registers[313] ));
 sg13g2_dfrbp_1 _13853_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net4589),
    .D(_00775_),
    .Q_N(_06640_),
    .Q(\cpu.keccak_alu.registers[314] ));
 sg13g2_dfrbp_1 _13854_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net4594),
    .D(_00776_),
    .Q_N(_06639_),
    .Q(\cpu.keccak_alu.registers[315] ));
 sg13g2_dfrbp_1 _13855_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net4607),
    .D(_00777_),
    .Q_N(_06638_),
    .Q(\cpu.keccak_alu.registers[316] ));
 sg13g2_dfrbp_1 _13856_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net4597),
    .D(_00778_),
    .Q_N(_06637_),
    .Q(\cpu.keccak_alu.registers[317] ));
 sg13g2_dfrbp_1 _13857_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net4594),
    .D(_00779_),
    .Q_N(_06636_),
    .Q(\cpu.keccak_alu.registers[318] ));
 sg13g2_dfrbp_1 _13858_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net4602),
    .D(_00780_),
    .Q_N(_06975_),
    .Q(\cpu.keccak_alu.registers[319] ));
 sg13g2_dfrbp_1 _13859_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net4642),
    .D(_06992_),
    .Q_N(_06976_),
    .Q(\cpu.registers[1][0] ));
 sg13g2_dfrbp_1 _13860_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4642),
    .D(net879),
    .Q_N(_00152_),
    .Q(\cpu.registers[1][1] ));
 sg13g2_dfrbp_1 _13861_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4635),
    .D(_00781_),
    .Q_N(_06635_),
    .Q(\memory_controller.register_enable ));
 sg13g2_dfrbp_1 _13862_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4633),
    .D(_00782_),
    .Q_N(_06634_),
    .Q(\memory_controller.upper_bit ));
 sg13g2_dfrbp_1 _13863_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4633),
    .D(net382),
    .Q_N(_06633_),
    .Q(\memory_controller.write_enable ));
 sg13g2_dfrbp_1 _13864_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4633),
    .D(_00784_),
    .Q_N(_06632_),
    .Q(lower_bit));
 sg13g2_dfrbp_1 _13865_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4645),
    .D(_00785_),
    .Q_N(_00130_),
    .Q(\cpu.memory_in[0] ));
 sg13g2_dfrbp_1 _13866_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4643),
    .D(_00786_),
    .Q_N(_00131_),
    .Q(\cpu.memory_in[1] ));
 sg13g2_dfrbp_1 _13867_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4647),
    .D(_00787_),
    .Q_N(_00132_),
    .Q(\cpu.memory_in[2] ));
 sg13g2_dfrbp_1 _13868_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net4645),
    .D(_00788_),
    .Q_N(_00133_),
    .Q(\cpu.memory_in[3] ));
 sg13g2_dfrbp_1 _13869_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4643),
    .D(_00789_),
    .Q_N(_00134_),
    .Q(\cpu.memory_in[4] ));
 sg13g2_dfrbp_1 _13870_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4647),
    .D(_00790_),
    .Q_N(_00135_),
    .Q(\cpu.memory_in[5] ));
 sg13g2_dfrbp_1 _13871_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4644),
    .D(_00791_),
    .Q_N(_00136_),
    .Q(\cpu.memory_in[6] ));
 sg13g2_dfrbp_1 _13872_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4643),
    .D(_00792_),
    .Q_N(_00137_),
    .Q(\cpu.memory_in[7] ));
 sg13g2_dfrbp_1 _13873_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4631),
    .D(net315),
    .Q_N(_00020_),
    .Q(\cpu.write_complete ));
 sg13g2_dfrbp_1 _13874_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4629),
    .D(net21),
    .Q_N(_06977_),
    .Q(\memory_controller.state[0] ));
 sg13g2_dfrbp_1 _13875_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4629),
    .D(net19),
    .Q_N(_06978_),
    .Q(\memory_controller.state[1] ));
 sg13g2_dfrbp_1 _13876_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net4631),
    .D(net22),
    .Q_N(_06979_),
    .Q(\memory_controller.state[2] ));
 sg13g2_dfrbp_1 _13877_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4631),
    .D(net20),
    .Q_N(_06980_),
    .Q(\memory_controller.state[3] ));
 sg13g2_dfrbp_1 _13878_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4634),
    .D(net23),
    .Q_N(_00019_),
    .Q(\memory_controller.state[4] ));
 sg13g2_dfrbp_1 _13879_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4631),
    .D(_00794_),
    .Q_N(_00022_),
    .Q(\cpu.memory_ready ));
 sg13g2_dfrbp_1 _13880_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4627),
    .D(_00010_),
    .Q_N(_06981_),
    .Q(\memory_controller.wait_counter[0] ));
 sg13g2_dfrbp_1 _13881_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4627),
    .D(_00011_),
    .Q_N(_06982_),
    .Q(\memory_controller.wait_counter[1] ));
 sg13g2_dfrbp_1 _13882_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4627),
    .D(net170),
    .Q_N(_06983_),
    .Q(\memory_controller.wait_counter[2] ));
 sg13g2_dfrbp_1 _13883_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4627),
    .D(_00013_),
    .Q_N(_06984_),
    .Q(\memory_controller.wait_counter[3] ));
 sg13g2_dfrbp_1 _13884_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4627),
    .D(_00014_),
    .Q_N(_06985_),
    .Q(\memory_controller.wait_counter[4] ));
 sg13g2_dfrbp_1 _13885_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net4627),
    .D(_00015_),
    .Q_N(_06631_),
    .Q(\memory_controller.wait_counter[5] ));
 sg13g2_dfrbp_1 _13886_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net4633),
    .D(_00795_),
    .Q_N(_06630_),
    .Q(uio_oe[7]));
 sg13g2_dfrbp_1 _13887_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net4633),
    .D(_00796_),
    .Q_N(_06629_),
    .Q(\memory_controller.read_enable ));
 sg13g2_dfrbp_1 _13888_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net4629),
    .D(net794),
    .Q_N(_06628_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _13889_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4629),
    .D(net721),
    .Q_N(_06627_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _13890_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net4630),
    .D(_00799_),
    .Q_N(_06626_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _13891_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4629),
    .D(net750),
    .Q_N(_06625_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _13892_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4629),
    .D(_00801_),
    .Q_N(_06624_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _13893_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net4630),
    .D(_00802_),
    .Q_N(_06623_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _13894_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net4630),
    .D(_00803_),
    .Q_N(_06622_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _13895_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net4629),
    .D(net723),
    .Q_N(_06621_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _13896_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4699),
    .D(net259),
    .Q_N(_06620_),
    .Q(\cpu.uart.data_sending[0] ));
 sg13g2_dfrbp_1 _13897_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4698),
    .D(net253),
    .Q_N(_06619_),
    .Q(\cpu.uart.data_sending[1] ));
 sg13g2_dfrbp_1 _13898_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4698),
    .D(net246),
    .Q_N(_06618_),
    .Q(\cpu.uart.data_sending[2] ));
 sg13g2_dfrbp_1 _13899_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4698),
    .D(net234),
    .Q_N(_06617_),
    .Q(\cpu.uart.data_sending[3] ));
 sg13g2_dfrbp_1 _13900_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net4698),
    .D(net215),
    .Q_N(_06616_),
    .Q(\cpu.uart.data_sending[4] ));
 sg13g2_dfrbp_1 _13901_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4697),
    .D(_00810_),
    .Q_N(_06615_),
    .Q(\cpu.uart.data_sending[5] ));
 sg13g2_dfrbp_1 _13902_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4696),
    .D(net345),
    .Q_N(_06614_),
    .Q(\cpu.uart.data_sending[6] ));
 sg13g2_dfrbp_1 _13903_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4697),
    .D(net213),
    .Q_N(_06613_),
    .Q(\cpu.uart.data_sending[7] ));
 sg13g2_dfrbp_1 _13904_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4651),
    .D(net46),
    .Q_N(\cpu.execution_stage[0] ),
    .Q(_00251_));
 sg13g2_dfrbp_1 _13905_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4648),
    .D(net934),
    .Q_N(_00045_),
    .Q(\cpu.execution_stage[1] ));
 sg13g2_dfrbp_1 _13906_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4643),
    .D(_00002_),
    .Q_N(_00016_),
    .Q(\cpu.execution_stage[2] ));
 sg13g2_dfrbp_1 _13907_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net4648),
    .D(_00003_),
    .Q_N(_00018_),
    .Q(\cpu.execution_stage[3] ));
 sg13g2_dfrbp_1 _13908_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net4684),
    .D(net4024),
    .Q_N(_06986_),
    .Q(\cpu.execution_stage[4] ));
 sg13g2_dfrbp_1 _13909_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net4642),
    .D(net832),
    .Q_N(_00021_),
    .Q(\cpu.execution_stage[5] ));
 sg13g2_dfrbp_1 _13910_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net4676),
    .D(net240),
    .Q_N(_00168_),
    .Q(\cpu.registers[1][5] ));
 sg13g2_dfrbp_1 _13911_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4679),
    .D(net256),
    .Q_N(_00172_),
    .Q(\cpu.registers[1][6] ));
 sg13g2_dfrbp_1 _13912_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net4676),
    .D(net291),
    .Q_N(_00176_),
    .Q(\cpu.registers[1][7] ));
 sg13g2_dfrbp_1 _13913_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4624),
    .D(net354),
    .Q_N(_00180_),
    .Q(\cpu.registers[1][8] ));
 sg13g2_dfrbp_1 _13914_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4637),
    .D(net228),
    .Q_N(_00184_),
    .Q(\cpu.registers[1][9] ));
 sg13g2_dfrbp_1 _13915_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4620),
    .D(net303),
    .Q_N(_00188_),
    .Q(\cpu.registers[1][10] ));
 sg13g2_dfrbp_1 _13916_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net4626),
    .D(net287),
    .Q_N(_00192_),
    .Q(\cpu.registers[1][11] ));
 sg13g2_dfrbp_1 _13917_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net4637),
    .D(net371),
    .Q_N(_00196_),
    .Q(\cpu.registers[1][12] ));
 sg13g2_dfrbp_1 _13918_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4622),
    .D(net363),
    .Q_N(_00200_),
    .Q(\cpu.registers[1][13] ));
 sg13g2_dfrbp_1 _13919_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4622),
    .D(net285),
    .Q_N(_00205_),
    .Q(\cpu.registers[1][14] ));
 sg13g2_dfrbp_1 _13920_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net4622),
    .D(net446),
    .Q_N(_00209_),
    .Q(\cpu.registers[1][15] ));
 sg13g2_dfrbp_1 _13921_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net4644),
    .D(_00824_),
    .Q_N(_00138_),
    .Q(\cpu.memory_in[8] ));
 sg13g2_dfrbp_1 _13922_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4638),
    .D(_00825_),
    .Q_N(_00139_),
    .Q(\cpu.memory_in[9] ));
 sg13g2_dfrbp_1 _13923_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4646),
    .D(_00826_),
    .Q_N(_00140_),
    .Q(\cpu.memory_in[10] ));
 sg13g2_dfrbp_1 _13924_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net4646),
    .D(_00827_),
    .Q_N(_00141_),
    .Q(\cpu.memory_in[11] ));
 sg13g2_dfrbp_1 _13925_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4644),
    .D(_00828_),
    .Q_N(_00142_),
    .Q(\cpu.memory_in[12] ));
 sg13g2_dfrbp_1 _13926_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net4646),
    .D(_00829_),
    .Q_N(_00143_),
    .Q(\cpu.memory_in[13] ));
 sg13g2_dfrbp_1 _13927_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net4638),
    .D(_00830_),
    .Q_N(_00144_),
    .Q(\cpu.memory_in[14] ));
 sg13g2_dfrbp_1 _13928_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net4644),
    .D(_00831_),
    .Q_N(_00145_),
    .Q(\cpu.memory_in[15] ));
 sg13g2_dfrbp_1 _13929_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net18),
    .D(_00832_),
    .Q_N(_06612_),
    .Q(\memory_controller.next_state[4] ));
 sg13g2_dfrbp_1 _13930_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net17),
    .D(_00833_),
    .Q_N(_06611_),
    .Q(\memory_controller.next_state[3] ));
 sg13g2_dfrbp_1 _13931_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net16),
    .D(_00834_),
    .Q_N(_06610_),
    .Q(\memory_controller.next_state[2] ));
 sg13g2_dfrbp_1 _13932_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net15),
    .D(_00835_),
    .Q_N(_06609_),
    .Q(\memory_controller.next_state[1] ));
 sg13g2_dfrbp_1 _13933_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net14),
    .D(_00836_),
    .Q_N(_06608_),
    .Q(\memory_controller.next_state[0] ));
 sg13g2_dfrbp_1 _13934_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4692),
    .D(net31),
    .Q_N(\cpu.uart.stage[0] ),
    .Q(_00252_));
 sg13g2_dfrbp_1 _13935_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4696),
    .D(net818),
    .Q_N(_00007_),
    .Q(\cpu.uart.stage[1] ));
 sg13g2_dfrbp_1 _13936_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4696),
    .D(_00006_),
    .Q_N(_00028_),
    .Q(\cpu.uart.stage[2] ));
 sg13g2_dfrbp_1 _13937_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4696),
    .D(net589),
    .Q_N(_00023_),
    .Q(\cpu.uart.busy ));
 sg13g2_dfrbp_1 _13938_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4640),
    .D(net348),
    .Q_N(_00243_),
    .Q(\cpu.registers[7][0] ));
 sg13g2_dfrbp_1 _13939_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4680),
    .D(net51),
    .Q_N(_00031_),
    .Q(\cpu.registers[7][1] ));
 sg13g2_dfrbp_1 _13940_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net4641),
    .D(_00840_),
    .Q_N(_00032_),
    .Q(\cpu.registers[7][2] ));
 sg13g2_dfrbp_1 _13941_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4680),
    .D(_00841_),
    .Q_N(_00033_),
    .Q(\cpu.registers[7][3] ));
 sg13g2_dfrbp_1 _13942_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net4681),
    .D(_00842_),
    .Q_N(_00034_),
    .Q(\cpu.registers[7][4] ));
 sg13g2_dfrbp_1 _13943_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net4677),
    .D(_00843_),
    .Q_N(_00035_),
    .Q(\cpu.registers[7][5] ));
 sg13g2_dfrbp_1 _13944_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net4679),
    .D(_00844_),
    .Q_N(_00036_),
    .Q(\cpu.registers[7][6] ));
 sg13g2_dfrbp_1 _13945_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net4676),
    .D(_00845_),
    .Q_N(_00037_),
    .Q(\cpu.registers[7][7] ));
 sg13g2_dfrbp_1 _13946_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4624),
    .D(_00846_),
    .Q_N(_00038_),
    .Q(\cpu.registers[7][8] ));
 sg13g2_dfrbp_1 _13947_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4639),
    .D(_00847_),
    .Q_N(_00039_),
    .Q(\cpu.registers[7][9] ));
 sg13g2_dfrbp_1 _13948_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net4623),
    .D(_00848_),
    .Q_N(_00040_),
    .Q(\cpu.registers[7][10] ));
 sg13g2_dfrbp_1 _13949_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net4626),
    .D(_00849_),
    .Q_N(_00041_),
    .Q(\cpu.registers[7][11] ));
 sg13g2_dfrbp_1 _13950_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net4637),
    .D(_00850_),
    .Q_N(_00042_),
    .Q(\cpu.registers[7][12] ));
 sg13g2_dfrbp_1 _13951_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4621),
    .D(_00851_),
    .Q_N(_00046_),
    .Q(\cpu.registers[7][13] ));
 sg13g2_dfrbp_1 _13952_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net4621),
    .D(_00852_),
    .Q_N(_00047_),
    .Q(\cpu.registers[7][14] ));
 sg13g2_dfrbp_1 _13953_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net4621),
    .D(_00853_),
    .Q_N(_00048_),
    .Q(\cpu.registers[7][15] ));
 sg13g2_dfrbp_1 _13954_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4694),
    .D(net392),
    .Q_N(_06607_),
    .Q(\cpu.uart.cycle_counter[0] ));
 sg13g2_dfrbp_1 _13955_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4694),
    .D(net266),
    .Q_N(_06606_),
    .Q(\cpu.uart.cycle_counter[1] ));
 sg13g2_dfrbp_1 _13956_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4694),
    .D(_00856_),
    .Q_N(_06605_),
    .Q(\cpu.uart.cycle_counter[2] ));
 sg13g2_dfrbp_1 _13957_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4694),
    .D(net119),
    .Q_N(_06604_),
    .Q(\cpu.uart.cycle_counter[3] ));
 sg13g2_dfrbp_1 _13958_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4694),
    .D(_00858_),
    .Q_N(_06603_),
    .Q(\cpu.uart.cycle_counter[4] ));
 sg13g2_dfrbp_1 _13959_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4694),
    .D(_00859_),
    .Q_N(_06602_),
    .Q(\cpu.uart.cycle_counter[5] ));
 sg13g2_dfrbp_1 _13960_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4695),
    .D(_00860_),
    .Q_N(_06601_),
    .Q(\cpu.uart.cycle_counter[6] ));
 sg13g2_dfrbp_1 _13961_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4695),
    .D(net115),
    .Q_N(_06600_),
    .Q(\cpu.uart.cycle_counter[7] ));
 sg13g2_dfrbp_1 _13962_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4690),
    .D(_00862_),
    .Q_N(_06599_),
    .Q(\cpu.uart.cycle_counter[8] ));
 sg13g2_dfrbp_1 _13963_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4690),
    .D(net280),
    .Q_N(_06598_),
    .Q(\cpu.uart.cycle_counter[9] ));
 sg13g2_dfrbp_1 _13964_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4690),
    .D(_00864_),
    .Q_N(_06597_),
    .Q(\cpu.uart.cycle_counter[10] ));
 sg13g2_dfrbp_1 _13965_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4690),
    .D(_00865_),
    .Q_N(_06596_),
    .Q(\cpu.uart.cycle_counter[11] ));
 sg13g2_dfrbp_1 _13966_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4690),
    .D(_00866_),
    .Q_N(_06595_),
    .Q(\cpu.uart.cycle_counter[12] ));
 sg13g2_dfrbp_1 _13967_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4695),
    .D(net185),
    .Q_N(_06594_),
    .Q(\cpu.uart.cycles_per_bit[0] ));
 sg13g2_dfrbp_1 _13968_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4691),
    .D(net29),
    .Q_N(\cpu.uart.cycles_per_bit[1] ),
    .Q(_00253_));
 sg13g2_dfrbp_1 _13969_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4694),
    .D(net199),
    .Q_N(_06593_),
    .Q(\cpu.uart.cycles_per_bit[2] ));
 sg13g2_dfrbp_1 _13970_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4695),
    .D(net27),
    .Q_N(\cpu.uart.cycles_per_bit[3] ),
    .Q(_00254_));
 sg13g2_dfrbp_1 _13971_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4694),
    .D(net188),
    .Q_N(_06592_),
    .Q(\cpu.uart.cycles_per_bit[4] ));
 sg13g2_dfrbp_1 _13972_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4693),
    .D(net38),
    .Q_N(\cpu.uart.cycles_per_bit[5] ),
    .Q(_00255_));
 sg13g2_dfrbp_1 _13973_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4691),
    .D(net33),
    .Q_N(\cpu.uart.cycles_per_bit[6] ),
    .Q(_00256_));
 sg13g2_dfrbp_1 _13974_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net4691),
    .D(net289),
    .Q_N(_06591_),
    .Q(\cpu.uart.cycles_per_bit[7] ));
 sg13g2_dfrbp_1 _13975_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net4691),
    .D(net230),
    .Q_N(_06590_),
    .Q(\cpu.uart.cycles_per_bit[8] ));
 sg13g2_dfrbp_1 _13976_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4689),
    .D(_00876_),
    .Q_N(_06589_),
    .Q(\cpu.uart.cycles_per_bit[9] ));
 sg13g2_dfrbp_1 _13977_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4689),
    .D(net377),
    .Q_N(_06588_),
    .Q(\cpu.uart.cycles_per_bit[10] ));
 sg13g2_dfrbp_1 _13978_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net4691),
    .D(net25),
    .Q_N(\cpu.uart.cycles_per_bit[11] ),
    .Q(_00257_));
 sg13g2_dfrbp_1 _13979_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net4690),
    .D(net40),
    .Q_N(\cpu.uart.cycles_per_bit[12] ),
    .Q(_00258_));
 sg13g2_dfrbp_1 _13980_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net4696),
    .D(net36),
    .Q_N(\cpu.tx ),
    .Q(_00259_));
 sg13g2_dfrbp_1 _13981_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4697),
    .D(net919),
    .Q_N(_06587_),
    .Q(\cpu.uart.bit_counter[0] ));
 sg13g2_dfrbp_1 _13982_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net4697),
    .D(net845),
    .Q_N(_06586_),
    .Q(\cpu.uart.bit_counter[1] ));
 sg13g2_dfrbp_1 _13983_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net4696),
    .D(net581),
    .Q_N(_00029_),
    .Q(\cpu.uart.bit_counter[2] ));
 sg13g2_tiehi _13932__15 (.L_HI(net15));
 sg13g2_tiehi _13931__16 (.L_HI(net16));
 sg13g2_tiehi _13930__17 (.L_HI(net17));
 sg13g2_tiehi _13929__18 (.L_HI(net18));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_zoom_zoom_13 (.L_LO(net13));
 sg13g2_tiehi _13933__14 (.L_HI(net14));
 sg13g2_buf_1 _13991_ (.A(uio_oe[7]),
    .X(uio_oe[0]));
 sg13g2_buf_1 _13992_ (.A(uio_oe[7]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _13993_ (.A(uio_oe[7]),
    .X(uio_oe[2]));
 sg13g2_buf_2 _13994_ (.A(uio_oe[7]),
    .X(uio_oe[3]));
 sg13g2_buf_2 _13995_ (.A(uio_oe[7]),
    .X(uio_oe[4]));
 sg13g2_buf_2 _13996_ (.A(uio_oe[7]),
    .X(uio_oe[5]));
 sg13g2_buf_2 _13997_ (.A(uio_oe[7]),
    .X(uio_oe[6]));
 sg13g2_buf_1 _13998_ (.A(\memory_controller.write_enable ),
    .X(uo_out[0]));
 sg13g2_buf_1 _13999_ (.A(\memory_controller.register_enable ),
    .X(uo_out[1]));
 sg13g2_buf_1 _14000_ (.A(\memory_controller.read_enable ),
    .X(uo_out[2]));
 sg13g2_buf_1 _14001_ (.A(lower_bit),
    .X(uo_out[3]));
 sg13g2_buf_4 _14002_ (.X(uo_out[4]),
    .A(\cpu.tx ));
 sg13g2_buf_1 _14003_ (.A(\memory_controller.upper_bit ),
    .X(uo_out[5]));
 sg13g2_inv_1 \uart_receiver/_334_  (.Y(\uart_receiver/_108_ ),
    .A(\uart_receiver/bit_counter[2] ));
 sg13g2_inv_1 \uart_receiver/_335_  (.Y(\uart_receiver/_109_ ),
    .A(net154));
 sg13g2_inv_1 \uart_receiver/_336_  (.Y(\uart_receiver/_110_ ),
    .A(net821));
 sg13g2_inv_1 \uart_receiver/_337_  (.Y(\uart_receiver/_111_ ),
    .A(net806));
 sg13g2_inv_1 \uart_receiver/_338_  (.Y(\uart_receiver/_112_ ),
    .A(\uart_receiver/cycle_counter[10] ));
 sg13g2_inv_1 \uart_receiver/_339_  (.Y(\uart_receiver/_113_ ),
    .A(net709));
 sg13g2_inv_1 \uart_receiver/_340_  (.Y(\uart_receiver/_114_ ),
    .A(net781));
 sg13g2_inv_1 \uart_receiver/_341_  (.Y(\uart_receiver/_115_ ),
    .A(net698));
 sg13g2_inv_1 \uart_receiver/_342_  (.Y(\uart_receiver/_116_ ),
    .A(net795));
 sg13g2_inv_1 \uart_receiver/_343_  (.Y(\uart_receiver/_117_ ),
    .A(\uart_receiver/cycle_counter[5] ));
 sg13g2_inv_1 \uart_receiver/_344_  (.Y(\uart_receiver/_118_ ),
    .A(\uart_receiver/cycle_counter[4] ));
 sg13g2_inv_1 \uart_receiver/_345_  (.Y(\uart_receiver/_119_ ),
    .A(net701));
 sg13g2_inv_1 \uart_receiver/_346_  (.Y(\uart_receiver/_120_ ),
    .A(net881));
 sg13g2_inv_1 \uart_receiver/_347_  (.Y(\uart_receiver/_121_ ),
    .A(net835));
 sg13g2_inv_1 \uart_receiver/_348_  (.Y(\uart_receiver/_122_ ),
    .A(net826));
 sg13g2_inv_1 \uart_receiver/_349_  (.Y(\uart_receiver/_123_ ),
    .A(\uart_receiver/cycles_per_bit[10] ));
 sg13g2_inv_1 \uart_receiver/_350_  (.Y(\uart_receiver/_124_ ),
    .A(\uart_receiver/cycles_per_bit[4] ));
 sg13g2_inv_1 \uart_receiver/_351_  (.Y(\uart_receiver/_125_ ),
    .A(\uart_receiver/cycles_per_bit[2] ));
 sg13g2_inv_1 \uart_receiver/_352_  (.Y(\uart_receiver/_126_ ),
    .A(\uart_receiver/stage[1] ));
 sg13g2_inv_1 \uart_receiver/_353_  (.Y(\uart_receiver/_127_ ),
    .A(\uart_receiver/stage[2] ));
 sg13g2_inv_1 \uart_receiver/_354_  (.Y(\uart_receiver/_012_ ),
    .A(net4581));
 sg13g2_o21ai_1 \uart_receiver/_355_  (.B1(net521),
    .Y(\uart_receiver/_128_ ),
    .A1(net4481),
    .A2(net3));
 sg13g2_nor2b_1 \uart_receiver/_356_  (.A(\uart_receiver/cycles_per_bit[11] ),
    .B_N(\uart_receiver/cycle_counter[11] ),
    .Y(\uart_receiver/_129_ ));
 sg13g2_xor2_1 \uart_receiver/_357_  (.B(\uart_receiver/cycles_per_bit[12] ),
    .A(\uart_receiver/cycle_counter[12] ),
    .X(\uart_receiver/_130_ ));
 sg13g2_xor2_1 \uart_receiver/_358_  (.B(\uart_receiver/cycles_per_bit[3] ),
    .A(\uart_receiver/cycle_counter[3] ),
    .X(\uart_receiver/_131_ ));
 sg13g2_xor2_1 \uart_receiver/_359_  (.B(\uart_receiver/cycles_per_bit[8] ),
    .A(\uart_receiver/cycle_counter[8] ),
    .X(\uart_receiver/_132_ ));
 sg13g2_xor2_1 \uart_receiver/_360_  (.B(\uart_receiver/cycles_per_bit[5] ),
    .A(\uart_receiver/cycle_counter[5] ),
    .X(\uart_receiver/_133_ ));
 sg13g2_nor2_1 \uart_receiver/_361_  (.A(\uart_receiver/_132_ ),
    .B(\uart_receiver/_133_ ),
    .Y(\uart_receiver/_134_ ));
 sg13g2_xnor2_1 \uart_receiver/_362_  (.Y(\uart_receiver/_135_ ),
    .A(\uart_receiver/cycle_counter[0] ),
    .B(\uart_receiver/cycles_per_bit[0] ));
 sg13g2_xor2_1 \uart_receiver/_363_  (.B(\uart_receiver/cycles_per_bit[4] ),
    .A(\uart_receiver/cycle_counter[4] ),
    .X(\uart_receiver/_136_ ));
 sg13g2_a22oi_1 \uart_receiver/_364_  (.Y(\uart_receiver/_137_ ),
    .B1(\uart_receiver/cycles_per_bit[6] ),
    .B2(\uart_receiver/_116_ ),
    .A2(\uart_receiver/cycles_per_bit[10] ),
    .A1(\uart_receiver/_112_ ));
 sg13g2_nor2b_1 \uart_receiver/_365_  (.A(\uart_receiver/cycles_per_bit[6] ),
    .B_N(\uart_receiver/cycle_counter[6] ),
    .Y(\uart_receiver/_138_ ));
 sg13g2_xnor2_1 \uart_receiver/_366_  (.Y(\uart_receiver/_139_ ),
    .A(\uart_receiver/cycle_counter[9] ),
    .B(\uart_receiver/cycles_per_bit[9] ));
 sg13g2_xor2_1 \uart_receiver/_367_  (.B(\uart_receiver/cycles_per_bit[7] ),
    .A(\uart_receiver/cycle_counter[7] ),
    .X(\uart_receiver/_140_ ));
 sg13g2_xor2_1 \uart_receiver/_368_  (.B(\uart_receiver/cycles_per_bit[1] ),
    .A(\uart_receiver/cycle_counter[1] ),
    .X(\uart_receiver/_141_ ));
 sg13g2_a221oi_1 \uart_receiver/_369_  (.B2(\uart_receiver/_111_ ),
    .C1(\uart_receiver/_140_ ),
    .B1(\uart_receiver/cycles_per_bit[11] ),
    .A1(\uart_receiver/cycle_counter[2] ),
    .Y(\uart_receiver/_142_ ),
    .A2(\uart_receiver/_125_ ));
 sg13g2_and4_2 \uart_receiver/_370_  (.A(\uart_receiver/_134_ ),
    .B(\uart_receiver/_135_ ),
    .C(\uart_receiver/_139_ ),
    .D(\uart_receiver/_142_ ),
    .X(\uart_receiver/_143_ ));
 sg13g2_nor2_1 \uart_receiver/_371_  (.A(\uart_receiver/_130_ ),
    .B(\uart_receiver/_136_ ),
    .Y(\uart_receiver/_144_ ));
 sg13g2_a22oi_1 \uart_receiver/_372_  (.Y(\uart_receiver/_145_ ),
    .B1(\uart_receiver/cycles_per_bit[2] ),
    .B2(\uart_receiver/_120_ ),
    .A2(\uart_receiver/_123_ ),
    .A1(\uart_receiver/cycle_counter[10] ));
 sg13g2_nor4_1 \uart_receiver/_373_  (.A(\uart_receiver/_129_ ),
    .B(\uart_receiver/_131_ ),
    .C(\uart_receiver/_138_ ),
    .D(\uart_receiver/_141_ ),
    .Y(\uart_receiver/_146_ ));
 sg13g2_and4_2 \uart_receiver/_374_  (.A(\uart_receiver/_137_ ),
    .B(\uart_receiver/_144_ ),
    .C(\uart_receiver/_145_ ),
    .D(\uart_receiver/_146_ ),
    .X(\uart_receiver/_147_ ));
 sg13g2_and2_1 \uart_receiver/_375_  (.A(\uart_receiver/_143_ ),
    .B(\uart_receiver/_147_ ),
    .X(\uart_receiver/_148_ ));
 sg13g2_nand2_2 \uart_receiver/_376_  (.Y(\uart_receiver/_149_ ),
    .A(\uart_receiver/_143_ ),
    .B(\uart_receiver/_147_ ));
 sg13g2_nor3_2 \uart_receiver/_377_  (.A(net4481),
    .B(\uart_receiver/_126_ ),
    .C(\uart_receiver/_149_ ),
    .Y(\uart_receiver/_150_ ));
 sg13g2_nor2_2 \uart_receiver/_378_  (.A(net4481),
    .B(\uart_receiver/_149_ ),
    .Y(\uart_receiver/_151_ ));
 sg13g2_nor2b_1 \uart_receiver/_379_  (.A(net3717),
    .B_N(\uart_receiver/_128_ ),
    .Y(\uart_receiver/_058_ ));
 sg13g2_nand2_2 \uart_receiver/_380_  (.Y(\uart_receiver/_152_ ),
    .A(\uart_receiver/bit_counter[1] ),
    .B(\uart_receiver/bit_counter[0] ));
 sg13g2_nor2_1 \uart_receiver/_381_  (.A(\uart_receiver/_002_ ),
    .B(\uart_receiver/_152_ ),
    .Y(\uart_receiver/_153_ ));
 sg13g2_nor3_2 \uart_receiver/_382_  (.A(net4083),
    .B(net813),
    .C(\uart_receiver/_152_ ),
    .Y(\uart_receiver/_154_ ));
 sg13g2_a21oi_1 \uart_receiver/_383_  (.A1(\uart_receiver/stage[0] ),
    .A2(net3),
    .Y(\uart_receiver/_155_ ),
    .B1(net4481));
 sg13g2_o21ai_1 \uart_receiver/_384_  (.B1(\uart_receiver/_155_ ),
    .Y(\uart_receiver/_156_ ),
    .A1(net951),
    .A2(\uart_receiver/stage[2] ));
 sg13g2_a21oi_2 \uart_receiver/_385_  (.B1(\uart_receiver/_156_ ),
    .Y(\uart_receiver/_157_ ),
    .A2(\uart_receiver/_149_ ),
    .A1(\uart_receiver/stage[2] ));
 sg13g2_a21o_1 \uart_receiver/_386_  (.A2(\uart_receiver/_149_ ),
    .A1(\uart_receiver/stage[2] ),
    .B1(\uart_receiver/_156_ ),
    .X(\uart_receiver/_158_ ));
 sg13g2_nor2_1 \uart_receiver/_387_  (.A(\uart_receiver/_154_ ),
    .B(net3716),
    .Y(\uart_receiver/_159_ ));
 sg13g2_nand2b_1 \uart_receiver/_388_  (.Y(\uart_receiver/_160_ ),
    .B(\uart_receiver/_108_ ),
    .A_N(\uart_receiver/_152_ ));
 sg13g2_xnor2_1 \uart_receiver/_389_  (.Y(\uart_receiver/_161_ ),
    .A(net4084),
    .B(\uart_receiver/_152_ ));
 sg13g2_or4_1 \uart_receiver/_390_  (.A(net4083),
    .B(\uart_receiver/_154_ ),
    .C(net3716),
    .D(\uart_receiver/_161_ ),
    .X(\uart_receiver/_162_ ));
 sg13g2_o21ai_1 \uart_receiver/_391_  (.B1(\uart_receiver/_162_ ),
    .Y(\uart_receiver/_107_ ),
    .A1(net4084),
    .A2(\uart_receiver/_159_ ));
 sg13g2_a21oi_1 \uart_receiver/_392_  (.A1(\uart_receiver/bit_counter[0] ),
    .A2(\uart_receiver/_157_ ),
    .Y(\uart_receiver/_163_ ),
    .B1(\uart_receiver/bit_counter[1] ));
 sg13g2_nand2b_1 \uart_receiver/_393_  (.Y(\uart_receiver/_164_ ),
    .B(\uart_receiver/_152_ ),
    .A_N(net707));
 sg13g2_a21oi_1 \uart_receiver/_394_  (.A1(\uart_receiver/_159_ ),
    .A2(\uart_receiver/_164_ ),
    .Y(\uart_receiver/_106_ ),
    .B1(\uart_receiver/_163_ ));
 sg13g2_a21oi_1 \uart_receiver/_395_  (.A1(net183),
    .A2(\uart_receiver/_157_ ),
    .Y(\uart_receiver/_165_ ),
    .B1(net761));
 sg13g2_a21oi_1 \uart_receiver/_396_  (.A1(net761),
    .A2(\uart_receiver/_159_ ),
    .Y(\uart_receiver/_105_ ),
    .B1(\uart_receiver/_165_ ));
 sg13g2_nand3_1 \uart_receiver/_397_  (.B(\uart_receiver/bit_counter[1] ),
    .C(\uart_receiver/bit_counter[0] ),
    .A(\uart_receiver/bit_counter[2] ),
    .Y(\uart_receiver/_166_ ));
 sg13g2_or2_1 \uart_receiver/_398_  (.X(\uart_receiver/_167_ ),
    .B(\uart_receiver/_166_ ),
    .A(\uart_receiver/_158_ ));
 sg13g2_o21ai_1 \uart_receiver/_399_  (.B1(\uart_receiver/stage[2] ),
    .Y(\uart_receiver/_168_ ),
    .A1(net3),
    .A2(\uart_receiver/_166_ ));
 sg13g2_a22oi_1 \uart_receiver/_400_  (.Y(\uart_receiver/_104_ ),
    .B1(\uart_receiver/_168_ ),
    .B2(\uart_receiver/_157_ ),
    .A2(\uart_receiver/_167_ ),
    .A1(\uart_receiver/_109_ ));
 sg13g2_nor2b_1 \uart_receiver/_401_  (.A(net950),
    .B_N(\uart_receiver/bit_counter[1] ),
    .Y(\uart_receiver/_169_ ));
 sg13g2_nand2_1 \uart_receiver/_402_  (.Y(\uart_receiver/_170_ ),
    .A(\uart_receiver/bit_counter[2] ),
    .B(\uart_receiver/_169_ ));
 sg13g2_a21oi_1 \uart_receiver/_403_  (.A1(\uart_receiver/bit_counter[2] ),
    .A2(\uart_receiver/_169_ ),
    .Y(\uart_receiver/_171_ ),
    .B1(net4083));
 sg13g2_o21ai_1 \uart_receiver/_404_  (.B1(net85),
    .Y(\uart_receiver/_172_ ),
    .A1(net3716),
    .A2(\uart_receiver/_171_ ));
 sg13g2_nand2_2 \uart_receiver/_405_  (.Y(\uart_receiver/_173_ ),
    .A(net3),
    .B(\uart_receiver/_157_ ));
 sg13g2_o21ai_1 \uart_receiver/_406_  (.B1(\uart_receiver/_172_ ),
    .Y(\uart_receiver/_103_ ),
    .A1(\uart_receiver/_170_ ),
    .A2(\uart_receiver/_173_ ));
 sg13g2_nor2b_2 \uart_receiver/_407_  (.A(\uart_receiver/bit_counter[1] ),
    .B_N(\uart_receiver/bit_counter[0] ),
    .Y(\uart_receiver/_174_ ));
 sg13g2_nand2_1 \uart_receiver/_408_  (.Y(\uart_receiver/_175_ ),
    .A(\uart_receiver/bit_counter[2] ),
    .B(\uart_receiver/_174_ ));
 sg13g2_a21oi_1 \uart_receiver/_409_  (.A1(\uart_receiver/bit_counter[2] ),
    .A2(\uart_receiver/_174_ ),
    .Y(\uart_receiver/_176_ ),
    .B1(net4083));
 sg13g2_o21ai_1 \uart_receiver/_410_  (.B1(net98),
    .Y(\uart_receiver/_177_ ),
    .A1(net3716),
    .A2(\uart_receiver/_176_ ));
 sg13g2_o21ai_1 \uart_receiver/_411_  (.B1(\uart_receiver/_177_ ),
    .Y(\uart_receiver/_102_ ),
    .A1(\uart_receiver/_173_ ),
    .A2(\uart_receiver/_175_ ));
 sg13g2_nor2_1 \uart_receiver/_412_  (.A(\uart_receiver/bit_counter[1] ),
    .B(\uart_receiver/bit_counter[0] ),
    .Y(\uart_receiver/_178_ ));
 sg13g2_nand2_1 \uart_receiver/_413_  (.Y(\uart_receiver/_179_ ),
    .A(\uart_receiver/bit_counter[2] ),
    .B(\uart_receiver/_178_ ));
 sg13g2_a21oi_1 \uart_receiver/_414_  (.A1(\uart_receiver/bit_counter[2] ),
    .A2(\uart_receiver/_178_ ),
    .Y(\uart_receiver/_180_ ),
    .B1(net4083));
 sg13g2_o21ai_1 \uart_receiver/_415_  (.B1(net147),
    .Y(\uart_receiver/_181_ ),
    .A1(net3716),
    .A2(\uart_receiver/_180_ ));
 sg13g2_o21ai_1 \uart_receiver/_416_  (.B1(net148),
    .Y(\uart_receiver/_101_ ),
    .A1(\uart_receiver/_173_ ),
    .A2(\uart_receiver/_179_ ));
 sg13g2_nand2_1 \uart_receiver/_417_  (.Y(\uart_receiver/_182_ ),
    .A(\uart_receiver/stage[2] ),
    .B(\uart_receiver/_160_ ));
 sg13g2_inv_1 \uart_receiver/_418_  (.Y(\uart_receiver/_183_ ),
    .A(\uart_receiver/_182_ ));
 sg13g2_o21ai_1 \uart_receiver/_419_  (.B1(net102),
    .Y(\uart_receiver/_184_ ),
    .A1(\uart_receiver/_158_ ),
    .A2(\uart_receiver/_183_ ));
 sg13g2_o21ai_1 \uart_receiver/_420_  (.B1(\uart_receiver/_184_ ),
    .Y(\uart_receiver/_100_ ),
    .A1(\uart_receiver/_160_ ),
    .A2(\uart_receiver/_173_ ));
 sg13g2_nand2_1 \uart_receiver/_421_  (.Y(\uart_receiver/_185_ ),
    .A(net4084),
    .B(\uart_receiver/_169_ ));
 sg13g2_a21oi_1 \uart_receiver/_422_  (.A1(net4084),
    .A2(\uart_receiver/_169_ ),
    .Y(\uart_receiver/_186_ ),
    .B1(net4083));
 sg13g2_o21ai_1 \uart_receiver/_423_  (.B1(net150),
    .Y(\uart_receiver/_187_ ),
    .A1(net3716),
    .A2(\uart_receiver/_186_ ));
 sg13g2_o21ai_1 \uart_receiver/_424_  (.B1(\uart_receiver/_187_ ),
    .Y(\uart_receiver/_099_ ),
    .A1(\uart_receiver/_173_ ),
    .A2(\uart_receiver/_185_ ));
 sg13g2_nand2_1 \uart_receiver/_425_  (.Y(\uart_receiver/_188_ ),
    .A(net4084),
    .B(\uart_receiver/_174_ ));
 sg13g2_a21oi_1 \uart_receiver/_426_  (.A1(net4084),
    .A2(\uart_receiver/_174_ ),
    .Y(\uart_receiver/_189_ ),
    .B1(net4083));
 sg13g2_o21ai_1 \uart_receiver/_427_  (.B1(net82),
    .Y(\uart_receiver/_190_ ),
    .A1(net3716),
    .A2(\uart_receiver/_189_ ));
 sg13g2_o21ai_1 \uart_receiver/_428_  (.B1(\uart_receiver/_190_ ),
    .Y(\uart_receiver/_098_ ),
    .A1(\uart_receiver/_173_ ),
    .A2(\uart_receiver/_188_ ));
 sg13g2_nand2_1 \uart_receiver/_429_  (.Y(\uart_receiver/_191_ ),
    .A(net4084),
    .B(\uart_receiver/_178_ ));
 sg13g2_a21oi_1 \uart_receiver/_430_  (.A1(net4084),
    .A2(\uart_receiver/_178_ ),
    .Y(\uart_receiver/_192_ ),
    .B1(net4083));
 sg13g2_o21ai_1 \uart_receiver/_431_  (.B1(net176),
    .Y(\uart_receiver/_193_ ),
    .A1(net3716),
    .A2(\uart_receiver/_192_ ));
 sg13g2_o21ai_1 \uart_receiver/_432_  (.B1(\uart_receiver/_193_ ),
    .Y(\uart_receiver/_097_ ),
    .A1(\uart_receiver/_173_ ),
    .A2(\uart_receiver/_191_ ));
 sg13g2_nor2_1 \uart_receiver/_433_  (.A(\uart_receiver/stage[1] ),
    .B(\uart_receiver/stage[0] ),
    .Y(\uart_receiver/_194_ ));
 sg13g2_nand2_1 \uart_receiver/_434_  (.Y(\uart_receiver/_195_ ),
    .A(\uart_receiver/_004_ ),
    .B(\uart_receiver/_194_ ));
 sg13g2_nand2_2 \uart_receiver/_435_  (.Y(\uart_receiver/_196_ ),
    .A(\uart_receiver/_155_ ),
    .B(\uart_receiver/_195_ ));
 sg13g2_a21oi_2 \uart_receiver/_436_  (.B1(\uart_receiver/_196_ ),
    .Y(\uart_receiver/_197_ ),
    .A2(\uart_receiver/_148_ ),
    .A1(\uart_receiver/stage[1] ));
 sg13g2_a21o_1 \uart_receiver/_437_  (.A2(\uart_receiver/_148_ ),
    .A1(\uart_receiver/stage[1] ),
    .B1(\uart_receiver/_196_ ),
    .X(\uart_receiver/_198_ ));
 sg13g2_nand3_1 \uart_receiver/_438_  (.B(\uart_receiver/cycle_counter[1] ),
    .C(\uart_receiver/cycle_counter[0] ),
    .A(\uart_receiver/cycle_counter[2] ),
    .Y(\uart_receiver/_199_ ));
 sg13g2_nand4_1 \uart_receiver/_439_  (.B(\uart_receiver/cycle_counter[2] ),
    .C(\uart_receiver/cycle_counter[1] ),
    .A(\uart_receiver/cycle_counter[3] ),
    .Y(\uart_receiver/_200_ ),
    .D(\uart_receiver/cycle_counter[0] ));
 sg13g2_nor4_2 \uart_receiver/_440_  (.A(\uart_receiver/_116_ ),
    .B(\uart_receiver/_117_ ),
    .C(\uart_receiver/_118_ ),
    .Y(\uart_receiver/_201_ ),
    .D(\uart_receiver/_200_ ));
 sg13g2_nand2_1 \uart_receiver/_441_  (.Y(\uart_receiver/_202_ ),
    .A(\uart_receiver/cycle_counter[7] ),
    .B(\uart_receiver/_201_ ));
 sg13g2_and4_2 \uart_receiver/_442_  (.A(\uart_receiver/cycle_counter[9] ),
    .B(\uart_receiver/cycle_counter[8] ),
    .C(\uart_receiver/cycle_counter[7] ),
    .D(\uart_receiver/_201_ ),
    .X(\uart_receiver/_203_ ));
 sg13g2_nand3_1 \uart_receiver/_443_  (.B(\uart_receiver/cycle_counter[10] ),
    .C(\uart_receiver/_203_ ),
    .A(\uart_receiver/cycle_counter[11] ),
    .Y(\uart_receiver/_204_ ));
 sg13g2_a21oi_1 \uart_receiver/_444_  (.A1(\uart_receiver/_143_ ),
    .A2(\uart_receiver/_147_ ),
    .Y(\uart_receiver/_205_ ),
    .B1(\uart_receiver/_126_ ));
 sg13g2_nor2_1 \uart_receiver/_445_  (.A(\uart_receiver/stage[1] ),
    .B(\uart_receiver/stage[2] ),
    .Y(\uart_receiver/_206_ ));
 sg13g2_a21oi_2 \uart_receiver/_446_  (.B1(net4081),
    .Y(\uart_receiver/_207_ ),
    .A2(\uart_receiver/_147_ ),
    .A1(\uart_receiver/_143_ ));
 sg13g2_nand2_1 \uart_receiver/_447_  (.Y(\uart_receiver/_208_ ),
    .A(\uart_receiver/_204_ ),
    .B(net3768));
 sg13g2_a21oi_1 \uart_receiver/_448_  (.A1(\uart_receiver/_197_ ),
    .A2(\uart_receiver/_208_ ),
    .Y(\uart_receiver/_209_ ),
    .B1(\uart_receiver/_110_ ));
 sg13g2_or2_1 \uart_receiver/_449_  (.X(\uart_receiver/_210_ ),
    .B(\uart_receiver/cycles_per_bit[0] ),
    .A(\uart_receiver/cycles_per_bit[1] ));
 sg13g2_or4_2 \uart_receiver/_450_  (.A(\uart_receiver/cycles_per_bit[2] ),
    .B(\uart_receiver/cycles_per_bit[1] ),
    .C(\uart_receiver/cycles_per_bit[0] ),
    .D(\uart_receiver/cycles_per_bit[3] ),
    .X(\uart_receiver/_211_ ));
 sg13g2_nand2b_1 \uart_receiver/_451_  (.Y(\uart_receiver/_212_ ),
    .B(\uart_receiver/_124_ ),
    .A_N(\uart_receiver/_211_ ));
 sg13g2_nor2_1 \uart_receiver/_452_  (.A(\uart_receiver/cycles_per_bit[5] ),
    .B(\uart_receiver/_212_ ),
    .Y(\uart_receiver/_213_ ));
 sg13g2_nor3_1 \uart_receiver/_453_  (.A(\uart_receiver/cycles_per_bit[7] ),
    .B(\uart_receiver/cycles_per_bit[5] ),
    .C(\uart_receiver/cycles_per_bit[6] ),
    .Y(\uart_receiver/_214_ ));
 sg13g2_nand3b_1 \uart_receiver/_454_  (.B(\uart_receiver/_214_ ),
    .C(\uart_receiver/_124_ ),
    .Y(\uart_receiver/_215_ ),
    .A_N(\uart_receiver/_211_ ));
 sg13g2_nor4_1 \uart_receiver/_455_  (.A(\uart_receiver/cycles_per_bit[10] ),
    .B(\uart_receiver/cycles_per_bit[9] ),
    .C(\uart_receiver/cycles_per_bit[8] ),
    .D(\uart_receiver/cycles_per_bit[11] ),
    .Y(\uart_receiver/_216_ ));
 sg13g2_nand2b_1 \uart_receiver/_456_  (.Y(\uart_receiver/_217_ ),
    .B(\uart_receiver/_216_ ),
    .A_N(\uart_receiver/_215_ ));
 sg13g2_o21ai_1 \uart_receiver/_457_  (.B1(net4081),
    .Y(\uart_receiver/_218_ ),
    .A1(\uart_receiver/cycles_per_bit[12] ),
    .A2(\uart_receiver/_217_ ));
 sg13g2_a21oi_1 \uart_receiver/_458_  (.A1(\uart_receiver/cycles_per_bit[12] ),
    .A2(\uart_receiver/_217_ ),
    .Y(\uart_receiver/_219_ ),
    .B1(\uart_receiver/_218_ ));
 sg13g2_nor2_1 \uart_receiver/_459_  (.A(\uart_receiver/cycle_counter[12] ),
    .B(\uart_receiver/_204_ ),
    .Y(\uart_receiver/_220_ ));
 sg13g2_a21o_1 \uart_receiver/_460_  (.A2(\uart_receiver/_220_ ),
    .A1(net3768),
    .B1(\uart_receiver/_219_ ),
    .X(\uart_receiver/_221_ ));
 sg13g2_a21o_1 \uart_receiver/_461_  (.A2(\uart_receiver/_221_ ),
    .A1(\uart_receiver/_197_ ),
    .B1(\uart_receiver/_209_ ),
    .X(\uart_receiver/_096_ ));
 sg13g2_a21oi_1 \uart_receiver/_462_  (.A1(\uart_receiver/cycle_counter[10] ),
    .A2(\uart_receiver/_203_ ),
    .Y(\uart_receiver/_222_ ),
    .B1(net806));
 sg13g2_a21o_1 \uart_receiver/_463_  (.A2(\uart_receiver/_208_ ),
    .A1(\uart_receiver/_197_ ),
    .B1(\uart_receiver/_222_ ),
    .X(\uart_receiver/_223_ ));
 sg13g2_nor3_1 \uart_receiver/_464_  (.A(\uart_receiver/cycles_per_bit[9] ),
    .B(\uart_receiver/cycles_per_bit[8] ),
    .C(\uart_receiver/_215_ ),
    .Y(\uart_receiver/_224_ ));
 sg13g2_nand2_1 \uart_receiver/_465_  (.Y(\uart_receiver/_225_ ),
    .A(net765),
    .B(\uart_receiver/_224_ ));
 sg13g2_xor2_1 \uart_receiver/_466_  (.B(\uart_receiver/_225_ ),
    .A(\uart_receiver/cycles_per_bit[11] ),
    .X(\uart_receiver/_226_ ));
 sg13g2_nand2b_1 \uart_receiver/_467_  (.Y(\uart_receiver/_227_ ),
    .B(\uart_receiver/_226_ ),
    .A_N(\uart_receiver/_218_ ));
 sg13g2_a22oi_1 \uart_receiver/_468_  (.Y(\uart_receiver/_095_ ),
    .B1(\uart_receiver/_223_ ),
    .B2(\uart_receiver/_227_ ),
    .A2(net3715),
    .A1(\uart_receiver/_111_ ));
 sg13g2_or2_1 \uart_receiver/_469_  (.X(\uart_receiver/_228_ ),
    .B(\uart_receiver/_203_ ),
    .A(\uart_receiver/cycle_counter[10] ));
 sg13g2_a221oi_1 \uart_receiver/_470_  (.B2(\uart_receiver/cycle_counter[10] ),
    .C1(net4081),
    .B1(\uart_receiver/_203_ ),
    .A1(\uart_receiver/_143_ ),
    .Y(\uart_receiver/_229_ ),
    .A2(\uart_receiver/_147_ ));
 sg13g2_o21ai_1 \uart_receiver/_471_  (.B1(\uart_receiver/_228_ ),
    .Y(\uart_receiver/_230_ ),
    .A1(net3715),
    .A2(\uart_receiver/_229_ ));
 sg13g2_or2_1 \uart_receiver/_472_  (.X(\uart_receiver/_231_ ),
    .B(\uart_receiver/_224_ ),
    .A(net765));
 sg13g2_nand3b_1 \uart_receiver/_473_  (.B(\uart_receiver/_225_ ),
    .C(\uart_receiver/_231_ ),
    .Y(\uart_receiver/_232_ ),
    .A_N(\uart_receiver/_218_ ));
 sg13g2_a22oi_1 \uart_receiver/_474_  (.Y(\uart_receiver/_094_ ),
    .B1(\uart_receiver/_230_ ),
    .B2(\uart_receiver/_232_ ),
    .A2(net3715),
    .A1(\uart_receiver/_112_ ));
 sg13g2_o21ai_1 \uart_receiver/_475_  (.B1(\uart_receiver/_113_ ),
    .Y(\uart_receiver/_233_ ),
    .A1(\uart_receiver/_114_ ),
    .A2(\uart_receiver/_202_ ));
 sg13g2_nor2b_1 \uart_receiver/_476_  (.A(\uart_receiver/_203_ ),
    .B_N(net3768),
    .Y(\uart_receiver/_234_ ));
 sg13g2_o21ai_1 \uart_receiver/_477_  (.B1(\uart_receiver/_233_ ),
    .Y(\uart_receiver/_235_ ),
    .A1(net3715),
    .A2(\uart_receiver/_234_ ));
 sg13g2_o21ai_1 \uart_receiver/_478_  (.B1(net495),
    .Y(\uart_receiver/_236_ ),
    .A1(\uart_receiver/cycles_per_bit[8] ),
    .A2(\uart_receiver/_215_ ));
 sg13g2_nand3b_1 \uart_receiver/_479_  (.B(\uart_receiver/_236_ ),
    .C(net4081),
    .Y(\uart_receiver/_237_ ),
    .A_N(\uart_receiver/_224_ ));
 sg13g2_a22oi_1 \uart_receiver/_480_  (.Y(\uart_receiver/_093_ ),
    .B1(\uart_receiver/_235_ ),
    .B2(\uart_receiver/_237_ ),
    .A2(net3715),
    .A1(\uart_receiver/_113_ ));
 sg13g2_xor2_1 \uart_receiver/_481_  (.B(\uart_receiver/_215_ ),
    .A(\uart_receiver/cycles_per_bit[8] ),
    .X(\uart_receiver/_238_ ));
 sg13g2_xnor2_1 \uart_receiver/_482_  (.Y(\uart_receiver/_239_ ),
    .A(net781),
    .B(\uart_receiver/_202_ ));
 sg13g2_a221oi_1 \uart_receiver/_483_  (.B2(net3768),
    .C1(net3715),
    .B1(\uart_receiver/_239_ ),
    .A1(net4081),
    .Y(\uart_receiver/_240_ ),
    .A2(\uart_receiver/_238_ ));
 sg13g2_a21oi_1 \uart_receiver/_484_  (.A1(\uart_receiver/_114_ ),
    .A2(net3715),
    .Y(\uart_receiver/_092_ ),
    .B1(\uart_receiver/_240_ ));
 sg13g2_nand2_1 \uart_receiver/_485_  (.Y(\uart_receiver/_241_ ),
    .A(\uart_receiver/_202_ ),
    .B(net3768));
 sg13g2_nor2_1 \uart_receiver/_486_  (.A(net698),
    .B(\uart_receiver/_201_ ),
    .Y(\uart_receiver/_242_ ));
 sg13g2_a21o_1 \uart_receiver/_487_  (.A2(\uart_receiver/_241_ ),
    .A1(\uart_receiver/_197_ ),
    .B1(\uart_receiver/_242_ ),
    .X(\uart_receiver/_243_ ));
 sg13g2_nand2b_1 \uart_receiver/_488_  (.Y(\uart_receiver/_244_ ),
    .B(\uart_receiver/_213_ ),
    .A_N(\uart_receiver/cycles_per_bit[6] ));
 sg13g2_nand2_1 \uart_receiver/_489_  (.Y(\uart_receiver/_245_ ),
    .A(net640),
    .B(\uart_receiver/_244_ ));
 sg13g2_nand3_1 \uart_receiver/_490_  (.B(\uart_receiver/_215_ ),
    .C(\uart_receiver/_245_ ),
    .A(net4081),
    .Y(\uart_receiver/_246_ ));
 sg13g2_a22oi_1 \uart_receiver/_491_  (.Y(\uart_receiver/_091_ ),
    .B1(\uart_receiver/_243_ ),
    .B2(\uart_receiver/_246_ ),
    .A2(net3715),
    .A1(\uart_receiver/_115_ ));
 sg13g2_xnor2_1 \uart_receiver/_492_  (.Y(\uart_receiver/_247_ ),
    .A(\uart_receiver/cycles_per_bit[6] ),
    .B(\uart_receiver/_213_ ));
 sg13g2_nor2_1 \uart_receiver/_493_  (.A(\uart_receiver/_118_ ),
    .B(\uart_receiver/_200_ ),
    .Y(\uart_receiver/_248_ ));
 sg13g2_a21oi_1 \uart_receiver/_494_  (.A1(\uart_receiver/cycle_counter[5] ),
    .A2(\uart_receiver/_248_ ),
    .Y(\uart_receiver/_249_ ),
    .B1(net795));
 sg13g2_nor2_1 \uart_receiver/_495_  (.A(\uart_receiver/_201_ ),
    .B(\uart_receiver/_249_ ),
    .Y(\uart_receiver/_250_ ));
 sg13g2_a221oi_1 \uart_receiver/_496_  (.B2(net3768),
    .C1(net3713),
    .B1(\uart_receiver/_250_ ),
    .A1(net4082),
    .Y(\uart_receiver/_251_ ),
    .A2(\uart_receiver/_247_ ));
 sg13g2_a21oi_1 \uart_receiver/_497_  (.A1(\uart_receiver/_116_ ),
    .A2(net3713),
    .Y(\uart_receiver/_090_ ),
    .B1(\uart_receiver/_251_ ));
 sg13g2_a221oi_1 \uart_receiver/_498_  (.B2(\uart_receiver/cycle_counter[5] ),
    .C1(net4081),
    .B1(\uart_receiver/_248_ ),
    .A1(\uart_receiver/_143_ ),
    .Y(\uart_receiver/_252_ ),
    .A2(\uart_receiver/_147_ ));
 sg13g2_o21ai_1 \uart_receiver/_499_  (.B1(\uart_receiver/_117_ ),
    .Y(\uart_receiver/_253_ ),
    .A1(\uart_receiver/_118_ ),
    .A2(\uart_receiver/_200_ ));
 sg13g2_o21ai_1 \uart_receiver/_500_  (.B1(\uart_receiver/_253_ ),
    .Y(\uart_receiver/_254_ ),
    .A1(net3713),
    .A2(\uart_receiver/_252_ ));
 sg13g2_nand2_1 \uart_receiver/_501_  (.Y(\uart_receiver/_255_ ),
    .A(net840),
    .B(\uart_receiver/_212_ ));
 sg13g2_nand3b_1 \uart_receiver/_502_  (.B(\uart_receiver/_255_ ),
    .C(net4081),
    .Y(\uart_receiver/_256_ ),
    .A_N(\uart_receiver/_213_ ));
 sg13g2_a22oi_1 \uart_receiver/_503_  (.Y(\uart_receiver/_089_ ),
    .B1(\uart_receiver/_254_ ),
    .B2(\uart_receiver/_256_ ),
    .A2(net3713),
    .A1(\uart_receiver/_117_ ));
 sg13g2_nand2_1 \uart_receiver/_504_  (.Y(\uart_receiver/_257_ ),
    .A(net858),
    .B(\uart_receiver/_211_ ));
 sg13g2_nand3_1 \uart_receiver/_505_  (.B(\uart_receiver/_212_ ),
    .C(net859),
    .A(net4082),
    .Y(\uart_receiver/_258_ ));
 sg13g2_xnor2_1 \uart_receiver/_506_  (.Y(\uart_receiver/_259_ ),
    .A(\uart_receiver/cycle_counter[4] ),
    .B(\uart_receiver/_200_ ));
 sg13g2_a21oi_1 \uart_receiver/_507_  (.A1(\uart_receiver/_207_ ),
    .A2(\uart_receiver/_259_ ),
    .Y(\uart_receiver/_260_ ),
    .B1(net3713));
 sg13g2_a22oi_1 \uart_receiver/_508_  (.Y(\uart_receiver/_088_ ),
    .B1(\uart_receiver/_258_ ),
    .B2(\uart_receiver/_260_ ),
    .A2(net3713),
    .A1(\uart_receiver/_118_ ));
 sg13g2_and2_1 \uart_receiver/_509_  (.A(\uart_receiver/_200_ ),
    .B(\uart_receiver/_207_ ),
    .X(\uart_receiver/_261_ ));
 sg13g2_nand2_1 \uart_receiver/_510_  (.Y(\uart_receiver/_262_ ),
    .A(\uart_receiver/_119_ ),
    .B(\uart_receiver/_199_ ));
 sg13g2_o21ai_1 \uart_receiver/_511_  (.B1(\uart_receiver/_262_ ),
    .Y(\uart_receiver/_263_ ),
    .A1(net3714),
    .A2(\uart_receiver/_261_ ));
 sg13g2_o21ai_1 \uart_receiver/_512_  (.B1(\uart_receiver/cycles_per_bit[3] ),
    .Y(\uart_receiver/_264_ ),
    .A1(\uart_receiver/cycles_per_bit[2] ),
    .A2(\uart_receiver/_210_ ));
 sg13g2_nand3_1 \uart_receiver/_513_  (.B(\uart_receiver/_211_ ),
    .C(\uart_receiver/_264_ ),
    .A(net4082),
    .Y(\uart_receiver/_265_ ));
 sg13g2_a22oi_1 \uart_receiver/_514_  (.Y(\uart_receiver/_087_ ),
    .B1(\uart_receiver/_263_ ),
    .B2(\uart_receiver/_265_ ),
    .A2(net3714),
    .A1(\uart_receiver/_119_ ));
 sg13g2_o21ai_1 \uart_receiver/_515_  (.B1(net4082),
    .Y(\uart_receiver/_266_ ),
    .A1(net812),
    .A2(\uart_receiver/_210_ ));
 sg13g2_a21o_1 \uart_receiver/_516_  (.A2(\uart_receiver/_210_ ),
    .A1(net812),
    .B1(\uart_receiver/_266_ ),
    .X(\uart_receiver/_267_ ));
 sg13g2_o21ai_1 \uart_receiver/_517_  (.B1(\uart_receiver/_120_ ),
    .Y(\uart_receiver/_268_ ),
    .A1(\uart_receiver/_121_ ),
    .A2(\uart_receiver/_122_ ));
 sg13g2_and2_1 \uart_receiver/_518_  (.A(\uart_receiver/_199_ ),
    .B(\uart_receiver/_268_ ),
    .X(\uart_receiver/_269_ ));
 sg13g2_a21oi_1 \uart_receiver/_519_  (.A1(net3768),
    .A2(\uart_receiver/_269_ ),
    .Y(\uart_receiver/_270_ ),
    .B1(net3714));
 sg13g2_a22oi_1 \uart_receiver/_520_  (.Y(\uart_receiver/_086_ ),
    .B1(\uart_receiver/_267_ ),
    .B2(\uart_receiver/_270_ ),
    .A2(net3714),
    .A1(\uart_receiver/_120_ ));
 sg13g2_xor2_1 \uart_receiver/_521_  (.B(\uart_receiver/cycle_counter[0] ),
    .A(\uart_receiver/cycle_counter[1] ),
    .X(\uart_receiver/_271_ ));
 sg13g2_nand2_1 \uart_receiver/_522_  (.Y(\uart_receiver/_272_ ),
    .A(net645),
    .B(\uart_receiver/cycles_per_bit[0] ));
 sg13g2_nand3_1 \uart_receiver/_523_  (.B(\uart_receiver/_210_ ),
    .C(\uart_receiver/_272_ ),
    .A(net4082),
    .Y(\uart_receiver/_273_ ));
 sg13g2_a21oi_1 \uart_receiver/_524_  (.A1(net3768),
    .A2(\uart_receiver/_271_ ),
    .Y(\uart_receiver/_274_ ),
    .B1(net3713));
 sg13g2_a22oi_1 \uart_receiver/_525_  (.Y(\uart_receiver/_085_ ),
    .B1(\uart_receiver/_273_ ),
    .B2(\uart_receiver/_274_ ),
    .A2(net3714),
    .A1(\uart_receiver/_121_ ));
 sg13g2_a221oi_1 \uart_receiver/_526_  (.B2(\uart_receiver/_122_ ),
    .C1(net3713),
    .B1(\uart_receiver/_207_ ),
    .A1(\uart_receiver/cycles_per_bit[0] ),
    .Y(\uart_receiver/_275_ ),
    .A2(net4082));
 sg13g2_a21oi_1 \uart_receiver/_527_  (.A1(\uart_receiver/_122_ ),
    .A2(net3714),
    .Y(\uart_receiver/_084_ ),
    .B1(\uart_receiver/_275_ ));
 sg13g2_nor2_1 \uart_receiver/_528_  (.A(\uart_receiver/_010_ ),
    .B(net4478),
    .Y(\uart_receiver/_276_ ));
 sg13g2_a21oi_1 \uart_receiver/_529_  (.A1(net4478),
    .A2(net41),
    .Y(\uart_receiver/_083_ ),
    .B1(\uart_receiver/_276_ ));
 sg13g2_nor2_1 \uart_receiver/_530_  (.A(net4478),
    .B(net59),
    .Y(\uart_receiver/_277_ ));
 sg13g2_a21oi_1 \uart_receiver/_531_  (.A1(net4478),
    .A2(\cpu.rx_speed[11] ),
    .Y(\uart_receiver/_082_ ),
    .B1(\uart_receiver/_277_ ));
 sg13g2_mux2_1 \uart_receiver/_532_  (.A0(net569),
    .A1(net409),
    .S(net4478),
    .X(\uart_receiver/_081_ ));
 sg13g2_mux2_1 \uart_receiver/_533_  (.A0(net495),
    .A1(net248),
    .S(net4478),
    .X(\uart_receiver/_080_ ));
 sg13g2_mux2_1 \uart_receiver/_534_  (.A0(net650),
    .A1(net270),
    .S(net4478),
    .X(\uart_receiver/_079_ ));
 sg13g2_mux2_1 \uart_receiver/_535_  (.A0(net640),
    .A1(\cpu.rx_speed[7] ),
    .S(net4480),
    .X(\uart_receiver/_078_ ));
 sg13g2_nor2_1 \uart_receiver/_536_  (.A(net4478),
    .B(net62),
    .Y(\uart_receiver/_278_ ));
 sg13g2_a21oi_1 \uart_receiver/_537_  (.A1(net4480),
    .A2(\cpu.rx_speed[6] ),
    .Y(\uart_receiver/_077_ ),
    .B1(\uart_receiver/_278_ ));
 sg13g2_nor2_1 \uart_receiver/_538_  (.A(net4479),
    .B(net48),
    .Y(\uart_receiver/_279_ ));
 sg13g2_a21oi_1 \uart_receiver/_539_  (.A1(net4479),
    .A2(\cpu.rx_speed[5] ),
    .Y(\uart_receiver/_076_ ),
    .B1(\uart_receiver/_279_ ));
 sg13g2_nand2_1 \uart_receiver/_540_  (.Y(\uart_receiver/_280_ ),
    .A(net4479),
    .B(net578));
 sg13g2_o21ai_1 \uart_receiver/_541_  (.B1(\uart_receiver/_280_ ),
    .Y(\uart_receiver/_075_ ),
    .A1(net4479),
    .A2(\uart_receiver/_124_ ));
 sg13g2_nor2_1 \uart_receiver/_542_  (.A(net4480),
    .B(net43),
    .Y(\uart_receiver/_281_ ));
 sg13g2_a21oi_1 \uart_receiver/_543_  (.A1(net4479),
    .A2(\cpu.rx_speed[3] ),
    .Y(\uart_receiver/_074_ ),
    .B1(\uart_receiver/_281_ ));
 sg13g2_mux2_1 \uart_receiver/_544_  (.A0(net812),
    .A1(net633),
    .S(net4480),
    .X(\uart_receiver/_073_ ));
 sg13g2_mux2_1 \uart_receiver/_545_  (.A0(net645),
    .A1(net311),
    .S(net4479),
    .X(\uart_receiver/_072_ ));
 sg13g2_nor2_1 \uart_receiver/_546_  (.A(net4479),
    .B(net57),
    .Y(\uart_receiver/_282_ ));
 sg13g2_a21oi_1 \uart_receiver/_547_  (.A1(net4479),
    .A2(\cpu.rx_speed[0] ),
    .Y(\uart_receiver/_071_ ),
    .B1(\uart_receiver/_282_ ));
 sg13g2_nor3_1 \uart_receiver/_548_  (.A(net4481),
    .B(\uart_receiver/_194_ ),
    .C(\uart_receiver/_205_ ),
    .Y(\uart_receiver/_283_ ));
 sg13g2_nor2b_1 \uart_receiver/_549_  (.A(net3712),
    .B_N(\data_received[7] ),
    .Y(\uart_receiver/_284_ ));
 sg13g2_a21o_1 \uart_receiver/_550_  (.A2(\uart_receiver/_150_ ),
    .A1(net154),
    .B1(\uart_receiver/_284_ ),
    .X(\uart_receiver/_070_ ));
 sg13g2_nor2b_1 \uart_receiver/_551_  (.A(net3712),
    .B_N(net151),
    .Y(\uart_receiver/_285_ ));
 sg13g2_a21o_1 \uart_receiver/_552_  (.A2(net3717),
    .A1(net85),
    .B1(\uart_receiver/_285_ ),
    .X(\uart_receiver/_069_ ));
 sg13g2_nor2b_1 \uart_receiver/_553_  (.A(net3712),
    .B_N(net206),
    .Y(\uart_receiver/_286_ ));
 sg13g2_a21o_1 \uart_receiver/_554_  (.A2(net3717),
    .A1(net98),
    .B1(\uart_receiver/_286_ ),
    .X(\uart_receiver/_068_ ));
 sg13g2_nor2b_1 \uart_receiver/_555_  (.A(net3712),
    .B_N(net374),
    .Y(\uart_receiver/_287_ ));
 sg13g2_a21o_1 \uart_receiver/_556_  (.A2(net3717),
    .A1(net147),
    .B1(\uart_receiver/_287_ ),
    .X(\uart_receiver/_067_ ));
 sg13g2_nor2b_1 \uart_receiver/_557_  (.A(net3712),
    .B_N(net190),
    .Y(\uart_receiver/_288_ ));
 sg13g2_a21o_1 \uart_receiver/_558_  (.A2(net3717),
    .A1(net102),
    .B1(\uart_receiver/_288_ ),
    .X(\uart_receiver/_066_ ));
 sg13g2_nor2b_1 \uart_receiver/_559_  (.A(net3712),
    .B_N(net197),
    .Y(\uart_receiver/_289_ ));
 sg13g2_a21o_1 \uart_receiver/_560_  (.A2(net3717),
    .A1(net150),
    .B1(\uart_receiver/_289_ ),
    .X(\uart_receiver/_065_ ));
 sg13g2_nor2b_1 \uart_receiver/_561_  (.A(net3712),
    .B_N(net139),
    .Y(\uart_receiver/_290_ ));
 sg13g2_a21o_1 \uart_receiver/_562_  (.A2(net3717),
    .A1(net82),
    .B1(\uart_receiver/_290_ ),
    .X(\uart_receiver/_064_ ));
 sg13g2_nor2b_1 \uart_receiver/_563_  (.A(net3712),
    .B_N(net339),
    .Y(\uart_receiver/_291_ ));
 sg13g2_a21o_1 \uart_receiver/_564_  (.A2(net3717),
    .A1(net176),
    .B1(\uart_receiver/_291_ ),
    .X(\uart_receiver/_063_ ));
 sg13g2_nand2b_1 \uart_receiver/_565_  (.Y(\uart_receiver/_292_ ),
    .B(net182),
    .A_N(\uart_receiver/_283_ ));
 sg13g2_nand2b_1 \uart_receiver/_566_  (.Y(\uart_receiver/_062_ ),
    .B(\uart_receiver/_292_ ),
    .A_N(\uart_receiver/_150_ ));
 sg13g2_a21o_1 \uart_receiver/_567_  (.A2(\uart_receiver/_153_ ),
    .A1(\uart_receiver/_151_ ),
    .B1(\uart_receiver/_127_ ),
    .X(\uart_receiver/_293_ ));
 sg13g2_nand2b_1 \uart_receiver/_568_  (.Y(\uart_receiver/_294_ ),
    .B(net521),
    .A_N(net4481));
 sg13g2_o21ai_1 \uart_receiver/_569_  (.B1(\uart_receiver/_293_ ),
    .Y(\uart_receiver/_001_ ),
    .A1(net3),
    .A2(\uart_receiver/_294_ ));
 sg13g2_mux2_1 \uart_receiver/_570_  (.A0(\uart_receiver/stage[1] ),
    .A1(\uart_receiver/_154_ ),
    .S(\uart_receiver/_151_ ),
    .X(\uart_receiver/_000_ ));
 sg13g2_inv_1 \uart_receiver/_571_  (.Y(\uart_receiver/_013_ ),
    .A(net4577));
 sg13g2_inv_1 \uart_receiver/_572_  (.Y(\uart_receiver/_014_ ),
    .A(net4577));
 sg13g2_inv_1 \uart_receiver/_573_  (.Y(\uart_receiver/_015_ ),
    .A(net4577));
 sg13g2_inv_1 \uart_receiver/_574_  (.Y(\uart_receiver/_016_ ),
    .A(net4578));
 sg13g2_inv_1 \uart_receiver/_575_  (.Y(\uart_receiver/_017_ ),
    .A(net4579));
 sg13g2_inv_1 \uart_receiver/_576_  (.Y(\uart_receiver/_018_ ),
    .A(net4577));
 sg13g2_inv_1 \uart_receiver/_577_  (.Y(\uart_receiver/_019_ ),
    .A(net4577));
 sg13g2_inv_1 \uart_receiver/_578_  (.Y(\uart_receiver/_020_ ),
    .A(net4581));
 sg13g2_inv_1 \uart_receiver/_579_  (.Y(\uart_receiver/_021_ ),
    .A(net4582));
 sg13g2_inv_1 \uart_receiver/_580_  (.Y(\uart_receiver/_022_ ),
    .A(net4582));
 sg13g2_inv_1 \uart_receiver/_581_  (.Y(\uart_receiver/_023_ ),
    .A(net4582));
 sg13g2_inv_1 \uart_receiver/_582_  (.Y(\uart_receiver/_024_ ),
    .A(net4582));
 sg13g2_inv_1 \uart_receiver/_583_  (.Y(\uart_receiver/_025_ ),
    .A(net4582));
 sg13g2_inv_1 \uart_receiver/_584_  (.Y(\uart_receiver/_026_ ),
    .A(net4582));
 sg13g2_inv_1 \uart_receiver/_585_  (.Y(\uart_receiver/_027_ ),
    .A(net4584));
 sg13g2_inv_1 \uart_receiver/_586_  (.Y(\uart_receiver/_028_ ),
    .A(net4584));
 sg13g2_inv_1 \uart_receiver/_587_  (.Y(\uart_receiver/_029_ ),
    .A(net4585));
 sg13g2_inv_1 \uart_receiver/_588_  (.Y(\uart_receiver/_030_ ),
    .A(net4585));
 sg13g2_inv_1 \uart_receiver/_589_  (.Y(\uart_receiver/_031_ ),
    .A(net4584));
 sg13g2_inv_1 \uart_receiver/_590_  (.Y(\uart_receiver/_032_ ),
    .A(net4585));
 sg13g2_inv_1 \uart_receiver/_591_  (.Y(\uart_receiver/_033_ ),
    .A(net4585));
 sg13g2_inv_1 \uart_receiver/_592_  (.Y(\uart_receiver/_034_ ),
    .A(net4583));
 sg13g2_inv_1 \uart_receiver/_593_  (.Y(\uart_receiver/_035_ ),
    .A(net4583));
 sg13g2_inv_1 \uart_receiver/_594_  (.Y(\uart_receiver/_036_ ),
    .A(net4582));
 sg13g2_inv_1 \uart_receiver/_595_  (.Y(\uart_receiver/_037_ ),
    .A(net4582));
 sg13g2_inv_1 \uart_receiver/_596_  (.Y(\uart_receiver/_038_ ),
    .A(net4583));
 sg13g2_inv_1 \uart_receiver/_597_  (.Y(\uart_receiver/_039_ ),
    .A(net4583));
 sg13g2_inv_1 \uart_receiver/_598_  (.Y(\uart_receiver/_040_ ),
    .A(net4584));
 sg13g2_inv_1 \uart_receiver/_599_  (.Y(\uart_receiver/_041_ ),
    .A(net4584));
 sg13g2_inv_1 \uart_receiver/_600_  (.Y(\uart_receiver/_042_ ),
    .A(net4585));
 sg13g2_inv_1 \uart_receiver/_601_  (.Y(\uart_receiver/_043_ ),
    .A(net4585));
 sg13g2_inv_1 \uart_receiver/_602_  (.Y(\uart_receiver/_044_ ),
    .A(net4584));
 sg13g2_inv_1 \uart_receiver/_603_  (.Y(\uart_receiver/_045_ ),
    .A(net4584));
 sg13g2_inv_1 \uart_receiver/_604_  (.Y(\uart_receiver/_046_ ),
    .A(net4585));
 sg13g2_inv_1 \uart_receiver/_605_  (.Y(\uart_receiver/_047_ ),
    .A(net4578));
 sg13g2_inv_1 \uart_receiver/_606_  (.Y(\uart_receiver/_048_ ),
    .A(net4577));
 sg13g2_inv_1 \uart_receiver/_607_  (.Y(\uart_receiver/_049_ ),
    .A(net4578));
 sg13g2_inv_1 \uart_receiver/_608_  (.Y(\uart_receiver/_050_ ),
    .A(net4578));
 sg13g2_inv_1 \uart_receiver/_609_  (.Y(\uart_receiver/_051_ ),
    .A(net4578));
 sg13g2_inv_1 \uart_receiver/_610_  (.Y(\uart_receiver/_052_ ),
    .A(net4577));
 sg13g2_inv_1 \uart_receiver/_611_  (.Y(\uart_receiver/_053_ ),
    .A(net4577));
 sg13g2_inv_1 \uart_receiver/_612_  (.Y(\uart_receiver/_054_ ),
    .A(net4581));
 sg13g2_inv_1 \uart_receiver/_613_  (.Y(\uart_receiver/_055_ ),
    .A(net4578));
 sg13g2_inv_1 \uart_receiver/_614_  (.Y(\uart_receiver/_056_ ),
    .A(net4578));
 sg13g2_inv_1 \uart_receiver/_615_  (.Y(\uart_receiver/_057_ ),
    .A(net4578));
 sg13g2_inv_1 \uart_receiver/_616_  (.Y(\uart_receiver/_059_ ),
    .A(net4581));
 sg13g2_inv_1 \uart_receiver/_617_  (.Y(\uart_receiver/_060_ ),
    .A(net4581));
 sg13g2_inv_1 \uart_receiver/_618_  (.Y(\uart_receiver/_061_ ),
    .A(net4581));
 sg13g2_dfrbp_1 \uart_receiver/_619_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(\uart_receiver/_012_ ),
    .D(\uart_receiver/_062_ ),
    .Q_N(\uart_receiver/_333_ ),
    .Q(\cpu.uart_inbound ));
 sg13g2_dfrbp_1 \uart_receiver/_620_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(\uart_receiver/_013_ ),
    .D(\uart_receiver/_063_ ),
    .Q_N(\uart_receiver/_332_ ),
    .Q(\data_received[0] ));
 sg13g2_dfrbp_1 \uart_receiver/_621_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(\uart_receiver/_014_ ),
    .D(\uart_receiver/_064_ ),
    .Q_N(\uart_receiver/_331_ ),
    .Q(\data_received[1] ));
 sg13g2_dfrbp_1 \uart_receiver/_622_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(\uart_receiver/_015_ ),
    .D(\uart_receiver/_065_ ),
    .Q_N(\uart_receiver/_330_ ),
    .Q(\data_received[2] ));
 sg13g2_dfrbp_1 \uart_receiver/_623_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(\uart_receiver/_016_ ),
    .D(\uart_receiver/_066_ ),
    .Q_N(\uart_receiver/_329_ ),
    .Q(\data_received[3] ));
 sg13g2_dfrbp_1 \uart_receiver/_624_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(\uart_receiver/_017_ ),
    .D(\uart_receiver/_067_ ),
    .Q_N(\uart_receiver/_328_ ),
    .Q(\data_received[4] ));
 sg13g2_dfrbp_1 \uart_receiver/_625_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(\uart_receiver/_018_ ),
    .D(\uart_receiver/_068_ ),
    .Q_N(\uart_receiver/_327_ ),
    .Q(\data_received[5] ));
 sg13g2_dfrbp_1 \uart_receiver/_626_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(\uart_receiver/_019_ ),
    .D(\uart_receiver/_069_ ),
    .Q_N(\uart_receiver/_326_ ),
    .Q(\data_received[6] ));
 sg13g2_dfrbp_1 \uart_receiver/_627_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(\uart_receiver/_020_ ),
    .D(net155),
    .Q_N(\uart_receiver/_325_ ),
    .Q(\data_received[7] ));
 sg13g2_dfrbp_1 \uart_receiver/_628_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(\uart_receiver/_021_ ),
    .D(net58),
    .Q_N(\uart_receiver/cycles_per_bit[0] ),
    .Q(\uart_receiver/_005_ ));
 sg13g2_dfrbp_1 \uart_receiver/_629_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(\uart_receiver/_022_ ),
    .D(\uart_receiver/_072_ ),
    .Q_N(\uart_receiver/_324_ ),
    .Q(\uart_receiver/cycles_per_bit[1] ));
 sg13g2_dfrbp_1 \uart_receiver/_630_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(\uart_receiver/_023_ ),
    .D(\uart_receiver/_073_ ),
    .Q_N(\uart_receiver/_323_ ),
    .Q(\uart_receiver/cycles_per_bit[2] ));
 sg13g2_dfrbp_1 \uart_receiver/_631_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(\uart_receiver/_024_ ),
    .D(net44),
    .Q_N(\uart_receiver/cycles_per_bit[3] ),
    .Q(\uart_receiver/_006_ ));
 sg13g2_dfrbp_1 \uart_receiver/_632_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(\uart_receiver/_025_ ),
    .D(net579),
    .Q_N(\uart_receiver/_322_ ),
    .Q(\uart_receiver/cycles_per_bit[4] ));
 sg13g2_dfrbp_1 \uart_receiver/_633_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(\uart_receiver/_026_ ),
    .D(net49),
    .Q_N(\uart_receiver/cycles_per_bit[5] ),
    .Q(\uart_receiver/_007_ ));
 sg13g2_dfrbp_1 \uart_receiver/_634_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(\uart_receiver/_027_ ),
    .D(net63),
    .Q_N(\uart_receiver/cycles_per_bit[6] ),
    .Q(\uart_receiver/_008_ ));
 sg13g2_dfrbp_1 \uart_receiver/_635_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(\uart_receiver/_028_ ),
    .D(net641),
    .Q_N(\uart_receiver/_321_ ),
    .Q(\uart_receiver/cycles_per_bit[7] ));
 sg13g2_dfrbp_1 \uart_receiver/_636_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(\uart_receiver/_029_ ),
    .D(\uart_receiver/_079_ ),
    .Q_N(\uart_receiver/_320_ ),
    .Q(\uart_receiver/cycles_per_bit[8] ));
 sg13g2_dfrbp_1 \uart_receiver/_637_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(\uart_receiver/_030_ ),
    .D(\uart_receiver/_080_ ),
    .Q_N(\uart_receiver/_319_ ),
    .Q(\uart_receiver/cycles_per_bit[9] ));
 sg13g2_dfrbp_1 \uart_receiver/_638_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(\uart_receiver/_031_ ),
    .D(\uart_receiver/_081_ ),
    .Q_N(\uart_receiver/_003_ ),
    .Q(\uart_receiver/cycles_per_bit[10] ));
 sg13g2_dfrbp_1 \uart_receiver/_639_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(\uart_receiver/_032_ ),
    .D(net60),
    .Q_N(\uart_receiver/cycles_per_bit[11] ),
    .Q(\uart_receiver/_009_ ));
 sg13g2_dfrbp_1 \uart_receiver/_640_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(\uart_receiver/_033_ ),
    .D(net42),
    .Q_N(\uart_receiver/cycles_per_bit[12] ),
    .Q(\uart_receiver/_010_ ));
 sg13g2_dfrbp_1 \uart_receiver/_641_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(\uart_receiver/_034_ ),
    .D(net827),
    .Q_N(\uart_receiver/_318_ ),
    .Q(\uart_receiver/cycle_counter[0] ));
 sg13g2_dfrbp_1 \uart_receiver/_642_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(\uart_receiver/_035_ ),
    .D(net836),
    .Q_N(\uart_receiver/_317_ ),
    .Q(\uart_receiver/cycle_counter[1] ));
 sg13g2_dfrbp_1 \uart_receiver/_643_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(\uart_receiver/_036_ ),
    .D(\uart_receiver/_086_ ),
    .Q_N(\uart_receiver/_316_ ),
    .Q(\uart_receiver/cycle_counter[2] ));
 sg13g2_dfrbp_1 \uart_receiver/_644_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(\uart_receiver/_037_ ),
    .D(net702),
    .Q_N(\uart_receiver/_315_ ),
    .Q(\uart_receiver/cycle_counter[3] ));
 sg13g2_dfrbp_1 \uart_receiver/_645_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(\uart_receiver/_038_ ),
    .D(net860),
    .Q_N(\uart_receiver/_314_ ),
    .Q(\uart_receiver/cycle_counter[4] ));
 sg13g2_dfrbp_1 \uart_receiver/_646_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(\uart_receiver/_039_ ),
    .D(net841),
    .Q_N(\uart_receiver/_313_ ),
    .Q(\uart_receiver/cycle_counter[5] ));
 sg13g2_dfrbp_1 \uart_receiver/_647_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(\uart_receiver/_040_ ),
    .D(net796),
    .Q_N(\uart_receiver/_312_ ),
    .Q(\uart_receiver/cycle_counter[6] ));
 sg13g2_dfrbp_1 \uart_receiver/_648_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(\uart_receiver/_041_ ),
    .D(\uart_receiver/_091_ ),
    .Q_N(\uart_receiver/_311_ ),
    .Q(\uart_receiver/cycle_counter[7] ));
 sg13g2_dfrbp_1 \uart_receiver/_649_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(\uart_receiver/_042_ ),
    .D(\uart_receiver/_092_ ),
    .Q_N(\uart_receiver/_310_ ),
    .Q(\uart_receiver/cycle_counter[8] ));
 sg13g2_dfrbp_1 \uart_receiver/_650_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(\uart_receiver/_043_ ),
    .D(net710),
    .Q_N(\uart_receiver/_309_ ),
    .Q(\uart_receiver/cycle_counter[9] ));
 sg13g2_dfrbp_1 \uart_receiver/_651_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(\uart_receiver/_044_ ),
    .D(net766),
    .Q_N(\uart_receiver/_308_ ),
    .Q(\uart_receiver/cycle_counter[10] ));
 sg13g2_dfrbp_1 \uart_receiver/_652_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(\uart_receiver/_045_ ),
    .D(net807),
    .Q_N(\uart_receiver/_307_ ),
    .Q(\uart_receiver/cycle_counter[11] ));
 sg13g2_dfrbp_1 \uart_receiver/_653_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(\uart_receiver/_046_ ),
    .D(\uart_receiver/_096_ ),
    .Q_N(\uart_receiver/_306_ ),
    .Q(\uart_receiver/cycle_counter[12] ));
 sg13g2_dfrbp_1 \uart_receiver/_654_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(\uart_receiver/_047_ ),
    .D(net177),
    .Q_N(\uart_receiver/_305_ ),
    .Q(\uart_receiver/data[0] ));
 sg13g2_dfrbp_1 \uart_receiver/_655_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(\uart_receiver/_048_ ),
    .D(net83),
    .Q_N(\uart_receiver/_304_ ),
    .Q(\uart_receiver/data[1] ));
 sg13g2_dfrbp_1 \uart_receiver/_656_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(\uart_receiver/_049_ ),
    .D(\uart_receiver/_099_ ),
    .Q_N(\uart_receiver/_303_ ),
    .Q(\uart_receiver/data[2] ));
 sg13g2_dfrbp_1 \uart_receiver/_657_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(\uart_receiver/_050_ ),
    .D(net103),
    .Q_N(\uart_receiver/_302_ ),
    .Q(\uart_receiver/data[3] ));
 sg13g2_dfrbp_1 \uart_receiver/_658_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(\uart_receiver/_051_ ),
    .D(net149),
    .Q_N(\uart_receiver/_301_ ),
    .Q(\uart_receiver/data[4] ));
 sg13g2_dfrbp_1 \uart_receiver/_659_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(\uart_receiver/_052_ ),
    .D(net99),
    .Q_N(\uart_receiver/_300_ ),
    .Q(\uart_receiver/data[5] ));
 sg13g2_dfrbp_1 \uart_receiver/_660_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(\uart_receiver/_053_ ),
    .D(net86),
    .Q_N(\uart_receiver/_299_ ),
    .Q(\uart_receiver/data[6] ));
 sg13g2_dfrbp_1 \uart_receiver/_661_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(\uart_receiver/_054_ ),
    .D(\uart_receiver/_104_ ),
    .Q_N(\uart_receiver/_298_ ),
    .Q(\uart_receiver/data[7] ));
 sg13g2_dfrbp_1 \uart_receiver/_662_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(\uart_receiver/_055_ ),
    .D(net762),
    .Q_N(\uart_receiver/_297_ ),
    .Q(\uart_receiver/bit_counter[0] ));
 sg13g2_dfrbp_1 \uart_receiver/_663_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(\uart_receiver/_056_ ),
    .D(net708),
    .Q_N(\uart_receiver/_296_ ),
    .Q(\uart_receiver/bit_counter[1] ));
 sg13g2_dfrbp_1 \uart_receiver/_664_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(\uart_receiver/_057_ ),
    .D(\uart_receiver/_107_ ),
    .Q_N(\uart_receiver/_002_ ),
    .Q(\uart_receiver/bit_counter[2] ));
 sg13g2_dfrbp_1 \uart_receiver/_665_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(\uart_receiver/_059_ ),
    .D(\uart_receiver/_058_ ),
    .Q_N(\uart_receiver/stage[0] ),
    .Q(\uart_receiver/_011_ ));
 sg13g2_dfrbp_1 \uart_receiver/_666_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(\uart_receiver/_060_ ),
    .D(net814),
    .Q_N(\uart_receiver/_295_ ),
    .Q(\uart_receiver/stage[1] ));
 sg13g2_dfrbp_1 \uart_receiver/_667_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(\uart_receiver/_061_ ),
    .D(net522),
    .Q_N(\uart_receiver/_004_ ),
    .Q(\uart_receiver/stage[2] ));
 sg13g2_buf_2 fanout3538 (.A(net3539),
    .X(net3538));
 sg13g2_buf_2 fanout3539 (.A(net3540),
    .X(net3539));
 sg13g2_buf_4 fanout3540 (.X(net3540),
    .A(_06334_));
 sg13g2_buf_2 fanout3541 (.A(net3542),
    .X(net3541));
 sg13g2_buf_1 fanout3542 (.A(_04132_),
    .X(net3542));
 sg13g2_buf_4 fanout3543 (.X(net3543),
    .A(net3544));
 sg13g2_buf_2 fanout3544 (.A(net3547),
    .X(net3544));
 sg13g2_buf_2 fanout3545 (.A(net3546),
    .X(net3545));
 sg13g2_buf_4 fanout3546 (.X(net3546),
    .A(net3547));
 sg13g2_buf_2 fanout3547 (.A(_06455_),
    .X(net3547));
 sg13g2_buf_2 fanout3548 (.A(net3551),
    .X(net3548));
 sg13g2_buf_2 fanout3549 (.A(net3551),
    .X(net3549));
 sg13g2_buf_1 fanout3550 (.A(net3551),
    .X(net3550));
 sg13g2_buf_2 fanout3551 (.A(_04130_),
    .X(net3551));
 sg13g2_buf_4 fanout3552 (.X(net3552),
    .A(net3553));
 sg13g2_buf_4 fanout3553 (.X(net3553),
    .A(net3555));
 sg13g2_buf_2 fanout3554 (.A(net3555),
    .X(net3554));
 sg13g2_buf_4 fanout3555 (.X(net3555),
    .A(_04130_));
 sg13g2_buf_2 fanout3556 (.A(net3557),
    .X(net3556));
 sg13g2_buf_1 fanout3557 (.A(net3558),
    .X(net3557));
 sg13g2_buf_2 fanout3558 (.A(_04129_),
    .X(net3558));
 sg13g2_buf_2 fanout3559 (.A(net3562),
    .X(net3559));
 sg13g2_buf_2 fanout3560 (.A(net3562),
    .X(net3560));
 sg13g2_buf_1 fanout3561 (.A(net3562),
    .X(net3561));
 sg13g2_buf_2 fanout3562 (.A(_04125_),
    .X(net3562));
 sg13g2_buf_4 fanout3563 (.X(net3563),
    .A(net3564));
 sg13g2_buf_4 fanout3564 (.X(net3564),
    .A(net3566));
 sg13g2_buf_2 fanout3565 (.A(net3566),
    .X(net3565));
 sg13g2_buf_2 fanout3566 (.A(_04125_),
    .X(net3566));
 sg13g2_buf_2 fanout3567 (.A(net3568),
    .X(net3567));
 sg13g2_buf_1 fanout3568 (.A(net3569),
    .X(net3568));
 sg13g2_buf_2 fanout3569 (.A(_04124_),
    .X(net3569));
 sg13g2_buf_2 fanout3570 (.A(net3572),
    .X(net3570));
 sg13g2_buf_2 fanout3571 (.A(net3572),
    .X(net3571));
 sg13g2_buf_2 fanout3572 (.A(net3573),
    .X(net3572));
 sg13g2_buf_4 fanout3573 (.X(net3573),
    .A(_04106_));
 sg13g2_buf_2 fanout3574 (.A(net3576),
    .X(net3574));
 sg13g2_buf_1 fanout3575 (.A(net3576),
    .X(net3575));
 sg13g2_buf_1 fanout3576 (.A(_04105_),
    .X(net3576));
 sg13g2_buf_2 fanout3577 (.A(net3578),
    .X(net3577));
 sg13g2_buf_2 fanout3578 (.A(_04105_),
    .X(net3578));
 sg13g2_buf_2 fanout3579 (.A(net3581),
    .X(net3579));
 sg13g2_buf_2 fanout3580 (.A(net3581),
    .X(net3580));
 sg13g2_buf_2 fanout3581 (.A(net3582),
    .X(net3581));
 sg13g2_buf_4 fanout3582 (.X(net3582),
    .A(_04065_));
 sg13g2_buf_2 fanout3583 (.A(net3585),
    .X(net3583));
 sg13g2_buf_1 fanout3584 (.A(net3585),
    .X(net3584));
 sg13g2_buf_1 fanout3585 (.A(_04064_),
    .X(net3585));
 sg13g2_buf_2 fanout3586 (.A(net3587),
    .X(net3586));
 sg13g2_buf_2 fanout3587 (.A(_04064_),
    .X(net3587));
 sg13g2_buf_2 fanout3588 (.A(net3590),
    .X(net3588));
 sg13g2_buf_1 fanout3589 (.A(net3590),
    .X(net3589));
 sg13g2_buf_1 fanout3590 (.A(_04058_),
    .X(net3590));
 sg13g2_buf_2 fanout3591 (.A(net3592),
    .X(net3591));
 sg13g2_buf_2 fanout3592 (.A(_04058_),
    .X(net3592));
 sg13g2_buf_2 fanout3593 (.A(net3594),
    .X(net3593));
 sg13g2_buf_2 fanout3594 (.A(_03783_),
    .X(net3594));
 sg13g2_buf_2 fanout3595 (.A(net3596),
    .X(net3595));
 sg13g2_buf_2 fanout3596 (.A(net3597),
    .X(net3596));
 sg13g2_buf_2 fanout3597 (.A(_03783_),
    .X(net3597));
 sg13g2_buf_2 fanout3598 (.A(net3599),
    .X(net3598));
 sg13g2_buf_2 fanout3599 (.A(_03700_),
    .X(net3599));
 sg13g2_buf_2 fanout3600 (.A(net3601),
    .X(net3600));
 sg13g2_buf_4 fanout3601 (.X(net3601),
    .A(_03700_));
 sg13g2_buf_2 fanout3602 (.A(net3603),
    .X(net3602));
 sg13g2_buf_4 fanout3603 (.X(net3603),
    .A(net3604));
 sg13g2_buf_4 fanout3604 (.X(net3604),
    .A(_02590_));
 sg13g2_buf_2 fanout3605 (.A(net3606),
    .X(net3605));
 sg13g2_buf_4 fanout3606 (.X(net3606),
    .A(_02590_));
 sg13g2_buf_2 fanout3607 (.A(net3609),
    .X(net3607));
 sg13g2_buf_1 fanout3608 (.A(net3609),
    .X(net3608));
 sg13g2_buf_4 fanout3609 (.X(net3609),
    .A(_02440_));
 sg13g2_buf_2 fanout3610 (.A(net3611),
    .X(net3610));
 sg13g2_buf_2 fanout3611 (.A(_02440_),
    .X(net3611));
 sg13g2_buf_2 fanout3612 (.A(net3613),
    .X(net3612));
 sg13g2_buf_2 fanout3613 (.A(net3614),
    .X(net3613));
 sg13g2_buf_1 fanout3614 (.A(_02018_),
    .X(net3614));
 sg13g2_buf_2 fanout3615 (.A(net3616),
    .X(net3615));
 sg13g2_buf_4 fanout3616 (.X(net3616),
    .A(_02018_));
 sg13g2_buf_2 fanout3617 (.A(net3618),
    .X(net3617));
 sg13g2_buf_2 fanout3618 (.A(net3621),
    .X(net3618));
 sg13g2_buf_2 fanout3619 (.A(net3620),
    .X(net3619));
 sg13g2_buf_2 fanout3620 (.A(net3621),
    .X(net3620));
 sg13g2_buf_2 fanout3621 (.A(_01930_),
    .X(net3621));
 sg13g2_buf_2 fanout3622 (.A(net3624),
    .X(net3622));
 sg13g2_buf_1 fanout3623 (.A(net3624),
    .X(net3623));
 sg13g2_buf_2 fanout3624 (.A(_01440_),
    .X(net3624));
 sg13g2_buf_4 fanout3625 (.X(net3625),
    .A(net3626));
 sg13g2_buf_4 fanout3626 (.X(net3626),
    .A(_01440_));
 sg13g2_buf_2 fanout3627 (.A(_06544_),
    .X(net3627));
 sg13g2_buf_1 fanout3628 (.A(_06544_),
    .X(net3628));
 sg13g2_buf_2 fanout3629 (.A(net3630),
    .X(net3629));
 sg13g2_buf_4 fanout3630 (.X(net3630),
    .A(net3631));
 sg13g2_buf_4 fanout3631 (.X(net3631),
    .A(_05895_));
 sg13g2_buf_4 fanout3632 (.X(net3632),
    .A(_05895_));
 sg13g2_buf_2 fanout3633 (.A(_05895_),
    .X(net3633));
 sg13g2_buf_4 fanout3634 (.X(net3634),
    .A(net3635));
 sg13g2_buf_4 fanout3635 (.X(net3635),
    .A(_05505_));
 sg13g2_buf_4 fanout3636 (.X(net3636),
    .A(_04059_));
 sg13g2_buf_2 fanout3637 (.A(net3639),
    .X(net3637));
 sg13g2_buf_2 fanout3638 (.A(net3639),
    .X(net3638));
 sg13g2_buf_4 fanout3639 (.X(net3639),
    .A(_04059_));
 sg13g2_buf_2 fanout3640 (.A(net3641),
    .X(net3640));
 sg13g2_buf_2 fanout3641 (.A(_03272_),
    .X(net3641));
 sg13g2_buf_2 fanout3642 (.A(net3644),
    .X(net3642));
 sg13g2_buf_1 fanout3643 (.A(net3644),
    .X(net3643));
 sg13g2_buf_2 fanout3644 (.A(_03272_),
    .X(net3644));
 sg13g2_buf_2 fanout3645 (.A(net3646),
    .X(net3645));
 sg13g2_buf_4 fanout3646 (.X(net3646),
    .A(_02573_));
 sg13g2_buf_4 fanout3647 (.X(net3647),
    .A(_02573_));
 sg13g2_buf_2 fanout3648 (.A(_02573_),
    .X(net3648));
 sg13g2_buf_4 fanout3649 (.X(net3649),
    .A(net3650));
 sg13g2_buf_4 fanout3650 (.X(net3650),
    .A(_02555_));
 sg13g2_buf_4 fanout3651 (.X(net3651),
    .A(_02555_));
 sg13g2_buf_2 fanout3652 (.A(_02555_),
    .X(net3652));
 sg13g2_buf_4 fanout3653 (.X(net3653),
    .A(net3655));
 sg13g2_buf_2 fanout3654 (.A(net3655),
    .X(net3654));
 sg13g2_buf_4 fanout3655 (.X(net3655),
    .A(_02538_));
 sg13g2_buf_4 fanout3656 (.X(net3656),
    .A(_02538_));
 sg13g2_buf_2 fanout3657 (.A(_02538_),
    .X(net3657));
 sg13g2_buf_2 fanout3658 (.A(net3660),
    .X(net3658));
 sg13g2_buf_1 fanout3659 (.A(net3660),
    .X(net3659));
 sg13g2_buf_8 fanout3660 (.A(net3661),
    .X(net3660));
 sg13g2_buf_8 fanout3661 (.A(_02521_),
    .X(net3661));
 sg13g2_buf_4 fanout3662 (.X(net3662),
    .A(_02504_));
 sg13g2_buf_2 fanout3663 (.A(_02504_),
    .X(net3663));
 sg13g2_buf_2 fanout3664 (.A(net3666),
    .X(net3664));
 sg13g2_buf_1 fanout3665 (.A(net3666),
    .X(net3665));
 sg13g2_buf_2 fanout3666 (.A(net3667),
    .X(net3666));
 sg13g2_buf_2 fanout3667 (.A(net3668),
    .X(net3667));
 sg13g2_buf_4 fanout3668 (.X(net3668),
    .A(_02458_));
 sg13g2_buf_2 fanout3669 (.A(net3670),
    .X(net3669));
 sg13g2_buf_4 fanout3670 (.X(net3670),
    .A(net3673));
 sg13g2_buf_2 fanout3671 (.A(net3672),
    .X(net3671));
 sg13g2_buf_2 fanout3672 (.A(net3673),
    .X(net3672));
 sg13g2_buf_2 fanout3673 (.A(_02419_),
    .X(net3673));
 sg13g2_buf_2 fanout3674 (.A(net3676),
    .X(net3674));
 sg13g2_buf_2 fanout3675 (.A(net3676),
    .X(net3675));
 sg13g2_buf_4 fanout3676 (.X(net3676),
    .A(_02401_));
 sg13g2_buf_4 fanout3677 (.X(net3677),
    .A(_02401_));
 sg13g2_buf_2 fanout3678 (.A(_02401_),
    .X(net3678));
 sg13g2_buf_4 fanout3679 (.X(net3679),
    .A(net3680));
 sg13g2_buf_4 fanout3680 (.X(net3680),
    .A(net3683));
 sg13g2_buf_4 fanout3681 (.X(net3681),
    .A(net3682));
 sg13g2_buf_4 fanout3682 (.X(net3682),
    .A(net3683));
 sg13g2_buf_4 fanout3683 (.X(net3683),
    .A(_02384_));
 sg13g2_buf_2 fanout3684 (.A(net3686),
    .X(net3684));
 sg13g2_buf_1 fanout3685 (.A(net3686),
    .X(net3685));
 sg13g2_buf_4 fanout3686 (.X(net3686),
    .A(_02362_));
 sg13g2_buf_2 fanout3687 (.A(_02362_),
    .X(net3687));
 sg13g2_buf_1 fanout3688 (.A(_02362_),
    .X(net3688));
 sg13g2_buf_4 fanout3689 (.X(net3689),
    .A(net3691));
 sg13g2_buf_4 fanout3690 (.X(net3690),
    .A(net3691));
 sg13g2_buf_2 fanout3691 (.A(_02329_),
    .X(net3691));
 sg13g2_buf_4 fanout3692 (.X(net3692),
    .A(net3694));
 sg13g2_buf_4 fanout3693 (.X(net3693),
    .A(net3694));
 sg13g2_buf_2 fanout3694 (.A(_02292_),
    .X(net3694));
 sg13g2_buf_4 fanout3695 (.X(net3695),
    .A(net3696));
 sg13g2_buf_4 fanout3696 (.X(net3696),
    .A(_05085_));
 sg13g2_buf_4 fanout3697 (.X(net3697),
    .A(net3698));
 sg13g2_buf_8 fanout3698 (.A(_04325_),
    .X(net3698));
 sg13g2_buf_4 fanout3699 (.X(net3699),
    .A(net3700));
 sg13g2_buf_4 fanout3700 (.X(net3700),
    .A(_02486_));
 sg13g2_buf_4 fanout3701 (.X(net3701),
    .A(net3705));
 sg13g2_buf_2 fanout3702 (.A(net3705),
    .X(net3702));
 sg13g2_buf_2 fanout3703 (.A(net3705),
    .X(net3703));
 sg13g2_buf_4 fanout3704 (.X(net3704),
    .A(net3705));
 sg13g2_buf_2 fanout3705 (.A(net3706),
    .X(net3705));
 sg13g2_buf_4 fanout3706 (.X(net3706),
    .A(_02484_));
 sg13g2_buf_4 fanout3707 (.X(net3707),
    .A(net3709));
 sg13g2_buf_4 fanout3708 (.X(net3708),
    .A(net3709));
 sg13g2_buf_4 fanout3709 (.X(net3709),
    .A(_02291_));
 sg13g2_buf_4 fanout3710 (.X(net3710),
    .A(net3711));
 sg13g2_buf_4 fanout3711 (.X(net3711),
    .A(_02290_));
 sg13g2_buf_4 fanout3712 (.X(net3712),
    .A(\uart_receiver/_283_ ));
 sg13g2_buf_2 fanout3713 (.A(\uart_receiver/_198_ ),
    .X(net3713));
 sg13g2_buf_1 fanout3714 (.A(\uart_receiver/_198_ ),
    .X(net3714));
 sg13g2_buf_2 fanout3715 (.A(\uart_receiver/_198_ ),
    .X(net3715));
 sg13g2_buf_2 fanout3716 (.A(\uart_receiver/_158_ ),
    .X(net3716));
 sg13g2_buf_4 fanout3717 (.X(net3717),
    .A(\uart_receiver/_150_ ));
 sg13g2_buf_4 fanout3718 (.X(net3718),
    .A(_05083_));
 sg13g2_buf_2 fanout3719 (.A(net3721),
    .X(net3719));
 sg13g2_buf_1 fanout3720 (.A(net3721),
    .X(net3720));
 sg13g2_buf_2 fanout3721 (.A(net3722),
    .X(net3721));
 sg13g2_buf_4 fanout3722 (.X(net3722),
    .A(net3725));
 sg13g2_buf_2 fanout3723 (.A(net3724),
    .X(net3723));
 sg13g2_buf_4 fanout3724 (.X(net3724),
    .A(net3725));
 sg13g2_buf_2 fanout3725 (.A(_03863_),
    .X(net3725));
 sg13g2_buf_4 fanout3726 (.X(net3726),
    .A(net3729));
 sg13g2_buf_4 fanout3727 (.X(net3727),
    .A(net3729));
 sg13g2_buf_2 fanout3728 (.A(net3729),
    .X(net3728));
 sg13g2_buf_2 fanout3729 (.A(_03863_),
    .X(net3729));
 sg13g2_buf_2 fanout3730 (.A(net3731),
    .X(net3730));
 sg13g2_buf_1 fanout3731 (.A(net3737),
    .X(net3731));
 sg13g2_buf_2 fanout3732 (.A(net3737),
    .X(net3732));
 sg13g2_buf_2 fanout3733 (.A(net3735),
    .X(net3733));
 sg13g2_buf_2 fanout3734 (.A(net3735),
    .X(net3734));
 sg13g2_buf_2 fanout3735 (.A(net3736),
    .X(net3735));
 sg13g2_buf_2 fanout3736 (.A(net3737),
    .X(net3736));
 sg13g2_buf_2 fanout3737 (.A(_03863_),
    .X(net3737));
 sg13g2_buf_4 fanout3738 (.X(net3738),
    .A(_03862_));
 sg13g2_buf_4 fanout3739 (.X(net3739),
    .A(_03862_));
 sg13g2_buf_2 fanout3740 (.A(net3741),
    .X(net3740));
 sg13g2_buf_4 fanout3741 (.X(net3741),
    .A(_02879_));
 sg13g2_buf_2 fanout3742 (.A(net3743),
    .X(net3742));
 sg13g2_buf_4 fanout3743 (.X(net3743),
    .A(_02876_));
 sg13g2_buf_4 fanout3744 (.X(net3744),
    .A(_02744_));
 sg13g2_buf_4 fanout3745 (.X(net3745),
    .A(_02744_));
 sg13g2_buf_2 fanout3746 (.A(_02743_),
    .X(net3746));
 sg13g2_buf_4 fanout3747 (.X(net3747),
    .A(_02743_));
 sg13g2_buf_2 fanout3748 (.A(net3749),
    .X(net3748));
 sg13g2_buf_4 fanout3749 (.X(net3749),
    .A(_02628_));
 sg13g2_buf_2 fanout3750 (.A(net3753),
    .X(net3750));
 sg13g2_buf_2 fanout3751 (.A(net3752),
    .X(net3751));
 sg13g2_buf_4 fanout3752 (.X(net3752),
    .A(net3753));
 sg13g2_buf_2 fanout3753 (.A(_02624_),
    .X(net3753));
 sg13g2_buf_4 fanout3754 (.X(net3754),
    .A(_02482_));
 sg13g2_buf_4 fanout3755 (.X(net3755),
    .A(_02457_));
 sg13g2_buf_2 fanout3756 (.A(net3757),
    .X(net3756));
 sg13g2_buf_2 fanout3757 (.A(net3758),
    .X(net3757));
 sg13g2_buf_2 fanout3758 (.A(net3759),
    .X(net3758));
 sg13g2_buf_4 fanout3759 (.X(net3759),
    .A(net3760));
 sg13g2_buf_4 fanout3760 (.X(net3760),
    .A(_02327_));
 sg13g2_buf_4 fanout3761 (.X(net3761),
    .A(net3762));
 sg13g2_buf_4 fanout3762 (.X(net3762),
    .A(_02288_));
 sg13g2_buf_2 fanout3763 (.A(net3765),
    .X(net3763));
 sg13g2_buf_2 fanout3764 (.A(net3765),
    .X(net3764));
 sg13g2_buf_4 fanout3765 (.X(net3765),
    .A(_02261_));
 sg13g2_buf_4 fanout3766 (.X(net3766),
    .A(_02261_));
 sg13g2_buf_2 fanout3767 (.A(_02261_),
    .X(net3767));
 sg13g2_buf_2 fanout3768 (.A(\uart_receiver/_207_ ),
    .X(net3768));
 sg13g2_buf_2 fanout3769 (.A(_06262_),
    .X(net3769));
 sg13g2_buf_4 fanout3770 (.X(net3770),
    .A(net3771));
 sg13g2_buf_4 fanout3771 (.X(net3771),
    .A(_05081_));
 sg13g2_buf_2 fanout3772 (.A(net3773),
    .X(net3772));
 sg13g2_buf_2 fanout3773 (.A(net3775),
    .X(net3773));
 sg13g2_buf_4 fanout3774 (.X(net3774),
    .A(net3775));
 sg13g2_buf_2 fanout3775 (.A(net3779),
    .X(net3775));
 sg13g2_buf_2 fanout3776 (.A(net3779),
    .X(net3776));
 sg13g2_buf_2 fanout3777 (.A(net3778),
    .X(net3777));
 sg13g2_buf_2 fanout3778 (.A(net3779),
    .X(net3778));
 sg13g2_buf_2 fanout3779 (.A(_04258_),
    .X(net3779));
 sg13g2_buf_2 fanout3780 (.A(_03930_),
    .X(net3780));
 sg13g2_buf_2 fanout3781 (.A(net3782),
    .X(net3781));
 sg13g2_buf_4 fanout3782 (.X(net3782),
    .A(net3784));
 sg13g2_buf_4 fanout3783 (.X(net3783),
    .A(net3784));
 sg13g2_buf_2 fanout3784 (.A(_03882_),
    .X(net3784));
 sg13g2_buf_2 fanout3785 (.A(net3787),
    .X(net3785));
 sg13g2_buf_4 fanout3786 (.X(net3786),
    .A(net3787));
 sg13g2_buf_2 fanout3787 (.A(_03882_),
    .X(net3787));
 sg13g2_buf_4 fanout3788 (.X(net3788),
    .A(net3790));
 sg13g2_buf_2 fanout3789 (.A(net3790),
    .X(net3789));
 sg13g2_buf_4 fanout3790 (.X(net3790),
    .A(net3794));
 sg13g2_buf_2 fanout3791 (.A(net3792),
    .X(net3791));
 sg13g2_buf_4 fanout3792 (.X(net3792),
    .A(net3794));
 sg13g2_buf_4 fanout3793 (.X(net3793),
    .A(net3794));
 sg13g2_buf_2 fanout3794 (.A(_03881_),
    .X(net3794));
 sg13g2_buf_4 fanout3795 (.X(net3795),
    .A(_03293_));
 sg13g2_buf_2 fanout3796 (.A(net3797),
    .X(net3796));
 sg13g2_buf_4 fanout3797 (.X(net3797),
    .A(net3800));
 sg13g2_buf_4 fanout3798 (.X(net3798),
    .A(net3799));
 sg13g2_buf_4 fanout3799 (.X(net3799),
    .A(net3800));
 sg13g2_buf_2 fanout3800 (.A(_02623_),
    .X(net3800));
 sg13g2_buf_2 fanout3801 (.A(net3804),
    .X(net3801));
 sg13g2_buf_1 fanout3802 (.A(net3804),
    .X(net3802));
 sg13g2_buf_4 fanout3803 (.X(net3803),
    .A(net3804));
 sg13g2_buf_2 fanout3804 (.A(_02622_),
    .X(net3804));
 sg13g2_buf_4 fanout3805 (.X(net3805),
    .A(_01291_));
 sg13g2_buf_2 fanout3806 (.A(_01291_),
    .X(net3806));
 sg13g2_buf_2 fanout3807 (.A(_06395_),
    .X(net3807));
 sg13g2_buf_4 fanout3808 (.X(net3808),
    .A(_06275_));
 sg13g2_buf_2 fanout3809 (.A(_06273_),
    .X(net3809));
 sg13g2_buf_2 fanout3810 (.A(_06267_),
    .X(net3810));
 sg13g2_buf_4 fanout3811 (.X(net3811),
    .A(net3812));
 sg13g2_buf_4 fanout3812 (.X(net3812),
    .A(_04324_));
 sg13g2_buf_4 fanout3813 (.X(net3813),
    .A(net3814));
 sg13g2_buf_4 fanout3814 (.X(net3814),
    .A(_04324_));
 sg13g2_buf_2 fanout3815 (.A(net3816),
    .X(net3815));
 sg13g2_buf_2 fanout3816 (.A(net3817),
    .X(net3816));
 sg13g2_buf_2 fanout3817 (.A(net3818),
    .X(net3817));
 sg13g2_buf_4 fanout3818 (.X(net3818),
    .A(net3820));
 sg13g2_buf_4 fanout3819 (.X(net3819),
    .A(net3820));
 sg13g2_buf_4 fanout3820 (.X(net3820),
    .A(_04323_));
 sg13g2_buf_2 fanout3821 (.A(net3826),
    .X(net3821));
 sg13g2_buf_1 fanout3822 (.A(net3826),
    .X(net3822));
 sg13g2_buf_2 fanout3823 (.A(net3825),
    .X(net3823));
 sg13g2_buf_1 fanout3824 (.A(net3825),
    .X(net3824));
 sg13g2_buf_2 fanout3825 (.A(net3826),
    .X(net3825));
 sg13g2_buf_4 fanout3826 (.X(net3826),
    .A(_04302_));
 sg13g2_buf_2 fanout3827 (.A(_04301_),
    .X(net3827));
 sg13g2_buf_2 fanout3828 (.A(net3830),
    .X(net3828));
 sg13g2_buf_1 fanout3829 (.A(net3830),
    .X(net3829));
 sg13g2_buf_2 fanout3830 (.A(net3831),
    .X(net3830));
 sg13g2_buf_2 fanout3831 (.A(net3832),
    .X(net3831));
 sg13g2_buf_2 fanout3832 (.A(_04301_),
    .X(net3832));
 sg13g2_buf_2 fanout3833 (.A(_04259_),
    .X(net3833));
 sg13g2_buf_4 fanout3834 (.X(net3834),
    .A(_04259_));
 sg13g2_buf_2 fanout3835 (.A(_03939_),
    .X(net3835));
 sg13g2_buf_2 fanout3836 (.A(net3837),
    .X(net3836));
 sg13g2_buf_1 fanout3837 (.A(net3838),
    .X(net3837));
 sg13g2_buf_4 fanout3838 (.X(net3838),
    .A(_03875_));
 sg13g2_buf_2 fanout3839 (.A(net3840),
    .X(net3839));
 sg13g2_buf_2 fanout3840 (.A(_03875_),
    .X(net3840));
 sg13g2_buf_4 fanout3841 (.X(net3841),
    .A(net3845));
 sg13g2_buf_2 fanout3842 (.A(net3845),
    .X(net3842));
 sg13g2_buf_4 fanout3843 (.X(net3843),
    .A(net3845));
 sg13g2_buf_2 fanout3844 (.A(net3845),
    .X(net3844));
 sg13g2_buf_2 fanout3845 (.A(_03694_),
    .X(net3845));
 sg13g2_buf_4 fanout3846 (.X(net3846),
    .A(net3847));
 sg13g2_buf_4 fanout3847 (.X(net3847),
    .A(_02901_));
 sg13g2_buf_4 fanout3848 (.X(net3848),
    .A(net3849));
 sg13g2_buf_2 fanout3849 (.A(_01413_),
    .X(net3849));
 sg13g2_buf_4 fanout3850 (.X(net3850),
    .A(net3851));
 sg13g2_buf_4 fanout3851 (.X(net3851),
    .A(_01413_));
 sg13g2_buf_4 fanout3852 (.X(net3852),
    .A(_01340_));
 sg13g2_buf_2 fanout3853 (.A(_01340_),
    .X(net3853));
 sg13g2_buf_4 fanout3854 (.X(net3854),
    .A(net3855));
 sg13g2_buf_4 fanout3855 (.X(net3855),
    .A(_01339_));
 sg13g2_buf_2 fanout3856 (.A(net3857),
    .X(net3856));
 sg13g2_buf_2 fanout3857 (.A(net3859),
    .X(net3857));
 sg13g2_buf_2 fanout3858 (.A(net3859),
    .X(net3858));
 sg13g2_buf_2 fanout3859 (.A(_01269_),
    .X(net3859));
 sg13g2_buf_2 fanout3860 (.A(_01254_),
    .X(net3860));
 sg13g2_buf_4 fanout3861 (.X(net3861),
    .A(_01254_));
 sg13g2_buf_4 fanout3862 (.X(net3862),
    .A(net3864));
 sg13g2_buf_2 fanout3863 (.A(net3864),
    .X(net3863));
 sg13g2_buf_4 fanout3864 (.X(net3864),
    .A(_01243_));
 sg13g2_buf_4 fanout3865 (.X(net3865),
    .A(net3869));
 sg13g2_buf_2 fanout3866 (.A(net3869),
    .X(net3866));
 sg13g2_buf_2 fanout3867 (.A(net3868),
    .X(net3867));
 sg13g2_buf_4 fanout3868 (.X(net3868),
    .A(net3869));
 sg13g2_buf_2 fanout3869 (.A(_01243_),
    .X(net3869));
 sg13g2_buf_4 fanout3870 (.X(net3870),
    .A(_06285_));
 sg13g2_buf_2 fanout3871 (.A(net3872),
    .X(net3871));
 sg13g2_buf_1 fanout3872 (.A(net3873),
    .X(net3872));
 sg13g2_buf_1 fanout3873 (.A(net3876),
    .X(net3873));
 sg13g2_buf_2 fanout3874 (.A(net3876),
    .X(net3874));
 sg13g2_buf_1 fanout3875 (.A(net3876),
    .X(net3875));
 sg13g2_buf_1 fanout3876 (.A(_05588_),
    .X(net3876));
 sg13g2_buf_4 fanout3877 (.X(net3877),
    .A(net3878));
 sg13g2_buf_4 fanout3878 (.X(net3878),
    .A(net3879));
 sg13g2_buf_4 fanout3879 (.X(net3879),
    .A(net3882));
 sg13g2_buf_4 fanout3880 (.X(net3880),
    .A(net3881));
 sg13g2_buf_4 fanout3881 (.X(net3881),
    .A(net3882));
 sg13g2_buf_2 fanout3882 (.A(_03888_),
    .X(net3882));
 sg13g2_buf_4 fanout3883 (.X(net3883),
    .A(net3885));
 sg13g2_buf_4 fanout3884 (.X(net3884),
    .A(net3885));
 sg13g2_buf_2 fanout3885 (.A(_03888_),
    .X(net3885));
 sg13g2_buf_4 fanout3886 (.X(net3886),
    .A(net3889));
 sg13g2_buf_4 fanout3887 (.X(net3887),
    .A(net3889));
 sg13g2_buf_1 fanout3888 (.A(net3889),
    .X(net3888));
 sg13g2_buf_2 fanout3889 (.A(_03887_),
    .X(net3889));
 sg13g2_buf_4 fanout3890 (.X(net3890),
    .A(net3891));
 sg13g2_buf_2 fanout3891 (.A(net3892),
    .X(net3891));
 sg13g2_buf_4 fanout3892 (.X(net3892),
    .A(_03887_));
 sg13g2_buf_4 fanout3893 (.X(net3893),
    .A(net3894));
 sg13g2_buf_2 fanout3894 (.A(net3895),
    .X(net3894));
 sg13g2_buf_4 fanout3895 (.X(net3895),
    .A(net3896));
 sg13g2_buf_2 fanout3896 (.A(_03887_),
    .X(net3896));
 sg13g2_buf_4 fanout3897 (.X(net3897),
    .A(net3898));
 sg13g2_buf_4 fanout3898 (.X(net3898),
    .A(net3901));
 sg13g2_buf_4 fanout3899 (.X(net3899),
    .A(net3901));
 sg13g2_buf_2 fanout3900 (.A(net3901),
    .X(net3900));
 sg13g2_buf_2 fanout3901 (.A(_03884_),
    .X(net3901));
 sg13g2_buf_4 fanout3902 (.X(net3902),
    .A(net3904));
 sg13g2_buf_2 fanout3903 (.A(_03884_),
    .X(net3903));
 sg13g2_buf_2 fanout3904 (.A(_03884_),
    .X(net3904));
 sg13g2_buf_4 fanout3905 (.X(net3905),
    .A(net3906));
 sg13g2_buf_4 fanout3906 (.X(net3906),
    .A(net3907));
 sg13g2_buf_4 fanout3907 (.X(net3907),
    .A(net3912));
 sg13g2_buf_4 fanout3908 (.X(net3908),
    .A(net3909));
 sg13g2_buf_4 fanout3909 (.X(net3909),
    .A(net3912));
 sg13g2_buf_4 fanout3910 (.X(net3910),
    .A(net3911));
 sg13g2_buf_4 fanout3911 (.X(net3911),
    .A(net3912));
 sg13g2_buf_4 fanout3912 (.X(net3912),
    .A(_03883_));
 sg13g2_buf_2 fanout3913 (.A(net3915),
    .X(net3913));
 sg13g2_buf_1 fanout3914 (.A(net3915),
    .X(net3914));
 sg13g2_buf_2 fanout3915 (.A(net3917),
    .X(net3915));
 sg13g2_buf_2 fanout3916 (.A(net3917),
    .X(net3916));
 sg13g2_buf_2 fanout3917 (.A(_03877_),
    .X(net3917));
 sg13g2_buf_2 fanout3918 (.A(net3919),
    .X(net3918));
 sg13g2_buf_2 fanout3919 (.A(net3920),
    .X(net3919));
 sg13g2_buf_1 fanout3920 (.A(net3922),
    .X(net3920));
 sg13g2_buf_2 fanout3921 (.A(net3922),
    .X(net3921));
 sg13g2_buf_2 fanout3922 (.A(_03877_),
    .X(net3922));
 sg13g2_buf_4 fanout3923 (.X(net3923),
    .A(net3924));
 sg13g2_buf_2 fanout3924 (.A(net3925),
    .X(net3924));
 sg13g2_buf_2 fanout3925 (.A(net3930),
    .X(net3925));
 sg13g2_buf_4 fanout3926 (.X(net3926),
    .A(net3927));
 sg13g2_buf_1 fanout3927 (.A(net3930),
    .X(net3927));
 sg13g2_buf_2 fanout3928 (.A(net3930),
    .X(net3928));
 sg13g2_buf_1 fanout3929 (.A(net3930),
    .X(net3929));
 sg13g2_buf_2 fanout3930 (.A(_03876_),
    .X(net3930));
 sg13g2_buf_2 fanout3931 (.A(net3933),
    .X(net3931));
 sg13g2_buf_1 fanout3932 (.A(net3933),
    .X(net3932));
 sg13g2_buf_2 fanout3933 (.A(_03872_),
    .X(net3933));
 sg13g2_buf_2 fanout3934 (.A(net3937),
    .X(net3934));
 sg13g2_buf_2 fanout3935 (.A(net3936),
    .X(net3935));
 sg13g2_buf_2 fanout3936 (.A(net3937),
    .X(net3936));
 sg13g2_buf_1 fanout3937 (.A(_03870_),
    .X(net3937));
 sg13g2_buf_4 fanout3938 (.X(net3938),
    .A(net3942));
 sg13g2_buf_2 fanout3939 (.A(net3942),
    .X(net3939));
 sg13g2_buf_4 fanout3940 (.X(net3940),
    .A(net3942));
 sg13g2_buf_2 fanout3941 (.A(net3942),
    .X(net3941));
 sg13g2_buf_2 fanout3942 (.A(_03778_),
    .X(net3942));
 sg13g2_buf_4 fanout3943 (.X(net3943),
    .A(_03255_));
 sg13g2_buf_2 fanout3944 (.A(_03255_),
    .X(net3944));
 sg13g2_buf_2 fanout3945 (.A(net3946),
    .X(net3945));
 sg13g2_buf_4 fanout3946 (.X(net3946),
    .A(_03254_));
 sg13g2_buf_4 fanout3947 (.X(net3947),
    .A(_02618_));
 sg13g2_buf_2 fanout3948 (.A(_02618_),
    .X(net3948));
 sg13g2_buf_4 fanout3949 (.X(net3949),
    .A(_02617_));
 sg13g2_buf_4 fanout3950 (.X(net3950),
    .A(_02617_));
 sg13g2_buf_4 fanout3951 (.X(net3951),
    .A(_02615_));
 sg13g2_buf_4 fanout3952 (.X(net3952),
    .A(_02615_));
 sg13g2_buf_4 fanout3953 (.X(net3953),
    .A(_02614_));
 sg13g2_buf_4 fanout3954 (.X(net3954),
    .A(_02614_));
 sg13g2_buf_4 fanout3955 (.X(net3955),
    .A(_02612_));
 sg13g2_buf_4 fanout3956 (.X(net3956),
    .A(_02612_));
 sg13g2_buf_4 fanout3957 (.X(net3957),
    .A(_02610_));
 sg13g2_buf_4 fanout3958 (.X(net3958),
    .A(_02610_));
 sg13g2_buf_2 fanout3959 (.A(net3960),
    .X(net3959));
 sg13g2_buf_4 fanout3960 (.X(net3960),
    .A(net3961));
 sg13g2_buf_4 fanout3961 (.X(net3961),
    .A(_02301_));
 sg13g2_buf_4 fanout3962 (.X(net3962),
    .A(net3963));
 sg13g2_buf_4 fanout3963 (.X(net3963),
    .A(_02301_));
 sg13g2_buf_4 fanout3964 (.X(net3964),
    .A(net3965));
 sg13g2_buf_4 fanout3965 (.X(net3965),
    .A(_02300_));
 sg13g2_buf_4 fanout3966 (.X(net3966),
    .A(_02283_));
 sg13g2_buf_4 fanout3967 (.X(net3967),
    .A(_02282_));
 sg13g2_buf_2 fanout3968 (.A(_02282_),
    .X(net3968));
 sg13g2_buf_4 fanout3969 (.X(net3969),
    .A(_02158_));
 sg13g2_buf_4 fanout3970 (.X(net3970),
    .A(_02158_));
 sg13g2_buf_4 fanout3971 (.X(net3971),
    .A(_02157_));
 sg13g2_buf_4 fanout3972 (.X(net3972),
    .A(_02157_));
 sg13g2_buf_4 fanout3973 (.X(net3973),
    .A(net3974));
 sg13g2_buf_4 fanout3974 (.X(net3974),
    .A(_02153_));
 sg13g2_buf_4 fanout3975 (.X(net3975),
    .A(_02152_));
 sg13g2_buf_4 fanout3976 (.X(net3976),
    .A(_02152_));
 sg13g2_buf_4 fanout3977 (.X(net3977),
    .A(_02149_));
 sg13g2_buf_4 fanout3978 (.X(net3978),
    .A(_02149_));
 sg13g2_buf_4 fanout3979 (.X(net3979),
    .A(_02148_));
 sg13g2_buf_4 fanout3980 (.X(net3980),
    .A(_02148_));
 sg13g2_buf_4 fanout3981 (.X(net3981),
    .A(_02143_));
 sg13g2_buf_4 fanout3982 (.X(net3982),
    .A(_02143_));
 sg13g2_buf_4 fanout3983 (.X(net3983),
    .A(net3985));
 sg13g2_buf_4 fanout3984 (.X(net3984),
    .A(net3985));
 sg13g2_buf_2 fanout3985 (.A(_02137_),
    .X(net3985));
 sg13g2_buf_4 fanout3986 (.X(net3986),
    .A(_02134_));
 sg13g2_buf_2 fanout3987 (.A(_02134_),
    .X(net3987));
 sg13g2_buf_4 fanout3988 (.X(net3988),
    .A(net3990));
 sg13g2_buf_4 fanout3989 (.X(net3989),
    .A(net3990));
 sg13g2_buf_2 fanout3990 (.A(_02015_),
    .X(net3990));
 sg13g2_buf_4 fanout3991 (.X(net3991),
    .A(net3992));
 sg13g2_buf_2 fanout3992 (.A(_02011_),
    .X(net3992));
 sg13g2_buf_2 fanout3993 (.A(net3994),
    .X(net3993));
 sg13g2_buf_4 fanout3994 (.X(net3994),
    .A(_02011_));
 sg13g2_buf_4 fanout3995 (.X(net3995),
    .A(_01924_));
 sg13g2_buf_4 fanout3996 (.X(net3996),
    .A(_01924_));
 sg13g2_buf_4 fanout3997 (.X(net3997),
    .A(net3999));
 sg13g2_buf_4 fanout3998 (.X(net3998),
    .A(net3999));
 sg13g2_buf_2 fanout3999 (.A(_01435_),
    .X(net3999));
 sg13g2_buf_2 fanout4000 (.A(net4001),
    .X(net4000));
 sg13g2_buf_2 fanout4001 (.A(net4002),
    .X(net4001));
 sg13g2_buf_2 fanout4002 (.A(net4003),
    .X(net4002));
 sg13g2_buf_4 fanout4003 (.X(net4003),
    .A(_01412_));
 sg13g2_buf_4 fanout4004 (.X(net4004),
    .A(net4008));
 sg13g2_buf_4 fanout4005 (.X(net4005),
    .A(net4007));
 sg13g2_buf_2 fanout4006 (.A(net4008),
    .X(net4006));
 sg13g2_buf_2 fanout4007 (.A(net4008),
    .X(net4007));
 sg13g2_buf_2 fanout4008 (.A(_01412_),
    .X(net4008));
 sg13g2_buf_2 fanout4009 (.A(net4010),
    .X(net4009));
 sg13g2_buf_4 fanout4010 (.X(net4010),
    .A(net4011));
 sg13g2_buf_2 fanout4011 (.A(net4013),
    .X(net4011));
 sg13g2_buf_2 fanout4012 (.A(net4013),
    .X(net4012));
 sg13g2_buf_2 fanout4013 (.A(net4021),
    .X(net4013));
 sg13g2_buf_4 fanout4014 (.X(net4014),
    .A(net4015));
 sg13g2_buf_4 fanout4015 (.X(net4015),
    .A(net4021));
 sg13g2_buf_2 fanout4016 (.A(net4017),
    .X(net4016));
 sg13g2_buf_2 fanout4017 (.A(net4018),
    .X(net4017));
 sg13g2_buf_2 fanout4018 (.A(net4021),
    .X(net4018));
 sg13g2_buf_2 fanout4019 (.A(net4021),
    .X(net4019));
 sg13g2_buf_1 fanout4020 (.A(net4021),
    .X(net4020));
 sg13g2_buf_4 fanout4021 (.X(net4021),
    .A(_01411_));
 sg13g2_buf_4 fanout4022 (.X(net4022),
    .A(net4024));
 sg13g2_buf_2 fanout4023 (.A(net4024),
    .X(net4023));
 sg13g2_buf_2 fanout4024 (.A(_00000_),
    .X(net4024));
 sg13g2_buf_2 fanout4025 (.A(_01391_),
    .X(net4025));
 sg13g2_buf_2 fanout4026 (.A(net4027),
    .X(net4026));
 sg13g2_buf_2 fanout4027 (.A(_01386_),
    .X(net4027));
 sg13g2_buf_4 fanout4028 (.X(net4028),
    .A(_01353_));
 sg13g2_buf_2 fanout4029 (.A(_01343_),
    .X(net4029));
 sg13g2_buf_2 fanout4030 (.A(_01343_),
    .X(net4030));
 sg13g2_buf_4 fanout4031 (.X(net4031),
    .A(net4032));
 sg13g2_buf_4 fanout4032 (.X(net4032),
    .A(net4034));
 sg13g2_buf_4 fanout4033 (.X(net4033),
    .A(net4034));
 sg13g2_buf_2 fanout4034 (.A(_01265_),
    .X(net4034));
 sg13g2_buf_4 fanout4035 (.X(net4035),
    .A(net4037));
 sg13g2_buf_4 fanout4036 (.X(net4036),
    .A(net4037));
 sg13g2_buf_4 fanout4037 (.X(net4037),
    .A(_01259_));
 sg13g2_buf_4 fanout4038 (.X(net4038),
    .A(net4039));
 sg13g2_buf_4 fanout4039 (.X(net4039),
    .A(_01258_));
 sg13g2_buf_2 fanout4040 (.A(net4043),
    .X(net4040));
 sg13g2_buf_2 fanout4041 (.A(net4043),
    .X(net4041));
 sg13g2_buf_1 fanout4042 (.A(net4043),
    .X(net4042));
 sg13g2_buf_2 fanout4043 (.A(net4059),
    .X(net4043));
 sg13g2_buf_2 fanout4044 (.A(net4045),
    .X(net4044));
 sg13g2_buf_2 fanout4045 (.A(net4059),
    .X(net4045));
 sg13g2_buf_2 fanout4046 (.A(net4050),
    .X(net4046));
 sg13g2_buf_4 fanout4047 (.X(net4047),
    .A(net4049));
 sg13g2_buf_2 fanout4048 (.A(net4049),
    .X(net4048));
 sg13g2_buf_2 fanout4049 (.A(net4050),
    .X(net4049));
 sg13g2_buf_2 fanout4050 (.A(net4059),
    .X(net4050));
 sg13g2_buf_2 fanout4051 (.A(net4053),
    .X(net4051));
 sg13g2_buf_2 fanout4052 (.A(net4053),
    .X(net4052));
 sg13g2_buf_2 fanout4053 (.A(net4059),
    .X(net4053));
 sg13g2_buf_2 fanout4054 (.A(net4058),
    .X(net4054));
 sg13g2_buf_2 fanout4055 (.A(net4058),
    .X(net4055));
 sg13g2_buf_4 fanout4056 (.X(net4056),
    .A(net4058));
 sg13g2_buf_2 fanout4057 (.A(net4058),
    .X(net4057));
 sg13g2_buf_2 fanout4058 (.A(net4059),
    .X(net4058));
 sg13g2_buf_4 fanout4059 (.X(net4059),
    .A(_01242_));
 sg13g2_buf_2 fanout4060 (.A(net4061),
    .X(net4060));
 sg13g2_buf_2 fanout4061 (.A(net4066),
    .X(net4061));
 sg13g2_buf_4 fanout4062 (.X(net4062),
    .A(net4066));
 sg13g2_buf_4 fanout4063 (.X(net4063),
    .A(net4064));
 sg13g2_buf_2 fanout4064 (.A(net4065),
    .X(net4064));
 sg13g2_buf_4 fanout4065 (.X(net4065),
    .A(net4066));
 sg13g2_buf_2 fanout4066 (.A(_01238_),
    .X(net4066));
 sg13g2_buf_4 fanout4067 (.X(net4067),
    .A(_01237_));
 sg13g2_buf_4 fanout4068 (.X(net4068),
    .A(net4069));
 sg13g2_buf_4 fanout4069 (.X(net4069),
    .A(_01232_));
 sg13g2_buf_4 fanout4070 (.X(net4070),
    .A(net4073));
 sg13g2_buf_2 fanout4071 (.A(net4073),
    .X(net4071));
 sg13g2_buf_4 fanout4072 (.X(net4072),
    .A(net4073));
 sg13g2_buf_2 fanout4073 (.A(_01232_),
    .X(net4073));
 sg13g2_buf_4 fanout4074 (.X(net4074),
    .A(_01231_));
 sg13g2_buf_2 fanout4075 (.A(_01231_),
    .X(net4075));
 sg13g2_buf_4 fanout4076 (.X(net4076),
    .A(_01231_));
 sg13g2_buf_2 fanout4077 (.A(net4080),
    .X(net4077));
 sg13g2_buf_2 fanout4078 (.A(net4080),
    .X(net4078));
 sg13g2_buf_2 fanout4079 (.A(net4080),
    .X(net4079));
 sg13g2_buf_2 fanout4080 (.A(_01228_),
    .X(net4080));
 sg13g2_buf_2 fanout4081 (.A(\uart_receiver/_206_ ),
    .X(net4081));
 sg13g2_buf_2 fanout4082 (.A(\uart_receiver/_206_ ),
    .X(net4082));
 sg13g2_buf_2 fanout4083 (.A(\uart_receiver/_127_ ),
    .X(net4083));
 sg13g2_buf_2 fanout4084 (.A(\uart_receiver/_108_ ),
    .X(net4084));
 sg13g2_buf_4 fanout4085 (.X(net4085),
    .A(_06448_));
 sg13g2_buf_2 fanout4086 (.A(_06448_),
    .X(net4086));
 sg13g2_buf_2 fanout4087 (.A(net4088),
    .X(net4087));
 sg13g2_buf_4 fanout4088 (.X(net4088),
    .A(_06448_));
 sg13g2_buf_2 fanout4089 (.A(net4090),
    .X(net4089));
 sg13g2_buf_4 fanout4090 (.X(net4090),
    .A(_03871_));
 sg13g2_buf_2 fanout4091 (.A(net4092),
    .X(net4091));
 sg13g2_buf_2 fanout4092 (.A(_03869_),
    .X(net4092));
 sg13g2_buf_2 fanout4093 (.A(net4094),
    .X(net4093));
 sg13g2_buf_4 fanout4094 (.X(net4094),
    .A(_03867_));
 sg13g2_buf_4 fanout4095 (.X(net4095),
    .A(_02607_));
 sg13g2_buf_4 fanout4096 (.X(net4096),
    .A(_02607_));
 sg13g2_buf_2 fanout4097 (.A(net4098),
    .X(net4097));
 sg13g2_buf_2 fanout4098 (.A(net4099),
    .X(net4098));
 sg13g2_buf_2 fanout4099 (.A(net4101),
    .X(net4099));
 sg13g2_buf_4 fanout4100 (.X(net4100),
    .A(net4101));
 sg13g2_buf_2 fanout4101 (.A(net4109),
    .X(net4101));
 sg13g2_buf_4 fanout4102 (.X(net4102),
    .A(net4109));
 sg13g2_buf_2 fanout4103 (.A(net4109),
    .X(net4103));
 sg13g2_buf_4 fanout4104 (.X(net4104),
    .A(net4105));
 sg13g2_buf_2 fanout4105 (.A(net4109),
    .X(net4105));
 sg13g2_buf_4 fanout4106 (.X(net4106),
    .A(net4107));
 sg13g2_buf_4 fanout4107 (.X(net4107),
    .A(net4108));
 sg13g2_buf_2 fanout4108 (.A(net4109),
    .X(net4108));
 sg13g2_buf_4 fanout4109 (.X(net4109),
    .A(_02325_));
 sg13g2_buf_2 fanout4110 (.A(net4111),
    .X(net4110));
 sg13g2_buf_2 fanout4111 (.A(net4112),
    .X(net4111));
 sg13g2_buf_2 fanout4112 (.A(net4114),
    .X(net4112));
 sg13g2_buf_2 fanout4113 (.A(net4114),
    .X(net4113));
 sg13g2_buf_2 fanout4114 (.A(net4122),
    .X(net4114));
 sg13g2_buf_4 fanout4115 (.X(net4115),
    .A(net4116));
 sg13g2_buf_4 fanout4116 (.X(net4116),
    .A(net4122));
 sg13g2_buf_2 fanout4117 (.A(net4118),
    .X(net4117));
 sg13g2_buf_2 fanout4118 (.A(net4122),
    .X(net4118));
 sg13g2_buf_2 fanout4119 (.A(net4120),
    .X(net4119));
 sg13g2_buf_2 fanout4120 (.A(net4121),
    .X(net4120));
 sg13g2_buf_2 fanout4121 (.A(net4122),
    .X(net4121));
 sg13g2_buf_4 fanout4122 (.X(net4122),
    .A(_02281_));
 sg13g2_buf_4 fanout4123 (.X(net4123),
    .A(net4124));
 sg13g2_buf_4 fanout4124 (.X(net4124),
    .A(_02156_));
 sg13g2_buf_4 fanout4125 (.X(net4125),
    .A(net4127));
 sg13g2_buf_4 fanout4126 (.X(net4126),
    .A(net4127));
 sg13g2_buf_8 fanout4127 (.A(_02155_),
    .X(net4127));
 sg13g2_buf_8 fanout4128 (.A(net4129),
    .X(net4128));
 sg13g2_buf_8 fanout4129 (.A(_02151_),
    .X(net4129));
 sg13g2_buf_4 fanout4130 (.X(net4130),
    .A(net4131));
 sg13g2_buf_4 fanout4131 (.X(net4131),
    .A(_02146_));
 sg13g2_buf_8 fanout4132 (.A(net4133),
    .X(net4132));
 sg13g2_buf_8 fanout4133 (.A(_02142_),
    .X(net4133));
 sg13g2_buf_4 fanout4134 (.X(net4134),
    .A(_01920_));
 sg13g2_buf_2 fanout4135 (.A(_01920_),
    .X(net4135));
 sg13g2_buf_4 fanout4136 (.X(net4136),
    .A(net4137));
 sg13g2_buf_2 fanout4137 (.A(_01920_),
    .X(net4137));
 sg13g2_buf_2 fanout4138 (.A(net4139),
    .X(net4138));
 sg13g2_buf_2 fanout4139 (.A(_01408_),
    .X(net4139));
 sg13g2_buf_4 fanout4140 (.X(net4140),
    .A(net4141));
 sg13g2_buf_2 fanout4141 (.A(_01408_),
    .X(net4141));
 sg13g2_buf_2 fanout4142 (.A(net4143),
    .X(net4142));
 sg13g2_buf_4 fanout4143 (.X(net4143),
    .A(_01408_));
 sg13g2_buf_2 fanout4144 (.A(_01382_),
    .X(net4144));
 sg13g2_buf_2 fanout4145 (.A(_01382_),
    .X(net4145));
 sg13g2_buf_2 fanout4146 (.A(_01369_),
    .X(net4146));
 sg13g2_buf_2 fanout4147 (.A(_01369_),
    .X(net4147));
 sg13g2_buf_4 fanout4148 (.X(net4148),
    .A(net4149));
 sg13g2_buf_4 fanout4149 (.X(net4149),
    .A(_01362_));
 sg13g2_buf_4 fanout4150 (.X(net4150),
    .A(_01281_));
 sg13g2_buf_4 fanout4151 (.X(net4151),
    .A(_01179_));
 sg13g2_buf_4 fanout4152 (.X(net4152),
    .A(_01178_));
 sg13g2_buf_4 fanout4153 (.X(net4153),
    .A(_01177_));
 sg13g2_buf_4 fanout4154 (.X(net4154),
    .A(_01176_));
 sg13g2_buf_4 fanout4155 (.X(net4155),
    .A(_01174_));
 sg13g2_buf_4 fanout4156 (.X(net4156),
    .A(_01172_));
 sg13g2_buf_2 fanout4157 (.A(net4158),
    .X(net4157));
 sg13g2_buf_2 fanout4158 (.A(_01046_),
    .X(net4158));
 sg13g2_buf_2 fanout4159 (.A(net4160),
    .X(net4159));
 sg13g2_buf_1 fanout4160 (.A(_01046_),
    .X(net4160));
 sg13g2_buf_2 fanout4161 (.A(net4162),
    .X(net4161));
 sg13g2_buf_2 fanout4162 (.A(net4163),
    .X(net4162));
 sg13g2_buf_4 fanout4163 (.X(net4163),
    .A(_01036_));
 sg13g2_buf_2 fanout4164 (.A(net4165),
    .X(net4164));
 sg13g2_buf_2 fanout4165 (.A(net4166),
    .X(net4165));
 sg13g2_buf_1 fanout4166 (.A(net4167),
    .X(net4166));
 sg13g2_buf_2 fanout4167 (.A(_01028_),
    .X(net4167));
 sg13g2_buf_2 fanout4168 (.A(net4170),
    .X(net4168));
 sg13g2_buf_2 fanout4169 (.A(net4170),
    .X(net4169));
 sg13g2_buf_2 fanout4170 (.A(_01028_),
    .X(net4170));
 sg13g2_buf_4 fanout4171 (.X(net4171),
    .A(net4173));
 sg13g2_buf_4 fanout4172 (.X(net4172),
    .A(net4173));
 sg13g2_buf_2 fanout4173 (.A(net4179),
    .X(net4173));
 sg13g2_buf_4 fanout4174 (.X(net4174),
    .A(net4176));
 sg13g2_buf_4 fanout4175 (.X(net4175),
    .A(net4176));
 sg13g2_buf_2 fanout4176 (.A(net4178),
    .X(net4176));
 sg13g2_buf_4 fanout4177 (.X(net4177),
    .A(net4178));
 sg13g2_buf_1 fanout4178 (.A(net4179),
    .X(net4178));
 sg13g2_buf_2 fanout4179 (.A(_01019_),
    .X(net4179));
 sg13g2_buf_4 fanout4180 (.X(net4180),
    .A(net4190));
 sg13g2_buf_2 fanout4181 (.A(net4190),
    .X(net4181));
 sg13g2_buf_4 fanout4182 (.X(net4182),
    .A(net4183));
 sg13g2_buf_2 fanout4183 (.A(net4184),
    .X(net4183));
 sg13g2_buf_1 fanout4184 (.A(net4190),
    .X(net4184));
 sg13g2_buf_2 fanout4185 (.A(net4187),
    .X(net4185));
 sg13g2_buf_1 fanout4186 (.A(net4187),
    .X(net4186));
 sg13g2_buf_4 fanout4187 (.X(net4187),
    .A(net4189));
 sg13g2_buf_4 fanout4188 (.X(net4188),
    .A(net4189));
 sg13g2_buf_2 fanout4189 (.A(net4190),
    .X(net4189));
 sg13g2_buf_2 fanout4190 (.A(_01011_),
    .X(net4190));
 sg13g2_buf_2 fanout4191 (.A(net4193),
    .X(net4191));
 sg13g2_buf_1 fanout4192 (.A(net4193),
    .X(net4192));
 sg13g2_buf_2 fanout4193 (.A(net4196),
    .X(net4193));
 sg13g2_buf_2 fanout4194 (.A(net4195),
    .X(net4194));
 sg13g2_buf_2 fanout4195 (.A(net4196),
    .X(net4195));
 sg13g2_buf_2 fanout4196 (.A(_01003_),
    .X(net4196));
 sg13g2_buf_2 fanout4197 (.A(net4198),
    .X(net4197));
 sg13g2_buf_2 fanout4198 (.A(net4199),
    .X(net4198));
 sg13g2_buf_1 fanout4199 (.A(net4200),
    .X(net4199));
 sg13g2_buf_4 fanout4200 (.X(net4200),
    .A(_01003_));
 sg13g2_buf_8 fanout4201 (.A(_00906_),
    .X(net4201));
 sg13g2_buf_4 fanout4202 (.X(net4202),
    .A(net4203));
 sg13g2_buf_2 fanout4203 (.A(_00895_),
    .X(net4203));
 sg13g2_buf_2 fanout4204 (.A(net4205),
    .X(net4204));
 sg13g2_buf_2 fanout4205 (.A(_00895_),
    .X(net4205));
 sg13g2_buf_4 fanout4206 (.X(net4206),
    .A(net4207));
 sg13g2_buf_8 fanout4207 (.A(net4212),
    .X(net4207));
 sg13g2_buf_4 fanout4208 (.X(net4208),
    .A(net4212));
 sg13g2_buf_4 fanout4209 (.X(net4209),
    .A(net4212));
 sg13g2_buf_2 fanout4210 (.A(net4211),
    .X(net4210));
 sg13g2_buf_4 fanout4211 (.X(net4211),
    .A(net4212));
 sg13g2_buf_4 fanout4212 (.X(net4212),
    .A(_00893_));
 sg13g2_buf_4 fanout4213 (.X(net4213),
    .A(net4215));
 sg13g2_buf_2 fanout4214 (.A(net4215),
    .X(net4214));
 sg13g2_buf_4 fanout4215 (.X(net4215),
    .A(net4217));
 sg13g2_buf_8 fanout4216 (.A(net4217),
    .X(net4216));
 sg13g2_buf_2 fanout4217 (.A(_00892_),
    .X(net4217));
 sg13g2_buf_2 fanout4218 (.A(net4219),
    .X(net4218));
 sg13g2_buf_4 fanout4219 (.X(net4219),
    .A(net4220));
 sg13g2_buf_4 fanout4220 (.X(net4220),
    .A(_00892_));
 sg13g2_buf_2 fanout4221 (.A(net4224),
    .X(net4221));
 sg13g2_buf_2 fanout4222 (.A(net4224),
    .X(net4222));
 sg13g2_buf_1 fanout4223 (.A(net4224),
    .X(net4223));
 sg13g2_buf_2 fanout4224 (.A(net4230),
    .X(net4224));
 sg13g2_buf_2 fanout4225 (.A(net4226),
    .X(net4225));
 sg13g2_buf_2 fanout4226 (.A(net4230),
    .X(net4226));
 sg13g2_buf_2 fanout4227 (.A(net4230),
    .X(net4227));
 sg13g2_buf_2 fanout4228 (.A(net4230),
    .X(net4228));
 sg13g2_buf_2 fanout4229 (.A(net4230),
    .X(net4229));
 sg13g2_buf_2 fanout4230 (.A(_00889_),
    .X(net4230));
 sg13g2_buf_2 fanout4231 (.A(net4232),
    .X(net4231));
 sg13g2_buf_2 fanout4232 (.A(net4233),
    .X(net4232));
 sg13g2_buf_2 fanout4233 (.A(_00889_),
    .X(net4233));
 sg13g2_buf_4 fanout4234 (.X(net4234),
    .A(net4236));
 sg13g2_buf_4 fanout4235 (.X(net4235),
    .A(net4236));
 sg13g2_buf_2 fanout4236 (.A(_00889_),
    .X(net4236));
 sg13g2_buf_2 fanout4237 (.A(net4238),
    .X(net4237));
 sg13g2_buf_2 fanout4238 (.A(net4239),
    .X(net4238));
 sg13g2_buf_4 fanout4239 (.X(net4239),
    .A(net4241));
 sg13g2_buf_2 fanout4240 (.A(net4241),
    .X(net4240));
 sg13g2_buf_2 fanout4241 (.A(_00887_),
    .X(net4241));
 sg13g2_buf_4 fanout4242 (.X(net4242),
    .A(_00886_));
 sg13g2_buf_2 fanout4243 (.A(_00886_),
    .X(net4243));
 sg13g2_buf_4 fanout4244 (.X(net4244),
    .A(net4254));
 sg13g2_buf_2 fanout4245 (.A(net4254),
    .X(net4245));
 sg13g2_buf_2 fanout4246 (.A(net4250),
    .X(net4246));
 sg13g2_buf_2 fanout4247 (.A(net4249),
    .X(net4247));
 sg13g2_buf_1 fanout4248 (.A(net4249),
    .X(net4248));
 sg13g2_buf_2 fanout4249 (.A(net4250),
    .X(net4249));
 sg13g2_buf_2 fanout4250 (.A(net4254),
    .X(net4250));
 sg13g2_buf_4 fanout4251 (.X(net4251),
    .A(net4253));
 sg13g2_buf_2 fanout4252 (.A(net4253),
    .X(net4252));
 sg13g2_buf_2 fanout4253 (.A(net4254),
    .X(net4253));
 sg13g2_buf_2 fanout4254 (.A(_00885_),
    .X(net4254));
 sg13g2_buf_2 fanout4255 (.A(net4256),
    .X(net4255));
 sg13g2_buf_4 fanout4256 (.X(net4256),
    .A(net4257));
 sg13g2_buf_2 fanout4257 (.A(net4258),
    .X(net4257));
 sg13g2_buf_2 fanout4258 (.A(_00885_),
    .X(net4258));
 sg13g2_buf_2 fanout4259 (.A(net4261),
    .X(net4259));
 sg13g2_buf_2 fanout4260 (.A(net4261),
    .X(net4260));
 sg13g2_buf_2 fanout4261 (.A(net4262),
    .X(net4261));
 sg13g2_buf_4 fanout4262 (.X(net4262),
    .A(net4263));
 sg13g2_buf_4 fanout4263 (.X(net4263),
    .A(net4266));
 sg13g2_buf_4 fanout4264 (.X(net4264),
    .A(net4266));
 sg13g2_buf_2 fanout4265 (.A(net4266),
    .X(net4265));
 sg13g2_buf_4 fanout4266 (.X(net4266),
    .A(_00885_));
 sg13g2_buf_2 fanout4267 (.A(net918),
    .X(net4267));
 sg13g2_buf_4 fanout4268 (.X(net4268),
    .A(_00145_));
 sg13g2_buf_4 fanout4269 (.X(net4269),
    .A(net4271));
 sg13g2_buf_2 fanout4270 (.A(net4271),
    .X(net4270));
 sg13g2_buf_2 fanout4271 (.A(_00145_),
    .X(net4271));
 sg13g2_buf_4 fanout4272 (.X(net4272),
    .A(net4273));
 sg13g2_buf_4 fanout4273 (.X(net4273),
    .A(net4274));
 sg13g2_buf_4 fanout4274 (.X(net4274),
    .A(net497));
 sg13g2_buf_4 fanout4275 (.X(net4275),
    .A(net4276));
 sg13g2_buf_4 fanout4276 (.X(net4276),
    .A(_00143_));
 sg13g2_buf_2 fanout4277 (.A(net4278),
    .X(net4277));
 sg13g2_buf_2 fanout4278 (.A(net4279),
    .X(net4278));
 sg13g2_buf_4 fanout4279 (.X(net4279),
    .A(_00142_));
 sg13g2_buf_2 fanout4280 (.A(_00142_),
    .X(net4280));
 sg13g2_buf_2 fanout4281 (.A(net4282),
    .X(net4281));
 sg13g2_buf_2 fanout4282 (.A(net4283),
    .X(net4282));
 sg13g2_buf_2 fanout4283 (.A(net4285),
    .X(net4283));
 sg13g2_buf_2 fanout4284 (.A(net4285),
    .X(net4284));
 sg13g2_buf_2 fanout4285 (.A(_00141_),
    .X(net4285));
 sg13g2_buf_4 fanout4286 (.X(net4286),
    .A(net4287));
 sg13g2_buf_2 fanout4287 (.A(net4288),
    .X(net4287));
 sg13g2_buf_4 fanout4288 (.X(net4288),
    .A(net4289));
 sg13g2_buf_4 fanout4289 (.X(net4289),
    .A(_00140_));
 sg13g2_buf_4 fanout4290 (.X(net4290),
    .A(net4291));
 sg13g2_buf_2 fanout4291 (.A(net4292),
    .X(net4291));
 sg13g2_buf_2 fanout4292 (.A(net4293),
    .X(net4292));
 sg13g2_buf_4 fanout4293 (.X(net4293),
    .A(_00139_));
 sg13g2_buf_2 fanout4294 (.A(net4295),
    .X(net4294));
 sg13g2_buf_2 fanout4295 (.A(net4296),
    .X(net4295));
 sg13g2_buf_2 fanout4296 (.A(net4298),
    .X(net4296));
 sg13g2_buf_4 fanout4297 (.X(net4297),
    .A(net4298));
 sg13g2_buf_4 fanout4298 (.X(net4298),
    .A(_00138_));
 sg13g2_buf_4 fanout4299 (.X(net4299),
    .A(net4301));
 sg13g2_buf_4 fanout4300 (.X(net4300),
    .A(\cpu.execution_stage[5] ));
 sg13g2_buf_4 fanout4301 (.X(net4301),
    .A(\cpu.execution_stage[5] ));
 sg13g2_buf_4 fanout4302 (.X(net4302),
    .A(\cpu.execution_stage[4] ));
 sg13g2_buf_2 fanout4303 (.A(\cpu.execution_stage[4] ),
    .X(net4303));
 sg13g2_buf_2 fanout4304 (.A(net4305),
    .X(net4304));
 sg13g2_buf_4 fanout4305 (.X(net4305),
    .A(net4308));
 sg13g2_buf_2 fanout4306 (.A(net4307),
    .X(net4306));
 sg13g2_buf_2 fanout4307 (.A(net4308),
    .X(net4307));
 sg13g2_buf_2 fanout4308 (.A(\cpu.execution_stage[3] ),
    .X(net4308));
 sg13g2_buf_4 fanout4309 (.X(net4309),
    .A(net4311));
 sg13g2_buf_2 fanout4310 (.A(net4311),
    .X(net4310));
 sg13g2_buf_2 fanout4311 (.A(net398),
    .X(net4311));
 sg13g2_buf_4 fanout4312 (.X(net4312),
    .A(_00016_));
 sg13g2_buf_4 fanout4313 (.X(net4313),
    .A(net4314));
 sg13g2_buf_4 fanout4314 (.X(net4314),
    .A(\cpu.execution_stage[2] ));
 sg13g2_buf_4 fanout4315 (.X(net4315),
    .A(net4318));
 sg13g2_buf_2 fanout4316 (.A(net4317),
    .X(net4316));
 sg13g2_buf_2 fanout4317 (.A(net4318),
    .X(net4317));
 sg13g2_buf_4 fanout4318 (.X(net4318),
    .A(\cpu.execution_stage[2] ));
 sg13g2_buf_4 fanout4319 (.X(net4319),
    .A(net4320));
 sg13g2_buf_2 fanout4320 (.A(net4321),
    .X(net4320));
 sg13g2_buf_4 fanout4321 (.X(net4321),
    .A(\cpu.execution_stage[2] ));
 sg13g2_buf_2 fanout4322 (.A(net4324),
    .X(net4322));
 sg13g2_buf_2 fanout4323 (.A(net4324),
    .X(net4323));
 sg13g2_buf_2 fanout4324 (.A(net4325),
    .X(net4324));
 sg13g2_buf_2 fanout4325 (.A(\cpu.memory_ready ),
    .X(net4325));
 sg13g2_buf_2 fanout4326 (.A(net4330),
    .X(net4326));
 sg13g2_buf_2 fanout4327 (.A(net4328),
    .X(net4327));
 sg13g2_buf_2 fanout4328 (.A(net4330),
    .X(net4328));
 sg13g2_buf_2 fanout4329 (.A(net4330),
    .X(net4329));
 sg13g2_buf_4 fanout4330 (.X(net4330),
    .A(\cpu.memory_ready ));
 sg13g2_buf_2 fanout4331 (.A(net314),
    .X(net4331));
 sg13g2_buf_2 fanout4332 (.A(\memory_controller.state[4] ),
    .X(net4332));
 sg13g2_buf_2 fanout4333 (.A(\memory_controller.state[0] ),
    .X(net4333));
 sg13g2_buf_4 fanout4334 (.X(net4334),
    .A(\cpu.write_complete ));
 sg13g2_buf_4 fanout4335 (.X(net4335),
    .A(\cpu.write_complete ));
 sg13g2_buf_2 fanout4336 (.A(net4337),
    .X(net4336));
 sg13g2_buf_4 fanout4337 (.X(net4337),
    .A(net4338));
 sg13g2_buf_4 fanout4338 (.X(net4338),
    .A(_00137_));
 sg13g2_buf_4 fanout4339 (.X(net4339),
    .A(net4341));
 sg13g2_buf_2 fanout4340 (.A(net4341),
    .X(net4340));
 sg13g2_buf_2 fanout4341 (.A(net4342),
    .X(net4341));
 sg13g2_buf_4 fanout4342 (.X(net4342),
    .A(net846));
 sg13g2_buf_4 fanout4343 (.X(net4343),
    .A(net4345));
 sg13g2_buf_2 fanout4344 (.A(net4345),
    .X(net4344));
 sg13g2_buf_4 fanout4345 (.X(net4345),
    .A(net4346));
 sg13g2_buf_4 fanout4346 (.X(net4346),
    .A(net922));
 sg13g2_buf_4 fanout4347 (.X(net4347),
    .A(net4348));
 sg13g2_buf_4 fanout4348 (.X(net4348),
    .A(net4349));
 sg13g2_buf_2 fanout4349 (.A(net851),
    .X(net4349));
 sg13g2_buf_4 fanout4350 (.X(net4350),
    .A(net4352));
 sg13g2_buf_4 fanout4351 (.X(net4351),
    .A(net4352));
 sg13g2_buf_4 fanout4352 (.X(net4352),
    .A(net787));
 sg13g2_buf_4 fanout4353 (.X(net4353),
    .A(net4357));
 sg13g2_buf_2 fanout4354 (.A(net4357),
    .X(net4354));
 sg13g2_buf_4 fanout4355 (.X(net4355),
    .A(net4357));
 sg13g2_buf_4 fanout4356 (.X(net4356),
    .A(net4357));
 sg13g2_buf_4 fanout4357 (.X(net4357),
    .A(_00132_));
 sg13g2_buf_4 fanout4358 (.X(net4358),
    .A(net4359));
 sg13g2_buf_2 fanout4359 (.A(net4360),
    .X(net4359));
 sg13g2_buf_2 fanout4360 (.A(net4361),
    .X(net4360));
 sg13g2_buf_4 fanout4361 (.X(net4361),
    .A(_00131_));
 sg13g2_buf_4 fanout4362 (.X(net4362),
    .A(net937));
 sg13g2_buf_4 fanout4363 (.X(net4363),
    .A(net4365));
 sg13g2_buf_2 fanout4364 (.A(net4365),
    .X(net4364));
 sg13g2_buf_8 fanout4365 (.A(net642),
    .X(net4365));
 sg13g2_buf_4 fanout4366 (.X(net4366),
    .A(net4367));
 sg13g2_buf_4 fanout4367 (.X(net4367),
    .A(net4368));
 sg13g2_buf_4 fanout4368 (.X(net4368),
    .A(net4370));
 sg13g2_buf_4 fanout4369 (.X(net4369),
    .A(net4370));
 sg13g2_buf_8 fanout4370 (.A(\cpu.current_instruction[15] ),
    .X(net4370));
 sg13g2_buf_2 fanout4371 (.A(net4373),
    .X(net4371));
 sg13g2_buf_2 fanout4372 (.A(net4373),
    .X(net4372));
 sg13g2_buf_2 fanout4373 (.A(net4375),
    .X(net4373));
 sg13g2_buf_2 fanout4374 (.A(net4375),
    .X(net4374));
 sg13g2_buf_2 fanout4375 (.A(net4381),
    .X(net4375));
 sg13g2_buf_4 fanout4376 (.X(net4376),
    .A(net4381));
 sg13g2_buf_4 fanout4377 (.X(net4377),
    .A(net4379));
 sg13g2_buf_2 fanout4378 (.A(net4379),
    .X(net4378));
 sg13g2_buf_4 fanout4379 (.X(net4379),
    .A(net4380));
 sg13g2_buf_2 fanout4380 (.A(net4381),
    .X(net4380));
 sg13g2_buf_2 fanout4381 (.A(\cpu.current_instruction[14] ),
    .X(net4381));
 sg13g2_buf_4 fanout4382 (.X(net4382),
    .A(net4383));
 sg13g2_buf_4 fanout4383 (.X(net4383),
    .A(net4387));
 sg13g2_buf_4 fanout4384 (.X(net4384),
    .A(net4386));
 sg13g2_buf_4 fanout4385 (.X(net4385),
    .A(net4386));
 sg13g2_buf_2 fanout4386 (.A(net4387),
    .X(net4386));
 sg13g2_buf_2 fanout4387 (.A(\cpu.current_instruction[14] ),
    .X(net4387));
 sg13g2_buf_2 fanout4388 (.A(net4389),
    .X(net4388));
 sg13g2_buf_2 fanout4389 (.A(net4390),
    .X(net4389));
 sg13g2_buf_2 fanout4390 (.A(net4395),
    .X(net4390));
 sg13g2_buf_2 fanout4391 (.A(net4395),
    .X(net4391));
 sg13g2_buf_2 fanout4392 (.A(net4395),
    .X(net4392));
 sg13g2_buf_4 fanout4393 (.X(net4393),
    .A(net4394));
 sg13g2_buf_4 fanout4394 (.X(net4394),
    .A(net4395));
 sg13g2_buf_4 fanout4395 (.X(net4395),
    .A(net4402));
 sg13g2_buf_8 fanout4396 (.A(net4402),
    .X(net4396));
 sg13g2_buf_2 fanout4397 (.A(net4398),
    .X(net4397));
 sg13g2_buf_2 fanout4398 (.A(net4402),
    .X(net4398));
 sg13g2_buf_2 fanout4399 (.A(net4401),
    .X(net4399));
 sg13g2_buf_2 fanout4400 (.A(net4401),
    .X(net4400));
 sg13g2_buf_2 fanout4401 (.A(net4402),
    .X(net4401));
 sg13g2_buf_8 fanout4402 (.A(net202),
    .X(net4402));
 sg13g2_buf_2 fanout4403 (.A(net4406),
    .X(net4403));
 sg13g2_buf_2 fanout4404 (.A(net4406),
    .X(net4404));
 sg13g2_buf_1 fanout4405 (.A(net4406),
    .X(net4405));
 sg13g2_buf_2 fanout4406 (.A(net4407),
    .X(net4406));
 sg13g2_buf_1 fanout4407 (.A(net4411),
    .X(net4407));
 sg13g2_buf_2 fanout4408 (.A(net4411),
    .X(net4408));
 sg13g2_buf_2 fanout4409 (.A(net4410),
    .X(net4409));
 sg13g2_buf_2 fanout4410 (.A(net4411),
    .X(net4410));
 sg13g2_buf_4 fanout4411 (.X(net4411),
    .A(net4412));
 sg13g2_buf_4 fanout4412 (.X(net4412),
    .A(net4429));
 sg13g2_buf_2 fanout4413 (.A(net4414),
    .X(net4413));
 sg13g2_buf_2 fanout4414 (.A(net4417),
    .X(net4414));
 sg13g2_buf_2 fanout4415 (.A(net4416),
    .X(net4415));
 sg13g2_buf_2 fanout4416 (.A(net4417),
    .X(net4416));
 sg13g2_buf_2 fanout4417 (.A(net4418),
    .X(net4417));
 sg13g2_buf_4 fanout4418 (.X(net4418),
    .A(net4429));
 sg13g2_buf_2 fanout4419 (.A(net4422),
    .X(net4419));
 sg13g2_buf_2 fanout4420 (.A(net4422),
    .X(net4420));
 sg13g2_buf_2 fanout4421 (.A(net4422),
    .X(net4421));
 sg13g2_buf_2 fanout4422 (.A(net4429),
    .X(net4422));
 sg13g2_buf_2 fanout4423 (.A(net4425),
    .X(net4423));
 sg13g2_buf_2 fanout4424 (.A(net4425),
    .X(net4424));
 sg13g2_buf_2 fanout4425 (.A(net4426),
    .X(net4425));
 sg13g2_buf_2 fanout4426 (.A(net4428),
    .X(net4426));
 sg13g2_buf_2 fanout4427 (.A(net4428),
    .X(net4427));
 sg13g2_buf_2 fanout4428 (.A(net4429),
    .X(net4428));
 sg13g2_buf_2 fanout4429 (.A(\cpu.current_instruction[12] ),
    .X(net4429));
 sg13g2_buf_2 fanout4430 (.A(net4431),
    .X(net4430));
 sg13g2_buf_4 fanout4431 (.X(net4431),
    .A(net194));
 sg13g2_buf_4 fanout4432 (.X(net4432),
    .A(net4433));
 sg13g2_buf_4 fanout4433 (.X(net4433),
    .A(net191));
 sg13g2_buf_2 fanout4434 (.A(net4436),
    .X(net4434));
 sg13g2_buf_1 fanout4435 (.A(net4436),
    .X(net4435));
 sg13g2_buf_4 fanout4436 (.X(net4436),
    .A(\cpu.current_instruction[9] ));
 sg13g2_buf_4 fanout4437 (.X(net4437),
    .A(\cpu.current_instruction[9] ));
 sg13g2_buf_2 fanout4438 (.A(\cpu.current_instruction[9] ),
    .X(net4438));
 sg13g2_buf_4 fanout4439 (.X(net4439),
    .A(net4440));
 sg13g2_buf_4 fanout4440 (.X(net4440),
    .A(net207));
 sg13g2_buf_4 fanout4441 (.X(net4441),
    .A(net4442));
 sg13g2_buf_2 fanout4442 (.A(\cpu.current_instruction[8] ),
    .X(net4442));
 sg13g2_buf_4 fanout4443 (.X(net4443),
    .A(net4444));
 sg13g2_buf_4 fanout4444 (.X(net4444),
    .A(net4445));
 sg13g2_buf_2 fanout4445 (.A(net4446),
    .X(net4445));
 sg13g2_buf_4 fanout4446 (.X(net4446),
    .A(net4447));
 sg13g2_buf_4 fanout4447 (.X(net4447),
    .A(net385));
 sg13g2_buf_2 fanout4448 (.A(net4449),
    .X(net4448));
 sg13g2_buf_2 fanout4449 (.A(\cpu.current_instruction[5] ),
    .X(net4449));
 sg13g2_buf_4 fanout4450 (.X(net4450),
    .A(net4451));
 sg13g2_buf_4 fanout4451 (.X(net4451),
    .A(net4452));
 sg13g2_buf_4 fanout4452 (.X(net4452),
    .A(\cpu.current_instruction[4] ));
 sg13g2_buf_4 fanout4453 (.X(net4453),
    .A(net838));
 sg13g2_buf_4 fanout4454 (.X(net4454),
    .A(\cpu.ALU.a[6] ));
 sg13g2_buf_4 fanout4455 (.X(net4455),
    .A(net822));
 sg13g2_buf_1 fanout4456 (.A(\cpu.ALU.a[5] ),
    .X(net4456));
 sg13g2_buf_4 fanout4457 (.X(net4457),
    .A(\cpu.ALU.a[4] ));
 sg13g2_buf_2 fanout4458 (.A(net842),
    .X(net4458));
 sg13g2_buf_4 fanout4459 (.X(net4459),
    .A(\cpu.ALU.a[3] ));
 sg13g2_buf_2 fanout4460 (.A(net883),
    .X(net4460));
 sg13g2_buf_2 fanout4461 (.A(net887),
    .X(net4461));
 sg13g2_buf_2 fanout4462 (.A(\cpu.ALU.a[2] ),
    .X(net4462));
 sg13g2_buf_4 fanout4463 (.X(net4463),
    .A(net849));
 sg13g2_buf_2 fanout4464 (.A(\cpu.ALU.a[1] ),
    .X(net4464));
 sg13g2_buf_4 fanout4465 (.X(net4465),
    .A(net856));
 sg13g2_buf_2 fanout4466 (.A(\cpu.ALU.a[0] ),
    .X(net4466));
 sg13g2_buf_4 fanout4467 (.X(net4467),
    .A(net894));
 sg13g2_buf_4 fanout4468 (.X(net4468),
    .A(net874));
 sg13g2_buf_4 fanout4469 (.X(net4469),
    .A(net889));
 sg13g2_buf_2 fanout4470 (.A(net899),
    .X(net4470));
 sg13g2_buf_2 fanout4471 (.A(net4472),
    .X(net4471));
 sg13g2_buf_4 fanout4472 (.X(net4472),
    .A(net802));
 sg13g2_buf_2 fanout4473 (.A(net4474),
    .X(net4473));
 sg13g2_buf_4 fanout4474 (.X(net4474),
    .A(net865));
 sg13g2_buf_4 fanout4475 (.X(net4475),
    .A(net4477));
 sg13g2_buf_4 fanout4476 (.X(net4476),
    .A(net4477));
 sg13g2_buf_2 fanout4477 (.A(net4481),
    .X(net4477));
 sg13g2_buf_2 fanout4478 (.A(net4480),
    .X(net4478));
 sg13g2_buf_2 fanout4479 (.A(net4480),
    .X(net4479));
 sg13g2_buf_2 fanout4480 (.A(net4481),
    .X(net4480));
 sg13g2_buf_4 fanout4481 (.X(net4481),
    .A(\cpu.set_rx_speed ));
 sg13g2_buf_4 fanout4482 (.X(net4482),
    .A(net936));
 sg13g2_buf_4 fanout4483 (.X(net4483),
    .A(net908));
 sg13g2_buf_4 fanout4484 (.X(net4484),
    .A(net895));
 sg13g2_buf_4 fanout4485 (.X(net4485),
    .A(\cpu.keccak_alu.registers[182] ));
 sg13g2_buf_4 fanout4486 (.X(net4486),
    .A(\cpu.keccak_alu.registers[181] ));
 sg13g2_buf_4 fanout4487 (.X(net4487),
    .A(\cpu.keccak_alu.registers[180] ));
 sg13g2_buf_4 fanout4488 (.X(net4488),
    .A(net931));
 sg13g2_buf_4 fanout4489 (.X(net4489),
    .A(\cpu.keccak_alu.registers[172] ));
 sg13g2_buf_2 fanout4490 (.A(net909),
    .X(net4490));
 sg13g2_buf_2 fanout4491 (.A(\cpu.keccak_alu.registers[171] ),
    .X(net4491));
 sg13g2_buf_4 fanout4492 (.X(net4492),
    .A(net898));
 sg13g2_buf_4 fanout4493 (.X(net4493),
    .A(\cpu.keccak_alu.registers[165] ));
 sg13g2_buf_4 fanout4494 (.X(net4494),
    .A(net941));
 sg13g2_buf_4 fanout4495 (.X(net4495),
    .A(\cpu.keccak_alu.registers[163] ));
 sg13g2_buf_4 fanout4496 (.X(net4496),
    .A(\cpu.keccak_alu.registers[161] ));
 sg13g2_buf_4 fanout4497 (.X(net4497),
    .A(\cpu.keccak_alu.registers[160] ));
 sg13g2_buf_4 fanout4498 (.X(net4498),
    .A(net943));
 sg13g2_buf_4 fanout4499 (.X(net4499),
    .A(net876));
 sg13g2_buf_4 fanout4500 (.X(net4500),
    .A(net917));
 sg13g2_buf_4 fanout4501 (.X(net4501),
    .A(net945));
 sg13g2_buf_4 fanout4502 (.X(net4502),
    .A(net905));
 sg13g2_buf_4 fanout4503 (.X(net4503),
    .A(net739));
 sg13g2_buf_4 fanout4504 (.X(net4504),
    .A(net896));
 sg13g2_buf_4 fanout4505 (.X(net4505),
    .A(\cpu.keccak_alu.registers[142] ));
 sg13g2_buf_4 fanout4506 (.X(net4506),
    .A(net902));
 sg13g2_buf_4 fanout4507 (.X(net4507),
    .A(net829));
 sg13g2_buf_2 fanout4508 (.A(\cpu.keccak_alu.registers[140] ),
    .X(net4508));
 sg13g2_buf_4 fanout4509 (.X(net4509),
    .A(net927));
 sg13g2_buf_2 fanout4510 (.A(net873),
    .X(net4510));
 sg13g2_buf_2 fanout4511 (.A(\cpu.keccak_alu.registers[136] ),
    .X(net4511));
 sg13g2_buf_2 fanout4512 (.A(\cpu.keccak_alu.registers[135] ),
    .X(net4512));
 sg13g2_buf_2 fanout4513 (.A(net4516),
    .X(net4513));
 sg13g2_buf_2 fanout4514 (.A(net4516),
    .X(net4514));
 sg13g2_buf_4 fanout4515 (.X(net4515),
    .A(net4516));
 sg13g2_buf_2 fanout4516 (.A(\cpu.keccak_alu.registers[134] ),
    .X(net4516));
 sg13g2_buf_2 fanout4517 (.A(net4518),
    .X(net4517));
 sg13g2_buf_2 fanout4518 (.A(\cpu.keccak_alu.registers[133] ),
    .X(net4518));
 sg13g2_buf_2 fanout4519 (.A(net4520),
    .X(net4519));
 sg13g2_buf_2 fanout4520 (.A(\cpu.keccak_alu.registers[133] ),
    .X(net4520));
 sg13g2_buf_4 fanout4521 (.X(net4521),
    .A(\cpu.keccak_alu.registers[132] ));
 sg13g2_buf_1 fanout4522 (.A(net914),
    .X(net4522));
 sg13g2_buf_2 fanout4523 (.A(net4524),
    .X(net4523));
 sg13g2_buf_1 fanout4524 (.A(\cpu.keccak_alu.registers[132] ),
    .X(net4524));
 sg13g2_buf_2 fanout4525 (.A(net4526),
    .X(net4525));
 sg13g2_buf_2 fanout4526 (.A(net4527),
    .X(net4526));
 sg13g2_buf_4 fanout4527 (.X(net4527),
    .A(\cpu.keccak_alu.registers[131] ));
 sg13g2_buf_4 fanout4528 (.X(net4528),
    .A(net4529));
 sg13g2_buf_1 fanout4529 (.A(net4530),
    .X(net4529));
 sg13g2_buf_4 fanout4530 (.X(net4530),
    .A(net870));
 sg13g2_buf_4 fanout4531 (.X(net4531),
    .A(net4534));
 sg13g2_buf_2 fanout4532 (.A(net4533),
    .X(net4532));
 sg13g2_buf_2 fanout4533 (.A(net4534),
    .X(net4533));
 sg13g2_buf_2 fanout4534 (.A(\cpu.keccak_alu.registers[130] ),
    .X(net4534));
 sg13g2_buf_2 fanout4535 (.A(net4536),
    .X(net4535));
 sg13g2_buf_2 fanout4536 (.A(net4537),
    .X(net4536));
 sg13g2_buf_4 fanout4537 (.X(net4537),
    .A(\cpu.keccak_alu.registers[129] ));
 sg13g2_buf_2 fanout4538 (.A(net4540),
    .X(net4538));
 sg13g2_buf_1 fanout4539 (.A(net4540),
    .X(net4539));
 sg13g2_buf_2 fanout4540 (.A(\cpu.keccak_alu.registers[129] ),
    .X(net4540));
 sg13g2_buf_2 fanout4541 (.A(net4543),
    .X(net4541));
 sg13g2_buf_2 fanout4542 (.A(net4543),
    .X(net4542));
 sg13g2_buf_1 fanout4543 (.A(net4547),
    .X(net4543));
 sg13g2_buf_2 fanout4544 (.A(net4546),
    .X(net4544));
 sg13g2_buf_1 fanout4545 (.A(net4546),
    .X(net4545));
 sg13g2_buf_4 fanout4546 (.X(net4546),
    .A(net4547));
 sg13g2_buf_2 fanout4547 (.A(net939),
    .X(net4547));
 sg13g2_buf_2 fanout4548 (.A(net4549),
    .X(net4548));
 sg13g2_buf_2 fanout4549 (.A(net4550),
    .X(net4549));
 sg13g2_buf_2 fanout4550 (.A(net4551),
    .X(net4550));
 sg13g2_buf_2 fanout4551 (.A(net4555),
    .X(net4551));
 sg13g2_buf_2 fanout4552 (.A(net4553),
    .X(net4552));
 sg13g2_buf_2 fanout4553 (.A(net4555),
    .X(net4553));
 sg13g2_buf_2 fanout4554 (.A(net4555),
    .X(net4554));
 sg13g2_buf_1 fanout4555 (.A(net4575),
    .X(net4555));
 sg13g2_buf_2 fanout4556 (.A(net4557),
    .X(net4556));
 sg13g2_buf_2 fanout4557 (.A(net4561),
    .X(net4557));
 sg13g2_buf_2 fanout4558 (.A(net4559),
    .X(net4558));
 sg13g2_buf_2 fanout4559 (.A(net4560),
    .X(net4559));
 sg13g2_buf_2 fanout4560 (.A(net4561),
    .X(net4560));
 sg13g2_buf_2 fanout4561 (.A(net4575),
    .X(net4561));
 sg13g2_buf_2 fanout4562 (.A(net4566),
    .X(net4562));
 sg13g2_buf_1 fanout4563 (.A(net4566),
    .X(net4563));
 sg13g2_buf_2 fanout4564 (.A(net4565),
    .X(net4564));
 sg13g2_buf_2 fanout4565 (.A(net4566),
    .X(net4565));
 sg13g2_buf_2 fanout4566 (.A(net4567),
    .X(net4566));
 sg13g2_buf_2 fanout4567 (.A(net4575),
    .X(net4567));
 sg13g2_buf_2 fanout4568 (.A(net4573),
    .X(net4568));
 sg13g2_buf_2 fanout4569 (.A(net4570),
    .X(net4569));
 sg13g2_buf_1 fanout4570 (.A(net4571),
    .X(net4570));
 sg13g2_buf_1 fanout4571 (.A(net4572),
    .X(net4571));
 sg13g2_buf_2 fanout4572 (.A(net4573),
    .X(net4572));
 sg13g2_buf_2 fanout4573 (.A(net4574),
    .X(net4573));
 sg13g2_buf_2 fanout4574 (.A(net4575),
    .X(net4574));
 sg13g2_buf_4 fanout4575 (.X(net4575),
    .A(\cpu.keccak_alu.registers[128] ));
 sg13g2_buf_4 fanout4576 (.X(net4576),
    .A(_00129_));
 sg13g2_buf_2 fanout4577 (.A(net4579),
    .X(net4577));
 sg13g2_buf_2 fanout4578 (.A(net4579),
    .X(net4578));
 sg13g2_buf_1 fanout4579 (.A(net4580),
    .X(net4579));
 sg13g2_buf_2 fanout4580 (.A(net4581),
    .X(net4580));
 sg13g2_buf_2 fanout4581 (.A(\cpu.reset ),
    .X(net4581));
 sg13g2_buf_2 fanout4582 (.A(\cpu.reset ),
    .X(net4582));
 sg13g2_buf_1 fanout4583 (.A(net4584),
    .X(net4583));
 sg13g2_buf_2 fanout4584 (.A(net4585),
    .X(net4584));
 sg13g2_buf_2 fanout4585 (.A(\cpu.reset ),
    .X(net4585));
 sg13g2_buf_4 fanout4586 (.X(net4586),
    .A(net4590));
 sg13g2_buf_4 fanout4587 (.X(net4587),
    .A(net4590));
 sg13g2_buf_4 fanout4588 (.X(net4588),
    .A(net4590));
 sg13g2_buf_4 fanout4589 (.X(net4589),
    .A(net4590));
 sg13g2_buf_2 fanout4590 (.A(net4619),
    .X(net4590));
 sg13g2_buf_4 fanout4591 (.X(net4591),
    .A(net4594));
 sg13g2_buf_4 fanout4592 (.X(net4592),
    .A(net4594));
 sg13g2_buf_4 fanout4593 (.X(net4593),
    .A(net4594));
 sg13g2_buf_4 fanout4594 (.X(net4594),
    .A(net4619));
 sg13g2_buf_4 fanout4595 (.X(net4595),
    .A(net4597));
 sg13g2_buf_2 fanout4596 (.A(net4597),
    .X(net4596));
 sg13g2_buf_4 fanout4597 (.X(net4597),
    .A(net4603));
 sg13g2_buf_4 fanout4598 (.X(net4598),
    .A(net4600));
 sg13g2_buf_4 fanout4599 (.X(net4599),
    .A(net4600));
 sg13g2_buf_2 fanout4600 (.A(net4603),
    .X(net4600));
 sg13g2_buf_4 fanout4601 (.X(net4601),
    .A(net4603));
 sg13g2_buf_4 fanout4602 (.X(net4602),
    .A(net4603));
 sg13g2_buf_2 fanout4603 (.A(net4619),
    .X(net4603));
 sg13g2_buf_4 fanout4604 (.X(net4604),
    .A(net4605));
 sg13g2_buf_4 fanout4605 (.X(net4605),
    .A(net4606));
 sg13g2_buf_4 fanout4606 (.X(net4606),
    .A(net4610));
 sg13g2_buf_4 fanout4607 (.X(net4607),
    .A(net4609));
 sg13g2_buf_2 fanout4608 (.A(net4609),
    .X(net4608));
 sg13g2_buf_4 fanout4609 (.X(net4609),
    .A(net4610));
 sg13g2_buf_2 fanout4610 (.A(net4619),
    .X(net4610));
 sg13g2_buf_4 fanout4611 (.X(net4611),
    .A(net4614));
 sg13g2_buf_4 fanout4612 (.X(net4612),
    .A(net4614));
 sg13g2_buf_4 fanout4613 (.X(net4613),
    .A(net4614));
 sg13g2_buf_2 fanout4614 (.A(net4619),
    .X(net4614));
 sg13g2_buf_4 fanout4615 (.X(net4615),
    .A(net4618));
 sg13g2_buf_4 fanout4616 (.X(net4616),
    .A(net4617));
 sg13g2_buf_4 fanout4617 (.X(net4617),
    .A(net4618));
 sg13g2_buf_2 fanout4618 (.A(net4619),
    .X(net4618));
 sg13g2_buf_4 fanout4619 (.X(net4619),
    .A(net4701));
 sg13g2_buf_4 fanout4620 (.X(net4620),
    .A(net4623));
 sg13g2_buf_4 fanout4621 (.X(net4621),
    .A(net4623));
 sg13g2_buf_2 fanout4622 (.A(net4623),
    .X(net4622));
 sg13g2_buf_4 fanout4623 (.X(net4623),
    .A(net4653));
 sg13g2_buf_4 fanout4624 (.X(net4624),
    .A(net4626));
 sg13g2_buf_4 fanout4625 (.X(net4625),
    .A(net4626));
 sg13g2_buf_4 fanout4626 (.X(net4626),
    .A(net4653));
 sg13g2_buf_4 fanout4627 (.X(net4627),
    .A(net4636));
 sg13g2_buf_4 fanout4628 (.X(net4628),
    .A(net4636));
 sg13g2_buf_4 fanout4629 (.X(net4629),
    .A(net4630));
 sg13g2_buf_4 fanout4630 (.X(net4630),
    .A(net4636));
 sg13g2_buf_4 fanout4631 (.X(net4631),
    .A(net4635));
 sg13g2_buf_4 fanout4632 (.X(net4632),
    .A(net4635));
 sg13g2_buf_4 fanout4633 (.X(net4633),
    .A(net4634));
 sg13g2_buf_4 fanout4634 (.X(net4634),
    .A(net4635));
 sg13g2_buf_2 fanout4635 (.A(net4636),
    .X(net4635));
 sg13g2_buf_2 fanout4636 (.A(net4653),
    .X(net4636));
 sg13g2_buf_4 fanout4637 (.X(net4637),
    .A(net4639));
 sg13g2_buf_4 fanout4638 (.X(net4638),
    .A(net4639));
 sg13g2_buf_4 fanout4639 (.X(net4639),
    .A(net4652));
 sg13g2_buf_4 fanout4640 (.X(net4640),
    .A(net4642));
 sg13g2_buf_2 fanout4641 (.A(net4642),
    .X(net4641));
 sg13g2_buf_4 fanout4642 (.X(net4642),
    .A(net4652));
 sg13g2_buf_4 fanout4643 (.X(net4643),
    .A(net4644));
 sg13g2_buf_4 fanout4644 (.X(net4644),
    .A(net4647));
 sg13g2_buf_4 fanout4645 (.X(net4645),
    .A(net4646));
 sg13g2_buf_4 fanout4646 (.X(net4646),
    .A(net4647));
 sg13g2_buf_2 fanout4647 (.A(net4651),
    .X(net4647));
 sg13g2_buf_4 fanout4648 (.X(net4648),
    .A(net4651));
 sg13g2_buf_4 fanout4649 (.X(net4649),
    .A(net4650));
 sg13g2_buf_2 fanout4650 (.A(net4651),
    .X(net4650));
 sg13g2_buf_2 fanout4651 (.A(net4652),
    .X(net4651));
 sg13g2_buf_2 fanout4652 (.A(net4653),
    .X(net4652));
 sg13g2_buf_2 fanout4653 (.A(net4701),
    .X(net4653));
 sg13g2_buf_4 fanout4654 (.X(net4654),
    .A(net4655));
 sg13g2_buf_4 fanout4655 (.X(net4655),
    .A(net4662));
 sg13g2_buf_4 fanout4656 (.X(net4656),
    .A(net4662));
 sg13g2_buf_4 fanout4657 (.X(net4657),
    .A(net4662));
 sg13g2_buf_4 fanout4658 (.X(net4658),
    .A(net4661));
 sg13g2_buf_2 fanout4659 (.A(net4661),
    .X(net4659));
 sg13g2_buf_4 fanout4660 (.X(net4660),
    .A(net4661));
 sg13g2_buf_2 fanout4661 (.A(net4662),
    .X(net4661));
 sg13g2_buf_2 fanout4662 (.A(net4675),
    .X(net4662));
 sg13g2_buf_4 fanout4663 (.X(net4663),
    .A(net4674));
 sg13g2_buf_2 fanout4664 (.A(net4674),
    .X(net4664));
 sg13g2_buf_4 fanout4665 (.X(net4665),
    .A(net4666));
 sg13g2_buf_4 fanout4666 (.X(net4666),
    .A(net4673));
 sg13g2_buf_4 fanout4667 (.X(net4667),
    .A(net4673));
 sg13g2_buf_2 fanout4668 (.A(net4673),
    .X(net4668));
 sg13g2_buf_8 fanout4669 (.A(net4673),
    .X(net4669));
 sg13g2_buf_4 fanout4670 (.X(net4670),
    .A(net4673));
 sg13g2_buf_4 fanout4671 (.X(net4671),
    .A(net4672));
 sg13g2_buf_4 fanout4672 (.X(net4672),
    .A(net4673));
 sg13g2_buf_4 fanout4673 (.X(net4673),
    .A(net4674));
 sg13g2_buf_2 fanout4674 (.A(net4675),
    .X(net4674));
 sg13g2_buf_2 fanout4675 (.A(net4701),
    .X(net4675));
 sg13g2_buf_4 fanout4676 (.X(net4676),
    .A(net4678));
 sg13g2_buf_2 fanout4677 (.A(net4678),
    .X(net4677));
 sg13g2_buf_4 fanout4678 (.X(net4678),
    .A(net4683));
 sg13g2_buf_4 fanout4679 (.X(net4679),
    .A(net4682));
 sg13g2_buf_4 fanout4680 (.X(net4680),
    .A(net4681));
 sg13g2_buf_4 fanout4681 (.X(net4681),
    .A(net4682));
 sg13g2_buf_2 fanout4682 (.A(net4683),
    .X(net4682));
 sg13g2_buf_2 fanout4683 (.A(net4700),
    .X(net4683));
 sg13g2_buf_4 fanout4684 (.X(net4684),
    .A(net4686));
 sg13g2_buf_2 fanout4685 (.A(net4686),
    .X(net4685));
 sg13g2_buf_2 fanout4686 (.A(net4700),
    .X(net4686));
 sg13g2_buf_4 fanout4687 (.X(net4687),
    .A(net4688));
 sg13g2_buf_2 fanout4688 (.A(net4700),
    .X(net4688));
 sg13g2_buf_4 fanout4689 (.X(net4689),
    .A(net4693));
 sg13g2_buf_4 fanout4690 (.X(net4690),
    .A(net4693));
 sg13g2_buf_4 fanout4691 (.X(net4691),
    .A(net4692));
 sg13g2_buf_4 fanout4692 (.X(net4692),
    .A(net4693));
 sg13g2_buf_2 fanout4693 (.A(net4699),
    .X(net4693));
 sg13g2_buf_4 fanout4694 (.X(net4694),
    .A(net4695));
 sg13g2_buf_2 fanout4695 (.A(net4699),
    .X(net4695));
 sg13g2_buf_4 fanout4696 (.X(net4696),
    .A(net4698));
 sg13g2_buf_2 fanout4697 (.A(net4698),
    .X(net4697));
 sg13g2_buf_4 fanout4698 (.X(net4698),
    .A(net4699));
 sg13g2_buf_2 fanout4699 (.A(net4700),
    .X(net4699));
 sg13g2_buf_2 fanout4700 (.A(net4701),
    .X(net4700));
 sg13g2_buf_4 fanout4701 (.X(net4701),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(uio_in[0]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(uio_in[1]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[2]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[3]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[4]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[5]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[6]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[7]),
    .X(net11));
 sg13g2_tielo tt_um_zoom_zoom_12 (.L_LO(net12));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_leaf_91_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_2 clkbuf_leaf_92_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_2 clkbuf_leaf_93_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_2 clkbuf_leaf_94_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_2 clkbuf_leaf_95_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_2 clkbuf_leaf_96_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_4_8_0_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_4_9_0_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_4_10_0_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_buf_2 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_buf_2 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_buf_2 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_92_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_4_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_91_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_9_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_11_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_84_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_85_clk));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_18_clk));
 sg13g2_inv_4 clkload23 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_38_clk));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_12_clk));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_43_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_77_clk));
 sg13g2_inv_4 clkload29 (.A(clknet_leaf_39_clk));
 sg13g2_inv_4 clkload30 (.A(clknet_leaf_42_clk));
 sg13g2_inv_4 clkload31 (.A(clknet_leaf_44_clk));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_64_clk));
 sg13g2_inv_4 clkload33 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload34 (.A(clknet_leaf_46_clk));
 sg13g2_inv_4 clkload35 (.A(clknet_leaf_60_clk));
 sg13g2_inv_4 clkload36 (.A(clknet_leaf_51_clk));
 sg13g2_inv_8 clkload37 (.A(clknet_leaf_53_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\memory_controller.next_state[1] ),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold2 (.A(\memory_controller.next_state[3] ),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold3 (.A(\memory_controller.next_state[0] ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold4 (.A(\memory_controller.next_state[2] ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold5 (.A(\memory_controller.next_state[4] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold6 (.A(_00245_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold7 (.A(_00878_),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold8 (.A(_00248_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold9 (.A(_00870_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold10 (.A(_00249_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold11 (.A(_00868_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cpu.uart.stage[0] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold13 (.A(_00262_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold14 (.A(_00246_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold15 (.A(_00873_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold16 (.A(_00259_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold17 (.A(_06568_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold18 (.A(_00880_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold19 (.A(_00247_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold20 (.A(_00872_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold21 (.A(_00244_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold22 (.A(_00879_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold23 (.A(\cpu.rx_speed[12] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold24 (.A(\uart_receiver/_083_ ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold25 (.A(\uart_receiver/_006_ ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold26 (.A(\uart_receiver/_074_ ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cpu.execution_stage[0] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold28 (.A(_00261_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cpu.registers[7][3] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold30 (.A(\uart_receiver/_007_ ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold31 (.A(\uart_receiver/_076_ ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cpu.registers[7][1] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold33 (.A(_00839_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cpu.memory_in[2] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cpu.memory_in[9] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold36 (.A(\cpu.memory_in[4] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold37 (.A(\memory_controller.wait_counter[0] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold38 (.A(\cpu.registers[7][2] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold39 (.A(\uart_receiver/_005_ ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold40 (.A(\uart_receiver/_071_ ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold41 (.A(\uart_receiver/_009_ ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold42 (.A(\uart_receiver/_082_ ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cpu.memory_in[8] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold44 (.A(\uart_receiver/_008_ ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold45 (.A(\uart_receiver/_077_ ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold46 (.A(\cpu.memory_in[11] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cpu.memory_in[5] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold48 (.A(_06292_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold49 (.A(\cpu.memory_in[3] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cpu.ALU.mode[2] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold51 (.A(_00618_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cpu.data_out[12] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold53 (.A(\cpu.memory_in[10] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cpu.data_out[5] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cpu.memory_in[0] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cpu.data_out[10] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold57 (.A(\cpu.memory_in[1] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cpu.data_out[15] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold59 (.A(_00666_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold60 (.A(\cpu.memory_in[13] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold61 (.A(\cpu.memory_in[6] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold62 (.A(\cpu.request ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold63 (.A(_06433_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold64 (.A(\uart_receiver/data[1] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold65 (.A(\uart_receiver/_098_ ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold66 (.A(\cpu.registers[7][8] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold67 (.A(\uart_receiver/data[6] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold68 (.A(\uart_receiver/_103_ ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold69 (.A(\cpu.data_out[11] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold70 (.A(_00662_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cpu.registers[7][10] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold72 (.A(\cpu.registers[7][5] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cpu.memory_in[7] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold74 (.A(\cpu.memory_in[15] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cpu.registers[7][6] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold76 (.A(\cpu.keccak_alu.registers[273] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold77 (.A(\cpu.registers[7][7] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cpu.registers[7][9] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold79 (.A(\cpu.data_out[4] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold80 (.A(\uart_receiver/data[5] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold81 (.A(\uart_receiver/_102_ ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cpu.registers[7][4] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cpu.keccak_alu.registers[276] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold84 (.A(\uart_receiver/data[3] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold85 (.A(\uart_receiver/_100_ ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold86 (.A(\cpu.registers[7][13] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold87 (.A(\cpu.data_out[13] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold88 (.A(\cpu.registers[7][11] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cpu.data_out[14] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cpu.keccak_alu.registers[291] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cpu.registers[7][12] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cpu.data_out[9] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cpu.data_out[2] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold94 (.A(_00653_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cpu.uart.cycle_counter[7] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold96 (.A(_06555_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold97 (.A(_00861_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cpu.keccak_alu.registers[275] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cpu.uart.cycle_counter[3] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold100 (.A(_06549_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold101 (.A(_00857_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cpu.memory_in[12] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cpu.current_instruction[5] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cpu.keccak_alu.registers[317] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cpu.keccak_alu.registers[181] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold106 (.A(_00509_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cpu.keccak_alu.registers[296] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cpu.registers[7][15] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cpu.rx_speed[11] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cpu.keccak_alu.registers[314] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cpu.keccak_alu.registers[298] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cpu.current_address[9] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold113 (.A(_00644_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cpu.keccak_alu.registers[306] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cpu.registers[7][14] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold116 (.A(lower_bit),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cpu.ALU.b[14] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cpu.current_address[4] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold119 (.A(_00639_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cpu.keccak_alu.registers[302] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold121 (.A(\data_received[1] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cpu.current_address[14] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold123 (.A(_00649_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cpu.current_address[6] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold125 (.A(_00641_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cpu.keccak_alu.registers[299] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold127 (.A(\cpu.current_address[3] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold128 (.A(_00638_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold129 (.A(\uart_receiver/data[4] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold130 (.A(\uart_receiver/_181_ ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold131 (.A(\uart_receiver/_101_ ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold132 (.A(\uart_receiver/data[2] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold133 (.A(\data_received[6] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cpu.keccak_alu.registers[315] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold135 (.A(\cpu.keccak_alu.registers[288] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold136 (.A(\uart_receiver/data[7] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold137 (.A(\uart_receiver/_070_ ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold138 (.A(\cpu.keccak_alu.registers[263] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cpu.keccak_alu.registers[312] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cpu.current_address[5] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold141 (.A(_00640_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cpu.registers[6][1] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold143 (.A(_00702_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cpu.registers[6][2] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold145 (.A(_00703_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cpu.keccak_alu.registers[309] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold147 (.A(\cpu.keccak_alu.registers[285] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold148 (.A(\cpu.keccak_alu.registers[318] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cpu.keccak_alu.registers[294] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold150 (.A(\memory_controller.wait_counter[2] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold151 (.A(_01327_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold152 (.A(_00012_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cpu.keccak_alu.registers[305] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cpu.keccak_alu.registers[304] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cpu.keccak_alu.registers[311] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold156 (.A(\memory_controller.wait_counter[2] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold157 (.A(_06414_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold158 (.A(\uart_receiver/data[0] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold159 (.A(\uart_receiver/_097_ ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold160 (.A(\cpu.keccak_alu.registers[18] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold161 (.A(\cpu.registers[1][3] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cpu.keccak_alu.registers[307] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cpu.keccak_alu.registers[261] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cpu.uart_inbound ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold165 (.A(\uart_receiver/stage[2] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cpu.uart.cycles_per_bit[0] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold167 (.A(_00867_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold168 (.A(\cpu.data_out[6] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cpu.uart.cycles_per_bit[4] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold170 (.A(_00871_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold171 (.A(\cpu.keccak_alu.registers[316] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold172 (.A(\data_received[3] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cpu.current_instruction[10] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold174 (.A(\memory_controller.uart_memory_address[10] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cpu.keccak_alu.registers[290] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold176 (.A(\cpu.current_instruction[11] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold177 (.A(\cpu.keccak_alu.registers[310] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cpu.keccak_alu.registers[287] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold179 (.A(\data_received[2] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cpu.uart.cycles_per_bit[2] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold181 (.A(_00869_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cpu.registers[4][2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold183 (.A(_00265_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold184 (.A(\cpu.current_instruction[13] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold185 (.A(\cpu.current_instruction[0] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold186 (.A(\cpu.jump_con ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold187 (.A(_00314_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold188 (.A(\data_received[5] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold189 (.A(\cpu.current_instruction[8] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold190 (.A(\cpu.current_instruction[3] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold191 (.A(\cpu.keccak_alu.registers[297] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold192 (.A(\cpu.keccak_alu.registers[289] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cpu.request_type ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold194 (.A(\cpu.uart.data_sending[7] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold195 (.A(_00812_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold196 (.A(\cpu.uart.data_sending[4] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold197 (.A(_00809_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cpu.data_out[8] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold199 (.A(_00659_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold200 (.A(\cpu.keccak_alu.registers[293] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold201 (.A(\cpu.registers[6][3] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold202 (.A(_00704_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold203 (.A(\cpu.keccak_alu.registers[277] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold204 (.A(\cpu.registers[4][9] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold205 (.A(_00272_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold206 (.A(\cpu.registers[4][1] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold207 (.A(_00264_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold208 (.A(\cpu.keccak_alu.registers[72] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold209 (.A(\cpu.registers[1][9] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold210 (.A(_00817_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold211 (.A(\cpu.uart.cycles_per_bit[8] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold212 (.A(_00875_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold213 (.A(\cpu.keccak_alu.registers[274] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold214 (.A(\cpu.keccak_alu.registers[73] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold215 (.A(\cpu.uart.data_sending[3] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold216 (.A(_00808_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold217 (.A(\cpu.current_address[8] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold218 (.A(_00643_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold219 (.A(\cpu.keccak_alu.registers[313] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold220 (.A(\cpu.current_instruction[2] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold221 (.A(\cpu.registers[1][5] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold222 (.A(_00813_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold223 (.A(\cpu.memory_in[14] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold224 (.A(\cpu.rx_speed[5] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold225 (.A(\cpu.registers[6][9] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold226 (.A(_00710_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold227 (.A(\cpu.uart.data_sending[2] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold228 (.A(_00807_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold229 (.A(\cpu.keccak_alu.registers[172] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold230 (.A(\cpu.rx_speed[9] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold231 (.A(_00324_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold232 (.A(\cpu.registers[4][6] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold233 (.A(\cpu.keccak_alu.registers[262] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold234 (.A(\cpu.uart.data_sending[1] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold235 (.A(_00806_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold236 (.A(\cpu.keccak_alu.registers[272] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold237 (.A(\cpu.registers[1][6] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold238 (.A(_00814_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold239 (.A(\cpu.keccak_alu.registers[91] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold240 (.A(\cpu.uart.data_sending[0] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold241 (.A(_00805_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold242 (.A(\cpu.keccak_alu.registers[193] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold243 (.A(\cpu.keccak_alu.registers[90] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold244 (.A(\cpu.keccak_alu.registers[78] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold245 (.A(_00406_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold246 (.A(\cpu.uart.cycle_counter[1] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold247 (.A(_06545_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold248 (.A(_00855_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold249 (.A(\cpu.keccak_alu.registers[256] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold250 (.A(\cpu.current_instruction[1] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold251 (.A(\cpu.keccak_alu.registers[301] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold252 (.A(\cpu.rx_speed[8] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold253 (.A(\cpu.registers[4][3] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold254 (.A(_00266_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold255 (.A(\cpu.keccak_alu.registers[229] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold256 (.A(\cpu.registers[4][7] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold257 (.A(_00270_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold258 (.A(\cpu.keccak_alu.registers[295] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold259 (.A(\cpu.keccak_alu.registers[270] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold260 (.A(\cpu.uart.cycle_counter[9] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold261 (.A(_06558_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold262 (.A(_00863_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold263 (.A(\cpu.keccak_alu.registers[215] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold264 (.A(\cpu.keccak_alu.registers[258] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold265 (.A(\cpu.keccak_alu.registers[267] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold266 (.A(\cpu.registers[1][14] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold267 (.A(_00822_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold268 (.A(\cpu.registers[1][11] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold269 (.A(_00819_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold270 (.A(\cpu.uart.cycles_per_bit[7] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold271 (.A(_00874_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold272 (.A(\cpu.registers[1][7] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold273 (.A(_00815_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold274 (.A(\cpu.registers[4][5] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold275 (.A(_00268_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold276 (.A(\cpu.registers[4][12] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold277 (.A(_00275_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold278 (.A(\cpu.keccak_alu.registers[303] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold279 (.A(\cpu.keccak_alu.registers[77] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold280 (.A(\cpu.registers[6][4] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold281 (.A(_00705_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold282 (.A(\cpu.keccak_alu.registers[210] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold283 (.A(\cpu.keccak_alu.registers[88] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold284 (.A(\cpu.registers[1][10] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold285 (.A(_00818_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold286 (.A(\cpu.keccak_alu.registers[95] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold287 (.A(\cpu.uart.data_sending[5] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold288 (.A(\cpu.data_out[7] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold289 (.A(_00658_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold290 (.A(\cpu.registers[6][0] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold291 (.A(_00701_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold292 (.A(\cpu.keccak_alu.registers[265] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold293 (.A(\cpu.rx_speed[1] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold294 (.A(\cpu.registers[4][10] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold295 (.A(_00273_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold296 (.A(_00019_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold297 (.A(_00793_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold298 (.A(\cpu.keccak_alu.registers[239] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold299 (.A(\cpu.current_address[12] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold300 (.A(_00647_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold301 (.A(\cpu.current_address[11] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold302 (.A(_00646_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold303 (.A(\cpu.registers[2][2] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold304 (.A(_00297_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold305 (.A(\cpu.keccak_alu.registers[199] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold306 (.A(\cpu.current_address[13] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold307 (.A(_00648_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold308 (.A(\cpu.registers[2][15] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold309 (.A(_00310_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold310 (.A(\cpu.keccak_alu.registers[225] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold311 (.A(\cpu.registers[4][14] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold312 (.A(_00277_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold313 (.A(\cpu.keccak_alu.registers[1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold314 (.A(\cpu.keccak_alu.registers[308] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold315 (.A(\cpu.keccak_alu.registers[74] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold316 (.A(\cpu.registers[6][8] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold317 (.A(_00709_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold318 (.A(\cpu.registers[6][12] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold319 (.A(_00713_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold320 (.A(\cpu.keccak_alu.registers[266] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold321 (.A(\data_received[0] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold322 (.A(\cpu.registers[4][11] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold323 (.A(_00274_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold324 (.A(\cpu.uart.busy ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold325 (.A(_00008_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold326 (.A(\cpu.uart.data_sending[6] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold327 (.A(_00811_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold328 (.A(\cpu.keccak_alu.registers[280] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold329 (.A(\cpu.registers[7][0] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold330 (.A(_00838_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold331 (.A(\cpu.keccak_alu.registers[226] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold332 (.A(\cpu.registers[1][4] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold333 (.A(\cpu.current_instruction[6] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold334 (.A(\cpu.uart.cycles_per_bit[9] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold335 (.A(\cpu.registers[1][8] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold336 (.A(_00816_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold337 (.A(\cpu.current_address[10] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold338 (.A(_00645_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold339 (.A(\cpu.request_address[15] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold340 (.A(\cpu.keccak_alu.registers[247] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold341 (.A(\cpu.keccak_alu.registers[217] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold342 (.A(\cpu.registers[3][4] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold343 (.A(_00283_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold344 (.A(\cpu.registers[1][13] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold345 (.A(_00821_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold346 (.A(\cpu.registers[6][5] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold347 (.A(_00706_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold348 (.A(\cpu.registers[6][11] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold349 (.A(_00712_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold350 (.A(\cpu.uart.cycle_counter[10] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold351 (.A(_06560_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold352 (.A(\cpu.registers[1][12] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold353 (.A(_00820_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold354 (.A(\cpu.registers[6][7] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold355 (.A(_00708_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold356 (.A(\data_received[4] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold357 (.A(\cpu.keccak_alu.registers[230] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold358 (.A(\cpu.uart.cycles_per_bit[10] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold359 (.A(_00877_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold360 (.A(\cpu.uart.cycle_counter[11] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold361 (.A(\memory_controller.wait_counter[3] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold362 (.A(_01329_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold363 (.A(\memory_controller.write_enable ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold364 (.A(_00783_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold365 (.A(\cpu.keccak_alu.registers[202] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold366 (.A(\cpu.keccak_alu.registers[194] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold367 (.A(\cpu.current_instruction[7] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold368 (.A(\cpu.keccak_alu.registers[269] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold369 (.A(\cpu.keccak_alu.registers[208] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold370 (.A(_00536_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold371 (.A(\cpu.keccak_alu.registers[257] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold372 (.A(\cpu.keccak_alu.registers[292] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold373 (.A(\cpu.uart.cycle_counter[0] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold374 (.A(_00854_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold375 (.A(\cpu.data_out[1] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold376 (.A(_00652_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold377 (.A(\cpu.keccak_alu.registers[34] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold378 (.A(\cpu.registers[4][13] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold379 (.A(_00276_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold380 (.A(\cpu.execution_stage[3] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold381 (.A(\cpu.registers[4][15] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold382 (.A(_00278_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold383 (.A(\cpu.keccak_alu.registers[237] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold384 (.A(\cpu.registers[4][8] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold385 (.A(_00271_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold386 (.A(\cpu.keccak_alu.registers[253] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold387 (.A(\cpu.rx_speed[6] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold388 (.A(\cpu.registers[6][13] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold389 (.A(_00714_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold390 (.A(\cpu.keccak_alu.registers[93] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold391 (.A(\cpu.rx_speed[10] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold392 (.A(\cpu.registers[4][4] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold393 (.A(\cpu.keccak_alu.registers[252] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold394 (.A(\cpu.keccak_alu.registers[192] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold395 (.A(_00520_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold396 (.A(\cpu.keccak_alu.registers[227] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold397 (.A(\cpu.keccak_alu.registers[212] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold398 (.A(\cpu.keccak_alu.registers[5] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold399 (.A(\cpu.keccak_alu.registers[200] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold400 (.A(\cpu.registers[4][0] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold401 (.A(_00263_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold402 (.A(\cpu.keccak_alu.registers[224] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold403 (.A(\cpu.keccak_alu.registers[82] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold404 (.A(\cpu.registers[5][1] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold405 (.A(_00686_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold406 (.A(\cpu.keccak_alu.registers[209] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold407 (.A(\cpu.keccak_alu.registers[94] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold408 (.A(\cpu.keccak_alu.registers[198] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold409 (.A(\cpu.ALU.a[6] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold410 (.A(_00606_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold411 (.A(\cpu.ALU.b[12] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold412 (.A(\cpu.keccak_alu.registers[250] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold413 (.A(\cpu.keccak_alu.registers[319] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold414 (.A(\cpu.registers[3][1] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold415 (.A(_00280_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold416 (.A(\cpu.keccak_alu.registers[108] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold417 (.A(\cpu.keccak_alu.registers[255] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold418 (.A(_00583_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold419 (.A(\cpu.keccak_alu.registers[22] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold420 (.A(_02306_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold421 (.A(\cpu.registers[6][15] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold422 (.A(_00716_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold423 (.A(\cpu.keccak_alu.registers[11] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold424 (.A(\cpu.keccak_alu.registers[223] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold425 (.A(\cpu.keccak_alu.registers[195] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold426 (.A(\cpu.keccak_alu.registers[278] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold427 (.A(\cpu.registers[1][15] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold428 (.A(_00823_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold429 (.A(\cpu.registers[5][2] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold430 (.A(_00687_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold431 (.A(\cpu.keccak_alu.registers[234] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold432 (.A(\memory_controller.wait_counter[1] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold433 (.A(\cpu.ALU.b[15] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold434 (.A(\cpu.keccak_alu.registers[92] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold435 (.A(\cpu.keccak_alu.registers[259] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold436 (.A(\cpu.keccak_alu.registers[264] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold437 (.A(\cpu.keccak_alu.registers[109] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold438 (.A(\cpu.uart.cycle_counter[5] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold439 (.A(_06552_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold440 (.A(\cpu.keccak_alu.registers[142] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold441 (.A(\cpu.keccak_alu.registers[236] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold442 (.A(\cpu.rx_speed[0] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold443 (.A(\cpu.keccak_alu.registers[206] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold444 (.A(\cpu.registers[2][9] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold445 (.A(_00304_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold446 (.A(\cpu.keccak_alu.registers[33] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold447 (.A(\cpu.keccak_alu.registers[222] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold448 (.A(\cpu.current_address[2] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold449 (.A(_00637_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold450 (.A(\cpu.data_out[3] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold451 (.A(_00654_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold452 (.A(\cpu.current_address[15] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold453 (.A(\cpu.registers[5][6] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold454 (.A(_00691_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold455 (.A(\cpu.keccak_alu.registers[220] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold456 (.A(_00548_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold457 (.A(\cpu.registers[3][6] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold458 (.A(_00285_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold459 (.A(\cpu.keccak_alu.registers[81] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold460 (.A(\cpu.keccak_alu.registers[204] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold461 (.A(\cpu.keccak_alu.registers[197] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold462 (.A(\cpu.registers[2][10] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold463 (.A(_00305_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold464 (.A(\cpu.registers[6][10] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold465 (.A(_00711_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold466 (.A(\cpu.keccak_alu.registers[260] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold467 (.A(\cpu.registers[3][2] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold468 (.A(_00281_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold469 (.A(\cpu.keccak_alu.registers[218] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold470 (.A(\cpu.keccak_alu.registers[105] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold471 (.A(_00433_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold472 (.A(\cpu.keccak_alu.registers[249] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold473 (.A(\cpu.registers[1][2] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold474 (.A(_00311_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold475 (.A(\cpu.keccak_alu.registers[29] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold476 (.A(\cpu.keccak_alu.registers[231] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold477 (.A(\uart_receiver/cycles_per_bit[9] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold478 (.A(\cpu.keccak_alu.registers[85] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold479 (.A(_00144_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold480 (.A(_00566_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold481 (.A(\cpu.keccak_alu.registers[283] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold482 (.A(\cpu.registers[3][5] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold483 (.A(_00284_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold484 (.A(\cpu.keccak_alu.registers[214] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold485 (.A(\cpu.keccak_alu.registers[75] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold486 (.A(\cpu.keccak_alu.registers[245] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold487 (.A(\cpu.keccak_alu.registers[203] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold488 (.A(\cpu.uart.cycle_counter[4] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold489 (.A(_06550_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold490 (.A(\cpu.registers[5][5] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold491 (.A(_00690_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold492 (.A(\cpu.keccak_alu.registers[240] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold493 (.A(\cpu.keccak_alu.registers[286] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold494 (.A(\cpu.registers[6][14] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold495 (.A(_00715_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold496 (.A(\cpu.registers[2][13] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold497 (.A(_00308_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold498 (.A(\memory_controller.read_enable ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold499 (.A(\cpu.keccak_alu.registers[87] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold500 (.A(\cpu.registers[2][0] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold501 (.A(_00295_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold502 (.A(\cpu.keccak_alu.registers[76] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold503 (.A(\uart_receiver/stage[0] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold504 (.A(\uart_receiver/_001_ ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold505 (.A(\cpu.keccak_alu.registers[2] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold506 (.A(\cpu.registers[5][9] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold507 (.A(_00694_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold508 (.A(\cpu.registers[3][7] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold509 (.A(_00286_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold510 (.A(\cpu.keccak_alu.registers[20] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold511 (.A(\cpu.keccak_alu.registers[127] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold512 (.A(\cpu.registers[2][8] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold513 (.A(_00303_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold514 (.A(\cpu.keccak_alu.registers[243] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold515 (.A(\cpu.keccak_alu.registers[254] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold516 (.A(\cpu.registers[2][1] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold517 (.A(_00296_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold518 (.A(\cpu.registers[2][14] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold519 (.A(_00309_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold520 (.A(\cpu.keccak_alu.registers[196] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold521 (.A(\cpu.keccak_alu.registers[232] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold522 (.A(\cpu.keccak_alu.registers[207] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold523 (.A(\cpu.current_address[7] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold524 (.A(_00642_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold525 (.A(\cpu.keccak_alu.registers[69] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold526 (.A(\cpu.registers[2][12] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold527 (.A(_00307_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold528 (.A(\cpu.keccak_alu.registers[284] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold529 (.A(\cpu.keccak_alu.registers[233] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold530 (.A(\cpu.keccak_alu.registers[120] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold531 (.A(\cpu.keccak_alu.registers[106] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold532 (.A(_00434_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold533 (.A(\cpu.keccak_alu.registers[50] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold534 (.A(\cpu.keccak_alu.registers[118] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold535 (.A(\cpu.registers[2][11] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold536 (.A(_00306_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold537 (.A(\cpu.keccak_alu.registers[65] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold538 (.A(\cpu.keccak_alu.registers[279] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold539 (.A(\cpu.keccak_alu.registers[10] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold540 (.A(\cpu.keccak_alu.registers[31] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold541 (.A(\cpu.keccak_alu.registers[51] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold542 (.A(\cpu.keccak_alu.registers[219] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold543 (.A(\cpu.keccak_alu.registers[98] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold544 (.A(\cpu.keccak_alu.registers[281] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold545 (.A(\cpu.keccak_alu.registers[246] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold546 (.A(\cpu.keccak_alu.registers[14] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold547 (.A(\cpu.ALU.b[11] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold548 (.A(\memory_controller.wait_counter[4] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold549 (.A(\cpu.keccak_alu.registers[125] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold550 (.A(_00453_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold551 (.A(\uart_receiver/cycles_per_bit[10] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold552 (.A(\cpu.registers[2][5] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold553 (.A(_00300_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold554 (.A(\cpu.keccak_alu.registers[110] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold555 (.A(\cpu.keccak_alu.registers[201] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold556 (.A(\cpu.keccak_alu.registers[7] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold557 (.A(\cpu.keccak_alu.registers[48] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold558 (.A(\cpu.registers[2][7] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold559 (.A(_00302_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold560 (.A(\cpu.rx_speed[4] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold561 (.A(\uart_receiver/_075_ ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold562 (.A(\cpu.uart.bit_counter[2] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold563 (.A(_00883_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold564 (.A(\cpu.keccak_alu.registers[12] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold565 (.A(\cpu.registers[6][6] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold566 (.A(\cpu.request_address[11] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold567 (.A(\cpu.keccak_alu.registers[9] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold568 (.A(\cpu.keccak_alu.registers[25] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold569 (.A(\cpu.keccak_alu.registers[248] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold570 (.A(_00027_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold571 (.A(_00837_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold572 (.A(\cpu.keccak_alu.registers[103] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold573 (.A(\cpu.registers[5][7] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold574 (.A(_00692_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold575 (.A(\cpu.registers[2][4] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold576 (.A(_00299_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold577 (.A(\cpu.registers[5][4] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold578 (.A(_00689_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold579 (.A(\cpu.keccak_alu.registers[241] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold580 (.A(_00569_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold581 (.A(\cpu.keccak_alu.registers[30] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold582 (.A(\cpu.keccak_alu.registers[84] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold583 (.A(\cpu.registers[3][11] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold584 (.A(_00290_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold585 (.A(\cpu.keccak_alu.registers[71] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold586 (.A(\cpu.keccak_alu.registers[135] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold587 (.A(\cpu.ALU.b[10] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold588 (.A(\cpu.keccak_alu.registers[271] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold589 (.A(\cpu.keccak_alu.registers[114] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold590 (.A(\cpu.keccak_alu.registers[268] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold591 (.A(\cpu.keccak_alu.registers[54] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold592 (.A(\cpu.keccak_alu.registers[66] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold593 (.A(\cpu.request_address[12] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold594 (.A(\cpu.keccak_alu.registers[13] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold595 (.A(\cpu.keccak_alu.registers[8] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold596 (.A(\cpu.keccak_alu.registers[251] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold597 (.A(\cpu.keccak_alu.registers[221] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold598 (.A(\cpu.keccak_alu.registers[97] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold599 (.A(\cpu.keccak_alu.registers[107] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold600 (.A(\cpu.keccak_alu.registers[86] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold601 (.A(\cpu.registers[3][0] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold602 (.A(_00279_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold603 (.A(\cpu.keccak_alu.registers[80] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold604 (.A(\cpu.registers[3][14] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold605 (.A(_00293_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold606 (.A(\cpu.keccak_alu.registers[4] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold607 (.A(\cpu.keccak_alu.registers[211] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold608 (.A(\cpu.registers[2][6] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold609 (.A(_00301_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold610 (.A(\cpu.keccak_alu.registers[35] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold611 (.A(\cpu.registers[3][3] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold612 (.A(_00282_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold613 (.A(\cpu.rx_speed[3] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold614 (.A(\cpu.keccak_alu.registers[117] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold615 (.A(\cpu.rx_speed[2] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold616 (.A(\cpu.ALU.b[13] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold617 (.A(\cpu.keccak_alu.registers[68] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold618 (.A(\cpu.keccak_alu.registers[23] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold619 (.A(\cpu.keccak_alu.registers[104] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold620 (.A(\cpu.keccak_alu.registers[67] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold621 (.A(\cpu.keccak_alu.registers[17] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold622 (.A(\uart_receiver/cycles_per_bit[7] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold623 (.A(\uart_receiver/_078_ ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold624 (.A(_00130_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold625 (.A(_00488_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold626 (.A(\cpu.keccak_alu.registers[52] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold627 (.A(\uart_receiver/cycles_per_bit[1] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold628 (.A(\cpu.registers[3][12] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold629 (.A(_00291_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold630 (.A(\cpu.keccak_alu.registers[102] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold631 (.A(\cpu.keccak_alu.registers[205] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold632 (.A(\uart_receiver/cycles_per_bit[8] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold633 (.A(\cpu.keccak_alu.registers[6] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold634 (.A(\cpu.registers[3][13] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold635 (.A(_00292_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold636 (.A(\cpu.keccak_alu.registers[119] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold637 (.A(\cpu.keccak_alu.registers[63] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold638 (.A(\cpu.registers[5][15] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold639 (.A(_00700_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold640 (.A(\cpu.keccak_alu.registers[38] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold641 (.A(_02341_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold642 (.A(\cpu.keccak_alu.registers[49] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold643 (.A(\cpu.keccak_alu.registers[57] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold644 (.A(\cpu.keccak_alu.registers[32] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold645 (.A(\cpu.ALU.a[14] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold646 (.A(_00614_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold647 (.A(\cpu.keccak_alu.registers[0] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold648 (.A(\cpu.keccak_alu.registers[124] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold649 (.A(\memory_controller.wait_counter[5] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold650 (.A(\cpu.registers[5][12] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold651 (.A(_00697_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold652 (.A(\cpu.keccak_alu.registers[40] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold653 (.A(\cpu.keccak_alu.registers[26] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold654 (.A(\cpu.keccak_alu.registers[300] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold655 (.A(_00761_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold656 (.A(\cpu.keccak_alu.registers[228] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold657 (.A(\cpu.keccak_alu.registers[115] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold658 (.A(\cpu.keccak_alu.registers[37] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold659 (.A(\cpu.current_address[0] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold660 (.A(_00635_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold661 (.A(\cpu.uart.cycle_counter[8] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold662 (.A(_06557_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold663 (.A(\cpu.rx_speed[7] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold664 (.A(_00322_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold665 (.A(\cpu.keccak_alu.registers[235] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold666 (.A(\cpu.keccak_alu.registers[15] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold667 (.A(\cpu.keccak_alu.registers[3] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold668 (.A(\cpu.registers[3][9] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold669 (.A(_00288_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold670 (.A(\cpu.keccak_alu.registers[46] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold671 (.A(\cpu.keccak_alu.registers[36] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold672 (.A(_02337_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold673 (.A(\cpu.registers[5][14] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold674 (.A(_00699_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold675 (.A(\cpu.keccak_alu.registers[244] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold676 (.A(\cpu.data_out[0] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold677 (.A(_00651_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold678 (.A(\cpu.keccak_alu.registers[99] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold679 (.A(\cpu.keccak_alu.registers[282] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold680 (.A(\uart_receiver/cycle_counter[7] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold681 (.A(\cpu.keccak_alu.registers[28] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold682 (.A(\cpu.keccak_alu.registers[112] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold683 (.A(\uart_receiver/cycle_counter[3] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold684 (.A(\uart_receiver/_087_ ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold685 (.A(\cpu.registers[3][10] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold686 (.A(_00289_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold687 (.A(\cpu.keccak_alu.registers[111] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold688 (.A(\cpu.uart.cycle_counter[12] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold689 (.A(\uart_receiver/_004_ ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold690 (.A(\uart_receiver/_106_ ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold691 (.A(\uart_receiver/cycle_counter[9] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold692 (.A(\uart_receiver/_093_ ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold693 (.A(\cpu.registers[3][15] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold694 (.A(_00294_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold695 (.A(\cpu.registers[5][11] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold696 (.A(_00696_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold697 (.A(\cpu.keccak_alu.registers[113] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold698 (.A(\cpu.keccak_alu.registers[60] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold699 (.A(\cpu.request_address[10] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold700 (.A(_00678_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold701 (.A(\cpu.keccak_alu.registers[83] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold702 (.A(uio_out[1]),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold703 (.A(_00798_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold704 (.A(\data_received[7] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold705 (.A(_00804_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold706 (.A(\cpu.uart.cycle_counter[2] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold707 (.A(\cpu.keccak_alu.registers[24] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold708 (.A(\cpu.registers[5][3] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold709 (.A(_00688_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold710 (.A(\cpu.keccak_alu.registers[116] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold711 (.A(\cpu.keccak_alu.registers[126] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold712 (.A(\cpu.registers[5][8] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold713 (.A(_00693_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold714 (.A(\cpu.registers[5][13] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold715 (.A(_00698_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold716 (.A(\cpu.keccak_alu.registers[89] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold717 (.A(\cpu.keccak_alu.registers[61] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold718 (.A(uio_out[4]),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold719 (.A(\cpu.keccak_alu.registers[55] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold720 (.A(\cpu.uart.cycle_counter[6] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold721 (.A(\cpu.keccak_alu.registers[144] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold722 (.A(\cpu.keccak_alu.registers[79] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold723 (.A(\cpu.keccak_alu.registers[27] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold724 (.A(\cpu.keccak_alu.registers[58] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold725 (.A(\cpu.request_address[9] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold726 (.A(\cpu.ALU.a[12] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold727 (.A(_00612_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold728 (.A(\cpu.registers[5][0] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold729 (.A(_00685_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold730 (.A(\cpu.keccak_alu.registers[242] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold731 (.A(uio_out[3]),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold732 (.A(_00800_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold733 (.A(\cpu.keccak_alu.registers[123] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold734 (.A(\cpu.registers[2][3] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold735 (.A(_00298_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold736 (.A(\cpu.keccak_alu.registers[96] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold737 (.A(\cpu.keccak_alu.registers[43] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold738 (.A(\cpu.ALU.b[9] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold739 (.A(\cpu.keccak_alu.registers[16] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold740 (.A(\cpu.keccak_alu.registers[42] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold741 (.A(\cpu.keccak_alu.registers[121] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold742 (.A(_00449_),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold743 (.A(\uart_receiver/bit_counter[0] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold744 (.A(\uart_receiver/_105_ ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold745 (.A(\cpu.request_address[13] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold746 (.A(_00681_),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold747 (.A(\uart_receiver/_003_ ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold748 (.A(\uart_receiver/_094_ ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold749 (.A(\cpu.keccak_alu.registers[59] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold750 (.A(\cpu.keccak_alu.registers[47] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold751 (.A(\cpu.keccak_alu.registers[70] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold752 (.A(\cpu.keccak_alu.registers[56] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold753 (.A(\cpu.registers[5][10] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold754 (.A(_00695_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold755 (.A(\cpu.keccak_alu.registers[216] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold756 (.A(\cpu.keccak_alu.registers[39] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold757 (.A(\cpu.keccak_alu.registers[45] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold758 (.A(\cpu.keccak_alu.registers[53] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold759 (.A(uio_out[5]),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold760 (.A(\cpu.keccak_alu.registers[213] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold761 (.A(_00541_),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold762 (.A(\memory_controller.register_enable ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold763 (.A(\uart_receiver/cycle_counter[8] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold764 (.A(uio_out[2]),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold765 (.A(\cpu.keccak_alu.registers[62] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold766 (.A(\cpu.keccak_alu.registers[19] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold767 (.A(\cpu.uart.stage[2] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold768 (.A(\cpu.keccak_alu.registers[21] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold769 (.A(_00133_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold770 (.A(\cpu.ALU.b[8] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold771 (.A(_00045_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold772 (.A(_02828_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold773 (.A(_00616_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold774 (.A(\cpu.ALU.mode[1] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold775 (.A(uio_out[0]),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold776 (.A(_00797_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold777 (.A(\uart_receiver/cycle_counter[6] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold778 (.A(\uart_receiver/_090_ ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold779 (.A(\cpu.registers[3][8] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold780 (.A(_00287_),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold781 (.A(\cpu.keccak_alu.registers[122] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold782 (.A(_00450_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold783 (.A(\cpu.keccak_alu.registers[41] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold784 (.A(\cpu.ALU.b[1] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold785 (.A(\cpu.ALU.a[15] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold786 (.A(_00615_),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold787 (.A(\cpu.request_address[14] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold788 (.A(\uart_receiver/cycle_counter[11] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold789 (.A(\uart_receiver/_095_ ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold790 (.A(\cpu.keccak_alu.registers[100] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold791 (.A(\cpu.execution_stage[1] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold792 (.A(uio_out[6]),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold793 (.A(\cpu.ALU.b[7] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold794 (.A(\uart_receiver/cycles_per_bit[2] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold795 (.A(\uart_receiver/_002_ ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold796 (.A(\uart_receiver/_000_ ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold797 (.A(\cpu.ALU.a[11] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold798 (.A(_00611_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold799 (.A(\cpu.uart.stage[1] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold800 (.A(_00005_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold801 (.A(\cpu.current_address[1] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold802 (.A(_00636_),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold803 (.A(\uart_receiver/cycle_counter[12] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold804 (.A(\cpu.ALU.a[5] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold805 (.A(_00605_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold806 (.A(\cpu.request_address[0] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold807 (.A(\cpu.keccak_alu.registers[44] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold808 (.A(\uart_receiver/cycle_counter[0] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold809 (.A(\uart_receiver/_084_ ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold810 (.A(\cpu.keccak_alu.registers[184] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold811 (.A(\cpu.keccak_alu.registers[140] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold812 (.A(_00468_),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold813 (.A(_00017_),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold814 (.A(_00004_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold815 (.A(\cpu.ALU.a[9] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold816 (.A(_00609_),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold817 (.A(\uart_receiver/cycle_counter[1] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold818 (.A(\uart_receiver/_085_ ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold819 (.A(\cpu.keccak_alu.registers[183] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold820 (.A(\cpu.ALU.a[7] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold821 (.A(_00607_),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold822 (.A(\uart_receiver/cycles_per_bit[5] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold823 (.A(\uart_receiver/_089_ ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold824 (.A(\cpu.ALU.a[4] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold825 (.A(_00604_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold826 (.A(\cpu.uart.bit_counter[1] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold827 (.A(_00882_),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold828 (.A(_00136_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold829 (.A(_00510_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold830 (.A(\cpu.keccak_alu.registers[138] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold831 (.A(\cpu.ALU.a[1] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold832 (.A(_00601_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold833 (.A(_00134_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold834 (.A(_00508_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold835 (.A(\cpu.ALU.a[13] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold836 (.A(_00613_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold837 (.A(\cpu.request_address[8] ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold838 (.A(\cpu.ALU.a[0] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold839 (.A(_00600_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold840 (.A(\uart_receiver/cycles_per_bit[4] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold841 (.A(\uart_receiver/_257_ ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold842 (.A(\uart_receiver/_088_ ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold843 (.A(\cpu.keccak_alu.registers[139] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold844 (.A(\cpu.keccak_alu.registers[101] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold845 (.A(\cpu.request_address[1] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold846 (.A(_00669_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold847 (.A(\cpu.ALU.b[0] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold848 (.A(_00584_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold849 (.A(\cpu.ALU.a[10] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold850 (.A(\cpu.ALU.a[8] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold851 (.A(_00608_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold852 (.A(\cpu.keccak_alu.registers[131] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold853 (.A(\cpu.keccak_alu.registers[190] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold854 (.A(\cpu.keccak_alu.registers[156] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold855 (.A(\cpu.keccak_alu.registers[136] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold856 (.A(\cpu.ALU.b[4] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold857 (.A(\cpu.request_address[2] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold858 (.A(\cpu.keccak_alu.registers[155] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold859 (.A(\cpu.request_address[7] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold860 (.A(\cpu.registers[1][1] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold861 (.A(_06993_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold862 (.A(\cpu.keccak_alu.registers[159] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold863 (.A(\uart_receiver/cycle_counter[2] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold864 (.A(\cpu.keccak_alu.registers[154] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold865 (.A(\cpu.ALU.a[3] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold866 (.A(_00603_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold867 (.A(\cpu.keccak_alu.registers[191] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold868 (.A(_00519_),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold869 (.A(\cpu.ALU.a[2] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold870 (.A(_00602_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold871 (.A(\cpu.ALU.b[3] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold872 (.A(uio_oe[7]),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold873 (.A(_00161_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold874 (.A(_00671_),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold875 (.A(\memory_controller.upper_bit ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold876 (.A(\cpu.ALU.b[5] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold877 (.A(\cpu.keccak_alu.registers[187] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold878 (.A(\cpu.keccak_alu.registers[143] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold879 (.A(\cpu.keccak_alu.registers[149] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold880 (.A(\cpu.keccak_alu.registers[170] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold881 (.A(\cpu.ALU.b[2] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold882 (.A(\cpu.keccak_alu.registers[168] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold883 (.A(\cpu.ALU.b[6] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold884 (.A(\cpu.keccak_alu.registers[141] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold885 (.A(_00469_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold886 (.A(\cpu.request_address[5] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold887 (.A(\cpu.keccak_alu.registers[151] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold888 (.A(\cpu.keccak_alu.registers[148] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold889 (.A(\cpu.keccak_alu.registers[185] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold890 (.A(\cpu.keccak_alu.registers[188] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold891 (.A(\cpu.keccak_alu.registers[171] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold892 (.A(\cpu.keccak_alu.registers[178] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold893 (.A(\cpu.keccak_alu.registers[158] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold894 (.A(\cpu.keccak_alu.registers[174] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold895 (.A(\cpu.request_address[4] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold896 (.A(\cpu.keccak_alu.registers[132] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold897 (.A(\cpu.keccak_alu.registers[186] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold898 (.A(\cpu.keccak_alu.registers[166] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold899 (.A(\cpu.keccak_alu.registers[153] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold900 (.A(\cpu.uart.bit_counter[0] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold901 (.A(_00881_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold902 (.A(\cpu.keccak_alu.registers[169] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold903 (.A(\cpu.keccak_alu.registers[150] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold904 (.A(_00135_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold905 (.A(_00493_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold906 (.A(\cpu.keccak_alu.registers[145] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold907 (.A(_00473_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold908 (.A(\cpu.keccak_alu.registers[162] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold909 (.A(\cpu.keccak_alu.registers[137] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold910 (.A(_00465_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold911 (.A(\cpu.request_address[6] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold912 (.A(\cpu.keccak_alu.registers[177] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold913 (.A(\cpu.keccak_alu.registers[173] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold914 (.A(\cpu.keccak_alu.registers[179] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold915 (.A(_00023_),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold916 (.A(_00001_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold917 (.A(\cpu.keccak_alu.registers[175] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold918 (.A(\cpu.keccak_alu.registers[189] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold919 (.A(_00131_),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold920 (.A(_00489_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold921 (.A(\cpu.keccak_alu.registers[129] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold922 (.A(\cpu.keccak_alu.registers[146] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold923 (.A(\cpu.keccak_alu.registers[164] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold924 (.A(\cpu.keccak_alu.registers[167] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold925 (.A(\cpu.keccak_alu.registers[157] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold926 (.A(\cpu.registers[1][0] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold927 (.A(\cpu.keccak_alu.registers[152] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold928 (.A(_00019_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold929 (.A(\memory_controller.wait_counter[4] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold930 (.A(_06414_),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold931 (.A(\cpu.keccak_alu.registers[63] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold932 (.A(\uart_receiver/bit_counter[0] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold933 (.A(\uart_receiver/stage[0] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold934 (.A(\cpu.keccak_alu.registers[30] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold935 (.A(\cpu.keccak_alu.registers[13] ),
    .X(net953));
 sg13g2_antennanp ANTENNA_1 (.A(_00076_));
 sg13g2_antennanp ANTENNA_2 (.A(_00076_));
 sg13g2_antennanp ANTENNA_3 (.A(_00076_));
 sg13g2_antennanp ANTENNA_4 (.A(_00076_));
 sg13g2_antennanp ANTENNA_5 (.A(_00092_));
 sg13g2_antennanp ANTENNA_6 (.A(_00092_));
 sg13g2_antennanp ANTENNA_7 (.A(_00092_));
 sg13g2_antennanp ANTENNA_8 (.A(_00092_));
 sg13g2_antennanp ANTENNA_9 (.A(_00096_));
 sg13g2_antennanp ANTENNA_10 (.A(_00096_));
 sg13g2_antennanp ANTENNA_11 (.A(_00260_));
 sg13g2_antennanp ANTENNA_12 (.A(_01413_));
 sg13g2_antennanp ANTENNA_13 (.A(_01413_));
 sg13g2_antennanp ANTENNA_14 (.A(_01413_));
 sg13g2_antennanp ANTENNA_15 (.A(_01413_));
 sg13g2_antennanp ANTENNA_16 (.A(_01413_));
 sg13g2_antennanp ANTENNA_17 (.A(_02977_));
 sg13g2_antennanp ANTENNA_18 (.A(_03001_));
 sg13g2_antennanp ANTENNA_19 (.A(_03025_));
 sg13g2_antennanp ANTENNA_20 (.A(_04794_));
 sg13g2_antennanp ANTENNA_21 (.A(_04858_));
 sg13g2_antennanp ANTENNA_22 (.A(_04890_));
 sg13g2_antennanp ANTENNA_23 (.A(_04988_));
 sg13g2_antennanp ANTENNA_24 (.A(_05018_));
 sg13g2_antennanp ANTENNA_25 (.A(_05045_));
 sg13g2_antennanp ANTENNA_26 (.A(_05313_));
 sg13g2_antennanp ANTENNA_27 (.A(_05341_));
 sg13g2_antennanp ANTENNA_28 (.A(_05424_));
 sg13g2_antennanp ANTENNA_29 (.A(_05445_));
 sg13g2_antennanp ANTENNA_30 (.A(_05472_));
 sg13g2_antennanp ANTENNA_31 (.A(_05723_));
 sg13g2_antennanp ANTENNA_32 (.A(_05770_));
 sg13g2_antennanp ANTENNA_33 (.A(_05814_));
 sg13g2_antennanp ANTENNA_34 (.A(_06102_));
 sg13g2_antennanp ANTENNA_35 (.A(_06197_));
 sg13g2_antennanp ANTENNA_36 (.A(_06243_));
 sg13g2_antennanp ANTENNA_37 (.A(clk));
 sg13g2_antennanp ANTENNA_38 (.A(_00074_));
 sg13g2_antennanp ANTENNA_39 (.A(_00074_));
 sg13g2_antennanp ANTENNA_40 (.A(_00076_));
 sg13g2_antennanp ANTENNA_41 (.A(_00076_));
 sg13g2_antennanp ANTENNA_42 (.A(_00076_));
 sg13g2_antennanp ANTENNA_43 (.A(_00076_));
 sg13g2_antennanp ANTENNA_44 (.A(_00096_));
 sg13g2_antennanp ANTENNA_45 (.A(_00096_));
 sg13g2_antennanp ANTENNA_46 (.A(_00096_));
 sg13g2_antennanp ANTENNA_47 (.A(_00096_));
 sg13g2_antennanp ANTENNA_48 (.A(_00260_));
 sg13g2_antennanp ANTENNA_49 (.A(_02977_));
 sg13g2_antennanp ANTENNA_50 (.A(_03001_));
 sg13g2_antennanp ANTENNA_51 (.A(_03025_));
 sg13g2_antennanp ANTENNA_52 (.A(_04858_));
 sg13g2_antennanp ANTENNA_53 (.A(_04890_));
 sg13g2_antennanp ANTENNA_54 (.A(_04988_));
 sg13g2_antennanp ANTENNA_55 (.A(_05018_));
 sg13g2_antennanp ANTENNA_56 (.A(_05045_));
 sg13g2_antennanp ANTENNA_57 (.A(_05313_));
 sg13g2_antennanp ANTENNA_58 (.A(_05341_));
 sg13g2_antennanp ANTENNA_59 (.A(_05424_));
 sg13g2_antennanp ANTENNA_60 (.A(_05445_));
 sg13g2_antennanp ANTENNA_61 (.A(_05472_));
 sg13g2_antennanp ANTENNA_62 (.A(_05723_));
 sg13g2_antennanp ANTENNA_63 (.A(_05770_));
 sg13g2_antennanp ANTENNA_64 (.A(_05814_));
 sg13g2_antennanp ANTENNA_65 (.A(_06102_));
 sg13g2_antennanp ANTENNA_66 (.A(_06197_));
 sg13g2_antennanp ANTENNA_67 (.A(_06243_));
 sg13g2_antennanp ANTENNA_68 (.A(clk));
 sg13g2_antennanp ANTENNA_69 (.A(clk));
 sg13g2_antennanp ANTENNA_70 (.A(_00096_));
 sg13g2_antennanp ANTENNA_71 (.A(_00096_));
 sg13g2_antennanp ANTENNA_72 (.A(_02977_));
 sg13g2_antennanp ANTENNA_73 (.A(_03001_));
 sg13g2_antennanp ANTENNA_74 (.A(_03025_));
 sg13g2_antennanp ANTENNA_75 (.A(_04858_));
 sg13g2_antennanp ANTENNA_76 (.A(_04890_));
 sg13g2_antennanp ANTENNA_77 (.A(_04988_));
 sg13g2_antennanp ANTENNA_78 (.A(_05018_));
 sg13g2_antennanp ANTENNA_79 (.A(_05045_));
 sg13g2_antennanp ANTENNA_80 (.A(_05313_));
 sg13g2_antennanp ANTENNA_81 (.A(_05341_));
 sg13g2_antennanp ANTENNA_82 (.A(_05424_));
 sg13g2_antennanp ANTENNA_83 (.A(_05445_));
 sg13g2_antennanp ANTENNA_84 (.A(_05472_));
 sg13g2_antennanp ANTENNA_85 (.A(_05723_));
 sg13g2_antennanp ANTENNA_86 (.A(_05770_));
 sg13g2_antennanp ANTENNA_87 (.A(_05814_));
 sg13g2_antennanp ANTENNA_88 (.A(_06102_));
 sg13g2_antennanp ANTENNA_89 (.A(_06197_));
 sg13g2_antennanp ANTENNA_90 (.A(_06243_));
 sg13g2_antennanp ANTENNA_91 (.A(clk));
 sg13g2_antennanp ANTENNA_92 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_583 ();
 sg13g2_decap_8 FILLER_0_610 ();
 sg13g2_decap_8 FILLER_0_617 ();
 sg13g2_fill_1 FILLER_0_624 ();
 sg13g2_decap_8 FILLER_0_654 ();
 sg13g2_decap_4 FILLER_0_661 ();
 sg13g2_fill_1 FILLER_0_665 ();
 sg13g2_fill_2 FILLER_0_676 ();
 sg13g2_decap_8 FILLER_0_699 ();
 sg13g2_decap_8 FILLER_0_706 ();
 sg13g2_decap_4 FILLER_0_713 ();
 sg13g2_decap_4 FILLER_0_725 ();
 sg13g2_fill_2 FILLER_0_729 ();
 sg13g2_fill_1 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_fill_1 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_fill_1 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_802 ();
 sg13g2_decap_8 FILLER_0_809 ();
 sg13g2_decap_8 FILLER_0_816 ();
 sg13g2_decap_8 FILLER_0_823 ();
 sg13g2_decap_8 FILLER_0_830 ();
 sg13g2_fill_1 FILLER_0_837 ();
 sg13g2_decap_4 FILLER_0_856 ();
 sg13g2_fill_2 FILLER_0_860 ();
 sg13g2_decap_8 FILLER_0_881 ();
 sg13g2_decap_8 FILLER_0_888 ();
 sg13g2_decap_4 FILLER_0_895 ();
 sg13g2_fill_1 FILLER_0_899 ();
 sg13g2_decap_8 FILLER_0_939 ();
 sg13g2_decap_8 FILLER_0_946 ();
 sg13g2_fill_2 FILLER_0_953 ();
 sg13g2_fill_1 FILLER_0_955 ();
 sg13g2_decap_4 FILLER_0_964 ();
 sg13g2_fill_2 FILLER_0_978 ();
 sg13g2_fill_1 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_989 ();
 sg13g2_decap_8 FILLER_0_996 ();
 sg13g2_decap_8 FILLER_0_1003 ();
 sg13g2_fill_2 FILLER_0_1020 ();
 sg13g2_decap_8 FILLER_0_1032 ();
 sg13g2_decap_8 FILLER_0_1039 ();
 sg13g2_decap_8 FILLER_0_1046 ();
 sg13g2_decap_8 FILLER_0_1053 ();
 sg13g2_decap_8 FILLER_0_1060 ();
 sg13g2_decap_8 FILLER_0_1067 ();
 sg13g2_decap_8 FILLER_0_1074 ();
 sg13g2_decap_8 FILLER_0_1081 ();
 sg13g2_decap_8 FILLER_0_1088 ();
 sg13g2_decap_8 FILLER_0_1095 ();
 sg13g2_decap_8 FILLER_0_1102 ();
 sg13g2_decap_8 FILLER_0_1109 ();
 sg13g2_decap_8 FILLER_0_1116 ();
 sg13g2_decap_8 FILLER_0_1123 ();
 sg13g2_decap_8 FILLER_0_1130 ();
 sg13g2_decap_8 FILLER_0_1137 ();
 sg13g2_decap_8 FILLER_0_1144 ();
 sg13g2_decap_8 FILLER_0_1151 ();
 sg13g2_decap_8 FILLER_0_1158 ();
 sg13g2_decap_8 FILLER_0_1165 ();
 sg13g2_decap_8 FILLER_0_1172 ();
 sg13g2_decap_8 FILLER_0_1179 ();
 sg13g2_decap_8 FILLER_0_1186 ();
 sg13g2_decap_8 FILLER_0_1193 ();
 sg13g2_decap_8 FILLER_0_1200 ();
 sg13g2_decap_8 FILLER_0_1207 ();
 sg13g2_decap_8 FILLER_0_1214 ();
 sg13g2_decap_8 FILLER_0_1221 ();
 sg13g2_decap_8 FILLER_0_1228 ();
 sg13g2_decap_8 FILLER_0_1235 ();
 sg13g2_decap_8 FILLER_0_1242 ();
 sg13g2_decap_8 FILLER_0_1249 ();
 sg13g2_decap_8 FILLER_0_1256 ();
 sg13g2_decap_8 FILLER_0_1263 ();
 sg13g2_decap_8 FILLER_0_1270 ();
 sg13g2_decap_8 FILLER_0_1277 ();
 sg13g2_decap_8 FILLER_0_1284 ();
 sg13g2_decap_8 FILLER_0_1291 ();
 sg13g2_decap_8 FILLER_0_1298 ();
 sg13g2_decap_8 FILLER_0_1305 ();
 sg13g2_decap_8 FILLER_0_1312 ();
 sg13g2_decap_8 FILLER_0_1319 ();
 sg13g2_decap_8 FILLER_0_1326 ();
 sg13g2_decap_8 FILLER_0_1333 ();
 sg13g2_decap_8 FILLER_0_1340 ();
 sg13g2_decap_8 FILLER_0_1347 ();
 sg13g2_decap_8 FILLER_0_1354 ();
 sg13g2_decap_8 FILLER_0_1361 ();
 sg13g2_decap_8 FILLER_0_1368 ();
 sg13g2_decap_8 FILLER_0_1375 ();
 sg13g2_decap_8 FILLER_0_1382 ();
 sg13g2_decap_8 FILLER_0_1389 ();
 sg13g2_decap_8 FILLER_0_1396 ();
 sg13g2_decap_8 FILLER_0_1403 ();
 sg13g2_decap_8 FILLER_0_1410 ();
 sg13g2_decap_8 FILLER_0_1417 ();
 sg13g2_decap_8 FILLER_0_1424 ();
 sg13g2_decap_8 FILLER_0_1431 ();
 sg13g2_decap_8 FILLER_0_1438 ();
 sg13g2_decap_8 FILLER_0_1445 ();
 sg13g2_decap_8 FILLER_0_1452 ();
 sg13g2_decap_8 FILLER_0_1459 ();
 sg13g2_decap_8 FILLER_0_1466 ();
 sg13g2_decap_8 FILLER_0_1473 ();
 sg13g2_decap_8 FILLER_0_1480 ();
 sg13g2_decap_8 FILLER_0_1487 ();
 sg13g2_decap_8 FILLER_0_1494 ();
 sg13g2_decap_8 FILLER_0_1501 ();
 sg13g2_decap_8 FILLER_0_1508 ();
 sg13g2_decap_8 FILLER_0_1515 ();
 sg13g2_decap_8 FILLER_0_1522 ();
 sg13g2_decap_8 FILLER_0_1529 ();
 sg13g2_decap_8 FILLER_0_1536 ();
 sg13g2_decap_8 FILLER_0_1543 ();
 sg13g2_decap_8 FILLER_0_1550 ();
 sg13g2_decap_8 FILLER_0_1557 ();
 sg13g2_decap_8 FILLER_0_1564 ();
 sg13g2_decap_8 FILLER_0_1571 ();
 sg13g2_decap_8 FILLER_0_1578 ();
 sg13g2_decap_8 FILLER_0_1585 ();
 sg13g2_decap_8 FILLER_0_1592 ();
 sg13g2_decap_8 FILLER_0_1599 ();
 sg13g2_decap_8 FILLER_0_1606 ();
 sg13g2_decap_8 FILLER_0_1613 ();
 sg13g2_decap_8 FILLER_0_1620 ();
 sg13g2_decap_8 FILLER_0_1627 ();
 sg13g2_decap_8 FILLER_0_1634 ();
 sg13g2_decap_8 FILLER_0_1641 ();
 sg13g2_decap_8 FILLER_0_1648 ();
 sg13g2_decap_8 FILLER_0_1655 ();
 sg13g2_decap_8 FILLER_0_1662 ();
 sg13g2_decap_8 FILLER_0_1669 ();
 sg13g2_decap_8 FILLER_0_1676 ();
 sg13g2_decap_8 FILLER_0_1683 ();
 sg13g2_decap_8 FILLER_0_1690 ();
 sg13g2_decap_8 FILLER_0_1697 ();
 sg13g2_decap_8 FILLER_0_1704 ();
 sg13g2_decap_8 FILLER_0_1711 ();
 sg13g2_decap_8 FILLER_0_1718 ();
 sg13g2_decap_8 FILLER_0_1725 ();
 sg13g2_decap_8 FILLER_0_1732 ();
 sg13g2_decap_8 FILLER_0_1739 ();
 sg13g2_decap_8 FILLER_0_1746 ();
 sg13g2_decap_8 FILLER_0_1753 ();
 sg13g2_decap_8 FILLER_0_1760 ();
 sg13g2_fill_1 FILLER_0_1767 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_4 FILLER_1_546 ();
 sg13g2_fill_2 FILLER_1_550 ();
 sg13g2_decap_4 FILLER_1_590 ();
 sg13g2_fill_1 FILLER_1_594 ();
 sg13g2_decap_8 FILLER_1_625 ();
 sg13g2_decap_4 FILLER_1_632 ();
 sg13g2_decap_4 FILLER_1_682 ();
 sg13g2_fill_1 FILLER_1_707 ();
 sg13g2_decap_4 FILLER_1_716 ();
 sg13g2_decap_4 FILLER_1_736 ();
 sg13g2_fill_1 FILLER_1_740 ();
 sg13g2_fill_2 FILLER_1_768 ();
 sg13g2_decap_8 FILLER_1_811 ();
 sg13g2_fill_1 FILLER_1_818 ();
 sg13g2_decap_4 FILLER_1_832 ();
 sg13g2_decap_4 FILLER_1_841 ();
 sg13g2_fill_2 FILLER_1_845 ();
 sg13g2_fill_1 FILLER_1_857 ();
 sg13g2_decap_4 FILLER_1_910 ();
 sg13g2_fill_2 FILLER_1_914 ();
 sg13g2_fill_2 FILLER_1_995 ();
 sg13g2_fill_1 FILLER_1_997 ();
 sg13g2_fill_2 FILLER_1_1050 ();
 sg13g2_decap_4 FILLER_1_1060 ();
 sg13g2_decap_8 FILLER_1_1072 ();
 sg13g2_decap_8 FILLER_1_1084 ();
 sg13g2_decap_8 FILLER_1_1091 ();
 sg13g2_decap_8 FILLER_1_1098 ();
 sg13g2_decap_8 FILLER_1_1105 ();
 sg13g2_decap_8 FILLER_1_1112 ();
 sg13g2_decap_8 FILLER_1_1119 ();
 sg13g2_decap_8 FILLER_1_1126 ();
 sg13g2_decap_8 FILLER_1_1133 ();
 sg13g2_decap_8 FILLER_1_1140 ();
 sg13g2_decap_8 FILLER_1_1147 ();
 sg13g2_decap_8 FILLER_1_1154 ();
 sg13g2_decap_8 FILLER_1_1161 ();
 sg13g2_decap_8 FILLER_1_1168 ();
 sg13g2_decap_8 FILLER_1_1175 ();
 sg13g2_decap_8 FILLER_1_1182 ();
 sg13g2_decap_8 FILLER_1_1189 ();
 sg13g2_decap_8 FILLER_1_1196 ();
 sg13g2_decap_8 FILLER_1_1203 ();
 sg13g2_decap_8 FILLER_1_1210 ();
 sg13g2_decap_8 FILLER_1_1217 ();
 sg13g2_decap_8 FILLER_1_1224 ();
 sg13g2_decap_8 FILLER_1_1231 ();
 sg13g2_decap_8 FILLER_1_1238 ();
 sg13g2_decap_8 FILLER_1_1245 ();
 sg13g2_decap_8 FILLER_1_1252 ();
 sg13g2_decap_8 FILLER_1_1259 ();
 sg13g2_decap_8 FILLER_1_1266 ();
 sg13g2_decap_8 FILLER_1_1273 ();
 sg13g2_decap_8 FILLER_1_1280 ();
 sg13g2_decap_8 FILLER_1_1287 ();
 sg13g2_decap_8 FILLER_1_1294 ();
 sg13g2_decap_8 FILLER_1_1301 ();
 sg13g2_decap_8 FILLER_1_1308 ();
 sg13g2_decap_8 FILLER_1_1315 ();
 sg13g2_decap_8 FILLER_1_1322 ();
 sg13g2_decap_8 FILLER_1_1329 ();
 sg13g2_decap_8 FILLER_1_1336 ();
 sg13g2_decap_8 FILLER_1_1343 ();
 sg13g2_decap_8 FILLER_1_1350 ();
 sg13g2_decap_8 FILLER_1_1357 ();
 sg13g2_decap_8 FILLER_1_1364 ();
 sg13g2_decap_8 FILLER_1_1371 ();
 sg13g2_decap_8 FILLER_1_1378 ();
 sg13g2_decap_8 FILLER_1_1385 ();
 sg13g2_decap_8 FILLER_1_1392 ();
 sg13g2_decap_8 FILLER_1_1399 ();
 sg13g2_decap_8 FILLER_1_1406 ();
 sg13g2_decap_8 FILLER_1_1413 ();
 sg13g2_decap_8 FILLER_1_1420 ();
 sg13g2_decap_8 FILLER_1_1427 ();
 sg13g2_decap_8 FILLER_1_1434 ();
 sg13g2_decap_8 FILLER_1_1441 ();
 sg13g2_decap_8 FILLER_1_1448 ();
 sg13g2_decap_8 FILLER_1_1455 ();
 sg13g2_decap_8 FILLER_1_1462 ();
 sg13g2_decap_8 FILLER_1_1469 ();
 sg13g2_decap_8 FILLER_1_1476 ();
 sg13g2_decap_8 FILLER_1_1483 ();
 sg13g2_decap_8 FILLER_1_1490 ();
 sg13g2_decap_8 FILLER_1_1497 ();
 sg13g2_decap_8 FILLER_1_1504 ();
 sg13g2_decap_8 FILLER_1_1511 ();
 sg13g2_decap_8 FILLER_1_1518 ();
 sg13g2_decap_8 FILLER_1_1525 ();
 sg13g2_decap_8 FILLER_1_1532 ();
 sg13g2_decap_8 FILLER_1_1539 ();
 sg13g2_decap_8 FILLER_1_1546 ();
 sg13g2_decap_8 FILLER_1_1553 ();
 sg13g2_decap_8 FILLER_1_1560 ();
 sg13g2_decap_8 FILLER_1_1567 ();
 sg13g2_decap_8 FILLER_1_1574 ();
 sg13g2_decap_8 FILLER_1_1581 ();
 sg13g2_decap_8 FILLER_1_1588 ();
 sg13g2_decap_8 FILLER_1_1595 ();
 sg13g2_decap_8 FILLER_1_1602 ();
 sg13g2_decap_8 FILLER_1_1609 ();
 sg13g2_decap_8 FILLER_1_1616 ();
 sg13g2_decap_8 FILLER_1_1623 ();
 sg13g2_decap_8 FILLER_1_1630 ();
 sg13g2_decap_8 FILLER_1_1637 ();
 sg13g2_decap_8 FILLER_1_1644 ();
 sg13g2_decap_8 FILLER_1_1651 ();
 sg13g2_decap_8 FILLER_1_1658 ();
 sg13g2_decap_8 FILLER_1_1665 ();
 sg13g2_decap_8 FILLER_1_1672 ();
 sg13g2_decap_8 FILLER_1_1679 ();
 sg13g2_decap_8 FILLER_1_1686 ();
 sg13g2_decap_8 FILLER_1_1693 ();
 sg13g2_decap_8 FILLER_1_1700 ();
 sg13g2_decap_8 FILLER_1_1707 ();
 sg13g2_decap_8 FILLER_1_1714 ();
 sg13g2_decap_8 FILLER_1_1721 ();
 sg13g2_decap_8 FILLER_1_1728 ();
 sg13g2_decap_8 FILLER_1_1735 ();
 sg13g2_decap_8 FILLER_1_1742 ();
 sg13g2_decap_8 FILLER_1_1749 ();
 sg13g2_decap_8 FILLER_1_1756 ();
 sg13g2_decap_4 FILLER_1_1763 ();
 sg13g2_fill_1 FILLER_1_1767 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_fill_1 FILLER_2_539 ();
 sg13g2_fill_1 FILLER_2_561 ();
 sg13g2_fill_1 FILLER_2_589 ();
 sg13g2_fill_1 FILLER_2_598 ();
 sg13g2_fill_1 FILLER_2_617 ();
 sg13g2_fill_2 FILLER_2_639 ();
 sg13g2_fill_1 FILLER_2_641 ();
 sg13g2_fill_2 FILLER_2_663 ();
 sg13g2_fill_1 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_687 ();
 sg13g2_decap_4 FILLER_2_694 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_fill_2 FILLER_2_718 ();
 sg13g2_fill_1 FILLER_2_720 ();
 sg13g2_fill_2 FILLER_2_755 ();
 sg13g2_fill_1 FILLER_2_757 ();
 sg13g2_fill_1 FILLER_2_772 ();
 sg13g2_fill_2 FILLER_2_779 ();
 sg13g2_fill_1 FILLER_2_793 ();
 sg13g2_decap_8 FILLER_2_804 ();
 sg13g2_decap_8 FILLER_2_811 ();
 sg13g2_fill_2 FILLER_2_818 ();
 sg13g2_fill_2 FILLER_2_850 ();
 sg13g2_decap_4 FILLER_2_861 ();
 sg13g2_fill_2 FILLER_2_865 ();
 sg13g2_decap_4 FILLER_2_889 ();
 sg13g2_decap_8 FILLER_2_925 ();
 sg13g2_fill_1 FILLER_2_932 ();
 sg13g2_fill_2 FILLER_2_954 ();
 sg13g2_fill_1 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_965 ();
 sg13g2_fill_2 FILLER_2_972 ();
 sg13g2_fill_1 FILLER_2_974 ();
 sg13g2_fill_2 FILLER_2_983 ();
 sg13g2_fill_1 FILLER_2_1011 ();
 sg13g2_fill_2 FILLER_2_1033 ();
 sg13g2_fill_1 FILLER_2_1035 ();
 sg13g2_decap_8 FILLER_2_1046 ();
 sg13g2_fill_2 FILLER_2_1053 ();
 sg13g2_fill_1 FILLER_2_1055 ();
 sg13g2_decap_8 FILLER_2_1064 ();
 sg13g2_fill_2 FILLER_2_1081 ();
 sg13g2_fill_1 FILLER_2_1083 ();
 sg13g2_decap_8 FILLER_2_1090 ();
 sg13g2_decap_8 FILLER_2_1097 ();
 sg13g2_decap_8 FILLER_2_1112 ();
 sg13g2_decap_8 FILLER_2_1119 ();
 sg13g2_decap_8 FILLER_2_1126 ();
 sg13g2_decap_8 FILLER_2_1133 ();
 sg13g2_decap_8 FILLER_2_1140 ();
 sg13g2_decap_8 FILLER_2_1147 ();
 sg13g2_decap_8 FILLER_2_1154 ();
 sg13g2_decap_8 FILLER_2_1161 ();
 sg13g2_decap_8 FILLER_2_1168 ();
 sg13g2_decap_8 FILLER_2_1175 ();
 sg13g2_decap_8 FILLER_2_1182 ();
 sg13g2_decap_8 FILLER_2_1189 ();
 sg13g2_decap_8 FILLER_2_1196 ();
 sg13g2_decap_8 FILLER_2_1203 ();
 sg13g2_decap_8 FILLER_2_1210 ();
 sg13g2_decap_8 FILLER_2_1217 ();
 sg13g2_decap_8 FILLER_2_1224 ();
 sg13g2_decap_8 FILLER_2_1231 ();
 sg13g2_decap_8 FILLER_2_1238 ();
 sg13g2_decap_8 FILLER_2_1245 ();
 sg13g2_decap_8 FILLER_2_1252 ();
 sg13g2_decap_8 FILLER_2_1259 ();
 sg13g2_decap_8 FILLER_2_1266 ();
 sg13g2_decap_8 FILLER_2_1273 ();
 sg13g2_decap_8 FILLER_2_1280 ();
 sg13g2_decap_8 FILLER_2_1287 ();
 sg13g2_decap_8 FILLER_2_1294 ();
 sg13g2_decap_8 FILLER_2_1301 ();
 sg13g2_decap_8 FILLER_2_1308 ();
 sg13g2_decap_8 FILLER_2_1315 ();
 sg13g2_decap_8 FILLER_2_1322 ();
 sg13g2_decap_8 FILLER_2_1329 ();
 sg13g2_decap_8 FILLER_2_1336 ();
 sg13g2_decap_8 FILLER_2_1343 ();
 sg13g2_decap_8 FILLER_2_1350 ();
 sg13g2_decap_8 FILLER_2_1357 ();
 sg13g2_decap_8 FILLER_2_1364 ();
 sg13g2_decap_8 FILLER_2_1371 ();
 sg13g2_decap_8 FILLER_2_1378 ();
 sg13g2_decap_8 FILLER_2_1385 ();
 sg13g2_decap_8 FILLER_2_1392 ();
 sg13g2_decap_8 FILLER_2_1399 ();
 sg13g2_decap_8 FILLER_2_1406 ();
 sg13g2_decap_8 FILLER_2_1413 ();
 sg13g2_decap_8 FILLER_2_1420 ();
 sg13g2_decap_8 FILLER_2_1427 ();
 sg13g2_decap_8 FILLER_2_1434 ();
 sg13g2_decap_8 FILLER_2_1441 ();
 sg13g2_decap_8 FILLER_2_1448 ();
 sg13g2_decap_8 FILLER_2_1455 ();
 sg13g2_decap_8 FILLER_2_1462 ();
 sg13g2_decap_8 FILLER_2_1469 ();
 sg13g2_decap_8 FILLER_2_1476 ();
 sg13g2_decap_8 FILLER_2_1483 ();
 sg13g2_decap_8 FILLER_2_1490 ();
 sg13g2_decap_8 FILLER_2_1497 ();
 sg13g2_decap_8 FILLER_2_1504 ();
 sg13g2_decap_8 FILLER_2_1511 ();
 sg13g2_decap_8 FILLER_2_1518 ();
 sg13g2_decap_8 FILLER_2_1525 ();
 sg13g2_decap_8 FILLER_2_1532 ();
 sg13g2_decap_8 FILLER_2_1539 ();
 sg13g2_decap_8 FILLER_2_1546 ();
 sg13g2_decap_8 FILLER_2_1553 ();
 sg13g2_decap_8 FILLER_2_1560 ();
 sg13g2_decap_8 FILLER_2_1567 ();
 sg13g2_decap_8 FILLER_2_1574 ();
 sg13g2_decap_8 FILLER_2_1581 ();
 sg13g2_decap_8 FILLER_2_1588 ();
 sg13g2_decap_8 FILLER_2_1595 ();
 sg13g2_decap_8 FILLER_2_1602 ();
 sg13g2_decap_8 FILLER_2_1609 ();
 sg13g2_decap_8 FILLER_2_1616 ();
 sg13g2_decap_8 FILLER_2_1623 ();
 sg13g2_decap_8 FILLER_2_1630 ();
 sg13g2_decap_8 FILLER_2_1637 ();
 sg13g2_decap_8 FILLER_2_1644 ();
 sg13g2_decap_8 FILLER_2_1651 ();
 sg13g2_decap_8 FILLER_2_1658 ();
 sg13g2_decap_8 FILLER_2_1665 ();
 sg13g2_decap_8 FILLER_2_1672 ();
 sg13g2_decap_8 FILLER_2_1679 ();
 sg13g2_decap_8 FILLER_2_1686 ();
 sg13g2_decap_8 FILLER_2_1693 ();
 sg13g2_decap_8 FILLER_2_1700 ();
 sg13g2_decap_8 FILLER_2_1707 ();
 sg13g2_decap_8 FILLER_2_1714 ();
 sg13g2_decap_8 FILLER_2_1721 ();
 sg13g2_decap_8 FILLER_2_1728 ();
 sg13g2_decap_8 FILLER_2_1735 ();
 sg13g2_decap_8 FILLER_2_1742 ();
 sg13g2_decap_8 FILLER_2_1749 ();
 sg13g2_decap_8 FILLER_2_1756 ();
 sg13g2_decap_4 FILLER_2_1763 ();
 sg13g2_fill_1 FILLER_2_1767 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_fill_1 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_561 ();
 sg13g2_decap_8 FILLER_3_625 ();
 sg13g2_decap_8 FILLER_3_632 ();
 sg13g2_fill_2 FILLER_3_639 ();
 sg13g2_decap_8 FILLER_3_662 ();
 sg13g2_decap_4 FILLER_3_669 ();
 sg13g2_decap_8 FILLER_3_694 ();
 sg13g2_decap_8 FILLER_3_701 ();
 sg13g2_decap_8 FILLER_3_723 ();
 sg13g2_decap_8 FILLER_3_730 ();
 sg13g2_fill_2 FILLER_3_737 ();
 sg13g2_fill_1 FILLER_3_766 ();
 sg13g2_fill_1 FILLER_3_775 ();
 sg13g2_decap_8 FILLER_3_785 ();
 sg13g2_fill_2 FILLER_3_792 ();
 sg13g2_fill_1 FILLER_3_794 ();
 sg13g2_decap_4 FILLER_3_816 ();
 sg13g2_fill_2 FILLER_3_820 ();
 sg13g2_decap_8 FILLER_3_830 ();
 sg13g2_decap_8 FILLER_3_843 ();
 sg13g2_fill_2 FILLER_3_854 ();
 sg13g2_fill_2 FILLER_3_872 ();
 sg13g2_decap_4 FILLER_3_895 ();
 sg13g2_fill_2 FILLER_3_920 ();
 sg13g2_fill_1 FILLER_3_922 ();
 sg13g2_fill_2 FILLER_3_946 ();
 sg13g2_fill_2 FILLER_3_979 ();
 sg13g2_fill_1 FILLER_3_999 ();
 sg13g2_fill_2 FILLER_3_1054 ();
 sg13g2_decap_4 FILLER_3_1077 ();
 sg13g2_decap_4 FILLER_3_1103 ();
 sg13g2_fill_1 FILLER_3_1107 ();
 sg13g2_decap_8 FILLER_3_1118 ();
 sg13g2_decap_8 FILLER_3_1125 ();
 sg13g2_decap_8 FILLER_3_1132 ();
 sg13g2_decap_8 FILLER_3_1139 ();
 sg13g2_decap_8 FILLER_3_1146 ();
 sg13g2_decap_8 FILLER_3_1153 ();
 sg13g2_decap_8 FILLER_3_1160 ();
 sg13g2_decap_8 FILLER_3_1167 ();
 sg13g2_decap_8 FILLER_3_1174 ();
 sg13g2_decap_8 FILLER_3_1181 ();
 sg13g2_decap_8 FILLER_3_1188 ();
 sg13g2_decap_8 FILLER_3_1195 ();
 sg13g2_decap_8 FILLER_3_1202 ();
 sg13g2_decap_8 FILLER_3_1209 ();
 sg13g2_decap_8 FILLER_3_1216 ();
 sg13g2_decap_8 FILLER_3_1223 ();
 sg13g2_decap_8 FILLER_3_1230 ();
 sg13g2_decap_8 FILLER_3_1237 ();
 sg13g2_decap_8 FILLER_3_1244 ();
 sg13g2_decap_8 FILLER_3_1251 ();
 sg13g2_decap_8 FILLER_3_1258 ();
 sg13g2_decap_8 FILLER_3_1265 ();
 sg13g2_decap_8 FILLER_3_1272 ();
 sg13g2_decap_8 FILLER_3_1279 ();
 sg13g2_decap_8 FILLER_3_1286 ();
 sg13g2_decap_8 FILLER_3_1293 ();
 sg13g2_decap_8 FILLER_3_1300 ();
 sg13g2_decap_8 FILLER_3_1307 ();
 sg13g2_decap_8 FILLER_3_1314 ();
 sg13g2_decap_8 FILLER_3_1321 ();
 sg13g2_decap_8 FILLER_3_1328 ();
 sg13g2_decap_8 FILLER_3_1335 ();
 sg13g2_decap_8 FILLER_3_1342 ();
 sg13g2_decap_8 FILLER_3_1349 ();
 sg13g2_decap_8 FILLER_3_1356 ();
 sg13g2_decap_8 FILLER_3_1363 ();
 sg13g2_decap_8 FILLER_3_1370 ();
 sg13g2_decap_8 FILLER_3_1377 ();
 sg13g2_decap_8 FILLER_3_1384 ();
 sg13g2_decap_8 FILLER_3_1391 ();
 sg13g2_decap_8 FILLER_3_1398 ();
 sg13g2_decap_8 FILLER_3_1405 ();
 sg13g2_decap_8 FILLER_3_1412 ();
 sg13g2_decap_8 FILLER_3_1419 ();
 sg13g2_decap_8 FILLER_3_1426 ();
 sg13g2_decap_8 FILLER_3_1433 ();
 sg13g2_decap_8 FILLER_3_1440 ();
 sg13g2_decap_8 FILLER_3_1447 ();
 sg13g2_decap_8 FILLER_3_1454 ();
 sg13g2_decap_8 FILLER_3_1461 ();
 sg13g2_decap_8 FILLER_3_1468 ();
 sg13g2_decap_8 FILLER_3_1475 ();
 sg13g2_decap_8 FILLER_3_1482 ();
 sg13g2_decap_8 FILLER_3_1489 ();
 sg13g2_decap_8 FILLER_3_1496 ();
 sg13g2_decap_8 FILLER_3_1503 ();
 sg13g2_decap_8 FILLER_3_1510 ();
 sg13g2_decap_8 FILLER_3_1517 ();
 sg13g2_decap_8 FILLER_3_1524 ();
 sg13g2_decap_8 FILLER_3_1531 ();
 sg13g2_decap_8 FILLER_3_1538 ();
 sg13g2_decap_8 FILLER_3_1545 ();
 sg13g2_decap_8 FILLER_3_1552 ();
 sg13g2_decap_8 FILLER_3_1559 ();
 sg13g2_decap_8 FILLER_3_1566 ();
 sg13g2_decap_8 FILLER_3_1573 ();
 sg13g2_decap_8 FILLER_3_1580 ();
 sg13g2_decap_8 FILLER_3_1587 ();
 sg13g2_decap_8 FILLER_3_1594 ();
 sg13g2_decap_8 FILLER_3_1601 ();
 sg13g2_decap_8 FILLER_3_1608 ();
 sg13g2_decap_8 FILLER_3_1615 ();
 sg13g2_decap_8 FILLER_3_1622 ();
 sg13g2_decap_8 FILLER_3_1629 ();
 sg13g2_decap_8 FILLER_3_1636 ();
 sg13g2_decap_8 FILLER_3_1643 ();
 sg13g2_decap_8 FILLER_3_1650 ();
 sg13g2_decap_8 FILLER_3_1657 ();
 sg13g2_decap_8 FILLER_3_1664 ();
 sg13g2_decap_8 FILLER_3_1671 ();
 sg13g2_decap_8 FILLER_3_1678 ();
 sg13g2_decap_8 FILLER_3_1685 ();
 sg13g2_decap_8 FILLER_3_1692 ();
 sg13g2_decap_8 FILLER_3_1699 ();
 sg13g2_decap_8 FILLER_3_1706 ();
 sg13g2_decap_8 FILLER_3_1713 ();
 sg13g2_decap_8 FILLER_3_1720 ();
 sg13g2_decap_8 FILLER_3_1727 ();
 sg13g2_decap_8 FILLER_3_1734 ();
 sg13g2_decap_8 FILLER_3_1741 ();
 sg13g2_decap_8 FILLER_3_1748 ();
 sg13g2_decap_8 FILLER_3_1755 ();
 sg13g2_decap_4 FILLER_3_1762 ();
 sg13g2_fill_2 FILLER_3_1766 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_fill_2 FILLER_4_287 ();
 sg13g2_fill_1 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_4 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_309 ();
 sg13g2_fill_1 FILLER_4_316 ();
 sg13g2_decap_8 FILLER_4_321 ();
 sg13g2_decap_8 FILLER_4_328 ();
 sg13g2_decap_8 FILLER_4_335 ();
 sg13g2_decap_8 FILLER_4_342 ();
 sg13g2_decap_8 FILLER_4_349 ();
 sg13g2_decap_4 FILLER_4_356 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_8 FILLER_4_430 ();
 sg13g2_decap_8 FILLER_4_437 ();
 sg13g2_decap_8 FILLER_4_444 ();
 sg13g2_decap_8 FILLER_4_451 ();
 sg13g2_decap_8 FILLER_4_458 ();
 sg13g2_decap_8 FILLER_4_465 ();
 sg13g2_decap_8 FILLER_4_472 ();
 sg13g2_decap_8 FILLER_4_479 ();
 sg13g2_decap_8 FILLER_4_486 ();
 sg13g2_decap_8 FILLER_4_493 ();
 sg13g2_decap_8 FILLER_4_500 ();
 sg13g2_decap_8 FILLER_4_507 ();
 sg13g2_decap_8 FILLER_4_514 ();
 sg13g2_decap_8 FILLER_4_521 ();
 sg13g2_decap_4 FILLER_4_528 ();
 sg13g2_fill_1 FILLER_4_532 ();
 sg13g2_decap_4 FILLER_4_545 ();
 sg13g2_decap_8 FILLER_4_559 ();
 sg13g2_decap_4 FILLER_4_566 ();
 sg13g2_fill_2 FILLER_4_570 ();
 sg13g2_decap_4 FILLER_4_596 ();
 sg13g2_decap_4 FILLER_4_608 ();
 sg13g2_decap_8 FILLER_4_627 ();
 sg13g2_decap_8 FILLER_4_634 ();
 sg13g2_fill_1 FILLER_4_641 ();
 sg13g2_fill_1 FILLER_4_663 ();
 sg13g2_fill_2 FILLER_4_711 ();
 sg13g2_fill_1 FILLER_4_713 ();
 sg13g2_decap_4 FILLER_4_735 ();
 sg13g2_fill_1 FILLER_4_739 ();
 sg13g2_decap_4 FILLER_4_762 ();
 sg13g2_fill_1 FILLER_4_766 ();
 sg13g2_fill_1 FILLER_4_777 ();
 sg13g2_fill_2 FILLER_4_794 ();
 sg13g2_fill_2 FILLER_4_832 ();
 sg13g2_fill_1 FILLER_4_834 ();
 sg13g2_fill_1 FILLER_4_851 ();
 sg13g2_fill_2 FILLER_4_870 ();
 sg13g2_fill_1 FILLER_4_893 ();
 sg13g2_fill_2 FILLER_4_923 ();
 sg13g2_fill_2 FILLER_4_954 ();
 sg13g2_fill_1 FILLER_4_956 ();
 sg13g2_fill_2 FILLER_4_978 ();
 sg13g2_fill_1 FILLER_4_980 ();
 sg13g2_fill_2 FILLER_4_998 ();
 sg13g2_fill_1 FILLER_4_1000 ();
 sg13g2_decap_8 FILLER_4_1016 ();
 sg13g2_decap_8 FILLER_4_1023 ();
 sg13g2_decap_4 FILLER_4_1030 ();
 sg13g2_fill_2 FILLER_4_1034 ();
 sg13g2_decap_8 FILLER_4_1042 ();
 sg13g2_decap_8 FILLER_4_1070 ();
 sg13g2_fill_1 FILLER_4_1077 ();
 sg13g2_fill_1 FILLER_4_1090 ();
 sg13g2_decap_8 FILLER_4_1122 ();
 sg13g2_decap_8 FILLER_4_1129 ();
 sg13g2_decap_8 FILLER_4_1136 ();
 sg13g2_decap_8 FILLER_4_1143 ();
 sg13g2_decap_8 FILLER_4_1150 ();
 sg13g2_decap_8 FILLER_4_1157 ();
 sg13g2_decap_8 FILLER_4_1164 ();
 sg13g2_decap_8 FILLER_4_1171 ();
 sg13g2_decap_8 FILLER_4_1178 ();
 sg13g2_decap_8 FILLER_4_1185 ();
 sg13g2_decap_8 FILLER_4_1192 ();
 sg13g2_decap_8 FILLER_4_1199 ();
 sg13g2_decap_8 FILLER_4_1206 ();
 sg13g2_decap_8 FILLER_4_1213 ();
 sg13g2_decap_8 FILLER_4_1220 ();
 sg13g2_decap_8 FILLER_4_1227 ();
 sg13g2_decap_8 FILLER_4_1234 ();
 sg13g2_decap_8 FILLER_4_1241 ();
 sg13g2_decap_8 FILLER_4_1248 ();
 sg13g2_decap_8 FILLER_4_1255 ();
 sg13g2_decap_8 FILLER_4_1262 ();
 sg13g2_decap_8 FILLER_4_1269 ();
 sg13g2_decap_8 FILLER_4_1276 ();
 sg13g2_decap_8 FILLER_4_1283 ();
 sg13g2_decap_8 FILLER_4_1290 ();
 sg13g2_decap_8 FILLER_4_1297 ();
 sg13g2_decap_8 FILLER_4_1304 ();
 sg13g2_decap_8 FILLER_4_1311 ();
 sg13g2_decap_8 FILLER_4_1318 ();
 sg13g2_decap_8 FILLER_4_1325 ();
 sg13g2_decap_8 FILLER_4_1332 ();
 sg13g2_decap_8 FILLER_4_1339 ();
 sg13g2_decap_8 FILLER_4_1346 ();
 sg13g2_decap_8 FILLER_4_1353 ();
 sg13g2_decap_8 FILLER_4_1360 ();
 sg13g2_decap_8 FILLER_4_1367 ();
 sg13g2_decap_8 FILLER_4_1374 ();
 sg13g2_decap_8 FILLER_4_1381 ();
 sg13g2_decap_8 FILLER_4_1388 ();
 sg13g2_decap_8 FILLER_4_1395 ();
 sg13g2_decap_8 FILLER_4_1402 ();
 sg13g2_decap_8 FILLER_4_1409 ();
 sg13g2_decap_8 FILLER_4_1416 ();
 sg13g2_decap_8 FILLER_4_1423 ();
 sg13g2_decap_8 FILLER_4_1430 ();
 sg13g2_decap_8 FILLER_4_1437 ();
 sg13g2_decap_8 FILLER_4_1444 ();
 sg13g2_decap_8 FILLER_4_1451 ();
 sg13g2_decap_8 FILLER_4_1458 ();
 sg13g2_decap_8 FILLER_4_1465 ();
 sg13g2_decap_8 FILLER_4_1472 ();
 sg13g2_decap_8 FILLER_4_1479 ();
 sg13g2_decap_8 FILLER_4_1486 ();
 sg13g2_decap_8 FILLER_4_1493 ();
 sg13g2_decap_8 FILLER_4_1500 ();
 sg13g2_decap_8 FILLER_4_1507 ();
 sg13g2_decap_8 FILLER_4_1514 ();
 sg13g2_decap_8 FILLER_4_1521 ();
 sg13g2_decap_8 FILLER_4_1528 ();
 sg13g2_decap_8 FILLER_4_1535 ();
 sg13g2_decap_8 FILLER_4_1542 ();
 sg13g2_decap_8 FILLER_4_1549 ();
 sg13g2_decap_8 FILLER_4_1556 ();
 sg13g2_decap_8 FILLER_4_1563 ();
 sg13g2_decap_8 FILLER_4_1570 ();
 sg13g2_decap_8 FILLER_4_1577 ();
 sg13g2_decap_8 FILLER_4_1584 ();
 sg13g2_decap_8 FILLER_4_1591 ();
 sg13g2_decap_8 FILLER_4_1598 ();
 sg13g2_decap_8 FILLER_4_1605 ();
 sg13g2_decap_8 FILLER_4_1612 ();
 sg13g2_decap_8 FILLER_4_1619 ();
 sg13g2_decap_8 FILLER_4_1626 ();
 sg13g2_decap_8 FILLER_4_1633 ();
 sg13g2_decap_8 FILLER_4_1640 ();
 sg13g2_decap_8 FILLER_4_1647 ();
 sg13g2_decap_8 FILLER_4_1654 ();
 sg13g2_decap_8 FILLER_4_1661 ();
 sg13g2_decap_8 FILLER_4_1668 ();
 sg13g2_decap_8 FILLER_4_1675 ();
 sg13g2_decap_8 FILLER_4_1682 ();
 sg13g2_decap_8 FILLER_4_1689 ();
 sg13g2_decap_8 FILLER_4_1696 ();
 sg13g2_decap_8 FILLER_4_1703 ();
 sg13g2_decap_8 FILLER_4_1710 ();
 sg13g2_decap_8 FILLER_4_1717 ();
 sg13g2_decap_8 FILLER_4_1724 ();
 sg13g2_decap_8 FILLER_4_1731 ();
 sg13g2_decap_8 FILLER_4_1738 ();
 sg13g2_decap_8 FILLER_4_1745 ();
 sg13g2_decap_8 FILLER_4_1752 ();
 sg13g2_decap_8 FILLER_4_1759 ();
 sg13g2_fill_2 FILLER_4_1766 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_4 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_202 ();
 sg13g2_decap_4 FILLER_5_209 ();
 sg13g2_fill_1 FILLER_5_213 ();
 sg13g2_decap_8 FILLER_5_227 ();
 sg13g2_decap_8 FILLER_5_234 ();
 sg13g2_fill_2 FILLER_5_241 ();
 sg13g2_decap_8 FILLER_5_258 ();
 sg13g2_decap_8 FILLER_5_265 ();
 sg13g2_decap_4 FILLER_5_276 ();
 sg13g2_fill_1 FILLER_5_280 ();
 sg13g2_fill_2 FILLER_5_312 ();
 sg13g2_fill_1 FILLER_5_314 ();
 sg13g2_decap_4 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_418 ();
 sg13g2_decap_8 FILLER_5_425 ();
 sg13g2_fill_2 FILLER_5_432 ();
 sg13g2_fill_2 FILLER_5_439 ();
 sg13g2_fill_1 FILLER_5_445 ();
 sg13g2_decap_8 FILLER_5_472 ();
 sg13g2_decap_8 FILLER_5_479 ();
 sg13g2_fill_2 FILLER_5_486 ();
 sg13g2_fill_1 FILLER_5_488 ();
 sg13g2_decap_8 FILLER_5_493 ();
 sg13g2_fill_2 FILLER_5_500 ();
 sg13g2_fill_1 FILLER_5_502 ();
 sg13g2_decap_8 FILLER_5_512 ();
 sg13g2_decap_8 FILLER_5_519 ();
 sg13g2_fill_1 FILLER_5_526 ();
 sg13g2_fill_1 FILLER_5_579 ();
 sg13g2_decap_4 FILLER_5_601 ();
 sg13g2_fill_1 FILLER_5_605 ();
 sg13g2_fill_1 FILLER_5_629 ();
 sg13g2_decap_4 FILLER_5_651 ();
 sg13g2_fill_2 FILLER_5_672 ();
 sg13g2_fill_2 FILLER_5_678 ();
 sg13g2_decap_4 FILLER_5_691 ();
 sg13g2_fill_1 FILLER_5_713 ();
 sg13g2_decap_8 FILLER_5_718 ();
 sg13g2_decap_4 FILLER_5_730 ();
 sg13g2_decap_4 FILLER_5_752 ();
 sg13g2_decap_8 FILLER_5_792 ();
 sg13g2_fill_1 FILLER_5_799 ();
 sg13g2_decap_8 FILLER_5_829 ();
 sg13g2_fill_2 FILLER_5_836 ();
 sg13g2_fill_1 FILLER_5_838 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_4 FILLER_5_858 ();
 sg13g2_fill_1 FILLER_5_862 ();
 sg13g2_decap_8 FILLER_5_868 ();
 sg13g2_fill_1 FILLER_5_903 ();
 sg13g2_fill_2 FILLER_5_915 ();
 sg13g2_fill_1 FILLER_5_917 ();
 sg13g2_decap_4 FILLER_5_940 ();
 sg13g2_fill_1 FILLER_5_944 ();
 sg13g2_decap_8 FILLER_5_955 ();
 sg13g2_decap_8 FILLER_5_962 ();
 sg13g2_decap_8 FILLER_5_974 ();
 sg13g2_decap_8 FILLER_5_981 ();
 sg13g2_fill_1 FILLER_5_988 ();
 sg13g2_fill_2 FILLER_5_998 ();
 sg13g2_fill_1 FILLER_5_1000 ();
 sg13g2_fill_1 FILLER_5_1016 ();
 sg13g2_fill_2 FILLER_5_1025 ();
 sg13g2_decap_8 FILLER_5_1048 ();
 sg13g2_decap_8 FILLER_5_1055 ();
 sg13g2_fill_2 FILLER_5_1062 ();
 sg13g2_fill_1 FILLER_5_1064 ();
 sg13g2_decap_4 FILLER_5_1075 ();
 sg13g2_decap_8 FILLER_5_1110 ();
 sg13g2_decap_4 FILLER_5_1117 ();
 sg13g2_fill_2 FILLER_5_1121 ();
 sg13g2_decap_8 FILLER_5_1131 ();
 sg13g2_decap_8 FILLER_5_1138 ();
 sg13g2_decap_8 FILLER_5_1145 ();
 sg13g2_decap_8 FILLER_5_1152 ();
 sg13g2_decap_8 FILLER_5_1159 ();
 sg13g2_decap_8 FILLER_5_1166 ();
 sg13g2_decap_8 FILLER_5_1173 ();
 sg13g2_decap_8 FILLER_5_1180 ();
 sg13g2_decap_8 FILLER_5_1187 ();
 sg13g2_decap_8 FILLER_5_1194 ();
 sg13g2_decap_8 FILLER_5_1201 ();
 sg13g2_decap_8 FILLER_5_1208 ();
 sg13g2_decap_8 FILLER_5_1215 ();
 sg13g2_decap_8 FILLER_5_1222 ();
 sg13g2_decap_8 FILLER_5_1229 ();
 sg13g2_decap_8 FILLER_5_1236 ();
 sg13g2_decap_8 FILLER_5_1243 ();
 sg13g2_decap_8 FILLER_5_1250 ();
 sg13g2_decap_8 FILLER_5_1257 ();
 sg13g2_decap_8 FILLER_5_1264 ();
 sg13g2_decap_8 FILLER_5_1271 ();
 sg13g2_decap_8 FILLER_5_1278 ();
 sg13g2_decap_8 FILLER_5_1285 ();
 sg13g2_decap_8 FILLER_5_1292 ();
 sg13g2_decap_8 FILLER_5_1299 ();
 sg13g2_decap_8 FILLER_5_1306 ();
 sg13g2_decap_8 FILLER_5_1313 ();
 sg13g2_decap_8 FILLER_5_1320 ();
 sg13g2_decap_8 FILLER_5_1327 ();
 sg13g2_decap_8 FILLER_5_1334 ();
 sg13g2_decap_8 FILLER_5_1341 ();
 sg13g2_decap_8 FILLER_5_1348 ();
 sg13g2_decap_8 FILLER_5_1355 ();
 sg13g2_decap_8 FILLER_5_1362 ();
 sg13g2_decap_8 FILLER_5_1369 ();
 sg13g2_decap_8 FILLER_5_1376 ();
 sg13g2_decap_8 FILLER_5_1383 ();
 sg13g2_decap_8 FILLER_5_1390 ();
 sg13g2_decap_8 FILLER_5_1397 ();
 sg13g2_decap_8 FILLER_5_1404 ();
 sg13g2_decap_8 FILLER_5_1411 ();
 sg13g2_decap_8 FILLER_5_1418 ();
 sg13g2_decap_8 FILLER_5_1425 ();
 sg13g2_decap_8 FILLER_5_1432 ();
 sg13g2_decap_8 FILLER_5_1439 ();
 sg13g2_decap_8 FILLER_5_1446 ();
 sg13g2_decap_8 FILLER_5_1453 ();
 sg13g2_decap_8 FILLER_5_1460 ();
 sg13g2_decap_8 FILLER_5_1467 ();
 sg13g2_decap_8 FILLER_5_1474 ();
 sg13g2_decap_8 FILLER_5_1481 ();
 sg13g2_decap_8 FILLER_5_1488 ();
 sg13g2_decap_8 FILLER_5_1495 ();
 sg13g2_decap_8 FILLER_5_1502 ();
 sg13g2_decap_8 FILLER_5_1509 ();
 sg13g2_decap_8 FILLER_5_1516 ();
 sg13g2_decap_8 FILLER_5_1523 ();
 sg13g2_decap_8 FILLER_5_1530 ();
 sg13g2_decap_8 FILLER_5_1537 ();
 sg13g2_decap_8 FILLER_5_1544 ();
 sg13g2_decap_8 FILLER_5_1551 ();
 sg13g2_decap_8 FILLER_5_1558 ();
 sg13g2_decap_8 FILLER_5_1565 ();
 sg13g2_decap_8 FILLER_5_1572 ();
 sg13g2_decap_8 FILLER_5_1579 ();
 sg13g2_decap_8 FILLER_5_1586 ();
 sg13g2_decap_8 FILLER_5_1593 ();
 sg13g2_decap_8 FILLER_5_1600 ();
 sg13g2_decap_8 FILLER_5_1607 ();
 sg13g2_decap_8 FILLER_5_1614 ();
 sg13g2_decap_8 FILLER_5_1621 ();
 sg13g2_decap_8 FILLER_5_1628 ();
 sg13g2_decap_8 FILLER_5_1635 ();
 sg13g2_decap_8 FILLER_5_1642 ();
 sg13g2_decap_8 FILLER_5_1649 ();
 sg13g2_decap_8 FILLER_5_1656 ();
 sg13g2_decap_8 FILLER_5_1663 ();
 sg13g2_decap_8 FILLER_5_1670 ();
 sg13g2_decap_8 FILLER_5_1677 ();
 sg13g2_decap_8 FILLER_5_1684 ();
 sg13g2_decap_8 FILLER_5_1691 ();
 sg13g2_decap_8 FILLER_5_1698 ();
 sg13g2_decap_8 FILLER_5_1705 ();
 sg13g2_decap_8 FILLER_5_1712 ();
 sg13g2_decap_8 FILLER_5_1719 ();
 sg13g2_decap_8 FILLER_5_1726 ();
 sg13g2_decap_8 FILLER_5_1733 ();
 sg13g2_decap_8 FILLER_5_1740 ();
 sg13g2_decap_8 FILLER_5_1747 ();
 sg13g2_decap_8 FILLER_5_1754 ();
 sg13g2_decap_8 FILLER_5_1761 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_fill_2 FILLER_6_154 ();
 sg13g2_fill_2 FILLER_6_165 ();
 sg13g2_fill_1 FILLER_6_245 ();
 sg13g2_fill_2 FILLER_6_294 ();
 sg13g2_fill_2 FILLER_6_319 ();
 sg13g2_fill_1 FILLER_6_321 ();
 sg13g2_fill_2 FILLER_6_365 ();
 sg13g2_fill_1 FILLER_6_367 ();
 sg13g2_fill_2 FILLER_6_443 ();
 sg13g2_decap_4 FILLER_6_476 ();
 sg13g2_fill_1 FILLER_6_519 ();
 sg13g2_decap_4 FILLER_6_544 ();
 sg13g2_fill_1 FILLER_6_548 ();
 sg13g2_decap_4 FILLER_6_563 ();
 sg13g2_fill_1 FILLER_6_567 ();
 sg13g2_decap_4 FILLER_6_589 ();
 sg13g2_fill_1 FILLER_6_593 ();
 sg13g2_decap_8 FILLER_6_646 ();
 sg13g2_fill_1 FILLER_6_653 ();
 sg13g2_fill_1 FILLER_6_676 ();
 sg13g2_fill_2 FILLER_6_685 ();
 sg13g2_fill_1 FILLER_6_687 ();
 sg13g2_decap_4 FILLER_6_713 ();
 sg13g2_fill_1 FILLER_6_717 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_fill_2 FILLER_6_746 ();
 sg13g2_fill_1 FILLER_6_748 ();
 sg13g2_decap_4 FILLER_6_772 ();
 sg13g2_fill_1 FILLER_6_776 ();
 sg13g2_fill_2 FILLER_6_798 ();
 sg13g2_fill_1 FILLER_6_800 ();
 sg13g2_fill_2 FILLER_6_829 ();
 sg13g2_fill_2 FILLER_6_849 ();
 sg13g2_fill_1 FILLER_6_851 ();
 sg13g2_fill_2 FILLER_6_865 ();
 sg13g2_fill_1 FILLER_6_867 ();
 sg13g2_decap_8 FILLER_6_878 ();
 sg13g2_decap_8 FILLER_6_885 ();
 sg13g2_fill_2 FILLER_6_892 ();
 sg13g2_decap_8 FILLER_6_904 ();
 sg13g2_fill_2 FILLER_6_911 ();
 sg13g2_decap_4 FILLER_6_934 ();
 sg13g2_decap_8 FILLER_6_958 ();
 sg13g2_fill_2 FILLER_6_965 ();
 sg13g2_fill_1 FILLER_6_967 ();
 sg13g2_decap_4 FILLER_6_991 ();
 sg13g2_fill_2 FILLER_6_995 ();
 sg13g2_fill_2 FILLER_6_1007 ();
 sg13g2_fill_1 FILLER_6_1009 ();
 sg13g2_decap_8 FILLER_6_1030 ();
 sg13g2_fill_2 FILLER_6_1058 ();
 sg13g2_decap_4 FILLER_6_1070 ();
 sg13g2_decap_8 FILLER_6_1100 ();
 sg13g2_fill_2 FILLER_6_1107 ();
 sg13g2_decap_8 FILLER_6_1130 ();
 sg13g2_decap_8 FILLER_6_1137 ();
 sg13g2_decap_8 FILLER_6_1144 ();
 sg13g2_decap_8 FILLER_6_1151 ();
 sg13g2_decap_8 FILLER_6_1158 ();
 sg13g2_decap_8 FILLER_6_1165 ();
 sg13g2_decap_8 FILLER_6_1172 ();
 sg13g2_decap_8 FILLER_6_1179 ();
 sg13g2_decap_8 FILLER_6_1186 ();
 sg13g2_decap_8 FILLER_6_1193 ();
 sg13g2_decap_8 FILLER_6_1200 ();
 sg13g2_decap_8 FILLER_6_1207 ();
 sg13g2_decap_8 FILLER_6_1214 ();
 sg13g2_decap_8 FILLER_6_1221 ();
 sg13g2_decap_8 FILLER_6_1228 ();
 sg13g2_decap_8 FILLER_6_1235 ();
 sg13g2_decap_8 FILLER_6_1242 ();
 sg13g2_decap_8 FILLER_6_1249 ();
 sg13g2_decap_8 FILLER_6_1256 ();
 sg13g2_decap_8 FILLER_6_1263 ();
 sg13g2_decap_8 FILLER_6_1270 ();
 sg13g2_decap_8 FILLER_6_1277 ();
 sg13g2_decap_8 FILLER_6_1284 ();
 sg13g2_decap_8 FILLER_6_1291 ();
 sg13g2_decap_8 FILLER_6_1298 ();
 sg13g2_decap_8 FILLER_6_1305 ();
 sg13g2_decap_8 FILLER_6_1312 ();
 sg13g2_decap_8 FILLER_6_1319 ();
 sg13g2_decap_8 FILLER_6_1326 ();
 sg13g2_decap_8 FILLER_6_1333 ();
 sg13g2_decap_8 FILLER_6_1340 ();
 sg13g2_decap_8 FILLER_6_1347 ();
 sg13g2_decap_8 FILLER_6_1354 ();
 sg13g2_decap_8 FILLER_6_1361 ();
 sg13g2_decap_8 FILLER_6_1368 ();
 sg13g2_decap_8 FILLER_6_1375 ();
 sg13g2_decap_8 FILLER_6_1382 ();
 sg13g2_decap_8 FILLER_6_1389 ();
 sg13g2_decap_8 FILLER_6_1396 ();
 sg13g2_decap_8 FILLER_6_1403 ();
 sg13g2_decap_8 FILLER_6_1410 ();
 sg13g2_decap_8 FILLER_6_1417 ();
 sg13g2_decap_8 FILLER_6_1424 ();
 sg13g2_decap_8 FILLER_6_1431 ();
 sg13g2_decap_8 FILLER_6_1438 ();
 sg13g2_decap_8 FILLER_6_1445 ();
 sg13g2_decap_8 FILLER_6_1452 ();
 sg13g2_decap_8 FILLER_6_1459 ();
 sg13g2_decap_8 FILLER_6_1466 ();
 sg13g2_decap_8 FILLER_6_1473 ();
 sg13g2_decap_8 FILLER_6_1480 ();
 sg13g2_decap_8 FILLER_6_1487 ();
 sg13g2_decap_8 FILLER_6_1494 ();
 sg13g2_decap_8 FILLER_6_1501 ();
 sg13g2_decap_8 FILLER_6_1508 ();
 sg13g2_decap_8 FILLER_6_1515 ();
 sg13g2_decap_8 FILLER_6_1522 ();
 sg13g2_decap_8 FILLER_6_1529 ();
 sg13g2_decap_8 FILLER_6_1536 ();
 sg13g2_decap_8 FILLER_6_1543 ();
 sg13g2_decap_8 FILLER_6_1550 ();
 sg13g2_decap_8 FILLER_6_1557 ();
 sg13g2_decap_8 FILLER_6_1564 ();
 sg13g2_decap_8 FILLER_6_1571 ();
 sg13g2_decap_8 FILLER_6_1578 ();
 sg13g2_decap_8 FILLER_6_1585 ();
 sg13g2_decap_8 FILLER_6_1592 ();
 sg13g2_decap_8 FILLER_6_1599 ();
 sg13g2_decap_8 FILLER_6_1606 ();
 sg13g2_decap_8 FILLER_6_1613 ();
 sg13g2_decap_8 FILLER_6_1620 ();
 sg13g2_decap_8 FILLER_6_1627 ();
 sg13g2_decap_8 FILLER_6_1634 ();
 sg13g2_decap_8 FILLER_6_1641 ();
 sg13g2_decap_8 FILLER_6_1648 ();
 sg13g2_decap_8 FILLER_6_1655 ();
 sg13g2_decap_8 FILLER_6_1662 ();
 sg13g2_decap_8 FILLER_6_1669 ();
 sg13g2_decap_8 FILLER_6_1676 ();
 sg13g2_decap_8 FILLER_6_1683 ();
 sg13g2_decap_8 FILLER_6_1690 ();
 sg13g2_decap_8 FILLER_6_1697 ();
 sg13g2_decap_8 FILLER_6_1704 ();
 sg13g2_decap_8 FILLER_6_1711 ();
 sg13g2_decap_8 FILLER_6_1718 ();
 sg13g2_decap_8 FILLER_6_1725 ();
 sg13g2_decap_8 FILLER_6_1732 ();
 sg13g2_decap_8 FILLER_6_1739 ();
 sg13g2_decap_8 FILLER_6_1746 ();
 sg13g2_decap_8 FILLER_6_1753 ();
 sg13g2_decap_8 FILLER_6_1760 ();
 sg13g2_fill_1 FILLER_6_1767 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_fill_2 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_fill_1 FILLER_7_190 ();
 sg13g2_fill_1 FILLER_7_204 ();
 sg13g2_fill_2 FILLER_7_210 ();
 sg13g2_fill_2 FILLER_7_267 ();
 sg13g2_fill_1 FILLER_7_269 ();
 sg13g2_fill_2 FILLER_7_327 ();
 sg13g2_fill_2 FILLER_7_348 ();
 sg13g2_fill_1 FILLER_7_382 ();
 sg13g2_fill_2 FILLER_7_392 ();
 sg13g2_fill_1 FILLER_7_394 ();
 sg13g2_fill_1 FILLER_7_430 ();
 sg13g2_fill_2 FILLER_7_436 ();
 sg13g2_fill_1 FILLER_7_438 ();
 sg13g2_fill_2 FILLER_7_507 ();
 sg13g2_fill_1 FILLER_7_509 ();
 sg13g2_decap_4 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_fill_2 FILLER_7_616 ();
 sg13g2_fill_1 FILLER_7_618 ();
 sg13g2_decap_4 FILLER_7_631 ();
 sg13g2_fill_1 FILLER_7_635 ();
 sg13g2_decap_4 FILLER_7_657 ();
 sg13g2_fill_1 FILLER_7_661 ();
 sg13g2_fill_1 FILLER_7_676 ();
 sg13g2_fill_1 FILLER_7_681 ();
 sg13g2_decap_4 FILLER_7_687 ();
 sg13g2_fill_1 FILLER_7_706 ();
 sg13g2_fill_2 FILLER_7_713 ();
 sg13g2_fill_2 FILLER_7_734 ();
 sg13g2_fill_2 FILLER_7_746 ();
 sg13g2_decap_8 FILLER_7_764 ();
 sg13g2_decap_8 FILLER_7_771 ();
 sg13g2_fill_1 FILLER_7_778 ();
 sg13g2_decap_8 FILLER_7_789 ();
 sg13g2_decap_8 FILLER_7_796 ();
 sg13g2_fill_1 FILLER_7_803 ();
 sg13g2_fill_2 FILLER_7_811 ();
 sg13g2_fill_1 FILLER_7_818 ();
 sg13g2_fill_2 FILLER_7_843 ();
 sg13g2_fill_2 FILLER_7_855 ();
 sg13g2_decap_8 FILLER_7_875 ();
 sg13g2_decap_8 FILLER_7_882 ();
 sg13g2_decap_4 FILLER_7_889 ();
 sg13g2_decap_8 FILLER_7_908 ();
 sg13g2_fill_2 FILLER_7_915 ();
 sg13g2_fill_1 FILLER_7_917 ();
 sg13g2_decap_4 FILLER_7_928 ();
 sg13g2_fill_1 FILLER_7_932 ();
 sg13g2_decap_8 FILLER_7_937 ();
 sg13g2_fill_1 FILLER_7_944 ();
 sg13g2_fill_2 FILLER_7_949 ();
 sg13g2_decap_8 FILLER_7_977 ();
 sg13g2_decap_4 FILLER_7_984 ();
 sg13g2_fill_1 FILLER_7_1063 ();
 sg13g2_decap_4 FILLER_7_1095 ();
 sg13g2_fill_1 FILLER_7_1099 ();
 sg13g2_fill_2 FILLER_7_1105 ();
 sg13g2_decap_8 FILLER_7_1136 ();
 sg13g2_decap_8 FILLER_7_1143 ();
 sg13g2_decap_8 FILLER_7_1150 ();
 sg13g2_decap_8 FILLER_7_1157 ();
 sg13g2_decap_8 FILLER_7_1164 ();
 sg13g2_decap_8 FILLER_7_1171 ();
 sg13g2_decap_8 FILLER_7_1178 ();
 sg13g2_decap_8 FILLER_7_1185 ();
 sg13g2_decap_8 FILLER_7_1192 ();
 sg13g2_decap_8 FILLER_7_1199 ();
 sg13g2_decap_8 FILLER_7_1206 ();
 sg13g2_decap_8 FILLER_7_1213 ();
 sg13g2_decap_8 FILLER_7_1220 ();
 sg13g2_decap_8 FILLER_7_1227 ();
 sg13g2_decap_8 FILLER_7_1234 ();
 sg13g2_decap_8 FILLER_7_1241 ();
 sg13g2_decap_8 FILLER_7_1248 ();
 sg13g2_decap_8 FILLER_7_1255 ();
 sg13g2_decap_8 FILLER_7_1262 ();
 sg13g2_decap_8 FILLER_7_1269 ();
 sg13g2_decap_8 FILLER_7_1276 ();
 sg13g2_decap_8 FILLER_7_1283 ();
 sg13g2_decap_8 FILLER_7_1290 ();
 sg13g2_decap_8 FILLER_7_1297 ();
 sg13g2_decap_8 FILLER_7_1304 ();
 sg13g2_decap_8 FILLER_7_1311 ();
 sg13g2_decap_8 FILLER_7_1318 ();
 sg13g2_decap_8 FILLER_7_1325 ();
 sg13g2_decap_8 FILLER_7_1332 ();
 sg13g2_decap_8 FILLER_7_1339 ();
 sg13g2_decap_8 FILLER_7_1346 ();
 sg13g2_decap_8 FILLER_7_1353 ();
 sg13g2_decap_8 FILLER_7_1360 ();
 sg13g2_decap_8 FILLER_7_1367 ();
 sg13g2_decap_8 FILLER_7_1374 ();
 sg13g2_decap_8 FILLER_7_1381 ();
 sg13g2_decap_8 FILLER_7_1388 ();
 sg13g2_decap_8 FILLER_7_1395 ();
 sg13g2_decap_8 FILLER_7_1402 ();
 sg13g2_decap_8 FILLER_7_1409 ();
 sg13g2_decap_8 FILLER_7_1416 ();
 sg13g2_decap_8 FILLER_7_1423 ();
 sg13g2_decap_8 FILLER_7_1430 ();
 sg13g2_decap_8 FILLER_7_1437 ();
 sg13g2_decap_8 FILLER_7_1444 ();
 sg13g2_decap_8 FILLER_7_1451 ();
 sg13g2_decap_8 FILLER_7_1458 ();
 sg13g2_decap_8 FILLER_7_1465 ();
 sg13g2_decap_8 FILLER_7_1472 ();
 sg13g2_decap_8 FILLER_7_1479 ();
 sg13g2_decap_8 FILLER_7_1486 ();
 sg13g2_decap_8 FILLER_7_1493 ();
 sg13g2_decap_8 FILLER_7_1500 ();
 sg13g2_decap_8 FILLER_7_1507 ();
 sg13g2_decap_8 FILLER_7_1514 ();
 sg13g2_decap_8 FILLER_7_1521 ();
 sg13g2_decap_8 FILLER_7_1528 ();
 sg13g2_decap_8 FILLER_7_1535 ();
 sg13g2_decap_8 FILLER_7_1542 ();
 sg13g2_decap_8 FILLER_7_1549 ();
 sg13g2_decap_8 FILLER_7_1556 ();
 sg13g2_decap_8 FILLER_7_1563 ();
 sg13g2_decap_8 FILLER_7_1570 ();
 sg13g2_decap_8 FILLER_7_1577 ();
 sg13g2_decap_8 FILLER_7_1584 ();
 sg13g2_decap_8 FILLER_7_1591 ();
 sg13g2_decap_8 FILLER_7_1598 ();
 sg13g2_decap_8 FILLER_7_1605 ();
 sg13g2_decap_8 FILLER_7_1612 ();
 sg13g2_decap_8 FILLER_7_1619 ();
 sg13g2_decap_8 FILLER_7_1626 ();
 sg13g2_decap_8 FILLER_7_1633 ();
 sg13g2_decap_8 FILLER_7_1640 ();
 sg13g2_decap_8 FILLER_7_1647 ();
 sg13g2_decap_8 FILLER_7_1654 ();
 sg13g2_decap_8 FILLER_7_1661 ();
 sg13g2_decap_8 FILLER_7_1668 ();
 sg13g2_decap_8 FILLER_7_1675 ();
 sg13g2_decap_8 FILLER_7_1682 ();
 sg13g2_decap_8 FILLER_7_1689 ();
 sg13g2_decap_8 FILLER_7_1696 ();
 sg13g2_decap_8 FILLER_7_1703 ();
 sg13g2_decap_8 FILLER_7_1710 ();
 sg13g2_decap_8 FILLER_7_1717 ();
 sg13g2_decap_8 FILLER_7_1724 ();
 sg13g2_decap_8 FILLER_7_1731 ();
 sg13g2_decap_8 FILLER_7_1738 ();
 sg13g2_decap_8 FILLER_7_1745 ();
 sg13g2_decap_8 FILLER_7_1752 ();
 sg13g2_decap_8 FILLER_7_1759 ();
 sg13g2_fill_2 FILLER_7_1766 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_4 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_151 ();
 sg13g2_fill_2 FILLER_8_162 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_fill_1 FILLER_8_175 ();
 sg13g2_fill_2 FILLER_8_246 ();
 sg13g2_fill_1 FILLER_8_248 ();
 sg13g2_fill_1 FILLER_8_283 ();
 sg13g2_fill_2 FILLER_8_312 ();
 sg13g2_fill_2 FILLER_8_478 ();
 sg13g2_fill_1 FILLER_8_480 ();
 sg13g2_decap_4 FILLER_8_551 ();
 sg13g2_fill_2 FILLER_8_555 ();
 sg13g2_fill_1 FILLER_8_562 ();
 sg13g2_fill_2 FILLER_8_568 ();
 sg13g2_decap_4 FILLER_8_586 ();
 sg13g2_fill_1 FILLER_8_590 ();
 sg13g2_decap_8 FILLER_8_625 ();
 sg13g2_decap_8 FILLER_8_632 ();
 sg13g2_decap_4 FILLER_8_639 ();
 sg13g2_decap_8 FILLER_8_668 ();
 sg13g2_fill_2 FILLER_8_675 ();
 sg13g2_fill_1 FILLER_8_677 ();
 sg13g2_fill_2 FILLER_8_693 ();
 sg13g2_fill_1 FILLER_8_695 ();
 sg13g2_fill_1 FILLER_8_711 ();
 sg13g2_fill_1 FILLER_8_716 ();
 sg13g2_fill_1 FILLER_8_726 ();
 sg13g2_decap_4 FILLER_8_745 ();
 sg13g2_fill_1 FILLER_8_749 ();
 sg13g2_fill_2 FILLER_8_760 ();
 sg13g2_decap_8 FILLER_8_809 ();
 sg13g2_decap_4 FILLER_8_821 ();
 sg13g2_fill_1 FILLER_8_825 ();
 sg13g2_fill_2 FILLER_8_836 ();
 sg13g2_fill_1 FILLER_8_838 ();
 sg13g2_decap_8 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_860 ();
 sg13g2_fill_2 FILLER_8_867 ();
 sg13g2_decap_4 FILLER_8_890 ();
 sg13g2_fill_2 FILLER_8_919 ();
 sg13g2_decap_4 FILLER_8_945 ();
 sg13g2_fill_2 FILLER_8_956 ();
 sg13g2_decap_8 FILLER_8_987 ();
 sg13g2_decap_4 FILLER_8_994 ();
 sg13g2_fill_2 FILLER_8_998 ();
 sg13g2_fill_1 FILLER_8_1005 ();
 sg13g2_decap_4 FILLER_8_1010 ();
 sg13g2_fill_1 FILLER_8_1014 ();
 sg13g2_decap_4 FILLER_8_1044 ();
 sg13g2_fill_2 FILLER_8_1048 ();
 sg13g2_decap_4 FILLER_8_1081 ();
 sg13g2_decap_4 FILLER_8_1099 ();
 sg13g2_fill_1 FILLER_8_1110 ();
 sg13g2_decap_8 FILLER_8_1134 ();
 sg13g2_decap_8 FILLER_8_1141 ();
 sg13g2_decap_8 FILLER_8_1148 ();
 sg13g2_decap_8 FILLER_8_1155 ();
 sg13g2_decap_8 FILLER_8_1162 ();
 sg13g2_decap_8 FILLER_8_1169 ();
 sg13g2_decap_8 FILLER_8_1176 ();
 sg13g2_decap_8 FILLER_8_1183 ();
 sg13g2_decap_8 FILLER_8_1190 ();
 sg13g2_decap_8 FILLER_8_1197 ();
 sg13g2_decap_8 FILLER_8_1204 ();
 sg13g2_decap_8 FILLER_8_1211 ();
 sg13g2_decap_8 FILLER_8_1218 ();
 sg13g2_decap_8 FILLER_8_1225 ();
 sg13g2_decap_8 FILLER_8_1232 ();
 sg13g2_decap_8 FILLER_8_1239 ();
 sg13g2_decap_8 FILLER_8_1246 ();
 sg13g2_decap_8 FILLER_8_1253 ();
 sg13g2_decap_8 FILLER_8_1260 ();
 sg13g2_decap_8 FILLER_8_1267 ();
 sg13g2_decap_8 FILLER_8_1274 ();
 sg13g2_decap_8 FILLER_8_1281 ();
 sg13g2_decap_8 FILLER_8_1288 ();
 sg13g2_decap_8 FILLER_8_1295 ();
 sg13g2_decap_8 FILLER_8_1302 ();
 sg13g2_decap_8 FILLER_8_1309 ();
 sg13g2_decap_8 FILLER_8_1316 ();
 sg13g2_decap_8 FILLER_8_1323 ();
 sg13g2_decap_8 FILLER_8_1330 ();
 sg13g2_decap_8 FILLER_8_1337 ();
 sg13g2_decap_8 FILLER_8_1344 ();
 sg13g2_decap_8 FILLER_8_1351 ();
 sg13g2_decap_8 FILLER_8_1358 ();
 sg13g2_decap_8 FILLER_8_1365 ();
 sg13g2_decap_8 FILLER_8_1372 ();
 sg13g2_decap_8 FILLER_8_1379 ();
 sg13g2_decap_8 FILLER_8_1386 ();
 sg13g2_decap_8 FILLER_8_1393 ();
 sg13g2_decap_8 FILLER_8_1400 ();
 sg13g2_decap_8 FILLER_8_1407 ();
 sg13g2_decap_8 FILLER_8_1414 ();
 sg13g2_decap_8 FILLER_8_1421 ();
 sg13g2_decap_8 FILLER_8_1428 ();
 sg13g2_decap_8 FILLER_8_1435 ();
 sg13g2_decap_8 FILLER_8_1442 ();
 sg13g2_decap_8 FILLER_8_1449 ();
 sg13g2_decap_8 FILLER_8_1456 ();
 sg13g2_decap_8 FILLER_8_1463 ();
 sg13g2_decap_8 FILLER_8_1470 ();
 sg13g2_decap_8 FILLER_8_1477 ();
 sg13g2_decap_8 FILLER_8_1484 ();
 sg13g2_decap_8 FILLER_8_1491 ();
 sg13g2_decap_8 FILLER_8_1498 ();
 sg13g2_decap_8 FILLER_8_1505 ();
 sg13g2_decap_8 FILLER_8_1512 ();
 sg13g2_decap_8 FILLER_8_1519 ();
 sg13g2_decap_8 FILLER_8_1526 ();
 sg13g2_decap_8 FILLER_8_1533 ();
 sg13g2_decap_8 FILLER_8_1540 ();
 sg13g2_decap_8 FILLER_8_1547 ();
 sg13g2_decap_8 FILLER_8_1554 ();
 sg13g2_decap_8 FILLER_8_1561 ();
 sg13g2_decap_8 FILLER_8_1568 ();
 sg13g2_decap_8 FILLER_8_1575 ();
 sg13g2_decap_8 FILLER_8_1582 ();
 sg13g2_decap_8 FILLER_8_1589 ();
 sg13g2_decap_8 FILLER_8_1596 ();
 sg13g2_decap_8 FILLER_8_1603 ();
 sg13g2_decap_8 FILLER_8_1610 ();
 sg13g2_decap_8 FILLER_8_1617 ();
 sg13g2_decap_8 FILLER_8_1624 ();
 sg13g2_decap_8 FILLER_8_1631 ();
 sg13g2_decap_8 FILLER_8_1638 ();
 sg13g2_decap_8 FILLER_8_1645 ();
 sg13g2_decap_8 FILLER_8_1652 ();
 sg13g2_decap_8 FILLER_8_1659 ();
 sg13g2_decap_8 FILLER_8_1666 ();
 sg13g2_decap_8 FILLER_8_1673 ();
 sg13g2_decap_8 FILLER_8_1680 ();
 sg13g2_decap_8 FILLER_8_1687 ();
 sg13g2_decap_8 FILLER_8_1694 ();
 sg13g2_decap_8 FILLER_8_1701 ();
 sg13g2_decap_8 FILLER_8_1708 ();
 sg13g2_decap_8 FILLER_8_1715 ();
 sg13g2_decap_8 FILLER_8_1722 ();
 sg13g2_decap_8 FILLER_8_1729 ();
 sg13g2_decap_8 FILLER_8_1736 ();
 sg13g2_decap_8 FILLER_8_1743 ();
 sg13g2_decap_8 FILLER_8_1750 ();
 sg13g2_decap_8 FILLER_8_1757 ();
 sg13g2_decap_4 FILLER_8_1764 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_66 ();
 sg13g2_decap_8 FILLER_9_73 ();
 sg13g2_fill_2 FILLER_9_80 ();
 sg13g2_fill_1 FILLER_9_82 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_fill_1 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_100 ();
 sg13g2_decap_8 FILLER_9_107 ();
 sg13g2_decap_8 FILLER_9_114 ();
 sg13g2_decap_8 FILLER_9_121 ();
 sg13g2_fill_2 FILLER_9_128 ();
 sg13g2_fill_1 FILLER_9_130 ();
 sg13g2_decap_4 FILLER_9_134 ();
 sg13g2_fill_1 FILLER_9_164 ();
 sg13g2_fill_2 FILLER_9_195 ();
 sg13g2_fill_2 FILLER_9_227 ();
 sg13g2_fill_1 FILLER_9_243 ();
 sg13g2_fill_1 FILLER_9_258 ();
 sg13g2_fill_1 FILLER_9_316 ();
 sg13g2_fill_2 FILLER_9_404 ();
 sg13g2_fill_2 FILLER_9_411 ();
 sg13g2_decap_4 FILLER_9_431 ();
 sg13g2_fill_1 FILLER_9_435 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_fill_2 FILLER_9_448 ();
 sg13g2_fill_2 FILLER_9_454 ();
 sg13g2_fill_1 FILLER_9_529 ();
 sg13g2_decap_8 FILLER_9_535 ();
 sg13g2_fill_1 FILLER_9_569 ();
 sg13g2_fill_1 FILLER_9_580 ();
 sg13g2_fill_2 FILLER_9_589 ();
 sg13g2_fill_1 FILLER_9_591 ();
 sg13g2_fill_2 FILLER_9_604 ();
 sg13g2_fill_1 FILLER_9_606 ();
 sg13g2_fill_2 FILLER_9_613 ();
 sg13g2_fill_2 FILLER_9_644 ();
 sg13g2_fill_1 FILLER_9_646 ();
 sg13g2_fill_1 FILLER_9_657 ();
 sg13g2_decap_4 FILLER_9_672 ();
 sg13g2_decap_4 FILLER_9_705 ();
 sg13g2_decap_8 FILLER_9_719 ();
 sg13g2_decap_4 FILLER_9_726 ();
 sg13g2_fill_1 FILLER_9_730 ();
 sg13g2_decap_4 FILLER_9_742 ();
 sg13g2_fill_2 FILLER_9_746 ();
 sg13g2_fill_1 FILLER_9_752 ();
 sg13g2_fill_1 FILLER_9_764 ();
 sg13g2_fill_2 FILLER_9_770 ();
 sg13g2_fill_1 FILLER_9_772 ();
 sg13g2_fill_2 FILLER_9_777 ();
 sg13g2_fill_2 FILLER_9_789 ();
 sg13g2_decap_4 FILLER_9_807 ();
 sg13g2_fill_1 FILLER_9_826 ();
 sg13g2_decap_4 FILLER_9_855 ();
 sg13g2_fill_2 FILLER_9_859 ();
 sg13g2_decap_8 FILLER_9_878 ();
 sg13g2_fill_1 FILLER_9_885 ();
 sg13g2_fill_2 FILLER_9_893 ();
 sg13g2_fill_1 FILLER_9_895 ();
 sg13g2_fill_2 FILLER_9_907 ();
 sg13g2_fill_1 FILLER_9_932 ();
 sg13g2_decap_8 FILLER_9_955 ();
 sg13g2_fill_2 FILLER_9_962 ();
 sg13g2_fill_1 FILLER_9_964 ();
 sg13g2_fill_1 FILLER_9_985 ();
 sg13g2_decap_8 FILLER_9_991 ();
 sg13g2_fill_2 FILLER_9_998 ();
 sg13g2_fill_1 FILLER_9_1000 ();
 sg13g2_fill_2 FILLER_9_1005 ();
 sg13g2_decap_4 FILLER_9_1023 ();
 sg13g2_fill_2 FILLER_9_1027 ();
 sg13g2_fill_2 FILLER_9_1042 ();
 sg13g2_decap_4 FILLER_9_1049 ();
 sg13g2_decap_4 FILLER_9_1062 ();
 sg13g2_fill_2 FILLER_9_1066 ();
 sg13g2_fill_2 FILLER_9_1073 ();
 sg13g2_fill_2 FILLER_9_1084 ();
 sg13g2_fill_1 FILLER_9_1086 ();
 sg13g2_decap_4 FILLER_9_1100 ();
 sg13g2_decap_8 FILLER_9_1134 ();
 sg13g2_decap_8 FILLER_9_1141 ();
 sg13g2_decap_8 FILLER_9_1148 ();
 sg13g2_decap_8 FILLER_9_1155 ();
 sg13g2_decap_8 FILLER_9_1162 ();
 sg13g2_decap_8 FILLER_9_1169 ();
 sg13g2_decap_8 FILLER_9_1176 ();
 sg13g2_decap_8 FILLER_9_1183 ();
 sg13g2_decap_8 FILLER_9_1190 ();
 sg13g2_decap_8 FILLER_9_1197 ();
 sg13g2_decap_8 FILLER_9_1204 ();
 sg13g2_decap_8 FILLER_9_1211 ();
 sg13g2_decap_8 FILLER_9_1218 ();
 sg13g2_decap_8 FILLER_9_1225 ();
 sg13g2_decap_8 FILLER_9_1232 ();
 sg13g2_decap_8 FILLER_9_1239 ();
 sg13g2_decap_8 FILLER_9_1246 ();
 sg13g2_decap_8 FILLER_9_1253 ();
 sg13g2_decap_8 FILLER_9_1260 ();
 sg13g2_decap_8 FILLER_9_1267 ();
 sg13g2_decap_8 FILLER_9_1274 ();
 sg13g2_decap_8 FILLER_9_1281 ();
 sg13g2_decap_8 FILLER_9_1288 ();
 sg13g2_decap_8 FILLER_9_1295 ();
 sg13g2_decap_8 FILLER_9_1302 ();
 sg13g2_decap_8 FILLER_9_1309 ();
 sg13g2_decap_8 FILLER_9_1316 ();
 sg13g2_decap_8 FILLER_9_1323 ();
 sg13g2_decap_8 FILLER_9_1330 ();
 sg13g2_decap_8 FILLER_9_1337 ();
 sg13g2_decap_8 FILLER_9_1344 ();
 sg13g2_decap_8 FILLER_9_1351 ();
 sg13g2_decap_8 FILLER_9_1358 ();
 sg13g2_decap_8 FILLER_9_1365 ();
 sg13g2_decap_8 FILLER_9_1372 ();
 sg13g2_decap_8 FILLER_9_1379 ();
 sg13g2_decap_8 FILLER_9_1386 ();
 sg13g2_decap_8 FILLER_9_1393 ();
 sg13g2_decap_8 FILLER_9_1400 ();
 sg13g2_decap_8 FILLER_9_1407 ();
 sg13g2_decap_8 FILLER_9_1414 ();
 sg13g2_decap_8 FILLER_9_1421 ();
 sg13g2_decap_8 FILLER_9_1428 ();
 sg13g2_decap_8 FILLER_9_1435 ();
 sg13g2_decap_8 FILLER_9_1442 ();
 sg13g2_decap_8 FILLER_9_1449 ();
 sg13g2_decap_8 FILLER_9_1456 ();
 sg13g2_decap_8 FILLER_9_1463 ();
 sg13g2_decap_8 FILLER_9_1470 ();
 sg13g2_decap_8 FILLER_9_1477 ();
 sg13g2_decap_8 FILLER_9_1484 ();
 sg13g2_decap_8 FILLER_9_1491 ();
 sg13g2_decap_8 FILLER_9_1498 ();
 sg13g2_decap_8 FILLER_9_1505 ();
 sg13g2_decap_8 FILLER_9_1512 ();
 sg13g2_decap_8 FILLER_9_1519 ();
 sg13g2_decap_8 FILLER_9_1526 ();
 sg13g2_decap_8 FILLER_9_1533 ();
 sg13g2_decap_8 FILLER_9_1540 ();
 sg13g2_decap_8 FILLER_9_1547 ();
 sg13g2_decap_8 FILLER_9_1554 ();
 sg13g2_decap_8 FILLER_9_1561 ();
 sg13g2_decap_8 FILLER_9_1568 ();
 sg13g2_decap_8 FILLER_9_1575 ();
 sg13g2_decap_8 FILLER_9_1582 ();
 sg13g2_decap_8 FILLER_9_1589 ();
 sg13g2_decap_8 FILLER_9_1596 ();
 sg13g2_decap_8 FILLER_9_1603 ();
 sg13g2_decap_8 FILLER_9_1610 ();
 sg13g2_decap_8 FILLER_9_1617 ();
 sg13g2_decap_8 FILLER_9_1624 ();
 sg13g2_decap_8 FILLER_9_1631 ();
 sg13g2_decap_8 FILLER_9_1638 ();
 sg13g2_decap_8 FILLER_9_1645 ();
 sg13g2_decap_8 FILLER_9_1652 ();
 sg13g2_decap_8 FILLER_9_1659 ();
 sg13g2_decap_8 FILLER_9_1666 ();
 sg13g2_decap_8 FILLER_9_1673 ();
 sg13g2_decap_8 FILLER_9_1680 ();
 sg13g2_decap_8 FILLER_9_1687 ();
 sg13g2_decap_8 FILLER_9_1694 ();
 sg13g2_decap_8 FILLER_9_1701 ();
 sg13g2_decap_8 FILLER_9_1708 ();
 sg13g2_decap_8 FILLER_9_1715 ();
 sg13g2_decap_8 FILLER_9_1722 ();
 sg13g2_decap_8 FILLER_9_1729 ();
 sg13g2_decap_8 FILLER_9_1736 ();
 sg13g2_decap_8 FILLER_9_1743 ();
 sg13g2_decap_8 FILLER_9_1750 ();
 sg13g2_decap_8 FILLER_9_1757 ();
 sg13g2_decap_4 FILLER_9_1764 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_49 ();
 sg13g2_fill_1 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_135 ();
 sg13g2_fill_2 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_180 ();
 sg13g2_fill_1 FILLER_10_182 ();
 sg13g2_fill_1 FILLER_10_188 ();
 sg13g2_fill_2 FILLER_10_224 ();
 sg13g2_fill_1 FILLER_10_226 ();
 sg13g2_fill_2 FILLER_10_299 ();
 sg13g2_fill_1 FILLER_10_301 ();
 sg13g2_fill_2 FILLER_10_307 ();
 sg13g2_fill_2 FILLER_10_336 ();
 sg13g2_fill_1 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_10_496 ();
 sg13g2_decap_8 FILLER_10_537 ();
 sg13g2_decap_4 FILLER_10_544 ();
 sg13g2_fill_1 FILLER_10_548 ();
 sg13g2_fill_2 FILLER_10_559 ();
 sg13g2_fill_2 FILLER_10_581 ();
 sg13g2_fill_2 FILLER_10_593 ();
 sg13g2_decap_4 FILLER_10_600 ();
 sg13g2_fill_1 FILLER_10_604 ();
 sg13g2_fill_1 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_619 ();
 sg13g2_fill_2 FILLER_10_626 ();
 sg13g2_fill_1 FILLER_10_628 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_fill_2 FILLER_10_648 ();
 sg13g2_fill_2 FILLER_10_662 ();
 sg13g2_fill_1 FILLER_10_685 ();
 sg13g2_fill_1 FILLER_10_710 ();
 sg13g2_fill_1 FILLER_10_723 ();
 sg13g2_fill_1 FILLER_10_773 ();
 sg13g2_fill_2 FILLER_10_785 ();
 sg13g2_fill_1 FILLER_10_787 ();
 sg13g2_fill_2 FILLER_10_804 ();
 sg13g2_fill_2 FILLER_10_821 ();
 sg13g2_fill_1 FILLER_10_823 ();
 sg13g2_fill_1 FILLER_10_841 ();
 sg13g2_decap_8 FILLER_10_852 ();
 sg13g2_decap_8 FILLER_10_859 ();
 sg13g2_decap_8 FILLER_10_866 ();
 sg13g2_decap_8 FILLER_10_873 ();
 sg13g2_decap_4 FILLER_10_880 ();
 sg13g2_fill_2 FILLER_10_884 ();
 sg13g2_decap_8 FILLER_10_914 ();
 sg13g2_fill_1 FILLER_10_921 ();
 sg13g2_fill_2 FILLER_10_926 ();
 sg13g2_decap_8 FILLER_10_933 ();
 sg13g2_decap_4 FILLER_10_949 ();
 sg13g2_fill_2 FILLER_10_953 ();
 sg13g2_fill_2 FILLER_10_965 ();
 sg13g2_fill_1 FILLER_10_967 ();
 sg13g2_fill_2 FILLER_10_978 ();
 sg13g2_fill_1 FILLER_10_980 ();
 sg13g2_decap_8 FILLER_10_1015 ();
 sg13g2_fill_1 FILLER_10_1022 ();
 sg13g2_decap_8 FILLER_10_1034 ();
 sg13g2_decap_4 FILLER_10_1041 ();
 sg13g2_fill_2 FILLER_10_1080 ();
 sg13g2_fill_2 FILLER_10_1087 ();
 sg13g2_fill_1 FILLER_10_1089 ();
 sg13g2_decap_4 FILLER_10_1095 ();
 sg13g2_fill_2 FILLER_10_1112 ();
 sg13g2_fill_1 FILLER_10_1114 ();
 sg13g2_decap_8 FILLER_10_1131 ();
 sg13g2_decap_8 FILLER_10_1138 ();
 sg13g2_decap_8 FILLER_10_1145 ();
 sg13g2_decap_8 FILLER_10_1152 ();
 sg13g2_decap_8 FILLER_10_1159 ();
 sg13g2_decap_8 FILLER_10_1166 ();
 sg13g2_decap_8 FILLER_10_1173 ();
 sg13g2_decap_8 FILLER_10_1180 ();
 sg13g2_decap_8 FILLER_10_1187 ();
 sg13g2_decap_8 FILLER_10_1194 ();
 sg13g2_decap_8 FILLER_10_1201 ();
 sg13g2_decap_8 FILLER_10_1208 ();
 sg13g2_decap_8 FILLER_10_1215 ();
 sg13g2_decap_8 FILLER_10_1222 ();
 sg13g2_decap_8 FILLER_10_1229 ();
 sg13g2_decap_8 FILLER_10_1236 ();
 sg13g2_decap_8 FILLER_10_1243 ();
 sg13g2_decap_8 FILLER_10_1250 ();
 sg13g2_decap_8 FILLER_10_1257 ();
 sg13g2_decap_8 FILLER_10_1264 ();
 sg13g2_decap_8 FILLER_10_1271 ();
 sg13g2_decap_8 FILLER_10_1278 ();
 sg13g2_decap_8 FILLER_10_1285 ();
 sg13g2_decap_8 FILLER_10_1292 ();
 sg13g2_decap_8 FILLER_10_1299 ();
 sg13g2_decap_8 FILLER_10_1306 ();
 sg13g2_decap_8 FILLER_10_1313 ();
 sg13g2_decap_8 FILLER_10_1320 ();
 sg13g2_decap_8 FILLER_10_1327 ();
 sg13g2_decap_8 FILLER_10_1334 ();
 sg13g2_decap_8 FILLER_10_1341 ();
 sg13g2_decap_8 FILLER_10_1348 ();
 sg13g2_decap_8 FILLER_10_1355 ();
 sg13g2_decap_8 FILLER_10_1362 ();
 sg13g2_decap_8 FILLER_10_1369 ();
 sg13g2_decap_8 FILLER_10_1376 ();
 sg13g2_decap_8 FILLER_10_1383 ();
 sg13g2_decap_8 FILLER_10_1390 ();
 sg13g2_decap_8 FILLER_10_1397 ();
 sg13g2_decap_8 FILLER_10_1404 ();
 sg13g2_decap_8 FILLER_10_1411 ();
 sg13g2_decap_8 FILLER_10_1418 ();
 sg13g2_decap_8 FILLER_10_1425 ();
 sg13g2_decap_8 FILLER_10_1432 ();
 sg13g2_decap_8 FILLER_10_1439 ();
 sg13g2_decap_8 FILLER_10_1446 ();
 sg13g2_decap_8 FILLER_10_1453 ();
 sg13g2_decap_8 FILLER_10_1460 ();
 sg13g2_decap_8 FILLER_10_1467 ();
 sg13g2_decap_8 FILLER_10_1474 ();
 sg13g2_decap_8 FILLER_10_1481 ();
 sg13g2_decap_8 FILLER_10_1488 ();
 sg13g2_decap_8 FILLER_10_1495 ();
 sg13g2_decap_8 FILLER_10_1502 ();
 sg13g2_decap_8 FILLER_10_1509 ();
 sg13g2_decap_8 FILLER_10_1516 ();
 sg13g2_decap_8 FILLER_10_1523 ();
 sg13g2_decap_8 FILLER_10_1530 ();
 sg13g2_decap_8 FILLER_10_1537 ();
 sg13g2_decap_8 FILLER_10_1544 ();
 sg13g2_decap_8 FILLER_10_1551 ();
 sg13g2_decap_8 FILLER_10_1558 ();
 sg13g2_decap_8 FILLER_10_1565 ();
 sg13g2_decap_8 FILLER_10_1572 ();
 sg13g2_decap_8 FILLER_10_1579 ();
 sg13g2_decap_8 FILLER_10_1586 ();
 sg13g2_decap_8 FILLER_10_1593 ();
 sg13g2_decap_8 FILLER_10_1600 ();
 sg13g2_decap_8 FILLER_10_1607 ();
 sg13g2_decap_8 FILLER_10_1614 ();
 sg13g2_decap_8 FILLER_10_1621 ();
 sg13g2_decap_8 FILLER_10_1628 ();
 sg13g2_decap_8 FILLER_10_1635 ();
 sg13g2_decap_8 FILLER_10_1642 ();
 sg13g2_decap_8 FILLER_10_1649 ();
 sg13g2_decap_8 FILLER_10_1656 ();
 sg13g2_decap_8 FILLER_10_1663 ();
 sg13g2_decap_8 FILLER_10_1670 ();
 sg13g2_decap_8 FILLER_10_1677 ();
 sg13g2_decap_8 FILLER_10_1684 ();
 sg13g2_decap_8 FILLER_10_1691 ();
 sg13g2_decap_8 FILLER_10_1698 ();
 sg13g2_decap_8 FILLER_10_1705 ();
 sg13g2_decap_8 FILLER_10_1712 ();
 sg13g2_decap_8 FILLER_10_1719 ();
 sg13g2_decap_8 FILLER_10_1726 ();
 sg13g2_decap_8 FILLER_10_1733 ();
 sg13g2_decap_8 FILLER_10_1740 ();
 sg13g2_decap_8 FILLER_10_1747 ();
 sg13g2_decap_8 FILLER_10_1754 ();
 sg13g2_decap_8 FILLER_10_1761 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_4 FILLER_11_42 ();
 sg13g2_fill_2 FILLER_11_46 ();
 sg13g2_fill_1 FILLER_11_66 ();
 sg13g2_fill_1 FILLER_11_85 ();
 sg13g2_fill_2 FILLER_11_118 ();
 sg13g2_fill_1 FILLER_11_186 ();
 sg13g2_fill_2 FILLER_11_237 ();
 sg13g2_fill_1 FILLER_11_239 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_fill_2 FILLER_11_291 ();
 sg13g2_fill_1 FILLER_11_324 ();
 sg13g2_fill_1 FILLER_11_407 ();
 sg13g2_fill_2 FILLER_11_413 ();
 sg13g2_fill_2 FILLER_11_514 ();
 sg13g2_fill_2 FILLER_11_524 ();
 sg13g2_decap_8 FILLER_11_557 ();
 sg13g2_decap_4 FILLER_11_564 ();
 sg13g2_decap_4 FILLER_11_585 ();
 sg13g2_decap_8 FILLER_11_596 ();
 sg13g2_fill_2 FILLER_11_618 ();
 sg13g2_fill_1 FILLER_11_620 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_fill_2 FILLER_11_644 ();
 sg13g2_decap_4 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_666 ();
 sg13g2_decap_4 FILLER_11_673 ();
 sg13g2_decap_4 FILLER_11_696 ();
 sg13g2_fill_1 FILLER_11_714 ();
 sg13g2_decap_4 FILLER_11_725 ();
 sg13g2_fill_1 FILLER_11_745 ();
 sg13g2_fill_2 FILLER_11_759 ();
 sg13g2_fill_1 FILLER_11_761 ();
 sg13g2_decap_4 FILLER_11_767 ();
 sg13g2_fill_1 FILLER_11_771 ();
 sg13g2_fill_2 FILLER_11_776 ();
 sg13g2_fill_1 FILLER_11_778 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_fill_2 FILLER_11_828 ();
 sg13g2_decap_8 FILLER_11_856 ();
 sg13g2_decap_8 FILLER_11_863 ();
 sg13g2_fill_2 FILLER_11_875 ();
 sg13g2_fill_1 FILLER_11_877 ();
 sg13g2_decap_4 FILLER_11_883 ();
 sg13g2_fill_1 FILLER_11_887 ();
 sg13g2_decap_8 FILLER_11_907 ();
 sg13g2_fill_1 FILLER_11_914 ();
 sg13g2_fill_2 FILLER_11_926 ();
 sg13g2_fill_1 FILLER_11_928 ();
 sg13g2_decap_4 FILLER_11_933 ();
 sg13g2_fill_1 FILLER_11_942 ();
 sg13g2_decap_8 FILLER_11_958 ();
 sg13g2_fill_1 FILLER_11_965 ();
 sg13g2_decap_8 FILLER_11_992 ();
 sg13g2_fill_1 FILLER_11_999 ();
 sg13g2_fill_1 FILLER_11_1016 ();
 sg13g2_decap_8 FILLER_11_1045 ();
 sg13g2_fill_2 FILLER_11_1052 ();
 sg13g2_fill_1 FILLER_11_1054 ();
 sg13g2_fill_1 FILLER_11_1065 ();
 sg13g2_decap_4 FILLER_11_1074 ();
 sg13g2_decap_8 FILLER_11_1098 ();
 sg13g2_decap_8 FILLER_11_1124 ();
 sg13g2_decap_8 FILLER_11_1131 ();
 sg13g2_decap_8 FILLER_11_1138 ();
 sg13g2_decap_8 FILLER_11_1145 ();
 sg13g2_decap_8 FILLER_11_1152 ();
 sg13g2_decap_8 FILLER_11_1159 ();
 sg13g2_decap_8 FILLER_11_1166 ();
 sg13g2_decap_8 FILLER_11_1173 ();
 sg13g2_decap_8 FILLER_11_1180 ();
 sg13g2_decap_8 FILLER_11_1187 ();
 sg13g2_decap_8 FILLER_11_1194 ();
 sg13g2_decap_8 FILLER_11_1201 ();
 sg13g2_decap_8 FILLER_11_1208 ();
 sg13g2_decap_8 FILLER_11_1215 ();
 sg13g2_decap_8 FILLER_11_1222 ();
 sg13g2_decap_8 FILLER_11_1229 ();
 sg13g2_decap_8 FILLER_11_1236 ();
 sg13g2_decap_8 FILLER_11_1243 ();
 sg13g2_decap_8 FILLER_11_1250 ();
 sg13g2_decap_8 FILLER_11_1257 ();
 sg13g2_decap_8 FILLER_11_1264 ();
 sg13g2_decap_8 FILLER_11_1271 ();
 sg13g2_decap_8 FILLER_11_1278 ();
 sg13g2_decap_8 FILLER_11_1285 ();
 sg13g2_decap_8 FILLER_11_1292 ();
 sg13g2_decap_8 FILLER_11_1299 ();
 sg13g2_decap_8 FILLER_11_1306 ();
 sg13g2_decap_8 FILLER_11_1313 ();
 sg13g2_decap_8 FILLER_11_1320 ();
 sg13g2_decap_8 FILLER_11_1327 ();
 sg13g2_decap_8 FILLER_11_1334 ();
 sg13g2_decap_8 FILLER_11_1341 ();
 sg13g2_decap_8 FILLER_11_1348 ();
 sg13g2_decap_8 FILLER_11_1355 ();
 sg13g2_decap_8 FILLER_11_1362 ();
 sg13g2_decap_8 FILLER_11_1369 ();
 sg13g2_decap_8 FILLER_11_1376 ();
 sg13g2_decap_8 FILLER_11_1383 ();
 sg13g2_decap_8 FILLER_11_1390 ();
 sg13g2_decap_8 FILLER_11_1397 ();
 sg13g2_decap_8 FILLER_11_1404 ();
 sg13g2_decap_8 FILLER_11_1411 ();
 sg13g2_decap_8 FILLER_11_1418 ();
 sg13g2_decap_8 FILLER_11_1425 ();
 sg13g2_decap_8 FILLER_11_1432 ();
 sg13g2_decap_8 FILLER_11_1439 ();
 sg13g2_decap_8 FILLER_11_1446 ();
 sg13g2_decap_8 FILLER_11_1453 ();
 sg13g2_decap_8 FILLER_11_1460 ();
 sg13g2_decap_8 FILLER_11_1467 ();
 sg13g2_decap_8 FILLER_11_1474 ();
 sg13g2_decap_8 FILLER_11_1481 ();
 sg13g2_decap_8 FILLER_11_1488 ();
 sg13g2_decap_8 FILLER_11_1495 ();
 sg13g2_decap_8 FILLER_11_1502 ();
 sg13g2_decap_8 FILLER_11_1509 ();
 sg13g2_decap_8 FILLER_11_1516 ();
 sg13g2_decap_8 FILLER_11_1523 ();
 sg13g2_decap_8 FILLER_11_1530 ();
 sg13g2_decap_8 FILLER_11_1537 ();
 sg13g2_decap_8 FILLER_11_1544 ();
 sg13g2_decap_8 FILLER_11_1551 ();
 sg13g2_decap_8 FILLER_11_1558 ();
 sg13g2_decap_8 FILLER_11_1565 ();
 sg13g2_decap_8 FILLER_11_1572 ();
 sg13g2_decap_8 FILLER_11_1579 ();
 sg13g2_decap_8 FILLER_11_1586 ();
 sg13g2_decap_8 FILLER_11_1593 ();
 sg13g2_decap_8 FILLER_11_1600 ();
 sg13g2_decap_8 FILLER_11_1607 ();
 sg13g2_decap_8 FILLER_11_1614 ();
 sg13g2_decap_8 FILLER_11_1621 ();
 sg13g2_decap_8 FILLER_11_1628 ();
 sg13g2_decap_8 FILLER_11_1635 ();
 sg13g2_decap_8 FILLER_11_1642 ();
 sg13g2_decap_8 FILLER_11_1649 ();
 sg13g2_decap_8 FILLER_11_1656 ();
 sg13g2_decap_8 FILLER_11_1663 ();
 sg13g2_decap_8 FILLER_11_1670 ();
 sg13g2_decap_8 FILLER_11_1677 ();
 sg13g2_decap_8 FILLER_11_1684 ();
 sg13g2_decap_8 FILLER_11_1691 ();
 sg13g2_decap_8 FILLER_11_1698 ();
 sg13g2_decap_8 FILLER_11_1705 ();
 sg13g2_decap_8 FILLER_11_1712 ();
 sg13g2_decap_8 FILLER_11_1719 ();
 sg13g2_decap_8 FILLER_11_1726 ();
 sg13g2_decap_8 FILLER_11_1733 ();
 sg13g2_decap_8 FILLER_11_1740 ();
 sg13g2_decap_8 FILLER_11_1747 ();
 sg13g2_decap_8 FILLER_11_1754 ();
 sg13g2_decap_8 FILLER_11_1761 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_4 FILLER_12_35 ();
 sg13g2_fill_1 FILLER_12_39 ();
 sg13g2_fill_1 FILLER_12_53 ();
 sg13g2_fill_1 FILLER_12_85 ();
 sg13g2_fill_1 FILLER_12_94 ();
 sg13g2_fill_2 FILLER_12_134 ();
 sg13g2_fill_1 FILLER_12_197 ();
 sg13g2_fill_2 FILLER_12_220 ();
 sg13g2_fill_2 FILLER_12_255 ();
 sg13g2_fill_1 FILLER_12_257 ();
 sg13g2_fill_2 FILLER_12_267 ();
 sg13g2_fill_1 FILLER_12_269 ();
 sg13g2_decap_4 FILLER_12_322 ();
 sg13g2_fill_1 FILLER_12_347 ();
 sg13g2_fill_2 FILLER_12_408 ();
 sg13g2_fill_2 FILLER_12_444 ();
 sg13g2_fill_1 FILLER_12_446 ();
 sg13g2_fill_1 FILLER_12_453 ();
 sg13g2_fill_2 FILLER_12_477 ();
 sg13g2_fill_1 FILLER_12_482 ();
 sg13g2_fill_2 FILLER_12_503 ();
 sg13g2_fill_2 FILLER_12_510 ();
 sg13g2_fill_1 FILLER_12_512 ();
 sg13g2_fill_2 FILLER_12_558 ();
 sg13g2_fill_2 FILLER_12_568 ();
 sg13g2_fill_1 FILLER_12_570 ();
 sg13g2_fill_2 FILLER_12_592 ();
 sg13g2_fill_1 FILLER_12_594 ();
 sg13g2_fill_2 FILLER_12_611 ();
 sg13g2_fill_1 FILLER_12_613 ();
 sg13g2_fill_2 FILLER_12_632 ();
 sg13g2_fill_2 FILLER_12_664 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_fill_2 FILLER_12_686 ();
 sg13g2_fill_2 FILLER_12_692 ();
 sg13g2_fill_1 FILLER_12_694 ();
 sg13g2_fill_2 FILLER_12_700 ();
 sg13g2_fill_1 FILLER_12_702 ();
 sg13g2_fill_2 FILLER_12_708 ();
 sg13g2_fill_1 FILLER_12_710 ();
 sg13g2_fill_2 FILLER_12_743 ();
 sg13g2_fill_1 FILLER_12_769 ();
 sg13g2_fill_1 FILLER_12_785 ();
 sg13g2_decap_8 FILLER_12_796 ();
 sg13g2_fill_1 FILLER_12_803 ();
 sg13g2_fill_1 FILLER_12_809 ();
 sg13g2_fill_1 FILLER_12_815 ();
 sg13g2_fill_2 FILLER_12_824 ();
 sg13g2_fill_2 FILLER_12_841 ();
 sg13g2_decap_8 FILLER_12_885 ();
 sg13g2_fill_2 FILLER_12_892 ();
 sg13g2_fill_1 FILLER_12_899 ();
 sg13g2_decap_4 FILLER_12_909 ();
 sg13g2_fill_2 FILLER_12_918 ();
 sg13g2_fill_1 FILLER_12_920 ();
 sg13g2_decap_4 FILLER_12_942 ();
 sg13g2_fill_2 FILLER_12_957 ();
 sg13g2_fill_1 FILLER_12_959 ();
 sg13g2_decap_4 FILLER_12_964 ();
 sg13g2_fill_1 FILLER_12_968 ();
 sg13g2_fill_2 FILLER_12_973 ();
 sg13g2_fill_1 FILLER_12_990 ();
 sg13g2_fill_2 FILLER_12_996 ();
 sg13g2_fill_1 FILLER_12_998 ();
 sg13g2_fill_2 FILLER_12_1008 ();
 sg13g2_decap_4 FILLER_12_1014 ();
 sg13g2_decap_4 FILLER_12_1023 ();
 sg13g2_fill_1 FILLER_12_1027 ();
 sg13g2_decap_4 FILLER_12_1034 ();
 sg13g2_fill_1 FILLER_12_1038 ();
 sg13g2_decap_4 FILLER_12_1057 ();
 sg13g2_fill_1 FILLER_12_1061 ();
 sg13g2_fill_2 FILLER_12_1084 ();
 sg13g2_fill_1 FILLER_12_1086 ();
 sg13g2_fill_1 FILLER_12_1106 ();
 sg13g2_decap_8 FILLER_12_1121 ();
 sg13g2_decap_8 FILLER_12_1128 ();
 sg13g2_decap_8 FILLER_12_1135 ();
 sg13g2_decap_8 FILLER_12_1142 ();
 sg13g2_decap_8 FILLER_12_1149 ();
 sg13g2_decap_8 FILLER_12_1156 ();
 sg13g2_decap_8 FILLER_12_1163 ();
 sg13g2_decap_8 FILLER_12_1170 ();
 sg13g2_decap_8 FILLER_12_1177 ();
 sg13g2_decap_8 FILLER_12_1184 ();
 sg13g2_decap_8 FILLER_12_1191 ();
 sg13g2_decap_8 FILLER_12_1198 ();
 sg13g2_decap_8 FILLER_12_1205 ();
 sg13g2_decap_8 FILLER_12_1212 ();
 sg13g2_decap_8 FILLER_12_1219 ();
 sg13g2_decap_8 FILLER_12_1226 ();
 sg13g2_decap_8 FILLER_12_1233 ();
 sg13g2_decap_8 FILLER_12_1240 ();
 sg13g2_decap_8 FILLER_12_1247 ();
 sg13g2_decap_8 FILLER_12_1254 ();
 sg13g2_decap_8 FILLER_12_1261 ();
 sg13g2_decap_8 FILLER_12_1268 ();
 sg13g2_decap_8 FILLER_12_1275 ();
 sg13g2_decap_8 FILLER_12_1282 ();
 sg13g2_decap_8 FILLER_12_1289 ();
 sg13g2_decap_8 FILLER_12_1296 ();
 sg13g2_decap_8 FILLER_12_1303 ();
 sg13g2_decap_8 FILLER_12_1310 ();
 sg13g2_decap_8 FILLER_12_1317 ();
 sg13g2_decap_8 FILLER_12_1324 ();
 sg13g2_decap_8 FILLER_12_1331 ();
 sg13g2_decap_8 FILLER_12_1338 ();
 sg13g2_decap_8 FILLER_12_1345 ();
 sg13g2_decap_8 FILLER_12_1352 ();
 sg13g2_decap_8 FILLER_12_1359 ();
 sg13g2_decap_8 FILLER_12_1366 ();
 sg13g2_decap_8 FILLER_12_1373 ();
 sg13g2_decap_8 FILLER_12_1380 ();
 sg13g2_decap_8 FILLER_12_1387 ();
 sg13g2_decap_8 FILLER_12_1394 ();
 sg13g2_decap_8 FILLER_12_1401 ();
 sg13g2_decap_8 FILLER_12_1408 ();
 sg13g2_decap_8 FILLER_12_1415 ();
 sg13g2_decap_8 FILLER_12_1422 ();
 sg13g2_decap_8 FILLER_12_1429 ();
 sg13g2_decap_8 FILLER_12_1436 ();
 sg13g2_decap_8 FILLER_12_1443 ();
 sg13g2_decap_8 FILLER_12_1450 ();
 sg13g2_decap_8 FILLER_12_1457 ();
 sg13g2_decap_8 FILLER_12_1464 ();
 sg13g2_decap_8 FILLER_12_1471 ();
 sg13g2_decap_8 FILLER_12_1478 ();
 sg13g2_decap_8 FILLER_12_1485 ();
 sg13g2_decap_8 FILLER_12_1492 ();
 sg13g2_decap_8 FILLER_12_1499 ();
 sg13g2_decap_8 FILLER_12_1506 ();
 sg13g2_decap_8 FILLER_12_1513 ();
 sg13g2_decap_8 FILLER_12_1520 ();
 sg13g2_decap_8 FILLER_12_1527 ();
 sg13g2_decap_8 FILLER_12_1534 ();
 sg13g2_decap_8 FILLER_12_1541 ();
 sg13g2_decap_8 FILLER_12_1548 ();
 sg13g2_decap_8 FILLER_12_1555 ();
 sg13g2_decap_8 FILLER_12_1562 ();
 sg13g2_decap_8 FILLER_12_1569 ();
 sg13g2_decap_8 FILLER_12_1576 ();
 sg13g2_decap_8 FILLER_12_1583 ();
 sg13g2_decap_8 FILLER_12_1590 ();
 sg13g2_decap_8 FILLER_12_1597 ();
 sg13g2_decap_8 FILLER_12_1604 ();
 sg13g2_decap_8 FILLER_12_1611 ();
 sg13g2_decap_8 FILLER_12_1618 ();
 sg13g2_decap_8 FILLER_12_1625 ();
 sg13g2_decap_8 FILLER_12_1632 ();
 sg13g2_decap_8 FILLER_12_1639 ();
 sg13g2_decap_8 FILLER_12_1646 ();
 sg13g2_decap_8 FILLER_12_1653 ();
 sg13g2_decap_8 FILLER_12_1660 ();
 sg13g2_decap_8 FILLER_12_1667 ();
 sg13g2_decap_8 FILLER_12_1674 ();
 sg13g2_decap_8 FILLER_12_1681 ();
 sg13g2_decap_8 FILLER_12_1688 ();
 sg13g2_decap_8 FILLER_12_1695 ();
 sg13g2_decap_8 FILLER_12_1702 ();
 sg13g2_decap_8 FILLER_12_1709 ();
 sg13g2_decap_8 FILLER_12_1716 ();
 sg13g2_decap_8 FILLER_12_1723 ();
 sg13g2_decap_8 FILLER_12_1730 ();
 sg13g2_decap_8 FILLER_12_1737 ();
 sg13g2_decap_8 FILLER_12_1744 ();
 sg13g2_decap_8 FILLER_12_1751 ();
 sg13g2_decap_8 FILLER_12_1758 ();
 sg13g2_fill_2 FILLER_12_1765 ();
 sg13g2_fill_1 FILLER_12_1767 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_32 ();
 sg13g2_fill_2 FILLER_13_60 ();
 sg13g2_fill_1 FILLER_13_62 ();
 sg13g2_fill_2 FILLER_13_92 ();
 sg13g2_fill_1 FILLER_13_106 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_fill_1 FILLER_13_131 ();
 sg13g2_decap_4 FILLER_13_158 ();
 sg13g2_fill_1 FILLER_13_162 ();
 sg13g2_fill_2 FILLER_13_170 ();
 sg13g2_fill_1 FILLER_13_172 ();
 sg13g2_decap_4 FILLER_13_180 ();
 sg13g2_decap_8 FILLER_13_279 ();
 sg13g2_fill_2 FILLER_13_286 ();
 sg13g2_fill_2 FILLER_13_300 ();
 sg13g2_fill_1 FILLER_13_302 ();
 sg13g2_fill_1 FILLER_13_347 ();
 sg13g2_fill_2 FILLER_13_356 ();
 sg13g2_fill_1 FILLER_13_382 ();
 sg13g2_fill_2 FILLER_13_432 ();
 sg13g2_fill_1 FILLER_13_434 ();
 sg13g2_decap_4 FILLER_13_463 ();
 sg13g2_fill_1 FILLER_13_480 ();
 sg13g2_decap_8 FILLER_13_486 ();
 sg13g2_decap_4 FILLER_13_493 ();
 sg13g2_decap_4 FILLER_13_502 ();
 sg13g2_fill_1 FILLER_13_506 ();
 sg13g2_fill_2 FILLER_13_512 ();
 sg13g2_fill_1 FILLER_13_514 ();
 sg13g2_fill_2 FILLER_13_526 ();
 sg13g2_decap_8 FILLER_13_555 ();
 sg13g2_fill_2 FILLER_13_562 ();
 sg13g2_decap_8 FILLER_13_576 ();
 sg13g2_decap_8 FILLER_13_583 ();
 sg13g2_decap_4 FILLER_13_590 ();
 sg13g2_fill_2 FILLER_13_620 ();
 sg13g2_fill_2 FILLER_13_638 ();
 sg13g2_decap_4 FILLER_13_655 ();
 sg13g2_fill_1 FILLER_13_659 ();
 sg13g2_decap_8 FILLER_13_668 ();
 sg13g2_fill_2 FILLER_13_675 ();
 sg13g2_decap_4 FILLER_13_685 ();
 sg13g2_fill_2 FILLER_13_689 ();
 sg13g2_decap_4 FILLER_13_765 ();
 sg13g2_decap_4 FILLER_13_782 ();
 sg13g2_fill_2 FILLER_13_786 ();
 sg13g2_fill_1 FILLER_13_793 ();
 sg13g2_decap_4 FILLER_13_801 ();
 sg13g2_fill_2 FILLER_13_805 ();
 sg13g2_fill_2 FILLER_13_825 ();
 sg13g2_fill_1 FILLER_13_851 ();
 sg13g2_decap_8 FILLER_13_857 ();
 sg13g2_decap_8 FILLER_13_864 ();
 sg13g2_fill_1 FILLER_13_871 ();
 sg13g2_fill_2 FILLER_13_894 ();
 sg13g2_fill_1 FILLER_13_896 ();
 sg13g2_fill_1 FILLER_13_917 ();
 sg13g2_decap_4 FILLER_13_924 ();
 sg13g2_fill_1 FILLER_13_949 ();
 sg13g2_fill_1 FILLER_13_955 ();
 sg13g2_fill_2 FILLER_13_968 ();
 sg13g2_decap_4 FILLER_13_985 ();
 sg13g2_decap_8 FILLER_13_1001 ();
 sg13g2_decap_4 FILLER_13_1008 ();
 sg13g2_fill_2 FILLER_13_1012 ();
 sg13g2_fill_2 FILLER_13_1038 ();
 sg13g2_fill_1 FILLER_13_1040 ();
 sg13g2_fill_1 FILLER_13_1062 ();
 sg13g2_decap_4 FILLER_13_1077 ();
 sg13g2_fill_2 FILLER_13_1089 ();
 sg13g2_fill_1 FILLER_13_1091 ();
 sg13g2_fill_1 FILLER_13_1099 ();
 sg13g2_decap_8 FILLER_13_1121 ();
 sg13g2_decap_8 FILLER_13_1128 ();
 sg13g2_decap_8 FILLER_13_1135 ();
 sg13g2_decap_8 FILLER_13_1142 ();
 sg13g2_decap_8 FILLER_13_1149 ();
 sg13g2_decap_8 FILLER_13_1156 ();
 sg13g2_decap_8 FILLER_13_1163 ();
 sg13g2_decap_8 FILLER_13_1170 ();
 sg13g2_decap_8 FILLER_13_1177 ();
 sg13g2_decap_8 FILLER_13_1184 ();
 sg13g2_decap_8 FILLER_13_1191 ();
 sg13g2_decap_8 FILLER_13_1198 ();
 sg13g2_decap_8 FILLER_13_1205 ();
 sg13g2_decap_8 FILLER_13_1212 ();
 sg13g2_decap_8 FILLER_13_1219 ();
 sg13g2_decap_8 FILLER_13_1226 ();
 sg13g2_decap_8 FILLER_13_1233 ();
 sg13g2_decap_8 FILLER_13_1240 ();
 sg13g2_decap_8 FILLER_13_1247 ();
 sg13g2_decap_8 FILLER_13_1254 ();
 sg13g2_decap_8 FILLER_13_1261 ();
 sg13g2_decap_8 FILLER_13_1268 ();
 sg13g2_decap_8 FILLER_13_1275 ();
 sg13g2_decap_8 FILLER_13_1282 ();
 sg13g2_decap_8 FILLER_13_1289 ();
 sg13g2_decap_8 FILLER_13_1296 ();
 sg13g2_decap_8 FILLER_13_1303 ();
 sg13g2_decap_8 FILLER_13_1310 ();
 sg13g2_decap_8 FILLER_13_1317 ();
 sg13g2_decap_8 FILLER_13_1324 ();
 sg13g2_decap_8 FILLER_13_1331 ();
 sg13g2_decap_8 FILLER_13_1338 ();
 sg13g2_decap_8 FILLER_13_1345 ();
 sg13g2_decap_8 FILLER_13_1352 ();
 sg13g2_decap_8 FILLER_13_1359 ();
 sg13g2_decap_8 FILLER_13_1366 ();
 sg13g2_decap_8 FILLER_13_1373 ();
 sg13g2_decap_8 FILLER_13_1380 ();
 sg13g2_decap_8 FILLER_13_1387 ();
 sg13g2_decap_8 FILLER_13_1394 ();
 sg13g2_decap_8 FILLER_13_1401 ();
 sg13g2_decap_8 FILLER_13_1408 ();
 sg13g2_decap_8 FILLER_13_1415 ();
 sg13g2_decap_8 FILLER_13_1422 ();
 sg13g2_decap_8 FILLER_13_1429 ();
 sg13g2_decap_8 FILLER_13_1436 ();
 sg13g2_decap_8 FILLER_13_1443 ();
 sg13g2_decap_8 FILLER_13_1450 ();
 sg13g2_decap_8 FILLER_13_1457 ();
 sg13g2_decap_8 FILLER_13_1464 ();
 sg13g2_decap_8 FILLER_13_1471 ();
 sg13g2_decap_8 FILLER_13_1478 ();
 sg13g2_decap_8 FILLER_13_1485 ();
 sg13g2_decap_8 FILLER_13_1492 ();
 sg13g2_decap_8 FILLER_13_1499 ();
 sg13g2_decap_8 FILLER_13_1506 ();
 sg13g2_decap_8 FILLER_13_1513 ();
 sg13g2_decap_8 FILLER_13_1520 ();
 sg13g2_decap_8 FILLER_13_1527 ();
 sg13g2_decap_8 FILLER_13_1534 ();
 sg13g2_decap_8 FILLER_13_1541 ();
 sg13g2_decap_8 FILLER_13_1548 ();
 sg13g2_decap_8 FILLER_13_1555 ();
 sg13g2_decap_8 FILLER_13_1562 ();
 sg13g2_decap_8 FILLER_13_1569 ();
 sg13g2_decap_8 FILLER_13_1576 ();
 sg13g2_decap_8 FILLER_13_1583 ();
 sg13g2_decap_8 FILLER_13_1590 ();
 sg13g2_decap_8 FILLER_13_1597 ();
 sg13g2_decap_8 FILLER_13_1604 ();
 sg13g2_decap_8 FILLER_13_1611 ();
 sg13g2_decap_8 FILLER_13_1618 ();
 sg13g2_decap_8 FILLER_13_1625 ();
 sg13g2_decap_8 FILLER_13_1632 ();
 sg13g2_decap_8 FILLER_13_1639 ();
 sg13g2_decap_8 FILLER_13_1646 ();
 sg13g2_decap_8 FILLER_13_1653 ();
 sg13g2_decap_8 FILLER_13_1660 ();
 sg13g2_decap_8 FILLER_13_1667 ();
 sg13g2_decap_8 FILLER_13_1674 ();
 sg13g2_decap_8 FILLER_13_1681 ();
 sg13g2_decap_8 FILLER_13_1688 ();
 sg13g2_decap_8 FILLER_13_1695 ();
 sg13g2_decap_8 FILLER_13_1702 ();
 sg13g2_decap_8 FILLER_13_1709 ();
 sg13g2_decap_8 FILLER_13_1716 ();
 sg13g2_decap_8 FILLER_13_1723 ();
 sg13g2_decap_8 FILLER_13_1730 ();
 sg13g2_decap_8 FILLER_13_1737 ();
 sg13g2_decap_8 FILLER_13_1744 ();
 sg13g2_decap_8 FILLER_13_1751 ();
 sg13g2_decap_8 FILLER_13_1758 ();
 sg13g2_fill_2 FILLER_13_1765 ();
 sg13g2_fill_1 FILLER_13_1767 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_fill_1 FILLER_14_42 ();
 sg13g2_fill_2 FILLER_14_93 ();
 sg13g2_fill_2 FILLER_14_100 ();
 sg13g2_fill_2 FILLER_14_129 ();
 sg13g2_fill_2 FILLER_14_144 ();
 sg13g2_fill_2 FILLER_14_183 ();
 sg13g2_decap_4 FILLER_14_190 ();
 sg13g2_fill_1 FILLER_14_194 ();
 sg13g2_fill_1 FILLER_14_200 ();
 sg13g2_fill_1 FILLER_14_224 ();
 sg13g2_fill_2 FILLER_14_254 ();
 sg13g2_decap_4 FILLER_14_265 ();
 sg13g2_fill_2 FILLER_14_269 ();
 sg13g2_fill_2 FILLER_14_302 ();
 sg13g2_fill_1 FILLER_14_304 ();
 sg13g2_fill_2 FILLER_14_323 ();
 sg13g2_fill_2 FILLER_14_362 ();
 sg13g2_fill_2 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_421 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_fill_2 FILLER_14_441 ();
 sg13g2_fill_1 FILLER_14_443 ();
 sg13g2_fill_2 FILLER_14_449 ();
 sg13g2_decap_4 FILLER_14_499 ();
 sg13g2_fill_2 FILLER_14_503 ();
 sg13g2_fill_2 FILLER_14_538 ();
 sg13g2_fill_1 FILLER_14_540 ();
 sg13g2_fill_2 FILLER_14_549 ();
 sg13g2_decap_8 FILLER_14_573 ();
 sg13g2_decap_8 FILLER_14_580 ();
 sg13g2_fill_2 FILLER_14_587 ();
 sg13g2_fill_1 FILLER_14_589 ();
 sg13g2_fill_1 FILLER_14_624 ();
 sg13g2_decap_8 FILLER_14_646 ();
 sg13g2_fill_2 FILLER_14_653 ();
 sg13g2_fill_2 FILLER_14_664 ();
 sg13g2_fill_1 FILLER_14_673 ();
 sg13g2_decap_8 FILLER_14_690 ();
 sg13g2_fill_1 FILLER_14_697 ();
 sg13g2_decap_8 FILLER_14_710 ();
 sg13g2_fill_2 FILLER_14_717 ();
 sg13g2_fill_1 FILLER_14_719 ();
 sg13g2_decap_4 FILLER_14_724 ();
 sg13g2_fill_2 FILLER_14_728 ();
 sg13g2_fill_2 FILLER_14_750 ();
 sg13g2_fill_2 FILLER_14_763 ();
 sg13g2_decap_4 FILLER_14_775 ();
 sg13g2_fill_1 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_fill_1 FILLER_14_805 ();
 sg13g2_fill_1 FILLER_14_813 ();
 sg13g2_fill_1 FILLER_14_829 ();
 sg13g2_decap_8 FILLER_14_852 ();
 sg13g2_decap_8 FILLER_14_863 ();
 sg13g2_decap_8 FILLER_14_888 ();
 sg13g2_fill_2 FILLER_14_895 ();
 sg13g2_fill_2 FILLER_14_966 ();
 sg13g2_decap_8 FILLER_14_978 ();
 sg13g2_decap_4 FILLER_14_990 ();
 sg13g2_fill_2 FILLER_14_994 ();
 sg13g2_fill_2 FILLER_14_1012 ();
 sg13g2_fill_1 FILLER_14_1014 ();
 sg13g2_fill_2 FILLER_14_1034 ();
 sg13g2_decap_8 FILLER_14_1067 ();
 sg13g2_fill_2 FILLER_14_1074 ();
 sg13g2_fill_1 FILLER_14_1085 ();
 sg13g2_fill_1 FILLER_14_1091 ();
 sg13g2_fill_1 FILLER_14_1097 ();
 sg13g2_decap_8 FILLER_14_1115 ();
 sg13g2_decap_8 FILLER_14_1122 ();
 sg13g2_decap_8 FILLER_14_1129 ();
 sg13g2_decap_8 FILLER_14_1136 ();
 sg13g2_decap_8 FILLER_14_1143 ();
 sg13g2_decap_8 FILLER_14_1150 ();
 sg13g2_decap_8 FILLER_14_1157 ();
 sg13g2_decap_8 FILLER_14_1164 ();
 sg13g2_decap_8 FILLER_14_1171 ();
 sg13g2_decap_8 FILLER_14_1178 ();
 sg13g2_decap_8 FILLER_14_1185 ();
 sg13g2_decap_8 FILLER_14_1192 ();
 sg13g2_decap_8 FILLER_14_1199 ();
 sg13g2_decap_8 FILLER_14_1206 ();
 sg13g2_decap_8 FILLER_14_1213 ();
 sg13g2_decap_8 FILLER_14_1220 ();
 sg13g2_decap_8 FILLER_14_1227 ();
 sg13g2_decap_8 FILLER_14_1234 ();
 sg13g2_decap_8 FILLER_14_1241 ();
 sg13g2_decap_8 FILLER_14_1248 ();
 sg13g2_decap_8 FILLER_14_1255 ();
 sg13g2_decap_8 FILLER_14_1262 ();
 sg13g2_decap_8 FILLER_14_1269 ();
 sg13g2_decap_8 FILLER_14_1276 ();
 sg13g2_decap_8 FILLER_14_1283 ();
 sg13g2_decap_8 FILLER_14_1290 ();
 sg13g2_decap_8 FILLER_14_1297 ();
 sg13g2_decap_8 FILLER_14_1304 ();
 sg13g2_decap_8 FILLER_14_1311 ();
 sg13g2_decap_8 FILLER_14_1318 ();
 sg13g2_decap_8 FILLER_14_1325 ();
 sg13g2_decap_8 FILLER_14_1332 ();
 sg13g2_decap_8 FILLER_14_1339 ();
 sg13g2_decap_8 FILLER_14_1346 ();
 sg13g2_decap_8 FILLER_14_1353 ();
 sg13g2_decap_8 FILLER_14_1360 ();
 sg13g2_decap_8 FILLER_14_1367 ();
 sg13g2_decap_8 FILLER_14_1374 ();
 sg13g2_decap_8 FILLER_14_1381 ();
 sg13g2_decap_8 FILLER_14_1388 ();
 sg13g2_decap_8 FILLER_14_1395 ();
 sg13g2_decap_8 FILLER_14_1402 ();
 sg13g2_decap_8 FILLER_14_1409 ();
 sg13g2_decap_8 FILLER_14_1416 ();
 sg13g2_decap_8 FILLER_14_1423 ();
 sg13g2_decap_8 FILLER_14_1430 ();
 sg13g2_decap_8 FILLER_14_1437 ();
 sg13g2_decap_8 FILLER_14_1444 ();
 sg13g2_decap_8 FILLER_14_1451 ();
 sg13g2_decap_8 FILLER_14_1458 ();
 sg13g2_decap_8 FILLER_14_1465 ();
 sg13g2_decap_8 FILLER_14_1472 ();
 sg13g2_decap_8 FILLER_14_1479 ();
 sg13g2_decap_8 FILLER_14_1486 ();
 sg13g2_decap_8 FILLER_14_1493 ();
 sg13g2_decap_8 FILLER_14_1500 ();
 sg13g2_decap_8 FILLER_14_1507 ();
 sg13g2_decap_8 FILLER_14_1514 ();
 sg13g2_decap_8 FILLER_14_1521 ();
 sg13g2_decap_8 FILLER_14_1528 ();
 sg13g2_decap_8 FILLER_14_1535 ();
 sg13g2_decap_8 FILLER_14_1542 ();
 sg13g2_decap_8 FILLER_14_1549 ();
 sg13g2_decap_8 FILLER_14_1556 ();
 sg13g2_decap_8 FILLER_14_1563 ();
 sg13g2_decap_8 FILLER_14_1570 ();
 sg13g2_decap_8 FILLER_14_1577 ();
 sg13g2_decap_8 FILLER_14_1584 ();
 sg13g2_decap_8 FILLER_14_1591 ();
 sg13g2_decap_8 FILLER_14_1598 ();
 sg13g2_decap_8 FILLER_14_1605 ();
 sg13g2_decap_8 FILLER_14_1612 ();
 sg13g2_decap_8 FILLER_14_1619 ();
 sg13g2_decap_8 FILLER_14_1626 ();
 sg13g2_decap_8 FILLER_14_1633 ();
 sg13g2_decap_8 FILLER_14_1640 ();
 sg13g2_decap_8 FILLER_14_1647 ();
 sg13g2_decap_8 FILLER_14_1654 ();
 sg13g2_decap_8 FILLER_14_1661 ();
 sg13g2_decap_8 FILLER_14_1668 ();
 sg13g2_decap_8 FILLER_14_1675 ();
 sg13g2_decap_8 FILLER_14_1682 ();
 sg13g2_decap_8 FILLER_14_1689 ();
 sg13g2_decap_8 FILLER_14_1696 ();
 sg13g2_decap_8 FILLER_14_1703 ();
 sg13g2_decap_8 FILLER_14_1710 ();
 sg13g2_decap_8 FILLER_14_1717 ();
 sg13g2_decap_8 FILLER_14_1724 ();
 sg13g2_decap_8 FILLER_14_1731 ();
 sg13g2_decap_8 FILLER_14_1738 ();
 sg13g2_decap_8 FILLER_14_1745 ();
 sg13g2_decap_8 FILLER_14_1752 ();
 sg13g2_decap_8 FILLER_14_1759 ();
 sg13g2_fill_2 FILLER_14_1766 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_109 ();
 sg13g2_fill_1 FILLER_15_118 ();
 sg13g2_fill_2 FILLER_15_124 ();
 sg13g2_fill_2 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_156 ();
 sg13g2_fill_1 FILLER_15_166 ();
 sg13g2_fill_2 FILLER_15_179 ();
 sg13g2_fill_1 FILLER_15_198 ();
 sg13g2_fill_2 FILLER_15_204 ();
 sg13g2_fill_1 FILLER_15_206 ();
 sg13g2_fill_2 FILLER_15_228 ();
 sg13g2_fill_1 FILLER_15_230 ();
 sg13g2_fill_2 FILLER_15_324 ();
 sg13g2_fill_1 FILLER_15_326 ();
 sg13g2_fill_2 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_334 ();
 sg13g2_fill_2 FILLER_15_359 ();
 sg13g2_fill_2 FILLER_15_366 ();
 sg13g2_fill_1 FILLER_15_368 ();
 sg13g2_decap_4 FILLER_15_408 ();
 sg13g2_fill_1 FILLER_15_412 ();
 sg13g2_decap_4 FILLER_15_448 ();
 sg13g2_fill_1 FILLER_15_467 ();
 sg13g2_fill_1 FILLER_15_471 ();
 sg13g2_fill_2 FILLER_15_487 ();
 sg13g2_decap_8 FILLER_15_505 ();
 sg13g2_decap_4 FILLER_15_512 ();
 sg13g2_fill_1 FILLER_15_516 ();
 sg13g2_decap_8 FILLER_15_527 ();
 sg13g2_decap_8 FILLER_15_534 ();
 sg13g2_decap_4 FILLER_15_541 ();
 sg13g2_fill_1 FILLER_15_545 ();
 sg13g2_fill_1 FILLER_15_578 ();
 sg13g2_decap_4 FILLER_15_587 ();
 sg13g2_fill_2 FILLER_15_602 ();
 sg13g2_fill_2 FILLER_15_618 ();
 sg13g2_fill_1 FILLER_15_620 ();
 sg13g2_fill_2 FILLER_15_636 ();
 sg13g2_fill_1 FILLER_15_638 ();
 sg13g2_decap_8 FILLER_15_652 ();
 sg13g2_fill_2 FILLER_15_701 ();
 sg13g2_decap_8 FILLER_15_726 ();
 sg13g2_fill_2 FILLER_15_733 ();
 sg13g2_fill_1 FILLER_15_735 ();
 sg13g2_fill_2 FILLER_15_740 ();
 sg13g2_decap_4 FILLER_15_754 ();
 sg13g2_decap_4 FILLER_15_762 ();
 sg13g2_decap_4 FILLER_15_775 ();
 sg13g2_fill_1 FILLER_15_779 ();
 sg13g2_fill_2 FILLER_15_790 ();
 sg13g2_decap_4 FILLER_15_837 ();
 sg13g2_fill_1 FILLER_15_855 ();
 sg13g2_fill_1 FILLER_15_863 ();
 sg13g2_fill_2 FILLER_15_879 ();
 sg13g2_fill_1 FILLER_15_881 ();
 sg13g2_fill_1 FILLER_15_926 ();
 sg13g2_fill_2 FILLER_15_938 ();
 sg13g2_fill_2 FILLER_15_944 ();
 sg13g2_fill_1 FILLER_15_961 ();
 sg13g2_decap_4 FILLER_15_971 ();
 sg13g2_fill_2 FILLER_15_975 ();
 sg13g2_fill_1 FILLER_15_981 ();
 sg13g2_fill_2 FILLER_15_997 ();
 sg13g2_decap_4 FILLER_15_1016 ();
 sg13g2_fill_1 FILLER_15_1020 ();
 sg13g2_fill_2 FILLER_15_1034 ();
 sg13g2_fill_1 FILLER_15_1036 ();
 sg13g2_fill_2 FILLER_15_1058 ();
 sg13g2_fill_1 FILLER_15_1060 ();
 sg13g2_fill_2 FILLER_15_1067 ();
 sg13g2_fill_1 FILLER_15_1069 ();
 sg13g2_fill_2 FILLER_15_1074 ();
 sg13g2_fill_1 FILLER_15_1096 ();
 sg13g2_decap_8 FILLER_15_1116 ();
 sg13g2_decap_8 FILLER_15_1123 ();
 sg13g2_decap_8 FILLER_15_1130 ();
 sg13g2_decap_8 FILLER_15_1137 ();
 sg13g2_decap_8 FILLER_15_1144 ();
 sg13g2_decap_8 FILLER_15_1151 ();
 sg13g2_decap_8 FILLER_15_1158 ();
 sg13g2_decap_8 FILLER_15_1165 ();
 sg13g2_decap_8 FILLER_15_1172 ();
 sg13g2_decap_8 FILLER_15_1179 ();
 sg13g2_decap_8 FILLER_15_1186 ();
 sg13g2_decap_8 FILLER_15_1193 ();
 sg13g2_decap_8 FILLER_15_1200 ();
 sg13g2_decap_8 FILLER_15_1207 ();
 sg13g2_decap_8 FILLER_15_1214 ();
 sg13g2_decap_8 FILLER_15_1221 ();
 sg13g2_decap_8 FILLER_15_1228 ();
 sg13g2_decap_8 FILLER_15_1235 ();
 sg13g2_decap_8 FILLER_15_1242 ();
 sg13g2_decap_8 FILLER_15_1249 ();
 sg13g2_decap_8 FILLER_15_1256 ();
 sg13g2_decap_8 FILLER_15_1263 ();
 sg13g2_decap_8 FILLER_15_1270 ();
 sg13g2_decap_8 FILLER_15_1277 ();
 sg13g2_decap_8 FILLER_15_1284 ();
 sg13g2_decap_8 FILLER_15_1291 ();
 sg13g2_decap_8 FILLER_15_1298 ();
 sg13g2_decap_8 FILLER_15_1305 ();
 sg13g2_decap_8 FILLER_15_1312 ();
 sg13g2_decap_8 FILLER_15_1319 ();
 sg13g2_decap_8 FILLER_15_1326 ();
 sg13g2_decap_8 FILLER_15_1333 ();
 sg13g2_decap_8 FILLER_15_1340 ();
 sg13g2_decap_8 FILLER_15_1347 ();
 sg13g2_decap_8 FILLER_15_1354 ();
 sg13g2_decap_8 FILLER_15_1361 ();
 sg13g2_decap_8 FILLER_15_1368 ();
 sg13g2_decap_8 FILLER_15_1375 ();
 sg13g2_decap_8 FILLER_15_1382 ();
 sg13g2_decap_8 FILLER_15_1389 ();
 sg13g2_decap_8 FILLER_15_1396 ();
 sg13g2_decap_8 FILLER_15_1403 ();
 sg13g2_decap_8 FILLER_15_1410 ();
 sg13g2_decap_8 FILLER_15_1417 ();
 sg13g2_decap_8 FILLER_15_1424 ();
 sg13g2_decap_8 FILLER_15_1431 ();
 sg13g2_decap_8 FILLER_15_1438 ();
 sg13g2_decap_8 FILLER_15_1445 ();
 sg13g2_decap_8 FILLER_15_1452 ();
 sg13g2_decap_8 FILLER_15_1459 ();
 sg13g2_decap_8 FILLER_15_1466 ();
 sg13g2_decap_8 FILLER_15_1473 ();
 sg13g2_decap_8 FILLER_15_1480 ();
 sg13g2_decap_8 FILLER_15_1487 ();
 sg13g2_decap_8 FILLER_15_1494 ();
 sg13g2_decap_8 FILLER_15_1501 ();
 sg13g2_decap_8 FILLER_15_1508 ();
 sg13g2_decap_8 FILLER_15_1515 ();
 sg13g2_decap_8 FILLER_15_1522 ();
 sg13g2_decap_8 FILLER_15_1529 ();
 sg13g2_decap_8 FILLER_15_1536 ();
 sg13g2_decap_8 FILLER_15_1543 ();
 sg13g2_decap_8 FILLER_15_1550 ();
 sg13g2_decap_8 FILLER_15_1557 ();
 sg13g2_decap_8 FILLER_15_1564 ();
 sg13g2_decap_8 FILLER_15_1571 ();
 sg13g2_decap_8 FILLER_15_1578 ();
 sg13g2_decap_8 FILLER_15_1585 ();
 sg13g2_decap_8 FILLER_15_1592 ();
 sg13g2_decap_8 FILLER_15_1599 ();
 sg13g2_decap_8 FILLER_15_1606 ();
 sg13g2_decap_8 FILLER_15_1613 ();
 sg13g2_decap_8 FILLER_15_1620 ();
 sg13g2_decap_8 FILLER_15_1627 ();
 sg13g2_decap_8 FILLER_15_1634 ();
 sg13g2_decap_8 FILLER_15_1641 ();
 sg13g2_decap_8 FILLER_15_1648 ();
 sg13g2_decap_8 FILLER_15_1655 ();
 sg13g2_decap_8 FILLER_15_1662 ();
 sg13g2_decap_8 FILLER_15_1669 ();
 sg13g2_decap_8 FILLER_15_1676 ();
 sg13g2_decap_8 FILLER_15_1683 ();
 sg13g2_decap_8 FILLER_15_1690 ();
 sg13g2_decap_8 FILLER_15_1697 ();
 sg13g2_decap_8 FILLER_15_1704 ();
 sg13g2_decap_8 FILLER_15_1711 ();
 sg13g2_decap_8 FILLER_15_1718 ();
 sg13g2_decap_8 FILLER_15_1725 ();
 sg13g2_decap_8 FILLER_15_1732 ();
 sg13g2_decap_8 FILLER_15_1739 ();
 sg13g2_decap_8 FILLER_15_1746 ();
 sg13g2_decap_8 FILLER_15_1753 ();
 sg13g2_decap_8 FILLER_15_1760 ();
 sg13g2_fill_1 FILLER_15_1767 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_23 ();
 sg13g2_fill_2 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_44 ();
 sg13g2_fill_2 FILLER_16_50 ();
 sg13g2_fill_1 FILLER_16_52 ();
 sg13g2_fill_2 FILLER_16_62 ();
 sg13g2_fill_1 FILLER_16_69 ();
 sg13g2_fill_2 FILLER_16_76 ();
 sg13g2_fill_1 FILLER_16_88 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_fill_2 FILLER_16_115 ();
 sg13g2_fill_2 FILLER_16_142 ();
 sg13g2_fill_2 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_216 ();
 sg13g2_fill_2 FILLER_16_230 ();
 sg13g2_fill_2 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_269 ();
 sg13g2_fill_1 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_decap_4 FILLER_16_305 ();
 sg13g2_fill_1 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_4 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_fill_2 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_365 ();
 sg13g2_decap_4 FILLER_16_397 ();
 sg13g2_fill_1 FILLER_16_401 ();
 sg13g2_fill_2 FILLER_16_418 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_451 ();
 sg13g2_decap_4 FILLER_16_458 ();
 sg13g2_decap_4 FILLER_16_482 ();
 sg13g2_fill_2 FILLER_16_512 ();
 sg13g2_fill_1 FILLER_16_519 ();
 sg13g2_decap_4 FILLER_16_544 ();
 sg13g2_fill_2 FILLER_16_548 ();
 sg13g2_fill_2 FILLER_16_560 ();
 sg13g2_fill_2 FILLER_16_571 ();
 sg13g2_decap_8 FILLER_16_586 ();
 sg13g2_decap_4 FILLER_16_593 ();
 sg13g2_fill_1 FILLER_16_597 ();
 sg13g2_fill_1 FILLER_16_618 ();
 sg13g2_decap_4 FILLER_16_628 ();
 sg13g2_fill_1 FILLER_16_632 ();
 sg13g2_fill_2 FILLER_16_647 ();
 sg13g2_fill_2 FILLER_16_662 ();
 sg13g2_fill_1 FILLER_16_664 ();
 sg13g2_decap_8 FILLER_16_670 ();
 sg13g2_decap_8 FILLER_16_699 ();
 sg13g2_decap_4 FILLER_16_706 ();
 sg13g2_fill_2 FILLER_16_750 ();
 sg13g2_decap_4 FILLER_16_756 ();
 sg13g2_fill_1 FILLER_16_760 ();
 sg13g2_decap_8 FILLER_16_769 ();
 sg13g2_fill_1 FILLER_16_776 ();
 sg13g2_fill_2 FILLER_16_815 ();
 sg13g2_decap_4 FILLER_16_835 ();
 sg13g2_fill_2 FILLER_16_869 ();
 sg13g2_fill_1 FILLER_16_871 ();
 sg13g2_decap_4 FILLER_16_893 ();
 sg13g2_decap_4 FILLER_16_901 ();
 sg13g2_fill_2 FILLER_16_905 ();
 sg13g2_decap_8 FILLER_16_917 ();
 sg13g2_decap_4 FILLER_16_924 ();
 sg13g2_fill_2 FILLER_16_928 ();
 sg13g2_decap_8 FILLER_16_944 ();
 sg13g2_fill_1 FILLER_16_951 ();
 sg13g2_fill_1 FILLER_16_1017 ();
 sg13g2_decap_8 FILLER_16_1023 ();
 sg13g2_decap_8 FILLER_16_1030 ();
 sg13g2_fill_1 FILLER_16_1037 ();
 sg13g2_decap_4 FILLER_16_1052 ();
 sg13g2_decap_8 FILLER_16_1080 ();
 sg13g2_fill_1 FILLER_16_1087 ();
 sg13g2_decap_8 FILLER_16_1108 ();
 sg13g2_decap_8 FILLER_16_1115 ();
 sg13g2_decap_8 FILLER_16_1122 ();
 sg13g2_decap_8 FILLER_16_1129 ();
 sg13g2_decap_8 FILLER_16_1136 ();
 sg13g2_decap_8 FILLER_16_1143 ();
 sg13g2_decap_8 FILLER_16_1150 ();
 sg13g2_decap_8 FILLER_16_1157 ();
 sg13g2_decap_8 FILLER_16_1164 ();
 sg13g2_decap_8 FILLER_16_1171 ();
 sg13g2_decap_8 FILLER_16_1178 ();
 sg13g2_decap_8 FILLER_16_1185 ();
 sg13g2_decap_8 FILLER_16_1192 ();
 sg13g2_decap_8 FILLER_16_1199 ();
 sg13g2_decap_8 FILLER_16_1206 ();
 sg13g2_decap_8 FILLER_16_1213 ();
 sg13g2_decap_8 FILLER_16_1220 ();
 sg13g2_decap_8 FILLER_16_1227 ();
 sg13g2_decap_8 FILLER_16_1234 ();
 sg13g2_decap_8 FILLER_16_1241 ();
 sg13g2_decap_8 FILLER_16_1248 ();
 sg13g2_decap_8 FILLER_16_1255 ();
 sg13g2_decap_8 FILLER_16_1262 ();
 sg13g2_decap_8 FILLER_16_1269 ();
 sg13g2_decap_8 FILLER_16_1276 ();
 sg13g2_decap_8 FILLER_16_1283 ();
 sg13g2_decap_8 FILLER_16_1290 ();
 sg13g2_decap_8 FILLER_16_1297 ();
 sg13g2_decap_8 FILLER_16_1304 ();
 sg13g2_decap_8 FILLER_16_1311 ();
 sg13g2_decap_8 FILLER_16_1318 ();
 sg13g2_decap_8 FILLER_16_1325 ();
 sg13g2_decap_8 FILLER_16_1332 ();
 sg13g2_decap_8 FILLER_16_1339 ();
 sg13g2_decap_8 FILLER_16_1346 ();
 sg13g2_decap_8 FILLER_16_1353 ();
 sg13g2_decap_8 FILLER_16_1360 ();
 sg13g2_decap_8 FILLER_16_1367 ();
 sg13g2_decap_8 FILLER_16_1374 ();
 sg13g2_decap_8 FILLER_16_1381 ();
 sg13g2_decap_8 FILLER_16_1388 ();
 sg13g2_decap_8 FILLER_16_1395 ();
 sg13g2_decap_8 FILLER_16_1402 ();
 sg13g2_decap_8 FILLER_16_1409 ();
 sg13g2_decap_8 FILLER_16_1416 ();
 sg13g2_decap_8 FILLER_16_1423 ();
 sg13g2_decap_8 FILLER_16_1430 ();
 sg13g2_decap_8 FILLER_16_1437 ();
 sg13g2_decap_8 FILLER_16_1444 ();
 sg13g2_decap_8 FILLER_16_1451 ();
 sg13g2_decap_8 FILLER_16_1458 ();
 sg13g2_decap_8 FILLER_16_1465 ();
 sg13g2_decap_8 FILLER_16_1472 ();
 sg13g2_decap_8 FILLER_16_1479 ();
 sg13g2_decap_8 FILLER_16_1486 ();
 sg13g2_decap_8 FILLER_16_1493 ();
 sg13g2_decap_8 FILLER_16_1500 ();
 sg13g2_decap_8 FILLER_16_1507 ();
 sg13g2_decap_8 FILLER_16_1514 ();
 sg13g2_decap_8 FILLER_16_1521 ();
 sg13g2_decap_8 FILLER_16_1528 ();
 sg13g2_decap_8 FILLER_16_1535 ();
 sg13g2_decap_8 FILLER_16_1542 ();
 sg13g2_decap_8 FILLER_16_1549 ();
 sg13g2_decap_8 FILLER_16_1556 ();
 sg13g2_decap_8 FILLER_16_1563 ();
 sg13g2_decap_8 FILLER_16_1570 ();
 sg13g2_decap_8 FILLER_16_1577 ();
 sg13g2_decap_8 FILLER_16_1584 ();
 sg13g2_decap_8 FILLER_16_1591 ();
 sg13g2_decap_8 FILLER_16_1598 ();
 sg13g2_decap_8 FILLER_16_1605 ();
 sg13g2_decap_8 FILLER_16_1612 ();
 sg13g2_decap_8 FILLER_16_1619 ();
 sg13g2_decap_8 FILLER_16_1626 ();
 sg13g2_decap_8 FILLER_16_1633 ();
 sg13g2_decap_8 FILLER_16_1640 ();
 sg13g2_decap_8 FILLER_16_1647 ();
 sg13g2_decap_8 FILLER_16_1654 ();
 sg13g2_decap_8 FILLER_16_1661 ();
 sg13g2_decap_8 FILLER_16_1668 ();
 sg13g2_decap_8 FILLER_16_1675 ();
 sg13g2_decap_8 FILLER_16_1682 ();
 sg13g2_decap_8 FILLER_16_1689 ();
 sg13g2_decap_8 FILLER_16_1696 ();
 sg13g2_decap_8 FILLER_16_1703 ();
 sg13g2_decap_8 FILLER_16_1710 ();
 sg13g2_decap_8 FILLER_16_1717 ();
 sg13g2_decap_8 FILLER_16_1724 ();
 sg13g2_decap_8 FILLER_16_1731 ();
 sg13g2_decap_8 FILLER_16_1738 ();
 sg13g2_decap_8 FILLER_16_1745 ();
 sg13g2_decap_8 FILLER_16_1752 ();
 sg13g2_decap_8 FILLER_16_1759 ();
 sg13g2_fill_2 FILLER_16_1766 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_53 ();
 sg13g2_fill_1 FILLER_17_99 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_fill_1 FILLER_17_173 ();
 sg13g2_fill_2 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_200 ();
 sg13g2_fill_2 FILLER_17_206 ();
 sg13g2_decap_8 FILLER_17_213 ();
 sg13g2_decap_4 FILLER_17_220 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_fill_2 FILLER_17_254 ();
 sg13g2_fill_1 FILLER_17_256 ();
 sg13g2_fill_2 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_327 ();
 sg13g2_decap_4 FILLER_17_331 ();
 sg13g2_fill_1 FILLER_17_335 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_decap_4 FILLER_17_348 ();
 sg13g2_fill_2 FILLER_17_355 ();
 sg13g2_fill_2 FILLER_17_362 ();
 sg13g2_fill_2 FILLER_17_382 ();
 sg13g2_fill_1 FILLER_17_384 ();
 sg13g2_decap_4 FILLER_17_390 ();
 sg13g2_fill_2 FILLER_17_394 ();
 sg13g2_decap_4 FILLER_17_401 ();
 sg13g2_fill_2 FILLER_17_421 ();
 sg13g2_fill_1 FILLER_17_423 ();
 sg13g2_fill_2 FILLER_17_445 ();
 sg13g2_fill_1 FILLER_17_447 ();
 sg13g2_fill_2 FILLER_17_453 ();
 sg13g2_fill_1 FILLER_17_464 ();
 sg13g2_fill_2 FILLER_17_489 ();
 sg13g2_fill_1 FILLER_17_491 ();
 sg13g2_fill_1 FILLER_17_497 ();
 sg13g2_fill_2 FILLER_17_501 ();
 sg13g2_fill_1 FILLER_17_503 ();
 sg13g2_fill_2 FILLER_17_509 ();
 sg13g2_fill_1 FILLER_17_511 ();
 sg13g2_decap_4 FILLER_17_522 ();
 sg13g2_decap_4 FILLER_17_531 ();
 sg13g2_fill_1 FILLER_17_535 ();
 sg13g2_decap_8 FILLER_17_541 ();
 sg13g2_fill_2 FILLER_17_548 ();
 sg13g2_fill_1 FILLER_17_550 ();
 sg13g2_fill_2 FILLER_17_570 ();
 sg13g2_fill_2 FILLER_17_580 ();
 sg13g2_fill_1 FILLER_17_596 ();
 sg13g2_decap_8 FILLER_17_601 ();
 sg13g2_fill_2 FILLER_17_623 ();
 sg13g2_fill_2 FILLER_17_648 ();
 sg13g2_fill_1 FILLER_17_659 ();
 sg13g2_decap_8 FILLER_17_669 ();
 sg13g2_fill_2 FILLER_17_676 ();
 sg13g2_fill_1 FILLER_17_678 ();
 sg13g2_fill_1 FILLER_17_704 ();
 sg13g2_fill_2 FILLER_17_710 ();
 sg13g2_fill_1 FILLER_17_712 ();
 sg13g2_fill_1 FILLER_17_725 ();
 sg13g2_decap_8 FILLER_17_746 ();
 sg13g2_fill_2 FILLER_17_753 ();
 sg13g2_decap_8 FILLER_17_765 ();
 sg13g2_fill_1 FILLER_17_772 ();
 sg13g2_fill_2 FILLER_17_785 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_4 FILLER_17_805 ();
 sg13g2_fill_2 FILLER_17_809 ();
 sg13g2_decap_8 FILLER_17_815 ();
 sg13g2_fill_2 FILLER_17_822 ();
 sg13g2_fill_2 FILLER_17_832 ();
 sg13g2_decap_8 FILLER_17_839 ();
 sg13g2_fill_2 FILLER_17_846 ();
 sg13g2_fill_2 FILLER_17_857 ();
 sg13g2_fill_1 FILLER_17_864 ();
 sg13g2_fill_1 FILLER_17_875 ();
 sg13g2_fill_2 FILLER_17_900 ();
 sg13g2_fill_1 FILLER_17_927 ();
 sg13g2_fill_1 FILLER_17_952 ();
 sg13g2_fill_2 FILLER_17_963 ();
 sg13g2_decap_8 FILLER_17_977 ();
 sg13g2_fill_2 FILLER_17_994 ();
 sg13g2_fill_1 FILLER_17_996 ();
 sg13g2_fill_2 FILLER_17_1007 ();
 sg13g2_decap_8 FILLER_17_1029 ();
 sg13g2_fill_2 FILLER_17_1036 ();
 sg13g2_decap_4 FILLER_17_1074 ();
 sg13g2_fill_1 FILLER_17_1078 ();
 sg13g2_fill_1 FILLER_17_1083 ();
 sg13g2_fill_2 FILLER_17_1088 ();
 sg13g2_decap_8 FILLER_17_1106 ();
 sg13g2_decap_8 FILLER_17_1113 ();
 sg13g2_decap_8 FILLER_17_1120 ();
 sg13g2_decap_8 FILLER_17_1127 ();
 sg13g2_decap_8 FILLER_17_1134 ();
 sg13g2_decap_8 FILLER_17_1141 ();
 sg13g2_decap_8 FILLER_17_1148 ();
 sg13g2_decap_8 FILLER_17_1155 ();
 sg13g2_decap_8 FILLER_17_1162 ();
 sg13g2_decap_8 FILLER_17_1169 ();
 sg13g2_decap_8 FILLER_17_1176 ();
 sg13g2_decap_8 FILLER_17_1183 ();
 sg13g2_decap_8 FILLER_17_1190 ();
 sg13g2_decap_8 FILLER_17_1197 ();
 sg13g2_decap_8 FILLER_17_1204 ();
 sg13g2_decap_8 FILLER_17_1211 ();
 sg13g2_decap_8 FILLER_17_1218 ();
 sg13g2_decap_8 FILLER_17_1225 ();
 sg13g2_decap_8 FILLER_17_1232 ();
 sg13g2_decap_8 FILLER_17_1239 ();
 sg13g2_decap_8 FILLER_17_1246 ();
 sg13g2_decap_8 FILLER_17_1253 ();
 sg13g2_decap_8 FILLER_17_1260 ();
 sg13g2_decap_8 FILLER_17_1267 ();
 sg13g2_decap_8 FILLER_17_1274 ();
 sg13g2_decap_8 FILLER_17_1281 ();
 sg13g2_decap_8 FILLER_17_1288 ();
 sg13g2_decap_8 FILLER_17_1295 ();
 sg13g2_decap_8 FILLER_17_1302 ();
 sg13g2_decap_8 FILLER_17_1309 ();
 sg13g2_decap_8 FILLER_17_1316 ();
 sg13g2_decap_8 FILLER_17_1323 ();
 sg13g2_decap_8 FILLER_17_1330 ();
 sg13g2_decap_8 FILLER_17_1337 ();
 sg13g2_decap_8 FILLER_17_1344 ();
 sg13g2_decap_8 FILLER_17_1351 ();
 sg13g2_decap_8 FILLER_17_1358 ();
 sg13g2_decap_8 FILLER_17_1365 ();
 sg13g2_decap_8 FILLER_17_1372 ();
 sg13g2_decap_8 FILLER_17_1379 ();
 sg13g2_decap_8 FILLER_17_1386 ();
 sg13g2_decap_8 FILLER_17_1393 ();
 sg13g2_decap_8 FILLER_17_1400 ();
 sg13g2_decap_8 FILLER_17_1407 ();
 sg13g2_decap_8 FILLER_17_1414 ();
 sg13g2_decap_8 FILLER_17_1421 ();
 sg13g2_decap_8 FILLER_17_1428 ();
 sg13g2_decap_8 FILLER_17_1435 ();
 sg13g2_decap_8 FILLER_17_1442 ();
 sg13g2_decap_8 FILLER_17_1449 ();
 sg13g2_decap_8 FILLER_17_1456 ();
 sg13g2_decap_8 FILLER_17_1463 ();
 sg13g2_decap_8 FILLER_17_1470 ();
 sg13g2_decap_8 FILLER_17_1477 ();
 sg13g2_decap_8 FILLER_17_1484 ();
 sg13g2_decap_8 FILLER_17_1491 ();
 sg13g2_decap_8 FILLER_17_1498 ();
 sg13g2_decap_8 FILLER_17_1505 ();
 sg13g2_decap_8 FILLER_17_1512 ();
 sg13g2_decap_8 FILLER_17_1519 ();
 sg13g2_decap_8 FILLER_17_1526 ();
 sg13g2_decap_8 FILLER_17_1533 ();
 sg13g2_decap_8 FILLER_17_1540 ();
 sg13g2_decap_8 FILLER_17_1547 ();
 sg13g2_decap_8 FILLER_17_1554 ();
 sg13g2_decap_8 FILLER_17_1561 ();
 sg13g2_decap_8 FILLER_17_1568 ();
 sg13g2_decap_8 FILLER_17_1575 ();
 sg13g2_decap_8 FILLER_17_1582 ();
 sg13g2_decap_8 FILLER_17_1589 ();
 sg13g2_decap_8 FILLER_17_1596 ();
 sg13g2_decap_8 FILLER_17_1603 ();
 sg13g2_decap_8 FILLER_17_1610 ();
 sg13g2_decap_8 FILLER_17_1617 ();
 sg13g2_decap_8 FILLER_17_1624 ();
 sg13g2_decap_8 FILLER_17_1631 ();
 sg13g2_decap_8 FILLER_17_1638 ();
 sg13g2_decap_8 FILLER_17_1645 ();
 sg13g2_decap_8 FILLER_17_1652 ();
 sg13g2_decap_8 FILLER_17_1659 ();
 sg13g2_decap_8 FILLER_17_1666 ();
 sg13g2_decap_8 FILLER_17_1673 ();
 sg13g2_decap_8 FILLER_17_1680 ();
 sg13g2_decap_8 FILLER_17_1687 ();
 sg13g2_decap_8 FILLER_17_1694 ();
 sg13g2_decap_8 FILLER_17_1701 ();
 sg13g2_decap_8 FILLER_17_1708 ();
 sg13g2_decap_8 FILLER_17_1715 ();
 sg13g2_decap_8 FILLER_17_1722 ();
 sg13g2_decap_8 FILLER_17_1729 ();
 sg13g2_decap_8 FILLER_17_1736 ();
 sg13g2_decap_8 FILLER_17_1743 ();
 sg13g2_decap_8 FILLER_17_1750 ();
 sg13g2_decap_8 FILLER_17_1757 ();
 sg13g2_decap_4 FILLER_17_1764 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_25 ();
 sg13g2_fill_2 FILLER_18_66 ();
 sg13g2_fill_2 FILLER_18_73 ();
 sg13g2_decap_4 FILLER_18_89 ();
 sg13g2_fill_2 FILLER_18_93 ();
 sg13g2_fill_2 FILLER_18_125 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_147 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_decap_8 FILLER_18_178 ();
 sg13g2_fill_2 FILLER_18_185 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_2 FILLER_18_201 ();
 sg13g2_fill_1 FILLER_18_214 ();
 sg13g2_decap_4 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_240 ();
 sg13g2_fill_1 FILLER_18_242 ();
 sg13g2_decap_4 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_258 ();
 sg13g2_decap_4 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_299 ();
 sg13g2_decap_4 FILLER_18_306 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_fill_2 FILLER_18_333 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_358 ();
 sg13g2_decap_4 FILLER_18_364 ();
 sg13g2_fill_2 FILLER_18_374 ();
 sg13g2_fill_1 FILLER_18_386 ();
 sg13g2_fill_2 FILLER_18_393 ();
 sg13g2_fill_1 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_412 ();
 sg13g2_decap_4 FILLER_18_419 ();
 sg13g2_decap_4 FILLER_18_458 ();
 sg13g2_fill_2 FILLER_18_467 ();
 sg13g2_fill_1 FILLER_18_474 ();
 sg13g2_decap_8 FILLER_18_486 ();
 sg13g2_fill_1 FILLER_18_497 ();
 sg13g2_fill_2 FILLER_18_502 ();
 sg13g2_decap_4 FILLER_18_512 ();
 sg13g2_fill_2 FILLER_18_536 ();
 sg13g2_fill_2 FILLER_18_541 ();
 sg13g2_fill_2 FILLER_18_555 ();
 sg13g2_fill_1 FILLER_18_557 ();
 sg13g2_fill_2 FILLER_18_564 ();
 sg13g2_fill_1 FILLER_18_566 ();
 sg13g2_decap_8 FILLER_18_607 ();
 sg13g2_decap_4 FILLER_18_614 ();
 sg13g2_fill_2 FILLER_18_618 ();
 sg13g2_decap_8 FILLER_18_640 ();
 sg13g2_decap_4 FILLER_18_647 ();
 sg13g2_fill_2 FILLER_18_674 ();
 sg13g2_fill_1 FILLER_18_681 ();
 sg13g2_fill_1 FILLER_18_689 ();
 sg13g2_fill_2 FILLER_18_705 ();
 sg13g2_fill_1 FILLER_18_707 ();
 sg13g2_decap_4 FILLER_18_713 ();
 sg13g2_decap_4 FILLER_18_747 ();
 sg13g2_fill_1 FILLER_18_751 ();
 sg13g2_fill_1 FILLER_18_802 ();
 sg13g2_fill_2 FILLER_18_823 ();
 sg13g2_decap_8 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_863 ();
 sg13g2_decap_4 FILLER_18_870 ();
 sg13g2_fill_2 FILLER_18_874 ();
 sg13g2_fill_1 FILLER_18_895 ();
 sg13g2_decap_8 FILLER_18_900 ();
 sg13g2_decap_8 FILLER_18_907 ();
 sg13g2_decap_8 FILLER_18_914 ();
 sg13g2_decap_8 FILLER_18_921 ();
 sg13g2_decap_4 FILLER_18_928 ();
 sg13g2_fill_1 FILLER_18_932 ();
 sg13g2_fill_2 FILLER_18_942 ();
 sg13g2_fill_1 FILLER_18_944 ();
 sg13g2_decap_8 FILLER_18_969 ();
 sg13g2_fill_2 FILLER_18_1014 ();
 sg13g2_fill_2 FILLER_18_1036 ();
 sg13g2_decap_8 FILLER_18_1048 ();
 sg13g2_fill_1 FILLER_18_1060 ();
 sg13g2_fill_2 FILLER_18_1066 ();
 sg13g2_fill_2 FILLER_18_1081 ();
 sg13g2_decap_8 FILLER_18_1106 ();
 sg13g2_decap_8 FILLER_18_1113 ();
 sg13g2_decap_8 FILLER_18_1120 ();
 sg13g2_decap_8 FILLER_18_1127 ();
 sg13g2_decap_8 FILLER_18_1134 ();
 sg13g2_decap_8 FILLER_18_1141 ();
 sg13g2_decap_8 FILLER_18_1148 ();
 sg13g2_decap_8 FILLER_18_1155 ();
 sg13g2_decap_8 FILLER_18_1162 ();
 sg13g2_decap_8 FILLER_18_1169 ();
 sg13g2_decap_8 FILLER_18_1176 ();
 sg13g2_decap_8 FILLER_18_1183 ();
 sg13g2_decap_8 FILLER_18_1190 ();
 sg13g2_decap_8 FILLER_18_1197 ();
 sg13g2_decap_8 FILLER_18_1204 ();
 sg13g2_decap_8 FILLER_18_1211 ();
 sg13g2_decap_8 FILLER_18_1218 ();
 sg13g2_decap_8 FILLER_18_1225 ();
 sg13g2_decap_8 FILLER_18_1232 ();
 sg13g2_decap_8 FILLER_18_1239 ();
 sg13g2_decap_8 FILLER_18_1246 ();
 sg13g2_decap_8 FILLER_18_1253 ();
 sg13g2_decap_8 FILLER_18_1260 ();
 sg13g2_decap_8 FILLER_18_1267 ();
 sg13g2_decap_8 FILLER_18_1274 ();
 sg13g2_decap_8 FILLER_18_1281 ();
 sg13g2_decap_8 FILLER_18_1288 ();
 sg13g2_decap_8 FILLER_18_1295 ();
 sg13g2_decap_8 FILLER_18_1302 ();
 sg13g2_decap_8 FILLER_18_1309 ();
 sg13g2_decap_8 FILLER_18_1316 ();
 sg13g2_decap_8 FILLER_18_1323 ();
 sg13g2_decap_8 FILLER_18_1330 ();
 sg13g2_decap_8 FILLER_18_1337 ();
 sg13g2_decap_8 FILLER_18_1344 ();
 sg13g2_decap_8 FILLER_18_1351 ();
 sg13g2_decap_8 FILLER_18_1358 ();
 sg13g2_decap_8 FILLER_18_1365 ();
 sg13g2_decap_8 FILLER_18_1372 ();
 sg13g2_decap_8 FILLER_18_1379 ();
 sg13g2_decap_8 FILLER_18_1386 ();
 sg13g2_decap_8 FILLER_18_1393 ();
 sg13g2_decap_8 FILLER_18_1400 ();
 sg13g2_decap_8 FILLER_18_1407 ();
 sg13g2_decap_8 FILLER_18_1414 ();
 sg13g2_decap_8 FILLER_18_1421 ();
 sg13g2_decap_8 FILLER_18_1428 ();
 sg13g2_decap_8 FILLER_18_1435 ();
 sg13g2_decap_8 FILLER_18_1442 ();
 sg13g2_decap_8 FILLER_18_1449 ();
 sg13g2_decap_8 FILLER_18_1456 ();
 sg13g2_decap_8 FILLER_18_1463 ();
 sg13g2_decap_8 FILLER_18_1470 ();
 sg13g2_decap_8 FILLER_18_1477 ();
 sg13g2_decap_8 FILLER_18_1484 ();
 sg13g2_decap_8 FILLER_18_1491 ();
 sg13g2_decap_8 FILLER_18_1498 ();
 sg13g2_decap_8 FILLER_18_1505 ();
 sg13g2_decap_8 FILLER_18_1512 ();
 sg13g2_decap_8 FILLER_18_1519 ();
 sg13g2_decap_8 FILLER_18_1526 ();
 sg13g2_decap_8 FILLER_18_1533 ();
 sg13g2_decap_8 FILLER_18_1540 ();
 sg13g2_decap_8 FILLER_18_1547 ();
 sg13g2_decap_8 FILLER_18_1554 ();
 sg13g2_decap_8 FILLER_18_1561 ();
 sg13g2_decap_8 FILLER_18_1568 ();
 sg13g2_decap_8 FILLER_18_1575 ();
 sg13g2_decap_8 FILLER_18_1582 ();
 sg13g2_decap_8 FILLER_18_1589 ();
 sg13g2_decap_8 FILLER_18_1596 ();
 sg13g2_decap_8 FILLER_18_1603 ();
 sg13g2_decap_8 FILLER_18_1610 ();
 sg13g2_decap_8 FILLER_18_1617 ();
 sg13g2_decap_8 FILLER_18_1624 ();
 sg13g2_decap_8 FILLER_18_1631 ();
 sg13g2_decap_8 FILLER_18_1638 ();
 sg13g2_decap_8 FILLER_18_1645 ();
 sg13g2_decap_8 FILLER_18_1652 ();
 sg13g2_decap_8 FILLER_18_1659 ();
 sg13g2_decap_8 FILLER_18_1666 ();
 sg13g2_decap_8 FILLER_18_1673 ();
 sg13g2_decap_8 FILLER_18_1680 ();
 sg13g2_decap_8 FILLER_18_1687 ();
 sg13g2_decap_8 FILLER_18_1694 ();
 sg13g2_decap_8 FILLER_18_1701 ();
 sg13g2_decap_8 FILLER_18_1708 ();
 sg13g2_decap_8 FILLER_18_1715 ();
 sg13g2_decap_8 FILLER_18_1722 ();
 sg13g2_decap_8 FILLER_18_1729 ();
 sg13g2_decap_8 FILLER_18_1736 ();
 sg13g2_decap_8 FILLER_18_1743 ();
 sg13g2_decap_8 FILLER_18_1750 ();
 sg13g2_decap_8 FILLER_18_1757 ();
 sg13g2_decap_4 FILLER_18_1764 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_4 FILLER_19_14 ();
 sg13g2_fill_1 FILLER_19_18 ();
 sg13g2_decap_4 FILLER_19_79 ();
 sg13g2_fill_1 FILLER_19_108 ();
 sg13g2_decap_8 FILLER_19_141 ();
 sg13g2_fill_2 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_160 ();
 sg13g2_decap_4 FILLER_19_172 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_fill_2 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_fill_2 FILLER_19_245 ();
 sg13g2_fill_2 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_fill_2 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_fill_1 FILLER_19_326 ();
 sg13g2_fill_2 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_366 ();
 sg13g2_fill_2 FILLER_19_375 ();
 sg13g2_fill_1 FILLER_19_377 ();
 sg13g2_fill_2 FILLER_19_393 ();
 sg13g2_fill_1 FILLER_19_395 ();
 sg13g2_fill_1 FILLER_19_440 ();
 sg13g2_decap_4 FILLER_19_449 ();
 sg13g2_decap_4 FILLER_19_510 ();
 sg13g2_fill_2 FILLER_19_538 ();
 sg13g2_fill_1 FILLER_19_540 ();
 sg13g2_decap_4 FILLER_19_550 ();
 sg13g2_fill_2 FILLER_19_554 ();
 sg13g2_fill_1 FILLER_19_566 ();
 sg13g2_fill_2 FILLER_19_571 ();
 sg13g2_fill_1 FILLER_19_573 ();
 sg13g2_fill_1 FILLER_19_588 ();
 sg13g2_decap_4 FILLER_19_592 ();
 sg13g2_fill_1 FILLER_19_596 ();
 sg13g2_decap_4 FILLER_19_601 ();
 sg13g2_fill_1 FILLER_19_605 ();
 sg13g2_fill_2 FILLER_19_626 ();
 sg13g2_fill_1 FILLER_19_628 ();
 sg13g2_fill_2 FILLER_19_639 ();
 sg13g2_decap_4 FILLER_19_650 ();
 sg13g2_fill_1 FILLER_19_654 ();
 sg13g2_fill_1 FILLER_19_665 ();
 sg13g2_fill_2 FILLER_19_703 ();
 sg13g2_fill_1 FILLER_19_705 ();
 sg13g2_decap_4 FILLER_19_726 ();
 sg13g2_fill_1 FILLER_19_730 ();
 sg13g2_decap_8 FILLER_19_736 ();
 sg13g2_decap_8 FILLER_19_743 ();
 sg13g2_fill_1 FILLER_19_750 ();
 sg13g2_decap_4 FILLER_19_786 ();
 sg13g2_fill_2 FILLER_19_810 ();
 sg13g2_fill_2 FILLER_19_822 ();
 sg13g2_decap_8 FILLER_19_862 ();
 sg13g2_fill_2 FILLER_19_872 ();
 sg13g2_decap_4 FILLER_19_880 ();
 sg13g2_fill_1 FILLER_19_884 ();
 sg13g2_decap_4 FILLER_19_918 ();
 sg13g2_fill_1 FILLER_19_922 ();
 sg13g2_fill_2 FILLER_19_953 ();
 sg13g2_fill_1 FILLER_19_955 ();
 sg13g2_fill_2 FILLER_19_966 ();
 sg13g2_decap_8 FILLER_19_988 ();
 sg13g2_decap_4 FILLER_19_995 ();
 sg13g2_fill_2 FILLER_19_999 ();
 sg13g2_decap_8 FILLER_19_1011 ();
 sg13g2_decap_8 FILLER_19_1038 ();
 sg13g2_fill_1 FILLER_19_1050 ();
 sg13g2_decap_4 FILLER_19_1081 ();
 sg13g2_decap_8 FILLER_19_1103 ();
 sg13g2_decap_8 FILLER_19_1110 ();
 sg13g2_decap_8 FILLER_19_1117 ();
 sg13g2_decap_8 FILLER_19_1124 ();
 sg13g2_decap_8 FILLER_19_1131 ();
 sg13g2_decap_8 FILLER_19_1138 ();
 sg13g2_decap_8 FILLER_19_1145 ();
 sg13g2_decap_8 FILLER_19_1152 ();
 sg13g2_decap_8 FILLER_19_1159 ();
 sg13g2_decap_8 FILLER_19_1166 ();
 sg13g2_decap_8 FILLER_19_1173 ();
 sg13g2_decap_8 FILLER_19_1180 ();
 sg13g2_decap_8 FILLER_19_1187 ();
 sg13g2_decap_8 FILLER_19_1194 ();
 sg13g2_decap_8 FILLER_19_1201 ();
 sg13g2_decap_8 FILLER_19_1208 ();
 sg13g2_decap_8 FILLER_19_1215 ();
 sg13g2_decap_8 FILLER_19_1222 ();
 sg13g2_decap_8 FILLER_19_1229 ();
 sg13g2_decap_8 FILLER_19_1236 ();
 sg13g2_decap_8 FILLER_19_1243 ();
 sg13g2_decap_8 FILLER_19_1250 ();
 sg13g2_decap_8 FILLER_19_1257 ();
 sg13g2_decap_8 FILLER_19_1264 ();
 sg13g2_decap_8 FILLER_19_1271 ();
 sg13g2_decap_8 FILLER_19_1278 ();
 sg13g2_decap_8 FILLER_19_1285 ();
 sg13g2_decap_8 FILLER_19_1292 ();
 sg13g2_decap_8 FILLER_19_1299 ();
 sg13g2_decap_8 FILLER_19_1306 ();
 sg13g2_decap_8 FILLER_19_1313 ();
 sg13g2_decap_8 FILLER_19_1320 ();
 sg13g2_decap_8 FILLER_19_1327 ();
 sg13g2_decap_8 FILLER_19_1334 ();
 sg13g2_decap_8 FILLER_19_1341 ();
 sg13g2_decap_8 FILLER_19_1348 ();
 sg13g2_decap_8 FILLER_19_1355 ();
 sg13g2_decap_8 FILLER_19_1362 ();
 sg13g2_decap_8 FILLER_19_1369 ();
 sg13g2_decap_8 FILLER_19_1376 ();
 sg13g2_decap_8 FILLER_19_1383 ();
 sg13g2_decap_8 FILLER_19_1390 ();
 sg13g2_decap_8 FILLER_19_1397 ();
 sg13g2_decap_8 FILLER_19_1404 ();
 sg13g2_decap_8 FILLER_19_1411 ();
 sg13g2_decap_8 FILLER_19_1418 ();
 sg13g2_decap_8 FILLER_19_1425 ();
 sg13g2_decap_8 FILLER_19_1432 ();
 sg13g2_decap_8 FILLER_19_1439 ();
 sg13g2_decap_8 FILLER_19_1446 ();
 sg13g2_decap_8 FILLER_19_1453 ();
 sg13g2_decap_8 FILLER_19_1460 ();
 sg13g2_decap_8 FILLER_19_1467 ();
 sg13g2_decap_8 FILLER_19_1474 ();
 sg13g2_decap_8 FILLER_19_1481 ();
 sg13g2_decap_8 FILLER_19_1488 ();
 sg13g2_decap_8 FILLER_19_1495 ();
 sg13g2_decap_8 FILLER_19_1502 ();
 sg13g2_decap_8 FILLER_19_1509 ();
 sg13g2_decap_8 FILLER_19_1516 ();
 sg13g2_decap_8 FILLER_19_1523 ();
 sg13g2_decap_8 FILLER_19_1530 ();
 sg13g2_decap_8 FILLER_19_1537 ();
 sg13g2_decap_8 FILLER_19_1544 ();
 sg13g2_decap_8 FILLER_19_1551 ();
 sg13g2_decap_8 FILLER_19_1558 ();
 sg13g2_decap_8 FILLER_19_1565 ();
 sg13g2_decap_8 FILLER_19_1572 ();
 sg13g2_decap_8 FILLER_19_1579 ();
 sg13g2_decap_8 FILLER_19_1586 ();
 sg13g2_decap_8 FILLER_19_1593 ();
 sg13g2_decap_8 FILLER_19_1600 ();
 sg13g2_decap_8 FILLER_19_1607 ();
 sg13g2_decap_8 FILLER_19_1614 ();
 sg13g2_decap_8 FILLER_19_1621 ();
 sg13g2_decap_8 FILLER_19_1628 ();
 sg13g2_decap_8 FILLER_19_1635 ();
 sg13g2_decap_8 FILLER_19_1642 ();
 sg13g2_decap_8 FILLER_19_1649 ();
 sg13g2_decap_8 FILLER_19_1656 ();
 sg13g2_decap_8 FILLER_19_1663 ();
 sg13g2_decap_8 FILLER_19_1670 ();
 sg13g2_decap_8 FILLER_19_1677 ();
 sg13g2_decap_8 FILLER_19_1684 ();
 sg13g2_decap_8 FILLER_19_1691 ();
 sg13g2_decap_8 FILLER_19_1698 ();
 sg13g2_decap_8 FILLER_19_1705 ();
 sg13g2_decap_8 FILLER_19_1712 ();
 sg13g2_decap_8 FILLER_19_1719 ();
 sg13g2_decap_8 FILLER_19_1726 ();
 sg13g2_decap_8 FILLER_19_1733 ();
 sg13g2_decap_8 FILLER_19_1740 ();
 sg13g2_decap_8 FILLER_19_1747 ();
 sg13g2_decap_8 FILLER_19_1754 ();
 sg13g2_decap_8 FILLER_19_1761 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_fill_1 FILLER_20_95 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_decap_8 FILLER_20_139 ();
 sg13g2_fill_2 FILLER_20_156 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_fill_2 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_197 ();
 sg13g2_fill_2 FILLER_20_204 ();
 sg13g2_fill_1 FILLER_20_215 ();
 sg13g2_decap_4 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_254 ();
 sg13g2_fill_2 FILLER_20_273 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_306 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_fill_2 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_387 ();
 sg13g2_decap_4 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_20_410 ();
 sg13g2_fill_2 FILLER_20_417 ();
 sg13g2_decap_4 FILLER_20_423 ();
 sg13g2_fill_2 FILLER_20_441 ();
 sg13g2_fill_1 FILLER_20_443 ();
 sg13g2_fill_2 FILLER_20_450 ();
 sg13g2_fill_1 FILLER_20_457 ();
 sg13g2_fill_2 FILLER_20_472 ();
 sg13g2_fill_1 FILLER_20_474 ();
 sg13g2_fill_1 FILLER_20_481 ();
 sg13g2_fill_1 FILLER_20_485 ();
 sg13g2_fill_2 FILLER_20_507 ();
 sg13g2_fill_1 FILLER_20_515 ();
 sg13g2_fill_2 FILLER_20_533 ();
 sg13g2_decap_8 FILLER_20_540 ();
 sg13g2_decap_4 FILLER_20_547 ();
 sg13g2_fill_2 FILLER_20_577 ();
 sg13g2_fill_2 FILLER_20_597 ();
 sg13g2_fill_1 FILLER_20_599 ();
 sg13g2_decap_8 FILLER_20_612 ();
 sg13g2_fill_2 FILLER_20_633 ();
 sg13g2_fill_1 FILLER_20_635 ();
 sg13g2_fill_2 FILLER_20_645 ();
 sg13g2_fill_2 FILLER_20_652 ();
 sg13g2_decap_8 FILLER_20_668 ();
 sg13g2_fill_2 FILLER_20_675 ();
 sg13g2_fill_1 FILLER_20_677 ();
 sg13g2_fill_1 FILLER_20_695 ();
 sg13g2_fill_1 FILLER_20_713 ();
 sg13g2_decap_8 FILLER_20_718 ();
 sg13g2_fill_2 FILLER_20_725 ();
 sg13g2_fill_1 FILLER_20_727 ();
 sg13g2_decap_4 FILLER_20_748 ();
 sg13g2_fill_2 FILLER_20_752 ();
 sg13g2_decap_8 FILLER_20_768 ();
 sg13g2_decap_8 FILLER_20_775 ();
 sg13g2_decap_4 FILLER_20_782 ();
 sg13g2_fill_1 FILLER_20_786 ();
 sg13g2_decap_4 FILLER_20_800 ();
 sg13g2_fill_1 FILLER_20_804 ();
 sg13g2_decap_4 FILLER_20_832 ();
 sg13g2_fill_2 FILLER_20_836 ();
 sg13g2_decap_8 FILLER_20_856 ();
 sg13g2_fill_1 FILLER_20_863 ();
 sg13g2_decap_8 FILLER_20_903 ();
 sg13g2_fill_2 FILLER_20_913 ();
 sg13g2_decap_4 FILLER_20_925 ();
 sg13g2_fill_2 FILLER_20_949 ();
 sg13g2_fill_1 FILLER_20_951 ();
 sg13g2_fill_1 FILLER_20_961 ();
 sg13g2_fill_1 FILLER_20_966 ();
 sg13g2_decap_4 FILLER_20_977 ();
 sg13g2_decap_4 FILLER_20_1018 ();
 sg13g2_fill_1 FILLER_20_1022 ();
 sg13g2_decap_8 FILLER_20_1033 ();
 sg13g2_fill_2 FILLER_20_1040 ();
 sg13g2_decap_8 FILLER_20_1072 ();
 sg13g2_decap_8 FILLER_20_1112 ();
 sg13g2_decap_8 FILLER_20_1119 ();
 sg13g2_decap_8 FILLER_20_1126 ();
 sg13g2_decap_8 FILLER_20_1133 ();
 sg13g2_decap_8 FILLER_20_1140 ();
 sg13g2_decap_8 FILLER_20_1147 ();
 sg13g2_decap_8 FILLER_20_1154 ();
 sg13g2_decap_8 FILLER_20_1161 ();
 sg13g2_decap_8 FILLER_20_1168 ();
 sg13g2_decap_8 FILLER_20_1175 ();
 sg13g2_decap_8 FILLER_20_1182 ();
 sg13g2_decap_8 FILLER_20_1189 ();
 sg13g2_decap_8 FILLER_20_1196 ();
 sg13g2_decap_8 FILLER_20_1203 ();
 sg13g2_decap_8 FILLER_20_1210 ();
 sg13g2_decap_8 FILLER_20_1217 ();
 sg13g2_decap_8 FILLER_20_1224 ();
 sg13g2_decap_8 FILLER_20_1231 ();
 sg13g2_decap_8 FILLER_20_1238 ();
 sg13g2_decap_8 FILLER_20_1245 ();
 sg13g2_decap_8 FILLER_20_1252 ();
 sg13g2_decap_8 FILLER_20_1259 ();
 sg13g2_decap_8 FILLER_20_1266 ();
 sg13g2_decap_8 FILLER_20_1273 ();
 sg13g2_decap_8 FILLER_20_1280 ();
 sg13g2_decap_8 FILLER_20_1287 ();
 sg13g2_decap_8 FILLER_20_1294 ();
 sg13g2_decap_8 FILLER_20_1301 ();
 sg13g2_decap_8 FILLER_20_1308 ();
 sg13g2_decap_8 FILLER_20_1315 ();
 sg13g2_decap_8 FILLER_20_1322 ();
 sg13g2_decap_8 FILLER_20_1329 ();
 sg13g2_decap_8 FILLER_20_1336 ();
 sg13g2_decap_8 FILLER_20_1343 ();
 sg13g2_decap_8 FILLER_20_1350 ();
 sg13g2_decap_8 FILLER_20_1357 ();
 sg13g2_decap_8 FILLER_20_1364 ();
 sg13g2_decap_8 FILLER_20_1371 ();
 sg13g2_decap_8 FILLER_20_1378 ();
 sg13g2_decap_8 FILLER_20_1385 ();
 sg13g2_decap_8 FILLER_20_1392 ();
 sg13g2_decap_8 FILLER_20_1399 ();
 sg13g2_decap_8 FILLER_20_1406 ();
 sg13g2_decap_8 FILLER_20_1413 ();
 sg13g2_decap_8 FILLER_20_1420 ();
 sg13g2_decap_8 FILLER_20_1427 ();
 sg13g2_decap_8 FILLER_20_1434 ();
 sg13g2_decap_8 FILLER_20_1441 ();
 sg13g2_decap_8 FILLER_20_1448 ();
 sg13g2_decap_8 FILLER_20_1455 ();
 sg13g2_decap_8 FILLER_20_1462 ();
 sg13g2_decap_8 FILLER_20_1469 ();
 sg13g2_decap_8 FILLER_20_1476 ();
 sg13g2_decap_8 FILLER_20_1483 ();
 sg13g2_decap_8 FILLER_20_1490 ();
 sg13g2_decap_8 FILLER_20_1497 ();
 sg13g2_decap_8 FILLER_20_1504 ();
 sg13g2_decap_8 FILLER_20_1511 ();
 sg13g2_decap_8 FILLER_20_1518 ();
 sg13g2_decap_8 FILLER_20_1525 ();
 sg13g2_decap_8 FILLER_20_1532 ();
 sg13g2_decap_8 FILLER_20_1539 ();
 sg13g2_decap_8 FILLER_20_1546 ();
 sg13g2_decap_8 FILLER_20_1553 ();
 sg13g2_decap_8 FILLER_20_1560 ();
 sg13g2_decap_8 FILLER_20_1567 ();
 sg13g2_decap_8 FILLER_20_1574 ();
 sg13g2_decap_8 FILLER_20_1581 ();
 sg13g2_decap_8 FILLER_20_1588 ();
 sg13g2_decap_8 FILLER_20_1595 ();
 sg13g2_decap_8 FILLER_20_1602 ();
 sg13g2_decap_8 FILLER_20_1609 ();
 sg13g2_decap_8 FILLER_20_1616 ();
 sg13g2_decap_8 FILLER_20_1623 ();
 sg13g2_decap_8 FILLER_20_1630 ();
 sg13g2_decap_8 FILLER_20_1637 ();
 sg13g2_decap_8 FILLER_20_1644 ();
 sg13g2_decap_8 FILLER_20_1651 ();
 sg13g2_decap_8 FILLER_20_1658 ();
 sg13g2_decap_8 FILLER_20_1665 ();
 sg13g2_decap_8 FILLER_20_1672 ();
 sg13g2_decap_8 FILLER_20_1679 ();
 sg13g2_decap_8 FILLER_20_1686 ();
 sg13g2_decap_8 FILLER_20_1693 ();
 sg13g2_decap_8 FILLER_20_1700 ();
 sg13g2_decap_8 FILLER_20_1707 ();
 sg13g2_decap_8 FILLER_20_1714 ();
 sg13g2_decap_8 FILLER_20_1721 ();
 sg13g2_decap_8 FILLER_20_1728 ();
 sg13g2_decap_8 FILLER_20_1735 ();
 sg13g2_decap_8 FILLER_20_1742 ();
 sg13g2_decap_8 FILLER_20_1749 ();
 sg13g2_decap_8 FILLER_20_1756 ();
 sg13g2_decap_4 FILLER_20_1763 ();
 sg13g2_fill_1 FILLER_20_1767 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_21 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_decap_4 FILLER_21_106 ();
 sg13g2_fill_1 FILLER_21_115 ();
 sg13g2_fill_1 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_190 ();
 sg13g2_fill_2 FILLER_21_210 ();
 sg13g2_fill_1 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_311 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_4 FILLER_21_357 ();
 sg13g2_decap_4 FILLER_21_366 ();
 sg13g2_decap_4 FILLER_21_382 ();
 sg13g2_fill_2 FILLER_21_386 ();
 sg13g2_fill_2 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_412 ();
 sg13g2_fill_1 FILLER_21_418 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_fill_2 FILLER_21_451 ();
 sg13g2_decap_4 FILLER_21_469 ();
 sg13g2_fill_1 FILLER_21_473 ();
 sg13g2_fill_1 FILLER_21_488 ();
 sg13g2_fill_1 FILLER_21_510 ();
 sg13g2_fill_1 FILLER_21_521 ();
 sg13g2_fill_1 FILLER_21_544 ();
 sg13g2_decap_8 FILLER_21_565 ();
 sg13g2_fill_1 FILLER_21_572 ();
 sg13g2_fill_2 FILLER_21_589 ();
 sg13g2_fill_2 FILLER_21_600 ();
 sg13g2_fill_2 FILLER_21_657 ();
 sg13g2_fill_1 FILLER_21_659 ();
 sg13g2_fill_2 FILLER_21_669 ();
 sg13g2_fill_1 FILLER_21_686 ();
 sg13g2_fill_1 FILLER_21_691 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_fill_2 FILLER_21_707 ();
 sg13g2_fill_1 FILLER_21_709 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_fill_2 FILLER_21_756 ();
 sg13g2_fill_1 FILLER_21_758 ();
 sg13g2_fill_1 FILLER_21_769 ();
 sg13g2_decap_4 FILLER_21_805 ();
 sg13g2_fill_1 FILLER_21_809 ();
 sg13g2_decap_4 FILLER_21_831 ();
 sg13g2_fill_2 FILLER_21_835 ();
 sg13g2_fill_1 FILLER_21_860 ();
 sg13g2_decap_8 FILLER_21_875 ();
 sg13g2_decap_8 FILLER_21_882 ();
 sg13g2_fill_1 FILLER_21_889 ();
 sg13g2_decap_8 FILLER_21_898 ();
 sg13g2_decap_4 FILLER_21_905 ();
 sg13g2_fill_2 FILLER_21_909 ();
 sg13g2_fill_1 FILLER_21_920 ();
 sg13g2_decap_4 FILLER_21_926 ();
 sg13g2_decap_8 FILLER_21_951 ();
 sg13g2_fill_2 FILLER_21_972 ();
 sg13g2_fill_1 FILLER_21_982 ();
 sg13g2_decap_4 FILLER_21_993 ();
 sg13g2_fill_1 FILLER_21_997 ();
 sg13g2_fill_2 FILLER_21_1008 ();
 sg13g2_fill_2 FILLER_21_1018 ();
 sg13g2_decap_4 FILLER_21_1034 ();
 sg13g2_decap_8 FILLER_21_1052 ();
 sg13g2_fill_1 FILLER_21_1075 ();
 sg13g2_decap_8 FILLER_21_1104 ();
 sg13g2_decap_8 FILLER_21_1111 ();
 sg13g2_decap_8 FILLER_21_1118 ();
 sg13g2_decap_8 FILLER_21_1125 ();
 sg13g2_decap_8 FILLER_21_1132 ();
 sg13g2_decap_8 FILLER_21_1139 ();
 sg13g2_decap_8 FILLER_21_1146 ();
 sg13g2_decap_8 FILLER_21_1153 ();
 sg13g2_decap_8 FILLER_21_1160 ();
 sg13g2_decap_8 FILLER_21_1167 ();
 sg13g2_decap_8 FILLER_21_1174 ();
 sg13g2_decap_8 FILLER_21_1181 ();
 sg13g2_decap_8 FILLER_21_1188 ();
 sg13g2_decap_8 FILLER_21_1195 ();
 sg13g2_decap_8 FILLER_21_1202 ();
 sg13g2_decap_8 FILLER_21_1209 ();
 sg13g2_decap_8 FILLER_21_1216 ();
 sg13g2_decap_8 FILLER_21_1223 ();
 sg13g2_decap_8 FILLER_21_1230 ();
 sg13g2_decap_8 FILLER_21_1237 ();
 sg13g2_decap_8 FILLER_21_1244 ();
 sg13g2_decap_8 FILLER_21_1251 ();
 sg13g2_decap_8 FILLER_21_1258 ();
 sg13g2_decap_8 FILLER_21_1265 ();
 sg13g2_decap_8 FILLER_21_1272 ();
 sg13g2_decap_8 FILLER_21_1279 ();
 sg13g2_decap_8 FILLER_21_1286 ();
 sg13g2_decap_8 FILLER_21_1293 ();
 sg13g2_decap_8 FILLER_21_1300 ();
 sg13g2_decap_8 FILLER_21_1307 ();
 sg13g2_decap_8 FILLER_21_1314 ();
 sg13g2_decap_8 FILLER_21_1321 ();
 sg13g2_decap_8 FILLER_21_1328 ();
 sg13g2_decap_8 FILLER_21_1335 ();
 sg13g2_decap_8 FILLER_21_1342 ();
 sg13g2_decap_8 FILLER_21_1349 ();
 sg13g2_decap_8 FILLER_21_1356 ();
 sg13g2_decap_8 FILLER_21_1363 ();
 sg13g2_decap_8 FILLER_21_1370 ();
 sg13g2_decap_8 FILLER_21_1377 ();
 sg13g2_decap_8 FILLER_21_1384 ();
 sg13g2_decap_8 FILLER_21_1391 ();
 sg13g2_decap_8 FILLER_21_1398 ();
 sg13g2_decap_8 FILLER_21_1405 ();
 sg13g2_decap_8 FILLER_21_1412 ();
 sg13g2_decap_8 FILLER_21_1419 ();
 sg13g2_decap_8 FILLER_21_1426 ();
 sg13g2_decap_8 FILLER_21_1433 ();
 sg13g2_decap_8 FILLER_21_1440 ();
 sg13g2_decap_8 FILLER_21_1447 ();
 sg13g2_decap_8 FILLER_21_1454 ();
 sg13g2_decap_8 FILLER_21_1461 ();
 sg13g2_decap_8 FILLER_21_1468 ();
 sg13g2_decap_8 FILLER_21_1475 ();
 sg13g2_decap_8 FILLER_21_1482 ();
 sg13g2_decap_8 FILLER_21_1489 ();
 sg13g2_decap_8 FILLER_21_1496 ();
 sg13g2_decap_8 FILLER_21_1503 ();
 sg13g2_decap_8 FILLER_21_1510 ();
 sg13g2_decap_8 FILLER_21_1517 ();
 sg13g2_decap_8 FILLER_21_1524 ();
 sg13g2_decap_8 FILLER_21_1531 ();
 sg13g2_decap_8 FILLER_21_1538 ();
 sg13g2_decap_8 FILLER_21_1545 ();
 sg13g2_decap_8 FILLER_21_1552 ();
 sg13g2_decap_8 FILLER_21_1559 ();
 sg13g2_decap_8 FILLER_21_1566 ();
 sg13g2_decap_8 FILLER_21_1573 ();
 sg13g2_decap_8 FILLER_21_1580 ();
 sg13g2_decap_8 FILLER_21_1587 ();
 sg13g2_decap_8 FILLER_21_1594 ();
 sg13g2_decap_8 FILLER_21_1601 ();
 sg13g2_decap_8 FILLER_21_1608 ();
 sg13g2_decap_8 FILLER_21_1615 ();
 sg13g2_decap_8 FILLER_21_1622 ();
 sg13g2_decap_8 FILLER_21_1629 ();
 sg13g2_decap_8 FILLER_21_1636 ();
 sg13g2_decap_8 FILLER_21_1643 ();
 sg13g2_decap_8 FILLER_21_1650 ();
 sg13g2_decap_8 FILLER_21_1657 ();
 sg13g2_decap_8 FILLER_21_1664 ();
 sg13g2_decap_8 FILLER_21_1671 ();
 sg13g2_decap_8 FILLER_21_1678 ();
 sg13g2_decap_8 FILLER_21_1685 ();
 sg13g2_decap_8 FILLER_21_1692 ();
 sg13g2_decap_8 FILLER_21_1699 ();
 sg13g2_decap_8 FILLER_21_1706 ();
 sg13g2_decap_8 FILLER_21_1713 ();
 sg13g2_decap_8 FILLER_21_1720 ();
 sg13g2_decap_8 FILLER_21_1727 ();
 sg13g2_decap_8 FILLER_21_1734 ();
 sg13g2_decap_8 FILLER_21_1741 ();
 sg13g2_decap_8 FILLER_21_1748 ();
 sg13g2_decap_8 FILLER_21_1755 ();
 sg13g2_decap_4 FILLER_21_1762 ();
 sg13g2_fill_2 FILLER_21_1766 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_95 ();
 sg13g2_fill_1 FILLER_22_99 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_fill_2 FILLER_22_213 ();
 sg13g2_fill_1 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_255 ();
 sg13g2_fill_1 FILLER_22_281 ();
 sg13g2_fill_1 FILLER_22_303 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_fill_2 FILLER_22_331 ();
 sg13g2_fill_1 FILLER_22_333 ();
 sg13g2_fill_1 FILLER_22_360 ();
 sg13g2_fill_2 FILLER_22_387 ();
 sg13g2_fill_1 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_fill_1 FILLER_22_409 ();
 sg13g2_decap_8 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_22_435 ();
 sg13g2_fill_1 FILLER_22_447 ();
 sg13g2_fill_2 FILLER_22_465 ();
 sg13g2_fill_1 FILLER_22_467 ();
 sg13g2_fill_1 FILLER_22_484 ();
 sg13g2_decap_4 FILLER_22_513 ();
 sg13g2_fill_1 FILLER_22_530 ();
 sg13g2_decap_8 FILLER_22_543 ();
 sg13g2_fill_2 FILLER_22_550 ();
 sg13g2_fill_1 FILLER_22_552 ();
 sg13g2_decap_4 FILLER_22_573 ();
 sg13g2_fill_1 FILLER_22_577 ();
 sg13g2_decap_4 FILLER_22_583 ();
 sg13g2_fill_2 FILLER_22_587 ();
 sg13g2_fill_1 FILLER_22_593 ();
 sg13g2_decap_4 FILLER_22_602 ();
 sg13g2_fill_2 FILLER_22_606 ();
 sg13g2_decap_8 FILLER_22_622 ();
 sg13g2_decap_8 FILLER_22_629 ();
 sg13g2_fill_2 FILLER_22_636 ();
 sg13g2_fill_2 FILLER_22_642 ();
 sg13g2_fill_2 FILLER_22_676 ();
 sg13g2_fill_1 FILLER_22_678 ();
 sg13g2_fill_2 FILLER_22_711 ();
 sg13g2_fill_2 FILLER_22_730 ();
 sg13g2_fill_1 FILLER_22_732 ();
 sg13g2_fill_2 FILLER_22_745 ();
 sg13g2_fill_2 FILLER_22_761 ();
 sg13g2_decap_8 FILLER_22_781 ();
 sg13g2_decap_4 FILLER_22_788 ();
 sg13g2_fill_2 FILLER_22_792 ();
 sg13g2_decap_8 FILLER_22_803 ();
 sg13g2_decap_8 FILLER_22_836 ();
 sg13g2_fill_2 FILLER_22_852 ();
 sg13g2_fill_1 FILLER_22_854 ();
 sg13g2_fill_1 FILLER_22_868 ();
 sg13g2_fill_2 FILLER_22_881 ();
 sg13g2_fill_1 FILLER_22_888 ();
 sg13g2_fill_2 FILLER_22_938 ();
 sg13g2_decap_8 FILLER_22_950 ();
 sg13g2_fill_2 FILLER_22_994 ();
 sg13g2_fill_2 FILLER_22_1008 ();
 sg13g2_fill_1 FILLER_22_1010 ();
 sg13g2_decap_8 FILLER_22_1025 ();
 sg13g2_fill_2 FILLER_22_1032 ();
 sg13g2_fill_1 FILLER_22_1034 ();
 sg13g2_decap_8 FILLER_22_1110 ();
 sg13g2_decap_8 FILLER_22_1117 ();
 sg13g2_decap_8 FILLER_22_1124 ();
 sg13g2_decap_8 FILLER_22_1131 ();
 sg13g2_decap_8 FILLER_22_1138 ();
 sg13g2_decap_8 FILLER_22_1145 ();
 sg13g2_decap_8 FILLER_22_1152 ();
 sg13g2_decap_8 FILLER_22_1159 ();
 sg13g2_decap_8 FILLER_22_1166 ();
 sg13g2_decap_8 FILLER_22_1173 ();
 sg13g2_decap_8 FILLER_22_1180 ();
 sg13g2_decap_8 FILLER_22_1187 ();
 sg13g2_decap_8 FILLER_22_1194 ();
 sg13g2_decap_8 FILLER_22_1201 ();
 sg13g2_decap_8 FILLER_22_1208 ();
 sg13g2_decap_8 FILLER_22_1215 ();
 sg13g2_decap_8 FILLER_22_1222 ();
 sg13g2_decap_8 FILLER_22_1229 ();
 sg13g2_decap_8 FILLER_22_1236 ();
 sg13g2_decap_8 FILLER_22_1243 ();
 sg13g2_decap_8 FILLER_22_1250 ();
 sg13g2_decap_8 FILLER_22_1257 ();
 sg13g2_decap_8 FILLER_22_1264 ();
 sg13g2_decap_8 FILLER_22_1271 ();
 sg13g2_decap_8 FILLER_22_1278 ();
 sg13g2_decap_8 FILLER_22_1285 ();
 sg13g2_decap_8 FILLER_22_1292 ();
 sg13g2_decap_8 FILLER_22_1299 ();
 sg13g2_decap_8 FILLER_22_1306 ();
 sg13g2_decap_8 FILLER_22_1313 ();
 sg13g2_decap_8 FILLER_22_1320 ();
 sg13g2_decap_8 FILLER_22_1327 ();
 sg13g2_decap_8 FILLER_22_1334 ();
 sg13g2_decap_8 FILLER_22_1341 ();
 sg13g2_decap_8 FILLER_22_1348 ();
 sg13g2_decap_8 FILLER_22_1355 ();
 sg13g2_decap_8 FILLER_22_1362 ();
 sg13g2_decap_8 FILLER_22_1369 ();
 sg13g2_decap_8 FILLER_22_1376 ();
 sg13g2_decap_8 FILLER_22_1383 ();
 sg13g2_decap_8 FILLER_22_1390 ();
 sg13g2_decap_8 FILLER_22_1397 ();
 sg13g2_decap_8 FILLER_22_1404 ();
 sg13g2_decap_8 FILLER_22_1411 ();
 sg13g2_decap_8 FILLER_22_1418 ();
 sg13g2_decap_8 FILLER_22_1425 ();
 sg13g2_decap_8 FILLER_22_1432 ();
 sg13g2_decap_8 FILLER_22_1439 ();
 sg13g2_decap_8 FILLER_22_1446 ();
 sg13g2_decap_8 FILLER_22_1453 ();
 sg13g2_decap_8 FILLER_22_1460 ();
 sg13g2_decap_8 FILLER_22_1467 ();
 sg13g2_decap_8 FILLER_22_1474 ();
 sg13g2_decap_8 FILLER_22_1481 ();
 sg13g2_decap_8 FILLER_22_1488 ();
 sg13g2_decap_8 FILLER_22_1495 ();
 sg13g2_decap_8 FILLER_22_1502 ();
 sg13g2_decap_8 FILLER_22_1509 ();
 sg13g2_decap_8 FILLER_22_1516 ();
 sg13g2_decap_8 FILLER_22_1523 ();
 sg13g2_decap_8 FILLER_22_1530 ();
 sg13g2_decap_8 FILLER_22_1537 ();
 sg13g2_decap_8 FILLER_22_1544 ();
 sg13g2_decap_8 FILLER_22_1551 ();
 sg13g2_decap_8 FILLER_22_1558 ();
 sg13g2_decap_8 FILLER_22_1565 ();
 sg13g2_decap_8 FILLER_22_1572 ();
 sg13g2_decap_8 FILLER_22_1579 ();
 sg13g2_decap_8 FILLER_22_1586 ();
 sg13g2_decap_8 FILLER_22_1593 ();
 sg13g2_decap_8 FILLER_22_1600 ();
 sg13g2_decap_8 FILLER_22_1607 ();
 sg13g2_decap_8 FILLER_22_1614 ();
 sg13g2_decap_8 FILLER_22_1621 ();
 sg13g2_decap_8 FILLER_22_1628 ();
 sg13g2_decap_8 FILLER_22_1635 ();
 sg13g2_decap_8 FILLER_22_1642 ();
 sg13g2_decap_8 FILLER_22_1649 ();
 sg13g2_decap_8 FILLER_22_1656 ();
 sg13g2_decap_8 FILLER_22_1663 ();
 sg13g2_decap_8 FILLER_22_1670 ();
 sg13g2_decap_8 FILLER_22_1677 ();
 sg13g2_decap_8 FILLER_22_1684 ();
 sg13g2_decap_8 FILLER_22_1691 ();
 sg13g2_decap_8 FILLER_22_1698 ();
 sg13g2_decap_8 FILLER_22_1705 ();
 sg13g2_decap_8 FILLER_22_1712 ();
 sg13g2_decap_8 FILLER_22_1719 ();
 sg13g2_decap_8 FILLER_22_1726 ();
 sg13g2_decap_8 FILLER_22_1733 ();
 sg13g2_decap_8 FILLER_22_1740 ();
 sg13g2_decap_8 FILLER_22_1747 ();
 sg13g2_decap_8 FILLER_22_1754 ();
 sg13g2_decap_8 FILLER_22_1761 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_78 ();
 sg13g2_fill_2 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_111 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_169 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_decap_4 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_339 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_fill_2 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_442 ();
 sg13g2_decap_8 FILLER_23_449 ();
 sg13g2_fill_1 FILLER_23_488 ();
 sg13g2_decap_4 FILLER_23_499 ();
 sg13g2_fill_1 FILLER_23_503 ();
 sg13g2_decap_4 FILLER_23_510 ();
 sg13g2_fill_1 FILLER_23_524 ();
 sg13g2_fill_1 FILLER_23_589 ();
 sg13g2_decap_4 FILLER_23_623 ();
 sg13g2_fill_2 FILLER_23_635 ();
 sg13g2_fill_1 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_643 ();
 sg13g2_decap_8 FILLER_23_650 ();
 sg13g2_fill_2 FILLER_23_657 ();
 sg13g2_fill_1 FILLER_23_659 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_4 FILLER_23_679 ();
 sg13g2_fill_1 FILLER_23_683 ();
 sg13g2_fill_1 FILLER_23_694 ();
 sg13g2_fill_2 FILLER_23_705 ();
 sg13g2_fill_1 FILLER_23_734 ();
 sg13g2_fill_2 FILLER_23_740 ();
 sg13g2_fill_1 FILLER_23_742 ();
 sg13g2_fill_2 FILLER_23_758 ();
 sg13g2_fill_1 FILLER_23_760 ();
 sg13g2_fill_1 FILLER_23_767 ();
 sg13g2_decap_4 FILLER_23_807 ();
 sg13g2_decap_8 FILLER_23_830 ();
 sg13g2_decap_8 FILLER_23_837 ();
 sg13g2_fill_1 FILLER_23_844 ();
 sg13g2_fill_2 FILLER_23_861 ();
 sg13g2_fill_2 FILLER_23_872 ();
 sg13g2_decap_8 FILLER_23_896 ();
 sg13g2_fill_2 FILLER_23_903 ();
 sg13g2_fill_1 FILLER_23_905 ();
 sg13g2_fill_2 FILLER_23_920 ();
 sg13g2_decap_4 FILLER_23_946 ();
 sg13g2_decap_4 FILLER_23_954 ();
 sg13g2_fill_2 FILLER_23_958 ();
 sg13g2_decap_4 FILLER_23_971 ();
 sg13g2_fill_1 FILLER_23_975 ();
 sg13g2_decap_4 FILLER_23_981 ();
 sg13g2_decap_8 FILLER_23_989 ();
 sg13g2_decap_4 FILLER_23_996 ();
 sg13g2_fill_1 FILLER_23_1008 ();
 sg13g2_fill_2 FILLER_23_1022 ();
 sg13g2_fill_1 FILLER_23_1028 ();
 sg13g2_decap_8 FILLER_23_1054 ();
 sg13g2_decap_4 FILLER_23_1061 ();
 sg13g2_decap_4 FILLER_23_1075 ();
 sg13g2_fill_2 FILLER_23_1079 ();
 sg13g2_decap_4 FILLER_23_1100 ();
 sg13g2_fill_1 FILLER_23_1104 ();
 sg13g2_decap_8 FILLER_23_1114 ();
 sg13g2_decap_8 FILLER_23_1121 ();
 sg13g2_decap_8 FILLER_23_1128 ();
 sg13g2_decap_8 FILLER_23_1135 ();
 sg13g2_decap_8 FILLER_23_1142 ();
 sg13g2_decap_8 FILLER_23_1149 ();
 sg13g2_decap_8 FILLER_23_1156 ();
 sg13g2_decap_8 FILLER_23_1163 ();
 sg13g2_decap_8 FILLER_23_1170 ();
 sg13g2_decap_8 FILLER_23_1177 ();
 sg13g2_decap_8 FILLER_23_1184 ();
 sg13g2_decap_8 FILLER_23_1191 ();
 sg13g2_decap_8 FILLER_23_1198 ();
 sg13g2_decap_8 FILLER_23_1205 ();
 sg13g2_decap_8 FILLER_23_1212 ();
 sg13g2_decap_8 FILLER_23_1219 ();
 sg13g2_decap_8 FILLER_23_1226 ();
 sg13g2_decap_8 FILLER_23_1233 ();
 sg13g2_decap_8 FILLER_23_1240 ();
 sg13g2_decap_8 FILLER_23_1247 ();
 sg13g2_decap_8 FILLER_23_1254 ();
 sg13g2_decap_8 FILLER_23_1261 ();
 sg13g2_decap_8 FILLER_23_1268 ();
 sg13g2_decap_8 FILLER_23_1275 ();
 sg13g2_decap_8 FILLER_23_1282 ();
 sg13g2_decap_8 FILLER_23_1289 ();
 sg13g2_decap_8 FILLER_23_1296 ();
 sg13g2_decap_8 FILLER_23_1303 ();
 sg13g2_decap_8 FILLER_23_1310 ();
 sg13g2_decap_8 FILLER_23_1317 ();
 sg13g2_decap_8 FILLER_23_1324 ();
 sg13g2_decap_8 FILLER_23_1331 ();
 sg13g2_decap_8 FILLER_23_1338 ();
 sg13g2_decap_8 FILLER_23_1345 ();
 sg13g2_decap_8 FILLER_23_1352 ();
 sg13g2_decap_8 FILLER_23_1359 ();
 sg13g2_decap_8 FILLER_23_1366 ();
 sg13g2_decap_8 FILLER_23_1373 ();
 sg13g2_decap_8 FILLER_23_1380 ();
 sg13g2_decap_8 FILLER_23_1387 ();
 sg13g2_decap_8 FILLER_23_1394 ();
 sg13g2_decap_8 FILLER_23_1401 ();
 sg13g2_decap_8 FILLER_23_1408 ();
 sg13g2_decap_8 FILLER_23_1415 ();
 sg13g2_decap_8 FILLER_23_1422 ();
 sg13g2_decap_8 FILLER_23_1429 ();
 sg13g2_decap_8 FILLER_23_1436 ();
 sg13g2_decap_8 FILLER_23_1443 ();
 sg13g2_decap_8 FILLER_23_1450 ();
 sg13g2_decap_8 FILLER_23_1457 ();
 sg13g2_decap_8 FILLER_23_1464 ();
 sg13g2_decap_8 FILLER_23_1471 ();
 sg13g2_decap_8 FILLER_23_1478 ();
 sg13g2_decap_8 FILLER_23_1485 ();
 sg13g2_decap_8 FILLER_23_1492 ();
 sg13g2_decap_8 FILLER_23_1499 ();
 sg13g2_decap_8 FILLER_23_1506 ();
 sg13g2_decap_8 FILLER_23_1513 ();
 sg13g2_decap_8 FILLER_23_1520 ();
 sg13g2_decap_8 FILLER_23_1527 ();
 sg13g2_decap_8 FILLER_23_1534 ();
 sg13g2_decap_8 FILLER_23_1541 ();
 sg13g2_decap_8 FILLER_23_1548 ();
 sg13g2_decap_8 FILLER_23_1555 ();
 sg13g2_decap_8 FILLER_23_1562 ();
 sg13g2_decap_8 FILLER_23_1569 ();
 sg13g2_decap_8 FILLER_23_1576 ();
 sg13g2_decap_8 FILLER_23_1583 ();
 sg13g2_decap_8 FILLER_23_1590 ();
 sg13g2_decap_8 FILLER_23_1597 ();
 sg13g2_decap_8 FILLER_23_1604 ();
 sg13g2_decap_8 FILLER_23_1611 ();
 sg13g2_decap_8 FILLER_23_1618 ();
 sg13g2_decap_8 FILLER_23_1625 ();
 sg13g2_decap_8 FILLER_23_1632 ();
 sg13g2_decap_8 FILLER_23_1639 ();
 sg13g2_decap_8 FILLER_23_1646 ();
 sg13g2_decap_8 FILLER_23_1653 ();
 sg13g2_decap_8 FILLER_23_1660 ();
 sg13g2_decap_8 FILLER_23_1667 ();
 sg13g2_decap_8 FILLER_23_1674 ();
 sg13g2_decap_8 FILLER_23_1681 ();
 sg13g2_decap_8 FILLER_23_1688 ();
 sg13g2_decap_8 FILLER_23_1695 ();
 sg13g2_decap_8 FILLER_23_1702 ();
 sg13g2_decap_8 FILLER_23_1709 ();
 sg13g2_decap_8 FILLER_23_1716 ();
 sg13g2_decap_8 FILLER_23_1723 ();
 sg13g2_decap_8 FILLER_23_1730 ();
 sg13g2_decap_8 FILLER_23_1737 ();
 sg13g2_decap_8 FILLER_23_1744 ();
 sg13g2_decap_8 FILLER_23_1751 ();
 sg13g2_decap_8 FILLER_23_1758 ();
 sg13g2_fill_2 FILLER_23_1765 ();
 sg13g2_fill_1 FILLER_23_1767 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_44 ();
 sg13g2_fill_1 FILLER_24_80 ();
 sg13g2_fill_1 FILLER_24_107 ();
 sg13g2_fill_2 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_decap_4 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_144 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_216 ();
 sg13g2_fill_1 FILLER_24_244 ();
 sg13g2_decap_4 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_319 ();
 sg13g2_fill_2 FILLER_24_332 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_fill_2 FILLER_24_412 ();
 sg13g2_fill_1 FILLER_24_414 ();
 sg13g2_fill_1 FILLER_24_430 ();
 sg13g2_decap_8 FILLER_24_439 ();
 sg13g2_fill_2 FILLER_24_446 ();
 sg13g2_decap_4 FILLER_24_474 ();
 sg13g2_fill_1 FILLER_24_478 ();
 sg13g2_fill_2 FILLER_24_488 ();
 sg13g2_fill_1 FILLER_24_502 ();
 sg13g2_fill_2 FILLER_24_526 ();
 sg13g2_fill_1 FILLER_24_528 ();
 sg13g2_fill_1 FILLER_24_544 ();
 sg13g2_decap_4 FILLER_24_551 ();
 sg13g2_fill_2 FILLER_24_555 ();
 sg13g2_decap_4 FILLER_24_574 ();
 sg13g2_fill_2 FILLER_24_590 ();
 sg13g2_fill_1 FILLER_24_592 ();
 sg13g2_fill_1 FILLER_24_649 ();
 sg13g2_fill_2 FILLER_24_676 ();
 sg13g2_fill_1 FILLER_24_678 ();
 sg13g2_fill_2 FILLER_24_699 ();
 sg13g2_fill_2 FILLER_24_713 ();
 sg13g2_fill_1 FILLER_24_715 ();
 sg13g2_fill_2 FILLER_24_744 ();
 sg13g2_fill_1 FILLER_24_746 ();
 sg13g2_fill_2 FILLER_24_772 ();
 sg13g2_fill_1 FILLER_24_774 ();
 sg13g2_fill_2 FILLER_24_783 ();
 sg13g2_decap_4 FILLER_24_790 ();
 sg13g2_fill_1 FILLER_24_794 ();
 sg13g2_decap_8 FILLER_24_841 ();
 sg13g2_decap_4 FILLER_24_848 ();
 sg13g2_fill_2 FILLER_24_852 ();
 sg13g2_fill_1 FILLER_24_876 ();
 sg13g2_decap_8 FILLER_24_881 ();
 sg13g2_fill_1 FILLER_24_888 ();
 sg13g2_fill_2 FILLER_24_897 ();
 sg13g2_decap_8 FILLER_24_911 ();
 sg13g2_fill_2 FILLER_24_918 ();
 sg13g2_fill_2 FILLER_24_937 ();
 sg13g2_fill_1 FILLER_24_939 ();
 sg13g2_fill_1 FILLER_24_950 ();
 sg13g2_fill_2 FILLER_24_970 ();
 sg13g2_decap_8 FILLER_24_977 ();
 sg13g2_fill_1 FILLER_24_998 ();
 sg13g2_fill_2 FILLER_24_1023 ();
 sg13g2_decap_8 FILLER_24_1037 ();
 sg13g2_fill_1 FILLER_24_1044 ();
 sg13g2_fill_1 FILLER_24_1058 ();
 sg13g2_decap_4 FILLER_24_1064 ();
 sg13g2_decap_8 FILLER_24_1074 ();
 sg13g2_fill_1 FILLER_24_1081 ();
 sg13g2_fill_1 FILLER_24_1095 ();
 sg13g2_decap_8 FILLER_24_1122 ();
 sg13g2_decap_8 FILLER_24_1129 ();
 sg13g2_decap_8 FILLER_24_1136 ();
 sg13g2_decap_8 FILLER_24_1143 ();
 sg13g2_decap_8 FILLER_24_1150 ();
 sg13g2_decap_8 FILLER_24_1157 ();
 sg13g2_decap_8 FILLER_24_1164 ();
 sg13g2_decap_8 FILLER_24_1171 ();
 sg13g2_decap_8 FILLER_24_1178 ();
 sg13g2_decap_8 FILLER_24_1185 ();
 sg13g2_decap_8 FILLER_24_1192 ();
 sg13g2_decap_8 FILLER_24_1199 ();
 sg13g2_decap_8 FILLER_24_1206 ();
 sg13g2_decap_8 FILLER_24_1213 ();
 sg13g2_decap_8 FILLER_24_1220 ();
 sg13g2_decap_8 FILLER_24_1227 ();
 sg13g2_decap_8 FILLER_24_1234 ();
 sg13g2_decap_8 FILLER_24_1241 ();
 sg13g2_decap_8 FILLER_24_1248 ();
 sg13g2_decap_8 FILLER_24_1255 ();
 sg13g2_decap_8 FILLER_24_1262 ();
 sg13g2_decap_8 FILLER_24_1269 ();
 sg13g2_decap_8 FILLER_24_1276 ();
 sg13g2_decap_8 FILLER_24_1283 ();
 sg13g2_decap_8 FILLER_24_1290 ();
 sg13g2_decap_8 FILLER_24_1297 ();
 sg13g2_decap_8 FILLER_24_1304 ();
 sg13g2_decap_8 FILLER_24_1311 ();
 sg13g2_decap_8 FILLER_24_1318 ();
 sg13g2_decap_8 FILLER_24_1325 ();
 sg13g2_decap_8 FILLER_24_1332 ();
 sg13g2_decap_8 FILLER_24_1339 ();
 sg13g2_decap_8 FILLER_24_1346 ();
 sg13g2_decap_8 FILLER_24_1353 ();
 sg13g2_decap_8 FILLER_24_1360 ();
 sg13g2_decap_8 FILLER_24_1367 ();
 sg13g2_decap_8 FILLER_24_1374 ();
 sg13g2_decap_8 FILLER_24_1381 ();
 sg13g2_decap_8 FILLER_24_1388 ();
 sg13g2_decap_8 FILLER_24_1395 ();
 sg13g2_decap_8 FILLER_24_1402 ();
 sg13g2_decap_8 FILLER_24_1409 ();
 sg13g2_decap_8 FILLER_24_1416 ();
 sg13g2_decap_8 FILLER_24_1423 ();
 sg13g2_decap_8 FILLER_24_1430 ();
 sg13g2_decap_8 FILLER_24_1437 ();
 sg13g2_decap_8 FILLER_24_1444 ();
 sg13g2_decap_8 FILLER_24_1451 ();
 sg13g2_decap_8 FILLER_24_1458 ();
 sg13g2_decap_8 FILLER_24_1465 ();
 sg13g2_decap_8 FILLER_24_1472 ();
 sg13g2_decap_8 FILLER_24_1479 ();
 sg13g2_decap_8 FILLER_24_1486 ();
 sg13g2_decap_8 FILLER_24_1493 ();
 sg13g2_decap_8 FILLER_24_1500 ();
 sg13g2_decap_8 FILLER_24_1507 ();
 sg13g2_decap_8 FILLER_24_1514 ();
 sg13g2_decap_8 FILLER_24_1521 ();
 sg13g2_decap_8 FILLER_24_1528 ();
 sg13g2_decap_8 FILLER_24_1535 ();
 sg13g2_decap_8 FILLER_24_1542 ();
 sg13g2_decap_8 FILLER_24_1549 ();
 sg13g2_decap_8 FILLER_24_1556 ();
 sg13g2_decap_8 FILLER_24_1563 ();
 sg13g2_decap_8 FILLER_24_1570 ();
 sg13g2_decap_8 FILLER_24_1577 ();
 sg13g2_decap_8 FILLER_24_1584 ();
 sg13g2_decap_8 FILLER_24_1591 ();
 sg13g2_decap_8 FILLER_24_1598 ();
 sg13g2_decap_8 FILLER_24_1605 ();
 sg13g2_decap_8 FILLER_24_1612 ();
 sg13g2_decap_8 FILLER_24_1619 ();
 sg13g2_decap_8 FILLER_24_1626 ();
 sg13g2_decap_8 FILLER_24_1633 ();
 sg13g2_decap_8 FILLER_24_1640 ();
 sg13g2_decap_8 FILLER_24_1647 ();
 sg13g2_decap_8 FILLER_24_1654 ();
 sg13g2_decap_8 FILLER_24_1661 ();
 sg13g2_decap_8 FILLER_24_1668 ();
 sg13g2_decap_8 FILLER_24_1675 ();
 sg13g2_decap_8 FILLER_24_1682 ();
 sg13g2_decap_8 FILLER_24_1689 ();
 sg13g2_decap_8 FILLER_24_1696 ();
 sg13g2_decap_8 FILLER_24_1703 ();
 sg13g2_decap_8 FILLER_24_1710 ();
 sg13g2_decap_8 FILLER_24_1717 ();
 sg13g2_decap_8 FILLER_24_1724 ();
 sg13g2_decap_8 FILLER_24_1731 ();
 sg13g2_decap_8 FILLER_24_1738 ();
 sg13g2_decap_8 FILLER_24_1745 ();
 sg13g2_decap_8 FILLER_24_1752 ();
 sg13g2_decap_8 FILLER_24_1759 ();
 sg13g2_fill_2 FILLER_24_1766 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_4 FILLER_25_49 ();
 sg13g2_fill_1 FILLER_25_53 ();
 sg13g2_fill_2 FILLER_25_80 ();
 sg13g2_fill_1 FILLER_25_82 ();
 sg13g2_decap_4 FILLER_25_157 ();
 sg13g2_decap_4 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_195 ();
 sg13g2_fill_1 FILLER_25_197 ();
 sg13g2_decap_8 FILLER_25_216 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_fill_2 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_decap_4 FILLER_25_283 ();
 sg13g2_fill_2 FILLER_25_287 ();
 sg13g2_fill_1 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_383 ();
 sg13g2_fill_1 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_fill_2 FILLER_25_429 ();
 sg13g2_fill_1 FILLER_25_448 ();
 sg13g2_fill_2 FILLER_25_465 ();
 sg13g2_fill_1 FILLER_25_467 ();
 sg13g2_decap_4 FILLER_25_473 ();
 sg13g2_decap_8 FILLER_25_482 ();
 sg13g2_fill_1 FILLER_25_489 ();
 sg13g2_fill_1 FILLER_25_514 ();
 sg13g2_fill_2 FILLER_25_542 ();
 sg13g2_decap_8 FILLER_25_552 ();
 sg13g2_fill_2 FILLER_25_559 ();
 sg13g2_fill_1 FILLER_25_561 ();
 sg13g2_decap_4 FILLER_25_566 ();
 sg13g2_fill_2 FILLER_25_570 ();
 sg13g2_fill_1 FILLER_25_634 ();
 sg13g2_decap_8 FILLER_25_664 ();
 sg13g2_decap_8 FILLER_25_671 ();
 sg13g2_decap_4 FILLER_25_678 ();
 sg13g2_fill_2 FILLER_25_682 ();
 sg13g2_decap_8 FILLER_25_689 ();
 sg13g2_decap_8 FILLER_25_696 ();
 sg13g2_fill_2 FILLER_25_703 ();
 sg13g2_decap_8 FILLER_25_710 ();
 sg13g2_fill_1 FILLER_25_717 ();
 sg13g2_decap_8 FILLER_25_729 ();
 sg13g2_fill_1 FILLER_25_736 ();
 sg13g2_decap_4 FILLER_25_745 ();
 sg13g2_fill_2 FILLER_25_749 ();
 sg13g2_fill_2 FILLER_25_756 ();
 sg13g2_fill_2 FILLER_25_762 ();
 sg13g2_decap_8 FILLER_25_768 ();
 sg13g2_fill_2 FILLER_25_775 ();
 sg13g2_fill_1 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_4 FILLER_25_800 ();
 sg13g2_fill_1 FILLER_25_804 ();
 sg13g2_fill_2 FILLER_25_820 ();
 sg13g2_fill_1 FILLER_25_822 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_fill_2 FILLER_25_842 ();
 sg13g2_fill_1 FILLER_25_848 ();
 sg13g2_decap_4 FILLER_25_875 ();
 sg13g2_decap_4 FILLER_25_899 ();
 sg13g2_fill_1 FILLER_25_903 ();
 sg13g2_fill_2 FILLER_25_937 ();
 sg13g2_fill_1 FILLER_25_939 ();
 sg13g2_decap_4 FILLER_25_957 ();
 sg13g2_fill_2 FILLER_25_961 ();
 sg13g2_fill_2 FILLER_25_985 ();
 sg13g2_fill_1 FILLER_25_1004 ();
 sg13g2_decap_8 FILLER_25_1040 ();
 sg13g2_fill_1 FILLER_25_1047 ();
 sg13g2_fill_2 FILLER_25_1072 ();
 sg13g2_fill_1 FILLER_25_1074 ();
 sg13g2_decap_8 FILLER_25_1112 ();
 sg13g2_decap_8 FILLER_25_1119 ();
 sg13g2_decap_8 FILLER_25_1126 ();
 sg13g2_decap_8 FILLER_25_1133 ();
 sg13g2_decap_8 FILLER_25_1140 ();
 sg13g2_decap_8 FILLER_25_1147 ();
 sg13g2_decap_8 FILLER_25_1154 ();
 sg13g2_decap_8 FILLER_25_1161 ();
 sg13g2_decap_8 FILLER_25_1168 ();
 sg13g2_decap_8 FILLER_25_1175 ();
 sg13g2_decap_8 FILLER_25_1182 ();
 sg13g2_decap_8 FILLER_25_1189 ();
 sg13g2_decap_8 FILLER_25_1196 ();
 sg13g2_decap_8 FILLER_25_1203 ();
 sg13g2_decap_8 FILLER_25_1210 ();
 sg13g2_decap_8 FILLER_25_1217 ();
 sg13g2_decap_8 FILLER_25_1224 ();
 sg13g2_decap_8 FILLER_25_1231 ();
 sg13g2_decap_8 FILLER_25_1238 ();
 sg13g2_decap_8 FILLER_25_1245 ();
 sg13g2_decap_8 FILLER_25_1252 ();
 sg13g2_decap_8 FILLER_25_1259 ();
 sg13g2_decap_8 FILLER_25_1266 ();
 sg13g2_decap_8 FILLER_25_1273 ();
 sg13g2_decap_8 FILLER_25_1280 ();
 sg13g2_decap_8 FILLER_25_1287 ();
 sg13g2_decap_8 FILLER_25_1294 ();
 sg13g2_decap_8 FILLER_25_1301 ();
 sg13g2_decap_8 FILLER_25_1308 ();
 sg13g2_decap_8 FILLER_25_1315 ();
 sg13g2_decap_8 FILLER_25_1322 ();
 sg13g2_decap_8 FILLER_25_1329 ();
 sg13g2_decap_8 FILLER_25_1336 ();
 sg13g2_decap_8 FILLER_25_1343 ();
 sg13g2_decap_8 FILLER_25_1350 ();
 sg13g2_decap_8 FILLER_25_1357 ();
 sg13g2_decap_8 FILLER_25_1364 ();
 sg13g2_decap_8 FILLER_25_1371 ();
 sg13g2_decap_8 FILLER_25_1378 ();
 sg13g2_decap_8 FILLER_25_1385 ();
 sg13g2_decap_8 FILLER_25_1392 ();
 sg13g2_decap_8 FILLER_25_1399 ();
 sg13g2_decap_8 FILLER_25_1406 ();
 sg13g2_decap_8 FILLER_25_1413 ();
 sg13g2_decap_8 FILLER_25_1420 ();
 sg13g2_decap_8 FILLER_25_1427 ();
 sg13g2_decap_8 FILLER_25_1434 ();
 sg13g2_decap_8 FILLER_25_1441 ();
 sg13g2_decap_8 FILLER_25_1448 ();
 sg13g2_decap_8 FILLER_25_1455 ();
 sg13g2_decap_8 FILLER_25_1462 ();
 sg13g2_decap_8 FILLER_25_1469 ();
 sg13g2_decap_8 FILLER_25_1476 ();
 sg13g2_decap_8 FILLER_25_1483 ();
 sg13g2_decap_8 FILLER_25_1490 ();
 sg13g2_decap_8 FILLER_25_1497 ();
 sg13g2_decap_8 FILLER_25_1504 ();
 sg13g2_decap_8 FILLER_25_1511 ();
 sg13g2_decap_8 FILLER_25_1518 ();
 sg13g2_decap_8 FILLER_25_1525 ();
 sg13g2_decap_8 FILLER_25_1532 ();
 sg13g2_decap_8 FILLER_25_1539 ();
 sg13g2_decap_8 FILLER_25_1546 ();
 sg13g2_decap_8 FILLER_25_1553 ();
 sg13g2_decap_8 FILLER_25_1560 ();
 sg13g2_decap_8 FILLER_25_1567 ();
 sg13g2_decap_8 FILLER_25_1574 ();
 sg13g2_decap_8 FILLER_25_1581 ();
 sg13g2_decap_8 FILLER_25_1588 ();
 sg13g2_decap_8 FILLER_25_1595 ();
 sg13g2_decap_8 FILLER_25_1602 ();
 sg13g2_decap_8 FILLER_25_1609 ();
 sg13g2_decap_8 FILLER_25_1616 ();
 sg13g2_decap_8 FILLER_25_1623 ();
 sg13g2_decap_8 FILLER_25_1630 ();
 sg13g2_decap_8 FILLER_25_1637 ();
 sg13g2_decap_8 FILLER_25_1644 ();
 sg13g2_decap_8 FILLER_25_1651 ();
 sg13g2_decap_8 FILLER_25_1658 ();
 sg13g2_decap_8 FILLER_25_1665 ();
 sg13g2_decap_8 FILLER_25_1672 ();
 sg13g2_decap_8 FILLER_25_1679 ();
 sg13g2_decap_8 FILLER_25_1686 ();
 sg13g2_decap_8 FILLER_25_1693 ();
 sg13g2_decap_8 FILLER_25_1700 ();
 sg13g2_decap_8 FILLER_25_1707 ();
 sg13g2_decap_8 FILLER_25_1714 ();
 sg13g2_decap_8 FILLER_25_1721 ();
 sg13g2_decap_8 FILLER_25_1728 ();
 sg13g2_decap_8 FILLER_25_1735 ();
 sg13g2_decap_8 FILLER_25_1742 ();
 sg13g2_decap_8 FILLER_25_1749 ();
 sg13g2_decap_8 FILLER_25_1756 ();
 sg13g2_decap_4 FILLER_25_1763 ();
 sg13g2_fill_1 FILLER_25_1767 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_108 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_decap_8 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_141 ();
 sg13g2_decap_4 FILLER_26_204 ();
 sg13g2_fill_2 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_222 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_fill_2 FILLER_26_304 ();
 sg13g2_fill_2 FILLER_26_319 ();
 sg13g2_fill_2 FILLER_26_337 ();
 sg13g2_fill_2 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_440 ();
 sg13g2_fill_2 FILLER_26_447 ();
 sg13g2_fill_1 FILLER_26_479 ();
 sg13g2_fill_1 FILLER_26_506 ();
 sg13g2_decap_4 FILLER_26_517 ();
 sg13g2_fill_2 FILLER_26_531 ();
 sg13g2_fill_1 FILLER_26_533 ();
 sg13g2_decap_4 FILLER_26_578 ();
 sg13g2_fill_1 FILLER_26_582 ();
 sg13g2_fill_1 FILLER_26_596 ();
 sg13g2_fill_2 FILLER_26_616 ();
 sg13g2_fill_1 FILLER_26_618 ();
 sg13g2_fill_2 FILLER_26_649 ();
 sg13g2_fill_2 FILLER_26_659 ();
 sg13g2_decap_8 FILLER_26_713 ();
 sg13g2_decap_4 FILLER_26_720 ();
 sg13g2_fill_1 FILLER_26_724 ();
 sg13g2_fill_2 FILLER_26_738 ();
 sg13g2_fill_1 FILLER_26_745 ();
 sg13g2_fill_1 FILLER_26_772 ();
 sg13g2_decap_8 FILLER_26_778 ();
 sg13g2_fill_2 FILLER_26_789 ();
 sg13g2_fill_1 FILLER_26_838 ();
 sg13g2_fill_2 FILLER_26_846 ();
 sg13g2_decap_8 FILLER_26_874 ();
 sg13g2_decap_4 FILLER_26_881 ();
 sg13g2_fill_1 FILLER_26_885 ();
 sg13g2_fill_2 FILLER_26_895 ();
 sg13g2_fill_1 FILLER_26_897 ();
 sg13g2_decap_8 FILLER_26_903 ();
 sg13g2_fill_1 FILLER_26_910 ();
 sg13g2_fill_2 FILLER_26_916 ();
 sg13g2_fill_1 FILLER_26_918 ();
 sg13g2_fill_2 FILLER_26_927 ();
 sg13g2_decap_4 FILLER_26_937 ();
 sg13g2_fill_2 FILLER_26_941 ();
 sg13g2_fill_2 FILLER_26_951 ();
 sg13g2_fill_2 FILLER_26_965 ();
 sg13g2_fill_2 FILLER_26_971 ();
 sg13g2_decap_4 FILLER_26_981 ();
 sg13g2_fill_2 FILLER_26_985 ();
 sg13g2_fill_2 FILLER_26_990 ();
 sg13g2_fill_2 FILLER_26_1004 ();
 sg13g2_fill_2 FILLER_26_1018 ();
 sg13g2_fill_1 FILLER_26_1020 ();
 sg13g2_decap_8 FILLER_26_1026 ();
 sg13g2_decap_8 FILLER_26_1033 ();
 sg13g2_decap_8 FILLER_26_1040 ();
 sg13g2_fill_2 FILLER_26_1047 ();
 sg13g2_fill_1 FILLER_26_1049 ();
 sg13g2_decap_4 FILLER_26_1065 ();
 sg13g2_fill_1 FILLER_26_1069 ();
 sg13g2_fill_1 FILLER_26_1079 ();
 sg13g2_fill_2 FILLER_26_1091 ();
 sg13g2_decap_8 FILLER_26_1119 ();
 sg13g2_decap_8 FILLER_26_1126 ();
 sg13g2_decap_8 FILLER_26_1133 ();
 sg13g2_decap_8 FILLER_26_1140 ();
 sg13g2_decap_8 FILLER_26_1147 ();
 sg13g2_decap_8 FILLER_26_1154 ();
 sg13g2_decap_8 FILLER_26_1161 ();
 sg13g2_decap_8 FILLER_26_1168 ();
 sg13g2_decap_8 FILLER_26_1175 ();
 sg13g2_decap_8 FILLER_26_1182 ();
 sg13g2_decap_8 FILLER_26_1189 ();
 sg13g2_decap_8 FILLER_26_1196 ();
 sg13g2_decap_8 FILLER_26_1203 ();
 sg13g2_decap_8 FILLER_26_1210 ();
 sg13g2_decap_8 FILLER_26_1217 ();
 sg13g2_decap_8 FILLER_26_1224 ();
 sg13g2_decap_8 FILLER_26_1231 ();
 sg13g2_decap_8 FILLER_26_1238 ();
 sg13g2_decap_8 FILLER_26_1245 ();
 sg13g2_decap_8 FILLER_26_1252 ();
 sg13g2_decap_8 FILLER_26_1259 ();
 sg13g2_decap_8 FILLER_26_1266 ();
 sg13g2_decap_8 FILLER_26_1273 ();
 sg13g2_decap_8 FILLER_26_1280 ();
 sg13g2_decap_8 FILLER_26_1287 ();
 sg13g2_decap_8 FILLER_26_1294 ();
 sg13g2_decap_8 FILLER_26_1301 ();
 sg13g2_decap_8 FILLER_26_1308 ();
 sg13g2_decap_8 FILLER_26_1315 ();
 sg13g2_decap_8 FILLER_26_1322 ();
 sg13g2_decap_8 FILLER_26_1329 ();
 sg13g2_decap_8 FILLER_26_1336 ();
 sg13g2_decap_8 FILLER_26_1343 ();
 sg13g2_decap_8 FILLER_26_1350 ();
 sg13g2_decap_8 FILLER_26_1357 ();
 sg13g2_decap_8 FILLER_26_1364 ();
 sg13g2_decap_8 FILLER_26_1371 ();
 sg13g2_decap_8 FILLER_26_1378 ();
 sg13g2_decap_8 FILLER_26_1385 ();
 sg13g2_decap_8 FILLER_26_1392 ();
 sg13g2_decap_8 FILLER_26_1399 ();
 sg13g2_decap_8 FILLER_26_1406 ();
 sg13g2_decap_8 FILLER_26_1413 ();
 sg13g2_decap_8 FILLER_26_1420 ();
 sg13g2_decap_8 FILLER_26_1427 ();
 sg13g2_decap_8 FILLER_26_1434 ();
 sg13g2_decap_8 FILLER_26_1441 ();
 sg13g2_decap_8 FILLER_26_1448 ();
 sg13g2_decap_8 FILLER_26_1455 ();
 sg13g2_decap_8 FILLER_26_1462 ();
 sg13g2_decap_8 FILLER_26_1469 ();
 sg13g2_decap_8 FILLER_26_1476 ();
 sg13g2_decap_8 FILLER_26_1483 ();
 sg13g2_decap_8 FILLER_26_1490 ();
 sg13g2_decap_8 FILLER_26_1497 ();
 sg13g2_decap_8 FILLER_26_1504 ();
 sg13g2_decap_8 FILLER_26_1511 ();
 sg13g2_decap_8 FILLER_26_1518 ();
 sg13g2_decap_8 FILLER_26_1525 ();
 sg13g2_decap_8 FILLER_26_1532 ();
 sg13g2_decap_8 FILLER_26_1539 ();
 sg13g2_decap_8 FILLER_26_1546 ();
 sg13g2_decap_8 FILLER_26_1553 ();
 sg13g2_decap_8 FILLER_26_1560 ();
 sg13g2_decap_8 FILLER_26_1567 ();
 sg13g2_decap_8 FILLER_26_1574 ();
 sg13g2_decap_8 FILLER_26_1581 ();
 sg13g2_decap_8 FILLER_26_1588 ();
 sg13g2_decap_8 FILLER_26_1595 ();
 sg13g2_decap_8 FILLER_26_1602 ();
 sg13g2_decap_8 FILLER_26_1609 ();
 sg13g2_decap_8 FILLER_26_1616 ();
 sg13g2_decap_8 FILLER_26_1623 ();
 sg13g2_decap_8 FILLER_26_1630 ();
 sg13g2_decap_8 FILLER_26_1637 ();
 sg13g2_decap_8 FILLER_26_1644 ();
 sg13g2_decap_8 FILLER_26_1651 ();
 sg13g2_decap_8 FILLER_26_1658 ();
 sg13g2_decap_8 FILLER_26_1665 ();
 sg13g2_decap_8 FILLER_26_1672 ();
 sg13g2_decap_8 FILLER_26_1679 ();
 sg13g2_decap_8 FILLER_26_1686 ();
 sg13g2_decap_8 FILLER_26_1693 ();
 sg13g2_decap_8 FILLER_26_1700 ();
 sg13g2_decap_8 FILLER_26_1707 ();
 sg13g2_decap_8 FILLER_26_1714 ();
 sg13g2_decap_8 FILLER_26_1721 ();
 sg13g2_decap_8 FILLER_26_1728 ();
 sg13g2_decap_8 FILLER_26_1735 ();
 sg13g2_decap_8 FILLER_26_1742 ();
 sg13g2_decap_8 FILLER_26_1749 ();
 sg13g2_decap_8 FILLER_26_1756 ();
 sg13g2_decap_4 FILLER_26_1763 ();
 sg13g2_fill_1 FILLER_26_1767 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_4 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_46 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_247 ();
 sg13g2_decap_4 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_fill_1 FILLER_27_348 ();
 sg13g2_fill_2 FILLER_27_391 ();
 sg13g2_fill_1 FILLER_27_393 ();
 sg13g2_fill_1 FILLER_27_428 ();
 sg13g2_decap_4 FILLER_27_466 ();
 sg13g2_fill_2 FILLER_27_485 ();
 sg13g2_fill_1 FILLER_27_487 ();
 sg13g2_decap_4 FILLER_27_496 ();
 sg13g2_fill_1 FILLER_27_506 ();
 sg13g2_decap_4 FILLER_27_547 ();
 sg13g2_fill_1 FILLER_27_551 ();
 sg13g2_fill_2 FILLER_27_598 ();
 sg13g2_fill_1 FILLER_27_600 ();
 sg13g2_fill_2 FILLER_27_606 ();
 sg13g2_fill_1 FILLER_27_654 ();
 sg13g2_fill_2 FILLER_27_660 ();
 sg13g2_decap_8 FILLER_27_667 ();
 sg13g2_decap_8 FILLER_27_674 ();
 sg13g2_fill_1 FILLER_27_681 ();
 sg13g2_fill_2 FILLER_27_739 ();
 sg13g2_fill_2 FILLER_27_751 ();
 sg13g2_fill_1 FILLER_27_758 ();
 sg13g2_fill_1 FILLER_27_803 ();
 sg13g2_fill_1 FILLER_27_815 ();
 sg13g2_fill_1 FILLER_27_845 ();
 sg13g2_fill_2 FILLER_27_856 ();
 sg13g2_decap_4 FILLER_27_867 ();
 sg13g2_fill_1 FILLER_27_871 ();
 sg13g2_decap_4 FILLER_27_876 ();
 sg13g2_decap_8 FILLER_27_939 ();
 sg13g2_fill_2 FILLER_27_946 ();
 sg13g2_fill_1 FILLER_27_948 ();
 sg13g2_fill_2 FILLER_27_975 ();
 sg13g2_fill_1 FILLER_27_977 ();
 sg13g2_fill_1 FILLER_27_1017 ();
 sg13g2_fill_2 FILLER_27_1049 ();
 sg13g2_fill_1 FILLER_27_1051 ();
 sg13g2_fill_2 FILLER_27_1083 ();
 sg13g2_fill_1 FILLER_27_1085 ();
 sg13g2_fill_2 FILLER_27_1091 ();
 sg13g2_fill_1 FILLER_27_1093 ();
 sg13g2_decap_8 FILLER_27_1124 ();
 sg13g2_decap_8 FILLER_27_1131 ();
 sg13g2_decap_8 FILLER_27_1138 ();
 sg13g2_decap_8 FILLER_27_1145 ();
 sg13g2_decap_8 FILLER_27_1152 ();
 sg13g2_decap_8 FILLER_27_1159 ();
 sg13g2_decap_8 FILLER_27_1166 ();
 sg13g2_decap_8 FILLER_27_1173 ();
 sg13g2_decap_8 FILLER_27_1180 ();
 sg13g2_decap_8 FILLER_27_1187 ();
 sg13g2_decap_8 FILLER_27_1194 ();
 sg13g2_decap_8 FILLER_27_1201 ();
 sg13g2_decap_8 FILLER_27_1208 ();
 sg13g2_decap_8 FILLER_27_1215 ();
 sg13g2_decap_8 FILLER_27_1222 ();
 sg13g2_decap_8 FILLER_27_1229 ();
 sg13g2_decap_8 FILLER_27_1236 ();
 sg13g2_decap_8 FILLER_27_1243 ();
 sg13g2_decap_8 FILLER_27_1250 ();
 sg13g2_decap_8 FILLER_27_1257 ();
 sg13g2_decap_8 FILLER_27_1264 ();
 sg13g2_decap_8 FILLER_27_1271 ();
 sg13g2_decap_8 FILLER_27_1278 ();
 sg13g2_decap_8 FILLER_27_1285 ();
 sg13g2_decap_8 FILLER_27_1292 ();
 sg13g2_decap_8 FILLER_27_1299 ();
 sg13g2_decap_8 FILLER_27_1306 ();
 sg13g2_decap_8 FILLER_27_1313 ();
 sg13g2_decap_8 FILLER_27_1320 ();
 sg13g2_decap_8 FILLER_27_1327 ();
 sg13g2_decap_8 FILLER_27_1334 ();
 sg13g2_decap_8 FILLER_27_1341 ();
 sg13g2_decap_8 FILLER_27_1348 ();
 sg13g2_decap_8 FILLER_27_1355 ();
 sg13g2_decap_8 FILLER_27_1362 ();
 sg13g2_decap_8 FILLER_27_1369 ();
 sg13g2_decap_8 FILLER_27_1376 ();
 sg13g2_decap_8 FILLER_27_1383 ();
 sg13g2_decap_8 FILLER_27_1390 ();
 sg13g2_decap_8 FILLER_27_1397 ();
 sg13g2_decap_8 FILLER_27_1404 ();
 sg13g2_decap_8 FILLER_27_1411 ();
 sg13g2_decap_8 FILLER_27_1418 ();
 sg13g2_decap_8 FILLER_27_1425 ();
 sg13g2_decap_8 FILLER_27_1432 ();
 sg13g2_decap_8 FILLER_27_1439 ();
 sg13g2_decap_8 FILLER_27_1446 ();
 sg13g2_decap_8 FILLER_27_1453 ();
 sg13g2_decap_8 FILLER_27_1460 ();
 sg13g2_decap_8 FILLER_27_1467 ();
 sg13g2_decap_8 FILLER_27_1474 ();
 sg13g2_decap_8 FILLER_27_1481 ();
 sg13g2_decap_8 FILLER_27_1488 ();
 sg13g2_decap_8 FILLER_27_1495 ();
 sg13g2_decap_8 FILLER_27_1502 ();
 sg13g2_decap_8 FILLER_27_1509 ();
 sg13g2_decap_8 FILLER_27_1516 ();
 sg13g2_decap_8 FILLER_27_1523 ();
 sg13g2_decap_8 FILLER_27_1530 ();
 sg13g2_decap_8 FILLER_27_1537 ();
 sg13g2_decap_8 FILLER_27_1544 ();
 sg13g2_decap_8 FILLER_27_1551 ();
 sg13g2_decap_8 FILLER_27_1558 ();
 sg13g2_decap_8 FILLER_27_1565 ();
 sg13g2_decap_8 FILLER_27_1572 ();
 sg13g2_decap_8 FILLER_27_1579 ();
 sg13g2_decap_8 FILLER_27_1586 ();
 sg13g2_decap_8 FILLER_27_1593 ();
 sg13g2_decap_8 FILLER_27_1600 ();
 sg13g2_decap_8 FILLER_27_1607 ();
 sg13g2_decap_8 FILLER_27_1614 ();
 sg13g2_decap_8 FILLER_27_1621 ();
 sg13g2_decap_8 FILLER_27_1628 ();
 sg13g2_decap_8 FILLER_27_1635 ();
 sg13g2_decap_8 FILLER_27_1642 ();
 sg13g2_decap_8 FILLER_27_1649 ();
 sg13g2_decap_8 FILLER_27_1656 ();
 sg13g2_decap_8 FILLER_27_1663 ();
 sg13g2_decap_8 FILLER_27_1670 ();
 sg13g2_decap_8 FILLER_27_1677 ();
 sg13g2_decap_8 FILLER_27_1684 ();
 sg13g2_decap_8 FILLER_27_1691 ();
 sg13g2_decap_8 FILLER_27_1698 ();
 sg13g2_decap_8 FILLER_27_1705 ();
 sg13g2_decap_8 FILLER_27_1712 ();
 sg13g2_decap_8 FILLER_27_1719 ();
 sg13g2_decap_8 FILLER_27_1726 ();
 sg13g2_decap_8 FILLER_27_1733 ();
 sg13g2_decap_8 FILLER_27_1740 ();
 sg13g2_decap_8 FILLER_27_1747 ();
 sg13g2_decap_8 FILLER_27_1754 ();
 sg13g2_decap_8 FILLER_27_1761 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_4 FILLER_28_56 ();
 sg13g2_fill_2 FILLER_28_86 ();
 sg13g2_fill_1 FILLER_28_88 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_2 FILLER_28_201 ();
 sg13g2_decap_4 FILLER_28_250 ();
 sg13g2_fill_1 FILLER_28_263 ();
 sg13g2_fill_1 FILLER_28_275 ();
 sg13g2_decap_4 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_343 ();
 sg13g2_fill_2 FILLER_28_393 ();
 sg13g2_fill_1 FILLER_28_395 ();
 sg13g2_fill_2 FILLER_28_404 ();
 sg13g2_decap_4 FILLER_28_429 ();
 sg13g2_fill_2 FILLER_28_433 ();
 sg13g2_fill_2 FILLER_28_450 ();
 sg13g2_fill_1 FILLER_28_452 ();
 sg13g2_decap_4 FILLER_28_484 ();
 sg13g2_fill_2 FILLER_28_488 ();
 sg13g2_fill_1 FILLER_28_522 ();
 sg13g2_decap_4 FILLER_28_547 ();
 sg13g2_fill_1 FILLER_28_551 ();
 sg13g2_fill_1 FILLER_28_589 ();
 sg13g2_fill_1 FILLER_28_663 ();
 sg13g2_fill_2 FILLER_28_669 ();
 sg13g2_fill_1 FILLER_28_671 ();
 sg13g2_fill_2 FILLER_28_681 ();
 sg13g2_fill_1 FILLER_28_683 ();
 sg13g2_fill_1 FILLER_28_728 ();
 sg13g2_fill_1 FILLER_28_778 ();
 sg13g2_fill_2 FILLER_28_810 ();
 sg13g2_fill_1 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_853 ();
 sg13g2_decap_4 FILLER_28_886 ();
 sg13g2_fill_2 FILLER_28_913 ();
 sg13g2_fill_2 FILLER_28_920 ();
 sg13g2_fill_2 FILLER_28_945 ();
 sg13g2_fill_1 FILLER_28_947 ();
 sg13g2_decap_4 FILLER_28_1002 ();
 sg13g2_fill_1 FILLER_28_1014 ();
 sg13g2_fill_2 FILLER_28_1050 ();
 sg13g2_decap_8 FILLER_28_1124 ();
 sg13g2_decap_8 FILLER_28_1131 ();
 sg13g2_decap_8 FILLER_28_1138 ();
 sg13g2_decap_8 FILLER_28_1145 ();
 sg13g2_decap_8 FILLER_28_1152 ();
 sg13g2_decap_8 FILLER_28_1159 ();
 sg13g2_decap_8 FILLER_28_1166 ();
 sg13g2_decap_8 FILLER_28_1173 ();
 sg13g2_decap_8 FILLER_28_1180 ();
 sg13g2_decap_8 FILLER_28_1187 ();
 sg13g2_decap_8 FILLER_28_1194 ();
 sg13g2_decap_8 FILLER_28_1201 ();
 sg13g2_decap_8 FILLER_28_1208 ();
 sg13g2_decap_8 FILLER_28_1215 ();
 sg13g2_decap_8 FILLER_28_1222 ();
 sg13g2_decap_8 FILLER_28_1229 ();
 sg13g2_decap_8 FILLER_28_1236 ();
 sg13g2_decap_8 FILLER_28_1243 ();
 sg13g2_decap_8 FILLER_28_1250 ();
 sg13g2_decap_8 FILLER_28_1257 ();
 sg13g2_decap_8 FILLER_28_1264 ();
 sg13g2_decap_8 FILLER_28_1271 ();
 sg13g2_decap_8 FILLER_28_1278 ();
 sg13g2_decap_8 FILLER_28_1285 ();
 sg13g2_decap_8 FILLER_28_1292 ();
 sg13g2_decap_8 FILLER_28_1299 ();
 sg13g2_decap_8 FILLER_28_1306 ();
 sg13g2_decap_8 FILLER_28_1313 ();
 sg13g2_decap_8 FILLER_28_1320 ();
 sg13g2_decap_8 FILLER_28_1327 ();
 sg13g2_decap_8 FILLER_28_1334 ();
 sg13g2_decap_8 FILLER_28_1341 ();
 sg13g2_decap_8 FILLER_28_1348 ();
 sg13g2_decap_8 FILLER_28_1355 ();
 sg13g2_decap_8 FILLER_28_1362 ();
 sg13g2_decap_8 FILLER_28_1369 ();
 sg13g2_decap_8 FILLER_28_1376 ();
 sg13g2_decap_8 FILLER_28_1383 ();
 sg13g2_decap_8 FILLER_28_1390 ();
 sg13g2_decap_8 FILLER_28_1397 ();
 sg13g2_decap_8 FILLER_28_1404 ();
 sg13g2_decap_8 FILLER_28_1411 ();
 sg13g2_decap_8 FILLER_28_1418 ();
 sg13g2_decap_8 FILLER_28_1425 ();
 sg13g2_decap_8 FILLER_28_1432 ();
 sg13g2_decap_8 FILLER_28_1439 ();
 sg13g2_decap_8 FILLER_28_1446 ();
 sg13g2_decap_8 FILLER_28_1453 ();
 sg13g2_decap_8 FILLER_28_1460 ();
 sg13g2_decap_8 FILLER_28_1467 ();
 sg13g2_decap_8 FILLER_28_1474 ();
 sg13g2_decap_8 FILLER_28_1481 ();
 sg13g2_decap_8 FILLER_28_1488 ();
 sg13g2_decap_8 FILLER_28_1495 ();
 sg13g2_decap_8 FILLER_28_1502 ();
 sg13g2_decap_8 FILLER_28_1509 ();
 sg13g2_decap_8 FILLER_28_1516 ();
 sg13g2_decap_8 FILLER_28_1523 ();
 sg13g2_decap_8 FILLER_28_1530 ();
 sg13g2_decap_8 FILLER_28_1537 ();
 sg13g2_decap_8 FILLER_28_1544 ();
 sg13g2_decap_8 FILLER_28_1551 ();
 sg13g2_decap_8 FILLER_28_1558 ();
 sg13g2_decap_8 FILLER_28_1565 ();
 sg13g2_decap_8 FILLER_28_1572 ();
 sg13g2_decap_8 FILLER_28_1579 ();
 sg13g2_decap_8 FILLER_28_1586 ();
 sg13g2_decap_8 FILLER_28_1593 ();
 sg13g2_decap_8 FILLER_28_1600 ();
 sg13g2_decap_8 FILLER_28_1607 ();
 sg13g2_decap_8 FILLER_28_1614 ();
 sg13g2_decap_8 FILLER_28_1621 ();
 sg13g2_decap_8 FILLER_28_1628 ();
 sg13g2_decap_8 FILLER_28_1635 ();
 sg13g2_decap_8 FILLER_28_1642 ();
 sg13g2_decap_8 FILLER_28_1649 ();
 sg13g2_decap_8 FILLER_28_1656 ();
 sg13g2_decap_8 FILLER_28_1663 ();
 sg13g2_decap_8 FILLER_28_1670 ();
 sg13g2_decap_8 FILLER_28_1677 ();
 sg13g2_decap_8 FILLER_28_1684 ();
 sg13g2_decap_8 FILLER_28_1691 ();
 sg13g2_decap_8 FILLER_28_1698 ();
 sg13g2_decap_8 FILLER_28_1705 ();
 sg13g2_decap_8 FILLER_28_1712 ();
 sg13g2_decap_8 FILLER_28_1719 ();
 sg13g2_decap_8 FILLER_28_1726 ();
 sg13g2_decap_8 FILLER_28_1733 ();
 sg13g2_decap_8 FILLER_28_1740 ();
 sg13g2_decap_8 FILLER_28_1747 ();
 sg13g2_decap_8 FILLER_28_1754 ();
 sg13g2_decap_8 FILLER_28_1761 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_56 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_decap_8 FILLER_29_162 ();
 sg13g2_decap_4 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_fill_2 FILLER_29_193 ();
 sg13g2_decap_4 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_379 ();
 sg13g2_fill_2 FILLER_29_389 ();
 sg13g2_fill_2 FILLER_29_430 ();
 sg13g2_fill_2 FILLER_29_486 ();
 sg13g2_fill_1 FILLER_29_488 ();
 sg13g2_decap_4 FILLER_29_495 ();
 sg13g2_fill_2 FILLER_29_499 ();
 sg13g2_fill_2 FILLER_29_516 ();
 sg13g2_fill_1 FILLER_29_564 ();
 sg13g2_fill_2 FILLER_29_605 ();
 sg13g2_fill_2 FILLER_29_642 ();
 sg13g2_fill_1 FILLER_29_644 ();
 sg13g2_fill_1 FILLER_29_736 ();
 sg13g2_fill_2 FILLER_29_750 ();
 sg13g2_fill_1 FILLER_29_752 ();
 sg13g2_fill_1 FILLER_29_762 ();
 sg13g2_fill_2 FILLER_29_805 ();
 sg13g2_fill_1 FILLER_29_807 ();
 sg13g2_fill_1 FILLER_29_816 ();
 sg13g2_fill_2 FILLER_29_874 ();
 sg13g2_fill_1 FILLER_29_876 ();
 sg13g2_fill_1 FILLER_29_948 ();
 sg13g2_fill_2 FILLER_29_977 ();
 sg13g2_fill_1 FILLER_29_979 ();
 sg13g2_decap_4 FILLER_29_998 ();
 sg13g2_fill_1 FILLER_29_1002 ();
 sg13g2_fill_2 FILLER_29_1011 ();
 sg13g2_fill_2 FILLER_29_1072 ();
 sg13g2_fill_2 FILLER_29_1083 ();
 sg13g2_fill_1 FILLER_29_1090 ();
 sg13g2_fill_2 FILLER_29_1100 ();
 sg13g2_decap_8 FILLER_29_1133 ();
 sg13g2_decap_8 FILLER_29_1140 ();
 sg13g2_decap_8 FILLER_29_1147 ();
 sg13g2_decap_8 FILLER_29_1154 ();
 sg13g2_decap_8 FILLER_29_1161 ();
 sg13g2_decap_8 FILLER_29_1168 ();
 sg13g2_decap_8 FILLER_29_1175 ();
 sg13g2_decap_8 FILLER_29_1182 ();
 sg13g2_decap_8 FILLER_29_1189 ();
 sg13g2_decap_8 FILLER_29_1196 ();
 sg13g2_decap_8 FILLER_29_1203 ();
 sg13g2_decap_8 FILLER_29_1210 ();
 sg13g2_decap_8 FILLER_29_1217 ();
 sg13g2_decap_8 FILLER_29_1224 ();
 sg13g2_decap_8 FILLER_29_1231 ();
 sg13g2_decap_8 FILLER_29_1238 ();
 sg13g2_decap_8 FILLER_29_1245 ();
 sg13g2_decap_8 FILLER_29_1252 ();
 sg13g2_decap_8 FILLER_29_1259 ();
 sg13g2_decap_8 FILLER_29_1266 ();
 sg13g2_decap_8 FILLER_29_1273 ();
 sg13g2_decap_8 FILLER_29_1280 ();
 sg13g2_decap_8 FILLER_29_1287 ();
 sg13g2_decap_8 FILLER_29_1294 ();
 sg13g2_decap_8 FILLER_29_1301 ();
 sg13g2_decap_8 FILLER_29_1308 ();
 sg13g2_decap_8 FILLER_29_1315 ();
 sg13g2_decap_8 FILLER_29_1322 ();
 sg13g2_decap_8 FILLER_29_1329 ();
 sg13g2_decap_8 FILLER_29_1336 ();
 sg13g2_decap_8 FILLER_29_1343 ();
 sg13g2_decap_8 FILLER_29_1350 ();
 sg13g2_decap_8 FILLER_29_1357 ();
 sg13g2_decap_8 FILLER_29_1364 ();
 sg13g2_decap_8 FILLER_29_1371 ();
 sg13g2_decap_8 FILLER_29_1378 ();
 sg13g2_decap_8 FILLER_29_1385 ();
 sg13g2_decap_8 FILLER_29_1392 ();
 sg13g2_decap_8 FILLER_29_1399 ();
 sg13g2_decap_8 FILLER_29_1406 ();
 sg13g2_decap_8 FILLER_29_1413 ();
 sg13g2_decap_8 FILLER_29_1420 ();
 sg13g2_decap_8 FILLER_29_1427 ();
 sg13g2_decap_8 FILLER_29_1434 ();
 sg13g2_decap_8 FILLER_29_1441 ();
 sg13g2_decap_8 FILLER_29_1448 ();
 sg13g2_decap_8 FILLER_29_1455 ();
 sg13g2_decap_8 FILLER_29_1462 ();
 sg13g2_decap_8 FILLER_29_1469 ();
 sg13g2_decap_8 FILLER_29_1476 ();
 sg13g2_decap_8 FILLER_29_1483 ();
 sg13g2_decap_8 FILLER_29_1490 ();
 sg13g2_decap_8 FILLER_29_1497 ();
 sg13g2_decap_8 FILLER_29_1504 ();
 sg13g2_decap_8 FILLER_29_1511 ();
 sg13g2_decap_8 FILLER_29_1518 ();
 sg13g2_decap_8 FILLER_29_1525 ();
 sg13g2_decap_8 FILLER_29_1532 ();
 sg13g2_decap_8 FILLER_29_1539 ();
 sg13g2_decap_8 FILLER_29_1546 ();
 sg13g2_decap_8 FILLER_29_1553 ();
 sg13g2_decap_8 FILLER_29_1560 ();
 sg13g2_decap_8 FILLER_29_1567 ();
 sg13g2_decap_8 FILLER_29_1574 ();
 sg13g2_decap_8 FILLER_29_1581 ();
 sg13g2_decap_8 FILLER_29_1588 ();
 sg13g2_decap_8 FILLER_29_1595 ();
 sg13g2_decap_8 FILLER_29_1602 ();
 sg13g2_decap_8 FILLER_29_1609 ();
 sg13g2_decap_8 FILLER_29_1616 ();
 sg13g2_decap_8 FILLER_29_1623 ();
 sg13g2_decap_8 FILLER_29_1630 ();
 sg13g2_decap_8 FILLER_29_1637 ();
 sg13g2_decap_8 FILLER_29_1644 ();
 sg13g2_decap_8 FILLER_29_1651 ();
 sg13g2_decap_8 FILLER_29_1658 ();
 sg13g2_decap_8 FILLER_29_1665 ();
 sg13g2_decap_8 FILLER_29_1672 ();
 sg13g2_decap_8 FILLER_29_1679 ();
 sg13g2_decap_8 FILLER_29_1686 ();
 sg13g2_decap_8 FILLER_29_1693 ();
 sg13g2_decap_8 FILLER_29_1700 ();
 sg13g2_decap_8 FILLER_29_1707 ();
 sg13g2_decap_8 FILLER_29_1714 ();
 sg13g2_decap_8 FILLER_29_1721 ();
 sg13g2_decap_8 FILLER_29_1728 ();
 sg13g2_decap_8 FILLER_29_1735 ();
 sg13g2_decap_8 FILLER_29_1742 ();
 sg13g2_decap_8 FILLER_29_1749 ();
 sg13g2_decap_8 FILLER_29_1756 ();
 sg13g2_decap_4 FILLER_29_1763 ();
 sg13g2_fill_1 FILLER_29_1767 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_120 ();
 sg13g2_fill_1 FILLER_30_206 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_224 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_235 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_247 ();
 sg13g2_decap_8 FILLER_30_261 ();
 sg13g2_decap_4 FILLER_30_280 ();
 sg13g2_fill_2 FILLER_30_284 ();
 sg13g2_decap_4 FILLER_30_309 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_decap_8 FILLER_30_330 ();
 sg13g2_decap_4 FILLER_30_337 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_355 ();
 sg13g2_fill_2 FILLER_30_392 ();
 sg13g2_fill_2 FILLER_30_403 ();
 sg13g2_fill_1 FILLER_30_405 ();
 sg13g2_fill_2 FILLER_30_411 ();
 sg13g2_fill_1 FILLER_30_413 ();
 sg13g2_fill_1 FILLER_30_458 ();
 sg13g2_fill_1 FILLER_30_501 ();
 sg13g2_fill_1 FILLER_30_523 ();
 sg13g2_fill_2 FILLER_30_537 ();
 sg13g2_decap_8 FILLER_30_565 ();
 sg13g2_decap_4 FILLER_30_572 ();
 sg13g2_fill_1 FILLER_30_576 ();
 sg13g2_fill_1 FILLER_30_595 ();
 sg13g2_fill_2 FILLER_30_639 ();
 sg13g2_fill_2 FILLER_30_651 ();
 sg13g2_fill_1 FILLER_30_653 ();
 sg13g2_fill_2 FILLER_30_659 ();
 sg13g2_decap_4 FILLER_30_720 ();
 sg13g2_decap_8 FILLER_30_729 ();
 sg13g2_decap_8 FILLER_30_744 ();
 sg13g2_fill_1 FILLER_30_751 ();
 sg13g2_fill_2 FILLER_30_812 ();
 sg13g2_fill_1 FILLER_30_814 ();
 sg13g2_fill_2 FILLER_30_829 ();
 sg13g2_fill_2 FILLER_30_840 ();
 sg13g2_fill_1 FILLER_30_842 ();
 sg13g2_fill_2 FILLER_30_856 ();
 sg13g2_fill_1 FILLER_30_858 ();
 sg13g2_fill_2 FILLER_30_890 ();
 sg13g2_decap_8 FILLER_30_896 ();
 sg13g2_fill_1 FILLER_30_903 ();
 sg13g2_fill_2 FILLER_30_952 ();
 sg13g2_fill_1 FILLER_30_954 ();
 sg13g2_decap_8 FILLER_30_980 ();
 sg13g2_fill_1 FILLER_30_992 ();
 sg13g2_decap_8 FILLER_30_1003 ();
 sg13g2_fill_1 FILLER_30_1010 ();
 sg13g2_fill_2 FILLER_30_1046 ();
 sg13g2_fill_1 FILLER_30_1095 ();
 sg13g2_fill_2 FILLER_30_1101 ();
 sg13g2_fill_1 FILLER_30_1103 ();
 sg13g2_decap_8 FILLER_30_1139 ();
 sg13g2_decap_8 FILLER_30_1146 ();
 sg13g2_decap_8 FILLER_30_1153 ();
 sg13g2_decap_8 FILLER_30_1160 ();
 sg13g2_decap_8 FILLER_30_1167 ();
 sg13g2_decap_8 FILLER_30_1174 ();
 sg13g2_decap_8 FILLER_30_1181 ();
 sg13g2_decap_8 FILLER_30_1188 ();
 sg13g2_decap_8 FILLER_30_1195 ();
 sg13g2_decap_8 FILLER_30_1202 ();
 sg13g2_decap_8 FILLER_30_1209 ();
 sg13g2_decap_8 FILLER_30_1216 ();
 sg13g2_decap_8 FILLER_30_1223 ();
 sg13g2_decap_8 FILLER_30_1230 ();
 sg13g2_decap_8 FILLER_30_1237 ();
 sg13g2_decap_8 FILLER_30_1244 ();
 sg13g2_decap_8 FILLER_30_1251 ();
 sg13g2_decap_8 FILLER_30_1258 ();
 sg13g2_decap_8 FILLER_30_1265 ();
 sg13g2_decap_8 FILLER_30_1272 ();
 sg13g2_decap_8 FILLER_30_1279 ();
 sg13g2_decap_8 FILLER_30_1286 ();
 sg13g2_decap_8 FILLER_30_1293 ();
 sg13g2_decap_8 FILLER_30_1300 ();
 sg13g2_decap_8 FILLER_30_1307 ();
 sg13g2_decap_8 FILLER_30_1314 ();
 sg13g2_decap_8 FILLER_30_1321 ();
 sg13g2_decap_8 FILLER_30_1328 ();
 sg13g2_decap_8 FILLER_30_1335 ();
 sg13g2_decap_8 FILLER_30_1342 ();
 sg13g2_decap_8 FILLER_30_1349 ();
 sg13g2_decap_8 FILLER_30_1356 ();
 sg13g2_decap_8 FILLER_30_1363 ();
 sg13g2_decap_8 FILLER_30_1370 ();
 sg13g2_decap_8 FILLER_30_1377 ();
 sg13g2_decap_8 FILLER_30_1384 ();
 sg13g2_decap_8 FILLER_30_1391 ();
 sg13g2_decap_8 FILLER_30_1398 ();
 sg13g2_decap_8 FILLER_30_1405 ();
 sg13g2_decap_8 FILLER_30_1412 ();
 sg13g2_decap_8 FILLER_30_1419 ();
 sg13g2_decap_8 FILLER_30_1426 ();
 sg13g2_decap_8 FILLER_30_1433 ();
 sg13g2_decap_8 FILLER_30_1440 ();
 sg13g2_decap_8 FILLER_30_1447 ();
 sg13g2_decap_8 FILLER_30_1454 ();
 sg13g2_decap_8 FILLER_30_1461 ();
 sg13g2_decap_8 FILLER_30_1468 ();
 sg13g2_decap_8 FILLER_30_1475 ();
 sg13g2_decap_8 FILLER_30_1482 ();
 sg13g2_decap_8 FILLER_30_1489 ();
 sg13g2_decap_8 FILLER_30_1496 ();
 sg13g2_decap_8 FILLER_30_1503 ();
 sg13g2_decap_8 FILLER_30_1510 ();
 sg13g2_decap_8 FILLER_30_1517 ();
 sg13g2_decap_8 FILLER_30_1524 ();
 sg13g2_decap_8 FILLER_30_1531 ();
 sg13g2_decap_8 FILLER_30_1538 ();
 sg13g2_decap_8 FILLER_30_1545 ();
 sg13g2_decap_8 FILLER_30_1552 ();
 sg13g2_decap_8 FILLER_30_1559 ();
 sg13g2_decap_8 FILLER_30_1566 ();
 sg13g2_decap_8 FILLER_30_1573 ();
 sg13g2_decap_8 FILLER_30_1580 ();
 sg13g2_decap_8 FILLER_30_1587 ();
 sg13g2_decap_8 FILLER_30_1594 ();
 sg13g2_decap_8 FILLER_30_1601 ();
 sg13g2_decap_8 FILLER_30_1608 ();
 sg13g2_decap_8 FILLER_30_1615 ();
 sg13g2_decap_8 FILLER_30_1622 ();
 sg13g2_decap_8 FILLER_30_1629 ();
 sg13g2_decap_8 FILLER_30_1636 ();
 sg13g2_decap_8 FILLER_30_1643 ();
 sg13g2_decap_8 FILLER_30_1650 ();
 sg13g2_decap_8 FILLER_30_1657 ();
 sg13g2_decap_8 FILLER_30_1664 ();
 sg13g2_decap_8 FILLER_30_1671 ();
 sg13g2_decap_8 FILLER_30_1678 ();
 sg13g2_decap_8 FILLER_30_1685 ();
 sg13g2_decap_8 FILLER_30_1692 ();
 sg13g2_decap_8 FILLER_30_1699 ();
 sg13g2_decap_8 FILLER_30_1706 ();
 sg13g2_decap_8 FILLER_30_1713 ();
 sg13g2_decap_8 FILLER_30_1720 ();
 sg13g2_decap_8 FILLER_30_1727 ();
 sg13g2_decap_8 FILLER_30_1734 ();
 sg13g2_decap_8 FILLER_30_1741 ();
 sg13g2_decap_8 FILLER_30_1748 ();
 sg13g2_decap_8 FILLER_30_1755 ();
 sg13g2_decap_4 FILLER_30_1762 ();
 sg13g2_fill_2 FILLER_30_1766 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_decap_4 FILLER_31_69 ();
 sg13g2_fill_2 FILLER_31_73 ();
 sg13g2_decap_4 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_122 ();
 sg13g2_decap_4 FILLER_31_164 ();
 sg13g2_fill_2 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_178 ();
 sg13g2_fill_1 FILLER_31_184 ();
 sg13g2_fill_2 FILLER_31_230 ();
 sg13g2_fill_1 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_339 ();
 sg13g2_fill_1 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_395 ();
 sg13g2_fill_2 FILLER_31_444 ();
 sg13g2_fill_1 FILLER_31_476 ();
 sg13g2_fill_1 FILLER_31_481 ();
 sg13g2_fill_1 FILLER_31_485 ();
 sg13g2_fill_1 FILLER_31_503 ();
 sg13g2_decap_4 FILLER_31_512 ();
 sg13g2_fill_2 FILLER_31_528 ();
 sg13g2_fill_1 FILLER_31_547 ();
 sg13g2_fill_2 FILLER_31_579 ();
 sg13g2_decap_8 FILLER_31_695 ();
 sg13g2_fill_2 FILLER_31_702 ();
 sg13g2_fill_1 FILLER_31_704 ();
 sg13g2_fill_2 FILLER_31_726 ();
 sg13g2_fill_1 FILLER_31_728 ();
 sg13g2_decap_4 FILLER_31_734 ();
 sg13g2_fill_1 FILLER_31_738 ();
 sg13g2_decap_4 FILLER_31_749 ();
 sg13g2_fill_2 FILLER_31_753 ();
 sg13g2_fill_1 FILLER_31_760 ();
 sg13g2_fill_2 FILLER_31_788 ();
 sg13g2_fill_2 FILLER_31_800 ();
 sg13g2_fill_2 FILLER_31_841 ();
 sg13g2_fill_2 FILLER_31_922 ();
 sg13g2_fill_2 FILLER_31_960 ();
 sg13g2_fill_1 FILLER_31_962 ();
 sg13g2_decap_4 FILLER_31_1045 ();
 sg13g2_decap_8 FILLER_31_1067 ();
 sg13g2_fill_2 FILLER_31_1074 ();
 sg13g2_fill_1 FILLER_31_1096 ();
 sg13g2_fill_2 FILLER_31_1106 ();
 sg13g2_fill_1 FILLER_31_1108 ();
 sg13g2_fill_2 FILLER_31_1114 ();
 sg13g2_fill_1 FILLER_31_1116 ();
 sg13g2_decap_8 FILLER_31_1126 ();
 sg13g2_decap_8 FILLER_31_1133 ();
 sg13g2_decap_8 FILLER_31_1140 ();
 sg13g2_decap_8 FILLER_31_1147 ();
 sg13g2_decap_8 FILLER_31_1154 ();
 sg13g2_decap_8 FILLER_31_1161 ();
 sg13g2_decap_8 FILLER_31_1168 ();
 sg13g2_decap_8 FILLER_31_1175 ();
 sg13g2_decap_8 FILLER_31_1182 ();
 sg13g2_decap_8 FILLER_31_1189 ();
 sg13g2_decap_8 FILLER_31_1196 ();
 sg13g2_decap_8 FILLER_31_1203 ();
 sg13g2_decap_8 FILLER_31_1210 ();
 sg13g2_decap_8 FILLER_31_1217 ();
 sg13g2_decap_8 FILLER_31_1224 ();
 sg13g2_decap_8 FILLER_31_1231 ();
 sg13g2_decap_8 FILLER_31_1238 ();
 sg13g2_decap_8 FILLER_31_1245 ();
 sg13g2_decap_8 FILLER_31_1252 ();
 sg13g2_decap_8 FILLER_31_1259 ();
 sg13g2_decap_8 FILLER_31_1266 ();
 sg13g2_decap_8 FILLER_31_1273 ();
 sg13g2_decap_8 FILLER_31_1280 ();
 sg13g2_decap_8 FILLER_31_1287 ();
 sg13g2_decap_8 FILLER_31_1294 ();
 sg13g2_decap_8 FILLER_31_1301 ();
 sg13g2_decap_8 FILLER_31_1308 ();
 sg13g2_decap_8 FILLER_31_1315 ();
 sg13g2_decap_8 FILLER_31_1322 ();
 sg13g2_decap_8 FILLER_31_1329 ();
 sg13g2_decap_8 FILLER_31_1336 ();
 sg13g2_decap_8 FILLER_31_1343 ();
 sg13g2_decap_8 FILLER_31_1350 ();
 sg13g2_decap_8 FILLER_31_1357 ();
 sg13g2_decap_8 FILLER_31_1364 ();
 sg13g2_decap_8 FILLER_31_1371 ();
 sg13g2_decap_8 FILLER_31_1378 ();
 sg13g2_decap_8 FILLER_31_1385 ();
 sg13g2_decap_8 FILLER_31_1392 ();
 sg13g2_decap_8 FILLER_31_1399 ();
 sg13g2_decap_8 FILLER_31_1406 ();
 sg13g2_decap_8 FILLER_31_1413 ();
 sg13g2_decap_8 FILLER_31_1420 ();
 sg13g2_decap_8 FILLER_31_1427 ();
 sg13g2_decap_8 FILLER_31_1434 ();
 sg13g2_decap_8 FILLER_31_1441 ();
 sg13g2_decap_8 FILLER_31_1448 ();
 sg13g2_decap_8 FILLER_31_1455 ();
 sg13g2_decap_8 FILLER_31_1462 ();
 sg13g2_decap_8 FILLER_31_1469 ();
 sg13g2_decap_8 FILLER_31_1476 ();
 sg13g2_decap_8 FILLER_31_1483 ();
 sg13g2_decap_8 FILLER_31_1490 ();
 sg13g2_decap_8 FILLER_31_1497 ();
 sg13g2_decap_8 FILLER_31_1504 ();
 sg13g2_decap_8 FILLER_31_1511 ();
 sg13g2_decap_8 FILLER_31_1518 ();
 sg13g2_decap_8 FILLER_31_1525 ();
 sg13g2_decap_8 FILLER_31_1532 ();
 sg13g2_decap_8 FILLER_31_1539 ();
 sg13g2_decap_8 FILLER_31_1546 ();
 sg13g2_decap_8 FILLER_31_1553 ();
 sg13g2_decap_8 FILLER_31_1560 ();
 sg13g2_decap_8 FILLER_31_1567 ();
 sg13g2_decap_8 FILLER_31_1574 ();
 sg13g2_decap_8 FILLER_31_1581 ();
 sg13g2_decap_8 FILLER_31_1588 ();
 sg13g2_decap_8 FILLER_31_1595 ();
 sg13g2_decap_8 FILLER_31_1602 ();
 sg13g2_decap_8 FILLER_31_1609 ();
 sg13g2_decap_8 FILLER_31_1616 ();
 sg13g2_decap_8 FILLER_31_1623 ();
 sg13g2_decap_8 FILLER_31_1630 ();
 sg13g2_decap_8 FILLER_31_1637 ();
 sg13g2_decap_8 FILLER_31_1644 ();
 sg13g2_decap_8 FILLER_31_1651 ();
 sg13g2_decap_8 FILLER_31_1658 ();
 sg13g2_decap_8 FILLER_31_1665 ();
 sg13g2_decap_8 FILLER_31_1672 ();
 sg13g2_decap_8 FILLER_31_1679 ();
 sg13g2_decap_8 FILLER_31_1686 ();
 sg13g2_decap_8 FILLER_31_1693 ();
 sg13g2_decap_8 FILLER_31_1700 ();
 sg13g2_decap_8 FILLER_31_1707 ();
 sg13g2_decap_8 FILLER_31_1714 ();
 sg13g2_decap_8 FILLER_31_1721 ();
 sg13g2_decap_8 FILLER_31_1728 ();
 sg13g2_decap_8 FILLER_31_1735 ();
 sg13g2_decap_8 FILLER_31_1742 ();
 sg13g2_decap_8 FILLER_31_1749 ();
 sg13g2_decap_8 FILLER_31_1756 ();
 sg13g2_decap_4 FILLER_31_1763 ();
 sg13g2_fill_1 FILLER_31_1767 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_4 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_67 ();
 sg13g2_fill_2 FILLER_32_121 ();
 sg13g2_fill_2 FILLER_32_131 ();
 sg13g2_fill_1 FILLER_32_151 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_fill_2 FILLER_32_211 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_245 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_fill_2 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_fill_2 FILLER_32_316 ();
 sg13g2_decap_4 FILLER_32_336 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_357 ();
 sg13g2_fill_1 FILLER_32_359 ();
 sg13g2_fill_2 FILLER_32_372 ();
 sg13g2_fill_1 FILLER_32_385 ();
 sg13g2_fill_2 FILLER_32_437 ();
 sg13g2_fill_1 FILLER_32_439 ();
 sg13g2_fill_2 FILLER_32_500 ();
 sg13g2_fill_1 FILLER_32_516 ();
 sg13g2_decap_8 FILLER_32_543 ();
 sg13g2_fill_1 FILLER_32_550 ();
 sg13g2_decap_8 FILLER_32_560 ();
 sg13g2_fill_1 FILLER_32_567 ();
 sg13g2_decap_4 FILLER_32_577 ();
 sg13g2_fill_2 FILLER_32_613 ();
 sg13g2_fill_1 FILLER_32_615 ();
 sg13g2_fill_2 FILLER_32_666 ();
 sg13g2_fill_2 FILLER_32_676 ();
 sg13g2_decap_8 FILLER_32_703 ();
 sg13g2_fill_2 FILLER_32_710 ();
 sg13g2_fill_1 FILLER_32_712 ();
 sg13g2_fill_2 FILLER_32_718 ();
 sg13g2_fill_1 FILLER_32_725 ();
 sg13g2_fill_2 FILLER_32_739 ();
 sg13g2_fill_1 FILLER_32_741 ();
 sg13g2_fill_2 FILLER_32_752 ();
 sg13g2_fill_1 FILLER_32_754 ();
 sg13g2_fill_2 FILLER_32_773 ();
 sg13g2_fill_1 FILLER_32_775 ();
 sg13g2_fill_2 FILLER_32_848 ();
 sg13g2_fill_1 FILLER_32_850 ();
 sg13g2_decap_8 FILLER_32_891 ();
 sg13g2_fill_1 FILLER_32_938 ();
 sg13g2_fill_2 FILLER_32_960 ();
 sg13g2_fill_1 FILLER_32_962 ();
 sg13g2_fill_2 FILLER_32_971 ();
 sg13g2_fill_2 FILLER_32_1006 ();
 sg13g2_fill_2 FILLER_32_1048 ();
 sg13g2_fill_1 FILLER_32_1050 ();
 sg13g2_fill_1 FILLER_32_1061 ();
 sg13g2_fill_2 FILLER_32_1111 ();
 sg13g2_decap_8 FILLER_32_1139 ();
 sg13g2_decap_8 FILLER_32_1146 ();
 sg13g2_decap_8 FILLER_32_1153 ();
 sg13g2_decap_8 FILLER_32_1160 ();
 sg13g2_decap_8 FILLER_32_1167 ();
 sg13g2_decap_8 FILLER_32_1174 ();
 sg13g2_decap_8 FILLER_32_1181 ();
 sg13g2_decap_8 FILLER_32_1188 ();
 sg13g2_decap_8 FILLER_32_1195 ();
 sg13g2_decap_8 FILLER_32_1202 ();
 sg13g2_decap_8 FILLER_32_1209 ();
 sg13g2_decap_8 FILLER_32_1216 ();
 sg13g2_decap_8 FILLER_32_1223 ();
 sg13g2_decap_8 FILLER_32_1230 ();
 sg13g2_decap_8 FILLER_32_1237 ();
 sg13g2_decap_8 FILLER_32_1244 ();
 sg13g2_decap_8 FILLER_32_1251 ();
 sg13g2_decap_8 FILLER_32_1258 ();
 sg13g2_decap_8 FILLER_32_1265 ();
 sg13g2_decap_8 FILLER_32_1272 ();
 sg13g2_decap_8 FILLER_32_1279 ();
 sg13g2_decap_8 FILLER_32_1286 ();
 sg13g2_decap_8 FILLER_32_1293 ();
 sg13g2_decap_8 FILLER_32_1300 ();
 sg13g2_decap_8 FILLER_32_1307 ();
 sg13g2_decap_8 FILLER_32_1314 ();
 sg13g2_decap_8 FILLER_32_1321 ();
 sg13g2_decap_8 FILLER_32_1328 ();
 sg13g2_decap_8 FILLER_32_1335 ();
 sg13g2_decap_8 FILLER_32_1342 ();
 sg13g2_decap_8 FILLER_32_1349 ();
 sg13g2_decap_8 FILLER_32_1356 ();
 sg13g2_decap_8 FILLER_32_1363 ();
 sg13g2_decap_8 FILLER_32_1370 ();
 sg13g2_decap_8 FILLER_32_1377 ();
 sg13g2_decap_8 FILLER_32_1384 ();
 sg13g2_decap_8 FILLER_32_1391 ();
 sg13g2_decap_8 FILLER_32_1398 ();
 sg13g2_decap_8 FILLER_32_1405 ();
 sg13g2_decap_8 FILLER_32_1412 ();
 sg13g2_decap_8 FILLER_32_1419 ();
 sg13g2_decap_8 FILLER_32_1426 ();
 sg13g2_decap_8 FILLER_32_1433 ();
 sg13g2_decap_8 FILLER_32_1440 ();
 sg13g2_decap_8 FILLER_32_1447 ();
 sg13g2_decap_8 FILLER_32_1454 ();
 sg13g2_decap_8 FILLER_32_1461 ();
 sg13g2_decap_8 FILLER_32_1468 ();
 sg13g2_decap_8 FILLER_32_1475 ();
 sg13g2_decap_8 FILLER_32_1482 ();
 sg13g2_decap_8 FILLER_32_1489 ();
 sg13g2_decap_8 FILLER_32_1496 ();
 sg13g2_decap_8 FILLER_32_1503 ();
 sg13g2_decap_8 FILLER_32_1510 ();
 sg13g2_decap_8 FILLER_32_1517 ();
 sg13g2_decap_8 FILLER_32_1524 ();
 sg13g2_decap_8 FILLER_32_1531 ();
 sg13g2_decap_8 FILLER_32_1538 ();
 sg13g2_decap_8 FILLER_32_1545 ();
 sg13g2_decap_8 FILLER_32_1552 ();
 sg13g2_decap_8 FILLER_32_1559 ();
 sg13g2_decap_8 FILLER_32_1566 ();
 sg13g2_decap_8 FILLER_32_1573 ();
 sg13g2_decap_8 FILLER_32_1580 ();
 sg13g2_decap_8 FILLER_32_1587 ();
 sg13g2_decap_8 FILLER_32_1594 ();
 sg13g2_decap_8 FILLER_32_1601 ();
 sg13g2_decap_8 FILLER_32_1608 ();
 sg13g2_decap_8 FILLER_32_1615 ();
 sg13g2_decap_8 FILLER_32_1622 ();
 sg13g2_decap_8 FILLER_32_1629 ();
 sg13g2_decap_8 FILLER_32_1636 ();
 sg13g2_decap_8 FILLER_32_1643 ();
 sg13g2_decap_8 FILLER_32_1650 ();
 sg13g2_decap_8 FILLER_32_1657 ();
 sg13g2_decap_8 FILLER_32_1664 ();
 sg13g2_decap_8 FILLER_32_1671 ();
 sg13g2_decap_8 FILLER_32_1678 ();
 sg13g2_decap_8 FILLER_32_1685 ();
 sg13g2_decap_8 FILLER_32_1692 ();
 sg13g2_decap_8 FILLER_32_1699 ();
 sg13g2_decap_8 FILLER_32_1706 ();
 sg13g2_decap_8 FILLER_32_1713 ();
 sg13g2_decap_8 FILLER_32_1720 ();
 sg13g2_decap_8 FILLER_32_1727 ();
 sg13g2_decap_8 FILLER_32_1734 ();
 sg13g2_decap_8 FILLER_32_1741 ();
 sg13g2_decap_8 FILLER_32_1748 ();
 sg13g2_decap_8 FILLER_32_1755 ();
 sg13g2_decap_4 FILLER_32_1762 ();
 sg13g2_fill_2 FILLER_32_1766 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_decap_8 FILLER_33_102 ();
 sg13g2_decap_4 FILLER_33_109 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_fill_2 FILLER_33_129 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_2 FILLER_33_142 ();
 sg13g2_fill_2 FILLER_33_170 ();
 sg13g2_fill_1 FILLER_33_172 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_219 ();
 sg13g2_decap_8 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_233 ();
 sg13g2_decap_4 FILLER_33_240 ();
 sg13g2_decap_4 FILLER_33_262 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_294 ();
 sg13g2_decap_4 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_330 ();
 sg13g2_fill_2 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_33_431 ();
 sg13g2_fill_2 FILLER_33_483 ();
 sg13g2_fill_2 FILLER_33_517 ();
 sg13g2_fill_1 FILLER_33_531 ();
 sg13g2_fill_2 FILLER_33_589 ();
 sg13g2_fill_1 FILLER_33_612 ();
 sg13g2_fill_2 FILLER_33_621 ();
 sg13g2_fill_1 FILLER_33_623 ();
 sg13g2_fill_1 FILLER_33_638 ();
 sg13g2_fill_2 FILLER_33_709 ();
 sg13g2_fill_1 FILLER_33_711 ();
 sg13g2_fill_1 FILLER_33_738 ();
 sg13g2_fill_2 FILLER_33_753 ();
 sg13g2_fill_1 FILLER_33_773 ();
 sg13g2_decap_4 FILLER_33_810 ();
 sg13g2_fill_1 FILLER_33_814 ();
 sg13g2_fill_2 FILLER_33_832 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_fill_1 FILLER_33_862 ();
 sg13g2_fill_1 FILLER_33_917 ();
 sg13g2_fill_1 FILLER_33_926 ();
 sg13g2_decap_4 FILLER_33_1000 ();
 sg13g2_fill_1 FILLER_33_1004 ();
 sg13g2_fill_1 FILLER_33_1008 ();
 sg13g2_decap_8 FILLER_33_1019 ();
 sg13g2_decap_4 FILLER_33_1026 ();
 sg13g2_fill_2 FILLER_33_1030 ();
 sg13g2_decap_8 FILLER_33_1050 ();
 sg13g2_decap_4 FILLER_33_1057 ();
 sg13g2_decap_4 FILLER_33_1079 ();
 sg13g2_fill_1 FILLER_33_1088 ();
 sg13g2_fill_1 FILLER_33_1099 ();
 sg13g2_decap_8 FILLER_33_1145 ();
 sg13g2_decap_8 FILLER_33_1152 ();
 sg13g2_decap_8 FILLER_33_1159 ();
 sg13g2_decap_8 FILLER_33_1166 ();
 sg13g2_decap_8 FILLER_33_1173 ();
 sg13g2_decap_8 FILLER_33_1180 ();
 sg13g2_decap_8 FILLER_33_1187 ();
 sg13g2_decap_8 FILLER_33_1194 ();
 sg13g2_decap_8 FILLER_33_1201 ();
 sg13g2_decap_8 FILLER_33_1208 ();
 sg13g2_decap_8 FILLER_33_1215 ();
 sg13g2_decap_8 FILLER_33_1222 ();
 sg13g2_decap_8 FILLER_33_1229 ();
 sg13g2_decap_8 FILLER_33_1236 ();
 sg13g2_decap_8 FILLER_33_1243 ();
 sg13g2_decap_8 FILLER_33_1250 ();
 sg13g2_decap_8 FILLER_33_1257 ();
 sg13g2_decap_8 FILLER_33_1264 ();
 sg13g2_decap_8 FILLER_33_1271 ();
 sg13g2_decap_8 FILLER_33_1278 ();
 sg13g2_decap_8 FILLER_33_1285 ();
 sg13g2_decap_8 FILLER_33_1292 ();
 sg13g2_decap_8 FILLER_33_1299 ();
 sg13g2_decap_8 FILLER_33_1306 ();
 sg13g2_decap_8 FILLER_33_1313 ();
 sg13g2_decap_8 FILLER_33_1320 ();
 sg13g2_decap_8 FILLER_33_1327 ();
 sg13g2_decap_8 FILLER_33_1334 ();
 sg13g2_decap_8 FILLER_33_1341 ();
 sg13g2_decap_8 FILLER_33_1348 ();
 sg13g2_decap_8 FILLER_33_1355 ();
 sg13g2_decap_8 FILLER_33_1362 ();
 sg13g2_decap_8 FILLER_33_1369 ();
 sg13g2_decap_8 FILLER_33_1376 ();
 sg13g2_decap_8 FILLER_33_1383 ();
 sg13g2_decap_8 FILLER_33_1390 ();
 sg13g2_decap_8 FILLER_33_1397 ();
 sg13g2_decap_8 FILLER_33_1404 ();
 sg13g2_decap_8 FILLER_33_1411 ();
 sg13g2_decap_8 FILLER_33_1418 ();
 sg13g2_decap_8 FILLER_33_1425 ();
 sg13g2_decap_8 FILLER_33_1432 ();
 sg13g2_decap_8 FILLER_33_1439 ();
 sg13g2_decap_8 FILLER_33_1446 ();
 sg13g2_decap_8 FILLER_33_1453 ();
 sg13g2_decap_8 FILLER_33_1460 ();
 sg13g2_decap_8 FILLER_33_1467 ();
 sg13g2_decap_8 FILLER_33_1474 ();
 sg13g2_decap_8 FILLER_33_1481 ();
 sg13g2_decap_8 FILLER_33_1488 ();
 sg13g2_decap_8 FILLER_33_1495 ();
 sg13g2_decap_8 FILLER_33_1502 ();
 sg13g2_decap_8 FILLER_33_1509 ();
 sg13g2_decap_8 FILLER_33_1516 ();
 sg13g2_decap_8 FILLER_33_1523 ();
 sg13g2_decap_8 FILLER_33_1530 ();
 sg13g2_decap_8 FILLER_33_1537 ();
 sg13g2_decap_8 FILLER_33_1544 ();
 sg13g2_decap_8 FILLER_33_1551 ();
 sg13g2_decap_8 FILLER_33_1558 ();
 sg13g2_decap_8 FILLER_33_1565 ();
 sg13g2_decap_8 FILLER_33_1572 ();
 sg13g2_decap_8 FILLER_33_1579 ();
 sg13g2_decap_8 FILLER_33_1586 ();
 sg13g2_decap_8 FILLER_33_1593 ();
 sg13g2_decap_8 FILLER_33_1600 ();
 sg13g2_decap_8 FILLER_33_1607 ();
 sg13g2_decap_8 FILLER_33_1614 ();
 sg13g2_decap_8 FILLER_33_1621 ();
 sg13g2_decap_8 FILLER_33_1628 ();
 sg13g2_decap_8 FILLER_33_1635 ();
 sg13g2_decap_8 FILLER_33_1642 ();
 sg13g2_decap_8 FILLER_33_1649 ();
 sg13g2_decap_8 FILLER_33_1656 ();
 sg13g2_decap_8 FILLER_33_1663 ();
 sg13g2_decap_8 FILLER_33_1670 ();
 sg13g2_decap_8 FILLER_33_1677 ();
 sg13g2_decap_8 FILLER_33_1684 ();
 sg13g2_decap_8 FILLER_33_1691 ();
 sg13g2_decap_8 FILLER_33_1698 ();
 sg13g2_decap_8 FILLER_33_1705 ();
 sg13g2_decap_8 FILLER_33_1712 ();
 sg13g2_decap_8 FILLER_33_1719 ();
 sg13g2_decap_8 FILLER_33_1726 ();
 sg13g2_decap_8 FILLER_33_1733 ();
 sg13g2_decap_8 FILLER_33_1740 ();
 sg13g2_decap_8 FILLER_33_1747 ();
 sg13g2_decap_8 FILLER_33_1754 ();
 sg13g2_decap_8 FILLER_33_1761 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_4 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_88 ();
 sg13g2_decap_4 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_decap_4 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_162 ();
 sg13g2_fill_2 FILLER_34_174 ();
 sg13g2_decap_4 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_288 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_fill_2 FILLER_34_340 ();
 sg13g2_fill_2 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_370 ();
 sg13g2_fill_1 FILLER_34_393 ();
 sg13g2_decap_4 FILLER_34_416 ();
 sg13g2_decap_4 FILLER_34_437 ();
 sg13g2_decap_8 FILLER_34_454 ();
 sg13g2_fill_2 FILLER_34_461 ();
 sg13g2_fill_1 FILLER_34_493 ();
 sg13g2_decap_4 FILLER_34_602 ();
 sg13g2_decap_4 FILLER_34_620 ();
 sg13g2_fill_2 FILLER_34_664 ();
 sg13g2_fill_2 FILLER_34_670 ();
 sg13g2_fill_1 FILLER_34_685 ();
 sg13g2_fill_1 FILLER_34_699 ();
 sg13g2_fill_2 FILLER_34_715 ();
 sg13g2_decap_4 FILLER_34_737 ();
 sg13g2_fill_2 FILLER_34_741 ();
 sg13g2_fill_2 FILLER_34_758 ();
 sg13g2_fill_1 FILLER_34_760 ();
 sg13g2_fill_2 FILLER_34_776 ();
 sg13g2_fill_1 FILLER_34_778 ();
 sg13g2_decap_4 FILLER_34_801 ();
 sg13g2_fill_1 FILLER_34_805 ();
 sg13g2_decap_4 FILLER_34_815 ();
 sg13g2_fill_1 FILLER_34_862 ();
 sg13g2_fill_2 FILLER_34_904 ();
 sg13g2_fill_1 FILLER_34_906 ();
 sg13g2_fill_2 FILLER_34_915 ();
 sg13g2_decap_8 FILLER_34_921 ();
 sg13g2_decap_8 FILLER_34_928 ();
 sg13g2_fill_1 FILLER_34_935 ();
 sg13g2_fill_2 FILLER_34_958 ();
 sg13g2_fill_1 FILLER_34_979 ();
 sg13g2_fill_2 FILLER_34_998 ();
 sg13g2_fill_1 FILLER_34_1008 ();
 sg13g2_fill_2 FILLER_34_1029 ();
 sg13g2_fill_2 FILLER_34_1057 ();
 sg13g2_fill_1 FILLER_34_1059 ();
 sg13g2_decap_8 FILLER_34_1134 ();
 sg13g2_decap_8 FILLER_34_1141 ();
 sg13g2_decap_8 FILLER_34_1148 ();
 sg13g2_decap_8 FILLER_34_1155 ();
 sg13g2_decap_8 FILLER_34_1162 ();
 sg13g2_decap_8 FILLER_34_1169 ();
 sg13g2_decap_8 FILLER_34_1176 ();
 sg13g2_decap_8 FILLER_34_1183 ();
 sg13g2_decap_8 FILLER_34_1190 ();
 sg13g2_decap_8 FILLER_34_1197 ();
 sg13g2_decap_8 FILLER_34_1204 ();
 sg13g2_decap_8 FILLER_34_1211 ();
 sg13g2_decap_8 FILLER_34_1218 ();
 sg13g2_decap_8 FILLER_34_1225 ();
 sg13g2_decap_8 FILLER_34_1232 ();
 sg13g2_decap_8 FILLER_34_1239 ();
 sg13g2_decap_8 FILLER_34_1246 ();
 sg13g2_decap_8 FILLER_34_1253 ();
 sg13g2_decap_8 FILLER_34_1260 ();
 sg13g2_decap_8 FILLER_34_1267 ();
 sg13g2_decap_8 FILLER_34_1274 ();
 sg13g2_decap_8 FILLER_34_1281 ();
 sg13g2_decap_8 FILLER_34_1288 ();
 sg13g2_decap_8 FILLER_34_1295 ();
 sg13g2_decap_8 FILLER_34_1302 ();
 sg13g2_decap_8 FILLER_34_1309 ();
 sg13g2_decap_8 FILLER_34_1316 ();
 sg13g2_decap_8 FILLER_34_1323 ();
 sg13g2_decap_8 FILLER_34_1330 ();
 sg13g2_decap_8 FILLER_34_1337 ();
 sg13g2_decap_8 FILLER_34_1344 ();
 sg13g2_decap_8 FILLER_34_1351 ();
 sg13g2_decap_8 FILLER_34_1358 ();
 sg13g2_decap_8 FILLER_34_1365 ();
 sg13g2_decap_8 FILLER_34_1372 ();
 sg13g2_decap_8 FILLER_34_1379 ();
 sg13g2_decap_8 FILLER_34_1386 ();
 sg13g2_decap_8 FILLER_34_1393 ();
 sg13g2_decap_8 FILLER_34_1400 ();
 sg13g2_decap_8 FILLER_34_1407 ();
 sg13g2_decap_8 FILLER_34_1414 ();
 sg13g2_decap_8 FILLER_34_1421 ();
 sg13g2_decap_8 FILLER_34_1428 ();
 sg13g2_decap_8 FILLER_34_1435 ();
 sg13g2_decap_8 FILLER_34_1442 ();
 sg13g2_decap_8 FILLER_34_1449 ();
 sg13g2_decap_8 FILLER_34_1456 ();
 sg13g2_decap_8 FILLER_34_1463 ();
 sg13g2_decap_8 FILLER_34_1470 ();
 sg13g2_decap_8 FILLER_34_1477 ();
 sg13g2_decap_8 FILLER_34_1484 ();
 sg13g2_decap_8 FILLER_34_1491 ();
 sg13g2_decap_8 FILLER_34_1498 ();
 sg13g2_decap_8 FILLER_34_1505 ();
 sg13g2_decap_8 FILLER_34_1512 ();
 sg13g2_decap_8 FILLER_34_1519 ();
 sg13g2_decap_8 FILLER_34_1526 ();
 sg13g2_decap_8 FILLER_34_1533 ();
 sg13g2_decap_8 FILLER_34_1540 ();
 sg13g2_decap_8 FILLER_34_1547 ();
 sg13g2_decap_8 FILLER_34_1554 ();
 sg13g2_decap_8 FILLER_34_1561 ();
 sg13g2_decap_8 FILLER_34_1568 ();
 sg13g2_decap_8 FILLER_34_1575 ();
 sg13g2_decap_8 FILLER_34_1582 ();
 sg13g2_decap_8 FILLER_34_1589 ();
 sg13g2_decap_8 FILLER_34_1596 ();
 sg13g2_decap_8 FILLER_34_1603 ();
 sg13g2_decap_8 FILLER_34_1610 ();
 sg13g2_decap_8 FILLER_34_1617 ();
 sg13g2_decap_8 FILLER_34_1624 ();
 sg13g2_decap_8 FILLER_34_1631 ();
 sg13g2_decap_8 FILLER_34_1638 ();
 sg13g2_decap_8 FILLER_34_1645 ();
 sg13g2_decap_8 FILLER_34_1652 ();
 sg13g2_decap_8 FILLER_34_1659 ();
 sg13g2_decap_8 FILLER_34_1666 ();
 sg13g2_decap_8 FILLER_34_1673 ();
 sg13g2_decap_8 FILLER_34_1680 ();
 sg13g2_decap_8 FILLER_34_1687 ();
 sg13g2_decap_8 FILLER_34_1694 ();
 sg13g2_decap_8 FILLER_34_1701 ();
 sg13g2_decap_8 FILLER_34_1708 ();
 sg13g2_decap_8 FILLER_34_1715 ();
 sg13g2_decap_8 FILLER_34_1722 ();
 sg13g2_decap_8 FILLER_34_1729 ();
 sg13g2_decap_8 FILLER_34_1736 ();
 sg13g2_decap_8 FILLER_34_1743 ();
 sg13g2_decap_8 FILLER_34_1750 ();
 sg13g2_decap_8 FILLER_34_1757 ();
 sg13g2_decap_4 FILLER_34_1764 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_105 ();
 sg13g2_fill_1 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_decap_4 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_206 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_decap_8 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_236 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_1 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_285 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_369 ();
 sg13g2_fill_1 FILLER_35_371 ();
 sg13g2_decap_4 FILLER_35_382 ();
 sg13g2_fill_1 FILLER_35_386 ();
 sg13g2_decap_4 FILLER_35_399 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_430 ();
 sg13g2_fill_1 FILLER_35_445 ();
 sg13g2_decap_4 FILLER_35_458 ();
 sg13g2_fill_1 FILLER_35_470 ();
 sg13g2_decap_8 FILLER_35_479 ();
 sg13g2_decap_8 FILLER_35_486 ();
 sg13g2_fill_2 FILLER_35_531 ();
 sg13g2_fill_1 FILLER_35_575 ();
 sg13g2_fill_1 FILLER_35_605 ();
 sg13g2_decap_8 FILLER_35_621 ();
 sg13g2_decap_4 FILLER_35_628 ();
 sg13g2_fill_1 FILLER_35_632 ();
 sg13g2_decap_4 FILLER_35_641 ();
 sg13g2_fill_2 FILLER_35_645 ();
 sg13g2_fill_1 FILLER_35_653 ();
 sg13g2_fill_2 FILLER_35_664 ();
 sg13g2_decap_4 FILLER_35_676 ();
 sg13g2_fill_2 FILLER_35_690 ();
 sg13g2_decap_4 FILLER_35_711 ();
 sg13g2_fill_2 FILLER_35_715 ();
 sg13g2_decap_4 FILLER_35_764 ();
 sg13g2_decap_8 FILLER_35_778 ();
 sg13g2_decap_4 FILLER_35_785 ();
 sg13g2_fill_1 FILLER_35_789 ();
 sg13g2_fill_1 FILLER_35_816 ();
 sg13g2_fill_1 FILLER_35_826 ();
 sg13g2_decap_4 FILLER_35_831 ();
 sg13g2_fill_1 FILLER_35_835 ();
 sg13g2_fill_2 FILLER_35_844 ();
 sg13g2_decap_4 FILLER_35_856 ();
 sg13g2_fill_2 FILLER_35_865 ();
 sg13g2_decap_8 FILLER_35_898 ();
 sg13g2_fill_2 FILLER_35_905 ();
 sg13g2_decap_4 FILLER_35_925 ();
 sg13g2_decap_4 FILLER_35_957 ();
 sg13g2_fill_1 FILLER_35_961 ();
 sg13g2_decap_8 FILLER_35_967 ();
 sg13g2_decap_4 FILLER_35_974 ();
 sg13g2_fill_2 FILLER_35_1041 ();
 sg13g2_fill_1 FILLER_35_1043 ();
 sg13g2_decap_8 FILLER_35_1054 ();
 sg13g2_fill_2 FILLER_35_1061 ();
 sg13g2_fill_2 FILLER_35_1083 ();
 sg13g2_fill_1 FILLER_35_1085 ();
 sg13g2_decap_8 FILLER_35_1092 ();
 sg13g2_fill_1 FILLER_35_1102 ();
 sg13g2_decap_8 FILLER_35_1140 ();
 sg13g2_decap_8 FILLER_35_1147 ();
 sg13g2_decap_8 FILLER_35_1154 ();
 sg13g2_decap_8 FILLER_35_1161 ();
 sg13g2_decap_8 FILLER_35_1168 ();
 sg13g2_decap_8 FILLER_35_1175 ();
 sg13g2_decap_8 FILLER_35_1182 ();
 sg13g2_decap_8 FILLER_35_1189 ();
 sg13g2_decap_8 FILLER_35_1196 ();
 sg13g2_decap_8 FILLER_35_1203 ();
 sg13g2_decap_8 FILLER_35_1210 ();
 sg13g2_decap_8 FILLER_35_1217 ();
 sg13g2_decap_8 FILLER_35_1224 ();
 sg13g2_decap_8 FILLER_35_1231 ();
 sg13g2_decap_8 FILLER_35_1238 ();
 sg13g2_decap_8 FILLER_35_1245 ();
 sg13g2_decap_8 FILLER_35_1252 ();
 sg13g2_decap_8 FILLER_35_1259 ();
 sg13g2_decap_8 FILLER_35_1266 ();
 sg13g2_decap_8 FILLER_35_1273 ();
 sg13g2_decap_8 FILLER_35_1280 ();
 sg13g2_decap_8 FILLER_35_1287 ();
 sg13g2_decap_8 FILLER_35_1294 ();
 sg13g2_decap_8 FILLER_35_1301 ();
 sg13g2_decap_8 FILLER_35_1308 ();
 sg13g2_decap_8 FILLER_35_1315 ();
 sg13g2_decap_8 FILLER_35_1322 ();
 sg13g2_decap_8 FILLER_35_1329 ();
 sg13g2_decap_8 FILLER_35_1336 ();
 sg13g2_decap_8 FILLER_35_1343 ();
 sg13g2_decap_8 FILLER_35_1350 ();
 sg13g2_decap_8 FILLER_35_1357 ();
 sg13g2_decap_8 FILLER_35_1364 ();
 sg13g2_decap_8 FILLER_35_1371 ();
 sg13g2_decap_8 FILLER_35_1378 ();
 sg13g2_decap_8 FILLER_35_1385 ();
 sg13g2_decap_8 FILLER_35_1392 ();
 sg13g2_decap_8 FILLER_35_1399 ();
 sg13g2_decap_8 FILLER_35_1406 ();
 sg13g2_decap_8 FILLER_35_1413 ();
 sg13g2_decap_8 FILLER_35_1420 ();
 sg13g2_decap_8 FILLER_35_1427 ();
 sg13g2_decap_8 FILLER_35_1434 ();
 sg13g2_decap_8 FILLER_35_1441 ();
 sg13g2_decap_8 FILLER_35_1448 ();
 sg13g2_decap_8 FILLER_35_1455 ();
 sg13g2_decap_8 FILLER_35_1462 ();
 sg13g2_decap_8 FILLER_35_1469 ();
 sg13g2_decap_8 FILLER_35_1476 ();
 sg13g2_decap_8 FILLER_35_1483 ();
 sg13g2_decap_8 FILLER_35_1490 ();
 sg13g2_decap_8 FILLER_35_1497 ();
 sg13g2_decap_8 FILLER_35_1504 ();
 sg13g2_decap_8 FILLER_35_1511 ();
 sg13g2_decap_8 FILLER_35_1518 ();
 sg13g2_decap_8 FILLER_35_1525 ();
 sg13g2_decap_8 FILLER_35_1532 ();
 sg13g2_decap_8 FILLER_35_1539 ();
 sg13g2_decap_8 FILLER_35_1546 ();
 sg13g2_decap_8 FILLER_35_1553 ();
 sg13g2_decap_8 FILLER_35_1560 ();
 sg13g2_decap_8 FILLER_35_1567 ();
 sg13g2_decap_8 FILLER_35_1574 ();
 sg13g2_decap_8 FILLER_35_1581 ();
 sg13g2_decap_8 FILLER_35_1588 ();
 sg13g2_decap_8 FILLER_35_1595 ();
 sg13g2_decap_8 FILLER_35_1602 ();
 sg13g2_decap_8 FILLER_35_1609 ();
 sg13g2_decap_8 FILLER_35_1616 ();
 sg13g2_decap_8 FILLER_35_1623 ();
 sg13g2_decap_8 FILLER_35_1630 ();
 sg13g2_decap_8 FILLER_35_1637 ();
 sg13g2_decap_8 FILLER_35_1644 ();
 sg13g2_decap_8 FILLER_35_1651 ();
 sg13g2_decap_8 FILLER_35_1658 ();
 sg13g2_decap_8 FILLER_35_1665 ();
 sg13g2_decap_8 FILLER_35_1672 ();
 sg13g2_decap_8 FILLER_35_1679 ();
 sg13g2_decap_8 FILLER_35_1686 ();
 sg13g2_decap_8 FILLER_35_1693 ();
 sg13g2_decap_8 FILLER_35_1700 ();
 sg13g2_decap_8 FILLER_35_1707 ();
 sg13g2_decap_8 FILLER_35_1714 ();
 sg13g2_decap_8 FILLER_35_1721 ();
 sg13g2_decap_8 FILLER_35_1728 ();
 sg13g2_decap_8 FILLER_35_1735 ();
 sg13g2_decap_8 FILLER_35_1742 ();
 sg13g2_decap_8 FILLER_35_1749 ();
 sg13g2_decap_8 FILLER_35_1756 ();
 sg13g2_decap_4 FILLER_35_1763 ();
 sg13g2_fill_1 FILLER_35_1767 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_4 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_130 ();
 sg13g2_decap_8 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_180 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_fill_2 FILLER_36_216 ();
 sg13g2_decap_4 FILLER_36_295 ();
 sg13g2_decap_8 FILLER_36_304 ();
 sg13g2_decap_4 FILLER_36_311 ();
 sg13g2_decap_4 FILLER_36_341 ();
 sg13g2_decap_4 FILLER_36_353 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_fill_1 FILLER_36_373 ();
 sg13g2_fill_2 FILLER_36_398 ();
 sg13g2_fill_2 FILLER_36_414 ();
 sg13g2_decap_8 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_450 ();
 sg13g2_fill_2 FILLER_36_465 ();
 sg13g2_fill_1 FILLER_36_467 ();
 sg13g2_fill_2 FILLER_36_490 ();
 sg13g2_fill_2 FILLER_36_501 ();
 sg13g2_fill_1 FILLER_36_503 ();
 sg13g2_decap_8 FILLER_36_523 ();
 sg13g2_decap_4 FILLER_36_530 ();
 sg13g2_fill_1 FILLER_36_555 ();
 sg13g2_decap_4 FILLER_36_593 ();
 sg13g2_fill_2 FILLER_36_626 ();
 sg13g2_fill_1 FILLER_36_641 ();
 sg13g2_fill_1 FILLER_36_656 ();
 sg13g2_decap_4 FILLER_36_669 ();
 sg13g2_fill_2 FILLER_36_673 ();
 sg13g2_decap_4 FILLER_36_711 ();
 sg13g2_fill_1 FILLER_36_715 ();
 sg13g2_fill_2 FILLER_36_728 ();
 sg13g2_decap_8 FILLER_36_751 ();
 sg13g2_fill_2 FILLER_36_758 ();
 sg13g2_fill_2 FILLER_36_809 ();
 sg13g2_fill_2 FILLER_36_864 ();
 sg13g2_fill_1 FILLER_36_866 ();
 sg13g2_decap_4 FILLER_36_907 ();
 sg13g2_fill_2 FILLER_36_911 ();
 sg13g2_decap_4 FILLER_36_921 ();
 sg13g2_fill_1 FILLER_36_925 ();
 sg13g2_fill_2 FILLER_36_938 ();
 sg13g2_decap_8 FILLER_36_950 ();
 sg13g2_decap_8 FILLER_36_957 ();
 sg13g2_fill_2 FILLER_36_964 ();
 sg13g2_fill_1 FILLER_36_966 ();
 sg13g2_fill_1 FILLER_36_978 ();
 sg13g2_fill_1 FILLER_36_1014 ();
 sg13g2_decap_4 FILLER_36_1041 ();
 sg13g2_decap_4 FILLER_36_1049 ();
 sg13g2_fill_1 FILLER_36_1053 ();
 sg13g2_fill_2 FILLER_36_1082 ();
 sg13g2_decap_8 FILLER_36_1147 ();
 sg13g2_decap_8 FILLER_36_1154 ();
 sg13g2_decap_8 FILLER_36_1161 ();
 sg13g2_decap_8 FILLER_36_1168 ();
 sg13g2_decap_8 FILLER_36_1175 ();
 sg13g2_decap_8 FILLER_36_1182 ();
 sg13g2_decap_8 FILLER_36_1189 ();
 sg13g2_decap_8 FILLER_36_1196 ();
 sg13g2_decap_8 FILLER_36_1203 ();
 sg13g2_decap_8 FILLER_36_1210 ();
 sg13g2_decap_8 FILLER_36_1217 ();
 sg13g2_decap_8 FILLER_36_1224 ();
 sg13g2_decap_8 FILLER_36_1231 ();
 sg13g2_decap_8 FILLER_36_1238 ();
 sg13g2_decap_8 FILLER_36_1245 ();
 sg13g2_decap_8 FILLER_36_1252 ();
 sg13g2_decap_8 FILLER_36_1259 ();
 sg13g2_decap_8 FILLER_36_1266 ();
 sg13g2_decap_8 FILLER_36_1273 ();
 sg13g2_decap_8 FILLER_36_1280 ();
 sg13g2_decap_8 FILLER_36_1287 ();
 sg13g2_decap_8 FILLER_36_1294 ();
 sg13g2_decap_8 FILLER_36_1301 ();
 sg13g2_decap_8 FILLER_36_1308 ();
 sg13g2_decap_8 FILLER_36_1315 ();
 sg13g2_decap_8 FILLER_36_1322 ();
 sg13g2_decap_8 FILLER_36_1329 ();
 sg13g2_decap_8 FILLER_36_1336 ();
 sg13g2_decap_8 FILLER_36_1343 ();
 sg13g2_decap_8 FILLER_36_1350 ();
 sg13g2_decap_8 FILLER_36_1357 ();
 sg13g2_decap_8 FILLER_36_1364 ();
 sg13g2_decap_8 FILLER_36_1371 ();
 sg13g2_decap_8 FILLER_36_1378 ();
 sg13g2_decap_8 FILLER_36_1385 ();
 sg13g2_decap_8 FILLER_36_1392 ();
 sg13g2_decap_8 FILLER_36_1399 ();
 sg13g2_decap_8 FILLER_36_1406 ();
 sg13g2_decap_8 FILLER_36_1413 ();
 sg13g2_decap_8 FILLER_36_1420 ();
 sg13g2_decap_8 FILLER_36_1427 ();
 sg13g2_decap_8 FILLER_36_1434 ();
 sg13g2_decap_8 FILLER_36_1441 ();
 sg13g2_decap_8 FILLER_36_1448 ();
 sg13g2_decap_8 FILLER_36_1455 ();
 sg13g2_decap_8 FILLER_36_1462 ();
 sg13g2_decap_8 FILLER_36_1469 ();
 sg13g2_decap_8 FILLER_36_1476 ();
 sg13g2_decap_8 FILLER_36_1483 ();
 sg13g2_decap_8 FILLER_36_1490 ();
 sg13g2_decap_8 FILLER_36_1497 ();
 sg13g2_decap_8 FILLER_36_1504 ();
 sg13g2_decap_8 FILLER_36_1511 ();
 sg13g2_decap_8 FILLER_36_1518 ();
 sg13g2_decap_8 FILLER_36_1525 ();
 sg13g2_decap_8 FILLER_36_1532 ();
 sg13g2_decap_8 FILLER_36_1539 ();
 sg13g2_decap_8 FILLER_36_1546 ();
 sg13g2_decap_8 FILLER_36_1553 ();
 sg13g2_decap_8 FILLER_36_1560 ();
 sg13g2_decap_8 FILLER_36_1567 ();
 sg13g2_decap_8 FILLER_36_1574 ();
 sg13g2_decap_8 FILLER_36_1581 ();
 sg13g2_decap_8 FILLER_36_1588 ();
 sg13g2_decap_8 FILLER_36_1595 ();
 sg13g2_decap_8 FILLER_36_1602 ();
 sg13g2_decap_8 FILLER_36_1609 ();
 sg13g2_decap_8 FILLER_36_1616 ();
 sg13g2_decap_8 FILLER_36_1623 ();
 sg13g2_decap_8 FILLER_36_1630 ();
 sg13g2_decap_8 FILLER_36_1637 ();
 sg13g2_decap_8 FILLER_36_1644 ();
 sg13g2_decap_8 FILLER_36_1651 ();
 sg13g2_decap_8 FILLER_36_1658 ();
 sg13g2_decap_8 FILLER_36_1665 ();
 sg13g2_decap_8 FILLER_36_1672 ();
 sg13g2_decap_8 FILLER_36_1679 ();
 sg13g2_decap_8 FILLER_36_1686 ();
 sg13g2_decap_8 FILLER_36_1693 ();
 sg13g2_decap_8 FILLER_36_1700 ();
 sg13g2_decap_8 FILLER_36_1707 ();
 sg13g2_decap_8 FILLER_36_1714 ();
 sg13g2_decap_8 FILLER_36_1721 ();
 sg13g2_decap_8 FILLER_36_1728 ();
 sg13g2_decap_8 FILLER_36_1735 ();
 sg13g2_decap_8 FILLER_36_1742 ();
 sg13g2_decap_8 FILLER_36_1749 ();
 sg13g2_decap_8 FILLER_36_1756 ();
 sg13g2_decap_4 FILLER_36_1763 ();
 sg13g2_fill_1 FILLER_36_1767 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_187 ();
 sg13g2_fill_2 FILLER_37_202 ();
 sg13g2_fill_1 FILLER_37_268 ();
 sg13g2_decap_8 FILLER_37_279 ();
 sg13g2_fill_1 FILLER_37_286 ();
 sg13g2_decap_4 FILLER_37_292 ();
 sg13g2_decap_4 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_4 FILLER_37_369 ();
 sg13g2_fill_1 FILLER_37_402 ();
 sg13g2_fill_2 FILLER_37_409 ();
 sg13g2_decap_8 FILLER_37_452 ();
 sg13g2_fill_2 FILLER_37_459 ();
 sg13g2_decap_4 FILLER_37_532 ();
 sg13g2_fill_2 FILLER_37_561 ();
 sg13g2_fill_1 FILLER_37_563 ();
 sg13g2_fill_1 FILLER_37_603 ();
 sg13g2_decap_4 FILLER_37_642 ();
 sg13g2_decap_4 FILLER_37_661 ();
 sg13g2_fill_1 FILLER_37_665 ();
 sg13g2_fill_2 FILLER_37_685 ();
 sg13g2_fill_1 FILLER_37_706 ();
 sg13g2_fill_2 FILLER_37_712 ();
 sg13g2_fill_1 FILLER_37_714 ();
 sg13g2_fill_1 FILLER_37_720 ();
 sg13g2_fill_1 FILLER_37_729 ();
 sg13g2_fill_1 FILLER_37_743 ();
 sg13g2_fill_2 FILLER_37_759 ();
 sg13g2_fill_1 FILLER_37_761 ();
 sg13g2_decap_8 FILLER_37_773 ();
 sg13g2_fill_1 FILLER_37_780 ();
 sg13g2_decap_4 FILLER_37_839 ();
 sg13g2_fill_2 FILLER_37_852 ();
 sg13g2_fill_2 FILLER_37_928 ();
 sg13g2_fill_1 FILLER_37_930 ();
 sg13g2_fill_2 FILLER_37_945 ();
 sg13g2_decap_4 FILLER_37_960 ();
 sg13g2_fill_1 FILLER_37_964 ();
 sg13g2_decap_4 FILLER_37_980 ();
 sg13g2_fill_1 FILLER_37_984 ();
 sg13g2_decap_8 FILLER_37_998 ();
 sg13g2_fill_1 FILLER_37_1005 ();
 sg13g2_decap_8 FILLER_37_1019 ();
 sg13g2_fill_2 FILLER_37_1026 ();
 sg13g2_fill_1 FILLER_37_1060 ();
 sg13g2_fill_2 FILLER_37_1072 ();
 sg13g2_decap_8 FILLER_37_1131 ();
 sg13g2_decap_8 FILLER_37_1138 ();
 sg13g2_decap_8 FILLER_37_1145 ();
 sg13g2_decap_8 FILLER_37_1152 ();
 sg13g2_decap_8 FILLER_37_1159 ();
 sg13g2_decap_8 FILLER_37_1166 ();
 sg13g2_decap_8 FILLER_37_1173 ();
 sg13g2_decap_8 FILLER_37_1180 ();
 sg13g2_decap_8 FILLER_37_1187 ();
 sg13g2_decap_8 FILLER_37_1194 ();
 sg13g2_decap_8 FILLER_37_1201 ();
 sg13g2_decap_8 FILLER_37_1208 ();
 sg13g2_decap_8 FILLER_37_1215 ();
 sg13g2_decap_8 FILLER_37_1222 ();
 sg13g2_decap_8 FILLER_37_1229 ();
 sg13g2_decap_8 FILLER_37_1236 ();
 sg13g2_decap_8 FILLER_37_1243 ();
 sg13g2_decap_8 FILLER_37_1250 ();
 sg13g2_decap_8 FILLER_37_1257 ();
 sg13g2_decap_8 FILLER_37_1264 ();
 sg13g2_decap_8 FILLER_37_1271 ();
 sg13g2_decap_8 FILLER_37_1278 ();
 sg13g2_decap_8 FILLER_37_1285 ();
 sg13g2_decap_8 FILLER_37_1292 ();
 sg13g2_decap_8 FILLER_37_1299 ();
 sg13g2_decap_8 FILLER_37_1306 ();
 sg13g2_decap_8 FILLER_37_1313 ();
 sg13g2_decap_8 FILLER_37_1320 ();
 sg13g2_decap_8 FILLER_37_1327 ();
 sg13g2_decap_8 FILLER_37_1334 ();
 sg13g2_decap_8 FILLER_37_1341 ();
 sg13g2_decap_8 FILLER_37_1348 ();
 sg13g2_decap_8 FILLER_37_1355 ();
 sg13g2_decap_8 FILLER_37_1362 ();
 sg13g2_decap_8 FILLER_37_1369 ();
 sg13g2_decap_8 FILLER_37_1376 ();
 sg13g2_decap_8 FILLER_37_1383 ();
 sg13g2_decap_8 FILLER_37_1390 ();
 sg13g2_decap_8 FILLER_37_1397 ();
 sg13g2_decap_8 FILLER_37_1404 ();
 sg13g2_decap_8 FILLER_37_1411 ();
 sg13g2_decap_8 FILLER_37_1418 ();
 sg13g2_decap_8 FILLER_37_1425 ();
 sg13g2_decap_8 FILLER_37_1432 ();
 sg13g2_decap_8 FILLER_37_1439 ();
 sg13g2_decap_8 FILLER_37_1446 ();
 sg13g2_decap_8 FILLER_37_1453 ();
 sg13g2_decap_8 FILLER_37_1460 ();
 sg13g2_decap_8 FILLER_37_1467 ();
 sg13g2_decap_8 FILLER_37_1474 ();
 sg13g2_decap_8 FILLER_37_1481 ();
 sg13g2_decap_8 FILLER_37_1488 ();
 sg13g2_decap_8 FILLER_37_1495 ();
 sg13g2_decap_8 FILLER_37_1502 ();
 sg13g2_decap_8 FILLER_37_1509 ();
 sg13g2_decap_8 FILLER_37_1516 ();
 sg13g2_decap_8 FILLER_37_1523 ();
 sg13g2_decap_8 FILLER_37_1530 ();
 sg13g2_decap_8 FILLER_37_1537 ();
 sg13g2_decap_8 FILLER_37_1544 ();
 sg13g2_decap_8 FILLER_37_1551 ();
 sg13g2_decap_8 FILLER_37_1558 ();
 sg13g2_decap_8 FILLER_37_1565 ();
 sg13g2_decap_8 FILLER_37_1572 ();
 sg13g2_decap_8 FILLER_37_1579 ();
 sg13g2_decap_8 FILLER_37_1586 ();
 sg13g2_decap_8 FILLER_37_1593 ();
 sg13g2_decap_8 FILLER_37_1600 ();
 sg13g2_decap_8 FILLER_37_1607 ();
 sg13g2_decap_8 FILLER_37_1614 ();
 sg13g2_decap_8 FILLER_37_1621 ();
 sg13g2_decap_8 FILLER_37_1628 ();
 sg13g2_decap_8 FILLER_37_1635 ();
 sg13g2_decap_8 FILLER_37_1642 ();
 sg13g2_decap_8 FILLER_37_1649 ();
 sg13g2_decap_8 FILLER_37_1656 ();
 sg13g2_decap_8 FILLER_37_1663 ();
 sg13g2_decap_8 FILLER_37_1670 ();
 sg13g2_decap_8 FILLER_37_1677 ();
 sg13g2_decap_8 FILLER_37_1684 ();
 sg13g2_decap_8 FILLER_37_1691 ();
 sg13g2_decap_8 FILLER_37_1698 ();
 sg13g2_decap_8 FILLER_37_1705 ();
 sg13g2_decap_8 FILLER_37_1712 ();
 sg13g2_decap_8 FILLER_37_1719 ();
 sg13g2_decap_8 FILLER_37_1726 ();
 sg13g2_decap_8 FILLER_37_1733 ();
 sg13g2_decap_8 FILLER_37_1740 ();
 sg13g2_decap_8 FILLER_37_1747 ();
 sg13g2_decap_8 FILLER_37_1754 ();
 sg13g2_decap_8 FILLER_37_1761 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_fill_2 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_138 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_fill_2 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_300 ();
 sg13g2_decap_4 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_325 ();
 sg13g2_decap_4 FILLER_38_351 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_fill_2 FILLER_38_371 ();
 sg13g2_fill_1 FILLER_38_427 ();
 sg13g2_decap_4 FILLER_38_446 ();
 sg13g2_fill_2 FILLER_38_450 ();
 sg13g2_fill_1 FILLER_38_477 ();
 sg13g2_fill_2 FILLER_38_486 ();
 sg13g2_decap_4 FILLER_38_517 ();
 sg13g2_decap_8 FILLER_38_530 ();
 sg13g2_decap_4 FILLER_38_537 ();
 sg13g2_fill_2 FILLER_38_550 ();
 sg13g2_decap_4 FILLER_38_566 ();
 sg13g2_fill_1 FILLER_38_570 ();
 sg13g2_fill_1 FILLER_38_598 ();
 sg13g2_decap_8 FILLER_38_643 ();
 sg13g2_decap_4 FILLER_38_650 ();
 sg13g2_fill_1 FILLER_38_662 ();
 sg13g2_fill_2 FILLER_38_709 ();
 sg13g2_fill_1 FILLER_38_721 ();
 sg13g2_fill_2 FILLER_38_740 ();
 sg13g2_fill_2 FILLER_38_747 ();
 sg13g2_decap_4 FILLER_38_772 ();
 sg13g2_fill_2 FILLER_38_786 ();
 sg13g2_fill_1 FILLER_38_788 ();
 sg13g2_fill_1 FILLER_38_798 ();
 sg13g2_fill_2 FILLER_38_805 ();
 sg13g2_fill_2 FILLER_38_827 ();
 sg13g2_fill_2 FILLER_38_860 ();
 sg13g2_decap_8 FILLER_38_867 ();
 sg13g2_decap_4 FILLER_38_874 ();
 sg13g2_fill_1 FILLER_38_878 ();
 sg13g2_decap_4 FILLER_38_888 ();
 sg13g2_fill_2 FILLER_38_892 ();
 sg13g2_decap_4 FILLER_38_898 ();
 sg13g2_fill_1 FILLER_38_902 ();
 sg13g2_fill_1 FILLER_38_908 ();
 sg13g2_decap_8 FILLER_38_923 ();
 sg13g2_decap_8 FILLER_38_957 ();
 sg13g2_decap_4 FILLER_38_964 ();
 sg13g2_fill_1 FILLER_38_968 ();
 sg13g2_fill_1 FILLER_38_981 ();
 sg13g2_decap_4 FILLER_38_1034 ();
 sg13g2_fill_1 FILLER_38_1038 ();
 sg13g2_decap_4 FILLER_38_1049 ();
 sg13g2_fill_2 FILLER_38_1053 ();
 sg13g2_fill_2 FILLER_38_1060 ();
 sg13g2_fill_1 FILLER_38_1062 ();
 sg13g2_fill_2 FILLER_38_1110 ();
 sg13g2_fill_1 FILLER_38_1112 ();
 sg13g2_decap_8 FILLER_38_1139 ();
 sg13g2_decap_8 FILLER_38_1146 ();
 sg13g2_decap_8 FILLER_38_1153 ();
 sg13g2_decap_8 FILLER_38_1160 ();
 sg13g2_decap_8 FILLER_38_1167 ();
 sg13g2_decap_8 FILLER_38_1174 ();
 sg13g2_decap_8 FILLER_38_1181 ();
 sg13g2_decap_8 FILLER_38_1188 ();
 sg13g2_decap_8 FILLER_38_1195 ();
 sg13g2_decap_8 FILLER_38_1202 ();
 sg13g2_decap_8 FILLER_38_1209 ();
 sg13g2_decap_8 FILLER_38_1216 ();
 sg13g2_decap_8 FILLER_38_1223 ();
 sg13g2_decap_8 FILLER_38_1230 ();
 sg13g2_decap_8 FILLER_38_1237 ();
 sg13g2_decap_8 FILLER_38_1244 ();
 sg13g2_decap_8 FILLER_38_1251 ();
 sg13g2_decap_8 FILLER_38_1258 ();
 sg13g2_decap_8 FILLER_38_1265 ();
 sg13g2_decap_8 FILLER_38_1272 ();
 sg13g2_decap_8 FILLER_38_1279 ();
 sg13g2_decap_8 FILLER_38_1286 ();
 sg13g2_decap_8 FILLER_38_1293 ();
 sg13g2_decap_8 FILLER_38_1300 ();
 sg13g2_decap_8 FILLER_38_1307 ();
 sg13g2_decap_8 FILLER_38_1314 ();
 sg13g2_decap_8 FILLER_38_1321 ();
 sg13g2_decap_8 FILLER_38_1328 ();
 sg13g2_decap_8 FILLER_38_1335 ();
 sg13g2_decap_8 FILLER_38_1342 ();
 sg13g2_decap_8 FILLER_38_1349 ();
 sg13g2_decap_8 FILLER_38_1356 ();
 sg13g2_decap_8 FILLER_38_1363 ();
 sg13g2_decap_8 FILLER_38_1370 ();
 sg13g2_decap_8 FILLER_38_1377 ();
 sg13g2_decap_8 FILLER_38_1384 ();
 sg13g2_decap_8 FILLER_38_1391 ();
 sg13g2_decap_8 FILLER_38_1398 ();
 sg13g2_decap_8 FILLER_38_1405 ();
 sg13g2_decap_8 FILLER_38_1412 ();
 sg13g2_decap_8 FILLER_38_1419 ();
 sg13g2_decap_8 FILLER_38_1426 ();
 sg13g2_decap_8 FILLER_38_1433 ();
 sg13g2_decap_8 FILLER_38_1440 ();
 sg13g2_decap_8 FILLER_38_1447 ();
 sg13g2_decap_8 FILLER_38_1454 ();
 sg13g2_decap_8 FILLER_38_1461 ();
 sg13g2_decap_8 FILLER_38_1468 ();
 sg13g2_decap_8 FILLER_38_1475 ();
 sg13g2_decap_8 FILLER_38_1482 ();
 sg13g2_decap_8 FILLER_38_1489 ();
 sg13g2_decap_8 FILLER_38_1496 ();
 sg13g2_decap_8 FILLER_38_1503 ();
 sg13g2_decap_8 FILLER_38_1510 ();
 sg13g2_decap_8 FILLER_38_1517 ();
 sg13g2_decap_8 FILLER_38_1524 ();
 sg13g2_decap_8 FILLER_38_1531 ();
 sg13g2_decap_8 FILLER_38_1538 ();
 sg13g2_decap_8 FILLER_38_1545 ();
 sg13g2_decap_8 FILLER_38_1552 ();
 sg13g2_decap_8 FILLER_38_1559 ();
 sg13g2_decap_8 FILLER_38_1566 ();
 sg13g2_decap_8 FILLER_38_1573 ();
 sg13g2_decap_8 FILLER_38_1580 ();
 sg13g2_decap_8 FILLER_38_1587 ();
 sg13g2_decap_8 FILLER_38_1594 ();
 sg13g2_decap_8 FILLER_38_1601 ();
 sg13g2_decap_8 FILLER_38_1608 ();
 sg13g2_decap_8 FILLER_38_1615 ();
 sg13g2_decap_8 FILLER_38_1622 ();
 sg13g2_decap_8 FILLER_38_1629 ();
 sg13g2_decap_8 FILLER_38_1636 ();
 sg13g2_decap_8 FILLER_38_1643 ();
 sg13g2_decap_8 FILLER_38_1650 ();
 sg13g2_decap_8 FILLER_38_1657 ();
 sg13g2_decap_8 FILLER_38_1664 ();
 sg13g2_decap_8 FILLER_38_1671 ();
 sg13g2_decap_8 FILLER_38_1678 ();
 sg13g2_decap_8 FILLER_38_1685 ();
 sg13g2_decap_8 FILLER_38_1692 ();
 sg13g2_decap_8 FILLER_38_1699 ();
 sg13g2_decap_8 FILLER_38_1706 ();
 sg13g2_decap_8 FILLER_38_1713 ();
 sg13g2_decap_8 FILLER_38_1720 ();
 sg13g2_decap_8 FILLER_38_1727 ();
 sg13g2_decap_8 FILLER_38_1734 ();
 sg13g2_decap_8 FILLER_38_1741 ();
 sg13g2_decap_8 FILLER_38_1748 ();
 sg13g2_decap_8 FILLER_38_1755 ();
 sg13g2_decap_4 FILLER_38_1762 ();
 sg13g2_fill_2 FILLER_38_1766 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_4 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_161 ();
 sg13g2_fill_2 FILLER_39_188 ();
 sg13g2_fill_2 FILLER_39_249 ();
 sg13g2_fill_1 FILLER_39_251 ();
 sg13g2_fill_2 FILLER_39_265 ();
 sg13g2_fill_2 FILLER_39_277 ();
 sg13g2_fill_1 FILLER_39_279 ();
 sg13g2_fill_2 FILLER_39_343 ();
 sg13g2_fill_1 FILLER_39_345 ();
 sg13g2_fill_2 FILLER_39_358 ();
 sg13g2_decap_4 FILLER_39_380 ();
 sg13g2_fill_2 FILLER_39_384 ();
 sg13g2_fill_2 FILLER_39_443 ();
 sg13g2_fill_1 FILLER_39_445 ();
 sg13g2_decap_8 FILLER_39_454 ();
 sg13g2_decap_4 FILLER_39_461 ();
 sg13g2_decap_4 FILLER_39_471 ();
 sg13g2_decap_4 FILLER_39_489 ();
 sg13g2_fill_2 FILLER_39_498 ();
 sg13g2_decap_8 FILLER_39_508 ();
 sg13g2_fill_2 FILLER_39_515 ();
 sg13g2_decap_8 FILLER_39_537 ();
 sg13g2_fill_2 FILLER_39_544 ();
 sg13g2_fill_2 FILLER_39_555 ();
 sg13g2_fill_1 FILLER_39_557 ();
 sg13g2_fill_2 FILLER_39_570 ();
 sg13g2_fill_1 FILLER_39_572 ();
 sg13g2_fill_2 FILLER_39_593 ();
 sg13g2_fill_2 FILLER_39_613 ();
 sg13g2_fill_2 FILLER_39_624 ();
 sg13g2_decap_4 FILLER_39_677 ();
 sg13g2_fill_2 FILLER_39_687 ();
 sg13g2_fill_2 FILLER_39_704 ();
 sg13g2_fill_1 FILLER_39_706 ();
 sg13g2_decap_8 FILLER_39_717 ();
 sg13g2_fill_2 FILLER_39_729 ();
 sg13g2_decap_4 FILLER_39_747 ();
 sg13g2_fill_2 FILLER_39_751 ();
 sg13g2_fill_2 FILLER_39_812 ();
 sg13g2_fill_1 FILLER_39_814 ();
 sg13g2_fill_2 FILLER_39_824 ();
 sg13g2_fill_1 FILLER_39_826 ();
 sg13g2_fill_2 FILLER_39_835 ();
 sg13g2_decap_4 FILLER_39_852 ();
 sg13g2_fill_1 FILLER_39_864 ();
 sg13g2_fill_1 FILLER_39_896 ();
 sg13g2_fill_1 FILLER_39_907 ();
 sg13g2_decap_4 FILLER_39_940 ();
 sg13g2_fill_2 FILLER_39_954 ();
 sg13g2_fill_1 FILLER_39_956 ();
 sg13g2_fill_1 FILLER_39_987 ();
 sg13g2_decap_8 FILLER_39_997 ();
 sg13g2_fill_1 FILLER_39_1004 ();
 sg13g2_fill_2 FILLER_39_1013 ();
 sg13g2_fill_1 FILLER_39_1015 ();
 sg13g2_fill_2 FILLER_39_1020 ();
 sg13g2_fill_1 FILLER_39_1022 ();
 sg13g2_fill_1 FILLER_39_1033 ();
 sg13g2_fill_1 FILLER_39_1056 ();
 sg13g2_fill_2 FILLER_39_1067 ();
 sg13g2_fill_1 FILLER_39_1088 ();
 sg13g2_decap_8 FILLER_39_1135 ();
 sg13g2_decap_8 FILLER_39_1142 ();
 sg13g2_decap_8 FILLER_39_1149 ();
 sg13g2_decap_8 FILLER_39_1156 ();
 sg13g2_decap_8 FILLER_39_1163 ();
 sg13g2_decap_8 FILLER_39_1170 ();
 sg13g2_decap_8 FILLER_39_1177 ();
 sg13g2_decap_8 FILLER_39_1184 ();
 sg13g2_decap_8 FILLER_39_1191 ();
 sg13g2_decap_8 FILLER_39_1198 ();
 sg13g2_decap_8 FILLER_39_1205 ();
 sg13g2_decap_8 FILLER_39_1212 ();
 sg13g2_decap_8 FILLER_39_1219 ();
 sg13g2_decap_8 FILLER_39_1226 ();
 sg13g2_decap_8 FILLER_39_1233 ();
 sg13g2_decap_8 FILLER_39_1240 ();
 sg13g2_decap_8 FILLER_39_1247 ();
 sg13g2_decap_8 FILLER_39_1254 ();
 sg13g2_decap_8 FILLER_39_1261 ();
 sg13g2_decap_8 FILLER_39_1268 ();
 sg13g2_decap_8 FILLER_39_1275 ();
 sg13g2_decap_8 FILLER_39_1282 ();
 sg13g2_decap_8 FILLER_39_1289 ();
 sg13g2_decap_8 FILLER_39_1296 ();
 sg13g2_decap_8 FILLER_39_1303 ();
 sg13g2_decap_8 FILLER_39_1310 ();
 sg13g2_decap_8 FILLER_39_1317 ();
 sg13g2_decap_8 FILLER_39_1324 ();
 sg13g2_decap_8 FILLER_39_1331 ();
 sg13g2_decap_8 FILLER_39_1338 ();
 sg13g2_decap_8 FILLER_39_1345 ();
 sg13g2_decap_8 FILLER_39_1352 ();
 sg13g2_decap_8 FILLER_39_1359 ();
 sg13g2_decap_8 FILLER_39_1366 ();
 sg13g2_decap_8 FILLER_39_1373 ();
 sg13g2_decap_8 FILLER_39_1380 ();
 sg13g2_decap_8 FILLER_39_1387 ();
 sg13g2_decap_8 FILLER_39_1394 ();
 sg13g2_decap_8 FILLER_39_1401 ();
 sg13g2_decap_8 FILLER_39_1408 ();
 sg13g2_decap_8 FILLER_39_1415 ();
 sg13g2_decap_8 FILLER_39_1422 ();
 sg13g2_decap_8 FILLER_39_1429 ();
 sg13g2_decap_8 FILLER_39_1436 ();
 sg13g2_decap_8 FILLER_39_1443 ();
 sg13g2_decap_8 FILLER_39_1450 ();
 sg13g2_decap_8 FILLER_39_1457 ();
 sg13g2_decap_8 FILLER_39_1464 ();
 sg13g2_decap_8 FILLER_39_1471 ();
 sg13g2_decap_8 FILLER_39_1478 ();
 sg13g2_decap_8 FILLER_39_1485 ();
 sg13g2_decap_8 FILLER_39_1492 ();
 sg13g2_decap_8 FILLER_39_1499 ();
 sg13g2_decap_8 FILLER_39_1506 ();
 sg13g2_decap_8 FILLER_39_1513 ();
 sg13g2_decap_8 FILLER_39_1520 ();
 sg13g2_decap_8 FILLER_39_1527 ();
 sg13g2_decap_8 FILLER_39_1534 ();
 sg13g2_decap_8 FILLER_39_1541 ();
 sg13g2_decap_8 FILLER_39_1548 ();
 sg13g2_decap_8 FILLER_39_1555 ();
 sg13g2_decap_8 FILLER_39_1562 ();
 sg13g2_decap_8 FILLER_39_1569 ();
 sg13g2_decap_8 FILLER_39_1576 ();
 sg13g2_decap_8 FILLER_39_1583 ();
 sg13g2_decap_8 FILLER_39_1590 ();
 sg13g2_decap_8 FILLER_39_1597 ();
 sg13g2_decap_8 FILLER_39_1604 ();
 sg13g2_decap_8 FILLER_39_1611 ();
 sg13g2_decap_8 FILLER_39_1618 ();
 sg13g2_decap_8 FILLER_39_1625 ();
 sg13g2_decap_8 FILLER_39_1632 ();
 sg13g2_decap_8 FILLER_39_1639 ();
 sg13g2_decap_8 FILLER_39_1646 ();
 sg13g2_decap_8 FILLER_39_1653 ();
 sg13g2_decap_8 FILLER_39_1660 ();
 sg13g2_decap_8 FILLER_39_1667 ();
 sg13g2_decap_8 FILLER_39_1674 ();
 sg13g2_decap_8 FILLER_39_1681 ();
 sg13g2_decap_8 FILLER_39_1688 ();
 sg13g2_decap_8 FILLER_39_1695 ();
 sg13g2_decap_8 FILLER_39_1702 ();
 sg13g2_decap_8 FILLER_39_1709 ();
 sg13g2_decap_8 FILLER_39_1716 ();
 sg13g2_decap_8 FILLER_39_1723 ();
 sg13g2_decap_8 FILLER_39_1730 ();
 sg13g2_decap_8 FILLER_39_1737 ();
 sg13g2_decap_8 FILLER_39_1744 ();
 sg13g2_decap_8 FILLER_39_1751 ();
 sg13g2_decap_8 FILLER_39_1758 ();
 sg13g2_fill_2 FILLER_39_1765 ();
 sg13g2_fill_1 FILLER_39_1767 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_4 FILLER_40_177 ();
 sg13g2_fill_1 FILLER_40_211 ();
 sg13g2_fill_2 FILLER_40_231 ();
 sg13g2_fill_1 FILLER_40_233 ();
 sg13g2_fill_2 FILLER_40_243 ();
 sg13g2_fill_1 FILLER_40_245 ();
 sg13g2_fill_2 FILLER_40_272 ();
 sg13g2_fill_1 FILLER_40_274 ();
 sg13g2_decap_4 FILLER_40_289 ();
 sg13g2_fill_1 FILLER_40_293 ();
 sg13g2_fill_1 FILLER_40_304 ();
 sg13g2_fill_1 FILLER_40_367 ();
 sg13g2_decap_8 FILLER_40_376 ();
 sg13g2_fill_1 FILLER_40_391 ();
 sg13g2_fill_1 FILLER_40_397 ();
 sg13g2_fill_1 FILLER_40_414 ();
 sg13g2_decap_4 FILLER_40_426 ();
 sg13g2_decap_4 FILLER_40_435 ();
 sg13g2_fill_1 FILLER_40_439 ();
 sg13g2_fill_2 FILLER_40_475 ();
 sg13g2_fill_1 FILLER_40_477 ();
 sg13g2_fill_2 FILLER_40_490 ();
 sg13g2_fill_2 FILLER_40_526 ();
 sg13g2_fill_2 FILLER_40_565 ();
 sg13g2_fill_1 FILLER_40_567 ();
 sg13g2_fill_2 FILLER_40_576 ();
 sg13g2_fill_1 FILLER_40_599 ();
 sg13g2_fill_2 FILLER_40_653 ();
 sg13g2_fill_1 FILLER_40_655 ();
 sg13g2_fill_1 FILLER_40_681 ();
 sg13g2_decap_4 FILLER_40_719 ();
 sg13g2_fill_2 FILLER_40_723 ();
 sg13g2_fill_1 FILLER_40_729 ();
 sg13g2_fill_2 FILLER_40_733 ();
 sg13g2_fill_1 FILLER_40_768 ();
 sg13g2_fill_2 FILLER_40_784 ();
 sg13g2_fill_1 FILLER_40_786 ();
 sg13g2_fill_2 FILLER_40_832 ();
 sg13g2_fill_1 FILLER_40_834 ();
 sg13g2_decap_8 FILLER_40_861 ();
 sg13g2_decap_4 FILLER_40_868 ();
 sg13g2_fill_1 FILLER_40_872 ();
 sg13g2_decap_8 FILLER_40_881 ();
 sg13g2_fill_2 FILLER_40_888 ();
 sg13g2_fill_2 FILLER_40_897 ();
 sg13g2_fill_2 FILLER_40_911 ();
 sg13g2_fill_1 FILLER_40_913 ();
 sg13g2_decap_4 FILLER_40_920 ();
 sg13g2_fill_1 FILLER_40_924 ();
 sg13g2_decap_8 FILLER_40_1006 ();
 sg13g2_fill_1 FILLER_40_1013 ();
 sg13g2_decap_8 FILLER_40_1042 ();
 sg13g2_decap_8 FILLER_40_1049 ();
 sg13g2_decap_8 FILLER_40_1056 ();
 sg13g2_fill_2 FILLER_40_1069 ();
 sg13g2_fill_1 FILLER_40_1071 ();
 sg13g2_fill_1 FILLER_40_1096 ();
 sg13g2_decap_8 FILLER_40_1145 ();
 sg13g2_decap_8 FILLER_40_1152 ();
 sg13g2_decap_8 FILLER_40_1159 ();
 sg13g2_decap_8 FILLER_40_1166 ();
 sg13g2_decap_8 FILLER_40_1173 ();
 sg13g2_decap_8 FILLER_40_1180 ();
 sg13g2_decap_8 FILLER_40_1187 ();
 sg13g2_decap_8 FILLER_40_1194 ();
 sg13g2_decap_8 FILLER_40_1201 ();
 sg13g2_decap_8 FILLER_40_1208 ();
 sg13g2_decap_8 FILLER_40_1215 ();
 sg13g2_decap_8 FILLER_40_1222 ();
 sg13g2_decap_8 FILLER_40_1229 ();
 sg13g2_decap_8 FILLER_40_1236 ();
 sg13g2_decap_8 FILLER_40_1243 ();
 sg13g2_decap_8 FILLER_40_1250 ();
 sg13g2_decap_8 FILLER_40_1257 ();
 sg13g2_decap_8 FILLER_40_1264 ();
 sg13g2_decap_8 FILLER_40_1271 ();
 sg13g2_decap_8 FILLER_40_1278 ();
 sg13g2_decap_8 FILLER_40_1285 ();
 sg13g2_decap_8 FILLER_40_1292 ();
 sg13g2_decap_8 FILLER_40_1299 ();
 sg13g2_decap_8 FILLER_40_1306 ();
 sg13g2_decap_8 FILLER_40_1313 ();
 sg13g2_decap_8 FILLER_40_1320 ();
 sg13g2_decap_8 FILLER_40_1327 ();
 sg13g2_decap_8 FILLER_40_1334 ();
 sg13g2_decap_8 FILLER_40_1341 ();
 sg13g2_decap_8 FILLER_40_1348 ();
 sg13g2_decap_8 FILLER_40_1355 ();
 sg13g2_decap_8 FILLER_40_1362 ();
 sg13g2_decap_8 FILLER_40_1369 ();
 sg13g2_decap_8 FILLER_40_1376 ();
 sg13g2_decap_8 FILLER_40_1383 ();
 sg13g2_decap_8 FILLER_40_1390 ();
 sg13g2_decap_8 FILLER_40_1397 ();
 sg13g2_decap_8 FILLER_40_1404 ();
 sg13g2_decap_8 FILLER_40_1411 ();
 sg13g2_decap_8 FILLER_40_1418 ();
 sg13g2_decap_8 FILLER_40_1425 ();
 sg13g2_decap_8 FILLER_40_1432 ();
 sg13g2_decap_8 FILLER_40_1439 ();
 sg13g2_decap_8 FILLER_40_1446 ();
 sg13g2_decap_8 FILLER_40_1453 ();
 sg13g2_decap_8 FILLER_40_1460 ();
 sg13g2_decap_8 FILLER_40_1467 ();
 sg13g2_decap_8 FILLER_40_1474 ();
 sg13g2_decap_8 FILLER_40_1481 ();
 sg13g2_decap_8 FILLER_40_1488 ();
 sg13g2_decap_8 FILLER_40_1495 ();
 sg13g2_decap_8 FILLER_40_1502 ();
 sg13g2_decap_8 FILLER_40_1509 ();
 sg13g2_decap_8 FILLER_40_1516 ();
 sg13g2_decap_8 FILLER_40_1523 ();
 sg13g2_decap_8 FILLER_40_1530 ();
 sg13g2_decap_8 FILLER_40_1537 ();
 sg13g2_decap_8 FILLER_40_1544 ();
 sg13g2_decap_8 FILLER_40_1551 ();
 sg13g2_decap_8 FILLER_40_1558 ();
 sg13g2_decap_8 FILLER_40_1565 ();
 sg13g2_decap_8 FILLER_40_1572 ();
 sg13g2_decap_8 FILLER_40_1579 ();
 sg13g2_decap_8 FILLER_40_1586 ();
 sg13g2_decap_8 FILLER_40_1593 ();
 sg13g2_decap_8 FILLER_40_1600 ();
 sg13g2_decap_8 FILLER_40_1607 ();
 sg13g2_decap_8 FILLER_40_1614 ();
 sg13g2_decap_8 FILLER_40_1621 ();
 sg13g2_decap_8 FILLER_40_1628 ();
 sg13g2_decap_8 FILLER_40_1635 ();
 sg13g2_decap_8 FILLER_40_1642 ();
 sg13g2_decap_8 FILLER_40_1649 ();
 sg13g2_decap_8 FILLER_40_1656 ();
 sg13g2_decap_8 FILLER_40_1663 ();
 sg13g2_decap_8 FILLER_40_1670 ();
 sg13g2_decap_8 FILLER_40_1677 ();
 sg13g2_decap_8 FILLER_40_1684 ();
 sg13g2_decap_8 FILLER_40_1691 ();
 sg13g2_decap_8 FILLER_40_1698 ();
 sg13g2_decap_8 FILLER_40_1705 ();
 sg13g2_decap_8 FILLER_40_1712 ();
 sg13g2_decap_8 FILLER_40_1719 ();
 sg13g2_decap_8 FILLER_40_1726 ();
 sg13g2_decap_8 FILLER_40_1733 ();
 sg13g2_decap_8 FILLER_40_1740 ();
 sg13g2_decap_8 FILLER_40_1747 ();
 sg13g2_decap_8 FILLER_40_1754 ();
 sg13g2_decap_8 FILLER_40_1761 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_4 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_71 ();
 sg13g2_decap_8 FILLER_41_78 ();
 sg13g2_decap_8 FILLER_41_85 ();
 sg13g2_decap_4 FILLER_41_92 ();
 sg13g2_decap_8 FILLER_41_108 ();
 sg13g2_decap_8 FILLER_41_115 ();
 sg13g2_decap_8 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_137 ();
 sg13g2_decap_4 FILLER_41_144 ();
 sg13g2_fill_1 FILLER_41_148 ();
 sg13g2_fill_1 FILLER_41_158 ();
 sg13g2_decap_4 FILLER_41_162 ();
 sg13g2_fill_2 FILLER_41_166 ();
 sg13g2_decap_8 FILLER_41_176 ();
 sg13g2_decap_8 FILLER_41_183 ();
 sg13g2_fill_1 FILLER_41_190 ();
 sg13g2_fill_2 FILLER_41_268 ();
 sg13g2_fill_1 FILLER_41_270 ();
 sg13g2_fill_1 FILLER_41_276 ();
 sg13g2_decap_8 FILLER_41_281 ();
 sg13g2_decap_8 FILLER_41_288 ();
 sg13g2_fill_2 FILLER_41_295 ();
 sg13g2_fill_1 FILLER_41_297 ();
 sg13g2_fill_1 FILLER_41_306 ();
 sg13g2_decap_8 FILLER_41_312 ();
 sg13g2_decap_8 FILLER_41_319 ();
 sg13g2_decap_8 FILLER_41_326 ();
 sg13g2_decap_8 FILLER_41_333 ();
 sg13g2_fill_2 FILLER_41_340 ();
 sg13g2_decap_4 FILLER_41_346 ();
 sg13g2_fill_2 FILLER_41_350 ();
 sg13g2_fill_1 FILLER_41_355 ();
 sg13g2_fill_2 FILLER_41_366 ();
 sg13g2_decap_4 FILLER_41_381 ();
 sg13g2_fill_1 FILLER_41_385 ();
 sg13g2_decap_4 FILLER_41_399 ();
 sg13g2_fill_1 FILLER_41_403 ();
 sg13g2_decap_8 FILLER_41_435 ();
 sg13g2_decap_4 FILLER_41_442 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_4 FILLER_41_497 ();
 sg13g2_decap_4 FILLER_41_509 ();
 sg13g2_fill_2 FILLER_41_513 ();
 sg13g2_fill_1 FILLER_41_523 ();
 sg13g2_fill_2 FILLER_41_529 ();
 sg13g2_fill_1 FILLER_41_531 ();
 sg13g2_fill_2 FILLER_41_536 ();
 sg13g2_fill_1 FILLER_41_538 ();
 sg13g2_decap_8 FILLER_41_568 ();
 sg13g2_fill_2 FILLER_41_575 ();
 sg13g2_fill_1 FILLER_41_577 ();
 sg13g2_fill_2 FILLER_41_589 ();
 sg13g2_fill_2 FILLER_41_613 ();
 sg13g2_decap_8 FILLER_41_622 ();
 sg13g2_fill_2 FILLER_41_629 ();
 sg13g2_fill_2 FILLER_41_666 ();
 sg13g2_fill_1 FILLER_41_683 ();
 sg13g2_fill_1 FILLER_41_703 ();
 sg13g2_fill_1 FILLER_41_730 ();
 sg13g2_fill_2 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_795 ();
 sg13g2_decap_8 FILLER_41_802 ();
 sg13g2_decap_4 FILLER_41_809 ();
 sg13g2_fill_1 FILLER_41_813 ();
 sg13g2_fill_2 FILLER_41_837 ();
 sg13g2_decap_4 FILLER_41_848 ();
 sg13g2_fill_1 FILLER_41_852 ();
 sg13g2_fill_2 FILLER_41_861 ();
 sg13g2_fill_1 FILLER_41_863 ();
 sg13g2_fill_2 FILLER_41_870 ();
 sg13g2_fill_1 FILLER_41_892 ();
 sg13g2_decap_4 FILLER_41_903 ();
 sg13g2_fill_2 FILLER_41_917 ();
 sg13g2_fill_1 FILLER_41_919 ();
 sg13g2_fill_2 FILLER_41_953 ();
 sg13g2_fill_2 FILLER_41_966 ();
 sg13g2_decap_8 FILLER_41_986 ();
 sg13g2_fill_2 FILLER_41_993 ();
 sg13g2_fill_1 FILLER_41_995 ();
 sg13g2_decap_4 FILLER_41_1002 ();
 sg13g2_fill_2 FILLER_41_1021 ();
 sg13g2_fill_1 FILLER_41_1023 ();
 sg13g2_decap_4 FILLER_41_1060 ();
 sg13g2_fill_1 FILLER_41_1064 ();
 sg13g2_fill_1 FILLER_41_1083 ();
 sg13g2_decap_8 FILLER_41_1123 ();
 sg13g2_decap_8 FILLER_41_1130 ();
 sg13g2_decap_8 FILLER_41_1137 ();
 sg13g2_decap_8 FILLER_41_1144 ();
 sg13g2_decap_8 FILLER_41_1151 ();
 sg13g2_decap_8 FILLER_41_1158 ();
 sg13g2_decap_8 FILLER_41_1165 ();
 sg13g2_decap_8 FILLER_41_1172 ();
 sg13g2_decap_8 FILLER_41_1179 ();
 sg13g2_decap_8 FILLER_41_1186 ();
 sg13g2_decap_8 FILLER_41_1193 ();
 sg13g2_decap_8 FILLER_41_1200 ();
 sg13g2_decap_8 FILLER_41_1207 ();
 sg13g2_decap_8 FILLER_41_1214 ();
 sg13g2_decap_8 FILLER_41_1221 ();
 sg13g2_decap_8 FILLER_41_1228 ();
 sg13g2_decap_8 FILLER_41_1235 ();
 sg13g2_decap_8 FILLER_41_1242 ();
 sg13g2_decap_8 FILLER_41_1249 ();
 sg13g2_decap_8 FILLER_41_1256 ();
 sg13g2_decap_8 FILLER_41_1263 ();
 sg13g2_decap_8 FILLER_41_1270 ();
 sg13g2_decap_8 FILLER_41_1277 ();
 sg13g2_decap_8 FILLER_41_1284 ();
 sg13g2_decap_8 FILLER_41_1291 ();
 sg13g2_decap_8 FILLER_41_1298 ();
 sg13g2_decap_8 FILLER_41_1305 ();
 sg13g2_decap_8 FILLER_41_1312 ();
 sg13g2_decap_8 FILLER_41_1319 ();
 sg13g2_decap_8 FILLER_41_1326 ();
 sg13g2_decap_8 FILLER_41_1333 ();
 sg13g2_decap_8 FILLER_41_1340 ();
 sg13g2_decap_8 FILLER_41_1347 ();
 sg13g2_decap_8 FILLER_41_1354 ();
 sg13g2_decap_8 FILLER_41_1361 ();
 sg13g2_decap_8 FILLER_41_1368 ();
 sg13g2_decap_8 FILLER_41_1375 ();
 sg13g2_decap_8 FILLER_41_1382 ();
 sg13g2_decap_8 FILLER_41_1389 ();
 sg13g2_decap_8 FILLER_41_1396 ();
 sg13g2_decap_8 FILLER_41_1403 ();
 sg13g2_decap_8 FILLER_41_1410 ();
 sg13g2_decap_8 FILLER_41_1417 ();
 sg13g2_decap_8 FILLER_41_1424 ();
 sg13g2_decap_8 FILLER_41_1431 ();
 sg13g2_decap_8 FILLER_41_1438 ();
 sg13g2_decap_8 FILLER_41_1445 ();
 sg13g2_decap_8 FILLER_41_1452 ();
 sg13g2_decap_8 FILLER_41_1459 ();
 sg13g2_decap_8 FILLER_41_1466 ();
 sg13g2_decap_8 FILLER_41_1473 ();
 sg13g2_decap_8 FILLER_41_1480 ();
 sg13g2_decap_8 FILLER_41_1487 ();
 sg13g2_decap_8 FILLER_41_1494 ();
 sg13g2_decap_8 FILLER_41_1501 ();
 sg13g2_decap_8 FILLER_41_1508 ();
 sg13g2_decap_8 FILLER_41_1515 ();
 sg13g2_decap_8 FILLER_41_1522 ();
 sg13g2_decap_8 FILLER_41_1529 ();
 sg13g2_decap_8 FILLER_41_1536 ();
 sg13g2_decap_8 FILLER_41_1543 ();
 sg13g2_decap_8 FILLER_41_1550 ();
 sg13g2_decap_8 FILLER_41_1557 ();
 sg13g2_decap_8 FILLER_41_1564 ();
 sg13g2_decap_8 FILLER_41_1571 ();
 sg13g2_decap_8 FILLER_41_1578 ();
 sg13g2_decap_8 FILLER_41_1585 ();
 sg13g2_decap_8 FILLER_41_1592 ();
 sg13g2_decap_8 FILLER_41_1599 ();
 sg13g2_decap_8 FILLER_41_1606 ();
 sg13g2_decap_8 FILLER_41_1613 ();
 sg13g2_decap_8 FILLER_41_1620 ();
 sg13g2_decap_8 FILLER_41_1627 ();
 sg13g2_decap_8 FILLER_41_1634 ();
 sg13g2_decap_8 FILLER_41_1641 ();
 sg13g2_decap_8 FILLER_41_1648 ();
 sg13g2_decap_8 FILLER_41_1655 ();
 sg13g2_decap_8 FILLER_41_1662 ();
 sg13g2_decap_8 FILLER_41_1669 ();
 sg13g2_decap_8 FILLER_41_1676 ();
 sg13g2_decap_8 FILLER_41_1683 ();
 sg13g2_decap_8 FILLER_41_1690 ();
 sg13g2_decap_8 FILLER_41_1697 ();
 sg13g2_decap_8 FILLER_41_1704 ();
 sg13g2_decap_8 FILLER_41_1711 ();
 sg13g2_decap_8 FILLER_41_1718 ();
 sg13g2_decap_8 FILLER_41_1725 ();
 sg13g2_decap_8 FILLER_41_1732 ();
 sg13g2_decap_8 FILLER_41_1739 ();
 sg13g2_decap_8 FILLER_41_1746 ();
 sg13g2_decap_8 FILLER_41_1753 ();
 sg13g2_decap_8 FILLER_41_1760 ();
 sg13g2_fill_1 FILLER_41_1767 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_fill_2 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_76 ();
 sg13g2_decap_8 FILLER_42_83 ();
 sg13g2_decap_4 FILLER_42_90 ();
 sg13g2_fill_1 FILLER_42_94 ();
 sg13g2_decap_4 FILLER_42_127 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_fill_1 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_198 ();
 sg13g2_fill_2 FILLER_42_235 ();
 sg13g2_fill_1 FILLER_42_237 ();
 sg13g2_fill_1 FILLER_42_242 ();
 sg13g2_decap_8 FILLER_42_253 ();
 sg13g2_fill_1 FILLER_42_260 ();
 sg13g2_fill_2 FILLER_42_291 ();
 sg13g2_fill_1 FILLER_42_311 ();
 sg13g2_fill_2 FILLER_42_373 ();
 sg13g2_fill_1 FILLER_42_375 ();
 sg13g2_decap_4 FILLER_42_379 ();
 sg13g2_decap_8 FILLER_42_409 ();
 sg13g2_fill_1 FILLER_42_416 ();
 sg13g2_decap_8 FILLER_42_448 ();
 sg13g2_decap_8 FILLER_42_455 ();
 sg13g2_fill_2 FILLER_42_462 ();
 sg13g2_fill_1 FILLER_42_464 ();
 sg13g2_fill_1 FILLER_42_473 ();
 sg13g2_decap_4 FILLER_42_486 ();
 sg13g2_fill_2 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_500 ();
 sg13g2_fill_1 FILLER_42_507 ();
 sg13g2_fill_1 FILLER_42_542 ();
 sg13g2_decap_4 FILLER_42_587 ();
 sg13g2_fill_2 FILLER_42_607 ();
 sg13g2_fill_1 FILLER_42_609 ();
 sg13g2_fill_2 FILLER_42_615 ();
 sg13g2_decap_4 FILLER_42_644 ();
 sg13g2_fill_2 FILLER_42_674 ();
 sg13g2_fill_1 FILLER_42_676 ();
 sg13g2_fill_1 FILLER_42_716 ();
 sg13g2_fill_1 FILLER_42_734 ();
 sg13g2_fill_2 FILLER_42_770 ();
 sg13g2_fill_2 FILLER_42_815 ();
 sg13g2_fill_1 FILLER_42_817 ();
 sg13g2_fill_2 FILLER_42_866 ();
 sg13g2_fill_1 FILLER_42_878 ();
 sg13g2_fill_2 FILLER_42_906 ();
 sg13g2_fill_1 FILLER_42_908 ();
 sg13g2_fill_1 FILLER_42_945 ();
 sg13g2_decap_8 FILLER_42_960 ();
 sg13g2_decap_4 FILLER_42_967 ();
 sg13g2_fill_2 FILLER_42_991 ();
 sg13g2_fill_1 FILLER_42_993 ();
 sg13g2_fill_1 FILLER_42_1022 ();
 sg13g2_decap_8 FILLER_42_1054 ();
 sg13g2_fill_2 FILLER_42_1061 ();
 sg13g2_fill_1 FILLER_42_1086 ();
 sg13g2_decap_8 FILLER_42_1113 ();
 sg13g2_decap_8 FILLER_42_1120 ();
 sg13g2_decap_8 FILLER_42_1127 ();
 sg13g2_decap_8 FILLER_42_1134 ();
 sg13g2_decap_8 FILLER_42_1141 ();
 sg13g2_decap_8 FILLER_42_1148 ();
 sg13g2_decap_8 FILLER_42_1155 ();
 sg13g2_decap_8 FILLER_42_1162 ();
 sg13g2_decap_8 FILLER_42_1169 ();
 sg13g2_decap_8 FILLER_42_1176 ();
 sg13g2_decap_8 FILLER_42_1183 ();
 sg13g2_decap_8 FILLER_42_1190 ();
 sg13g2_decap_8 FILLER_42_1197 ();
 sg13g2_decap_8 FILLER_42_1204 ();
 sg13g2_decap_8 FILLER_42_1211 ();
 sg13g2_decap_8 FILLER_42_1218 ();
 sg13g2_decap_8 FILLER_42_1225 ();
 sg13g2_decap_8 FILLER_42_1232 ();
 sg13g2_decap_8 FILLER_42_1239 ();
 sg13g2_decap_8 FILLER_42_1246 ();
 sg13g2_decap_8 FILLER_42_1253 ();
 sg13g2_decap_8 FILLER_42_1260 ();
 sg13g2_decap_8 FILLER_42_1267 ();
 sg13g2_decap_8 FILLER_42_1274 ();
 sg13g2_decap_8 FILLER_42_1281 ();
 sg13g2_decap_8 FILLER_42_1288 ();
 sg13g2_decap_8 FILLER_42_1295 ();
 sg13g2_decap_8 FILLER_42_1302 ();
 sg13g2_decap_8 FILLER_42_1309 ();
 sg13g2_decap_8 FILLER_42_1316 ();
 sg13g2_decap_8 FILLER_42_1323 ();
 sg13g2_decap_8 FILLER_42_1330 ();
 sg13g2_decap_8 FILLER_42_1337 ();
 sg13g2_decap_8 FILLER_42_1344 ();
 sg13g2_decap_8 FILLER_42_1351 ();
 sg13g2_decap_8 FILLER_42_1358 ();
 sg13g2_decap_8 FILLER_42_1365 ();
 sg13g2_decap_8 FILLER_42_1372 ();
 sg13g2_decap_8 FILLER_42_1379 ();
 sg13g2_decap_8 FILLER_42_1386 ();
 sg13g2_decap_8 FILLER_42_1393 ();
 sg13g2_decap_8 FILLER_42_1400 ();
 sg13g2_decap_8 FILLER_42_1407 ();
 sg13g2_decap_8 FILLER_42_1414 ();
 sg13g2_decap_8 FILLER_42_1421 ();
 sg13g2_decap_8 FILLER_42_1428 ();
 sg13g2_decap_8 FILLER_42_1435 ();
 sg13g2_decap_8 FILLER_42_1442 ();
 sg13g2_decap_8 FILLER_42_1449 ();
 sg13g2_decap_8 FILLER_42_1456 ();
 sg13g2_decap_8 FILLER_42_1463 ();
 sg13g2_decap_8 FILLER_42_1470 ();
 sg13g2_decap_8 FILLER_42_1477 ();
 sg13g2_decap_8 FILLER_42_1484 ();
 sg13g2_decap_8 FILLER_42_1491 ();
 sg13g2_decap_8 FILLER_42_1498 ();
 sg13g2_decap_8 FILLER_42_1505 ();
 sg13g2_decap_8 FILLER_42_1512 ();
 sg13g2_decap_8 FILLER_42_1519 ();
 sg13g2_decap_8 FILLER_42_1526 ();
 sg13g2_decap_8 FILLER_42_1533 ();
 sg13g2_decap_8 FILLER_42_1540 ();
 sg13g2_decap_8 FILLER_42_1547 ();
 sg13g2_decap_8 FILLER_42_1554 ();
 sg13g2_decap_8 FILLER_42_1561 ();
 sg13g2_decap_8 FILLER_42_1568 ();
 sg13g2_decap_8 FILLER_42_1575 ();
 sg13g2_decap_8 FILLER_42_1582 ();
 sg13g2_decap_8 FILLER_42_1589 ();
 sg13g2_decap_8 FILLER_42_1596 ();
 sg13g2_decap_8 FILLER_42_1603 ();
 sg13g2_decap_8 FILLER_42_1610 ();
 sg13g2_decap_8 FILLER_42_1617 ();
 sg13g2_decap_8 FILLER_42_1624 ();
 sg13g2_decap_8 FILLER_42_1631 ();
 sg13g2_decap_8 FILLER_42_1638 ();
 sg13g2_decap_8 FILLER_42_1645 ();
 sg13g2_decap_8 FILLER_42_1652 ();
 sg13g2_decap_8 FILLER_42_1659 ();
 sg13g2_decap_8 FILLER_42_1666 ();
 sg13g2_decap_8 FILLER_42_1673 ();
 sg13g2_decap_8 FILLER_42_1680 ();
 sg13g2_decap_8 FILLER_42_1687 ();
 sg13g2_decap_8 FILLER_42_1694 ();
 sg13g2_decap_8 FILLER_42_1701 ();
 sg13g2_decap_8 FILLER_42_1708 ();
 sg13g2_decap_8 FILLER_42_1715 ();
 sg13g2_decap_8 FILLER_42_1722 ();
 sg13g2_decap_8 FILLER_42_1729 ();
 sg13g2_decap_8 FILLER_42_1736 ();
 sg13g2_decap_8 FILLER_42_1743 ();
 sg13g2_decap_8 FILLER_42_1750 ();
 sg13g2_decap_8 FILLER_42_1757 ();
 sg13g2_decap_4 FILLER_42_1764 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_fill_1 FILLER_43_72 ();
 sg13g2_fill_2 FILLER_43_103 ();
 sg13g2_fill_1 FILLER_43_105 ();
 sg13g2_fill_2 FILLER_43_132 ();
 sg13g2_fill_1 FILLER_43_134 ();
 sg13g2_fill_2 FILLER_43_150 ();
 sg13g2_fill_1 FILLER_43_152 ();
 sg13g2_decap_8 FILLER_43_193 ();
 sg13g2_fill_2 FILLER_43_219 ();
 sg13g2_fill_1 FILLER_43_330 ();
 sg13g2_fill_2 FILLER_43_341 ();
 sg13g2_decap_4 FILLER_43_362 ();
 sg13g2_fill_2 FILLER_43_396 ();
 sg13g2_fill_1 FILLER_43_398 ();
 sg13g2_fill_2 FILLER_43_408 ();
 sg13g2_fill_1 FILLER_43_410 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_fill_2 FILLER_43_427 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_fill_2 FILLER_43_439 ();
 sg13g2_fill_2 FILLER_43_449 ();
 sg13g2_decap_4 FILLER_43_464 ();
 sg13g2_fill_1 FILLER_43_468 ();
 sg13g2_decap_8 FILLER_43_477 ();
 sg13g2_fill_1 FILLER_43_484 ();
 sg13g2_fill_1 FILLER_43_504 ();
 sg13g2_fill_2 FILLER_43_518 ();
 sg13g2_fill_1 FILLER_43_520 ();
 sg13g2_fill_1 FILLER_43_562 ();
 sg13g2_fill_2 FILLER_43_589 ();
 sg13g2_fill_2 FILLER_43_599 ();
 sg13g2_fill_1 FILLER_43_601 ();
 sg13g2_decap_8 FILLER_43_638 ();
 sg13g2_fill_1 FILLER_43_645 ();
 sg13g2_fill_1 FILLER_43_659 ();
 sg13g2_fill_2 FILLER_43_680 ();
 sg13g2_fill_2 FILLER_43_717 ();
 sg13g2_fill_1 FILLER_43_719 ();
 sg13g2_fill_2 FILLER_43_755 ();
 sg13g2_fill_1 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_801 ();
 sg13g2_decap_4 FILLER_43_808 ();
 sg13g2_fill_1 FILLER_43_812 ();
 sg13g2_fill_2 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_decap_4 FILLER_43_845 ();
 sg13g2_fill_1 FILLER_43_849 ();
 sg13g2_fill_1 FILLER_43_876 ();
 sg13g2_fill_2 FILLER_43_884 ();
 sg13g2_fill_1 FILLER_43_886 ();
 sg13g2_fill_1 FILLER_43_898 ();
 sg13g2_fill_2 FILLER_43_907 ();
 sg13g2_decap_4 FILLER_43_917 ();
 sg13g2_fill_2 FILLER_43_956 ();
 sg13g2_fill_2 FILLER_43_981 ();
 sg13g2_fill_1 FILLER_43_998 ();
 sg13g2_decap_4 FILLER_43_1004 ();
 sg13g2_fill_1 FILLER_43_1008 ();
 sg13g2_fill_1 FILLER_43_1027 ();
 sg13g2_fill_2 FILLER_43_1050 ();
 sg13g2_fill_2 FILLER_43_1066 ();
 sg13g2_fill_1 FILLER_43_1068 ();
 sg13g2_decap_8 FILLER_43_1106 ();
 sg13g2_decap_8 FILLER_43_1113 ();
 sg13g2_decap_8 FILLER_43_1120 ();
 sg13g2_decap_8 FILLER_43_1127 ();
 sg13g2_decap_8 FILLER_43_1134 ();
 sg13g2_decap_8 FILLER_43_1141 ();
 sg13g2_decap_8 FILLER_43_1148 ();
 sg13g2_decap_8 FILLER_43_1155 ();
 sg13g2_decap_8 FILLER_43_1162 ();
 sg13g2_decap_8 FILLER_43_1169 ();
 sg13g2_decap_8 FILLER_43_1176 ();
 sg13g2_decap_8 FILLER_43_1183 ();
 sg13g2_decap_8 FILLER_43_1190 ();
 sg13g2_decap_8 FILLER_43_1197 ();
 sg13g2_decap_8 FILLER_43_1204 ();
 sg13g2_decap_8 FILLER_43_1211 ();
 sg13g2_decap_8 FILLER_43_1218 ();
 sg13g2_decap_8 FILLER_43_1225 ();
 sg13g2_decap_8 FILLER_43_1232 ();
 sg13g2_decap_8 FILLER_43_1239 ();
 sg13g2_decap_8 FILLER_43_1246 ();
 sg13g2_decap_8 FILLER_43_1253 ();
 sg13g2_decap_8 FILLER_43_1260 ();
 sg13g2_decap_8 FILLER_43_1267 ();
 sg13g2_decap_8 FILLER_43_1274 ();
 sg13g2_decap_8 FILLER_43_1281 ();
 sg13g2_decap_8 FILLER_43_1288 ();
 sg13g2_decap_8 FILLER_43_1295 ();
 sg13g2_decap_8 FILLER_43_1302 ();
 sg13g2_decap_8 FILLER_43_1309 ();
 sg13g2_decap_8 FILLER_43_1316 ();
 sg13g2_decap_8 FILLER_43_1323 ();
 sg13g2_decap_8 FILLER_43_1330 ();
 sg13g2_decap_8 FILLER_43_1337 ();
 sg13g2_decap_8 FILLER_43_1344 ();
 sg13g2_decap_8 FILLER_43_1351 ();
 sg13g2_decap_8 FILLER_43_1358 ();
 sg13g2_decap_8 FILLER_43_1365 ();
 sg13g2_decap_8 FILLER_43_1372 ();
 sg13g2_decap_8 FILLER_43_1379 ();
 sg13g2_decap_8 FILLER_43_1386 ();
 sg13g2_decap_8 FILLER_43_1393 ();
 sg13g2_decap_8 FILLER_43_1400 ();
 sg13g2_decap_8 FILLER_43_1407 ();
 sg13g2_decap_8 FILLER_43_1414 ();
 sg13g2_decap_8 FILLER_43_1421 ();
 sg13g2_decap_8 FILLER_43_1428 ();
 sg13g2_decap_8 FILLER_43_1435 ();
 sg13g2_decap_8 FILLER_43_1442 ();
 sg13g2_decap_8 FILLER_43_1449 ();
 sg13g2_decap_8 FILLER_43_1456 ();
 sg13g2_decap_8 FILLER_43_1463 ();
 sg13g2_decap_8 FILLER_43_1470 ();
 sg13g2_decap_8 FILLER_43_1477 ();
 sg13g2_decap_8 FILLER_43_1484 ();
 sg13g2_decap_8 FILLER_43_1491 ();
 sg13g2_decap_8 FILLER_43_1498 ();
 sg13g2_decap_8 FILLER_43_1505 ();
 sg13g2_decap_8 FILLER_43_1512 ();
 sg13g2_decap_8 FILLER_43_1519 ();
 sg13g2_decap_8 FILLER_43_1526 ();
 sg13g2_decap_8 FILLER_43_1533 ();
 sg13g2_decap_8 FILLER_43_1540 ();
 sg13g2_decap_8 FILLER_43_1547 ();
 sg13g2_decap_8 FILLER_43_1554 ();
 sg13g2_decap_8 FILLER_43_1561 ();
 sg13g2_decap_8 FILLER_43_1568 ();
 sg13g2_decap_8 FILLER_43_1575 ();
 sg13g2_decap_8 FILLER_43_1582 ();
 sg13g2_decap_8 FILLER_43_1589 ();
 sg13g2_decap_8 FILLER_43_1596 ();
 sg13g2_decap_8 FILLER_43_1603 ();
 sg13g2_decap_8 FILLER_43_1610 ();
 sg13g2_decap_8 FILLER_43_1617 ();
 sg13g2_decap_8 FILLER_43_1624 ();
 sg13g2_decap_8 FILLER_43_1631 ();
 sg13g2_decap_8 FILLER_43_1638 ();
 sg13g2_decap_8 FILLER_43_1645 ();
 sg13g2_decap_8 FILLER_43_1652 ();
 sg13g2_decap_8 FILLER_43_1659 ();
 sg13g2_decap_8 FILLER_43_1666 ();
 sg13g2_decap_8 FILLER_43_1673 ();
 sg13g2_decap_8 FILLER_43_1680 ();
 sg13g2_decap_8 FILLER_43_1687 ();
 sg13g2_decap_8 FILLER_43_1694 ();
 sg13g2_decap_8 FILLER_43_1701 ();
 sg13g2_decap_8 FILLER_43_1708 ();
 sg13g2_decap_8 FILLER_43_1715 ();
 sg13g2_decap_8 FILLER_43_1722 ();
 sg13g2_decap_8 FILLER_43_1729 ();
 sg13g2_decap_8 FILLER_43_1736 ();
 sg13g2_decap_8 FILLER_43_1743 ();
 sg13g2_decap_8 FILLER_43_1750 ();
 sg13g2_decap_8 FILLER_43_1757 ();
 sg13g2_decap_4 FILLER_43_1764 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_fill_2 FILLER_44_35 ();
 sg13g2_fill_2 FILLER_44_66 ();
 sg13g2_fill_2 FILLER_44_77 ();
 sg13g2_fill_2 FILLER_44_106 ();
 sg13g2_fill_1 FILLER_44_125 ();
 sg13g2_fill_1 FILLER_44_153 ();
 sg13g2_fill_2 FILLER_44_217 ();
 sg13g2_fill_2 FILLER_44_243 ();
 sg13g2_fill_1 FILLER_44_303 ();
 sg13g2_fill_1 FILLER_44_314 ();
 sg13g2_fill_2 FILLER_44_320 ();
 sg13g2_fill_1 FILLER_44_325 ();
 sg13g2_fill_1 FILLER_44_339 ();
 sg13g2_fill_1 FILLER_44_345 ();
 sg13g2_fill_2 FILLER_44_352 ();
 sg13g2_fill_1 FILLER_44_379 ();
 sg13g2_fill_1 FILLER_44_453 ();
 sg13g2_decap_8 FILLER_44_485 ();
 sg13g2_fill_1 FILLER_44_492 ();
 sg13g2_decap_8 FILLER_44_498 ();
 sg13g2_fill_2 FILLER_44_505 ();
 sg13g2_fill_1 FILLER_44_507 ();
 sg13g2_decap_8 FILLER_44_537 ();
 sg13g2_fill_2 FILLER_44_544 ();
 sg13g2_fill_1 FILLER_44_546 ();
 sg13g2_fill_2 FILLER_44_555 ();
 sg13g2_fill_1 FILLER_44_557 ();
 sg13g2_fill_2 FILLER_44_572 ();
 sg13g2_decap_8 FILLER_44_600 ();
 sg13g2_decap_8 FILLER_44_615 ();
 sg13g2_decap_4 FILLER_44_622 ();
 sg13g2_fill_2 FILLER_44_626 ();
 sg13g2_fill_1 FILLER_44_692 ();
 sg13g2_fill_2 FILLER_44_734 ();
 sg13g2_fill_1 FILLER_44_736 ();
 sg13g2_decap_4 FILLER_44_756 ();
 sg13g2_fill_1 FILLER_44_760 ();
 sg13g2_fill_1 FILLER_44_787 ();
 sg13g2_fill_2 FILLER_44_793 ();
 sg13g2_decap_4 FILLER_44_800 ();
 sg13g2_fill_2 FILLER_44_804 ();
 sg13g2_fill_2 FILLER_44_814 ();
 sg13g2_fill_2 FILLER_44_821 ();
 sg13g2_fill_1 FILLER_44_823 ();
 sg13g2_decap_4 FILLER_44_837 ();
 sg13g2_fill_2 FILLER_44_841 ();
 sg13g2_fill_2 FILLER_44_863 ();
 sg13g2_fill_1 FILLER_44_865 ();
 sg13g2_decap_8 FILLER_44_885 ();
 sg13g2_decap_4 FILLER_44_901 ();
 sg13g2_fill_2 FILLER_44_905 ();
 sg13g2_decap_8 FILLER_44_920 ();
 sg13g2_decap_8 FILLER_44_927 ();
 sg13g2_decap_4 FILLER_44_934 ();
 sg13g2_decap_8 FILLER_44_995 ();
 sg13g2_fill_2 FILLER_44_1002 ();
 sg13g2_fill_1 FILLER_44_1004 ();
 sg13g2_decap_4 FILLER_44_1080 ();
 sg13g2_fill_1 FILLER_44_1084 ();
 sg13g2_fill_2 FILLER_44_1098 ();
 sg13g2_decap_8 FILLER_44_1109 ();
 sg13g2_decap_8 FILLER_44_1116 ();
 sg13g2_decap_8 FILLER_44_1123 ();
 sg13g2_decap_8 FILLER_44_1130 ();
 sg13g2_decap_8 FILLER_44_1137 ();
 sg13g2_decap_8 FILLER_44_1144 ();
 sg13g2_decap_8 FILLER_44_1151 ();
 sg13g2_decap_8 FILLER_44_1158 ();
 sg13g2_decap_8 FILLER_44_1165 ();
 sg13g2_decap_8 FILLER_44_1172 ();
 sg13g2_decap_8 FILLER_44_1179 ();
 sg13g2_decap_8 FILLER_44_1186 ();
 sg13g2_decap_8 FILLER_44_1193 ();
 sg13g2_decap_8 FILLER_44_1200 ();
 sg13g2_decap_8 FILLER_44_1207 ();
 sg13g2_decap_8 FILLER_44_1214 ();
 sg13g2_decap_8 FILLER_44_1221 ();
 sg13g2_decap_8 FILLER_44_1228 ();
 sg13g2_decap_8 FILLER_44_1235 ();
 sg13g2_decap_8 FILLER_44_1242 ();
 sg13g2_decap_8 FILLER_44_1249 ();
 sg13g2_decap_8 FILLER_44_1256 ();
 sg13g2_decap_8 FILLER_44_1263 ();
 sg13g2_decap_8 FILLER_44_1270 ();
 sg13g2_decap_8 FILLER_44_1277 ();
 sg13g2_decap_8 FILLER_44_1284 ();
 sg13g2_decap_8 FILLER_44_1291 ();
 sg13g2_decap_8 FILLER_44_1298 ();
 sg13g2_decap_8 FILLER_44_1305 ();
 sg13g2_decap_8 FILLER_44_1312 ();
 sg13g2_decap_8 FILLER_44_1319 ();
 sg13g2_decap_8 FILLER_44_1326 ();
 sg13g2_decap_8 FILLER_44_1333 ();
 sg13g2_decap_8 FILLER_44_1340 ();
 sg13g2_decap_8 FILLER_44_1347 ();
 sg13g2_decap_8 FILLER_44_1354 ();
 sg13g2_decap_8 FILLER_44_1361 ();
 sg13g2_decap_8 FILLER_44_1368 ();
 sg13g2_decap_8 FILLER_44_1375 ();
 sg13g2_decap_8 FILLER_44_1382 ();
 sg13g2_decap_8 FILLER_44_1389 ();
 sg13g2_decap_8 FILLER_44_1396 ();
 sg13g2_decap_8 FILLER_44_1403 ();
 sg13g2_decap_8 FILLER_44_1410 ();
 sg13g2_decap_8 FILLER_44_1417 ();
 sg13g2_decap_8 FILLER_44_1424 ();
 sg13g2_decap_8 FILLER_44_1431 ();
 sg13g2_decap_8 FILLER_44_1438 ();
 sg13g2_decap_8 FILLER_44_1445 ();
 sg13g2_decap_8 FILLER_44_1452 ();
 sg13g2_decap_8 FILLER_44_1459 ();
 sg13g2_decap_8 FILLER_44_1466 ();
 sg13g2_decap_8 FILLER_44_1473 ();
 sg13g2_decap_8 FILLER_44_1480 ();
 sg13g2_decap_8 FILLER_44_1487 ();
 sg13g2_decap_8 FILLER_44_1494 ();
 sg13g2_decap_8 FILLER_44_1501 ();
 sg13g2_decap_8 FILLER_44_1508 ();
 sg13g2_decap_8 FILLER_44_1515 ();
 sg13g2_decap_8 FILLER_44_1522 ();
 sg13g2_decap_8 FILLER_44_1529 ();
 sg13g2_decap_8 FILLER_44_1536 ();
 sg13g2_decap_8 FILLER_44_1543 ();
 sg13g2_decap_8 FILLER_44_1550 ();
 sg13g2_decap_8 FILLER_44_1557 ();
 sg13g2_decap_8 FILLER_44_1564 ();
 sg13g2_decap_8 FILLER_44_1571 ();
 sg13g2_decap_8 FILLER_44_1578 ();
 sg13g2_decap_8 FILLER_44_1585 ();
 sg13g2_decap_8 FILLER_44_1592 ();
 sg13g2_decap_8 FILLER_44_1599 ();
 sg13g2_decap_8 FILLER_44_1606 ();
 sg13g2_decap_8 FILLER_44_1613 ();
 sg13g2_decap_8 FILLER_44_1620 ();
 sg13g2_decap_8 FILLER_44_1627 ();
 sg13g2_decap_8 FILLER_44_1634 ();
 sg13g2_decap_8 FILLER_44_1641 ();
 sg13g2_decap_8 FILLER_44_1648 ();
 sg13g2_decap_8 FILLER_44_1655 ();
 sg13g2_decap_8 FILLER_44_1662 ();
 sg13g2_decap_8 FILLER_44_1669 ();
 sg13g2_decap_8 FILLER_44_1676 ();
 sg13g2_decap_8 FILLER_44_1683 ();
 sg13g2_decap_8 FILLER_44_1690 ();
 sg13g2_decap_8 FILLER_44_1697 ();
 sg13g2_decap_8 FILLER_44_1704 ();
 sg13g2_decap_8 FILLER_44_1711 ();
 sg13g2_decap_8 FILLER_44_1718 ();
 sg13g2_decap_8 FILLER_44_1725 ();
 sg13g2_decap_8 FILLER_44_1732 ();
 sg13g2_decap_8 FILLER_44_1739 ();
 sg13g2_decap_8 FILLER_44_1746 ();
 sg13g2_decap_8 FILLER_44_1753 ();
 sg13g2_decap_8 FILLER_44_1760 ();
 sg13g2_fill_1 FILLER_44_1767 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_4 FILLER_45_35 ();
 sg13g2_fill_2 FILLER_45_76 ();
 sg13g2_fill_2 FILLER_45_87 ();
 sg13g2_fill_1 FILLER_45_99 ();
 sg13g2_fill_2 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_198 ();
 sg13g2_fill_1 FILLER_45_208 ();
 sg13g2_fill_2 FILLER_45_215 ();
 sg13g2_fill_1 FILLER_45_222 ();
 sg13g2_fill_1 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_249 ();
 sg13g2_decap_8 FILLER_45_314 ();
 sg13g2_fill_2 FILLER_45_326 ();
 sg13g2_fill_1 FILLER_45_345 ();
 sg13g2_fill_1 FILLER_45_355 ();
 sg13g2_fill_1 FILLER_45_388 ();
 sg13g2_fill_1 FILLER_45_394 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_fill_2 FILLER_45_412 ();
 sg13g2_decap_4 FILLER_45_417 ();
 sg13g2_decap_4 FILLER_45_438 ();
 sg13g2_fill_2 FILLER_45_442 ();
 sg13g2_decap_8 FILLER_45_449 ();
 sg13g2_decap_8 FILLER_45_472 ();
 sg13g2_fill_2 FILLER_45_479 ();
 sg13g2_fill_2 FILLER_45_486 ();
 sg13g2_decap_8 FILLER_45_496 ();
 sg13g2_fill_1 FILLER_45_503 ();
 sg13g2_fill_1 FILLER_45_517 ();
 sg13g2_decap_4 FILLER_45_540 ();
 sg13g2_decap_4 FILLER_45_552 ();
 sg13g2_fill_2 FILLER_45_556 ();
 sg13g2_fill_2 FILLER_45_587 ();
 sg13g2_fill_1 FILLER_45_589 ();
 sg13g2_fill_1 FILLER_45_630 ();
 sg13g2_fill_1 FILLER_45_657 ();
 sg13g2_fill_2 FILLER_45_663 ();
 sg13g2_fill_2 FILLER_45_675 ();
 sg13g2_fill_1 FILLER_45_681 ();
 sg13g2_fill_1 FILLER_45_697 ();
 sg13g2_decap_4 FILLER_45_746 ();
 sg13g2_fill_2 FILLER_45_750 ();
 sg13g2_fill_2 FILLER_45_766 ();
 sg13g2_decap_8 FILLER_45_771 ();
 sg13g2_decap_4 FILLER_45_778 ();
 sg13g2_fill_1 FILLER_45_782 ();
 sg13g2_decap_4 FILLER_45_809 ();
 sg13g2_fill_2 FILLER_45_824 ();
 sg13g2_fill_1 FILLER_45_866 ();
 sg13g2_decap_4 FILLER_45_871 ();
 sg13g2_fill_2 FILLER_45_901 ();
 sg13g2_fill_1 FILLER_45_903 ();
 sg13g2_fill_1 FILLER_45_943 ();
 sg13g2_fill_1 FILLER_45_974 ();
 sg13g2_decap_4 FILLER_45_1018 ();
 sg13g2_decap_8 FILLER_45_1079 ();
 sg13g2_decap_8 FILLER_45_1086 ();
 sg13g2_decap_4 FILLER_45_1093 ();
 sg13g2_fill_1 FILLER_45_1097 ();
 sg13g2_decap_8 FILLER_45_1101 ();
 sg13g2_decap_8 FILLER_45_1108 ();
 sg13g2_decap_8 FILLER_45_1115 ();
 sg13g2_decap_8 FILLER_45_1122 ();
 sg13g2_decap_8 FILLER_45_1129 ();
 sg13g2_decap_8 FILLER_45_1136 ();
 sg13g2_decap_8 FILLER_45_1143 ();
 sg13g2_decap_8 FILLER_45_1150 ();
 sg13g2_decap_8 FILLER_45_1157 ();
 sg13g2_decap_8 FILLER_45_1164 ();
 sg13g2_decap_8 FILLER_45_1171 ();
 sg13g2_decap_8 FILLER_45_1178 ();
 sg13g2_decap_8 FILLER_45_1185 ();
 sg13g2_decap_8 FILLER_45_1192 ();
 sg13g2_decap_8 FILLER_45_1199 ();
 sg13g2_decap_8 FILLER_45_1206 ();
 sg13g2_decap_8 FILLER_45_1213 ();
 sg13g2_decap_8 FILLER_45_1220 ();
 sg13g2_decap_8 FILLER_45_1227 ();
 sg13g2_decap_8 FILLER_45_1234 ();
 sg13g2_decap_8 FILLER_45_1241 ();
 sg13g2_decap_8 FILLER_45_1248 ();
 sg13g2_decap_8 FILLER_45_1255 ();
 sg13g2_decap_8 FILLER_45_1262 ();
 sg13g2_decap_8 FILLER_45_1269 ();
 sg13g2_decap_8 FILLER_45_1276 ();
 sg13g2_decap_8 FILLER_45_1283 ();
 sg13g2_decap_8 FILLER_45_1290 ();
 sg13g2_decap_8 FILLER_45_1297 ();
 sg13g2_decap_8 FILLER_45_1304 ();
 sg13g2_decap_8 FILLER_45_1311 ();
 sg13g2_decap_8 FILLER_45_1318 ();
 sg13g2_decap_8 FILLER_45_1325 ();
 sg13g2_decap_8 FILLER_45_1332 ();
 sg13g2_decap_8 FILLER_45_1339 ();
 sg13g2_decap_8 FILLER_45_1346 ();
 sg13g2_decap_8 FILLER_45_1353 ();
 sg13g2_decap_8 FILLER_45_1360 ();
 sg13g2_decap_8 FILLER_45_1367 ();
 sg13g2_decap_8 FILLER_45_1374 ();
 sg13g2_decap_8 FILLER_45_1381 ();
 sg13g2_decap_8 FILLER_45_1388 ();
 sg13g2_decap_8 FILLER_45_1395 ();
 sg13g2_decap_8 FILLER_45_1402 ();
 sg13g2_decap_8 FILLER_45_1409 ();
 sg13g2_decap_8 FILLER_45_1416 ();
 sg13g2_decap_8 FILLER_45_1423 ();
 sg13g2_decap_8 FILLER_45_1430 ();
 sg13g2_decap_8 FILLER_45_1437 ();
 sg13g2_decap_8 FILLER_45_1444 ();
 sg13g2_decap_8 FILLER_45_1451 ();
 sg13g2_decap_8 FILLER_45_1458 ();
 sg13g2_decap_8 FILLER_45_1465 ();
 sg13g2_decap_8 FILLER_45_1472 ();
 sg13g2_decap_8 FILLER_45_1479 ();
 sg13g2_decap_8 FILLER_45_1486 ();
 sg13g2_decap_8 FILLER_45_1493 ();
 sg13g2_decap_8 FILLER_45_1500 ();
 sg13g2_decap_8 FILLER_45_1507 ();
 sg13g2_decap_8 FILLER_45_1514 ();
 sg13g2_decap_8 FILLER_45_1521 ();
 sg13g2_decap_8 FILLER_45_1528 ();
 sg13g2_decap_8 FILLER_45_1535 ();
 sg13g2_decap_8 FILLER_45_1542 ();
 sg13g2_decap_8 FILLER_45_1549 ();
 sg13g2_decap_8 FILLER_45_1556 ();
 sg13g2_decap_8 FILLER_45_1563 ();
 sg13g2_decap_8 FILLER_45_1570 ();
 sg13g2_decap_8 FILLER_45_1577 ();
 sg13g2_decap_8 FILLER_45_1584 ();
 sg13g2_decap_8 FILLER_45_1591 ();
 sg13g2_decap_8 FILLER_45_1598 ();
 sg13g2_decap_8 FILLER_45_1605 ();
 sg13g2_decap_8 FILLER_45_1612 ();
 sg13g2_decap_8 FILLER_45_1619 ();
 sg13g2_decap_8 FILLER_45_1626 ();
 sg13g2_decap_8 FILLER_45_1633 ();
 sg13g2_decap_8 FILLER_45_1640 ();
 sg13g2_decap_8 FILLER_45_1647 ();
 sg13g2_decap_8 FILLER_45_1654 ();
 sg13g2_decap_8 FILLER_45_1661 ();
 sg13g2_decap_8 FILLER_45_1668 ();
 sg13g2_decap_8 FILLER_45_1675 ();
 sg13g2_decap_8 FILLER_45_1682 ();
 sg13g2_decap_8 FILLER_45_1689 ();
 sg13g2_decap_8 FILLER_45_1696 ();
 sg13g2_decap_8 FILLER_45_1703 ();
 sg13g2_decap_8 FILLER_45_1710 ();
 sg13g2_decap_8 FILLER_45_1717 ();
 sg13g2_decap_8 FILLER_45_1724 ();
 sg13g2_decap_8 FILLER_45_1731 ();
 sg13g2_decap_8 FILLER_45_1738 ();
 sg13g2_decap_8 FILLER_45_1745 ();
 sg13g2_decap_8 FILLER_45_1752 ();
 sg13g2_decap_8 FILLER_45_1759 ();
 sg13g2_fill_2 FILLER_45_1766 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_fill_2 FILLER_46_35 ();
 sg13g2_fill_1 FILLER_46_37 ();
 sg13g2_fill_2 FILLER_46_71 ();
 sg13g2_fill_2 FILLER_46_81 ();
 sg13g2_fill_1 FILLER_46_109 ();
 sg13g2_fill_2 FILLER_46_133 ();
 sg13g2_fill_1 FILLER_46_171 ();
 sg13g2_fill_2 FILLER_46_197 ();
 sg13g2_fill_2 FILLER_46_225 ();
 sg13g2_fill_1 FILLER_46_262 ();
 sg13g2_fill_2 FILLER_46_303 ();
 sg13g2_fill_1 FILLER_46_314 ();
 sg13g2_fill_2 FILLER_46_320 ();
 sg13g2_fill_2 FILLER_46_368 ();
 sg13g2_fill_1 FILLER_46_370 ();
 sg13g2_fill_2 FILLER_46_387 ();
 sg13g2_fill_2 FILLER_46_424 ();
 sg13g2_fill_1 FILLER_46_426 ();
 sg13g2_decap_4 FILLER_46_432 ();
 sg13g2_fill_2 FILLER_46_436 ();
 sg13g2_fill_2 FILLER_46_443 ();
 sg13g2_decap_4 FILLER_46_449 ();
 sg13g2_fill_1 FILLER_46_453 ();
 sg13g2_fill_2 FILLER_46_485 ();
 sg13g2_fill_1 FILLER_46_503 ();
 sg13g2_fill_2 FILLER_46_522 ();
 sg13g2_decap_4 FILLER_46_529 ();
 sg13g2_fill_2 FILLER_46_533 ();
 sg13g2_fill_2 FILLER_46_556 ();
 sg13g2_fill_2 FILLER_46_571 ();
 sg13g2_fill_1 FILLER_46_573 ();
 sg13g2_fill_1 FILLER_46_609 ();
 sg13g2_fill_2 FILLER_46_636 ();
 sg13g2_fill_1 FILLER_46_655 ();
 sg13g2_fill_1 FILLER_46_693 ();
 sg13g2_fill_1 FILLER_46_698 ();
 sg13g2_fill_2 FILLER_46_741 ();
 sg13g2_fill_1 FILLER_46_743 ();
 sg13g2_fill_2 FILLER_46_802 ();
 sg13g2_fill_1 FILLER_46_804 ();
 sg13g2_fill_1 FILLER_46_847 ();
 sg13g2_fill_1 FILLER_46_879 ();
 sg13g2_decap_4 FILLER_46_897 ();
 sg13g2_fill_2 FILLER_46_901 ();
 sg13g2_fill_1 FILLER_46_911 ();
 sg13g2_fill_2 FILLER_46_916 ();
 sg13g2_fill_1 FILLER_46_918 ();
 sg13g2_fill_2 FILLER_46_933 ();
 sg13g2_fill_1 FILLER_46_935 ();
 sg13g2_fill_1 FILLER_46_952 ();
 sg13g2_decap_4 FILLER_46_1017 ();
 sg13g2_decap_8 FILLER_46_1047 ();
 sg13g2_decap_8 FILLER_46_1054 ();
 sg13g2_decap_4 FILLER_46_1061 ();
 sg13g2_decap_8 FILLER_46_1074 ();
 sg13g2_decap_8 FILLER_46_1081 ();
 sg13g2_decap_8 FILLER_46_1088 ();
 sg13g2_decap_8 FILLER_46_1095 ();
 sg13g2_decap_8 FILLER_46_1102 ();
 sg13g2_decap_8 FILLER_46_1109 ();
 sg13g2_decap_8 FILLER_46_1116 ();
 sg13g2_decap_8 FILLER_46_1123 ();
 sg13g2_decap_8 FILLER_46_1130 ();
 sg13g2_decap_8 FILLER_46_1137 ();
 sg13g2_decap_8 FILLER_46_1144 ();
 sg13g2_decap_8 FILLER_46_1151 ();
 sg13g2_decap_8 FILLER_46_1158 ();
 sg13g2_decap_8 FILLER_46_1165 ();
 sg13g2_decap_8 FILLER_46_1172 ();
 sg13g2_decap_8 FILLER_46_1179 ();
 sg13g2_decap_8 FILLER_46_1186 ();
 sg13g2_decap_8 FILLER_46_1193 ();
 sg13g2_decap_8 FILLER_46_1200 ();
 sg13g2_decap_8 FILLER_46_1207 ();
 sg13g2_decap_8 FILLER_46_1214 ();
 sg13g2_decap_8 FILLER_46_1221 ();
 sg13g2_decap_8 FILLER_46_1228 ();
 sg13g2_decap_8 FILLER_46_1235 ();
 sg13g2_decap_8 FILLER_46_1242 ();
 sg13g2_decap_8 FILLER_46_1249 ();
 sg13g2_decap_8 FILLER_46_1256 ();
 sg13g2_decap_8 FILLER_46_1263 ();
 sg13g2_decap_8 FILLER_46_1270 ();
 sg13g2_decap_8 FILLER_46_1277 ();
 sg13g2_decap_8 FILLER_46_1284 ();
 sg13g2_decap_8 FILLER_46_1291 ();
 sg13g2_decap_8 FILLER_46_1298 ();
 sg13g2_decap_8 FILLER_46_1305 ();
 sg13g2_decap_8 FILLER_46_1312 ();
 sg13g2_decap_8 FILLER_46_1319 ();
 sg13g2_decap_8 FILLER_46_1326 ();
 sg13g2_decap_8 FILLER_46_1333 ();
 sg13g2_decap_8 FILLER_46_1340 ();
 sg13g2_decap_8 FILLER_46_1347 ();
 sg13g2_decap_8 FILLER_46_1354 ();
 sg13g2_decap_8 FILLER_46_1361 ();
 sg13g2_decap_8 FILLER_46_1368 ();
 sg13g2_decap_8 FILLER_46_1375 ();
 sg13g2_decap_8 FILLER_46_1382 ();
 sg13g2_decap_8 FILLER_46_1389 ();
 sg13g2_decap_8 FILLER_46_1396 ();
 sg13g2_decap_8 FILLER_46_1403 ();
 sg13g2_decap_8 FILLER_46_1410 ();
 sg13g2_decap_8 FILLER_46_1417 ();
 sg13g2_decap_8 FILLER_46_1424 ();
 sg13g2_decap_8 FILLER_46_1431 ();
 sg13g2_decap_8 FILLER_46_1438 ();
 sg13g2_decap_8 FILLER_46_1445 ();
 sg13g2_decap_8 FILLER_46_1452 ();
 sg13g2_decap_8 FILLER_46_1459 ();
 sg13g2_decap_8 FILLER_46_1466 ();
 sg13g2_decap_8 FILLER_46_1473 ();
 sg13g2_decap_8 FILLER_46_1480 ();
 sg13g2_decap_8 FILLER_46_1487 ();
 sg13g2_decap_8 FILLER_46_1494 ();
 sg13g2_decap_8 FILLER_46_1501 ();
 sg13g2_decap_8 FILLER_46_1508 ();
 sg13g2_decap_8 FILLER_46_1515 ();
 sg13g2_decap_8 FILLER_46_1522 ();
 sg13g2_decap_8 FILLER_46_1529 ();
 sg13g2_decap_8 FILLER_46_1536 ();
 sg13g2_decap_8 FILLER_46_1543 ();
 sg13g2_decap_8 FILLER_46_1550 ();
 sg13g2_decap_8 FILLER_46_1557 ();
 sg13g2_decap_8 FILLER_46_1564 ();
 sg13g2_decap_8 FILLER_46_1571 ();
 sg13g2_decap_8 FILLER_46_1578 ();
 sg13g2_decap_8 FILLER_46_1585 ();
 sg13g2_decap_8 FILLER_46_1592 ();
 sg13g2_decap_8 FILLER_46_1599 ();
 sg13g2_decap_8 FILLER_46_1606 ();
 sg13g2_decap_8 FILLER_46_1613 ();
 sg13g2_decap_8 FILLER_46_1620 ();
 sg13g2_decap_8 FILLER_46_1627 ();
 sg13g2_decap_8 FILLER_46_1634 ();
 sg13g2_decap_8 FILLER_46_1641 ();
 sg13g2_decap_8 FILLER_46_1648 ();
 sg13g2_decap_8 FILLER_46_1655 ();
 sg13g2_decap_8 FILLER_46_1662 ();
 sg13g2_decap_8 FILLER_46_1669 ();
 sg13g2_decap_8 FILLER_46_1676 ();
 sg13g2_decap_8 FILLER_46_1683 ();
 sg13g2_decap_8 FILLER_46_1690 ();
 sg13g2_decap_8 FILLER_46_1697 ();
 sg13g2_decap_8 FILLER_46_1704 ();
 sg13g2_decap_8 FILLER_46_1711 ();
 sg13g2_decap_8 FILLER_46_1718 ();
 sg13g2_decap_8 FILLER_46_1725 ();
 sg13g2_decap_8 FILLER_46_1732 ();
 sg13g2_decap_8 FILLER_46_1739 ();
 sg13g2_decap_8 FILLER_46_1746 ();
 sg13g2_decap_8 FILLER_46_1753 ();
 sg13g2_decap_8 FILLER_46_1760 ();
 sg13g2_fill_1 FILLER_46_1767 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_4 FILLER_47_35 ();
 sg13g2_fill_2 FILLER_47_70 ();
 sg13g2_fill_2 FILLER_47_113 ();
 sg13g2_fill_2 FILLER_47_181 ();
 sg13g2_fill_2 FILLER_47_204 ();
 sg13g2_fill_1 FILLER_47_253 ();
 sg13g2_fill_2 FILLER_47_314 ();
 sg13g2_fill_1 FILLER_47_316 ();
 sg13g2_fill_1 FILLER_47_341 ();
 sg13g2_fill_2 FILLER_47_352 ();
 sg13g2_fill_2 FILLER_47_372 ();
 sg13g2_fill_1 FILLER_47_374 ();
 sg13g2_fill_2 FILLER_47_380 ();
 sg13g2_fill_1 FILLER_47_382 ();
 sg13g2_fill_2 FILLER_47_425 ();
 sg13g2_fill_2 FILLER_47_443 ();
 sg13g2_fill_2 FILLER_47_454 ();
 sg13g2_decap_8 FILLER_47_461 ();
 sg13g2_decap_8 FILLER_47_468 ();
 sg13g2_decap_4 FILLER_47_475 ();
 sg13g2_fill_1 FILLER_47_479 ();
 sg13g2_fill_2 FILLER_47_501 ();
 sg13g2_fill_1 FILLER_47_503 ();
 sg13g2_decap_4 FILLER_47_509 ();
 sg13g2_fill_2 FILLER_47_539 ();
 sg13g2_fill_1 FILLER_47_583 ();
 sg13g2_fill_2 FILLER_47_635 ();
 sg13g2_fill_2 FILLER_47_646 ();
 sg13g2_fill_2 FILLER_47_670 ();
 sg13g2_fill_1 FILLER_47_707 ();
 sg13g2_fill_2 FILLER_47_766 ();
 sg13g2_fill_1 FILLER_47_768 ();
 sg13g2_fill_2 FILLER_47_795 ();
 sg13g2_fill_1 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_817 ();
 sg13g2_fill_1 FILLER_47_824 ();
 sg13g2_decap_8 FILLER_47_846 ();
 sg13g2_decap_4 FILLER_47_853 ();
 sg13g2_fill_1 FILLER_47_857 ();
 sg13g2_fill_2 FILLER_47_863 ();
 sg13g2_fill_1 FILLER_47_865 ();
 sg13g2_decap_4 FILLER_47_897 ();
 sg13g2_fill_2 FILLER_47_963 ();
 sg13g2_decap_8 FILLER_47_974 ();
 sg13g2_decap_4 FILLER_47_990 ();
 sg13g2_fill_1 FILLER_47_994 ();
 sg13g2_fill_1 FILLER_47_1034 ();
 sg13g2_decap_8 FILLER_47_1043 ();
 sg13g2_decap_8 FILLER_47_1050 ();
 sg13g2_decap_8 FILLER_47_1057 ();
 sg13g2_decap_8 FILLER_47_1064 ();
 sg13g2_decap_8 FILLER_47_1071 ();
 sg13g2_decap_8 FILLER_47_1078 ();
 sg13g2_decap_8 FILLER_47_1085 ();
 sg13g2_decap_8 FILLER_47_1092 ();
 sg13g2_decap_8 FILLER_47_1099 ();
 sg13g2_decap_8 FILLER_47_1106 ();
 sg13g2_decap_8 FILLER_47_1113 ();
 sg13g2_decap_8 FILLER_47_1120 ();
 sg13g2_decap_8 FILLER_47_1127 ();
 sg13g2_decap_8 FILLER_47_1134 ();
 sg13g2_decap_8 FILLER_47_1141 ();
 sg13g2_decap_8 FILLER_47_1148 ();
 sg13g2_decap_8 FILLER_47_1155 ();
 sg13g2_decap_8 FILLER_47_1162 ();
 sg13g2_decap_8 FILLER_47_1169 ();
 sg13g2_decap_8 FILLER_47_1176 ();
 sg13g2_decap_8 FILLER_47_1183 ();
 sg13g2_decap_8 FILLER_47_1190 ();
 sg13g2_decap_8 FILLER_47_1197 ();
 sg13g2_decap_8 FILLER_47_1204 ();
 sg13g2_decap_8 FILLER_47_1211 ();
 sg13g2_decap_8 FILLER_47_1218 ();
 sg13g2_decap_8 FILLER_47_1225 ();
 sg13g2_decap_8 FILLER_47_1232 ();
 sg13g2_decap_8 FILLER_47_1239 ();
 sg13g2_decap_8 FILLER_47_1246 ();
 sg13g2_decap_8 FILLER_47_1253 ();
 sg13g2_decap_8 FILLER_47_1260 ();
 sg13g2_decap_8 FILLER_47_1267 ();
 sg13g2_decap_8 FILLER_47_1274 ();
 sg13g2_decap_8 FILLER_47_1281 ();
 sg13g2_decap_8 FILLER_47_1288 ();
 sg13g2_decap_8 FILLER_47_1295 ();
 sg13g2_decap_8 FILLER_47_1302 ();
 sg13g2_decap_8 FILLER_47_1309 ();
 sg13g2_decap_8 FILLER_47_1316 ();
 sg13g2_decap_8 FILLER_47_1323 ();
 sg13g2_decap_8 FILLER_47_1330 ();
 sg13g2_decap_8 FILLER_47_1337 ();
 sg13g2_decap_8 FILLER_47_1344 ();
 sg13g2_decap_8 FILLER_47_1351 ();
 sg13g2_decap_8 FILLER_47_1358 ();
 sg13g2_decap_8 FILLER_47_1365 ();
 sg13g2_decap_8 FILLER_47_1372 ();
 sg13g2_decap_8 FILLER_47_1379 ();
 sg13g2_decap_8 FILLER_47_1386 ();
 sg13g2_decap_8 FILLER_47_1393 ();
 sg13g2_decap_8 FILLER_47_1400 ();
 sg13g2_decap_8 FILLER_47_1407 ();
 sg13g2_decap_8 FILLER_47_1414 ();
 sg13g2_decap_8 FILLER_47_1421 ();
 sg13g2_decap_8 FILLER_47_1428 ();
 sg13g2_decap_8 FILLER_47_1435 ();
 sg13g2_decap_8 FILLER_47_1442 ();
 sg13g2_decap_8 FILLER_47_1449 ();
 sg13g2_decap_8 FILLER_47_1456 ();
 sg13g2_decap_8 FILLER_47_1463 ();
 sg13g2_decap_8 FILLER_47_1470 ();
 sg13g2_decap_8 FILLER_47_1477 ();
 sg13g2_decap_8 FILLER_47_1484 ();
 sg13g2_decap_8 FILLER_47_1491 ();
 sg13g2_decap_8 FILLER_47_1498 ();
 sg13g2_decap_8 FILLER_47_1505 ();
 sg13g2_decap_8 FILLER_47_1512 ();
 sg13g2_decap_8 FILLER_47_1519 ();
 sg13g2_decap_8 FILLER_47_1526 ();
 sg13g2_decap_8 FILLER_47_1533 ();
 sg13g2_decap_8 FILLER_47_1540 ();
 sg13g2_decap_8 FILLER_47_1547 ();
 sg13g2_decap_8 FILLER_47_1554 ();
 sg13g2_decap_8 FILLER_47_1561 ();
 sg13g2_decap_8 FILLER_47_1568 ();
 sg13g2_decap_8 FILLER_47_1575 ();
 sg13g2_decap_8 FILLER_47_1582 ();
 sg13g2_decap_8 FILLER_47_1589 ();
 sg13g2_decap_8 FILLER_47_1596 ();
 sg13g2_decap_8 FILLER_47_1603 ();
 sg13g2_decap_8 FILLER_47_1610 ();
 sg13g2_decap_8 FILLER_47_1617 ();
 sg13g2_decap_8 FILLER_47_1624 ();
 sg13g2_decap_8 FILLER_47_1631 ();
 sg13g2_decap_8 FILLER_47_1638 ();
 sg13g2_decap_8 FILLER_47_1645 ();
 sg13g2_decap_8 FILLER_47_1652 ();
 sg13g2_decap_8 FILLER_47_1659 ();
 sg13g2_decap_8 FILLER_47_1666 ();
 sg13g2_decap_8 FILLER_47_1673 ();
 sg13g2_decap_8 FILLER_47_1680 ();
 sg13g2_decap_8 FILLER_47_1687 ();
 sg13g2_decap_8 FILLER_47_1694 ();
 sg13g2_decap_8 FILLER_47_1701 ();
 sg13g2_decap_8 FILLER_47_1708 ();
 sg13g2_decap_8 FILLER_47_1715 ();
 sg13g2_decap_8 FILLER_47_1722 ();
 sg13g2_decap_8 FILLER_47_1729 ();
 sg13g2_decap_8 FILLER_47_1736 ();
 sg13g2_decap_8 FILLER_47_1743 ();
 sg13g2_decap_8 FILLER_47_1750 ();
 sg13g2_decap_8 FILLER_47_1757 ();
 sg13g2_decap_4 FILLER_47_1764 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_4 FILLER_48_14 ();
 sg13g2_fill_1 FILLER_48_18 ();
 sg13g2_fill_1 FILLER_48_68 ();
 sg13g2_fill_2 FILLER_48_139 ();
 sg13g2_fill_2 FILLER_48_156 ();
 sg13g2_fill_1 FILLER_48_163 ();
 sg13g2_fill_1 FILLER_48_191 ();
 sg13g2_decap_8 FILLER_48_253 ();
 sg13g2_decap_8 FILLER_48_260 ();
 sg13g2_fill_2 FILLER_48_267 ();
 sg13g2_fill_1 FILLER_48_269 ();
 sg13g2_decap_4 FILLER_48_320 ();
 sg13g2_fill_1 FILLER_48_385 ();
 sg13g2_fill_1 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_484 ();
 sg13g2_fill_1 FILLER_48_491 ();
 sg13g2_fill_1 FILLER_48_500 ();
 sg13g2_decap_8 FILLER_48_522 ();
 sg13g2_decap_4 FILLER_48_529 ();
 sg13g2_fill_2 FILLER_48_533 ();
 sg13g2_fill_1 FILLER_48_539 ();
 sg13g2_fill_2 FILLER_48_545 ();
 sg13g2_fill_1 FILLER_48_633 ();
 sg13g2_fill_2 FILLER_48_652 ();
 sg13g2_fill_2 FILLER_48_668 ();
 sg13g2_fill_1 FILLER_48_757 ();
 sg13g2_fill_1 FILLER_48_781 ();
 sg13g2_fill_2 FILLER_48_808 ();
 sg13g2_fill_2 FILLER_48_828 ();
 sg13g2_fill_1 FILLER_48_830 ();
 sg13g2_decap_8 FILLER_48_834 ();
 sg13g2_fill_2 FILLER_48_841 ();
 sg13g2_decap_4 FILLER_48_873 ();
 sg13g2_decap_8 FILLER_48_893 ();
 sg13g2_fill_2 FILLER_48_900 ();
 sg13g2_decap_4 FILLER_48_910 ();
 sg13g2_fill_2 FILLER_48_914 ();
 sg13g2_decap_4 FILLER_48_920 ();
 sg13g2_fill_1 FILLER_48_924 ();
 sg13g2_decap_4 FILLER_48_938 ();
 sg13g2_fill_2 FILLER_48_956 ();
 sg13g2_fill_2 FILLER_48_963 ();
 sg13g2_fill_1 FILLER_48_965 ();
 sg13g2_decap_8 FILLER_48_992 ();
 sg13g2_fill_2 FILLER_48_999 ();
 sg13g2_decap_8 FILLER_48_1027 ();
 sg13g2_decap_8 FILLER_48_1034 ();
 sg13g2_decap_8 FILLER_48_1041 ();
 sg13g2_decap_8 FILLER_48_1048 ();
 sg13g2_decap_8 FILLER_48_1055 ();
 sg13g2_decap_8 FILLER_48_1062 ();
 sg13g2_decap_8 FILLER_48_1069 ();
 sg13g2_decap_8 FILLER_48_1076 ();
 sg13g2_decap_8 FILLER_48_1083 ();
 sg13g2_decap_8 FILLER_48_1090 ();
 sg13g2_decap_8 FILLER_48_1097 ();
 sg13g2_decap_8 FILLER_48_1104 ();
 sg13g2_decap_8 FILLER_48_1111 ();
 sg13g2_decap_8 FILLER_48_1118 ();
 sg13g2_decap_8 FILLER_48_1125 ();
 sg13g2_decap_8 FILLER_48_1132 ();
 sg13g2_decap_8 FILLER_48_1139 ();
 sg13g2_decap_8 FILLER_48_1146 ();
 sg13g2_decap_8 FILLER_48_1153 ();
 sg13g2_decap_8 FILLER_48_1160 ();
 sg13g2_decap_8 FILLER_48_1167 ();
 sg13g2_decap_8 FILLER_48_1174 ();
 sg13g2_decap_8 FILLER_48_1181 ();
 sg13g2_decap_8 FILLER_48_1188 ();
 sg13g2_decap_8 FILLER_48_1195 ();
 sg13g2_decap_8 FILLER_48_1202 ();
 sg13g2_decap_8 FILLER_48_1209 ();
 sg13g2_decap_8 FILLER_48_1216 ();
 sg13g2_decap_8 FILLER_48_1223 ();
 sg13g2_decap_8 FILLER_48_1230 ();
 sg13g2_decap_8 FILLER_48_1237 ();
 sg13g2_decap_8 FILLER_48_1244 ();
 sg13g2_decap_8 FILLER_48_1251 ();
 sg13g2_decap_8 FILLER_48_1258 ();
 sg13g2_decap_8 FILLER_48_1265 ();
 sg13g2_decap_8 FILLER_48_1272 ();
 sg13g2_decap_8 FILLER_48_1279 ();
 sg13g2_decap_8 FILLER_48_1286 ();
 sg13g2_decap_8 FILLER_48_1293 ();
 sg13g2_decap_8 FILLER_48_1300 ();
 sg13g2_decap_8 FILLER_48_1307 ();
 sg13g2_decap_8 FILLER_48_1314 ();
 sg13g2_decap_8 FILLER_48_1321 ();
 sg13g2_decap_8 FILLER_48_1328 ();
 sg13g2_decap_8 FILLER_48_1335 ();
 sg13g2_decap_8 FILLER_48_1342 ();
 sg13g2_decap_8 FILLER_48_1349 ();
 sg13g2_decap_8 FILLER_48_1356 ();
 sg13g2_decap_8 FILLER_48_1363 ();
 sg13g2_decap_8 FILLER_48_1370 ();
 sg13g2_decap_8 FILLER_48_1377 ();
 sg13g2_decap_8 FILLER_48_1384 ();
 sg13g2_decap_8 FILLER_48_1391 ();
 sg13g2_decap_8 FILLER_48_1398 ();
 sg13g2_decap_8 FILLER_48_1405 ();
 sg13g2_decap_8 FILLER_48_1412 ();
 sg13g2_decap_8 FILLER_48_1419 ();
 sg13g2_decap_8 FILLER_48_1426 ();
 sg13g2_decap_8 FILLER_48_1433 ();
 sg13g2_decap_8 FILLER_48_1440 ();
 sg13g2_decap_8 FILLER_48_1447 ();
 sg13g2_decap_8 FILLER_48_1454 ();
 sg13g2_decap_8 FILLER_48_1461 ();
 sg13g2_decap_8 FILLER_48_1468 ();
 sg13g2_decap_8 FILLER_48_1475 ();
 sg13g2_decap_8 FILLER_48_1482 ();
 sg13g2_decap_8 FILLER_48_1489 ();
 sg13g2_decap_8 FILLER_48_1496 ();
 sg13g2_decap_8 FILLER_48_1503 ();
 sg13g2_decap_8 FILLER_48_1510 ();
 sg13g2_decap_8 FILLER_48_1517 ();
 sg13g2_decap_8 FILLER_48_1524 ();
 sg13g2_decap_8 FILLER_48_1531 ();
 sg13g2_decap_8 FILLER_48_1538 ();
 sg13g2_decap_8 FILLER_48_1545 ();
 sg13g2_decap_8 FILLER_48_1552 ();
 sg13g2_decap_8 FILLER_48_1559 ();
 sg13g2_decap_8 FILLER_48_1566 ();
 sg13g2_decap_8 FILLER_48_1573 ();
 sg13g2_decap_8 FILLER_48_1580 ();
 sg13g2_decap_8 FILLER_48_1587 ();
 sg13g2_decap_8 FILLER_48_1594 ();
 sg13g2_decap_8 FILLER_48_1601 ();
 sg13g2_decap_8 FILLER_48_1608 ();
 sg13g2_decap_8 FILLER_48_1615 ();
 sg13g2_decap_8 FILLER_48_1622 ();
 sg13g2_decap_8 FILLER_48_1629 ();
 sg13g2_decap_8 FILLER_48_1636 ();
 sg13g2_decap_8 FILLER_48_1643 ();
 sg13g2_decap_8 FILLER_48_1650 ();
 sg13g2_decap_8 FILLER_48_1657 ();
 sg13g2_decap_8 FILLER_48_1664 ();
 sg13g2_decap_8 FILLER_48_1671 ();
 sg13g2_decap_8 FILLER_48_1678 ();
 sg13g2_decap_8 FILLER_48_1685 ();
 sg13g2_decap_8 FILLER_48_1692 ();
 sg13g2_decap_8 FILLER_48_1699 ();
 sg13g2_decap_8 FILLER_48_1706 ();
 sg13g2_decap_8 FILLER_48_1713 ();
 sg13g2_decap_8 FILLER_48_1720 ();
 sg13g2_decap_8 FILLER_48_1727 ();
 sg13g2_decap_8 FILLER_48_1734 ();
 sg13g2_decap_8 FILLER_48_1741 ();
 sg13g2_decap_8 FILLER_48_1748 ();
 sg13g2_decap_8 FILLER_48_1755 ();
 sg13g2_decap_4 FILLER_48_1762 ();
 sg13g2_fill_2 FILLER_48_1766 ();
 sg13g2_fill_2 FILLER_49_26 ();
 sg13g2_fill_2 FILLER_49_37 ();
 sg13g2_fill_1 FILLER_49_49 ();
 sg13g2_fill_2 FILLER_49_60 ();
 sg13g2_fill_1 FILLER_49_73 ();
 sg13g2_fill_2 FILLER_49_106 ();
 sg13g2_fill_1 FILLER_49_108 ();
 sg13g2_fill_1 FILLER_49_113 ();
 sg13g2_fill_2 FILLER_49_118 ();
 sg13g2_fill_2 FILLER_49_192 ();
 sg13g2_fill_2 FILLER_49_202 ();
 sg13g2_fill_1 FILLER_49_233 ();
 sg13g2_decap_4 FILLER_49_253 ();
 sg13g2_fill_2 FILLER_49_283 ();
 sg13g2_fill_2 FILLER_49_316 ();
 sg13g2_fill_2 FILLER_49_343 ();
 sg13g2_fill_2 FILLER_49_366 ();
 sg13g2_fill_1 FILLER_49_401 ();
 sg13g2_fill_1 FILLER_49_419 ();
 sg13g2_decap_8 FILLER_49_452 ();
 sg13g2_decap_8 FILLER_49_459 ();
 sg13g2_fill_1 FILLER_49_466 ();
 sg13g2_fill_1 FILLER_49_475 ();
 sg13g2_fill_2 FILLER_49_482 ();
 sg13g2_decap_4 FILLER_49_494 ();
 sg13g2_decap_8 FILLER_49_506 ();
 sg13g2_fill_1 FILLER_49_513 ();
 sg13g2_fill_2 FILLER_49_550 ();
 sg13g2_fill_1 FILLER_49_552 ();
 sg13g2_fill_1 FILLER_49_569 ();
 sg13g2_fill_2 FILLER_49_596 ();
 sg13g2_decap_4 FILLER_49_643 ();
 sg13g2_fill_1 FILLER_49_647 ();
 sg13g2_fill_1 FILLER_49_663 ();
 sg13g2_fill_2 FILLER_49_678 ();
 sg13g2_fill_1 FILLER_49_735 ();
 sg13g2_fill_2 FILLER_49_771 ();
 sg13g2_fill_2 FILLER_49_796 ();
 sg13g2_fill_1 FILLER_49_798 ();
 sg13g2_fill_1 FILLER_49_871 ();
 sg13g2_fill_1 FILLER_49_910 ();
 sg13g2_decap_8 FILLER_49_928 ();
 sg13g2_decap_8 FILLER_49_935 ();
 sg13g2_decap_8 FILLER_49_942 ();
 sg13g2_decap_8 FILLER_49_949 ();
 sg13g2_decap_8 FILLER_49_965 ();
 sg13g2_fill_2 FILLER_49_972 ();
 sg13g2_fill_1 FILLER_49_974 ();
 sg13g2_decap_8 FILLER_49_984 ();
 sg13g2_decap_8 FILLER_49_991 ();
 sg13g2_decap_8 FILLER_49_998 ();
 sg13g2_decap_8 FILLER_49_1005 ();
 sg13g2_decap_8 FILLER_49_1012 ();
 sg13g2_decap_8 FILLER_49_1019 ();
 sg13g2_decap_8 FILLER_49_1026 ();
 sg13g2_decap_8 FILLER_49_1033 ();
 sg13g2_decap_8 FILLER_49_1040 ();
 sg13g2_decap_8 FILLER_49_1047 ();
 sg13g2_decap_8 FILLER_49_1054 ();
 sg13g2_decap_8 FILLER_49_1061 ();
 sg13g2_decap_8 FILLER_49_1068 ();
 sg13g2_decap_8 FILLER_49_1075 ();
 sg13g2_decap_8 FILLER_49_1082 ();
 sg13g2_decap_8 FILLER_49_1089 ();
 sg13g2_decap_8 FILLER_49_1096 ();
 sg13g2_decap_8 FILLER_49_1103 ();
 sg13g2_decap_8 FILLER_49_1110 ();
 sg13g2_decap_8 FILLER_49_1117 ();
 sg13g2_decap_8 FILLER_49_1124 ();
 sg13g2_decap_8 FILLER_49_1131 ();
 sg13g2_decap_8 FILLER_49_1138 ();
 sg13g2_decap_8 FILLER_49_1145 ();
 sg13g2_decap_8 FILLER_49_1152 ();
 sg13g2_decap_8 FILLER_49_1159 ();
 sg13g2_decap_8 FILLER_49_1166 ();
 sg13g2_decap_8 FILLER_49_1173 ();
 sg13g2_decap_8 FILLER_49_1180 ();
 sg13g2_decap_8 FILLER_49_1187 ();
 sg13g2_decap_8 FILLER_49_1194 ();
 sg13g2_decap_8 FILLER_49_1201 ();
 sg13g2_decap_8 FILLER_49_1208 ();
 sg13g2_decap_8 FILLER_49_1215 ();
 sg13g2_decap_8 FILLER_49_1222 ();
 sg13g2_decap_8 FILLER_49_1229 ();
 sg13g2_decap_8 FILLER_49_1236 ();
 sg13g2_decap_8 FILLER_49_1243 ();
 sg13g2_decap_8 FILLER_49_1250 ();
 sg13g2_decap_8 FILLER_49_1257 ();
 sg13g2_decap_8 FILLER_49_1264 ();
 sg13g2_decap_8 FILLER_49_1271 ();
 sg13g2_decap_8 FILLER_49_1278 ();
 sg13g2_decap_8 FILLER_49_1285 ();
 sg13g2_decap_8 FILLER_49_1292 ();
 sg13g2_decap_8 FILLER_49_1299 ();
 sg13g2_decap_8 FILLER_49_1306 ();
 sg13g2_decap_8 FILLER_49_1313 ();
 sg13g2_decap_8 FILLER_49_1320 ();
 sg13g2_decap_8 FILLER_49_1327 ();
 sg13g2_decap_8 FILLER_49_1334 ();
 sg13g2_decap_8 FILLER_49_1341 ();
 sg13g2_decap_8 FILLER_49_1348 ();
 sg13g2_decap_8 FILLER_49_1355 ();
 sg13g2_decap_8 FILLER_49_1362 ();
 sg13g2_decap_8 FILLER_49_1369 ();
 sg13g2_decap_8 FILLER_49_1376 ();
 sg13g2_decap_8 FILLER_49_1383 ();
 sg13g2_decap_8 FILLER_49_1390 ();
 sg13g2_decap_8 FILLER_49_1397 ();
 sg13g2_decap_8 FILLER_49_1404 ();
 sg13g2_decap_8 FILLER_49_1411 ();
 sg13g2_decap_8 FILLER_49_1418 ();
 sg13g2_decap_8 FILLER_49_1425 ();
 sg13g2_decap_8 FILLER_49_1432 ();
 sg13g2_decap_8 FILLER_49_1439 ();
 sg13g2_decap_8 FILLER_49_1446 ();
 sg13g2_decap_8 FILLER_49_1453 ();
 sg13g2_decap_8 FILLER_49_1460 ();
 sg13g2_decap_8 FILLER_49_1467 ();
 sg13g2_decap_8 FILLER_49_1474 ();
 sg13g2_decap_8 FILLER_49_1481 ();
 sg13g2_decap_8 FILLER_49_1488 ();
 sg13g2_decap_8 FILLER_49_1495 ();
 sg13g2_decap_8 FILLER_49_1502 ();
 sg13g2_decap_8 FILLER_49_1509 ();
 sg13g2_decap_8 FILLER_49_1516 ();
 sg13g2_decap_8 FILLER_49_1523 ();
 sg13g2_decap_8 FILLER_49_1530 ();
 sg13g2_decap_8 FILLER_49_1537 ();
 sg13g2_decap_8 FILLER_49_1544 ();
 sg13g2_decap_8 FILLER_49_1551 ();
 sg13g2_decap_8 FILLER_49_1558 ();
 sg13g2_decap_8 FILLER_49_1565 ();
 sg13g2_decap_8 FILLER_49_1572 ();
 sg13g2_decap_8 FILLER_49_1579 ();
 sg13g2_decap_8 FILLER_49_1586 ();
 sg13g2_decap_8 FILLER_49_1593 ();
 sg13g2_decap_8 FILLER_49_1600 ();
 sg13g2_decap_8 FILLER_49_1607 ();
 sg13g2_decap_8 FILLER_49_1614 ();
 sg13g2_decap_8 FILLER_49_1621 ();
 sg13g2_decap_8 FILLER_49_1628 ();
 sg13g2_decap_8 FILLER_49_1635 ();
 sg13g2_decap_8 FILLER_49_1642 ();
 sg13g2_decap_8 FILLER_49_1649 ();
 sg13g2_decap_8 FILLER_49_1656 ();
 sg13g2_decap_8 FILLER_49_1663 ();
 sg13g2_decap_8 FILLER_49_1670 ();
 sg13g2_decap_8 FILLER_49_1677 ();
 sg13g2_decap_8 FILLER_49_1684 ();
 sg13g2_decap_8 FILLER_49_1691 ();
 sg13g2_decap_8 FILLER_49_1698 ();
 sg13g2_decap_8 FILLER_49_1705 ();
 sg13g2_decap_8 FILLER_49_1712 ();
 sg13g2_decap_8 FILLER_49_1719 ();
 sg13g2_decap_8 FILLER_49_1726 ();
 sg13g2_decap_8 FILLER_49_1733 ();
 sg13g2_decap_8 FILLER_49_1740 ();
 sg13g2_decap_8 FILLER_49_1747 ();
 sg13g2_decap_8 FILLER_49_1754 ();
 sg13g2_decap_8 FILLER_49_1761 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_9 ();
 sg13g2_fill_1 FILLER_50_23 ();
 sg13g2_fill_1 FILLER_50_40 ();
 sg13g2_fill_1 FILLER_50_63 ();
 sg13g2_fill_2 FILLER_50_76 ();
 sg13g2_fill_1 FILLER_50_78 ();
 sg13g2_fill_1 FILLER_50_105 ();
 sg13g2_fill_1 FILLER_50_120 ();
 sg13g2_decap_4 FILLER_50_160 ();
 sg13g2_fill_1 FILLER_50_193 ();
 sg13g2_fill_2 FILLER_50_258 ();
 sg13g2_fill_1 FILLER_50_260 ();
 sg13g2_fill_2 FILLER_50_316 ();
 sg13g2_fill_1 FILLER_50_362 ();
 sg13g2_decap_8 FILLER_50_434 ();
 sg13g2_fill_2 FILLER_50_441 ();
 sg13g2_fill_1 FILLER_50_451 ();
 sg13g2_decap_8 FILLER_50_460 ();
 sg13g2_fill_2 FILLER_50_476 ();
 sg13g2_decap_8 FILLER_50_491 ();
 sg13g2_fill_2 FILLER_50_498 ();
 sg13g2_fill_1 FILLER_50_508 ();
 sg13g2_fill_2 FILLER_50_523 ();
 sg13g2_fill_1 FILLER_50_525 ();
 sg13g2_fill_2 FILLER_50_534 ();
 sg13g2_fill_1 FILLER_50_552 ();
 sg13g2_fill_2 FILLER_50_576 ();
 sg13g2_fill_1 FILLER_50_578 ();
 sg13g2_fill_1 FILLER_50_622 ();
 sg13g2_decap_8 FILLER_50_648 ();
 sg13g2_decap_4 FILLER_50_710 ();
 sg13g2_decap_4 FILLER_50_717 ();
 sg13g2_fill_2 FILLER_50_721 ();
 sg13g2_fill_1 FILLER_50_783 ();
 sg13g2_fill_2 FILLER_50_795 ();
 sg13g2_fill_2 FILLER_50_826 ();
 sg13g2_fill_2 FILLER_50_832 ();
 sg13g2_fill_2 FILLER_50_849 ();
 sg13g2_decap_4 FILLER_50_870 ();
 sg13g2_fill_1 FILLER_50_874 ();
 sg13g2_decap_4 FILLER_50_894 ();
 sg13g2_fill_2 FILLER_50_898 ();
 sg13g2_decap_8 FILLER_50_946 ();
 sg13g2_decap_8 FILLER_50_953 ();
 sg13g2_decap_8 FILLER_50_960 ();
 sg13g2_decap_8 FILLER_50_967 ();
 sg13g2_decap_8 FILLER_50_974 ();
 sg13g2_decap_8 FILLER_50_981 ();
 sg13g2_decap_8 FILLER_50_988 ();
 sg13g2_decap_8 FILLER_50_995 ();
 sg13g2_decap_4 FILLER_50_1002 ();
 sg13g2_decap_8 FILLER_50_1012 ();
 sg13g2_decap_8 FILLER_50_1019 ();
 sg13g2_decap_8 FILLER_50_1026 ();
 sg13g2_decap_8 FILLER_50_1033 ();
 sg13g2_decap_8 FILLER_50_1040 ();
 sg13g2_decap_8 FILLER_50_1047 ();
 sg13g2_decap_8 FILLER_50_1054 ();
 sg13g2_decap_8 FILLER_50_1061 ();
 sg13g2_decap_8 FILLER_50_1068 ();
 sg13g2_decap_8 FILLER_50_1075 ();
 sg13g2_decap_8 FILLER_50_1082 ();
 sg13g2_decap_8 FILLER_50_1089 ();
 sg13g2_decap_8 FILLER_50_1096 ();
 sg13g2_decap_8 FILLER_50_1103 ();
 sg13g2_decap_8 FILLER_50_1110 ();
 sg13g2_decap_8 FILLER_50_1117 ();
 sg13g2_decap_8 FILLER_50_1124 ();
 sg13g2_decap_8 FILLER_50_1131 ();
 sg13g2_decap_8 FILLER_50_1138 ();
 sg13g2_decap_8 FILLER_50_1145 ();
 sg13g2_decap_8 FILLER_50_1152 ();
 sg13g2_decap_8 FILLER_50_1159 ();
 sg13g2_decap_8 FILLER_50_1166 ();
 sg13g2_decap_8 FILLER_50_1173 ();
 sg13g2_decap_8 FILLER_50_1180 ();
 sg13g2_decap_8 FILLER_50_1187 ();
 sg13g2_decap_8 FILLER_50_1194 ();
 sg13g2_decap_8 FILLER_50_1201 ();
 sg13g2_decap_8 FILLER_50_1208 ();
 sg13g2_decap_8 FILLER_50_1215 ();
 sg13g2_decap_8 FILLER_50_1222 ();
 sg13g2_decap_8 FILLER_50_1229 ();
 sg13g2_decap_8 FILLER_50_1236 ();
 sg13g2_decap_8 FILLER_50_1243 ();
 sg13g2_decap_8 FILLER_50_1250 ();
 sg13g2_decap_8 FILLER_50_1257 ();
 sg13g2_decap_8 FILLER_50_1264 ();
 sg13g2_decap_8 FILLER_50_1271 ();
 sg13g2_decap_8 FILLER_50_1278 ();
 sg13g2_decap_8 FILLER_50_1285 ();
 sg13g2_decap_8 FILLER_50_1292 ();
 sg13g2_decap_8 FILLER_50_1299 ();
 sg13g2_decap_8 FILLER_50_1306 ();
 sg13g2_decap_8 FILLER_50_1313 ();
 sg13g2_decap_8 FILLER_50_1320 ();
 sg13g2_decap_8 FILLER_50_1327 ();
 sg13g2_decap_8 FILLER_50_1334 ();
 sg13g2_decap_8 FILLER_50_1341 ();
 sg13g2_decap_8 FILLER_50_1348 ();
 sg13g2_decap_8 FILLER_50_1355 ();
 sg13g2_decap_8 FILLER_50_1362 ();
 sg13g2_decap_8 FILLER_50_1369 ();
 sg13g2_decap_8 FILLER_50_1376 ();
 sg13g2_decap_8 FILLER_50_1383 ();
 sg13g2_decap_8 FILLER_50_1390 ();
 sg13g2_decap_8 FILLER_50_1397 ();
 sg13g2_decap_8 FILLER_50_1404 ();
 sg13g2_decap_8 FILLER_50_1411 ();
 sg13g2_decap_8 FILLER_50_1418 ();
 sg13g2_decap_8 FILLER_50_1425 ();
 sg13g2_decap_8 FILLER_50_1432 ();
 sg13g2_decap_8 FILLER_50_1439 ();
 sg13g2_decap_8 FILLER_50_1446 ();
 sg13g2_decap_8 FILLER_50_1453 ();
 sg13g2_decap_8 FILLER_50_1460 ();
 sg13g2_decap_8 FILLER_50_1467 ();
 sg13g2_decap_8 FILLER_50_1474 ();
 sg13g2_decap_8 FILLER_50_1481 ();
 sg13g2_decap_8 FILLER_50_1488 ();
 sg13g2_decap_8 FILLER_50_1495 ();
 sg13g2_decap_8 FILLER_50_1502 ();
 sg13g2_decap_8 FILLER_50_1509 ();
 sg13g2_decap_8 FILLER_50_1516 ();
 sg13g2_decap_8 FILLER_50_1523 ();
 sg13g2_decap_8 FILLER_50_1530 ();
 sg13g2_decap_8 FILLER_50_1537 ();
 sg13g2_decap_8 FILLER_50_1544 ();
 sg13g2_decap_8 FILLER_50_1551 ();
 sg13g2_decap_8 FILLER_50_1558 ();
 sg13g2_decap_8 FILLER_50_1565 ();
 sg13g2_decap_8 FILLER_50_1572 ();
 sg13g2_decap_8 FILLER_50_1579 ();
 sg13g2_decap_8 FILLER_50_1586 ();
 sg13g2_decap_8 FILLER_50_1593 ();
 sg13g2_decap_8 FILLER_50_1600 ();
 sg13g2_decap_8 FILLER_50_1607 ();
 sg13g2_decap_8 FILLER_50_1614 ();
 sg13g2_decap_8 FILLER_50_1621 ();
 sg13g2_decap_8 FILLER_50_1628 ();
 sg13g2_decap_8 FILLER_50_1635 ();
 sg13g2_decap_8 FILLER_50_1642 ();
 sg13g2_decap_8 FILLER_50_1649 ();
 sg13g2_decap_8 FILLER_50_1656 ();
 sg13g2_decap_8 FILLER_50_1663 ();
 sg13g2_decap_8 FILLER_50_1670 ();
 sg13g2_decap_8 FILLER_50_1677 ();
 sg13g2_decap_8 FILLER_50_1684 ();
 sg13g2_decap_8 FILLER_50_1691 ();
 sg13g2_decap_8 FILLER_50_1698 ();
 sg13g2_decap_8 FILLER_50_1705 ();
 sg13g2_decap_8 FILLER_50_1712 ();
 sg13g2_decap_8 FILLER_50_1719 ();
 sg13g2_decap_8 FILLER_50_1726 ();
 sg13g2_decap_8 FILLER_50_1733 ();
 sg13g2_decap_8 FILLER_50_1740 ();
 sg13g2_decap_8 FILLER_50_1747 ();
 sg13g2_decap_8 FILLER_50_1754 ();
 sg13g2_decap_8 FILLER_50_1761 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_35 ();
 sg13g2_fill_2 FILLER_51_42 ();
 sg13g2_fill_1 FILLER_51_81 ();
 sg13g2_fill_2 FILLER_51_112 ();
 sg13g2_fill_1 FILLER_51_114 ();
 sg13g2_fill_1 FILLER_51_124 ();
 sg13g2_fill_2 FILLER_51_129 ();
 sg13g2_fill_1 FILLER_51_131 ();
 sg13g2_fill_2 FILLER_51_145 ();
 sg13g2_fill_1 FILLER_51_147 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_fill_2 FILLER_51_161 ();
 sg13g2_fill_2 FILLER_51_169 ();
 sg13g2_fill_1 FILLER_51_171 ();
 sg13g2_fill_1 FILLER_51_231 ();
 sg13g2_fill_1 FILLER_51_244 ();
 sg13g2_fill_1 FILLER_51_261 ();
 sg13g2_fill_1 FILLER_51_270 ();
 sg13g2_fill_1 FILLER_51_287 ();
 sg13g2_decap_4 FILLER_51_318 ();
 sg13g2_fill_2 FILLER_51_322 ();
 sg13g2_fill_2 FILLER_51_338 ();
 sg13g2_fill_1 FILLER_51_395 ();
 sg13g2_decap_4 FILLER_51_435 ();
 sg13g2_fill_1 FILLER_51_439 ();
 sg13g2_fill_2 FILLER_51_448 ();
 sg13g2_fill_2 FILLER_51_467 ();
 sg13g2_fill_2 FILLER_51_492 ();
 sg13g2_decap_4 FILLER_51_498 ();
 sg13g2_fill_2 FILLER_51_502 ();
 sg13g2_decap_8 FILLER_51_532 ();
 sg13g2_fill_1 FILLER_51_565 ();
 sg13g2_fill_2 FILLER_51_607 ();
 sg13g2_fill_2 FILLER_51_635 ();
 sg13g2_fill_2 FILLER_51_651 ();
 sg13g2_fill_1 FILLER_51_653 ();
 sg13g2_fill_1 FILLER_51_693 ();
 sg13g2_fill_2 FILLER_51_715 ();
 sg13g2_fill_2 FILLER_51_725 ();
 sg13g2_fill_1 FILLER_51_727 ();
 sg13g2_fill_2 FILLER_51_744 ();
 sg13g2_fill_2 FILLER_51_774 ();
 sg13g2_fill_2 FILLER_51_790 ();
 sg13g2_fill_1 FILLER_51_862 ();
 sg13g2_fill_2 FILLER_51_923 ();
 sg13g2_fill_1 FILLER_51_925 ();
 sg13g2_decap_8 FILLER_51_957 ();
 sg13g2_decap_8 FILLER_51_964 ();
 sg13g2_decap_8 FILLER_51_971 ();
 sg13g2_decap_8 FILLER_51_978 ();
 sg13g2_decap_8 FILLER_51_985 ();
 sg13g2_decap_8 FILLER_51_992 ();
 sg13g2_decap_8 FILLER_51_999 ();
 sg13g2_decap_8 FILLER_51_1006 ();
 sg13g2_decap_8 FILLER_51_1013 ();
 sg13g2_decap_8 FILLER_51_1020 ();
 sg13g2_decap_8 FILLER_51_1027 ();
 sg13g2_decap_8 FILLER_51_1034 ();
 sg13g2_decap_8 FILLER_51_1041 ();
 sg13g2_decap_8 FILLER_51_1048 ();
 sg13g2_decap_8 FILLER_51_1055 ();
 sg13g2_decap_8 FILLER_51_1062 ();
 sg13g2_decap_8 FILLER_51_1069 ();
 sg13g2_decap_8 FILLER_51_1076 ();
 sg13g2_decap_8 FILLER_51_1083 ();
 sg13g2_decap_8 FILLER_51_1090 ();
 sg13g2_decap_8 FILLER_51_1097 ();
 sg13g2_decap_8 FILLER_51_1104 ();
 sg13g2_decap_8 FILLER_51_1111 ();
 sg13g2_decap_8 FILLER_51_1118 ();
 sg13g2_decap_8 FILLER_51_1125 ();
 sg13g2_decap_8 FILLER_51_1132 ();
 sg13g2_decap_8 FILLER_51_1139 ();
 sg13g2_decap_8 FILLER_51_1146 ();
 sg13g2_decap_8 FILLER_51_1153 ();
 sg13g2_decap_8 FILLER_51_1160 ();
 sg13g2_decap_8 FILLER_51_1167 ();
 sg13g2_decap_8 FILLER_51_1174 ();
 sg13g2_decap_8 FILLER_51_1181 ();
 sg13g2_decap_8 FILLER_51_1188 ();
 sg13g2_decap_8 FILLER_51_1195 ();
 sg13g2_decap_8 FILLER_51_1202 ();
 sg13g2_decap_8 FILLER_51_1209 ();
 sg13g2_decap_8 FILLER_51_1216 ();
 sg13g2_decap_8 FILLER_51_1223 ();
 sg13g2_decap_8 FILLER_51_1230 ();
 sg13g2_decap_8 FILLER_51_1237 ();
 sg13g2_decap_8 FILLER_51_1244 ();
 sg13g2_decap_8 FILLER_51_1251 ();
 sg13g2_decap_8 FILLER_51_1258 ();
 sg13g2_decap_8 FILLER_51_1265 ();
 sg13g2_decap_8 FILLER_51_1272 ();
 sg13g2_decap_8 FILLER_51_1279 ();
 sg13g2_decap_8 FILLER_51_1286 ();
 sg13g2_decap_8 FILLER_51_1293 ();
 sg13g2_decap_8 FILLER_51_1300 ();
 sg13g2_decap_8 FILLER_51_1307 ();
 sg13g2_decap_8 FILLER_51_1314 ();
 sg13g2_decap_8 FILLER_51_1321 ();
 sg13g2_decap_8 FILLER_51_1328 ();
 sg13g2_decap_8 FILLER_51_1335 ();
 sg13g2_decap_8 FILLER_51_1342 ();
 sg13g2_decap_8 FILLER_51_1349 ();
 sg13g2_decap_8 FILLER_51_1356 ();
 sg13g2_decap_8 FILLER_51_1363 ();
 sg13g2_decap_8 FILLER_51_1370 ();
 sg13g2_decap_8 FILLER_51_1377 ();
 sg13g2_decap_8 FILLER_51_1384 ();
 sg13g2_decap_8 FILLER_51_1391 ();
 sg13g2_decap_8 FILLER_51_1398 ();
 sg13g2_decap_8 FILLER_51_1405 ();
 sg13g2_decap_8 FILLER_51_1412 ();
 sg13g2_decap_8 FILLER_51_1419 ();
 sg13g2_decap_8 FILLER_51_1426 ();
 sg13g2_decap_8 FILLER_51_1433 ();
 sg13g2_decap_8 FILLER_51_1440 ();
 sg13g2_decap_8 FILLER_51_1447 ();
 sg13g2_decap_8 FILLER_51_1454 ();
 sg13g2_decap_8 FILLER_51_1461 ();
 sg13g2_decap_8 FILLER_51_1468 ();
 sg13g2_decap_8 FILLER_51_1475 ();
 sg13g2_decap_8 FILLER_51_1482 ();
 sg13g2_decap_8 FILLER_51_1489 ();
 sg13g2_decap_8 FILLER_51_1496 ();
 sg13g2_decap_8 FILLER_51_1503 ();
 sg13g2_decap_8 FILLER_51_1510 ();
 sg13g2_decap_8 FILLER_51_1517 ();
 sg13g2_decap_8 FILLER_51_1524 ();
 sg13g2_decap_8 FILLER_51_1531 ();
 sg13g2_decap_8 FILLER_51_1538 ();
 sg13g2_decap_8 FILLER_51_1545 ();
 sg13g2_decap_8 FILLER_51_1552 ();
 sg13g2_decap_8 FILLER_51_1559 ();
 sg13g2_decap_8 FILLER_51_1566 ();
 sg13g2_decap_8 FILLER_51_1573 ();
 sg13g2_decap_8 FILLER_51_1580 ();
 sg13g2_decap_8 FILLER_51_1587 ();
 sg13g2_decap_8 FILLER_51_1594 ();
 sg13g2_decap_8 FILLER_51_1601 ();
 sg13g2_decap_8 FILLER_51_1608 ();
 sg13g2_decap_8 FILLER_51_1615 ();
 sg13g2_decap_8 FILLER_51_1622 ();
 sg13g2_decap_8 FILLER_51_1629 ();
 sg13g2_decap_8 FILLER_51_1636 ();
 sg13g2_decap_8 FILLER_51_1643 ();
 sg13g2_decap_8 FILLER_51_1650 ();
 sg13g2_decap_8 FILLER_51_1657 ();
 sg13g2_decap_8 FILLER_51_1664 ();
 sg13g2_decap_8 FILLER_51_1671 ();
 sg13g2_decap_8 FILLER_51_1678 ();
 sg13g2_decap_8 FILLER_51_1685 ();
 sg13g2_decap_8 FILLER_51_1692 ();
 sg13g2_decap_8 FILLER_51_1699 ();
 sg13g2_decap_8 FILLER_51_1706 ();
 sg13g2_decap_8 FILLER_51_1713 ();
 sg13g2_decap_8 FILLER_51_1720 ();
 sg13g2_decap_8 FILLER_51_1727 ();
 sg13g2_decap_8 FILLER_51_1734 ();
 sg13g2_decap_8 FILLER_51_1741 ();
 sg13g2_decap_8 FILLER_51_1748 ();
 sg13g2_decap_8 FILLER_51_1755 ();
 sg13g2_decap_4 FILLER_51_1762 ();
 sg13g2_fill_2 FILLER_51_1766 ();
 sg13g2_fill_1 FILLER_52_115 ();
 sg13g2_fill_2 FILLER_52_120 ();
 sg13g2_fill_1 FILLER_52_122 ();
 sg13g2_fill_2 FILLER_52_131 ();
 sg13g2_fill_1 FILLER_52_163 ();
 sg13g2_fill_1 FILLER_52_182 ();
 sg13g2_decap_8 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_196 ();
 sg13g2_decap_4 FILLER_52_203 ();
 sg13g2_fill_1 FILLER_52_207 ();
 sg13g2_fill_2 FILLER_52_232 ();
 sg13g2_fill_2 FILLER_52_239 ();
 sg13g2_fill_1 FILLER_52_241 ();
 sg13g2_fill_2 FILLER_52_257 ();
 sg13g2_fill_1 FILLER_52_259 ();
 sg13g2_fill_2 FILLER_52_319 ();
 sg13g2_fill_1 FILLER_52_353 ();
 sg13g2_fill_2 FILLER_52_455 ();
 sg13g2_fill_2 FILLER_52_469 ();
 sg13g2_decap_4 FILLER_52_488 ();
 sg13g2_fill_1 FILLER_52_492 ();
 sg13g2_fill_2 FILLER_52_509 ();
 sg13g2_fill_2 FILLER_52_524 ();
 sg13g2_fill_1 FILLER_52_526 ();
 sg13g2_fill_2 FILLER_52_540 ();
 sg13g2_fill_1 FILLER_52_575 ();
 sg13g2_fill_1 FILLER_52_590 ();
 sg13g2_fill_1 FILLER_52_600 ();
 sg13g2_decap_8 FILLER_52_606 ();
 sg13g2_decap_8 FILLER_52_613 ();
 sg13g2_fill_1 FILLER_52_620 ();
 sg13g2_fill_1 FILLER_52_631 ();
 sg13g2_fill_2 FILLER_52_642 ();
 sg13g2_fill_2 FILLER_52_652 ();
 sg13g2_fill_1 FILLER_52_654 ();
 sg13g2_fill_2 FILLER_52_679 ();
 sg13g2_fill_2 FILLER_52_698 ();
 sg13g2_fill_2 FILLER_52_707 ();
 sg13g2_fill_1 FILLER_52_709 ();
 sg13g2_decap_4 FILLER_52_726 ();
 sg13g2_fill_1 FILLER_52_730 ();
 sg13g2_fill_1 FILLER_52_755 ();
 sg13g2_decap_4 FILLER_52_795 ();
 sg13g2_fill_1 FILLER_52_799 ();
 sg13g2_fill_1 FILLER_52_814 ();
 sg13g2_fill_2 FILLER_52_842 ();
 sg13g2_fill_1 FILLER_52_881 ();
 sg13g2_fill_1 FILLER_52_901 ();
 sg13g2_fill_1 FILLER_52_906 ();
 sg13g2_fill_1 FILLER_52_922 ();
 sg13g2_fill_1 FILLER_52_928 ();
 sg13g2_decap_8 FILLER_52_961 ();
 sg13g2_decap_8 FILLER_52_968 ();
 sg13g2_decap_8 FILLER_52_975 ();
 sg13g2_decap_8 FILLER_52_982 ();
 sg13g2_decap_8 FILLER_52_989 ();
 sg13g2_decap_8 FILLER_52_996 ();
 sg13g2_decap_8 FILLER_52_1003 ();
 sg13g2_decap_8 FILLER_52_1010 ();
 sg13g2_decap_8 FILLER_52_1017 ();
 sg13g2_decap_8 FILLER_52_1024 ();
 sg13g2_decap_8 FILLER_52_1031 ();
 sg13g2_decap_8 FILLER_52_1038 ();
 sg13g2_decap_8 FILLER_52_1045 ();
 sg13g2_decap_8 FILLER_52_1052 ();
 sg13g2_decap_8 FILLER_52_1059 ();
 sg13g2_decap_8 FILLER_52_1066 ();
 sg13g2_decap_8 FILLER_52_1073 ();
 sg13g2_decap_8 FILLER_52_1080 ();
 sg13g2_decap_8 FILLER_52_1087 ();
 sg13g2_decap_8 FILLER_52_1094 ();
 sg13g2_decap_8 FILLER_52_1101 ();
 sg13g2_decap_8 FILLER_52_1108 ();
 sg13g2_decap_8 FILLER_52_1115 ();
 sg13g2_decap_8 FILLER_52_1122 ();
 sg13g2_decap_8 FILLER_52_1129 ();
 sg13g2_decap_8 FILLER_52_1136 ();
 sg13g2_decap_8 FILLER_52_1143 ();
 sg13g2_decap_8 FILLER_52_1150 ();
 sg13g2_decap_8 FILLER_52_1157 ();
 sg13g2_decap_8 FILLER_52_1164 ();
 sg13g2_decap_8 FILLER_52_1171 ();
 sg13g2_decap_8 FILLER_52_1178 ();
 sg13g2_decap_8 FILLER_52_1185 ();
 sg13g2_decap_8 FILLER_52_1192 ();
 sg13g2_decap_8 FILLER_52_1199 ();
 sg13g2_decap_8 FILLER_52_1206 ();
 sg13g2_decap_8 FILLER_52_1213 ();
 sg13g2_decap_8 FILLER_52_1220 ();
 sg13g2_decap_8 FILLER_52_1227 ();
 sg13g2_decap_8 FILLER_52_1234 ();
 sg13g2_decap_8 FILLER_52_1241 ();
 sg13g2_decap_8 FILLER_52_1248 ();
 sg13g2_decap_8 FILLER_52_1255 ();
 sg13g2_decap_8 FILLER_52_1262 ();
 sg13g2_decap_8 FILLER_52_1269 ();
 sg13g2_decap_8 FILLER_52_1276 ();
 sg13g2_decap_8 FILLER_52_1283 ();
 sg13g2_decap_8 FILLER_52_1290 ();
 sg13g2_decap_8 FILLER_52_1297 ();
 sg13g2_decap_8 FILLER_52_1304 ();
 sg13g2_decap_8 FILLER_52_1311 ();
 sg13g2_decap_8 FILLER_52_1318 ();
 sg13g2_decap_8 FILLER_52_1325 ();
 sg13g2_decap_8 FILLER_52_1332 ();
 sg13g2_decap_8 FILLER_52_1339 ();
 sg13g2_decap_8 FILLER_52_1346 ();
 sg13g2_decap_8 FILLER_52_1353 ();
 sg13g2_decap_8 FILLER_52_1360 ();
 sg13g2_decap_8 FILLER_52_1367 ();
 sg13g2_decap_8 FILLER_52_1374 ();
 sg13g2_decap_8 FILLER_52_1381 ();
 sg13g2_decap_8 FILLER_52_1388 ();
 sg13g2_decap_8 FILLER_52_1395 ();
 sg13g2_decap_8 FILLER_52_1402 ();
 sg13g2_decap_8 FILLER_52_1409 ();
 sg13g2_decap_8 FILLER_52_1416 ();
 sg13g2_decap_8 FILLER_52_1423 ();
 sg13g2_decap_8 FILLER_52_1430 ();
 sg13g2_decap_8 FILLER_52_1437 ();
 sg13g2_decap_8 FILLER_52_1444 ();
 sg13g2_decap_8 FILLER_52_1451 ();
 sg13g2_decap_8 FILLER_52_1458 ();
 sg13g2_decap_8 FILLER_52_1465 ();
 sg13g2_decap_8 FILLER_52_1472 ();
 sg13g2_decap_8 FILLER_52_1479 ();
 sg13g2_decap_8 FILLER_52_1486 ();
 sg13g2_decap_8 FILLER_52_1493 ();
 sg13g2_decap_8 FILLER_52_1500 ();
 sg13g2_decap_8 FILLER_52_1507 ();
 sg13g2_decap_8 FILLER_52_1514 ();
 sg13g2_decap_8 FILLER_52_1521 ();
 sg13g2_decap_8 FILLER_52_1528 ();
 sg13g2_decap_8 FILLER_52_1535 ();
 sg13g2_decap_8 FILLER_52_1542 ();
 sg13g2_decap_8 FILLER_52_1549 ();
 sg13g2_decap_8 FILLER_52_1556 ();
 sg13g2_decap_8 FILLER_52_1563 ();
 sg13g2_decap_8 FILLER_52_1570 ();
 sg13g2_decap_8 FILLER_52_1577 ();
 sg13g2_decap_8 FILLER_52_1584 ();
 sg13g2_decap_8 FILLER_52_1591 ();
 sg13g2_decap_8 FILLER_52_1598 ();
 sg13g2_decap_8 FILLER_52_1605 ();
 sg13g2_decap_8 FILLER_52_1612 ();
 sg13g2_decap_8 FILLER_52_1619 ();
 sg13g2_decap_8 FILLER_52_1626 ();
 sg13g2_decap_8 FILLER_52_1633 ();
 sg13g2_decap_8 FILLER_52_1640 ();
 sg13g2_decap_8 FILLER_52_1647 ();
 sg13g2_decap_8 FILLER_52_1654 ();
 sg13g2_decap_8 FILLER_52_1661 ();
 sg13g2_decap_8 FILLER_52_1668 ();
 sg13g2_decap_8 FILLER_52_1675 ();
 sg13g2_decap_8 FILLER_52_1682 ();
 sg13g2_decap_8 FILLER_52_1689 ();
 sg13g2_decap_8 FILLER_52_1696 ();
 sg13g2_decap_8 FILLER_52_1703 ();
 sg13g2_decap_8 FILLER_52_1710 ();
 sg13g2_decap_8 FILLER_52_1717 ();
 sg13g2_decap_8 FILLER_52_1724 ();
 sg13g2_decap_8 FILLER_52_1731 ();
 sg13g2_decap_8 FILLER_52_1738 ();
 sg13g2_decap_8 FILLER_52_1745 ();
 sg13g2_decap_8 FILLER_52_1752 ();
 sg13g2_decap_8 FILLER_52_1759 ();
 sg13g2_fill_2 FILLER_52_1766 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_9 ();
 sg13g2_fill_1 FILLER_53_73 ();
 sg13g2_fill_1 FILLER_53_83 ();
 sg13g2_fill_2 FILLER_53_132 ();
 sg13g2_fill_1 FILLER_53_134 ();
 sg13g2_decap_4 FILLER_53_157 ();
 sg13g2_decap_4 FILLER_53_179 ();
 sg13g2_decap_8 FILLER_53_197 ();
 sg13g2_decap_4 FILLER_53_204 ();
 sg13g2_fill_1 FILLER_53_208 ();
 sg13g2_decap_8 FILLER_53_261 ();
 sg13g2_fill_2 FILLER_53_268 ();
 sg13g2_fill_1 FILLER_53_270 ();
 sg13g2_fill_2 FILLER_53_281 ();
 sg13g2_fill_1 FILLER_53_283 ();
 sg13g2_fill_2 FILLER_53_308 ();
 sg13g2_decap_8 FILLER_53_371 ();
 sg13g2_fill_2 FILLER_53_378 ();
 sg13g2_fill_1 FILLER_53_389 ();
 sg13g2_fill_2 FILLER_53_403 ();
 sg13g2_fill_1 FILLER_53_412 ();
 sg13g2_fill_2 FILLER_53_429 ();
 sg13g2_fill_2 FILLER_53_452 ();
 sg13g2_fill_2 FILLER_53_460 ();
 sg13g2_fill_1 FILLER_53_462 ();
 sg13g2_decap_8 FILLER_53_477 ();
 sg13g2_fill_2 FILLER_53_484 ();
 sg13g2_fill_1 FILLER_53_486 ();
 sg13g2_fill_2 FILLER_53_498 ();
 sg13g2_fill_1 FILLER_53_504 ();
 sg13g2_fill_2 FILLER_53_519 ();
 sg13g2_fill_1 FILLER_53_521 ();
 sg13g2_fill_2 FILLER_53_533 ();
 sg13g2_fill_1 FILLER_53_539 ();
 sg13g2_fill_1 FILLER_53_555 ();
 sg13g2_fill_1 FILLER_53_566 ();
 sg13g2_fill_2 FILLER_53_579 ();
 sg13g2_fill_2 FILLER_53_600 ();
 sg13g2_fill_2 FILLER_53_676 ();
 sg13g2_fill_2 FILLER_53_790 ();
 sg13g2_decap_8 FILLER_53_800 ();
 sg13g2_fill_2 FILLER_53_807 ();
 sg13g2_fill_2 FILLER_53_826 ();
 sg13g2_fill_1 FILLER_53_828 ();
 sg13g2_decap_4 FILLER_53_841 ();
 sg13g2_fill_2 FILLER_53_845 ();
 sg13g2_fill_1 FILLER_53_854 ();
 sg13g2_fill_2 FILLER_53_892 ();
 sg13g2_fill_1 FILLER_53_924 ();
 sg13g2_fill_2 FILLER_53_948 ();
 sg13g2_decap_8 FILLER_53_967 ();
 sg13g2_decap_8 FILLER_53_974 ();
 sg13g2_decap_8 FILLER_53_981 ();
 sg13g2_decap_8 FILLER_53_988 ();
 sg13g2_decap_8 FILLER_53_995 ();
 sg13g2_decap_8 FILLER_53_1002 ();
 sg13g2_decap_8 FILLER_53_1009 ();
 sg13g2_decap_8 FILLER_53_1016 ();
 sg13g2_decap_8 FILLER_53_1023 ();
 sg13g2_decap_8 FILLER_53_1030 ();
 sg13g2_decap_8 FILLER_53_1037 ();
 sg13g2_decap_8 FILLER_53_1044 ();
 sg13g2_decap_8 FILLER_53_1051 ();
 sg13g2_decap_8 FILLER_53_1058 ();
 sg13g2_decap_8 FILLER_53_1065 ();
 sg13g2_decap_8 FILLER_53_1072 ();
 sg13g2_decap_8 FILLER_53_1079 ();
 sg13g2_decap_8 FILLER_53_1086 ();
 sg13g2_decap_8 FILLER_53_1093 ();
 sg13g2_decap_8 FILLER_53_1100 ();
 sg13g2_decap_8 FILLER_53_1107 ();
 sg13g2_decap_8 FILLER_53_1114 ();
 sg13g2_decap_8 FILLER_53_1121 ();
 sg13g2_decap_8 FILLER_53_1128 ();
 sg13g2_decap_8 FILLER_53_1135 ();
 sg13g2_decap_8 FILLER_53_1142 ();
 sg13g2_decap_8 FILLER_53_1149 ();
 sg13g2_decap_8 FILLER_53_1156 ();
 sg13g2_decap_8 FILLER_53_1163 ();
 sg13g2_decap_8 FILLER_53_1170 ();
 sg13g2_decap_8 FILLER_53_1177 ();
 sg13g2_decap_8 FILLER_53_1184 ();
 sg13g2_decap_8 FILLER_53_1191 ();
 sg13g2_decap_8 FILLER_53_1198 ();
 sg13g2_decap_8 FILLER_53_1205 ();
 sg13g2_decap_8 FILLER_53_1212 ();
 sg13g2_decap_8 FILLER_53_1219 ();
 sg13g2_decap_8 FILLER_53_1226 ();
 sg13g2_decap_8 FILLER_53_1233 ();
 sg13g2_decap_8 FILLER_53_1240 ();
 sg13g2_decap_8 FILLER_53_1247 ();
 sg13g2_decap_8 FILLER_53_1254 ();
 sg13g2_decap_8 FILLER_53_1261 ();
 sg13g2_decap_8 FILLER_53_1268 ();
 sg13g2_decap_8 FILLER_53_1275 ();
 sg13g2_decap_8 FILLER_53_1282 ();
 sg13g2_decap_8 FILLER_53_1289 ();
 sg13g2_decap_8 FILLER_53_1296 ();
 sg13g2_decap_8 FILLER_53_1303 ();
 sg13g2_decap_8 FILLER_53_1310 ();
 sg13g2_decap_8 FILLER_53_1317 ();
 sg13g2_decap_8 FILLER_53_1324 ();
 sg13g2_decap_8 FILLER_53_1331 ();
 sg13g2_decap_8 FILLER_53_1338 ();
 sg13g2_decap_8 FILLER_53_1345 ();
 sg13g2_decap_8 FILLER_53_1352 ();
 sg13g2_decap_8 FILLER_53_1359 ();
 sg13g2_decap_8 FILLER_53_1366 ();
 sg13g2_decap_8 FILLER_53_1373 ();
 sg13g2_decap_8 FILLER_53_1380 ();
 sg13g2_decap_8 FILLER_53_1387 ();
 sg13g2_decap_8 FILLER_53_1394 ();
 sg13g2_decap_8 FILLER_53_1401 ();
 sg13g2_decap_8 FILLER_53_1408 ();
 sg13g2_decap_8 FILLER_53_1415 ();
 sg13g2_decap_8 FILLER_53_1422 ();
 sg13g2_decap_8 FILLER_53_1429 ();
 sg13g2_decap_8 FILLER_53_1436 ();
 sg13g2_decap_8 FILLER_53_1443 ();
 sg13g2_decap_8 FILLER_53_1450 ();
 sg13g2_decap_8 FILLER_53_1457 ();
 sg13g2_decap_8 FILLER_53_1464 ();
 sg13g2_decap_8 FILLER_53_1471 ();
 sg13g2_decap_8 FILLER_53_1478 ();
 sg13g2_decap_8 FILLER_53_1485 ();
 sg13g2_decap_8 FILLER_53_1492 ();
 sg13g2_decap_8 FILLER_53_1499 ();
 sg13g2_decap_8 FILLER_53_1506 ();
 sg13g2_decap_8 FILLER_53_1513 ();
 sg13g2_decap_8 FILLER_53_1520 ();
 sg13g2_decap_8 FILLER_53_1527 ();
 sg13g2_decap_8 FILLER_53_1534 ();
 sg13g2_decap_8 FILLER_53_1541 ();
 sg13g2_decap_8 FILLER_53_1548 ();
 sg13g2_decap_8 FILLER_53_1555 ();
 sg13g2_decap_8 FILLER_53_1562 ();
 sg13g2_decap_8 FILLER_53_1569 ();
 sg13g2_decap_8 FILLER_53_1576 ();
 sg13g2_decap_8 FILLER_53_1583 ();
 sg13g2_decap_8 FILLER_53_1590 ();
 sg13g2_decap_8 FILLER_53_1597 ();
 sg13g2_decap_8 FILLER_53_1604 ();
 sg13g2_decap_8 FILLER_53_1611 ();
 sg13g2_decap_8 FILLER_53_1618 ();
 sg13g2_decap_8 FILLER_53_1625 ();
 sg13g2_decap_8 FILLER_53_1632 ();
 sg13g2_decap_8 FILLER_53_1639 ();
 sg13g2_decap_8 FILLER_53_1646 ();
 sg13g2_decap_8 FILLER_53_1653 ();
 sg13g2_decap_8 FILLER_53_1660 ();
 sg13g2_decap_8 FILLER_53_1667 ();
 sg13g2_decap_8 FILLER_53_1674 ();
 sg13g2_decap_8 FILLER_53_1681 ();
 sg13g2_decap_8 FILLER_53_1688 ();
 sg13g2_decap_8 FILLER_53_1695 ();
 sg13g2_decap_8 FILLER_53_1702 ();
 sg13g2_decap_8 FILLER_53_1709 ();
 sg13g2_decap_8 FILLER_53_1716 ();
 sg13g2_decap_8 FILLER_53_1723 ();
 sg13g2_decap_8 FILLER_53_1730 ();
 sg13g2_decap_8 FILLER_53_1737 ();
 sg13g2_decap_8 FILLER_53_1744 ();
 sg13g2_decap_8 FILLER_53_1751 ();
 sg13g2_decap_8 FILLER_53_1758 ();
 sg13g2_fill_2 FILLER_53_1765 ();
 sg13g2_fill_1 FILLER_53_1767 ();
 sg13g2_fill_1 FILLER_54_69 ();
 sg13g2_fill_1 FILLER_54_120 ();
 sg13g2_fill_1 FILLER_54_126 ();
 sg13g2_fill_1 FILLER_54_168 ();
 sg13g2_decap_4 FILLER_54_204 ();
 sg13g2_fill_1 FILLER_54_208 ();
 sg13g2_fill_2 FILLER_54_214 ();
 sg13g2_fill_1 FILLER_54_216 ();
 sg13g2_fill_1 FILLER_54_234 ();
 sg13g2_fill_1 FILLER_54_252 ();
 sg13g2_fill_2 FILLER_54_293 ();
 sg13g2_fill_2 FILLER_54_385 ();
 sg13g2_fill_2 FILLER_54_397 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_fill_1 FILLER_54_409 ();
 sg13g2_fill_1 FILLER_54_424 ();
 sg13g2_fill_1 FILLER_54_453 ();
 sg13g2_decap_4 FILLER_54_469 ();
 sg13g2_fill_2 FILLER_54_473 ();
 sg13g2_fill_2 FILLER_54_480 ();
 sg13g2_fill_1 FILLER_54_482 ();
 sg13g2_decap_4 FILLER_54_503 ();
 sg13g2_fill_2 FILLER_54_507 ();
 sg13g2_fill_2 FILLER_54_525 ();
 sg13g2_fill_1 FILLER_54_527 ();
 sg13g2_fill_1 FILLER_54_581 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_2 FILLER_54_652 ();
 sg13g2_fill_1 FILLER_54_654 ();
 sg13g2_fill_1 FILLER_54_675 ();
 sg13g2_fill_2 FILLER_54_704 ();
 sg13g2_fill_1 FILLER_54_711 ();
 sg13g2_fill_1 FILLER_54_720 ();
 sg13g2_fill_2 FILLER_54_746 ();
 sg13g2_fill_2 FILLER_54_756 ();
 sg13g2_fill_1 FILLER_54_772 ();
 sg13g2_decap_8 FILLER_54_782 ();
 sg13g2_fill_1 FILLER_54_806 ();
 sg13g2_fill_1 FILLER_54_824 ();
 sg13g2_fill_2 FILLER_54_849 ();
 sg13g2_fill_1 FILLER_54_851 ();
 sg13g2_fill_2 FILLER_54_858 ();
 sg13g2_fill_2 FILLER_54_874 ();
 sg13g2_fill_1 FILLER_54_876 ();
 sg13g2_fill_2 FILLER_54_897 ();
 sg13g2_fill_1 FILLER_54_925 ();
 sg13g2_decap_8 FILLER_54_961 ();
 sg13g2_decap_8 FILLER_54_968 ();
 sg13g2_decap_8 FILLER_54_975 ();
 sg13g2_decap_8 FILLER_54_982 ();
 sg13g2_decap_8 FILLER_54_989 ();
 sg13g2_decap_8 FILLER_54_996 ();
 sg13g2_decap_8 FILLER_54_1003 ();
 sg13g2_decap_8 FILLER_54_1010 ();
 sg13g2_decap_8 FILLER_54_1017 ();
 sg13g2_decap_8 FILLER_54_1024 ();
 sg13g2_decap_8 FILLER_54_1031 ();
 sg13g2_decap_8 FILLER_54_1038 ();
 sg13g2_decap_8 FILLER_54_1045 ();
 sg13g2_decap_8 FILLER_54_1052 ();
 sg13g2_decap_8 FILLER_54_1059 ();
 sg13g2_decap_8 FILLER_54_1066 ();
 sg13g2_decap_8 FILLER_54_1073 ();
 sg13g2_decap_8 FILLER_54_1080 ();
 sg13g2_decap_8 FILLER_54_1087 ();
 sg13g2_decap_8 FILLER_54_1094 ();
 sg13g2_decap_8 FILLER_54_1101 ();
 sg13g2_decap_8 FILLER_54_1108 ();
 sg13g2_decap_8 FILLER_54_1115 ();
 sg13g2_decap_8 FILLER_54_1122 ();
 sg13g2_decap_8 FILLER_54_1129 ();
 sg13g2_decap_8 FILLER_54_1136 ();
 sg13g2_decap_8 FILLER_54_1143 ();
 sg13g2_decap_8 FILLER_54_1150 ();
 sg13g2_decap_8 FILLER_54_1157 ();
 sg13g2_decap_8 FILLER_54_1164 ();
 sg13g2_decap_8 FILLER_54_1171 ();
 sg13g2_decap_8 FILLER_54_1178 ();
 sg13g2_decap_8 FILLER_54_1185 ();
 sg13g2_decap_8 FILLER_54_1192 ();
 sg13g2_decap_8 FILLER_54_1199 ();
 sg13g2_decap_8 FILLER_54_1206 ();
 sg13g2_decap_8 FILLER_54_1213 ();
 sg13g2_decap_8 FILLER_54_1220 ();
 sg13g2_decap_8 FILLER_54_1227 ();
 sg13g2_decap_8 FILLER_54_1234 ();
 sg13g2_decap_8 FILLER_54_1241 ();
 sg13g2_decap_8 FILLER_54_1248 ();
 sg13g2_decap_8 FILLER_54_1255 ();
 sg13g2_decap_8 FILLER_54_1262 ();
 sg13g2_decap_8 FILLER_54_1269 ();
 sg13g2_decap_8 FILLER_54_1276 ();
 sg13g2_decap_8 FILLER_54_1283 ();
 sg13g2_decap_8 FILLER_54_1290 ();
 sg13g2_decap_8 FILLER_54_1297 ();
 sg13g2_decap_8 FILLER_54_1304 ();
 sg13g2_decap_8 FILLER_54_1311 ();
 sg13g2_decap_8 FILLER_54_1318 ();
 sg13g2_decap_8 FILLER_54_1325 ();
 sg13g2_decap_8 FILLER_54_1332 ();
 sg13g2_decap_8 FILLER_54_1339 ();
 sg13g2_decap_8 FILLER_54_1346 ();
 sg13g2_decap_8 FILLER_54_1353 ();
 sg13g2_decap_8 FILLER_54_1360 ();
 sg13g2_decap_8 FILLER_54_1367 ();
 sg13g2_decap_8 FILLER_54_1374 ();
 sg13g2_decap_8 FILLER_54_1381 ();
 sg13g2_decap_8 FILLER_54_1388 ();
 sg13g2_decap_8 FILLER_54_1395 ();
 sg13g2_decap_8 FILLER_54_1402 ();
 sg13g2_decap_8 FILLER_54_1409 ();
 sg13g2_decap_8 FILLER_54_1416 ();
 sg13g2_decap_8 FILLER_54_1423 ();
 sg13g2_decap_8 FILLER_54_1430 ();
 sg13g2_decap_8 FILLER_54_1437 ();
 sg13g2_decap_8 FILLER_54_1444 ();
 sg13g2_decap_8 FILLER_54_1451 ();
 sg13g2_decap_8 FILLER_54_1458 ();
 sg13g2_decap_8 FILLER_54_1465 ();
 sg13g2_decap_8 FILLER_54_1472 ();
 sg13g2_decap_8 FILLER_54_1479 ();
 sg13g2_decap_8 FILLER_54_1486 ();
 sg13g2_decap_8 FILLER_54_1493 ();
 sg13g2_decap_8 FILLER_54_1500 ();
 sg13g2_decap_8 FILLER_54_1507 ();
 sg13g2_decap_8 FILLER_54_1514 ();
 sg13g2_decap_8 FILLER_54_1521 ();
 sg13g2_decap_8 FILLER_54_1528 ();
 sg13g2_decap_8 FILLER_54_1535 ();
 sg13g2_decap_8 FILLER_54_1542 ();
 sg13g2_decap_8 FILLER_54_1549 ();
 sg13g2_decap_8 FILLER_54_1556 ();
 sg13g2_decap_8 FILLER_54_1563 ();
 sg13g2_decap_8 FILLER_54_1570 ();
 sg13g2_decap_8 FILLER_54_1577 ();
 sg13g2_decap_8 FILLER_54_1584 ();
 sg13g2_decap_8 FILLER_54_1591 ();
 sg13g2_decap_8 FILLER_54_1598 ();
 sg13g2_decap_8 FILLER_54_1605 ();
 sg13g2_decap_8 FILLER_54_1612 ();
 sg13g2_decap_8 FILLER_54_1619 ();
 sg13g2_decap_8 FILLER_54_1626 ();
 sg13g2_decap_8 FILLER_54_1633 ();
 sg13g2_decap_8 FILLER_54_1640 ();
 sg13g2_decap_8 FILLER_54_1647 ();
 sg13g2_decap_8 FILLER_54_1654 ();
 sg13g2_decap_8 FILLER_54_1661 ();
 sg13g2_decap_8 FILLER_54_1668 ();
 sg13g2_decap_8 FILLER_54_1675 ();
 sg13g2_decap_8 FILLER_54_1682 ();
 sg13g2_decap_8 FILLER_54_1689 ();
 sg13g2_decap_8 FILLER_54_1696 ();
 sg13g2_decap_8 FILLER_54_1703 ();
 sg13g2_decap_8 FILLER_54_1710 ();
 sg13g2_decap_8 FILLER_54_1717 ();
 sg13g2_decap_8 FILLER_54_1724 ();
 sg13g2_decap_8 FILLER_54_1731 ();
 sg13g2_decap_8 FILLER_54_1738 ();
 sg13g2_decap_8 FILLER_54_1745 ();
 sg13g2_decap_8 FILLER_54_1752 ();
 sg13g2_decap_8 FILLER_54_1759 ();
 sg13g2_fill_2 FILLER_54_1766 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_24 ();
 sg13g2_fill_1 FILLER_55_102 ();
 sg13g2_fill_1 FILLER_55_126 ();
 sg13g2_fill_2 FILLER_55_144 ();
 sg13g2_fill_2 FILLER_55_151 ();
 sg13g2_fill_1 FILLER_55_180 ();
 sg13g2_fill_1 FILLER_55_229 ();
 sg13g2_fill_1 FILLER_55_255 ();
 sg13g2_fill_2 FILLER_55_264 ();
 sg13g2_fill_1 FILLER_55_277 ();
 sg13g2_fill_2 FILLER_55_299 ();
 sg13g2_fill_1 FILLER_55_301 ();
 sg13g2_fill_2 FILLER_55_310 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_2 FILLER_55_378 ();
 sg13g2_fill_1 FILLER_55_380 ();
 sg13g2_decap_8 FILLER_55_423 ();
 sg13g2_fill_2 FILLER_55_430 ();
 sg13g2_fill_2 FILLER_55_460 ();
 sg13g2_fill_1 FILLER_55_493 ();
 sg13g2_decap_8 FILLER_55_507 ();
 sg13g2_fill_1 FILLER_55_535 ();
 sg13g2_fill_2 FILLER_55_556 ();
 sg13g2_fill_1 FILLER_55_558 ();
 sg13g2_fill_1 FILLER_55_597 ();
 sg13g2_fill_2 FILLER_55_601 ();
 sg13g2_fill_1 FILLER_55_603 ();
 sg13g2_fill_1 FILLER_55_632 ();
 sg13g2_fill_2 FILLER_55_645 ();
 sg13g2_fill_2 FILLER_55_663 ();
 sg13g2_fill_2 FILLER_55_695 ();
 sg13g2_fill_1 FILLER_55_743 ();
 sg13g2_fill_2 FILLER_55_848 ();
 sg13g2_fill_1 FILLER_55_856 ();
 sg13g2_fill_2 FILLER_55_869 ();
 sg13g2_decap_4 FILLER_55_899 ();
 sg13g2_fill_1 FILLER_55_903 ();
 sg13g2_fill_2 FILLER_55_934 ();
 sg13g2_fill_1 FILLER_55_936 ();
 sg13g2_decap_8 FILLER_55_966 ();
 sg13g2_decap_8 FILLER_55_973 ();
 sg13g2_decap_8 FILLER_55_980 ();
 sg13g2_decap_8 FILLER_55_987 ();
 sg13g2_decap_8 FILLER_55_994 ();
 sg13g2_decap_8 FILLER_55_1001 ();
 sg13g2_decap_8 FILLER_55_1008 ();
 sg13g2_decap_8 FILLER_55_1015 ();
 sg13g2_decap_8 FILLER_55_1022 ();
 sg13g2_decap_8 FILLER_55_1029 ();
 sg13g2_decap_8 FILLER_55_1036 ();
 sg13g2_decap_8 FILLER_55_1043 ();
 sg13g2_decap_8 FILLER_55_1050 ();
 sg13g2_decap_8 FILLER_55_1057 ();
 sg13g2_decap_8 FILLER_55_1064 ();
 sg13g2_decap_8 FILLER_55_1071 ();
 sg13g2_decap_8 FILLER_55_1078 ();
 sg13g2_decap_8 FILLER_55_1085 ();
 sg13g2_decap_8 FILLER_55_1092 ();
 sg13g2_decap_8 FILLER_55_1099 ();
 sg13g2_decap_8 FILLER_55_1106 ();
 sg13g2_decap_8 FILLER_55_1113 ();
 sg13g2_decap_8 FILLER_55_1120 ();
 sg13g2_decap_8 FILLER_55_1127 ();
 sg13g2_decap_8 FILLER_55_1134 ();
 sg13g2_decap_8 FILLER_55_1141 ();
 sg13g2_decap_8 FILLER_55_1148 ();
 sg13g2_decap_8 FILLER_55_1155 ();
 sg13g2_decap_8 FILLER_55_1162 ();
 sg13g2_decap_8 FILLER_55_1169 ();
 sg13g2_decap_8 FILLER_55_1176 ();
 sg13g2_decap_8 FILLER_55_1183 ();
 sg13g2_decap_8 FILLER_55_1190 ();
 sg13g2_decap_8 FILLER_55_1197 ();
 sg13g2_decap_8 FILLER_55_1204 ();
 sg13g2_decap_8 FILLER_55_1211 ();
 sg13g2_decap_8 FILLER_55_1218 ();
 sg13g2_decap_8 FILLER_55_1225 ();
 sg13g2_decap_8 FILLER_55_1232 ();
 sg13g2_decap_8 FILLER_55_1239 ();
 sg13g2_decap_8 FILLER_55_1246 ();
 sg13g2_decap_8 FILLER_55_1253 ();
 sg13g2_decap_8 FILLER_55_1260 ();
 sg13g2_decap_8 FILLER_55_1267 ();
 sg13g2_decap_8 FILLER_55_1274 ();
 sg13g2_decap_8 FILLER_55_1281 ();
 sg13g2_decap_8 FILLER_55_1288 ();
 sg13g2_decap_8 FILLER_55_1295 ();
 sg13g2_decap_8 FILLER_55_1302 ();
 sg13g2_decap_8 FILLER_55_1309 ();
 sg13g2_decap_8 FILLER_55_1316 ();
 sg13g2_decap_8 FILLER_55_1323 ();
 sg13g2_decap_8 FILLER_55_1330 ();
 sg13g2_decap_8 FILLER_55_1337 ();
 sg13g2_decap_8 FILLER_55_1344 ();
 sg13g2_decap_8 FILLER_55_1351 ();
 sg13g2_decap_8 FILLER_55_1358 ();
 sg13g2_decap_8 FILLER_55_1365 ();
 sg13g2_decap_8 FILLER_55_1372 ();
 sg13g2_decap_8 FILLER_55_1379 ();
 sg13g2_decap_8 FILLER_55_1386 ();
 sg13g2_decap_8 FILLER_55_1393 ();
 sg13g2_decap_8 FILLER_55_1400 ();
 sg13g2_decap_8 FILLER_55_1407 ();
 sg13g2_decap_8 FILLER_55_1414 ();
 sg13g2_decap_8 FILLER_55_1421 ();
 sg13g2_decap_8 FILLER_55_1428 ();
 sg13g2_decap_8 FILLER_55_1435 ();
 sg13g2_decap_8 FILLER_55_1442 ();
 sg13g2_decap_8 FILLER_55_1449 ();
 sg13g2_decap_8 FILLER_55_1456 ();
 sg13g2_decap_8 FILLER_55_1463 ();
 sg13g2_decap_8 FILLER_55_1470 ();
 sg13g2_decap_8 FILLER_55_1477 ();
 sg13g2_decap_8 FILLER_55_1484 ();
 sg13g2_decap_8 FILLER_55_1491 ();
 sg13g2_decap_8 FILLER_55_1498 ();
 sg13g2_decap_8 FILLER_55_1505 ();
 sg13g2_decap_8 FILLER_55_1512 ();
 sg13g2_decap_8 FILLER_55_1519 ();
 sg13g2_decap_8 FILLER_55_1526 ();
 sg13g2_decap_8 FILLER_55_1533 ();
 sg13g2_decap_8 FILLER_55_1540 ();
 sg13g2_decap_8 FILLER_55_1547 ();
 sg13g2_decap_8 FILLER_55_1554 ();
 sg13g2_decap_8 FILLER_55_1561 ();
 sg13g2_decap_8 FILLER_55_1568 ();
 sg13g2_decap_8 FILLER_55_1575 ();
 sg13g2_decap_8 FILLER_55_1582 ();
 sg13g2_decap_8 FILLER_55_1589 ();
 sg13g2_decap_8 FILLER_55_1596 ();
 sg13g2_decap_8 FILLER_55_1603 ();
 sg13g2_decap_8 FILLER_55_1610 ();
 sg13g2_decap_8 FILLER_55_1617 ();
 sg13g2_decap_8 FILLER_55_1624 ();
 sg13g2_decap_8 FILLER_55_1631 ();
 sg13g2_decap_8 FILLER_55_1638 ();
 sg13g2_decap_8 FILLER_55_1645 ();
 sg13g2_decap_8 FILLER_55_1652 ();
 sg13g2_decap_8 FILLER_55_1659 ();
 sg13g2_decap_8 FILLER_55_1666 ();
 sg13g2_decap_8 FILLER_55_1673 ();
 sg13g2_decap_8 FILLER_55_1680 ();
 sg13g2_decap_8 FILLER_55_1687 ();
 sg13g2_decap_8 FILLER_55_1694 ();
 sg13g2_decap_8 FILLER_55_1701 ();
 sg13g2_decap_8 FILLER_55_1708 ();
 sg13g2_decap_8 FILLER_55_1715 ();
 sg13g2_decap_8 FILLER_55_1722 ();
 sg13g2_decap_8 FILLER_55_1729 ();
 sg13g2_decap_8 FILLER_55_1736 ();
 sg13g2_decap_8 FILLER_55_1743 ();
 sg13g2_decap_8 FILLER_55_1750 ();
 sg13g2_decap_8 FILLER_55_1757 ();
 sg13g2_decap_4 FILLER_55_1764 ();
 sg13g2_fill_2 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_47 ();
 sg13g2_fill_1 FILLER_56_140 ();
 sg13g2_fill_2 FILLER_56_212 ();
 sg13g2_decap_4 FILLER_56_232 ();
 sg13g2_fill_1 FILLER_56_236 ();
 sg13g2_fill_2 FILLER_56_259 ();
 sg13g2_fill_1 FILLER_56_261 ();
 sg13g2_fill_2 FILLER_56_271 ();
 sg13g2_fill_1 FILLER_56_273 ();
 sg13g2_decap_4 FILLER_56_287 ();
 sg13g2_fill_2 FILLER_56_291 ();
 sg13g2_fill_2 FILLER_56_318 ();
 sg13g2_fill_2 FILLER_56_333 ();
 sg13g2_decap_4 FILLER_56_370 ();
 sg13g2_fill_2 FILLER_56_404 ();
 sg13g2_fill_2 FILLER_56_420 ();
 sg13g2_fill_1 FILLER_56_422 ();
 sg13g2_fill_1 FILLER_56_474 ();
 sg13g2_fill_2 FILLER_56_479 ();
 sg13g2_fill_2 FILLER_56_489 ();
 sg13g2_decap_8 FILLER_56_507 ();
 sg13g2_fill_1 FILLER_56_514 ();
 sg13g2_decap_8 FILLER_56_579 ();
 sg13g2_decap_4 FILLER_56_586 ();
 sg13g2_fill_2 FILLER_56_602 ();
 sg13g2_fill_2 FILLER_56_608 ();
 sg13g2_fill_2 FILLER_56_625 ();
 sg13g2_fill_1 FILLER_56_633 ();
 sg13g2_decap_4 FILLER_56_648 ();
 sg13g2_fill_1 FILLER_56_652 ();
 sg13g2_decap_8 FILLER_56_658 ();
 sg13g2_decap_4 FILLER_56_723 ();
 sg13g2_decap_4 FILLER_56_734 ();
 sg13g2_fill_1 FILLER_56_738 ();
 sg13g2_fill_1 FILLER_56_764 ();
 sg13g2_decap_4 FILLER_56_779 ();
 sg13g2_fill_2 FILLER_56_783 ();
 sg13g2_decap_4 FILLER_56_798 ();
 sg13g2_fill_2 FILLER_56_802 ();
 sg13g2_fill_1 FILLER_56_813 ();
 sg13g2_fill_1 FILLER_56_845 ();
 sg13g2_fill_1 FILLER_56_877 ();
 sg13g2_fill_2 FILLER_56_888 ();
 sg13g2_fill_2 FILLER_56_916 ();
 sg13g2_fill_1 FILLER_56_918 ();
 sg13g2_decap_8 FILLER_56_951 ();
 sg13g2_decap_4 FILLER_56_958 ();
 sg13g2_fill_2 FILLER_56_962 ();
 sg13g2_decap_8 FILLER_56_973 ();
 sg13g2_decap_8 FILLER_56_980 ();
 sg13g2_decap_8 FILLER_56_987 ();
 sg13g2_decap_8 FILLER_56_994 ();
 sg13g2_decap_8 FILLER_56_1001 ();
 sg13g2_decap_8 FILLER_56_1008 ();
 sg13g2_decap_8 FILLER_56_1015 ();
 sg13g2_decap_8 FILLER_56_1022 ();
 sg13g2_decap_8 FILLER_56_1029 ();
 sg13g2_decap_8 FILLER_56_1036 ();
 sg13g2_decap_8 FILLER_56_1043 ();
 sg13g2_decap_8 FILLER_56_1050 ();
 sg13g2_decap_8 FILLER_56_1057 ();
 sg13g2_decap_8 FILLER_56_1064 ();
 sg13g2_decap_8 FILLER_56_1071 ();
 sg13g2_decap_8 FILLER_56_1078 ();
 sg13g2_decap_8 FILLER_56_1085 ();
 sg13g2_decap_8 FILLER_56_1092 ();
 sg13g2_decap_8 FILLER_56_1099 ();
 sg13g2_decap_8 FILLER_56_1106 ();
 sg13g2_decap_8 FILLER_56_1113 ();
 sg13g2_decap_8 FILLER_56_1120 ();
 sg13g2_decap_8 FILLER_56_1127 ();
 sg13g2_decap_8 FILLER_56_1134 ();
 sg13g2_decap_8 FILLER_56_1141 ();
 sg13g2_decap_8 FILLER_56_1148 ();
 sg13g2_decap_8 FILLER_56_1155 ();
 sg13g2_decap_8 FILLER_56_1162 ();
 sg13g2_decap_8 FILLER_56_1169 ();
 sg13g2_decap_8 FILLER_56_1176 ();
 sg13g2_decap_8 FILLER_56_1183 ();
 sg13g2_decap_8 FILLER_56_1190 ();
 sg13g2_decap_8 FILLER_56_1197 ();
 sg13g2_decap_8 FILLER_56_1204 ();
 sg13g2_decap_8 FILLER_56_1211 ();
 sg13g2_decap_8 FILLER_56_1218 ();
 sg13g2_decap_8 FILLER_56_1225 ();
 sg13g2_decap_8 FILLER_56_1232 ();
 sg13g2_decap_8 FILLER_56_1239 ();
 sg13g2_decap_8 FILLER_56_1246 ();
 sg13g2_decap_8 FILLER_56_1253 ();
 sg13g2_decap_8 FILLER_56_1260 ();
 sg13g2_decap_8 FILLER_56_1267 ();
 sg13g2_decap_8 FILLER_56_1274 ();
 sg13g2_decap_8 FILLER_56_1281 ();
 sg13g2_decap_8 FILLER_56_1288 ();
 sg13g2_decap_8 FILLER_56_1295 ();
 sg13g2_decap_8 FILLER_56_1302 ();
 sg13g2_decap_8 FILLER_56_1309 ();
 sg13g2_decap_8 FILLER_56_1316 ();
 sg13g2_decap_8 FILLER_56_1323 ();
 sg13g2_decap_8 FILLER_56_1330 ();
 sg13g2_decap_8 FILLER_56_1337 ();
 sg13g2_decap_8 FILLER_56_1344 ();
 sg13g2_decap_8 FILLER_56_1351 ();
 sg13g2_decap_8 FILLER_56_1358 ();
 sg13g2_decap_8 FILLER_56_1365 ();
 sg13g2_decap_8 FILLER_56_1372 ();
 sg13g2_decap_8 FILLER_56_1379 ();
 sg13g2_decap_8 FILLER_56_1386 ();
 sg13g2_decap_8 FILLER_56_1393 ();
 sg13g2_decap_8 FILLER_56_1400 ();
 sg13g2_decap_8 FILLER_56_1407 ();
 sg13g2_decap_8 FILLER_56_1414 ();
 sg13g2_decap_8 FILLER_56_1421 ();
 sg13g2_decap_8 FILLER_56_1428 ();
 sg13g2_decap_8 FILLER_56_1435 ();
 sg13g2_decap_8 FILLER_56_1442 ();
 sg13g2_decap_8 FILLER_56_1449 ();
 sg13g2_decap_8 FILLER_56_1456 ();
 sg13g2_decap_8 FILLER_56_1463 ();
 sg13g2_decap_8 FILLER_56_1470 ();
 sg13g2_decap_8 FILLER_56_1477 ();
 sg13g2_decap_8 FILLER_56_1484 ();
 sg13g2_decap_8 FILLER_56_1491 ();
 sg13g2_decap_8 FILLER_56_1498 ();
 sg13g2_decap_8 FILLER_56_1505 ();
 sg13g2_decap_8 FILLER_56_1512 ();
 sg13g2_decap_8 FILLER_56_1519 ();
 sg13g2_decap_8 FILLER_56_1526 ();
 sg13g2_decap_8 FILLER_56_1533 ();
 sg13g2_decap_8 FILLER_56_1540 ();
 sg13g2_decap_8 FILLER_56_1547 ();
 sg13g2_decap_8 FILLER_56_1554 ();
 sg13g2_decap_8 FILLER_56_1561 ();
 sg13g2_decap_8 FILLER_56_1568 ();
 sg13g2_decap_8 FILLER_56_1575 ();
 sg13g2_decap_8 FILLER_56_1582 ();
 sg13g2_decap_8 FILLER_56_1589 ();
 sg13g2_decap_8 FILLER_56_1596 ();
 sg13g2_decap_8 FILLER_56_1603 ();
 sg13g2_decap_8 FILLER_56_1610 ();
 sg13g2_decap_8 FILLER_56_1617 ();
 sg13g2_decap_8 FILLER_56_1624 ();
 sg13g2_decap_8 FILLER_56_1631 ();
 sg13g2_decap_8 FILLER_56_1638 ();
 sg13g2_decap_8 FILLER_56_1645 ();
 sg13g2_decap_8 FILLER_56_1652 ();
 sg13g2_decap_8 FILLER_56_1659 ();
 sg13g2_decap_8 FILLER_56_1666 ();
 sg13g2_decap_8 FILLER_56_1673 ();
 sg13g2_decap_8 FILLER_56_1680 ();
 sg13g2_decap_8 FILLER_56_1687 ();
 sg13g2_decap_8 FILLER_56_1694 ();
 sg13g2_decap_8 FILLER_56_1701 ();
 sg13g2_decap_8 FILLER_56_1708 ();
 sg13g2_decap_8 FILLER_56_1715 ();
 sg13g2_decap_8 FILLER_56_1722 ();
 sg13g2_decap_8 FILLER_56_1729 ();
 sg13g2_decap_8 FILLER_56_1736 ();
 sg13g2_decap_8 FILLER_56_1743 ();
 sg13g2_decap_8 FILLER_56_1750 ();
 sg13g2_decap_8 FILLER_56_1757 ();
 sg13g2_decap_4 FILLER_56_1764 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_4 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_34 ();
 sg13g2_fill_2 FILLER_57_75 ();
 sg13g2_fill_1 FILLER_57_101 ();
 sg13g2_fill_2 FILLER_57_121 ();
 sg13g2_fill_2 FILLER_57_131 ();
 sg13g2_fill_2 FILLER_57_156 ();
 sg13g2_fill_1 FILLER_57_158 ();
 sg13g2_fill_2 FILLER_57_220 ();
 sg13g2_decap_4 FILLER_57_267 ();
 sg13g2_fill_2 FILLER_57_271 ();
 sg13g2_fill_2 FILLER_57_302 ();
 sg13g2_fill_1 FILLER_57_304 ();
 sg13g2_decap_8 FILLER_57_310 ();
 sg13g2_fill_1 FILLER_57_317 ();
 sg13g2_fill_1 FILLER_57_347 ();
 sg13g2_fill_1 FILLER_57_377 ();
 sg13g2_fill_1 FILLER_57_415 ();
 sg13g2_fill_2 FILLER_57_424 ();
 sg13g2_fill_1 FILLER_57_426 ();
 sg13g2_fill_1 FILLER_57_446 ();
 sg13g2_fill_1 FILLER_57_455 ();
 sg13g2_decap_4 FILLER_57_465 ();
 sg13g2_fill_2 FILLER_57_507 ();
 sg13g2_fill_1 FILLER_57_530 ();
 sg13g2_decap_8 FILLER_57_568 ();
 sg13g2_fill_2 FILLER_57_575 ();
 sg13g2_fill_2 FILLER_57_622 ();
 sg13g2_decap_8 FILLER_57_646 ();
 sg13g2_fill_1 FILLER_57_653 ();
 sg13g2_fill_2 FILLER_57_721 ();
 sg13g2_fill_1 FILLER_57_723 ();
 sg13g2_fill_1 FILLER_57_740 ();
 sg13g2_fill_1 FILLER_57_775 ();
 sg13g2_decap_4 FILLER_57_781 ();
 sg13g2_fill_2 FILLER_57_785 ();
 sg13g2_fill_2 FILLER_57_804 ();
 sg13g2_fill_1 FILLER_57_806 ();
 sg13g2_decap_4 FILLER_57_810 ();
 sg13g2_fill_2 FILLER_57_814 ();
 sg13g2_fill_2 FILLER_57_842 ();
 sg13g2_fill_2 FILLER_57_851 ();
 sg13g2_fill_1 FILLER_57_862 ();
 sg13g2_fill_1 FILLER_57_912 ();
 sg13g2_decap_8 FILLER_57_923 ();
 sg13g2_fill_2 FILLER_57_930 ();
 sg13g2_fill_2 FILLER_57_941 ();
 sg13g2_fill_2 FILLER_57_946 ();
 sg13g2_decap_8 FILLER_57_957 ();
 sg13g2_decap_8 FILLER_57_964 ();
 sg13g2_decap_8 FILLER_57_971 ();
 sg13g2_decap_8 FILLER_57_978 ();
 sg13g2_decap_8 FILLER_57_985 ();
 sg13g2_decap_8 FILLER_57_992 ();
 sg13g2_decap_8 FILLER_57_999 ();
 sg13g2_decap_8 FILLER_57_1006 ();
 sg13g2_decap_8 FILLER_57_1013 ();
 sg13g2_decap_8 FILLER_57_1020 ();
 sg13g2_decap_8 FILLER_57_1027 ();
 sg13g2_decap_8 FILLER_57_1034 ();
 sg13g2_fill_2 FILLER_57_1041 ();
 sg13g2_fill_1 FILLER_57_1043 ();
 sg13g2_decap_8 FILLER_57_1059 ();
 sg13g2_decap_8 FILLER_57_1066 ();
 sg13g2_fill_2 FILLER_57_1073 ();
 sg13g2_decap_8 FILLER_57_1101 ();
 sg13g2_decap_8 FILLER_57_1108 ();
 sg13g2_decap_8 FILLER_57_1115 ();
 sg13g2_decap_8 FILLER_57_1122 ();
 sg13g2_decap_8 FILLER_57_1129 ();
 sg13g2_decap_8 FILLER_57_1136 ();
 sg13g2_decap_8 FILLER_57_1143 ();
 sg13g2_decap_8 FILLER_57_1150 ();
 sg13g2_decap_8 FILLER_57_1157 ();
 sg13g2_decap_8 FILLER_57_1164 ();
 sg13g2_decap_8 FILLER_57_1171 ();
 sg13g2_decap_8 FILLER_57_1178 ();
 sg13g2_decap_8 FILLER_57_1185 ();
 sg13g2_decap_8 FILLER_57_1192 ();
 sg13g2_decap_8 FILLER_57_1199 ();
 sg13g2_decap_8 FILLER_57_1206 ();
 sg13g2_decap_8 FILLER_57_1213 ();
 sg13g2_decap_8 FILLER_57_1220 ();
 sg13g2_decap_8 FILLER_57_1227 ();
 sg13g2_decap_8 FILLER_57_1234 ();
 sg13g2_decap_8 FILLER_57_1241 ();
 sg13g2_decap_8 FILLER_57_1248 ();
 sg13g2_decap_8 FILLER_57_1255 ();
 sg13g2_decap_8 FILLER_57_1262 ();
 sg13g2_decap_8 FILLER_57_1269 ();
 sg13g2_decap_8 FILLER_57_1276 ();
 sg13g2_decap_8 FILLER_57_1283 ();
 sg13g2_decap_8 FILLER_57_1290 ();
 sg13g2_decap_8 FILLER_57_1297 ();
 sg13g2_decap_8 FILLER_57_1304 ();
 sg13g2_decap_8 FILLER_57_1311 ();
 sg13g2_decap_8 FILLER_57_1318 ();
 sg13g2_decap_8 FILLER_57_1325 ();
 sg13g2_decap_8 FILLER_57_1332 ();
 sg13g2_decap_8 FILLER_57_1339 ();
 sg13g2_decap_8 FILLER_57_1346 ();
 sg13g2_decap_8 FILLER_57_1353 ();
 sg13g2_decap_8 FILLER_57_1360 ();
 sg13g2_decap_8 FILLER_57_1367 ();
 sg13g2_decap_8 FILLER_57_1374 ();
 sg13g2_decap_8 FILLER_57_1381 ();
 sg13g2_decap_8 FILLER_57_1388 ();
 sg13g2_decap_8 FILLER_57_1395 ();
 sg13g2_decap_8 FILLER_57_1402 ();
 sg13g2_decap_8 FILLER_57_1409 ();
 sg13g2_decap_8 FILLER_57_1416 ();
 sg13g2_decap_8 FILLER_57_1423 ();
 sg13g2_decap_8 FILLER_57_1430 ();
 sg13g2_decap_8 FILLER_57_1437 ();
 sg13g2_decap_8 FILLER_57_1444 ();
 sg13g2_decap_8 FILLER_57_1451 ();
 sg13g2_decap_8 FILLER_57_1458 ();
 sg13g2_decap_8 FILLER_57_1465 ();
 sg13g2_decap_8 FILLER_57_1472 ();
 sg13g2_decap_8 FILLER_57_1479 ();
 sg13g2_decap_8 FILLER_57_1486 ();
 sg13g2_decap_8 FILLER_57_1493 ();
 sg13g2_decap_8 FILLER_57_1500 ();
 sg13g2_decap_8 FILLER_57_1507 ();
 sg13g2_decap_8 FILLER_57_1514 ();
 sg13g2_decap_8 FILLER_57_1521 ();
 sg13g2_decap_8 FILLER_57_1528 ();
 sg13g2_decap_8 FILLER_57_1535 ();
 sg13g2_decap_8 FILLER_57_1542 ();
 sg13g2_decap_8 FILLER_57_1549 ();
 sg13g2_decap_8 FILLER_57_1556 ();
 sg13g2_decap_8 FILLER_57_1563 ();
 sg13g2_decap_8 FILLER_57_1570 ();
 sg13g2_decap_8 FILLER_57_1577 ();
 sg13g2_decap_8 FILLER_57_1584 ();
 sg13g2_decap_8 FILLER_57_1591 ();
 sg13g2_decap_8 FILLER_57_1598 ();
 sg13g2_decap_8 FILLER_57_1605 ();
 sg13g2_decap_8 FILLER_57_1612 ();
 sg13g2_decap_8 FILLER_57_1619 ();
 sg13g2_decap_8 FILLER_57_1626 ();
 sg13g2_decap_8 FILLER_57_1633 ();
 sg13g2_decap_8 FILLER_57_1640 ();
 sg13g2_decap_8 FILLER_57_1647 ();
 sg13g2_decap_8 FILLER_57_1654 ();
 sg13g2_decap_8 FILLER_57_1661 ();
 sg13g2_decap_8 FILLER_57_1668 ();
 sg13g2_decap_8 FILLER_57_1675 ();
 sg13g2_decap_8 FILLER_57_1682 ();
 sg13g2_decap_8 FILLER_57_1689 ();
 sg13g2_decap_8 FILLER_57_1696 ();
 sg13g2_decap_8 FILLER_57_1703 ();
 sg13g2_decap_8 FILLER_57_1710 ();
 sg13g2_decap_8 FILLER_57_1717 ();
 sg13g2_decap_8 FILLER_57_1724 ();
 sg13g2_decap_8 FILLER_57_1731 ();
 sg13g2_decap_8 FILLER_57_1738 ();
 sg13g2_decap_8 FILLER_57_1745 ();
 sg13g2_decap_8 FILLER_57_1752 ();
 sg13g2_decap_8 FILLER_57_1759 ();
 sg13g2_fill_2 FILLER_57_1766 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_fill_2 FILLER_58_28 ();
 sg13g2_fill_1 FILLER_58_30 ();
 sg13g2_fill_1 FILLER_58_70 ();
 sg13g2_fill_1 FILLER_58_136 ();
 sg13g2_fill_1 FILLER_58_260 ();
 sg13g2_fill_2 FILLER_58_269 ();
 sg13g2_fill_1 FILLER_58_271 ();
 sg13g2_fill_1 FILLER_58_311 ();
 sg13g2_fill_2 FILLER_58_347 ();
 sg13g2_fill_1 FILLER_58_375 ();
 sg13g2_fill_2 FILLER_58_384 ();
 sg13g2_fill_2 FILLER_58_443 ();
 sg13g2_fill_2 FILLER_58_458 ();
 sg13g2_decap_4 FILLER_58_476 ();
 sg13g2_fill_1 FILLER_58_480 ();
 sg13g2_fill_2 FILLER_58_485 ();
 sg13g2_decap_8 FILLER_58_504 ();
 sg13g2_decap_4 FILLER_58_511 ();
 sg13g2_fill_2 FILLER_58_526 ();
 sg13g2_fill_1 FILLER_58_528 ();
 sg13g2_fill_1 FILLER_58_535 ();
 sg13g2_fill_2 FILLER_58_588 ();
 sg13g2_fill_2 FILLER_58_653 ();
 sg13g2_fill_2 FILLER_58_671 ();
 sg13g2_decap_4 FILLER_58_683 ();
 sg13g2_fill_2 FILLER_58_697 ();
 sg13g2_fill_1 FILLER_58_699 ();
 sg13g2_fill_2 FILLER_58_705 ();
 sg13g2_fill_1 FILLER_58_707 ();
 sg13g2_fill_2 FILLER_58_734 ();
 sg13g2_fill_2 FILLER_58_767 ();
 sg13g2_fill_1 FILLER_58_769 ();
 sg13g2_fill_2 FILLER_58_831 ();
 sg13g2_fill_1 FILLER_58_833 ();
 sg13g2_fill_1 FILLER_58_848 ();
 sg13g2_fill_1 FILLER_58_877 ();
 sg13g2_decap_8 FILLER_58_939 ();
 sg13g2_decap_4 FILLER_58_946 ();
 sg13g2_fill_2 FILLER_58_950 ();
 sg13g2_decap_8 FILLER_58_980 ();
 sg13g2_decap_8 FILLER_58_987 ();
 sg13g2_decap_8 FILLER_58_994 ();
 sg13g2_fill_2 FILLER_58_1001 ();
 sg13g2_fill_1 FILLER_58_1003 ();
 sg13g2_fill_1 FILLER_58_1017 ();
 sg13g2_decap_8 FILLER_58_1119 ();
 sg13g2_decap_8 FILLER_58_1126 ();
 sg13g2_decap_8 FILLER_58_1133 ();
 sg13g2_decap_8 FILLER_58_1140 ();
 sg13g2_decap_8 FILLER_58_1147 ();
 sg13g2_decap_8 FILLER_58_1154 ();
 sg13g2_decap_8 FILLER_58_1161 ();
 sg13g2_decap_8 FILLER_58_1168 ();
 sg13g2_decap_8 FILLER_58_1175 ();
 sg13g2_decap_8 FILLER_58_1182 ();
 sg13g2_decap_8 FILLER_58_1189 ();
 sg13g2_decap_8 FILLER_58_1196 ();
 sg13g2_decap_8 FILLER_58_1203 ();
 sg13g2_decap_8 FILLER_58_1210 ();
 sg13g2_decap_8 FILLER_58_1217 ();
 sg13g2_decap_8 FILLER_58_1224 ();
 sg13g2_decap_8 FILLER_58_1231 ();
 sg13g2_decap_8 FILLER_58_1238 ();
 sg13g2_decap_8 FILLER_58_1245 ();
 sg13g2_decap_8 FILLER_58_1252 ();
 sg13g2_decap_8 FILLER_58_1259 ();
 sg13g2_decap_8 FILLER_58_1266 ();
 sg13g2_decap_8 FILLER_58_1273 ();
 sg13g2_decap_8 FILLER_58_1280 ();
 sg13g2_decap_8 FILLER_58_1287 ();
 sg13g2_decap_8 FILLER_58_1294 ();
 sg13g2_decap_8 FILLER_58_1301 ();
 sg13g2_decap_8 FILLER_58_1308 ();
 sg13g2_decap_8 FILLER_58_1315 ();
 sg13g2_decap_8 FILLER_58_1322 ();
 sg13g2_decap_8 FILLER_58_1329 ();
 sg13g2_decap_8 FILLER_58_1336 ();
 sg13g2_decap_8 FILLER_58_1343 ();
 sg13g2_decap_8 FILLER_58_1350 ();
 sg13g2_decap_8 FILLER_58_1357 ();
 sg13g2_decap_8 FILLER_58_1364 ();
 sg13g2_decap_8 FILLER_58_1371 ();
 sg13g2_decap_8 FILLER_58_1378 ();
 sg13g2_decap_8 FILLER_58_1385 ();
 sg13g2_decap_8 FILLER_58_1392 ();
 sg13g2_decap_8 FILLER_58_1399 ();
 sg13g2_decap_8 FILLER_58_1406 ();
 sg13g2_decap_8 FILLER_58_1413 ();
 sg13g2_decap_8 FILLER_58_1420 ();
 sg13g2_decap_8 FILLER_58_1427 ();
 sg13g2_decap_8 FILLER_58_1434 ();
 sg13g2_decap_8 FILLER_58_1441 ();
 sg13g2_decap_8 FILLER_58_1448 ();
 sg13g2_decap_8 FILLER_58_1455 ();
 sg13g2_decap_8 FILLER_58_1462 ();
 sg13g2_decap_8 FILLER_58_1469 ();
 sg13g2_decap_8 FILLER_58_1476 ();
 sg13g2_decap_8 FILLER_58_1483 ();
 sg13g2_decap_8 FILLER_58_1490 ();
 sg13g2_decap_8 FILLER_58_1497 ();
 sg13g2_decap_8 FILLER_58_1504 ();
 sg13g2_decap_8 FILLER_58_1511 ();
 sg13g2_decap_8 FILLER_58_1518 ();
 sg13g2_decap_8 FILLER_58_1525 ();
 sg13g2_decap_8 FILLER_58_1532 ();
 sg13g2_decap_8 FILLER_58_1539 ();
 sg13g2_decap_8 FILLER_58_1546 ();
 sg13g2_decap_8 FILLER_58_1553 ();
 sg13g2_decap_8 FILLER_58_1560 ();
 sg13g2_decap_8 FILLER_58_1567 ();
 sg13g2_decap_8 FILLER_58_1574 ();
 sg13g2_decap_8 FILLER_58_1581 ();
 sg13g2_decap_8 FILLER_58_1588 ();
 sg13g2_decap_8 FILLER_58_1595 ();
 sg13g2_decap_8 FILLER_58_1602 ();
 sg13g2_decap_8 FILLER_58_1609 ();
 sg13g2_decap_8 FILLER_58_1616 ();
 sg13g2_decap_8 FILLER_58_1623 ();
 sg13g2_decap_8 FILLER_58_1630 ();
 sg13g2_decap_8 FILLER_58_1637 ();
 sg13g2_decap_8 FILLER_58_1644 ();
 sg13g2_decap_8 FILLER_58_1651 ();
 sg13g2_decap_8 FILLER_58_1658 ();
 sg13g2_decap_8 FILLER_58_1665 ();
 sg13g2_decap_8 FILLER_58_1672 ();
 sg13g2_decap_8 FILLER_58_1679 ();
 sg13g2_decap_8 FILLER_58_1686 ();
 sg13g2_decap_8 FILLER_58_1693 ();
 sg13g2_decap_8 FILLER_58_1700 ();
 sg13g2_decap_8 FILLER_58_1707 ();
 sg13g2_decap_8 FILLER_58_1714 ();
 sg13g2_decap_8 FILLER_58_1721 ();
 sg13g2_decap_8 FILLER_58_1728 ();
 sg13g2_decap_8 FILLER_58_1735 ();
 sg13g2_decap_8 FILLER_58_1742 ();
 sg13g2_decap_8 FILLER_58_1749 ();
 sg13g2_decap_8 FILLER_58_1756 ();
 sg13g2_decap_4 FILLER_58_1763 ();
 sg13g2_fill_1 FILLER_58_1767 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_39 ();
 sg13g2_fill_1 FILLER_59_46 ();
 sg13g2_fill_1 FILLER_59_58 ();
 sg13g2_fill_2 FILLER_59_68 ();
 sg13g2_fill_2 FILLER_59_100 ();
 sg13g2_fill_2 FILLER_59_166 ();
 sg13g2_fill_1 FILLER_59_168 ();
 sg13g2_fill_2 FILLER_59_174 ();
 sg13g2_fill_1 FILLER_59_179 ();
 sg13g2_fill_2 FILLER_59_195 ();
 sg13g2_fill_1 FILLER_59_197 ();
 sg13g2_fill_1 FILLER_59_231 ();
 sg13g2_fill_2 FILLER_59_261 ();
 sg13g2_fill_2 FILLER_59_307 ();
 sg13g2_fill_1 FILLER_59_309 ();
 sg13g2_decap_4 FILLER_59_315 ();
 sg13g2_fill_1 FILLER_59_319 ();
 sg13g2_fill_2 FILLER_59_346 ();
 sg13g2_fill_2 FILLER_59_440 ();
 sg13g2_fill_1 FILLER_59_459 ();
 sg13g2_fill_2 FILLER_59_474 ();
 sg13g2_fill_1 FILLER_59_476 ();
 sg13g2_fill_1 FILLER_59_508 ();
 sg13g2_fill_1 FILLER_59_514 ();
 sg13g2_fill_1 FILLER_59_520 ();
 sg13g2_fill_1 FILLER_59_532 ();
 sg13g2_decap_4 FILLER_59_537 ();
 sg13g2_fill_1 FILLER_59_541 ();
 sg13g2_fill_2 FILLER_59_554 ();
 sg13g2_fill_2 FILLER_59_561 ();
 sg13g2_fill_1 FILLER_59_563 ();
 sg13g2_fill_2 FILLER_59_574 ();
 sg13g2_fill_1 FILLER_59_576 ();
 sg13g2_fill_2 FILLER_59_586 ();
 sg13g2_fill_1 FILLER_59_588 ();
 sg13g2_fill_2 FILLER_59_631 ();
 sg13g2_fill_1 FILLER_59_657 ();
 sg13g2_fill_1 FILLER_59_700 ();
 sg13g2_decap_8 FILLER_59_783 ();
 sg13g2_decap_4 FILLER_59_790 ();
 sg13g2_fill_1 FILLER_59_794 ();
 sg13g2_fill_2 FILLER_59_815 ();
 sg13g2_fill_1 FILLER_59_861 ();
 sg13g2_fill_2 FILLER_59_888 ();
 sg13g2_decap_4 FILLER_59_902 ();
 sg13g2_decap_4 FILLER_59_954 ();
 sg13g2_fill_2 FILLER_59_989 ();
 sg13g2_decap_4 FILLER_59_999 ();
 sg13g2_fill_1 FILLER_59_1003 ();
 sg13g2_fill_2 FILLER_59_1111 ();
 sg13g2_fill_1 FILLER_59_1113 ();
 sg13g2_decap_8 FILLER_59_1140 ();
 sg13g2_decap_8 FILLER_59_1147 ();
 sg13g2_decap_8 FILLER_59_1154 ();
 sg13g2_decap_8 FILLER_59_1161 ();
 sg13g2_decap_8 FILLER_59_1168 ();
 sg13g2_decap_8 FILLER_59_1175 ();
 sg13g2_decap_8 FILLER_59_1182 ();
 sg13g2_decap_8 FILLER_59_1189 ();
 sg13g2_decap_8 FILLER_59_1196 ();
 sg13g2_decap_8 FILLER_59_1203 ();
 sg13g2_decap_8 FILLER_59_1210 ();
 sg13g2_decap_8 FILLER_59_1217 ();
 sg13g2_decap_8 FILLER_59_1224 ();
 sg13g2_decap_8 FILLER_59_1231 ();
 sg13g2_decap_8 FILLER_59_1238 ();
 sg13g2_decap_8 FILLER_59_1245 ();
 sg13g2_decap_8 FILLER_59_1252 ();
 sg13g2_decap_8 FILLER_59_1259 ();
 sg13g2_decap_8 FILLER_59_1266 ();
 sg13g2_decap_8 FILLER_59_1273 ();
 sg13g2_decap_8 FILLER_59_1280 ();
 sg13g2_decap_8 FILLER_59_1287 ();
 sg13g2_decap_8 FILLER_59_1294 ();
 sg13g2_decap_8 FILLER_59_1301 ();
 sg13g2_decap_8 FILLER_59_1308 ();
 sg13g2_decap_8 FILLER_59_1315 ();
 sg13g2_decap_8 FILLER_59_1322 ();
 sg13g2_decap_8 FILLER_59_1329 ();
 sg13g2_decap_8 FILLER_59_1336 ();
 sg13g2_decap_8 FILLER_59_1343 ();
 sg13g2_decap_8 FILLER_59_1350 ();
 sg13g2_decap_8 FILLER_59_1357 ();
 sg13g2_decap_8 FILLER_59_1364 ();
 sg13g2_decap_8 FILLER_59_1371 ();
 sg13g2_decap_8 FILLER_59_1378 ();
 sg13g2_decap_8 FILLER_59_1385 ();
 sg13g2_decap_8 FILLER_59_1392 ();
 sg13g2_decap_8 FILLER_59_1399 ();
 sg13g2_decap_8 FILLER_59_1406 ();
 sg13g2_decap_8 FILLER_59_1413 ();
 sg13g2_decap_8 FILLER_59_1420 ();
 sg13g2_decap_8 FILLER_59_1427 ();
 sg13g2_decap_8 FILLER_59_1434 ();
 sg13g2_decap_8 FILLER_59_1441 ();
 sg13g2_decap_8 FILLER_59_1448 ();
 sg13g2_decap_8 FILLER_59_1455 ();
 sg13g2_decap_8 FILLER_59_1462 ();
 sg13g2_decap_8 FILLER_59_1469 ();
 sg13g2_decap_8 FILLER_59_1476 ();
 sg13g2_decap_8 FILLER_59_1483 ();
 sg13g2_decap_8 FILLER_59_1490 ();
 sg13g2_decap_8 FILLER_59_1497 ();
 sg13g2_decap_8 FILLER_59_1504 ();
 sg13g2_decap_8 FILLER_59_1511 ();
 sg13g2_decap_8 FILLER_59_1518 ();
 sg13g2_decap_8 FILLER_59_1525 ();
 sg13g2_decap_8 FILLER_59_1532 ();
 sg13g2_decap_8 FILLER_59_1539 ();
 sg13g2_decap_8 FILLER_59_1546 ();
 sg13g2_decap_8 FILLER_59_1553 ();
 sg13g2_decap_8 FILLER_59_1560 ();
 sg13g2_decap_8 FILLER_59_1567 ();
 sg13g2_decap_8 FILLER_59_1574 ();
 sg13g2_decap_8 FILLER_59_1581 ();
 sg13g2_decap_8 FILLER_59_1588 ();
 sg13g2_decap_8 FILLER_59_1595 ();
 sg13g2_decap_8 FILLER_59_1602 ();
 sg13g2_decap_8 FILLER_59_1609 ();
 sg13g2_decap_8 FILLER_59_1616 ();
 sg13g2_decap_8 FILLER_59_1623 ();
 sg13g2_decap_8 FILLER_59_1630 ();
 sg13g2_decap_8 FILLER_59_1637 ();
 sg13g2_decap_8 FILLER_59_1644 ();
 sg13g2_decap_8 FILLER_59_1651 ();
 sg13g2_decap_8 FILLER_59_1658 ();
 sg13g2_decap_8 FILLER_59_1665 ();
 sg13g2_decap_8 FILLER_59_1672 ();
 sg13g2_decap_8 FILLER_59_1679 ();
 sg13g2_decap_8 FILLER_59_1686 ();
 sg13g2_decap_8 FILLER_59_1693 ();
 sg13g2_decap_8 FILLER_59_1700 ();
 sg13g2_decap_8 FILLER_59_1707 ();
 sg13g2_decap_8 FILLER_59_1714 ();
 sg13g2_decap_8 FILLER_59_1721 ();
 sg13g2_decap_8 FILLER_59_1728 ();
 sg13g2_decap_8 FILLER_59_1735 ();
 sg13g2_decap_8 FILLER_59_1742 ();
 sg13g2_decap_8 FILLER_59_1749 ();
 sg13g2_decap_8 FILLER_59_1756 ();
 sg13g2_decap_4 FILLER_59_1763 ();
 sg13g2_fill_1 FILLER_59_1767 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_fill_2 FILLER_60_54 ();
 sg13g2_decap_8 FILLER_60_64 ();
 sg13g2_decap_4 FILLER_60_71 ();
 sg13g2_fill_1 FILLER_60_75 ();
 sg13g2_fill_2 FILLER_60_110 ();
 sg13g2_fill_2 FILLER_60_125 ();
 sg13g2_fill_1 FILLER_60_140 ();
 sg13g2_fill_2 FILLER_60_145 ();
 sg13g2_fill_1 FILLER_60_147 ();
 sg13g2_fill_2 FILLER_60_163 ();
 sg13g2_fill_1 FILLER_60_165 ();
 sg13g2_fill_1 FILLER_60_198 ();
 sg13g2_fill_2 FILLER_60_207 ();
 sg13g2_fill_1 FILLER_60_209 ();
 sg13g2_decap_8 FILLER_60_225 ();
 sg13g2_fill_1 FILLER_60_232 ();
 sg13g2_fill_1 FILLER_60_265 ();
 sg13g2_fill_2 FILLER_60_271 ();
 sg13g2_fill_1 FILLER_60_273 ();
 sg13g2_fill_1 FILLER_60_287 ();
 sg13g2_fill_2 FILLER_60_311 ();
 sg13g2_fill_1 FILLER_60_313 ();
 sg13g2_decap_8 FILLER_60_323 ();
 sg13g2_fill_2 FILLER_60_330 ();
 sg13g2_fill_2 FILLER_60_359 ();
 sg13g2_fill_2 FILLER_60_399 ();
 sg13g2_fill_2 FILLER_60_450 ();
 sg13g2_fill_1 FILLER_60_452 ();
 sg13g2_fill_2 FILLER_60_479 ();
 sg13g2_fill_1 FILLER_60_481 ();
 sg13g2_fill_1 FILLER_60_495 ();
 sg13g2_fill_2 FILLER_60_504 ();
 sg13g2_fill_1 FILLER_60_506 ();
 sg13g2_fill_1 FILLER_60_530 ();
 sg13g2_fill_1 FILLER_60_540 ();
 sg13g2_fill_2 FILLER_60_584 ();
 sg13g2_fill_1 FILLER_60_586 ();
 sg13g2_fill_1 FILLER_60_592 ();
 sg13g2_fill_2 FILLER_60_604 ();
 sg13g2_fill_1 FILLER_60_606 ();
 sg13g2_fill_1 FILLER_60_612 ();
 sg13g2_fill_1 FILLER_60_672 ();
 sg13g2_fill_2 FILLER_60_697 ();
 sg13g2_fill_2 FILLER_60_733 ();
 sg13g2_fill_2 FILLER_60_772 ();
 sg13g2_fill_1 FILLER_60_774 ();
 sg13g2_fill_2 FILLER_60_788 ();
 sg13g2_fill_2 FILLER_60_795 ();
 sg13g2_fill_1 FILLER_60_797 ();
 sg13g2_decap_4 FILLER_60_817 ();
 sg13g2_fill_2 FILLER_60_821 ();
 sg13g2_decap_8 FILLER_60_852 ();
 sg13g2_fill_1 FILLER_60_859 ();
 sg13g2_fill_1 FILLER_60_886 ();
 sg13g2_decap_4 FILLER_60_903 ();
 sg13g2_fill_2 FILLER_60_952 ();
 sg13g2_fill_1 FILLER_60_954 ();
 sg13g2_fill_2 FILLER_60_1017 ();
 sg13g2_fill_2 FILLER_60_1101 ();
 sg13g2_fill_1 FILLER_60_1103 ();
 sg13g2_fill_1 FILLER_60_1130 ();
 sg13g2_decap_8 FILLER_60_1150 ();
 sg13g2_decap_8 FILLER_60_1157 ();
 sg13g2_decap_8 FILLER_60_1164 ();
 sg13g2_decap_8 FILLER_60_1171 ();
 sg13g2_decap_8 FILLER_60_1178 ();
 sg13g2_decap_8 FILLER_60_1185 ();
 sg13g2_decap_8 FILLER_60_1192 ();
 sg13g2_decap_8 FILLER_60_1199 ();
 sg13g2_decap_8 FILLER_60_1206 ();
 sg13g2_decap_8 FILLER_60_1213 ();
 sg13g2_decap_8 FILLER_60_1220 ();
 sg13g2_decap_8 FILLER_60_1227 ();
 sg13g2_decap_8 FILLER_60_1234 ();
 sg13g2_decap_8 FILLER_60_1241 ();
 sg13g2_decap_8 FILLER_60_1248 ();
 sg13g2_decap_8 FILLER_60_1255 ();
 sg13g2_decap_8 FILLER_60_1262 ();
 sg13g2_decap_8 FILLER_60_1269 ();
 sg13g2_decap_8 FILLER_60_1276 ();
 sg13g2_decap_8 FILLER_60_1283 ();
 sg13g2_decap_8 FILLER_60_1290 ();
 sg13g2_decap_8 FILLER_60_1297 ();
 sg13g2_decap_8 FILLER_60_1304 ();
 sg13g2_decap_8 FILLER_60_1311 ();
 sg13g2_decap_8 FILLER_60_1318 ();
 sg13g2_decap_8 FILLER_60_1325 ();
 sg13g2_decap_8 FILLER_60_1332 ();
 sg13g2_decap_8 FILLER_60_1339 ();
 sg13g2_decap_8 FILLER_60_1346 ();
 sg13g2_decap_8 FILLER_60_1353 ();
 sg13g2_decap_8 FILLER_60_1360 ();
 sg13g2_decap_8 FILLER_60_1367 ();
 sg13g2_decap_8 FILLER_60_1374 ();
 sg13g2_decap_8 FILLER_60_1381 ();
 sg13g2_decap_8 FILLER_60_1388 ();
 sg13g2_decap_8 FILLER_60_1395 ();
 sg13g2_decap_8 FILLER_60_1402 ();
 sg13g2_decap_8 FILLER_60_1409 ();
 sg13g2_decap_8 FILLER_60_1416 ();
 sg13g2_decap_8 FILLER_60_1423 ();
 sg13g2_decap_8 FILLER_60_1430 ();
 sg13g2_decap_8 FILLER_60_1437 ();
 sg13g2_decap_8 FILLER_60_1444 ();
 sg13g2_decap_8 FILLER_60_1451 ();
 sg13g2_decap_8 FILLER_60_1458 ();
 sg13g2_decap_8 FILLER_60_1465 ();
 sg13g2_decap_8 FILLER_60_1472 ();
 sg13g2_decap_8 FILLER_60_1479 ();
 sg13g2_decap_8 FILLER_60_1486 ();
 sg13g2_decap_8 FILLER_60_1493 ();
 sg13g2_decap_8 FILLER_60_1500 ();
 sg13g2_decap_8 FILLER_60_1507 ();
 sg13g2_decap_8 FILLER_60_1514 ();
 sg13g2_decap_8 FILLER_60_1521 ();
 sg13g2_decap_8 FILLER_60_1528 ();
 sg13g2_decap_8 FILLER_60_1535 ();
 sg13g2_decap_8 FILLER_60_1542 ();
 sg13g2_decap_8 FILLER_60_1549 ();
 sg13g2_decap_8 FILLER_60_1556 ();
 sg13g2_decap_8 FILLER_60_1563 ();
 sg13g2_decap_8 FILLER_60_1570 ();
 sg13g2_decap_8 FILLER_60_1577 ();
 sg13g2_decap_8 FILLER_60_1584 ();
 sg13g2_decap_8 FILLER_60_1591 ();
 sg13g2_decap_8 FILLER_60_1598 ();
 sg13g2_decap_8 FILLER_60_1605 ();
 sg13g2_decap_8 FILLER_60_1612 ();
 sg13g2_decap_8 FILLER_60_1619 ();
 sg13g2_decap_8 FILLER_60_1626 ();
 sg13g2_decap_8 FILLER_60_1633 ();
 sg13g2_decap_8 FILLER_60_1640 ();
 sg13g2_decap_8 FILLER_60_1647 ();
 sg13g2_decap_8 FILLER_60_1654 ();
 sg13g2_decap_8 FILLER_60_1661 ();
 sg13g2_decap_8 FILLER_60_1668 ();
 sg13g2_decap_8 FILLER_60_1675 ();
 sg13g2_decap_8 FILLER_60_1682 ();
 sg13g2_decap_8 FILLER_60_1689 ();
 sg13g2_decap_8 FILLER_60_1696 ();
 sg13g2_decap_8 FILLER_60_1703 ();
 sg13g2_decap_8 FILLER_60_1710 ();
 sg13g2_decap_8 FILLER_60_1717 ();
 sg13g2_decap_8 FILLER_60_1724 ();
 sg13g2_decap_8 FILLER_60_1731 ();
 sg13g2_decap_8 FILLER_60_1738 ();
 sg13g2_decap_8 FILLER_60_1745 ();
 sg13g2_decap_8 FILLER_60_1752 ();
 sg13g2_decap_8 FILLER_60_1759 ();
 sg13g2_fill_2 FILLER_60_1766 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_4 FILLER_61_28 ();
 sg13g2_fill_1 FILLER_61_69 ();
 sg13g2_fill_2 FILLER_61_146 ();
 sg13g2_decap_4 FILLER_61_153 ();
 sg13g2_fill_2 FILLER_61_157 ();
 sg13g2_fill_2 FILLER_61_164 ();
 sg13g2_fill_1 FILLER_61_166 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_fill_2 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_182 ();
 sg13g2_fill_2 FILLER_61_201 ();
 sg13g2_fill_1 FILLER_61_203 ();
 sg13g2_fill_2 FILLER_61_214 ();
 sg13g2_fill_1 FILLER_61_252 ();
 sg13g2_fill_2 FILLER_61_262 ();
 sg13g2_fill_2 FILLER_61_269 ();
 sg13g2_fill_1 FILLER_61_271 ();
 sg13g2_fill_1 FILLER_61_306 ();
 sg13g2_fill_2 FILLER_61_320 ();
 sg13g2_fill_1 FILLER_61_322 ();
 sg13g2_fill_2 FILLER_61_368 ();
 sg13g2_fill_2 FILLER_61_397 ();
 sg13g2_decap_8 FILLER_61_454 ();
 sg13g2_fill_2 FILLER_61_461 ();
 sg13g2_decap_8 FILLER_61_467 ();
 sg13g2_decap_4 FILLER_61_474 ();
 sg13g2_fill_1 FILLER_61_478 ();
 sg13g2_decap_8 FILLER_61_516 ();
 sg13g2_fill_1 FILLER_61_528 ();
 sg13g2_decap_4 FILLER_61_537 ();
 sg13g2_fill_1 FILLER_61_551 ();
 sg13g2_fill_2 FILLER_61_557 ();
 sg13g2_fill_1 FILLER_61_574 ();
 sg13g2_decap_4 FILLER_61_664 ();
 sg13g2_fill_2 FILLER_61_676 ();
 sg13g2_fill_1 FILLER_61_678 ();
 sg13g2_fill_1 FILLER_61_706 ();
 sg13g2_fill_2 FILLER_61_727 ();
 sg13g2_decap_4 FILLER_61_735 ();
 sg13g2_fill_1 FILLER_61_765 ();
 sg13g2_fill_1 FILLER_61_780 ();
 sg13g2_fill_1 FILLER_61_808 ();
 sg13g2_decap_4 FILLER_61_814 ();
 sg13g2_decap_4 FILLER_61_855 ();
 sg13g2_fill_2 FILLER_61_906 ();
 sg13g2_fill_2 FILLER_61_912 ();
 sg13g2_fill_2 FILLER_61_928 ();
 sg13g2_fill_2 FILLER_61_939 ();
 sg13g2_fill_2 FILLER_61_1032 ();
 sg13g2_fill_2 FILLER_61_1071 ();
 sg13g2_fill_1 FILLER_61_1147 ();
 sg13g2_decap_8 FILLER_61_1161 ();
 sg13g2_decap_8 FILLER_61_1168 ();
 sg13g2_decap_8 FILLER_61_1175 ();
 sg13g2_decap_8 FILLER_61_1182 ();
 sg13g2_decap_8 FILLER_61_1189 ();
 sg13g2_decap_8 FILLER_61_1196 ();
 sg13g2_decap_8 FILLER_61_1203 ();
 sg13g2_decap_8 FILLER_61_1210 ();
 sg13g2_decap_8 FILLER_61_1217 ();
 sg13g2_decap_8 FILLER_61_1224 ();
 sg13g2_decap_8 FILLER_61_1231 ();
 sg13g2_decap_8 FILLER_61_1238 ();
 sg13g2_decap_8 FILLER_61_1245 ();
 sg13g2_decap_8 FILLER_61_1252 ();
 sg13g2_decap_8 FILLER_61_1259 ();
 sg13g2_decap_8 FILLER_61_1266 ();
 sg13g2_decap_8 FILLER_61_1273 ();
 sg13g2_decap_8 FILLER_61_1280 ();
 sg13g2_decap_8 FILLER_61_1287 ();
 sg13g2_decap_8 FILLER_61_1294 ();
 sg13g2_decap_8 FILLER_61_1301 ();
 sg13g2_decap_8 FILLER_61_1308 ();
 sg13g2_decap_8 FILLER_61_1315 ();
 sg13g2_decap_8 FILLER_61_1322 ();
 sg13g2_decap_8 FILLER_61_1329 ();
 sg13g2_decap_8 FILLER_61_1336 ();
 sg13g2_decap_8 FILLER_61_1343 ();
 sg13g2_decap_8 FILLER_61_1350 ();
 sg13g2_decap_8 FILLER_61_1357 ();
 sg13g2_decap_8 FILLER_61_1364 ();
 sg13g2_decap_8 FILLER_61_1371 ();
 sg13g2_decap_8 FILLER_61_1378 ();
 sg13g2_decap_8 FILLER_61_1385 ();
 sg13g2_decap_8 FILLER_61_1392 ();
 sg13g2_decap_8 FILLER_61_1399 ();
 sg13g2_decap_8 FILLER_61_1406 ();
 sg13g2_decap_8 FILLER_61_1413 ();
 sg13g2_decap_8 FILLER_61_1420 ();
 sg13g2_decap_8 FILLER_61_1427 ();
 sg13g2_decap_8 FILLER_61_1434 ();
 sg13g2_decap_8 FILLER_61_1441 ();
 sg13g2_decap_8 FILLER_61_1448 ();
 sg13g2_decap_8 FILLER_61_1455 ();
 sg13g2_decap_8 FILLER_61_1462 ();
 sg13g2_decap_8 FILLER_61_1469 ();
 sg13g2_decap_8 FILLER_61_1476 ();
 sg13g2_decap_8 FILLER_61_1483 ();
 sg13g2_decap_8 FILLER_61_1490 ();
 sg13g2_decap_8 FILLER_61_1497 ();
 sg13g2_decap_8 FILLER_61_1504 ();
 sg13g2_decap_8 FILLER_61_1511 ();
 sg13g2_decap_8 FILLER_61_1518 ();
 sg13g2_decap_8 FILLER_61_1525 ();
 sg13g2_decap_8 FILLER_61_1532 ();
 sg13g2_decap_8 FILLER_61_1539 ();
 sg13g2_decap_8 FILLER_61_1546 ();
 sg13g2_decap_8 FILLER_61_1553 ();
 sg13g2_decap_8 FILLER_61_1560 ();
 sg13g2_decap_8 FILLER_61_1567 ();
 sg13g2_decap_8 FILLER_61_1574 ();
 sg13g2_decap_8 FILLER_61_1581 ();
 sg13g2_decap_8 FILLER_61_1588 ();
 sg13g2_decap_8 FILLER_61_1595 ();
 sg13g2_decap_8 FILLER_61_1602 ();
 sg13g2_decap_8 FILLER_61_1609 ();
 sg13g2_decap_8 FILLER_61_1616 ();
 sg13g2_decap_8 FILLER_61_1623 ();
 sg13g2_decap_8 FILLER_61_1630 ();
 sg13g2_decap_8 FILLER_61_1637 ();
 sg13g2_decap_8 FILLER_61_1644 ();
 sg13g2_decap_8 FILLER_61_1651 ();
 sg13g2_decap_8 FILLER_61_1658 ();
 sg13g2_decap_8 FILLER_61_1665 ();
 sg13g2_decap_8 FILLER_61_1672 ();
 sg13g2_decap_8 FILLER_61_1679 ();
 sg13g2_decap_8 FILLER_61_1686 ();
 sg13g2_decap_8 FILLER_61_1693 ();
 sg13g2_decap_8 FILLER_61_1700 ();
 sg13g2_decap_8 FILLER_61_1707 ();
 sg13g2_decap_8 FILLER_61_1714 ();
 sg13g2_decap_8 FILLER_61_1721 ();
 sg13g2_decap_8 FILLER_61_1728 ();
 sg13g2_decap_8 FILLER_61_1735 ();
 sg13g2_decap_8 FILLER_61_1742 ();
 sg13g2_decap_8 FILLER_61_1749 ();
 sg13g2_decap_8 FILLER_61_1756 ();
 sg13g2_decap_4 FILLER_61_1763 ();
 sg13g2_fill_1 FILLER_61_1767 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_14 ();
 sg13g2_fill_1 FILLER_62_42 ();
 sg13g2_fill_2 FILLER_62_100 ();
 sg13g2_fill_1 FILLER_62_172 ();
 sg13g2_fill_2 FILLER_62_196 ();
 sg13g2_fill_1 FILLER_62_198 ();
 sg13g2_fill_2 FILLER_62_229 ();
 sg13g2_fill_2 FILLER_62_250 ();
 sg13g2_fill_1 FILLER_62_261 ();
 sg13g2_fill_2 FILLER_62_275 ();
 sg13g2_fill_1 FILLER_62_277 ();
 sg13g2_fill_1 FILLER_62_283 ();
 sg13g2_fill_2 FILLER_62_313 ();
 sg13g2_fill_1 FILLER_62_315 ();
 sg13g2_decap_4 FILLER_62_322 ();
 sg13g2_fill_1 FILLER_62_326 ();
 sg13g2_fill_2 FILLER_62_355 ();
 sg13g2_decap_4 FILLER_62_381 ();
 sg13g2_fill_1 FILLER_62_404 ();
 sg13g2_fill_1 FILLER_62_440 ();
 sg13g2_decap_8 FILLER_62_455 ();
 sg13g2_fill_1 FILLER_62_462 ();
 sg13g2_decap_4 FILLER_62_477 ();
 sg13g2_fill_1 FILLER_62_489 ();
 sg13g2_fill_1 FILLER_62_495 ();
 sg13g2_fill_2 FILLER_62_501 ();
 sg13g2_fill_1 FILLER_62_503 ();
 sg13g2_fill_2 FILLER_62_517 ();
 sg13g2_fill_1 FILLER_62_519 ();
 sg13g2_fill_1 FILLER_62_532 ();
 sg13g2_decap_4 FILLER_62_538 ();
 sg13g2_fill_2 FILLER_62_542 ();
 sg13g2_fill_2 FILLER_62_554 ();
 sg13g2_fill_1 FILLER_62_562 ();
 sg13g2_fill_1 FILLER_62_573 ();
 sg13g2_fill_2 FILLER_62_577 ();
 sg13g2_fill_1 FILLER_62_579 ();
 sg13g2_fill_2 FILLER_62_607 ();
 sg13g2_decap_8 FILLER_62_621 ();
 sg13g2_fill_1 FILLER_62_628 ();
 sg13g2_fill_2 FILLER_62_636 ();
 sg13g2_fill_1 FILLER_62_638 ();
 sg13g2_decap_8 FILLER_62_652 ();
 sg13g2_decap_8 FILLER_62_659 ();
 sg13g2_decap_8 FILLER_62_666 ();
 sg13g2_fill_2 FILLER_62_673 ();
 sg13g2_decap_8 FILLER_62_693 ();
 sg13g2_decap_8 FILLER_62_700 ();
 sg13g2_fill_2 FILLER_62_707 ();
 sg13g2_fill_2 FILLER_62_722 ();
 sg13g2_decap_4 FILLER_62_734 ();
 sg13g2_fill_2 FILLER_62_738 ();
 sg13g2_fill_2 FILLER_62_747 ();
 sg13g2_decap_4 FILLER_62_817 ();
 sg13g2_fill_1 FILLER_62_839 ();
 sg13g2_decap_4 FILLER_62_858 ();
 sg13g2_fill_2 FILLER_62_862 ();
 sg13g2_fill_2 FILLER_62_989 ();
 sg13g2_fill_1 FILLER_62_991 ();
 sg13g2_decap_8 FILLER_62_1167 ();
 sg13g2_decap_8 FILLER_62_1174 ();
 sg13g2_decap_8 FILLER_62_1181 ();
 sg13g2_decap_8 FILLER_62_1188 ();
 sg13g2_decap_8 FILLER_62_1195 ();
 sg13g2_decap_8 FILLER_62_1202 ();
 sg13g2_decap_8 FILLER_62_1209 ();
 sg13g2_decap_8 FILLER_62_1216 ();
 sg13g2_decap_8 FILLER_62_1223 ();
 sg13g2_decap_8 FILLER_62_1230 ();
 sg13g2_decap_8 FILLER_62_1237 ();
 sg13g2_decap_8 FILLER_62_1244 ();
 sg13g2_decap_8 FILLER_62_1251 ();
 sg13g2_decap_8 FILLER_62_1258 ();
 sg13g2_decap_8 FILLER_62_1265 ();
 sg13g2_decap_8 FILLER_62_1272 ();
 sg13g2_decap_8 FILLER_62_1279 ();
 sg13g2_decap_8 FILLER_62_1286 ();
 sg13g2_decap_8 FILLER_62_1293 ();
 sg13g2_decap_8 FILLER_62_1300 ();
 sg13g2_decap_8 FILLER_62_1307 ();
 sg13g2_decap_8 FILLER_62_1314 ();
 sg13g2_decap_8 FILLER_62_1321 ();
 sg13g2_decap_8 FILLER_62_1328 ();
 sg13g2_decap_8 FILLER_62_1335 ();
 sg13g2_decap_8 FILLER_62_1342 ();
 sg13g2_decap_8 FILLER_62_1349 ();
 sg13g2_decap_8 FILLER_62_1356 ();
 sg13g2_decap_8 FILLER_62_1363 ();
 sg13g2_decap_8 FILLER_62_1370 ();
 sg13g2_decap_8 FILLER_62_1377 ();
 sg13g2_decap_8 FILLER_62_1384 ();
 sg13g2_decap_8 FILLER_62_1391 ();
 sg13g2_decap_8 FILLER_62_1398 ();
 sg13g2_decap_8 FILLER_62_1405 ();
 sg13g2_decap_8 FILLER_62_1412 ();
 sg13g2_decap_8 FILLER_62_1419 ();
 sg13g2_decap_8 FILLER_62_1426 ();
 sg13g2_decap_8 FILLER_62_1433 ();
 sg13g2_decap_8 FILLER_62_1440 ();
 sg13g2_decap_8 FILLER_62_1447 ();
 sg13g2_decap_8 FILLER_62_1454 ();
 sg13g2_decap_8 FILLER_62_1461 ();
 sg13g2_decap_8 FILLER_62_1468 ();
 sg13g2_decap_8 FILLER_62_1475 ();
 sg13g2_decap_8 FILLER_62_1482 ();
 sg13g2_decap_8 FILLER_62_1489 ();
 sg13g2_decap_8 FILLER_62_1496 ();
 sg13g2_decap_8 FILLER_62_1503 ();
 sg13g2_decap_8 FILLER_62_1510 ();
 sg13g2_decap_8 FILLER_62_1517 ();
 sg13g2_decap_8 FILLER_62_1524 ();
 sg13g2_decap_8 FILLER_62_1531 ();
 sg13g2_decap_8 FILLER_62_1538 ();
 sg13g2_decap_8 FILLER_62_1545 ();
 sg13g2_decap_8 FILLER_62_1552 ();
 sg13g2_decap_8 FILLER_62_1559 ();
 sg13g2_decap_8 FILLER_62_1566 ();
 sg13g2_decap_8 FILLER_62_1573 ();
 sg13g2_decap_8 FILLER_62_1580 ();
 sg13g2_decap_8 FILLER_62_1587 ();
 sg13g2_decap_8 FILLER_62_1594 ();
 sg13g2_decap_8 FILLER_62_1601 ();
 sg13g2_decap_8 FILLER_62_1608 ();
 sg13g2_decap_8 FILLER_62_1615 ();
 sg13g2_decap_8 FILLER_62_1622 ();
 sg13g2_decap_8 FILLER_62_1629 ();
 sg13g2_decap_8 FILLER_62_1636 ();
 sg13g2_decap_8 FILLER_62_1643 ();
 sg13g2_decap_8 FILLER_62_1650 ();
 sg13g2_decap_8 FILLER_62_1657 ();
 sg13g2_decap_8 FILLER_62_1664 ();
 sg13g2_decap_8 FILLER_62_1671 ();
 sg13g2_decap_8 FILLER_62_1678 ();
 sg13g2_decap_8 FILLER_62_1685 ();
 sg13g2_decap_8 FILLER_62_1692 ();
 sg13g2_decap_8 FILLER_62_1699 ();
 sg13g2_decap_8 FILLER_62_1706 ();
 sg13g2_decap_8 FILLER_62_1713 ();
 sg13g2_decap_8 FILLER_62_1720 ();
 sg13g2_decap_8 FILLER_62_1727 ();
 sg13g2_decap_8 FILLER_62_1734 ();
 sg13g2_decap_8 FILLER_62_1741 ();
 sg13g2_decap_8 FILLER_62_1748 ();
 sg13g2_decap_8 FILLER_62_1755 ();
 sg13g2_decap_4 FILLER_62_1762 ();
 sg13g2_fill_2 FILLER_62_1766 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_4 FILLER_63_14 ();
 sg13g2_fill_1 FILLER_63_18 ();
 sg13g2_fill_1 FILLER_63_77 ();
 sg13g2_fill_1 FILLER_63_201 ();
 sg13g2_fill_1 FILLER_63_212 ();
 sg13g2_fill_2 FILLER_63_231 ();
 sg13g2_fill_1 FILLER_63_233 ();
 sg13g2_fill_2 FILLER_63_243 ();
 sg13g2_fill_1 FILLER_63_245 ();
 sg13g2_fill_1 FILLER_63_254 ();
 sg13g2_fill_1 FILLER_63_270 ();
 sg13g2_decap_8 FILLER_63_281 ();
 sg13g2_decap_8 FILLER_63_288 ();
 sg13g2_fill_2 FILLER_63_295 ();
 sg13g2_fill_1 FILLER_63_297 ();
 sg13g2_fill_2 FILLER_63_317 ();
 sg13g2_fill_1 FILLER_63_319 ();
 sg13g2_fill_1 FILLER_63_330 ();
 sg13g2_fill_1 FILLER_63_345 ();
 sg13g2_fill_1 FILLER_63_367 ();
 sg13g2_decap_4 FILLER_63_376 ();
 sg13g2_decap_8 FILLER_63_386 ();
 sg13g2_fill_1 FILLER_63_393 ();
 sg13g2_fill_2 FILLER_63_439 ();
 sg13g2_fill_1 FILLER_63_441 ();
 sg13g2_fill_1 FILLER_63_477 ();
 sg13g2_decap_4 FILLER_63_515 ();
 sg13g2_fill_2 FILLER_63_532 ();
 sg13g2_fill_2 FILLER_63_551 ();
 sg13g2_fill_1 FILLER_63_568 ();
 sg13g2_fill_2 FILLER_63_575 ();
 sg13g2_fill_1 FILLER_63_577 ();
 sg13g2_fill_2 FILLER_63_586 ();
 sg13g2_fill_1 FILLER_63_606 ();
 sg13g2_fill_1 FILLER_63_617 ();
 sg13g2_decap_4 FILLER_63_624 ();
 sg13g2_fill_1 FILLER_63_655 ();
 sg13g2_decap_4 FILLER_63_667 ();
 sg13g2_fill_2 FILLER_63_681 ();
 sg13g2_fill_1 FILLER_63_688 ();
 sg13g2_fill_2 FILLER_63_698 ();
 sg13g2_fill_1 FILLER_63_700 ();
 sg13g2_fill_2 FILLER_63_722 ();
 sg13g2_fill_1 FILLER_63_724 ();
 sg13g2_decap_8 FILLER_63_730 ();
 sg13g2_fill_2 FILLER_63_737 ();
 sg13g2_fill_1 FILLER_63_739 ();
 sg13g2_fill_2 FILLER_63_763 ();
 sg13g2_fill_1 FILLER_63_765 ();
 sg13g2_fill_2 FILLER_63_780 ();
 sg13g2_fill_2 FILLER_63_802 ();
 sg13g2_fill_1 FILLER_63_804 ();
 sg13g2_fill_2 FILLER_63_809 ();
 sg13g2_fill_1 FILLER_63_811 ();
 sg13g2_fill_1 FILLER_63_829 ();
 sg13g2_fill_1 FILLER_63_839 ();
 sg13g2_fill_1 FILLER_63_914 ();
 sg13g2_fill_2 FILLER_63_933 ();
 sg13g2_fill_1 FILLER_63_935 ();
 sg13g2_fill_1 FILLER_63_950 ();
 sg13g2_fill_2 FILLER_63_977 ();
 sg13g2_fill_2 FILLER_63_992 ();
 sg13g2_fill_1 FILLER_63_994 ();
 sg13g2_fill_2 FILLER_63_1121 ();
 sg13g2_decap_8 FILLER_63_1177 ();
 sg13g2_decap_8 FILLER_63_1184 ();
 sg13g2_decap_8 FILLER_63_1191 ();
 sg13g2_decap_8 FILLER_63_1198 ();
 sg13g2_decap_8 FILLER_63_1205 ();
 sg13g2_decap_8 FILLER_63_1212 ();
 sg13g2_decap_8 FILLER_63_1219 ();
 sg13g2_decap_8 FILLER_63_1226 ();
 sg13g2_decap_8 FILLER_63_1233 ();
 sg13g2_decap_8 FILLER_63_1240 ();
 sg13g2_decap_8 FILLER_63_1247 ();
 sg13g2_decap_8 FILLER_63_1254 ();
 sg13g2_decap_8 FILLER_63_1261 ();
 sg13g2_decap_8 FILLER_63_1268 ();
 sg13g2_decap_8 FILLER_63_1275 ();
 sg13g2_decap_8 FILLER_63_1282 ();
 sg13g2_decap_8 FILLER_63_1289 ();
 sg13g2_decap_8 FILLER_63_1296 ();
 sg13g2_decap_8 FILLER_63_1303 ();
 sg13g2_decap_8 FILLER_63_1310 ();
 sg13g2_decap_8 FILLER_63_1317 ();
 sg13g2_decap_8 FILLER_63_1324 ();
 sg13g2_decap_8 FILLER_63_1331 ();
 sg13g2_decap_8 FILLER_63_1338 ();
 sg13g2_decap_8 FILLER_63_1345 ();
 sg13g2_decap_8 FILLER_63_1352 ();
 sg13g2_decap_8 FILLER_63_1359 ();
 sg13g2_decap_8 FILLER_63_1366 ();
 sg13g2_decap_8 FILLER_63_1373 ();
 sg13g2_decap_8 FILLER_63_1380 ();
 sg13g2_decap_8 FILLER_63_1387 ();
 sg13g2_decap_8 FILLER_63_1394 ();
 sg13g2_decap_8 FILLER_63_1401 ();
 sg13g2_decap_8 FILLER_63_1408 ();
 sg13g2_decap_8 FILLER_63_1415 ();
 sg13g2_decap_8 FILLER_63_1422 ();
 sg13g2_decap_8 FILLER_63_1429 ();
 sg13g2_decap_8 FILLER_63_1436 ();
 sg13g2_decap_8 FILLER_63_1443 ();
 sg13g2_decap_8 FILLER_63_1450 ();
 sg13g2_decap_8 FILLER_63_1457 ();
 sg13g2_decap_8 FILLER_63_1464 ();
 sg13g2_decap_8 FILLER_63_1471 ();
 sg13g2_decap_8 FILLER_63_1478 ();
 sg13g2_decap_8 FILLER_63_1485 ();
 sg13g2_decap_8 FILLER_63_1492 ();
 sg13g2_decap_8 FILLER_63_1499 ();
 sg13g2_decap_8 FILLER_63_1506 ();
 sg13g2_decap_8 FILLER_63_1513 ();
 sg13g2_decap_8 FILLER_63_1520 ();
 sg13g2_decap_8 FILLER_63_1527 ();
 sg13g2_decap_8 FILLER_63_1534 ();
 sg13g2_decap_8 FILLER_63_1541 ();
 sg13g2_decap_8 FILLER_63_1548 ();
 sg13g2_decap_8 FILLER_63_1555 ();
 sg13g2_decap_8 FILLER_63_1562 ();
 sg13g2_decap_8 FILLER_63_1569 ();
 sg13g2_decap_8 FILLER_63_1576 ();
 sg13g2_decap_8 FILLER_63_1583 ();
 sg13g2_decap_8 FILLER_63_1590 ();
 sg13g2_decap_8 FILLER_63_1597 ();
 sg13g2_decap_8 FILLER_63_1604 ();
 sg13g2_decap_8 FILLER_63_1611 ();
 sg13g2_decap_8 FILLER_63_1618 ();
 sg13g2_decap_8 FILLER_63_1625 ();
 sg13g2_decap_8 FILLER_63_1632 ();
 sg13g2_decap_8 FILLER_63_1639 ();
 sg13g2_decap_8 FILLER_63_1646 ();
 sg13g2_decap_8 FILLER_63_1653 ();
 sg13g2_decap_8 FILLER_63_1660 ();
 sg13g2_decap_8 FILLER_63_1667 ();
 sg13g2_decap_8 FILLER_63_1674 ();
 sg13g2_decap_8 FILLER_63_1681 ();
 sg13g2_decap_8 FILLER_63_1688 ();
 sg13g2_decap_8 FILLER_63_1695 ();
 sg13g2_decap_8 FILLER_63_1702 ();
 sg13g2_decap_8 FILLER_63_1709 ();
 sg13g2_decap_8 FILLER_63_1716 ();
 sg13g2_decap_8 FILLER_63_1723 ();
 sg13g2_decap_8 FILLER_63_1730 ();
 sg13g2_decap_8 FILLER_63_1737 ();
 sg13g2_decap_8 FILLER_63_1744 ();
 sg13g2_decap_8 FILLER_63_1751 ();
 sg13g2_decap_8 FILLER_63_1758 ();
 sg13g2_fill_2 FILLER_63_1765 ();
 sg13g2_fill_1 FILLER_63_1767 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_14 ();
 sg13g2_fill_1 FILLER_64_94 ();
 sg13g2_fill_1 FILLER_64_148 ();
 sg13g2_fill_1 FILLER_64_157 ();
 sg13g2_fill_2 FILLER_64_239 ();
 sg13g2_decap_4 FILLER_64_246 ();
 sg13g2_fill_2 FILLER_64_250 ();
 sg13g2_fill_1 FILLER_64_278 ();
 sg13g2_decap_4 FILLER_64_291 ();
 sg13g2_fill_1 FILLER_64_300 ();
 sg13g2_fill_2 FILLER_64_321 ();
 sg13g2_fill_1 FILLER_64_323 ();
 sg13g2_fill_2 FILLER_64_340 ();
 sg13g2_decap_8 FILLER_64_376 ();
 sg13g2_fill_1 FILLER_64_383 ();
 sg13g2_fill_2 FILLER_64_387 ();
 sg13g2_fill_1 FILLER_64_389 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_fill_1 FILLER_64_409 ();
 sg13g2_fill_1 FILLER_64_430 ();
 sg13g2_decap_8 FILLER_64_445 ();
 sg13g2_decap_8 FILLER_64_452 ();
 sg13g2_decap_8 FILLER_64_459 ();
 sg13g2_fill_2 FILLER_64_466 ();
 sg13g2_fill_1 FILLER_64_468 ();
 sg13g2_fill_2 FILLER_64_474 ();
 sg13g2_fill_1 FILLER_64_482 ();
 sg13g2_decap_4 FILLER_64_488 ();
 sg13g2_fill_1 FILLER_64_510 ();
 sg13g2_fill_1 FILLER_64_534 ();
 sg13g2_decap_8 FILLER_64_549 ();
 sg13g2_decap_4 FILLER_64_556 ();
 sg13g2_decap_4 FILLER_64_570 ();
 sg13g2_fill_2 FILLER_64_574 ();
 sg13g2_decap_8 FILLER_64_594 ();
 sg13g2_fill_1 FILLER_64_618 ();
 sg13g2_fill_1 FILLER_64_626 ();
 sg13g2_fill_1 FILLER_64_653 ();
 sg13g2_decap_4 FILLER_64_659 ();
 sg13g2_fill_1 FILLER_64_663 ();
 sg13g2_fill_1 FILLER_64_690 ();
 sg13g2_decap_8 FILLER_64_699 ();
 sg13g2_fill_2 FILLER_64_706 ();
 sg13g2_fill_1 FILLER_64_708 ();
 sg13g2_decap_4 FILLER_64_714 ();
 sg13g2_fill_2 FILLER_64_724 ();
 sg13g2_fill_1 FILLER_64_735 ();
 sg13g2_decap_4 FILLER_64_766 ();
 sg13g2_fill_2 FILLER_64_775 ();
 sg13g2_fill_2 FILLER_64_797 ();
 sg13g2_fill_1 FILLER_64_799 ();
 sg13g2_fill_2 FILLER_64_815 ();
 sg13g2_fill_1 FILLER_64_817 ();
 sg13g2_fill_2 FILLER_64_830 ();
 sg13g2_fill_1 FILLER_64_843 ();
 sg13g2_decap_4 FILLER_64_859 ();
 sg13g2_fill_2 FILLER_64_971 ();
 sg13g2_fill_1 FILLER_64_973 ();
 sg13g2_fill_1 FILLER_64_1009 ();
 sg13g2_fill_1 FILLER_64_1048 ();
 sg13g2_fill_2 FILLER_64_1095 ();
 sg13g2_decap_8 FILLER_64_1185 ();
 sg13g2_decap_8 FILLER_64_1192 ();
 sg13g2_decap_8 FILLER_64_1199 ();
 sg13g2_decap_8 FILLER_64_1206 ();
 sg13g2_decap_8 FILLER_64_1213 ();
 sg13g2_decap_8 FILLER_64_1220 ();
 sg13g2_decap_8 FILLER_64_1227 ();
 sg13g2_decap_8 FILLER_64_1234 ();
 sg13g2_decap_8 FILLER_64_1241 ();
 sg13g2_decap_8 FILLER_64_1248 ();
 sg13g2_decap_8 FILLER_64_1255 ();
 sg13g2_decap_8 FILLER_64_1262 ();
 sg13g2_decap_8 FILLER_64_1269 ();
 sg13g2_decap_8 FILLER_64_1276 ();
 sg13g2_decap_8 FILLER_64_1283 ();
 sg13g2_decap_8 FILLER_64_1290 ();
 sg13g2_decap_8 FILLER_64_1297 ();
 sg13g2_decap_8 FILLER_64_1304 ();
 sg13g2_decap_8 FILLER_64_1311 ();
 sg13g2_decap_8 FILLER_64_1318 ();
 sg13g2_decap_8 FILLER_64_1325 ();
 sg13g2_decap_8 FILLER_64_1332 ();
 sg13g2_decap_8 FILLER_64_1339 ();
 sg13g2_decap_8 FILLER_64_1346 ();
 sg13g2_decap_8 FILLER_64_1353 ();
 sg13g2_decap_8 FILLER_64_1360 ();
 sg13g2_decap_8 FILLER_64_1367 ();
 sg13g2_decap_8 FILLER_64_1374 ();
 sg13g2_decap_8 FILLER_64_1381 ();
 sg13g2_decap_8 FILLER_64_1388 ();
 sg13g2_decap_8 FILLER_64_1395 ();
 sg13g2_decap_8 FILLER_64_1402 ();
 sg13g2_decap_8 FILLER_64_1409 ();
 sg13g2_decap_8 FILLER_64_1416 ();
 sg13g2_decap_8 FILLER_64_1423 ();
 sg13g2_decap_8 FILLER_64_1430 ();
 sg13g2_decap_8 FILLER_64_1437 ();
 sg13g2_decap_8 FILLER_64_1444 ();
 sg13g2_decap_8 FILLER_64_1451 ();
 sg13g2_decap_8 FILLER_64_1458 ();
 sg13g2_decap_8 FILLER_64_1465 ();
 sg13g2_decap_8 FILLER_64_1472 ();
 sg13g2_decap_8 FILLER_64_1479 ();
 sg13g2_decap_8 FILLER_64_1486 ();
 sg13g2_decap_8 FILLER_64_1493 ();
 sg13g2_decap_8 FILLER_64_1500 ();
 sg13g2_decap_8 FILLER_64_1507 ();
 sg13g2_decap_8 FILLER_64_1514 ();
 sg13g2_decap_8 FILLER_64_1521 ();
 sg13g2_decap_8 FILLER_64_1528 ();
 sg13g2_decap_8 FILLER_64_1535 ();
 sg13g2_decap_8 FILLER_64_1542 ();
 sg13g2_decap_8 FILLER_64_1549 ();
 sg13g2_decap_8 FILLER_64_1556 ();
 sg13g2_decap_8 FILLER_64_1563 ();
 sg13g2_decap_8 FILLER_64_1570 ();
 sg13g2_decap_8 FILLER_64_1577 ();
 sg13g2_decap_8 FILLER_64_1584 ();
 sg13g2_decap_8 FILLER_64_1591 ();
 sg13g2_decap_8 FILLER_64_1598 ();
 sg13g2_decap_8 FILLER_64_1605 ();
 sg13g2_decap_8 FILLER_64_1612 ();
 sg13g2_decap_8 FILLER_64_1619 ();
 sg13g2_decap_8 FILLER_64_1626 ();
 sg13g2_decap_8 FILLER_64_1633 ();
 sg13g2_decap_8 FILLER_64_1640 ();
 sg13g2_decap_8 FILLER_64_1647 ();
 sg13g2_decap_8 FILLER_64_1654 ();
 sg13g2_decap_8 FILLER_64_1661 ();
 sg13g2_decap_8 FILLER_64_1668 ();
 sg13g2_decap_8 FILLER_64_1675 ();
 sg13g2_decap_8 FILLER_64_1682 ();
 sg13g2_decap_8 FILLER_64_1689 ();
 sg13g2_decap_8 FILLER_64_1696 ();
 sg13g2_decap_8 FILLER_64_1703 ();
 sg13g2_decap_8 FILLER_64_1710 ();
 sg13g2_decap_8 FILLER_64_1717 ();
 sg13g2_decap_8 FILLER_64_1724 ();
 sg13g2_decap_8 FILLER_64_1731 ();
 sg13g2_decap_8 FILLER_64_1738 ();
 sg13g2_decap_8 FILLER_64_1745 ();
 sg13g2_decap_8 FILLER_64_1752 ();
 sg13g2_decap_8 FILLER_64_1759 ();
 sg13g2_fill_2 FILLER_64_1766 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_fill_2 FILLER_65_28 ();
 sg13g2_fill_1 FILLER_65_30 ();
 sg13g2_fill_2 FILLER_65_69 ();
 sg13g2_fill_1 FILLER_65_71 ();
 sg13g2_fill_1 FILLER_65_134 ();
 sg13g2_fill_2 FILLER_65_140 ();
 sg13g2_fill_2 FILLER_65_151 ();
 sg13g2_fill_1 FILLER_65_179 ();
 sg13g2_fill_1 FILLER_65_221 ();
 sg13g2_fill_2 FILLER_65_229 ();
 sg13g2_fill_1 FILLER_65_231 ();
 sg13g2_fill_1 FILLER_65_252 ();
 sg13g2_fill_2 FILLER_65_287 ();
 sg13g2_fill_1 FILLER_65_289 ();
 sg13g2_fill_2 FILLER_65_311 ();
 sg13g2_fill_2 FILLER_65_322 ();
 sg13g2_decap_4 FILLER_65_353 ();
 sg13g2_fill_1 FILLER_65_377 ();
 sg13g2_decap_4 FILLER_65_450 ();
 sg13g2_decap_8 FILLER_65_476 ();
 sg13g2_decap_4 FILLER_65_483 ();
 sg13g2_fill_2 FILLER_65_492 ();
 sg13g2_fill_1 FILLER_65_494 ();
 sg13g2_fill_1 FILLER_65_500 ();
 sg13g2_fill_2 FILLER_65_511 ();
 sg13g2_fill_1 FILLER_65_513 ();
 sg13g2_fill_1 FILLER_65_524 ();
 sg13g2_fill_2 FILLER_65_530 ();
 sg13g2_fill_1 FILLER_65_532 ();
 sg13g2_decap_4 FILLER_65_553 ();
 sg13g2_fill_2 FILLER_65_557 ();
 sg13g2_fill_1 FILLER_65_571 ();
 sg13g2_fill_2 FILLER_65_595 ();
 sg13g2_fill_1 FILLER_65_597 ();
 sg13g2_decap_4 FILLER_65_604 ();
 sg13g2_decap_4 FILLER_65_613 ();
 sg13g2_decap_8 FILLER_65_627 ();
 sg13g2_decap_8 FILLER_65_634 ();
 sg13g2_fill_2 FILLER_65_669 ();
 sg13g2_fill_2 FILLER_65_699 ();
 sg13g2_fill_2 FILLER_65_715 ();
 sg13g2_fill_1 FILLER_65_717 ();
 sg13g2_fill_1 FILLER_65_728 ();
 sg13g2_fill_2 FILLER_65_734 ();
 sg13g2_fill_1 FILLER_65_736 ();
 sg13g2_decap_4 FILLER_65_763 ();
 sg13g2_fill_2 FILLER_65_767 ();
 sg13g2_decap_4 FILLER_65_799 ();
 sg13g2_fill_2 FILLER_65_817 ();
 sg13g2_fill_1 FILLER_65_824 ();
 sg13g2_decap_8 FILLER_65_856 ();
 sg13g2_decap_8 FILLER_65_863 ();
 sg13g2_decap_8 FILLER_65_870 ();
 sg13g2_fill_2 FILLER_65_877 ();
 sg13g2_fill_1 FILLER_65_888 ();
 sg13g2_fill_1 FILLER_65_952 ();
 sg13g2_fill_2 FILLER_65_981 ();
 sg13g2_fill_2 FILLER_65_1052 ();
 sg13g2_fill_1 FILLER_65_1088 ();
 sg13g2_fill_1 FILLER_65_1148 ();
 sg13g2_decap_8 FILLER_65_1180 ();
 sg13g2_decap_8 FILLER_65_1187 ();
 sg13g2_decap_8 FILLER_65_1194 ();
 sg13g2_decap_8 FILLER_65_1201 ();
 sg13g2_decap_8 FILLER_65_1208 ();
 sg13g2_decap_8 FILLER_65_1215 ();
 sg13g2_decap_8 FILLER_65_1222 ();
 sg13g2_decap_8 FILLER_65_1229 ();
 sg13g2_decap_8 FILLER_65_1236 ();
 sg13g2_decap_8 FILLER_65_1243 ();
 sg13g2_decap_8 FILLER_65_1250 ();
 sg13g2_decap_8 FILLER_65_1257 ();
 sg13g2_decap_8 FILLER_65_1264 ();
 sg13g2_decap_8 FILLER_65_1271 ();
 sg13g2_decap_8 FILLER_65_1278 ();
 sg13g2_decap_8 FILLER_65_1285 ();
 sg13g2_decap_8 FILLER_65_1292 ();
 sg13g2_decap_8 FILLER_65_1299 ();
 sg13g2_decap_8 FILLER_65_1306 ();
 sg13g2_decap_8 FILLER_65_1313 ();
 sg13g2_decap_8 FILLER_65_1320 ();
 sg13g2_decap_8 FILLER_65_1327 ();
 sg13g2_decap_8 FILLER_65_1334 ();
 sg13g2_decap_8 FILLER_65_1341 ();
 sg13g2_decap_8 FILLER_65_1348 ();
 sg13g2_decap_8 FILLER_65_1355 ();
 sg13g2_decap_8 FILLER_65_1362 ();
 sg13g2_decap_8 FILLER_65_1369 ();
 sg13g2_decap_8 FILLER_65_1376 ();
 sg13g2_decap_8 FILLER_65_1383 ();
 sg13g2_decap_8 FILLER_65_1390 ();
 sg13g2_decap_8 FILLER_65_1397 ();
 sg13g2_decap_8 FILLER_65_1404 ();
 sg13g2_decap_8 FILLER_65_1411 ();
 sg13g2_decap_8 FILLER_65_1418 ();
 sg13g2_decap_8 FILLER_65_1425 ();
 sg13g2_decap_8 FILLER_65_1432 ();
 sg13g2_decap_8 FILLER_65_1439 ();
 sg13g2_decap_8 FILLER_65_1446 ();
 sg13g2_decap_8 FILLER_65_1453 ();
 sg13g2_decap_8 FILLER_65_1460 ();
 sg13g2_decap_8 FILLER_65_1467 ();
 sg13g2_decap_8 FILLER_65_1474 ();
 sg13g2_decap_8 FILLER_65_1481 ();
 sg13g2_decap_8 FILLER_65_1488 ();
 sg13g2_decap_8 FILLER_65_1495 ();
 sg13g2_decap_8 FILLER_65_1502 ();
 sg13g2_decap_8 FILLER_65_1509 ();
 sg13g2_decap_8 FILLER_65_1516 ();
 sg13g2_decap_8 FILLER_65_1523 ();
 sg13g2_decap_8 FILLER_65_1530 ();
 sg13g2_decap_8 FILLER_65_1537 ();
 sg13g2_decap_8 FILLER_65_1544 ();
 sg13g2_decap_8 FILLER_65_1551 ();
 sg13g2_decap_8 FILLER_65_1558 ();
 sg13g2_decap_8 FILLER_65_1565 ();
 sg13g2_decap_8 FILLER_65_1572 ();
 sg13g2_decap_8 FILLER_65_1579 ();
 sg13g2_decap_8 FILLER_65_1586 ();
 sg13g2_decap_8 FILLER_65_1593 ();
 sg13g2_decap_8 FILLER_65_1600 ();
 sg13g2_decap_8 FILLER_65_1607 ();
 sg13g2_decap_8 FILLER_65_1614 ();
 sg13g2_decap_8 FILLER_65_1621 ();
 sg13g2_decap_8 FILLER_65_1628 ();
 sg13g2_decap_8 FILLER_65_1635 ();
 sg13g2_decap_8 FILLER_65_1642 ();
 sg13g2_decap_8 FILLER_65_1649 ();
 sg13g2_decap_8 FILLER_65_1656 ();
 sg13g2_decap_8 FILLER_65_1663 ();
 sg13g2_decap_8 FILLER_65_1670 ();
 sg13g2_decap_8 FILLER_65_1677 ();
 sg13g2_decap_8 FILLER_65_1684 ();
 sg13g2_decap_8 FILLER_65_1691 ();
 sg13g2_decap_8 FILLER_65_1698 ();
 sg13g2_decap_8 FILLER_65_1705 ();
 sg13g2_decap_8 FILLER_65_1712 ();
 sg13g2_decap_8 FILLER_65_1719 ();
 sg13g2_decap_8 FILLER_65_1726 ();
 sg13g2_decap_8 FILLER_65_1733 ();
 sg13g2_decap_8 FILLER_65_1740 ();
 sg13g2_decap_8 FILLER_65_1747 ();
 sg13g2_decap_8 FILLER_65_1754 ();
 sg13g2_decap_8 FILLER_65_1761 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_fill_1 FILLER_66_35 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_fill_2 FILLER_66_156 ();
 sg13g2_fill_1 FILLER_66_203 ();
 sg13g2_fill_2 FILLER_66_218 ();
 sg13g2_fill_1 FILLER_66_220 ();
 sg13g2_fill_2 FILLER_66_291 ();
 sg13g2_decap_4 FILLER_66_297 ();
 sg13g2_fill_2 FILLER_66_305 ();
 sg13g2_fill_1 FILLER_66_328 ();
 sg13g2_fill_1 FILLER_66_365 ();
 sg13g2_fill_2 FILLER_66_393 ();
 sg13g2_fill_1 FILLER_66_455 ();
 sg13g2_fill_2 FILLER_66_473 ();
 sg13g2_fill_1 FILLER_66_475 ();
 sg13g2_fill_1 FILLER_66_488 ();
 sg13g2_fill_1 FILLER_66_494 ();
 sg13g2_fill_1 FILLER_66_519 ();
 sg13g2_fill_2 FILLER_66_549 ();
 sg13g2_fill_1 FILLER_66_551 ();
 sg13g2_fill_1 FILLER_66_558 ();
 sg13g2_fill_1 FILLER_66_595 ();
 sg13g2_fill_2 FILLER_66_636 ();
 sg13g2_fill_2 FILLER_66_671 ();
 sg13g2_fill_1 FILLER_66_673 ();
 sg13g2_fill_2 FILLER_66_684 ();
 sg13g2_fill_1 FILLER_66_686 ();
 sg13g2_fill_2 FILLER_66_692 ();
 sg13g2_fill_2 FILLER_66_723 ();
 sg13g2_fill_1 FILLER_66_725 ();
 sg13g2_fill_2 FILLER_66_750 ();
 sg13g2_fill_1 FILLER_66_752 ();
 sg13g2_fill_1 FILLER_66_767 ();
 sg13g2_fill_2 FILLER_66_794 ();
 sg13g2_fill_1 FILLER_66_835 ();
 sg13g2_fill_2 FILLER_66_867 ();
 sg13g2_fill_2 FILLER_66_877 ();
 sg13g2_fill_1 FILLER_66_879 ();
 sg13g2_decap_4 FILLER_66_885 ();
 sg13g2_fill_1 FILLER_66_889 ();
 sg13g2_fill_1 FILLER_66_895 ();
 sg13g2_decap_8 FILLER_66_901 ();
 sg13g2_fill_2 FILLER_66_965 ();
 sg13g2_fill_2 FILLER_66_998 ();
 sg13g2_fill_2 FILLER_66_1037 ();
 sg13g2_fill_1 FILLER_66_1053 ();
 sg13g2_fill_1 FILLER_66_1063 ();
 sg13g2_fill_1 FILLER_66_1129 ();
 sg13g2_decap_8 FILLER_66_1179 ();
 sg13g2_decap_8 FILLER_66_1186 ();
 sg13g2_decap_8 FILLER_66_1193 ();
 sg13g2_decap_8 FILLER_66_1200 ();
 sg13g2_decap_8 FILLER_66_1207 ();
 sg13g2_decap_8 FILLER_66_1214 ();
 sg13g2_decap_8 FILLER_66_1221 ();
 sg13g2_decap_8 FILLER_66_1228 ();
 sg13g2_decap_8 FILLER_66_1235 ();
 sg13g2_decap_8 FILLER_66_1242 ();
 sg13g2_decap_8 FILLER_66_1249 ();
 sg13g2_decap_8 FILLER_66_1256 ();
 sg13g2_decap_8 FILLER_66_1263 ();
 sg13g2_decap_8 FILLER_66_1270 ();
 sg13g2_decap_8 FILLER_66_1277 ();
 sg13g2_decap_8 FILLER_66_1284 ();
 sg13g2_decap_8 FILLER_66_1291 ();
 sg13g2_decap_8 FILLER_66_1298 ();
 sg13g2_decap_8 FILLER_66_1305 ();
 sg13g2_decap_8 FILLER_66_1312 ();
 sg13g2_decap_8 FILLER_66_1319 ();
 sg13g2_decap_8 FILLER_66_1326 ();
 sg13g2_decap_8 FILLER_66_1333 ();
 sg13g2_decap_8 FILLER_66_1340 ();
 sg13g2_decap_8 FILLER_66_1347 ();
 sg13g2_decap_8 FILLER_66_1354 ();
 sg13g2_decap_8 FILLER_66_1361 ();
 sg13g2_decap_8 FILLER_66_1368 ();
 sg13g2_decap_8 FILLER_66_1375 ();
 sg13g2_decap_8 FILLER_66_1382 ();
 sg13g2_decap_8 FILLER_66_1389 ();
 sg13g2_decap_8 FILLER_66_1396 ();
 sg13g2_decap_8 FILLER_66_1403 ();
 sg13g2_decap_8 FILLER_66_1410 ();
 sg13g2_decap_8 FILLER_66_1417 ();
 sg13g2_decap_8 FILLER_66_1424 ();
 sg13g2_decap_8 FILLER_66_1431 ();
 sg13g2_decap_8 FILLER_66_1438 ();
 sg13g2_decap_8 FILLER_66_1445 ();
 sg13g2_decap_8 FILLER_66_1452 ();
 sg13g2_decap_8 FILLER_66_1459 ();
 sg13g2_decap_8 FILLER_66_1466 ();
 sg13g2_decap_8 FILLER_66_1473 ();
 sg13g2_decap_8 FILLER_66_1480 ();
 sg13g2_decap_8 FILLER_66_1487 ();
 sg13g2_decap_8 FILLER_66_1494 ();
 sg13g2_decap_8 FILLER_66_1501 ();
 sg13g2_decap_8 FILLER_66_1508 ();
 sg13g2_decap_8 FILLER_66_1515 ();
 sg13g2_decap_8 FILLER_66_1522 ();
 sg13g2_decap_8 FILLER_66_1529 ();
 sg13g2_decap_8 FILLER_66_1536 ();
 sg13g2_decap_8 FILLER_66_1543 ();
 sg13g2_decap_8 FILLER_66_1550 ();
 sg13g2_decap_8 FILLER_66_1557 ();
 sg13g2_decap_8 FILLER_66_1564 ();
 sg13g2_decap_8 FILLER_66_1571 ();
 sg13g2_decap_8 FILLER_66_1578 ();
 sg13g2_decap_8 FILLER_66_1585 ();
 sg13g2_decap_8 FILLER_66_1592 ();
 sg13g2_decap_8 FILLER_66_1599 ();
 sg13g2_decap_8 FILLER_66_1606 ();
 sg13g2_decap_8 FILLER_66_1613 ();
 sg13g2_decap_8 FILLER_66_1620 ();
 sg13g2_decap_8 FILLER_66_1627 ();
 sg13g2_decap_8 FILLER_66_1634 ();
 sg13g2_decap_8 FILLER_66_1641 ();
 sg13g2_decap_8 FILLER_66_1648 ();
 sg13g2_decap_8 FILLER_66_1655 ();
 sg13g2_decap_8 FILLER_66_1662 ();
 sg13g2_decap_8 FILLER_66_1669 ();
 sg13g2_decap_8 FILLER_66_1676 ();
 sg13g2_decap_8 FILLER_66_1683 ();
 sg13g2_decap_8 FILLER_66_1690 ();
 sg13g2_decap_8 FILLER_66_1697 ();
 sg13g2_decap_8 FILLER_66_1704 ();
 sg13g2_decap_8 FILLER_66_1711 ();
 sg13g2_decap_8 FILLER_66_1718 ();
 sg13g2_decap_8 FILLER_66_1725 ();
 sg13g2_decap_8 FILLER_66_1732 ();
 sg13g2_decap_8 FILLER_66_1739 ();
 sg13g2_decap_8 FILLER_66_1746 ();
 sg13g2_decap_8 FILLER_66_1753 ();
 sg13g2_decap_8 FILLER_66_1760 ();
 sg13g2_fill_1 FILLER_66_1767 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_fill_2 FILLER_67_42 ();
 sg13g2_fill_2 FILLER_67_124 ();
 sg13g2_fill_1 FILLER_67_126 ();
 sg13g2_fill_2 FILLER_67_201 ();
 sg13g2_fill_1 FILLER_67_203 ();
 sg13g2_fill_2 FILLER_67_244 ();
 sg13g2_fill_1 FILLER_67_246 ();
 sg13g2_fill_1 FILLER_67_290 ();
 sg13g2_fill_1 FILLER_67_317 ();
 sg13g2_fill_2 FILLER_67_331 ();
 sg13g2_fill_1 FILLER_67_333 ();
 sg13g2_fill_1 FILLER_67_353 ();
 sg13g2_fill_2 FILLER_67_439 ();
 sg13g2_fill_2 FILLER_67_465 ();
 sg13g2_fill_2 FILLER_67_534 ();
 sg13g2_decap_4 FILLER_67_556 ();
 sg13g2_fill_1 FILLER_67_560 ();
 sg13g2_fill_1 FILLER_67_576 ();
 sg13g2_decap_4 FILLER_67_594 ();
 sg13g2_fill_2 FILLER_67_598 ();
 sg13g2_decap_4 FILLER_67_608 ();
 sg13g2_fill_1 FILLER_67_620 ();
 sg13g2_decap_4 FILLER_67_660 ();
 sg13g2_fill_2 FILLER_67_672 ();
 sg13g2_fill_1 FILLER_67_674 ();
 sg13g2_fill_2 FILLER_67_722 ();
 sg13g2_fill_1 FILLER_67_724 ();
 sg13g2_fill_2 FILLER_67_762 ();
 sg13g2_decap_4 FILLER_67_774 ();
 sg13g2_fill_1 FILLER_67_783 ();
 sg13g2_fill_1 FILLER_67_818 ();
 sg13g2_decap_8 FILLER_67_876 ();
 sg13g2_decap_8 FILLER_67_883 ();
 sg13g2_fill_2 FILLER_67_890 ();
 sg13g2_decap_8 FILLER_67_895 ();
 sg13g2_fill_2 FILLER_67_902 ();
 sg13g2_fill_2 FILLER_67_948 ();
 sg13g2_fill_2 FILLER_67_976 ();
 sg13g2_fill_1 FILLER_67_978 ();
 sg13g2_fill_2 FILLER_67_1083 ();
 sg13g2_fill_2 FILLER_67_1109 ();
 sg13g2_fill_1 FILLER_67_1111 ();
 sg13g2_decap_8 FILLER_67_1184 ();
 sg13g2_decap_8 FILLER_67_1191 ();
 sg13g2_decap_8 FILLER_67_1198 ();
 sg13g2_decap_8 FILLER_67_1205 ();
 sg13g2_decap_8 FILLER_67_1212 ();
 sg13g2_decap_8 FILLER_67_1219 ();
 sg13g2_decap_8 FILLER_67_1226 ();
 sg13g2_decap_8 FILLER_67_1233 ();
 sg13g2_decap_8 FILLER_67_1240 ();
 sg13g2_decap_8 FILLER_67_1247 ();
 sg13g2_decap_8 FILLER_67_1254 ();
 sg13g2_decap_8 FILLER_67_1261 ();
 sg13g2_decap_8 FILLER_67_1268 ();
 sg13g2_decap_8 FILLER_67_1275 ();
 sg13g2_decap_8 FILLER_67_1282 ();
 sg13g2_decap_8 FILLER_67_1289 ();
 sg13g2_decap_8 FILLER_67_1296 ();
 sg13g2_decap_8 FILLER_67_1303 ();
 sg13g2_decap_8 FILLER_67_1310 ();
 sg13g2_decap_8 FILLER_67_1317 ();
 sg13g2_decap_8 FILLER_67_1324 ();
 sg13g2_decap_8 FILLER_67_1331 ();
 sg13g2_decap_8 FILLER_67_1338 ();
 sg13g2_decap_8 FILLER_67_1345 ();
 sg13g2_decap_8 FILLER_67_1352 ();
 sg13g2_decap_8 FILLER_67_1359 ();
 sg13g2_decap_8 FILLER_67_1366 ();
 sg13g2_decap_8 FILLER_67_1373 ();
 sg13g2_decap_8 FILLER_67_1380 ();
 sg13g2_decap_8 FILLER_67_1387 ();
 sg13g2_decap_8 FILLER_67_1394 ();
 sg13g2_decap_8 FILLER_67_1401 ();
 sg13g2_decap_8 FILLER_67_1408 ();
 sg13g2_decap_8 FILLER_67_1415 ();
 sg13g2_decap_8 FILLER_67_1422 ();
 sg13g2_decap_8 FILLER_67_1429 ();
 sg13g2_decap_8 FILLER_67_1436 ();
 sg13g2_decap_8 FILLER_67_1443 ();
 sg13g2_decap_8 FILLER_67_1450 ();
 sg13g2_decap_8 FILLER_67_1457 ();
 sg13g2_decap_8 FILLER_67_1464 ();
 sg13g2_decap_8 FILLER_67_1471 ();
 sg13g2_decap_8 FILLER_67_1478 ();
 sg13g2_decap_8 FILLER_67_1485 ();
 sg13g2_decap_8 FILLER_67_1492 ();
 sg13g2_decap_8 FILLER_67_1499 ();
 sg13g2_decap_8 FILLER_67_1506 ();
 sg13g2_decap_8 FILLER_67_1513 ();
 sg13g2_decap_8 FILLER_67_1520 ();
 sg13g2_decap_8 FILLER_67_1527 ();
 sg13g2_decap_8 FILLER_67_1534 ();
 sg13g2_decap_8 FILLER_67_1541 ();
 sg13g2_decap_8 FILLER_67_1548 ();
 sg13g2_decap_8 FILLER_67_1555 ();
 sg13g2_decap_8 FILLER_67_1562 ();
 sg13g2_decap_8 FILLER_67_1569 ();
 sg13g2_decap_8 FILLER_67_1576 ();
 sg13g2_decap_8 FILLER_67_1583 ();
 sg13g2_decap_8 FILLER_67_1590 ();
 sg13g2_decap_8 FILLER_67_1597 ();
 sg13g2_decap_8 FILLER_67_1604 ();
 sg13g2_decap_8 FILLER_67_1611 ();
 sg13g2_decap_8 FILLER_67_1618 ();
 sg13g2_decap_8 FILLER_67_1625 ();
 sg13g2_decap_8 FILLER_67_1632 ();
 sg13g2_decap_8 FILLER_67_1639 ();
 sg13g2_decap_8 FILLER_67_1646 ();
 sg13g2_decap_8 FILLER_67_1653 ();
 sg13g2_decap_8 FILLER_67_1660 ();
 sg13g2_decap_8 FILLER_67_1667 ();
 sg13g2_decap_8 FILLER_67_1674 ();
 sg13g2_decap_8 FILLER_67_1681 ();
 sg13g2_decap_8 FILLER_67_1688 ();
 sg13g2_decap_8 FILLER_67_1695 ();
 sg13g2_decap_8 FILLER_67_1702 ();
 sg13g2_decap_8 FILLER_67_1709 ();
 sg13g2_decap_8 FILLER_67_1716 ();
 sg13g2_decap_8 FILLER_67_1723 ();
 sg13g2_decap_8 FILLER_67_1730 ();
 sg13g2_decap_8 FILLER_67_1737 ();
 sg13g2_decap_8 FILLER_67_1744 ();
 sg13g2_decap_8 FILLER_67_1751 ();
 sg13g2_decap_8 FILLER_67_1758 ();
 sg13g2_fill_2 FILLER_67_1765 ();
 sg13g2_fill_1 FILLER_67_1767 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_fill_1 FILLER_68_56 ();
 sg13g2_fill_1 FILLER_68_87 ();
 sg13g2_fill_1 FILLER_68_103 ();
 sg13g2_fill_2 FILLER_68_116 ();
 sg13g2_fill_1 FILLER_68_118 ();
 sg13g2_fill_1 FILLER_68_134 ();
 sg13g2_fill_2 FILLER_68_144 ();
 sg13g2_fill_2 FILLER_68_152 ();
 sg13g2_fill_1 FILLER_68_180 ();
 sg13g2_fill_1 FILLER_68_196 ();
 sg13g2_fill_1 FILLER_68_217 ();
 sg13g2_fill_2 FILLER_68_273 ();
 sg13g2_fill_2 FILLER_68_308 ();
 sg13g2_fill_1 FILLER_68_346 ();
 sg13g2_fill_1 FILLER_68_373 ();
 sg13g2_fill_2 FILLER_68_383 ();
 sg13g2_fill_1 FILLER_68_385 ();
 sg13g2_fill_1 FILLER_68_427 ();
 sg13g2_fill_1 FILLER_68_456 ();
 sg13g2_fill_2 FILLER_68_497 ();
 sg13g2_fill_1 FILLER_68_528 ();
 sg13g2_fill_2 FILLER_68_534 ();
 sg13g2_fill_1 FILLER_68_536 ();
 sg13g2_fill_1 FILLER_68_567 ();
 sg13g2_fill_2 FILLER_68_575 ();
 sg13g2_fill_1 FILLER_68_577 ();
 sg13g2_fill_2 FILLER_68_591 ();
 sg13g2_fill_1 FILLER_68_593 ();
 sg13g2_fill_1 FILLER_68_615 ();
 sg13g2_fill_2 FILLER_68_621 ();
 sg13g2_fill_1 FILLER_68_623 ();
 sg13g2_decap_8 FILLER_68_656 ();
 sg13g2_fill_1 FILLER_68_663 ();
 sg13g2_fill_2 FILLER_68_690 ();
 sg13g2_fill_1 FILLER_68_709 ();
 sg13g2_fill_2 FILLER_68_779 ();
 sg13g2_fill_1 FILLER_68_786 ();
 sg13g2_fill_2 FILLER_68_824 ();
 sg13g2_fill_1 FILLER_68_875 ();
 sg13g2_fill_2 FILLER_68_911 ();
 sg13g2_fill_2 FILLER_68_949 ();
 sg13g2_fill_1 FILLER_68_977 ();
 sg13g2_fill_2 FILLER_68_1009 ();
 sg13g2_fill_2 FILLER_68_1133 ();
 sg13g2_fill_1 FILLER_68_1135 ();
 sg13g2_fill_1 FILLER_68_1146 ();
 sg13g2_decap_8 FILLER_68_1182 ();
 sg13g2_decap_8 FILLER_68_1189 ();
 sg13g2_decap_8 FILLER_68_1196 ();
 sg13g2_decap_8 FILLER_68_1203 ();
 sg13g2_decap_8 FILLER_68_1210 ();
 sg13g2_decap_8 FILLER_68_1217 ();
 sg13g2_decap_8 FILLER_68_1224 ();
 sg13g2_decap_8 FILLER_68_1231 ();
 sg13g2_decap_8 FILLER_68_1238 ();
 sg13g2_decap_8 FILLER_68_1245 ();
 sg13g2_decap_8 FILLER_68_1252 ();
 sg13g2_decap_8 FILLER_68_1259 ();
 sg13g2_decap_8 FILLER_68_1266 ();
 sg13g2_decap_8 FILLER_68_1273 ();
 sg13g2_decap_8 FILLER_68_1280 ();
 sg13g2_decap_8 FILLER_68_1287 ();
 sg13g2_decap_8 FILLER_68_1294 ();
 sg13g2_decap_8 FILLER_68_1301 ();
 sg13g2_decap_8 FILLER_68_1308 ();
 sg13g2_decap_8 FILLER_68_1315 ();
 sg13g2_decap_8 FILLER_68_1322 ();
 sg13g2_decap_8 FILLER_68_1329 ();
 sg13g2_decap_8 FILLER_68_1336 ();
 sg13g2_decap_8 FILLER_68_1343 ();
 sg13g2_decap_8 FILLER_68_1350 ();
 sg13g2_decap_8 FILLER_68_1357 ();
 sg13g2_decap_8 FILLER_68_1364 ();
 sg13g2_decap_8 FILLER_68_1371 ();
 sg13g2_decap_8 FILLER_68_1378 ();
 sg13g2_decap_8 FILLER_68_1385 ();
 sg13g2_decap_8 FILLER_68_1392 ();
 sg13g2_decap_8 FILLER_68_1399 ();
 sg13g2_decap_8 FILLER_68_1406 ();
 sg13g2_decap_8 FILLER_68_1413 ();
 sg13g2_decap_8 FILLER_68_1420 ();
 sg13g2_decap_8 FILLER_68_1427 ();
 sg13g2_decap_8 FILLER_68_1434 ();
 sg13g2_decap_8 FILLER_68_1441 ();
 sg13g2_decap_8 FILLER_68_1448 ();
 sg13g2_decap_8 FILLER_68_1455 ();
 sg13g2_decap_8 FILLER_68_1462 ();
 sg13g2_decap_8 FILLER_68_1469 ();
 sg13g2_decap_8 FILLER_68_1476 ();
 sg13g2_decap_8 FILLER_68_1483 ();
 sg13g2_decap_8 FILLER_68_1490 ();
 sg13g2_decap_8 FILLER_68_1497 ();
 sg13g2_decap_8 FILLER_68_1504 ();
 sg13g2_decap_8 FILLER_68_1511 ();
 sg13g2_decap_8 FILLER_68_1518 ();
 sg13g2_decap_8 FILLER_68_1525 ();
 sg13g2_decap_8 FILLER_68_1532 ();
 sg13g2_decap_8 FILLER_68_1539 ();
 sg13g2_decap_8 FILLER_68_1546 ();
 sg13g2_decap_8 FILLER_68_1553 ();
 sg13g2_decap_8 FILLER_68_1560 ();
 sg13g2_decap_8 FILLER_68_1567 ();
 sg13g2_decap_8 FILLER_68_1574 ();
 sg13g2_decap_8 FILLER_68_1581 ();
 sg13g2_decap_8 FILLER_68_1588 ();
 sg13g2_decap_8 FILLER_68_1595 ();
 sg13g2_decap_8 FILLER_68_1602 ();
 sg13g2_decap_8 FILLER_68_1609 ();
 sg13g2_decap_8 FILLER_68_1616 ();
 sg13g2_decap_8 FILLER_68_1623 ();
 sg13g2_decap_8 FILLER_68_1630 ();
 sg13g2_decap_8 FILLER_68_1637 ();
 sg13g2_decap_8 FILLER_68_1644 ();
 sg13g2_decap_8 FILLER_68_1651 ();
 sg13g2_decap_8 FILLER_68_1658 ();
 sg13g2_decap_8 FILLER_68_1665 ();
 sg13g2_decap_8 FILLER_68_1672 ();
 sg13g2_decap_8 FILLER_68_1679 ();
 sg13g2_decap_8 FILLER_68_1686 ();
 sg13g2_decap_8 FILLER_68_1693 ();
 sg13g2_decap_8 FILLER_68_1700 ();
 sg13g2_decap_8 FILLER_68_1707 ();
 sg13g2_decap_8 FILLER_68_1714 ();
 sg13g2_decap_8 FILLER_68_1721 ();
 sg13g2_decap_8 FILLER_68_1728 ();
 sg13g2_decap_8 FILLER_68_1735 ();
 sg13g2_decap_8 FILLER_68_1742 ();
 sg13g2_decap_8 FILLER_68_1749 ();
 sg13g2_decap_8 FILLER_68_1756 ();
 sg13g2_decap_4 FILLER_68_1763 ();
 sg13g2_fill_1 FILLER_68_1767 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_fill_1 FILLER_69_70 ();
 sg13g2_fill_1 FILLER_69_146 ();
 sg13g2_fill_2 FILLER_69_199 ();
 sg13g2_fill_2 FILLER_69_261 ();
 sg13g2_fill_1 FILLER_69_263 ();
 sg13g2_fill_2 FILLER_69_269 ();
 sg13g2_fill_1 FILLER_69_271 ();
 sg13g2_fill_2 FILLER_69_286 ();
 sg13g2_fill_1 FILLER_69_296 ();
 sg13g2_fill_2 FILLER_69_381 ();
 sg13g2_fill_1 FILLER_69_440 ();
 sg13g2_fill_2 FILLER_69_475 ();
 sg13g2_fill_2 FILLER_69_486 ();
 sg13g2_fill_2 FILLER_69_510 ();
 sg13g2_fill_1 FILLER_69_540 ();
 sg13g2_fill_2 FILLER_69_554 ();
 sg13g2_fill_1 FILLER_69_568 ();
 sg13g2_decap_4 FILLER_69_586 ();
 sg13g2_decap_4 FILLER_69_600 ();
 sg13g2_fill_2 FILLER_69_620 ();
 sg13g2_fill_1 FILLER_69_637 ();
 sg13g2_decap_8 FILLER_69_668 ();
 sg13g2_fill_1 FILLER_69_675 ();
 sg13g2_fill_2 FILLER_69_693 ();
 sg13g2_decap_8 FILLER_69_721 ();
 sg13g2_decap_8 FILLER_69_734 ();
 sg13g2_decap_4 FILLER_69_741 ();
 sg13g2_fill_1 FILLER_69_745 ();
 sg13g2_fill_1 FILLER_69_769 ();
 sg13g2_decap_4 FILLER_69_796 ();
 sg13g2_fill_2 FILLER_69_838 ();
 sg13g2_fill_1 FILLER_69_853 ();
 sg13g2_decap_8 FILLER_69_881 ();
 sg13g2_fill_2 FILLER_69_891 ();
 sg13g2_fill_2 FILLER_69_909 ();
 sg13g2_fill_2 FILLER_69_996 ();
 sg13g2_fill_2 FILLER_69_1125 ();
 sg13g2_decap_8 FILLER_69_1174 ();
 sg13g2_decap_8 FILLER_69_1181 ();
 sg13g2_decap_8 FILLER_69_1188 ();
 sg13g2_decap_8 FILLER_69_1195 ();
 sg13g2_decap_8 FILLER_69_1202 ();
 sg13g2_decap_8 FILLER_69_1209 ();
 sg13g2_decap_8 FILLER_69_1216 ();
 sg13g2_decap_8 FILLER_69_1223 ();
 sg13g2_decap_8 FILLER_69_1230 ();
 sg13g2_decap_8 FILLER_69_1237 ();
 sg13g2_decap_8 FILLER_69_1244 ();
 sg13g2_decap_8 FILLER_69_1251 ();
 sg13g2_decap_8 FILLER_69_1258 ();
 sg13g2_decap_8 FILLER_69_1265 ();
 sg13g2_decap_8 FILLER_69_1272 ();
 sg13g2_decap_8 FILLER_69_1279 ();
 sg13g2_decap_8 FILLER_69_1286 ();
 sg13g2_decap_8 FILLER_69_1293 ();
 sg13g2_decap_8 FILLER_69_1300 ();
 sg13g2_decap_8 FILLER_69_1307 ();
 sg13g2_decap_8 FILLER_69_1314 ();
 sg13g2_decap_8 FILLER_69_1321 ();
 sg13g2_decap_8 FILLER_69_1328 ();
 sg13g2_decap_8 FILLER_69_1335 ();
 sg13g2_decap_8 FILLER_69_1342 ();
 sg13g2_decap_8 FILLER_69_1349 ();
 sg13g2_decap_8 FILLER_69_1356 ();
 sg13g2_decap_8 FILLER_69_1363 ();
 sg13g2_decap_8 FILLER_69_1370 ();
 sg13g2_decap_8 FILLER_69_1377 ();
 sg13g2_decap_8 FILLER_69_1384 ();
 sg13g2_decap_8 FILLER_69_1391 ();
 sg13g2_decap_8 FILLER_69_1398 ();
 sg13g2_decap_8 FILLER_69_1405 ();
 sg13g2_decap_8 FILLER_69_1412 ();
 sg13g2_decap_8 FILLER_69_1419 ();
 sg13g2_decap_8 FILLER_69_1426 ();
 sg13g2_decap_8 FILLER_69_1433 ();
 sg13g2_decap_8 FILLER_69_1440 ();
 sg13g2_decap_8 FILLER_69_1447 ();
 sg13g2_decap_8 FILLER_69_1454 ();
 sg13g2_decap_8 FILLER_69_1461 ();
 sg13g2_decap_8 FILLER_69_1468 ();
 sg13g2_decap_8 FILLER_69_1475 ();
 sg13g2_decap_8 FILLER_69_1482 ();
 sg13g2_decap_8 FILLER_69_1489 ();
 sg13g2_decap_8 FILLER_69_1496 ();
 sg13g2_decap_8 FILLER_69_1503 ();
 sg13g2_decap_8 FILLER_69_1510 ();
 sg13g2_decap_8 FILLER_69_1517 ();
 sg13g2_decap_8 FILLER_69_1524 ();
 sg13g2_decap_8 FILLER_69_1531 ();
 sg13g2_decap_8 FILLER_69_1538 ();
 sg13g2_decap_8 FILLER_69_1545 ();
 sg13g2_decap_8 FILLER_69_1552 ();
 sg13g2_decap_8 FILLER_69_1559 ();
 sg13g2_decap_8 FILLER_69_1566 ();
 sg13g2_decap_8 FILLER_69_1573 ();
 sg13g2_decap_8 FILLER_69_1580 ();
 sg13g2_decap_8 FILLER_69_1587 ();
 sg13g2_decap_8 FILLER_69_1594 ();
 sg13g2_decap_8 FILLER_69_1601 ();
 sg13g2_decap_8 FILLER_69_1608 ();
 sg13g2_decap_8 FILLER_69_1615 ();
 sg13g2_decap_8 FILLER_69_1622 ();
 sg13g2_decap_8 FILLER_69_1629 ();
 sg13g2_decap_8 FILLER_69_1636 ();
 sg13g2_decap_8 FILLER_69_1643 ();
 sg13g2_decap_8 FILLER_69_1650 ();
 sg13g2_decap_8 FILLER_69_1657 ();
 sg13g2_decap_8 FILLER_69_1664 ();
 sg13g2_decap_8 FILLER_69_1671 ();
 sg13g2_decap_8 FILLER_69_1678 ();
 sg13g2_decap_8 FILLER_69_1685 ();
 sg13g2_decap_8 FILLER_69_1692 ();
 sg13g2_decap_8 FILLER_69_1699 ();
 sg13g2_decap_8 FILLER_69_1706 ();
 sg13g2_decap_8 FILLER_69_1713 ();
 sg13g2_decap_8 FILLER_69_1720 ();
 sg13g2_decap_8 FILLER_69_1727 ();
 sg13g2_decap_8 FILLER_69_1734 ();
 sg13g2_decap_8 FILLER_69_1741 ();
 sg13g2_decap_8 FILLER_69_1748 ();
 sg13g2_decap_8 FILLER_69_1755 ();
 sg13g2_decap_4 FILLER_69_1762 ();
 sg13g2_fill_2 FILLER_69_1766 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_fill_2 FILLER_70_14 ();
 sg13g2_fill_1 FILLER_70_16 ();
 sg13g2_fill_1 FILLER_70_43 ();
 sg13g2_fill_1 FILLER_70_47 ();
 sg13g2_decap_4 FILLER_70_56 ();
 sg13g2_fill_2 FILLER_70_60 ();
 sg13g2_fill_1 FILLER_70_126 ();
 sg13g2_fill_2 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_135 ();
 sg13g2_fill_1 FILLER_70_159 ();
 sg13g2_fill_2 FILLER_70_231 ();
 sg13g2_fill_1 FILLER_70_233 ();
 sg13g2_fill_2 FILLER_70_252 ();
 sg13g2_fill_1 FILLER_70_254 ();
 sg13g2_fill_2 FILLER_70_261 ();
 sg13g2_fill_2 FILLER_70_268 ();
 sg13g2_fill_2 FILLER_70_296 ();
 sg13g2_fill_1 FILLER_70_530 ();
 sg13g2_decap_4 FILLER_70_635 ();
 sg13g2_fill_2 FILLER_70_721 ();
 sg13g2_fill_1 FILLER_70_723 ();
 sg13g2_fill_2 FILLER_70_769 ();
 sg13g2_fill_1 FILLER_70_808 ();
 sg13g2_fill_1 FILLER_70_834 ();
 sg13g2_fill_1 FILLER_70_840 ();
 sg13g2_fill_2 FILLER_70_867 ();
 sg13g2_fill_1 FILLER_70_869 ();
 sg13g2_decap_4 FILLER_70_875 ();
 sg13g2_fill_2 FILLER_70_879 ();
 sg13g2_fill_2 FILLER_70_965 ();
 sg13g2_fill_1 FILLER_70_1060 ();
 sg13g2_fill_1 FILLER_70_1135 ();
 sg13g2_fill_2 FILLER_70_1146 ();
 sg13g2_fill_1 FILLER_70_1148 ();
 sg13g2_decap_8 FILLER_70_1180 ();
 sg13g2_decap_8 FILLER_70_1187 ();
 sg13g2_decap_8 FILLER_70_1194 ();
 sg13g2_decap_8 FILLER_70_1201 ();
 sg13g2_decap_8 FILLER_70_1208 ();
 sg13g2_decap_8 FILLER_70_1215 ();
 sg13g2_decap_8 FILLER_70_1222 ();
 sg13g2_decap_8 FILLER_70_1229 ();
 sg13g2_decap_8 FILLER_70_1236 ();
 sg13g2_decap_8 FILLER_70_1243 ();
 sg13g2_decap_8 FILLER_70_1250 ();
 sg13g2_decap_8 FILLER_70_1257 ();
 sg13g2_decap_8 FILLER_70_1264 ();
 sg13g2_decap_8 FILLER_70_1271 ();
 sg13g2_decap_8 FILLER_70_1278 ();
 sg13g2_decap_8 FILLER_70_1285 ();
 sg13g2_decap_8 FILLER_70_1292 ();
 sg13g2_decap_8 FILLER_70_1299 ();
 sg13g2_decap_8 FILLER_70_1306 ();
 sg13g2_decap_8 FILLER_70_1313 ();
 sg13g2_decap_8 FILLER_70_1320 ();
 sg13g2_decap_8 FILLER_70_1327 ();
 sg13g2_decap_8 FILLER_70_1334 ();
 sg13g2_decap_8 FILLER_70_1341 ();
 sg13g2_decap_8 FILLER_70_1348 ();
 sg13g2_decap_8 FILLER_70_1355 ();
 sg13g2_decap_8 FILLER_70_1362 ();
 sg13g2_decap_8 FILLER_70_1369 ();
 sg13g2_decap_8 FILLER_70_1376 ();
 sg13g2_decap_8 FILLER_70_1383 ();
 sg13g2_decap_8 FILLER_70_1390 ();
 sg13g2_decap_8 FILLER_70_1397 ();
 sg13g2_decap_8 FILLER_70_1404 ();
 sg13g2_decap_8 FILLER_70_1411 ();
 sg13g2_decap_8 FILLER_70_1418 ();
 sg13g2_decap_8 FILLER_70_1425 ();
 sg13g2_decap_8 FILLER_70_1432 ();
 sg13g2_decap_8 FILLER_70_1439 ();
 sg13g2_decap_8 FILLER_70_1446 ();
 sg13g2_decap_8 FILLER_70_1453 ();
 sg13g2_decap_8 FILLER_70_1460 ();
 sg13g2_decap_8 FILLER_70_1467 ();
 sg13g2_decap_8 FILLER_70_1474 ();
 sg13g2_decap_8 FILLER_70_1481 ();
 sg13g2_decap_8 FILLER_70_1488 ();
 sg13g2_decap_8 FILLER_70_1495 ();
 sg13g2_decap_8 FILLER_70_1502 ();
 sg13g2_decap_8 FILLER_70_1509 ();
 sg13g2_decap_8 FILLER_70_1516 ();
 sg13g2_decap_8 FILLER_70_1523 ();
 sg13g2_decap_8 FILLER_70_1530 ();
 sg13g2_decap_8 FILLER_70_1537 ();
 sg13g2_decap_8 FILLER_70_1544 ();
 sg13g2_decap_8 FILLER_70_1551 ();
 sg13g2_decap_8 FILLER_70_1558 ();
 sg13g2_decap_8 FILLER_70_1565 ();
 sg13g2_decap_8 FILLER_70_1572 ();
 sg13g2_decap_8 FILLER_70_1579 ();
 sg13g2_decap_8 FILLER_70_1586 ();
 sg13g2_decap_8 FILLER_70_1593 ();
 sg13g2_decap_8 FILLER_70_1600 ();
 sg13g2_decap_8 FILLER_70_1607 ();
 sg13g2_decap_8 FILLER_70_1614 ();
 sg13g2_decap_8 FILLER_70_1621 ();
 sg13g2_decap_8 FILLER_70_1628 ();
 sg13g2_decap_8 FILLER_70_1635 ();
 sg13g2_decap_8 FILLER_70_1642 ();
 sg13g2_decap_8 FILLER_70_1649 ();
 sg13g2_decap_8 FILLER_70_1656 ();
 sg13g2_decap_8 FILLER_70_1663 ();
 sg13g2_decap_8 FILLER_70_1670 ();
 sg13g2_decap_8 FILLER_70_1677 ();
 sg13g2_decap_8 FILLER_70_1684 ();
 sg13g2_decap_8 FILLER_70_1691 ();
 sg13g2_decap_8 FILLER_70_1698 ();
 sg13g2_decap_8 FILLER_70_1705 ();
 sg13g2_decap_8 FILLER_70_1712 ();
 sg13g2_decap_8 FILLER_70_1719 ();
 sg13g2_decap_8 FILLER_70_1726 ();
 sg13g2_decap_8 FILLER_70_1733 ();
 sg13g2_decap_8 FILLER_70_1740 ();
 sg13g2_decap_8 FILLER_70_1747 ();
 sg13g2_decap_8 FILLER_70_1754 ();
 sg13g2_decap_8 FILLER_70_1761 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_fill_2 FILLER_71_21 ();
 sg13g2_fill_1 FILLER_71_23 ();
 sg13g2_fill_1 FILLER_71_27 ();
 sg13g2_fill_1 FILLER_71_135 ();
 sg13g2_fill_2 FILLER_71_162 ();
 sg13g2_fill_1 FILLER_71_164 ();
 sg13g2_fill_1 FILLER_71_185 ();
 sg13g2_fill_1 FILLER_71_192 ();
 sg13g2_fill_2 FILLER_71_215 ();
 sg13g2_fill_1 FILLER_71_217 ();
 sg13g2_fill_2 FILLER_71_254 ();
 sg13g2_decap_8 FILLER_71_286 ();
 sg13g2_fill_1 FILLER_71_310 ();
 sg13g2_fill_2 FILLER_71_411 ();
 sg13g2_fill_1 FILLER_71_413 ();
 sg13g2_fill_2 FILLER_71_441 ();
 sg13g2_fill_2 FILLER_71_471 ();
 sg13g2_fill_1 FILLER_71_496 ();
 sg13g2_fill_1 FILLER_71_556 ();
 sg13g2_fill_1 FILLER_71_572 ();
 sg13g2_fill_1 FILLER_71_595 ();
 sg13g2_decap_4 FILLER_71_631 ();
 sg13g2_fill_1 FILLER_71_713 ();
 sg13g2_fill_1 FILLER_71_731 ();
 sg13g2_fill_2 FILLER_71_810 ();
 sg13g2_fill_2 FILLER_71_863 ();
 sg13g2_fill_1 FILLER_71_865 ();
 sg13g2_decap_8 FILLER_71_874 ();
 sg13g2_decap_8 FILLER_71_881 ();
 sg13g2_fill_2 FILLER_71_940 ();
 sg13g2_fill_2 FILLER_71_970 ();
 sg13g2_fill_2 FILLER_71_1037 ();
 sg13g2_fill_2 FILLER_71_1119 ();
 sg13g2_fill_1 FILLER_71_1146 ();
 sg13g2_decap_8 FILLER_71_1173 ();
 sg13g2_decap_8 FILLER_71_1180 ();
 sg13g2_decap_8 FILLER_71_1187 ();
 sg13g2_decap_8 FILLER_71_1194 ();
 sg13g2_decap_8 FILLER_71_1201 ();
 sg13g2_decap_8 FILLER_71_1208 ();
 sg13g2_decap_8 FILLER_71_1215 ();
 sg13g2_decap_8 FILLER_71_1222 ();
 sg13g2_decap_8 FILLER_71_1229 ();
 sg13g2_decap_8 FILLER_71_1236 ();
 sg13g2_decap_8 FILLER_71_1243 ();
 sg13g2_decap_8 FILLER_71_1250 ();
 sg13g2_decap_8 FILLER_71_1257 ();
 sg13g2_decap_8 FILLER_71_1264 ();
 sg13g2_decap_8 FILLER_71_1271 ();
 sg13g2_decap_8 FILLER_71_1278 ();
 sg13g2_decap_8 FILLER_71_1285 ();
 sg13g2_decap_8 FILLER_71_1292 ();
 sg13g2_decap_8 FILLER_71_1299 ();
 sg13g2_decap_8 FILLER_71_1306 ();
 sg13g2_decap_8 FILLER_71_1313 ();
 sg13g2_decap_8 FILLER_71_1320 ();
 sg13g2_decap_8 FILLER_71_1327 ();
 sg13g2_decap_8 FILLER_71_1334 ();
 sg13g2_decap_8 FILLER_71_1341 ();
 sg13g2_decap_8 FILLER_71_1348 ();
 sg13g2_decap_8 FILLER_71_1355 ();
 sg13g2_decap_8 FILLER_71_1362 ();
 sg13g2_decap_8 FILLER_71_1369 ();
 sg13g2_decap_8 FILLER_71_1376 ();
 sg13g2_decap_8 FILLER_71_1383 ();
 sg13g2_decap_8 FILLER_71_1390 ();
 sg13g2_decap_8 FILLER_71_1397 ();
 sg13g2_decap_8 FILLER_71_1404 ();
 sg13g2_decap_8 FILLER_71_1411 ();
 sg13g2_decap_8 FILLER_71_1418 ();
 sg13g2_decap_8 FILLER_71_1425 ();
 sg13g2_decap_8 FILLER_71_1432 ();
 sg13g2_decap_8 FILLER_71_1439 ();
 sg13g2_decap_8 FILLER_71_1446 ();
 sg13g2_decap_8 FILLER_71_1453 ();
 sg13g2_decap_8 FILLER_71_1460 ();
 sg13g2_decap_8 FILLER_71_1467 ();
 sg13g2_decap_8 FILLER_71_1474 ();
 sg13g2_decap_8 FILLER_71_1481 ();
 sg13g2_decap_8 FILLER_71_1488 ();
 sg13g2_decap_8 FILLER_71_1495 ();
 sg13g2_decap_8 FILLER_71_1502 ();
 sg13g2_decap_8 FILLER_71_1509 ();
 sg13g2_decap_8 FILLER_71_1516 ();
 sg13g2_decap_8 FILLER_71_1523 ();
 sg13g2_decap_8 FILLER_71_1530 ();
 sg13g2_decap_8 FILLER_71_1537 ();
 sg13g2_decap_8 FILLER_71_1544 ();
 sg13g2_decap_8 FILLER_71_1551 ();
 sg13g2_decap_8 FILLER_71_1558 ();
 sg13g2_decap_8 FILLER_71_1565 ();
 sg13g2_decap_8 FILLER_71_1572 ();
 sg13g2_decap_8 FILLER_71_1579 ();
 sg13g2_decap_8 FILLER_71_1586 ();
 sg13g2_decap_8 FILLER_71_1593 ();
 sg13g2_decap_8 FILLER_71_1600 ();
 sg13g2_decap_8 FILLER_71_1607 ();
 sg13g2_decap_8 FILLER_71_1614 ();
 sg13g2_decap_8 FILLER_71_1621 ();
 sg13g2_decap_8 FILLER_71_1628 ();
 sg13g2_decap_8 FILLER_71_1635 ();
 sg13g2_decap_8 FILLER_71_1642 ();
 sg13g2_decap_8 FILLER_71_1649 ();
 sg13g2_decap_8 FILLER_71_1656 ();
 sg13g2_decap_8 FILLER_71_1663 ();
 sg13g2_decap_8 FILLER_71_1670 ();
 sg13g2_decap_8 FILLER_71_1677 ();
 sg13g2_decap_8 FILLER_71_1684 ();
 sg13g2_decap_8 FILLER_71_1691 ();
 sg13g2_decap_8 FILLER_71_1698 ();
 sg13g2_decap_8 FILLER_71_1705 ();
 sg13g2_decap_8 FILLER_71_1712 ();
 sg13g2_decap_8 FILLER_71_1719 ();
 sg13g2_decap_8 FILLER_71_1726 ();
 sg13g2_decap_8 FILLER_71_1733 ();
 sg13g2_decap_8 FILLER_71_1740 ();
 sg13g2_decap_8 FILLER_71_1747 ();
 sg13g2_decap_8 FILLER_71_1754 ();
 sg13g2_decap_8 FILLER_71_1761 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_4 FILLER_72_14 ();
 sg13g2_fill_2 FILLER_72_18 ();
 sg13g2_decap_4 FILLER_72_23 ();
 sg13g2_fill_2 FILLER_72_27 ();
 sg13g2_fill_1 FILLER_72_36 ();
 sg13g2_fill_1 FILLER_72_51 ();
 sg13g2_fill_2 FILLER_72_143 ();
 sg13g2_fill_2 FILLER_72_202 ();
 sg13g2_fill_1 FILLER_72_209 ();
 sg13g2_fill_1 FILLER_72_215 ();
 sg13g2_fill_1 FILLER_72_238 ();
 sg13g2_fill_2 FILLER_72_344 ();
 sg13g2_fill_1 FILLER_72_346 ();
 sg13g2_fill_2 FILLER_72_430 ();
 sg13g2_fill_2 FILLER_72_492 ();
 sg13g2_fill_1 FILLER_72_494 ();
 sg13g2_fill_2 FILLER_72_547 ();
 sg13g2_fill_1 FILLER_72_549 ();
 sg13g2_fill_1 FILLER_72_624 ();
 sg13g2_decap_4 FILLER_72_651 ();
 sg13g2_fill_1 FILLER_72_726 ();
 sg13g2_fill_2 FILLER_72_769 ();
 sg13g2_fill_1 FILLER_72_771 ();
 sg13g2_fill_1 FILLER_72_815 ();
 sg13g2_decap_8 FILLER_72_868 ();
 sg13g2_decap_4 FILLER_72_875 ();
 sg13g2_fill_1 FILLER_72_882 ();
 sg13g2_fill_2 FILLER_72_909 ();
 sg13g2_fill_2 FILLER_72_980 ();
 sg13g2_fill_2 FILLER_72_1031 ();
 sg13g2_fill_1 FILLER_72_1056 ();
 sg13g2_fill_2 FILLER_72_1119 ();
 sg13g2_decap_8 FILLER_72_1174 ();
 sg13g2_decap_8 FILLER_72_1181 ();
 sg13g2_decap_8 FILLER_72_1188 ();
 sg13g2_decap_8 FILLER_72_1195 ();
 sg13g2_decap_8 FILLER_72_1202 ();
 sg13g2_decap_8 FILLER_72_1209 ();
 sg13g2_decap_8 FILLER_72_1216 ();
 sg13g2_decap_8 FILLER_72_1223 ();
 sg13g2_decap_8 FILLER_72_1230 ();
 sg13g2_decap_8 FILLER_72_1237 ();
 sg13g2_decap_8 FILLER_72_1244 ();
 sg13g2_decap_8 FILLER_72_1251 ();
 sg13g2_decap_8 FILLER_72_1258 ();
 sg13g2_decap_8 FILLER_72_1265 ();
 sg13g2_decap_8 FILLER_72_1272 ();
 sg13g2_decap_8 FILLER_72_1279 ();
 sg13g2_decap_8 FILLER_72_1286 ();
 sg13g2_decap_8 FILLER_72_1293 ();
 sg13g2_decap_8 FILLER_72_1300 ();
 sg13g2_decap_8 FILLER_72_1307 ();
 sg13g2_decap_8 FILLER_72_1314 ();
 sg13g2_decap_8 FILLER_72_1321 ();
 sg13g2_decap_8 FILLER_72_1328 ();
 sg13g2_decap_8 FILLER_72_1335 ();
 sg13g2_decap_8 FILLER_72_1342 ();
 sg13g2_decap_8 FILLER_72_1349 ();
 sg13g2_decap_8 FILLER_72_1356 ();
 sg13g2_decap_8 FILLER_72_1363 ();
 sg13g2_decap_8 FILLER_72_1370 ();
 sg13g2_decap_8 FILLER_72_1377 ();
 sg13g2_decap_8 FILLER_72_1384 ();
 sg13g2_decap_8 FILLER_72_1391 ();
 sg13g2_decap_8 FILLER_72_1398 ();
 sg13g2_decap_8 FILLER_72_1405 ();
 sg13g2_decap_8 FILLER_72_1412 ();
 sg13g2_decap_8 FILLER_72_1419 ();
 sg13g2_decap_8 FILLER_72_1426 ();
 sg13g2_decap_8 FILLER_72_1433 ();
 sg13g2_decap_8 FILLER_72_1440 ();
 sg13g2_decap_8 FILLER_72_1447 ();
 sg13g2_decap_8 FILLER_72_1454 ();
 sg13g2_decap_8 FILLER_72_1461 ();
 sg13g2_decap_8 FILLER_72_1468 ();
 sg13g2_decap_8 FILLER_72_1475 ();
 sg13g2_decap_8 FILLER_72_1482 ();
 sg13g2_decap_8 FILLER_72_1489 ();
 sg13g2_decap_8 FILLER_72_1496 ();
 sg13g2_decap_8 FILLER_72_1503 ();
 sg13g2_decap_8 FILLER_72_1510 ();
 sg13g2_decap_8 FILLER_72_1517 ();
 sg13g2_decap_8 FILLER_72_1524 ();
 sg13g2_decap_8 FILLER_72_1531 ();
 sg13g2_decap_8 FILLER_72_1538 ();
 sg13g2_decap_8 FILLER_72_1545 ();
 sg13g2_decap_8 FILLER_72_1552 ();
 sg13g2_decap_8 FILLER_72_1559 ();
 sg13g2_decap_8 FILLER_72_1566 ();
 sg13g2_decap_8 FILLER_72_1573 ();
 sg13g2_decap_8 FILLER_72_1580 ();
 sg13g2_decap_8 FILLER_72_1587 ();
 sg13g2_decap_8 FILLER_72_1594 ();
 sg13g2_decap_8 FILLER_72_1601 ();
 sg13g2_decap_8 FILLER_72_1608 ();
 sg13g2_decap_8 FILLER_72_1615 ();
 sg13g2_decap_8 FILLER_72_1622 ();
 sg13g2_decap_8 FILLER_72_1629 ();
 sg13g2_decap_8 FILLER_72_1636 ();
 sg13g2_decap_8 FILLER_72_1643 ();
 sg13g2_decap_8 FILLER_72_1650 ();
 sg13g2_decap_8 FILLER_72_1657 ();
 sg13g2_decap_8 FILLER_72_1664 ();
 sg13g2_decap_8 FILLER_72_1671 ();
 sg13g2_decap_8 FILLER_72_1678 ();
 sg13g2_decap_8 FILLER_72_1685 ();
 sg13g2_decap_8 FILLER_72_1692 ();
 sg13g2_decap_8 FILLER_72_1699 ();
 sg13g2_decap_8 FILLER_72_1706 ();
 sg13g2_decap_8 FILLER_72_1713 ();
 sg13g2_decap_8 FILLER_72_1720 ();
 sg13g2_decap_8 FILLER_72_1727 ();
 sg13g2_decap_8 FILLER_72_1734 ();
 sg13g2_decap_8 FILLER_72_1741 ();
 sg13g2_decap_8 FILLER_72_1748 ();
 sg13g2_decap_8 FILLER_72_1755 ();
 sg13g2_decap_4 FILLER_72_1762 ();
 sg13g2_fill_2 FILLER_72_1766 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_4 FILLER_73_7 ();
 sg13g2_fill_2 FILLER_73_11 ();
 sg13g2_fill_2 FILLER_73_39 ();
 sg13g2_fill_2 FILLER_73_67 ();
 sg13g2_fill_1 FILLER_73_91 ();
 sg13g2_fill_2 FILLER_73_158 ();
 sg13g2_fill_1 FILLER_73_178 ();
 sg13g2_fill_1 FILLER_73_199 ();
 sg13g2_fill_2 FILLER_73_206 ();
 sg13g2_fill_1 FILLER_73_208 ();
 sg13g2_fill_2 FILLER_73_241 ();
 sg13g2_fill_2 FILLER_73_253 ();
 sg13g2_fill_2 FILLER_73_302 ();
 sg13g2_fill_2 FILLER_73_453 ();
 sg13g2_fill_1 FILLER_73_455 ();
 sg13g2_fill_2 FILLER_73_465 ();
 sg13g2_fill_1 FILLER_73_467 ();
 sg13g2_fill_2 FILLER_73_472 ();
 sg13g2_fill_1 FILLER_73_474 ();
 sg13g2_fill_2 FILLER_73_490 ();
 sg13g2_fill_2 FILLER_73_508 ();
 sg13g2_fill_2 FILLER_73_539 ();
 sg13g2_decap_8 FILLER_73_567 ();
 sg13g2_decap_4 FILLER_73_574 ();
 sg13g2_fill_2 FILLER_73_578 ();
 sg13g2_fill_2 FILLER_73_589 ();
 sg13g2_decap_4 FILLER_73_599 ();
 sg13g2_fill_1 FILLER_73_621 ();
 sg13g2_decap_8 FILLER_73_631 ();
 sg13g2_fill_2 FILLER_73_661 ();
 sg13g2_fill_2 FILLER_73_677 ();
 sg13g2_fill_1 FILLER_73_683 ();
 sg13g2_fill_2 FILLER_73_706 ();
 sg13g2_fill_2 FILLER_73_724 ();
 sg13g2_fill_1 FILLER_73_726 ();
 sg13g2_fill_1 FILLER_73_748 ();
 sg13g2_fill_2 FILLER_73_776 ();
 sg13g2_fill_1 FILLER_73_778 ();
 sg13g2_fill_2 FILLER_73_797 ();
 sg13g2_fill_1 FILLER_73_799 ();
 sg13g2_fill_2 FILLER_73_870 ();
 sg13g2_fill_1 FILLER_73_879 ();
 sg13g2_fill_2 FILLER_73_887 ();
 sg13g2_fill_2 FILLER_73_900 ();
 sg13g2_fill_1 FILLER_73_944 ();
 sg13g2_fill_1 FILLER_73_954 ();
 sg13g2_fill_1 FILLER_73_1004 ();
 sg13g2_fill_2 FILLER_73_1039 ();
 sg13g2_fill_2 FILLER_73_1067 ();
 sg13g2_decap_8 FILLER_73_1152 ();
 sg13g2_decap_8 FILLER_73_1159 ();
 sg13g2_decap_8 FILLER_73_1166 ();
 sg13g2_decap_8 FILLER_73_1173 ();
 sg13g2_decap_8 FILLER_73_1180 ();
 sg13g2_decap_8 FILLER_73_1187 ();
 sg13g2_decap_8 FILLER_73_1194 ();
 sg13g2_decap_8 FILLER_73_1201 ();
 sg13g2_decap_8 FILLER_73_1208 ();
 sg13g2_decap_8 FILLER_73_1215 ();
 sg13g2_decap_8 FILLER_73_1222 ();
 sg13g2_decap_8 FILLER_73_1229 ();
 sg13g2_decap_8 FILLER_73_1236 ();
 sg13g2_decap_8 FILLER_73_1243 ();
 sg13g2_decap_8 FILLER_73_1250 ();
 sg13g2_decap_8 FILLER_73_1257 ();
 sg13g2_decap_8 FILLER_73_1264 ();
 sg13g2_decap_8 FILLER_73_1271 ();
 sg13g2_decap_8 FILLER_73_1278 ();
 sg13g2_decap_8 FILLER_73_1285 ();
 sg13g2_decap_8 FILLER_73_1292 ();
 sg13g2_decap_8 FILLER_73_1299 ();
 sg13g2_decap_8 FILLER_73_1306 ();
 sg13g2_decap_8 FILLER_73_1313 ();
 sg13g2_decap_8 FILLER_73_1320 ();
 sg13g2_decap_8 FILLER_73_1327 ();
 sg13g2_decap_8 FILLER_73_1334 ();
 sg13g2_decap_8 FILLER_73_1341 ();
 sg13g2_decap_8 FILLER_73_1348 ();
 sg13g2_decap_8 FILLER_73_1355 ();
 sg13g2_decap_8 FILLER_73_1362 ();
 sg13g2_decap_8 FILLER_73_1369 ();
 sg13g2_decap_8 FILLER_73_1376 ();
 sg13g2_decap_8 FILLER_73_1383 ();
 sg13g2_decap_8 FILLER_73_1390 ();
 sg13g2_decap_8 FILLER_73_1397 ();
 sg13g2_decap_8 FILLER_73_1404 ();
 sg13g2_decap_8 FILLER_73_1411 ();
 sg13g2_decap_8 FILLER_73_1418 ();
 sg13g2_decap_8 FILLER_73_1425 ();
 sg13g2_decap_8 FILLER_73_1432 ();
 sg13g2_decap_8 FILLER_73_1439 ();
 sg13g2_decap_8 FILLER_73_1446 ();
 sg13g2_decap_8 FILLER_73_1453 ();
 sg13g2_decap_8 FILLER_73_1460 ();
 sg13g2_decap_8 FILLER_73_1467 ();
 sg13g2_decap_8 FILLER_73_1474 ();
 sg13g2_decap_8 FILLER_73_1481 ();
 sg13g2_decap_8 FILLER_73_1488 ();
 sg13g2_decap_8 FILLER_73_1495 ();
 sg13g2_decap_8 FILLER_73_1502 ();
 sg13g2_decap_8 FILLER_73_1509 ();
 sg13g2_decap_8 FILLER_73_1516 ();
 sg13g2_decap_8 FILLER_73_1523 ();
 sg13g2_decap_8 FILLER_73_1530 ();
 sg13g2_decap_8 FILLER_73_1537 ();
 sg13g2_decap_8 FILLER_73_1544 ();
 sg13g2_decap_8 FILLER_73_1551 ();
 sg13g2_decap_8 FILLER_73_1558 ();
 sg13g2_decap_8 FILLER_73_1565 ();
 sg13g2_decap_8 FILLER_73_1572 ();
 sg13g2_decap_8 FILLER_73_1579 ();
 sg13g2_decap_8 FILLER_73_1586 ();
 sg13g2_decap_8 FILLER_73_1593 ();
 sg13g2_decap_8 FILLER_73_1600 ();
 sg13g2_decap_8 FILLER_73_1607 ();
 sg13g2_decap_8 FILLER_73_1614 ();
 sg13g2_decap_8 FILLER_73_1621 ();
 sg13g2_decap_8 FILLER_73_1628 ();
 sg13g2_decap_8 FILLER_73_1635 ();
 sg13g2_decap_8 FILLER_73_1642 ();
 sg13g2_decap_8 FILLER_73_1649 ();
 sg13g2_decap_8 FILLER_73_1656 ();
 sg13g2_decap_8 FILLER_73_1663 ();
 sg13g2_decap_8 FILLER_73_1670 ();
 sg13g2_decap_8 FILLER_73_1677 ();
 sg13g2_decap_8 FILLER_73_1684 ();
 sg13g2_decap_8 FILLER_73_1691 ();
 sg13g2_decap_8 FILLER_73_1698 ();
 sg13g2_decap_8 FILLER_73_1705 ();
 sg13g2_decap_8 FILLER_73_1712 ();
 sg13g2_decap_8 FILLER_73_1719 ();
 sg13g2_decap_8 FILLER_73_1726 ();
 sg13g2_decap_8 FILLER_73_1733 ();
 sg13g2_decap_8 FILLER_73_1740 ();
 sg13g2_decap_8 FILLER_73_1747 ();
 sg13g2_decap_8 FILLER_73_1754 ();
 sg13g2_decap_8 FILLER_73_1761 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_28 ();
 sg13g2_fill_1 FILLER_74_107 ();
 sg13g2_fill_1 FILLER_74_140 ();
 sg13g2_fill_2 FILLER_74_155 ();
 sg13g2_fill_1 FILLER_74_157 ();
 sg13g2_fill_1 FILLER_74_186 ();
 sg13g2_fill_1 FILLER_74_197 ();
 sg13g2_fill_2 FILLER_74_203 ();
 sg13g2_fill_1 FILLER_74_205 ();
 sg13g2_fill_2 FILLER_74_220 ();
 sg13g2_fill_2 FILLER_74_247 ();
 sg13g2_fill_2 FILLER_74_261 ();
 sg13g2_fill_2 FILLER_74_273 ();
 sg13g2_fill_1 FILLER_74_327 ();
 sg13g2_fill_1 FILLER_74_337 ();
 sg13g2_fill_1 FILLER_74_371 ();
 sg13g2_fill_2 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_74_460 ();
 sg13g2_fill_2 FILLER_74_467 ();
 sg13g2_fill_1 FILLER_74_469 ();
 sg13g2_fill_2 FILLER_74_509 ();
 sg13g2_fill_1 FILLER_74_511 ();
 sg13g2_fill_2 FILLER_74_557 ();
 sg13g2_fill_1 FILLER_74_563 ();
 sg13g2_decap_8 FILLER_74_567 ();
 sg13g2_fill_2 FILLER_74_599 ();
 sg13g2_decap_4 FILLER_74_646 ();
 sg13g2_fill_1 FILLER_74_650 ();
 sg13g2_decap_8 FILLER_74_666 ();
 sg13g2_fill_2 FILLER_74_694 ();
 sg13g2_decap_4 FILLER_74_701 ();
 sg13g2_fill_2 FILLER_74_705 ();
 sg13g2_fill_2 FILLER_74_725 ();
 sg13g2_fill_1 FILLER_74_773 ();
 sg13g2_fill_2 FILLER_74_802 ();
 sg13g2_fill_1 FILLER_74_827 ();
 sg13g2_fill_2 FILLER_74_851 ();
 sg13g2_fill_1 FILLER_74_879 ();
 sg13g2_fill_1 FILLER_74_900 ();
 sg13g2_fill_2 FILLER_74_909 ();
 sg13g2_fill_2 FILLER_74_963 ();
 sg13g2_fill_2 FILLER_74_1003 ();
 sg13g2_fill_1 FILLER_74_1051 ();
 sg13g2_fill_2 FILLER_74_1077 ();
 sg13g2_fill_1 FILLER_74_1079 ();
 sg13g2_fill_2 FILLER_74_1109 ();
 sg13g2_decap_4 FILLER_74_1116 ();
 sg13g2_fill_1 FILLER_74_1120 ();
 sg13g2_decap_8 FILLER_74_1141 ();
 sg13g2_decap_8 FILLER_74_1148 ();
 sg13g2_decap_8 FILLER_74_1155 ();
 sg13g2_decap_8 FILLER_74_1162 ();
 sg13g2_decap_8 FILLER_74_1169 ();
 sg13g2_decap_8 FILLER_74_1176 ();
 sg13g2_decap_8 FILLER_74_1183 ();
 sg13g2_decap_8 FILLER_74_1190 ();
 sg13g2_decap_8 FILLER_74_1197 ();
 sg13g2_decap_8 FILLER_74_1204 ();
 sg13g2_decap_8 FILLER_74_1211 ();
 sg13g2_decap_8 FILLER_74_1218 ();
 sg13g2_decap_8 FILLER_74_1225 ();
 sg13g2_decap_8 FILLER_74_1232 ();
 sg13g2_decap_8 FILLER_74_1239 ();
 sg13g2_decap_8 FILLER_74_1246 ();
 sg13g2_decap_8 FILLER_74_1253 ();
 sg13g2_decap_8 FILLER_74_1260 ();
 sg13g2_decap_8 FILLER_74_1267 ();
 sg13g2_decap_8 FILLER_74_1274 ();
 sg13g2_decap_8 FILLER_74_1281 ();
 sg13g2_decap_8 FILLER_74_1288 ();
 sg13g2_decap_8 FILLER_74_1295 ();
 sg13g2_decap_8 FILLER_74_1302 ();
 sg13g2_decap_8 FILLER_74_1309 ();
 sg13g2_decap_8 FILLER_74_1316 ();
 sg13g2_decap_8 FILLER_74_1323 ();
 sg13g2_decap_8 FILLER_74_1330 ();
 sg13g2_decap_8 FILLER_74_1337 ();
 sg13g2_decap_8 FILLER_74_1344 ();
 sg13g2_decap_8 FILLER_74_1351 ();
 sg13g2_decap_8 FILLER_74_1358 ();
 sg13g2_decap_8 FILLER_74_1365 ();
 sg13g2_decap_8 FILLER_74_1372 ();
 sg13g2_decap_8 FILLER_74_1379 ();
 sg13g2_decap_8 FILLER_74_1386 ();
 sg13g2_decap_8 FILLER_74_1393 ();
 sg13g2_decap_8 FILLER_74_1400 ();
 sg13g2_decap_8 FILLER_74_1407 ();
 sg13g2_decap_8 FILLER_74_1414 ();
 sg13g2_decap_8 FILLER_74_1421 ();
 sg13g2_decap_8 FILLER_74_1428 ();
 sg13g2_decap_8 FILLER_74_1435 ();
 sg13g2_decap_8 FILLER_74_1442 ();
 sg13g2_decap_8 FILLER_74_1449 ();
 sg13g2_decap_8 FILLER_74_1456 ();
 sg13g2_decap_8 FILLER_74_1463 ();
 sg13g2_decap_8 FILLER_74_1470 ();
 sg13g2_decap_8 FILLER_74_1477 ();
 sg13g2_decap_8 FILLER_74_1484 ();
 sg13g2_decap_8 FILLER_74_1491 ();
 sg13g2_decap_8 FILLER_74_1498 ();
 sg13g2_decap_8 FILLER_74_1505 ();
 sg13g2_decap_8 FILLER_74_1512 ();
 sg13g2_decap_8 FILLER_74_1519 ();
 sg13g2_decap_8 FILLER_74_1526 ();
 sg13g2_decap_8 FILLER_74_1533 ();
 sg13g2_decap_8 FILLER_74_1540 ();
 sg13g2_decap_8 FILLER_74_1547 ();
 sg13g2_decap_8 FILLER_74_1554 ();
 sg13g2_decap_8 FILLER_74_1561 ();
 sg13g2_decap_8 FILLER_74_1568 ();
 sg13g2_decap_8 FILLER_74_1575 ();
 sg13g2_decap_8 FILLER_74_1582 ();
 sg13g2_decap_8 FILLER_74_1589 ();
 sg13g2_decap_8 FILLER_74_1596 ();
 sg13g2_decap_8 FILLER_74_1603 ();
 sg13g2_decap_8 FILLER_74_1610 ();
 sg13g2_decap_8 FILLER_74_1617 ();
 sg13g2_decap_8 FILLER_74_1624 ();
 sg13g2_decap_8 FILLER_74_1631 ();
 sg13g2_decap_8 FILLER_74_1638 ();
 sg13g2_decap_8 FILLER_74_1645 ();
 sg13g2_decap_8 FILLER_74_1652 ();
 sg13g2_decap_8 FILLER_74_1659 ();
 sg13g2_decap_8 FILLER_74_1666 ();
 sg13g2_decap_8 FILLER_74_1673 ();
 sg13g2_decap_8 FILLER_74_1680 ();
 sg13g2_decap_8 FILLER_74_1687 ();
 sg13g2_decap_8 FILLER_74_1694 ();
 sg13g2_decap_8 FILLER_74_1701 ();
 sg13g2_decap_8 FILLER_74_1708 ();
 sg13g2_decap_8 FILLER_74_1715 ();
 sg13g2_decap_8 FILLER_74_1722 ();
 sg13g2_decap_8 FILLER_74_1729 ();
 sg13g2_decap_8 FILLER_74_1736 ();
 sg13g2_decap_8 FILLER_74_1743 ();
 sg13g2_decap_8 FILLER_74_1750 ();
 sg13g2_decap_8 FILLER_74_1757 ();
 sg13g2_decap_4 FILLER_74_1764 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_26 ();
 sg13g2_fill_2 FILLER_75_45 ();
 sg13g2_fill_2 FILLER_75_61 ();
 sg13g2_fill_1 FILLER_75_77 ();
 sg13g2_fill_1 FILLER_75_111 ();
 sg13g2_fill_1 FILLER_75_138 ();
 sg13g2_fill_2 FILLER_75_155 ();
 sg13g2_fill_1 FILLER_75_185 ();
 sg13g2_fill_2 FILLER_75_191 ();
 sg13g2_fill_2 FILLER_75_246 ();
 sg13g2_fill_2 FILLER_75_305 ();
 sg13g2_fill_2 FILLER_75_315 ();
 sg13g2_fill_2 FILLER_75_321 ();
 sg13g2_fill_1 FILLER_75_378 ();
 sg13g2_fill_2 FILLER_75_393 ();
 sg13g2_fill_2 FILLER_75_455 ();
 sg13g2_fill_2 FILLER_75_488 ();
 sg13g2_fill_1 FILLER_75_490 ();
 sg13g2_fill_2 FILLER_75_524 ();
 sg13g2_fill_1 FILLER_75_526 ();
 sg13g2_fill_2 FILLER_75_550 ();
 sg13g2_fill_2 FILLER_75_592 ();
 sg13g2_fill_1 FILLER_75_641 ();
 sg13g2_decap_4 FILLER_75_667 ();
 sg13g2_fill_1 FILLER_75_671 ();
 sg13g2_fill_2 FILLER_75_706 ();
 sg13g2_fill_1 FILLER_75_728 ();
 sg13g2_fill_1 FILLER_75_754 ();
 sg13g2_decap_8 FILLER_75_763 ();
 sg13g2_decap_8 FILLER_75_770 ();
 sg13g2_fill_2 FILLER_75_777 ();
 sg13g2_fill_2 FILLER_75_792 ();
 sg13g2_fill_1 FILLER_75_794 ();
 sg13g2_fill_2 FILLER_75_824 ();
 sg13g2_decap_4 FILLER_75_846 ();
 sg13g2_fill_2 FILLER_75_850 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_75_868 ();
 sg13g2_fill_2 FILLER_75_875 ();
 sg13g2_fill_1 FILLER_75_877 ();
 sg13g2_fill_2 FILLER_75_883 ();
 sg13g2_fill_1 FILLER_75_885 ();
 sg13g2_fill_1 FILLER_75_903 ();
 sg13g2_fill_1 FILLER_75_998 ();
 sg13g2_fill_2 FILLER_75_1070 ();
 sg13g2_fill_1 FILLER_75_1072 ();
 sg13g2_fill_2 FILLER_75_1089 ();
 sg13g2_fill_2 FILLER_75_1095 ();
 sg13g2_fill_1 FILLER_75_1097 ();
 sg13g2_decap_8 FILLER_75_1110 ();
 sg13g2_decap_8 FILLER_75_1117 ();
 sg13g2_decap_8 FILLER_75_1124 ();
 sg13g2_decap_8 FILLER_75_1131 ();
 sg13g2_decap_8 FILLER_75_1138 ();
 sg13g2_decap_8 FILLER_75_1145 ();
 sg13g2_decap_8 FILLER_75_1152 ();
 sg13g2_decap_8 FILLER_75_1159 ();
 sg13g2_decap_8 FILLER_75_1166 ();
 sg13g2_decap_8 FILLER_75_1173 ();
 sg13g2_decap_8 FILLER_75_1180 ();
 sg13g2_decap_8 FILLER_75_1187 ();
 sg13g2_decap_8 FILLER_75_1194 ();
 sg13g2_decap_8 FILLER_75_1201 ();
 sg13g2_decap_8 FILLER_75_1208 ();
 sg13g2_decap_8 FILLER_75_1215 ();
 sg13g2_decap_8 FILLER_75_1222 ();
 sg13g2_decap_8 FILLER_75_1229 ();
 sg13g2_decap_8 FILLER_75_1236 ();
 sg13g2_decap_8 FILLER_75_1243 ();
 sg13g2_decap_8 FILLER_75_1250 ();
 sg13g2_decap_8 FILLER_75_1257 ();
 sg13g2_decap_8 FILLER_75_1264 ();
 sg13g2_decap_8 FILLER_75_1271 ();
 sg13g2_decap_8 FILLER_75_1278 ();
 sg13g2_decap_8 FILLER_75_1285 ();
 sg13g2_decap_8 FILLER_75_1292 ();
 sg13g2_decap_8 FILLER_75_1299 ();
 sg13g2_decap_8 FILLER_75_1306 ();
 sg13g2_decap_8 FILLER_75_1313 ();
 sg13g2_decap_8 FILLER_75_1320 ();
 sg13g2_decap_8 FILLER_75_1327 ();
 sg13g2_decap_8 FILLER_75_1334 ();
 sg13g2_decap_8 FILLER_75_1341 ();
 sg13g2_decap_8 FILLER_75_1348 ();
 sg13g2_decap_8 FILLER_75_1355 ();
 sg13g2_decap_8 FILLER_75_1362 ();
 sg13g2_decap_8 FILLER_75_1369 ();
 sg13g2_decap_8 FILLER_75_1376 ();
 sg13g2_decap_8 FILLER_75_1383 ();
 sg13g2_decap_8 FILLER_75_1390 ();
 sg13g2_decap_8 FILLER_75_1397 ();
 sg13g2_decap_8 FILLER_75_1404 ();
 sg13g2_decap_8 FILLER_75_1411 ();
 sg13g2_decap_8 FILLER_75_1418 ();
 sg13g2_decap_8 FILLER_75_1425 ();
 sg13g2_decap_8 FILLER_75_1432 ();
 sg13g2_decap_8 FILLER_75_1439 ();
 sg13g2_decap_8 FILLER_75_1446 ();
 sg13g2_decap_8 FILLER_75_1453 ();
 sg13g2_decap_8 FILLER_75_1460 ();
 sg13g2_decap_8 FILLER_75_1467 ();
 sg13g2_decap_8 FILLER_75_1474 ();
 sg13g2_decap_8 FILLER_75_1481 ();
 sg13g2_decap_8 FILLER_75_1488 ();
 sg13g2_decap_8 FILLER_75_1495 ();
 sg13g2_decap_8 FILLER_75_1502 ();
 sg13g2_decap_8 FILLER_75_1509 ();
 sg13g2_decap_8 FILLER_75_1516 ();
 sg13g2_decap_8 FILLER_75_1523 ();
 sg13g2_decap_8 FILLER_75_1530 ();
 sg13g2_decap_8 FILLER_75_1537 ();
 sg13g2_decap_8 FILLER_75_1544 ();
 sg13g2_decap_8 FILLER_75_1551 ();
 sg13g2_decap_8 FILLER_75_1558 ();
 sg13g2_decap_8 FILLER_75_1565 ();
 sg13g2_decap_8 FILLER_75_1572 ();
 sg13g2_decap_8 FILLER_75_1579 ();
 sg13g2_decap_8 FILLER_75_1586 ();
 sg13g2_decap_8 FILLER_75_1593 ();
 sg13g2_decap_8 FILLER_75_1600 ();
 sg13g2_decap_8 FILLER_75_1607 ();
 sg13g2_decap_8 FILLER_75_1614 ();
 sg13g2_decap_8 FILLER_75_1621 ();
 sg13g2_decap_8 FILLER_75_1628 ();
 sg13g2_decap_8 FILLER_75_1635 ();
 sg13g2_decap_8 FILLER_75_1642 ();
 sg13g2_decap_8 FILLER_75_1649 ();
 sg13g2_decap_8 FILLER_75_1656 ();
 sg13g2_decap_8 FILLER_75_1663 ();
 sg13g2_decap_8 FILLER_75_1670 ();
 sg13g2_decap_8 FILLER_75_1677 ();
 sg13g2_decap_8 FILLER_75_1684 ();
 sg13g2_decap_8 FILLER_75_1691 ();
 sg13g2_decap_8 FILLER_75_1698 ();
 sg13g2_decap_8 FILLER_75_1705 ();
 sg13g2_decap_8 FILLER_75_1712 ();
 sg13g2_decap_8 FILLER_75_1719 ();
 sg13g2_decap_8 FILLER_75_1726 ();
 sg13g2_decap_8 FILLER_75_1733 ();
 sg13g2_decap_8 FILLER_75_1740 ();
 sg13g2_decap_8 FILLER_75_1747 ();
 sg13g2_decap_8 FILLER_75_1754 ();
 sg13g2_decap_8 FILLER_75_1761 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_37 ();
 sg13g2_fill_1 FILLER_76_48 ();
 sg13g2_fill_1 FILLER_76_101 ();
 sg13g2_fill_1 FILLER_76_146 ();
 sg13g2_fill_2 FILLER_76_184 ();
 sg13g2_fill_1 FILLER_76_209 ();
 sg13g2_fill_2 FILLER_76_339 ();
 sg13g2_fill_1 FILLER_76_421 ();
 sg13g2_fill_1 FILLER_76_437 ();
 sg13g2_decap_8 FILLER_76_458 ();
 sg13g2_decap_4 FILLER_76_465 ();
 sg13g2_fill_1 FILLER_76_469 ();
 sg13g2_decap_8 FILLER_76_477 ();
 sg13g2_fill_2 FILLER_76_484 ();
 sg13g2_fill_1 FILLER_76_486 ();
 sg13g2_fill_1 FILLER_76_500 ();
 sg13g2_decap_4 FILLER_76_531 ();
 sg13g2_fill_1 FILLER_76_545 ();
 sg13g2_fill_2 FILLER_76_551 ();
 sg13g2_fill_1 FILLER_76_553 ();
 sg13g2_fill_2 FILLER_76_600 ();
 sg13g2_decap_8 FILLER_76_623 ();
 sg13g2_decap_4 FILLER_76_630 ();
 sg13g2_fill_1 FILLER_76_654 ();
 sg13g2_fill_2 FILLER_76_674 ();
 sg13g2_fill_1 FILLER_76_676 ();
 sg13g2_fill_2 FILLER_76_691 ();
 sg13g2_fill_1 FILLER_76_693 ();
 sg13g2_decap_4 FILLER_76_714 ();
 sg13g2_fill_1 FILLER_76_718 ();
 sg13g2_fill_1 FILLER_76_727 ();
 sg13g2_fill_2 FILLER_76_736 ();
 sg13g2_fill_1 FILLER_76_742 ();
 sg13g2_fill_1 FILLER_76_751 ();
 sg13g2_decap_4 FILLER_76_756 ();
 sg13g2_fill_1 FILLER_76_760 ();
 sg13g2_fill_1 FILLER_76_772 ();
 sg13g2_decap_8 FILLER_76_794 ();
 sg13g2_fill_1 FILLER_76_801 ();
 sg13g2_fill_2 FILLER_76_822 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_fill_2 FILLER_76_856 ();
 sg13g2_fill_1 FILLER_76_884 ();
 sg13g2_fill_1 FILLER_76_906 ();
 sg13g2_fill_1 FILLER_76_937 ();
 sg13g2_fill_1 FILLER_76_969 ();
 sg13g2_fill_1 FILLER_76_1020 ();
 sg13g2_decap_8 FILLER_76_1079 ();
 sg13g2_decap_8 FILLER_76_1086 ();
 sg13g2_decap_8 FILLER_76_1093 ();
 sg13g2_decap_8 FILLER_76_1100 ();
 sg13g2_decap_8 FILLER_76_1107 ();
 sg13g2_decap_8 FILLER_76_1114 ();
 sg13g2_decap_8 FILLER_76_1121 ();
 sg13g2_decap_8 FILLER_76_1128 ();
 sg13g2_decap_8 FILLER_76_1135 ();
 sg13g2_decap_8 FILLER_76_1142 ();
 sg13g2_decap_8 FILLER_76_1149 ();
 sg13g2_decap_8 FILLER_76_1156 ();
 sg13g2_decap_8 FILLER_76_1163 ();
 sg13g2_decap_8 FILLER_76_1170 ();
 sg13g2_decap_8 FILLER_76_1177 ();
 sg13g2_decap_8 FILLER_76_1184 ();
 sg13g2_decap_8 FILLER_76_1191 ();
 sg13g2_decap_8 FILLER_76_1198 ();
 sg13g2_decap_8 FILLER_76_1205 ();
 sg13g2_decap_8 FILLER_76_1212 ();
 sg13g2_decap_8 FILLER_76_1219 ();
 sg13g2_decap_8 FILLER_76_1226 ();
 sg13g2_decap_8 FILLER_76_1233 ();
 sg13g2_decap_8 FILLER_76_1240 ();
 sg13g2_decap_8 FILLER_76_1247 ();
 sg13g2_decap_8 FILLER_76_1254 ();
 sg13g2_decap_8 FILLER_76_1261 ();
 sg13g2_decap_8 FILLER_76_1268 ();
 sg13g2_decap_8 FILLER_76_1275 ();
 sg13g2_decap_8 FILLER_76_1282 ();
 sg13g2_decap_8 FILLER_76_1289 ();
 sg13g2_decap_8 FILLER_76_1296 ();
 sg13g2_decap_8 FILLER_76_1303 ();
 sg13g2_decap_8 FILLER_76_1310 ();
 sg13g2_decap_8 FILLER_76_1317 ();
 sg13g2_decap_8 FILLER_76_1324 ();
 sg13g2_decap_8 FILLER_76_1331 ();
 sg13g2_decap_8 FILLER_76_1338 ();
 sg13g2_decap_8 FILLER_76_1345 ();
 sg13g2_decap_8 FILLER_76_1352 ();
 sg13g2_decap_8 FILLER_76_1359 ();
 sg13g2_decap_8 FILLER_76_1366 ();
 sg13g2_decap_8 FILLER_76_1373 ();
 sg13g2_decap_8 FILLER_76_1380 ();
 sg13g2_decap_8 FILLER_76_1387 ();
 sg13g2_decap_8 FILLER_76_1394 ();
 sg13g2_decap_8 FILLER_76_1401 ();
 sg13g2_decap_8 FILLER_76_1408 ();
 sg13g2_decap_8 FILLER_76_1415 ();
 sg13g2_decap_8 FILLER_76_1422 ();
 sg13g2_decap_8 FILLER_76_1429 ();
 sg13g2_decap_8 FILLER_76_1436 ();
 sg13g2_decap_8 FILLER_76_1443 ();
 sg13g2_decap_8 FILLER_76_1450 ();
 sg13g2_decap_8 FILLER_76_1457 ();
 sg13g2_decap_8 FILLER_76_1464 ();
 sg13g2_decap_8 FILLER_76_1471 ();
 sg13g2_decap_8 FILLER_76_1478 ();
 sg13g2_decap_8 FILLER_76_1485 ();
 sg13g2_decap_8 FILLER_76_1492 ();
 sg13g2_decap_8 FILLER_76_1499 ();
 sg13g2_decap_8 FILLER_76_1506 ();
 sg13g2_decap_8 FILLER_76_1513 ();
 sg13g2_decap_8 FILLER_76_1520 ();
 sg13g2_decap_8 FILLER_76_1527 ();
 sg13g2_decap_8 FILLER_76_1534 ();
 sg13g2_decap_8 FILLER_76_1541 ();
 sg13g2_decap_8 FILLER_76_1548 ();
 sg13g2_decap_8 FILLER_76_1555 ();
 sg13g2_decap_8 FILLER_76_1562 ();
 sg13g2_decap_8 FILLER_76_1569 ();
 sg13g2_decap_8 FILLER_76_1576 ();
 sg13g2_decap_8 FILLER_76_1583 ();
 sg13g2_decap_8 FILLER_76_1590 ();
 sg13g2_decap_8 FILLER_76_1597 ();
 sg13g2_decap_8 FILLER_76_1604 ();
 sg13g2_decap_8 FILLER_76_1611 ();
 sg13g2_decap_8 FILLER_76_1618 ();
 sg13g2_decap_8 FILLER_76_1625 ();
 sg13g2_decap_8 FILLER_76_1632 ();
 sg13g2_decap_8 FILLER_76_1639 ();
 sg13g2_decap_8 FILLER_76_1646 ();
 sg13g2_decap_8 FILLER_76_1653 ();
 sg13g2_decap_8 FILLER_76_1660 ();
 sg13g2_decap_8 FILLER_76_1667 ();
 sg13g2_decap_8 FILLER_76_1674 ();
 sg13g2_decap_8 FILLER_76_1681 ();
 sg13g2_decap_8 FILLER_76_1688 ();
 sg13g2_decap_8 FILLER_76_1695 ();
 sg13g2_decap_8 FILLER_76_1702 ();
 sg13g2_decap_8 FILLER_76_1709 ();
 sg13g2_decap_8 FILLER_76_1716 ();
 sg13g2_decap_8 FILLER_76_1723 ();
 sg13g2_decap_8 FILLER_76_1730 ();
 sg13g2_decap_8 FILLER_76_1737 ();
 sg13g2_decap_8 FILLER_76_1744 ();
 sg13g2_decap_8 FILLER_76_1751 ();
 sg13g2_decap_8 FILLER_76_1758 ();
 sg13g2_fill_2 FILLER_76_1765 ();
 sg13g2_fill_1 FILLER_76_1767 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_31 ();
 sg13g2_fill_1 FILLER_77_56 ();
 sg13g2_fill_2 FILLER_77_106 ();
 sg13g2_fill_2 FILLER_77_130 ();
 sg13g2_fill_2 FILLER_77_139 ();
 sg13g2_fill_1 FILLER_77_146 ();
 sg13g2_fill_2 FILLER_77_233 ();
 sg13g2_fill_1 FILLER_77_261 ();
 sg13g2_fill_1 FILLER_77_315 ();
 sg13g2_fill_1 FILLER_77_324 ();
 sg13g2_fill_2 FILLER_77_351 ();
 sg13g2_fill_1 FILLER_77_365 ();
 sg13g2_fill_2 FILLER_77_397 ();
 sg13g2_fill_1 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_424 ();
 sg13g2_fill_2 FILLER_77_439 ();
 sg13g2_fill_1 FILLER_77_441 ();
 sg13g2_decap_8 FILLER_77_452 ();
 sg13g2_fill_1 FILLER_77_459 ();
 sg13g2_decap_4 FILLER_77_487 ();
 sg13g2_fill_1 FILLER_77_491 ();
 sg13g2_decap_8 FILLER_77_550 ();
 sg13g2_decap_8 FILLER_77_557 ();
 sg13g2_decap_8 FILLER_77_564 ();
 sg13g2_decap_8 FILLER_77_575 ();
 sg13g2_fill_1 FILLER_77_582 ();
 sg13g2_decap_4 FILLER_77_587 ();
 sg13g2_fill_1 FILLER_77_591 ();
 sg13g2_decap_8 FILLER_77_597 ();
 sg13g2_fill_1 FILLER_77_604 ();
 sg13g2_decap_8 FILLER_77_613 ();
 sg13g2_fill_2 FILLER_77_649 ();
 sg13g2_fill_1 FILLER_77_651 ();
 sg13g2_decap_8 FILLER_77_674 ();
 sg13g2_decap_4 FILLER_77_681 ();
 sg13g2_decap_4 FILLER_77_691 ();
 sg13g2_fill_1 FILLER_77_695 ();
 sg13g2_fill_2 FILLER_77_710 ();
 sg13g2_fill_1 FILLER_77_712 ();
 sg13g2_fill_2 FILLER_77_749 ();
 sg13g2_fill_1 FILLER_77_751 ();
 sg13g2_fill_2 FILLER_77_773 ();
 sg13g2_fill_1 FILLER_77_775 ();
 sg13g2_fill_2 FILLER_77_802 ();
 sg13g2_decap_8 FILLER_77_847 ();
 sg13g2_fill_2 FILLER_77_854 ();
 sg13g2_fill_2 FILLER_77_925 ();
 sg13g2_fill_1 FILLER_77_927 ();
 sg13g2_fill_2 FILLER_77_949 ();
 sg13g2_fill_2 FILLER_77_1053 ();
 sg13g2_decap_8 FILLER_77_1074 ();
 sg13g2_decap_8 FILLER_77_1081 ();
 sg13g2_decap_8 FILLER_77_1088 ();
 sg13g2_decap_8 FILLER_77_1095 ();
 sg13g2_decap_8 FILLER_77_1102 ();
 sg13g2_decap_8 FILLER_77_1109 ();
 sg13g2_decap_8 FILLER_77_1116 ();
 sg13g2_decap_8 FILLER_77_1123 ();
 sg13g2_decap_8 FILLER_77_1130 ();
 sg13g2_decap_8 FILLER_77_1137 ();
 sg13g2_decap_8 FILLER_77_1144 ();
 sg13g2_decap_8 FILLER_77_1151 ();
 sg13g2_decap_8 FILLER_77_1158 ();
 sg13g2_decap_8 FILLER_77_1165 ();
 sg13g2_decap_8 FILLER_77_1172 ();
 sg13g2_decap_8 FILLER_77_1179 ();
 sg13g2_decap_8 FILLER_77_1186 ();
 sg13g2_decap_8 FILLER_77_1193 ();
 sg13g2_decap_8 FILLER_77_1200 ();
 sg13g2_decap_8 FILLER_77_1207 ();
 sg13g2_decap_8 FILLER_77_1214 ();
 sg13g2_decap_8 FILLER_77_1221 ();
 sg13g2_decap_8 FILLER_77_1228 ();
 sg13g2_decap_8 FILLER_77_1235 ();
 sg13g2_decap_8 FILLER_77_1242 ();
 sg13g2_decap_8 FILLER_77_1249 ();
 sg13g2_decap_8 FILLER_77_1256 ();
 sg13g2_decap_8 FILLER_77_1263 ();
 sg13g2_decap_8 FILLER_77_1270 ();
 sg13g2_decap_8 FILLER_77_1277 ();
 sg13g2_decap_8 FILLER_77_1284 ();
 sg13g2_decap_8 FILLER_77_1291 ();
 sg13g2_decap_8 FILLER_77_1298 ();
 sg13g2_decap_8 FILLER_77_1305 ();
 sg13g2_decap_8 FILLER_77_1312 ();
 sg13g2_decap_8 FILLER_77_1319 ();
 sg13g2_decap_8 FILLER_77_1326 ();
 sg13g2_decap_8 FILLER_77_1333 ();
 sg13g2_decap_8 FILLER_77_1340 ();
 sg13g2_decap_8 FILLER_77_1347 ();
 sg13g2_decap_8 FILLER_77_1354 ();
 sg13g2_decap_8 FILLER_77_1361 ();
 sg13g2_decap_8 FILLER_77_1368 ();
 sg13g2_decap_8 FILLER_77_1375 ();
 sg13g2_decap_8 FILLER_77_1382 ();
 sg13g2_decap_8 FILLER_77_1389 ();
 sg13g2_decap_8 FILLER_77_1396 ();
 sg13g2_decap_8 FILLER_77_1403 ();
 sg13g2_decap_8 FILLER_77_1410 ();
 sg13g2_decap_8 FILLER_77_1417 ();
 sg13g2_decap_8 FILLER_77_1424 ();
 sg13g2_decap_8 FILLER_77_1431 ();
 sg13g2_decap_8 FILLER_77_1438 ();
 sg13g2_decap_8 FILLER_77_1445 ();
 sg13g2_decap_8 FILLER_77_1452 ();
 sg13g2_decap_8 FILLER_77_1459 ();
 sg13g2_decap_8 FILLER_77_1466 ();
 sg13g2_decap_8 FILLER_77_1473 ();
 sg13g2_decap_8 FILLER_77_1480 ();
 sg13g2_decap_8 FILLER_77_1487 ();
 sg13g2_decap_8 FILLER_77_1494 ();
 sg13g2_decap_8 FILLER_77_1501 ();
 sg13g2_decap_8 FILLER_77_1508 ();
 sg13g2_decap_8 FILLER_77_1515 ();
 sg13g2_decap_8 FILLER_77_1522 ();
 sg13g2_decap_8 FILLER_77_1529 ();
 sg13g2_decap_8 FILLER_77_1536 ();
 sg13g2_decap_8 FILLER_77_1543 ();
 sg13g2_decap_8 FILLER_77_1550 ();
 sg13g2_decap_8 FILLER_77_1557 ();
 sg13g2_decap_8 FILLER_77_1564 ();
 sg13g2_decap_8 FILLER_77_1571 ();
 sg13g2_decap_8 FILLER_77_1578 ();
 sg13g2_decap_8 FILLER_77_1585 ();
 sg13g2_decap_8 FILLER_77_1592 ();
 sg13g2_decap_8 FILLER_77_1599 ();
 sg13g2_decap_8 FILLER_77_1606 ();
 sg13g2_decap_8 FILLER_77_1613 ();
 sg13g2_decap_8 FILLER_77_1620 ();
 sg13g2_decap_8 FILLER_77_1627 ();
 sg13g2_decap_8 FILLER_77_1634 ();
 sg13g2_decap_8 FILLER_77_1641 ();
 sg13g2_decap_8 FILLER_77_1648 ();
 sg13g2_decap_8 FILLER_77_1655 ();
 sg13g2_decap_8 FILLER_77_1662 ();
 sg13g2_decap_8 FILLER_77_1669 ();
 sg13g2_decap_8 FILLER_77_1676 ();
 sg13g2_decap_8 FILLER_77_1683 ();
 sg13g2_decap_8 FILLER_77_1690 ();
 sg13g2_decap_8 FILLER_77_1697 ();
 sg13g2_decap_8 FILLER_77_1704 ();
 sg13g2_decap_8 FILLER_77_1711 ();
 sg13g2_decap_8 FILLER_77_1718 ();
 sg13g2_decap_8 FILLER_77_1725 ();
 sg13g2_decap_8 FILLER_77_1732 ();
 sg13g2_decap_8 FILLER_77_1739 ();
 sg13g2_decap_8 FILLER_77_1746 ();
 sg13g2_decap_8 FILLER_77_1753 ();
 sg13g2_decap_8 FILLER_77_1760 ();
 sg13g2_fill_1 FILLER_77_1767 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_66 ();
 sg13g2_fill_1 FILLER_78_83 ();
 sg13g2_fill_2 FILLER_78_119 ();
 sg13g2_fill_2 FILLER_78_173 ();
 sg13g2_fill_1 FILLER_78_182 ();
 sg13g2_fill_1 FILLER_78_227 ();
 sg13g2_fill_1 FILLER_78_267 ();
 sg13g2_fill_2 FILLER_78_281 ();
 sg13g2_fill_2 FILLER_78_293 ();
 sg13g2_fill_1 FILLER_78_336 ();
 sg13g2_fill_2 FILLER_78_346 ();
 sg13g2_fill_2 FILLER_78_404 ();
 sg13g2_fill_2 FILLER_78_411 ();
 sg13g2_fill_2 FILLER_78_433 ();
 sg13g2_fill_1 FILLER_78_435 ();
 sg13g2_fill_2 FILLER_78_441 ();
 sg13g2_fill_1 FILLER_78_443 ();
 sg13g2_decap_4 FILLER_78_454 ();
 sg13g2_fill_2 FILLER_78_458 ();
 sg13g2_fill_1 FILLER_78_470 ();
 sg13g2_decap_4 FILLER_78_479 ();
 sg13g2_fill_2 FILLER_78_483 ();
 sg13g2_fill_2 FILLER_78_493 ();
 sg13g2_fill_1 FILLER_78_495 ();
 sg13g2_fill_2 FILLER_78_507 ();
 sg13g2_fill_2 FILLER_78_513 ();
 sg13g2_fill_1 FILLER_78_524 ();
 sg13g2_fill_2 FILLER_78_537 ();
 sg13g2_fill_1 FILLER_78_539 ();
 sg13g2_fill_1 FILLER_78_563 ();
 sg13g2_fill_1 FILLER_78_583 ();
 sg13g2_fill_1 FILLER_78_597 ();
 sg13g2_fill_2 FILLER_78_609 ();
 sg13g2_decap_8 FILLER_78_646 ();
 sg13g2_fill_1 FILLER_78_653 ();
 sg13g2_decap_4 FILLER_78_670 ();
 sg13g2_decap_8 FILLER_78_694 ();
 sg13g2_fill_1 FILLER_78_708 ();
 sg13g2_fill_1 FILLER_78_720 ();
 sg13g2_fill_2 FILLER_78_729 ();
 sg13g2_fill_1 FILLER_78_741 ();
 sg13g2_decap_8 FILLER_78_751 ();
 sg13g2_fill_2 FILLER_78_758 ();
 sg13g2_fill_1 FILLER_78_787 ();
 sg13g2_decap_4 FILLER_78_796 ();
 sg13g2_fill_1 FILLER_78_800 ();
 sg13g2_decap_8 FILLER_78_821 ();
 sg13g2_fill_2 FILLER_78_828 ();
 sg13g2_decap_8 FILLER_78_855 ();
 sg13g2_fill_1 FILLER_78_862 ();
 sg13g2_decap_8 FILLER_78_866 ();
 sg13g2_decap_4 FILLER_78_873 ();
 sg13g2_fill_2 FILLER_78_877 ();
 sg13g2_decap_8 FILLER_78_915 ();
 sg13g2_decap_4 FILLER_78_922 ();
 sg13g2_fill_1 FILLER_78_976 ();
 sg13g2_fill_2 FILLER_78_981 ();
 sg13g2_fill_2 FILLER_78_1023 ();
 sg13g2_decap_8 FILLER_78_1068 ();
 sg13g2_decap_8 FILLER_78_1075 ();
 sg13g2_decap_8 FILLER_78_1082 ();
 sg13g2_decap_8 FILLER_78_1089 ();
 sg13g2_decap_8 FILLER_78_1096 ();
 sg13g2_decap_8 FILLER_78_1103 ();
 sg13g2_decap_8 FILLER_78_1110 ();
 sg13g2_decap_8 FILLER_78_1117 ();
 sg13g2_decap_8 FILLER_78_1124 ();
 sg13g2_decap_8 FILLER_78_1131 ();
 sg13g2_decap_8 FILLER_78_1138 ();
 sg13g2_decap_8 FILLER_78_1145 ();
 sg13g2_decap_8 FILLER_78_1152 ();
 sg13g2_decap_8 FILLER_78_1159 ();
 sg13g2_decap_8 FILLER_78_1166 ();
 sg13g2_decap_8 FILLER_78_1173 ();
 sg13g2_decap_8 FILLER_78_1180 ();
 sg13g2_decap_8 FILLER_78_1187 ();
 sg13g2_decap_8 FILLER_78_1194 ();
 sg13g2_decap_8 FILLER_78_1201 ();
 sg13g2_decap_8 FILLER_78_1208 ();
 sg13g2_decap_8 FILLER_78_1215 ();
 sg13g2_decap_8 FILLER_78_1222 ();
 sg13g2_decap_8 FILLER_78_1229 ();
 sg13g2_decap_8 FILLER_78_1236 ();
 sg13g2_decap_8 FILLER_78_1243 ();
 sg13g2_decap_8 FILLER_78_1250 ();
 sg13g2_decap_8 FILLER_78_1257 ();
 sg13g2_decap_8 FILLER_78_1264 ();
 sg13g2_decap_8 FILLER_78_1271 ();
 sg13g2_decap_8 FILLER_78_1278 ();
 sg13g2_decap_8 FILLER_78_1285 ();
 sg13g2_decap_8 FILLER_78_1292 ();
 sg13g2_decap_8 FILLER_78_1299 ();
 sg13g2_decap_8 FILLER_78_1306 ();
 sg13g2_decap_8 FILLER_78_1313 ();
 sg13g2_decap_8 FILLER_78_1320 ();
 sg13g2_decap_8 FILLER_78_1327 ();
 sg13g2_decap_8 FILLER_78_1334 ();
 sg13g2_decap_8 FILLER_78_1341 ();
 sg13g2_decap_8 FILLER_78_1348 ();
 sg13g2_decap_8 FILLER_78_1355 ();
 sg13g2_decap_8 FILLER_78_1362 ();
 sg13g2_decap_8 FILLER_78_1369 ();
 sg13g2_decap_8 FILLER_78_1376 ();
 sg13g2_decap_8 FILLER_78_1383 ();
 sg13g2_decap_8 FILLER_78_1390 ();
 sg13g2_decap_8 FILLER_78_1397 ();
 sg13g2_decap_8 FILLER_78_1404 ();
 sg13g2_decap_8 FILLER_78_1411 ();
 sg13g2_decap_8 FILLER_78_1418 ();
 sg13g2_decap_8 FILLER_78_1425 ();
 sg13g2_decap_8 FILLER_78_1432 ();
 sg13g2_decap_8 FILLER_78_1439 ();
 sg13g2_decap_8 FILLER_78_1446 ();
 sg13g2_decap_8 FILLER_78_1453 ();
 sg13g2_decap_8 FILLER_78_1460 ();
 sg13g2_decap_8 FILLER_78_1467 ();
 sg13g2_decap_8 FILLER_78_1474 ();
 sg13g2_decap_8 FILLER_78_1481 ();
 sg13g2_decap_8 FILLER_78_1488 ();
 sg13g2_decap_8 FILLER_78_1495 ();
 sg13g2_decap_8 FILLER_78_1502 ();
 sg13g2_decap_8 FILLER_78_1509 ();
 sg13g2_decap_8 FILLER_78_1516 ();
 sg13g2_decap_8 FILLER_78_1523 ();
 sg13g2_decap_8 FILLER_78_1530 ();
 sg13g2_decap_8 FILLER_78_1537 ();
 sg13g2_decap_8 FILLER_78_1544 ();
 sg13g2_decap_8 FILLER_78_1551 ();
 sg13g2_decap_8 FILLER_78_1558 ();
 sg13g2_decap_8 FILLER_78_1565 ();
 sg13g2_decap_8 FILLER_78_1572 ();
 sg13g2_decap_8 FILLER_78_1579 ();
 sg13g2_decap_8 FILLER_78_1586 ();
 sg13g2_decap_8 FILLER_78_1593 ();
 sg13g2_decap_8 FILLER_78_1600 ();
 sg13g2_decap_8 FILLER_78_1607 ();
 sg13g2_decap_8 FILLER_78_1614 ();
 sg13g2_decap_8 FILLER_78_1621 ();
 sg13g2_decap_8 FILLER_78_1628 ();
 sg13g2_decap_8 FILLER_78_1635 ();
 sg13g2_decap_8 FILLER_78_1642 ();
 sg13g2_decap_8 FILLER_78_1649 ();
 sg13g2_decap_8 FILLER_78_1656 ();
 sg13g2_decap_8 FILLER_78_1663 ();
 sg13g2_decap_8 FILLER_78_1670 ();
 sg13g2_decap_8 FILLER_78_1677 ();
 sg13g2_decap_8 FILLER_78_1684 ();
 sg13g2_decap_8 FILLER_78_1691 ();
 sg13g2_decap_8 FILLER_78_1698 ();
 sg13g2_decap_8 FILLER_78_1705 ();
 sg13g2_decap_8 FILLER_78_1712 ();
 sg13g2_decap_8 FILLER_78_1719 ();
 sg13g2_decap_8 FILLER_78_1726 ();
 sg13g2_decap_8 FILLER_78_1733 ();
 sg13g2_decap_8 FILLER_78_1740 ();
 sg13g2_decap_8 FILLER_78_1747 ();
 sg13g2_decap_8 FILLER_78_1754 ();
 sg13g2_decap_8 FILLER_78_1761 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_53 ();
 sg13g2_fill_1 FILLER_79_95 ();
 sg13g2_fill_2 FILLER_79_129 ();
 sg13g2_fill_2 FILLER_79_136 ();
 sg13g2_fill_1 FILLER_79_147 ();
 sg13g2_fill_1 FILLER_79_217 ();
 sg13g2_fill_2 FILLER_79_289 ();
 sg13g2_fill_1 FILLER_79_357 ();
 sg13g2_fill_2 FILLER_79_390 ();
 sg13g2_fill_2 FILLER_79_439 ();
 sg13g2_fill_1 FILLER_79_483 ();
 sg13g2_fill_1 FILLER_79_523 ();
 sg13g2_fill_1 FILLER_79_589 ();
 sg13g2_fill_2 FILLER_79_600 ();
 sg13g2_fill_1 FILLER_79_623 ();
 sg13g2_fill_2 FILLER_79_647 ();
 sg13g2_fill_1 FILLER_79_672 ();
 sg13g2_fill_2 FILLER_79_681 ();
 sg13g2_fill_2 FILLER_79_696 ();
 sg13g2_fill_1 FILLER_79_698 ();
 sg13g2_decap_8 FILLER_79_717 ();
 sg13g2_fill_2 FILLER_79_724 ();
 sg13g2_fill_1 FILLER_79_758 ();
 sg13g2_fill_1 FILLER_79_797 ();
 sg13g2_fill_2 FILLER_79_831 ();
 sg13g2_fill_1 FILLER_79_833 ();
 sg13g2_decap_8 FILLER_79_852 ();
 sg13g2_decap_4 FILLER_79_883 ();
 sg13g2_decap_4 FILLER_79_892 ();
 sg13g2_fill_1 FILLER_79_903 ();
 sg13g2_fill_2 FILLER_79_920 ();
 sg13g2_fill_1 FILLER_79_922 ();
 sg13g2_fill_1 FILLER_79_956 ();
 sg13g2_fill_1 FILLER_79_994 ();
 sg13g2_decap_8 FILLER_79_1064 ();
 sg13g2_decap_8 FILLER_79_1071 ();
 sg13g2_decap_8 FILLER_79_1078 ();
 sg13g2_decap_8 FILLER_79_1085 ();
 sg13g2_decap_8 FILLER_79_1092 ();
 sg13g2_decap_8 FILLER_79_1099 ();
 sg13g2_decap_8 FILLER_79_1106 ();
 sg13g2_decap_8 FILLER_79_1113 ();
 sg13g2_decap_8 FILLER_79_1120 ();
 sg13g2_decap_8 FILLER_79_1127 ();
 sg13g2_decap_8 FILLER_79_1134 ();
 sg13g2_decap_8 FILLER_79_1141 ();
 sg13g2_decap_8 FILLER_79_1148 ();
 sg13g2_decap_8 FILLER_79_1155 ();
 sg13g2_decap_8 FILLER_79_1162 ();
 sg13g2_decap_8 FILLER_79_1169 ();
 sg13g2_decap_8 FILLER_79_1176 ();
 sg13g2_decap_8 FILLER_79_1183 ();
 sg13g2_decap_8 FILLER_79_1190 ();
 sg13g2_decap_8 FILLER_79_1197 ();
 sg13g2_decap_8 FILLER_79_1204 ();
 sg13g2_decap_8 FILLER_79_1211 ();
 sg13g2_decap_8 FILLER_79_1218 ();
 sg13g2_decap_8 FILLER_79_1225 ();
 sg13g2_decap_8 FILLER_79_1232 ();
 sg13g2_decap_8 FILLER_79_1239 ();
 sg13g2_decap_8 FILLER_79_1246 ();
 sg13g2_decap_8 FILLER_79_1253 ();
 sg13g2_decap_8 FILLER_79_1260 ();
 sg13g2_decap_8 FILLER_79_1267 ();
 sg13g2_decap_8 FILLER_79_1274 ();
 sg13g2_decap_8 FILLER_79_1281 ();
 sg13g2_decap_8 FILLER_79_1288 ();
 sg13g2_decap_8 FILLER_79_1295 ();
 sg13g2_decap_8 FILLER_79_1302 ();
 sg13g2_decap_8 FILLER_79_1309 ();
 sg13g2_decap_8 FILLER_79_1316 ();
 sg13g2_decap_8 FILLER_79_1323 ();
 sg13g2_decap_8 FILLER_79_1330 ();
 sg13g2_decap_8 FILLER_79_1337 ();
 sg13g2_decap_8 FILLER_79_1344 ();
 sg13g2_decap_8 FILLER_79_1351 ();
 sg13g2_decap_8 FILLER_79_1358 ();
 sg13g2_decap_8 FILLER_79_1365 ();
 sg13g2_decap_8 FILLER_79_1372 ();
 sg13g2_decap_8 FILLER_79_1379 ();
 sg13g2_decap_8 FILLER_79_1386 ();
 sg13g2_decap_8 FILLER_79_1393 ();
 sg13g2_decap_8 FILLER_79_1400 ();
 sg13g2_decap_8 FILLER_79_1407 ();
 sg13g2_decap_8 FILLER_79_1414 ();
 sg13g2_decap_8 FILLER_79_1421 ();
 sg13g2_decap_8 FILLER_79_1428 ();
 sg13g2_decap_8 FILLER_79_1435 ();
 sg13g2_decap_8 FILLER_79_1442 ();
 sg13g2_decap_8 FILLER_79_1449 ();
 sg13g2_decap_8 FILLER_79_1456 ();
 sg13g2_decap_8 FILLER_79_1463 ();
 sg13g2_decap_8 FILLER_79_1470 ();
 sg13g2_decap_8 FILLER_79_1477 ();
 sg13g2_decap_8 FILLER_79_1484 ();
 sg13g2_decap_8 FILLER_79_1491 ();
 sg13g2_decap_8 FILLER_79_1498 ();
 sg13g2_decap_8 FILLER_79_1505 ();
 sg13g2_decap_8 FILLER_79_1512 ();
 sg13g2_decap_8 FILLER_79_1519 ();
 sg13g2_decap_8 FILLER_79_1526 ();
 sg13g2_decap_8 FILLER_79_1533 ();
 sg13g2_decap_8 FILLER_79_1540 ();
 sg13g2_decap_8 FILLER_79_1547 ();
 sg13g2_decap_8 FILLER_79_1554 ();
 sg13g2_decap_8 FILLER_79_1561 ();
 sg13g2_decap_8 FILLER_79_1568 ();
 sg13g2_decap_8 FILLER_79_1575 ();
 sg13g2_decap_8 FILLER_79_1582 ();
 sg13g2_decap_8 FILLER_79_1589 ();
 sg13g2_decap_8 FILLER_79_1596 ();
 sg13g2_decap_8 FILLER_79_1603 ();
 sg13g2_decap_8 FILLER_79_1610 ();
 sg13g2_decap_8 FILLER_79_1617 ();
 sg13g2_decap_8 FILLER_79_1624 ();
 sg13g2_decap_8 FILLER_79_1631 ();
 sg13g2_decap_8 FILLER_79_1638 ();
 sg13g2_decap_8 FILLER_79_1645 ();
 sg13g2_decap_8 FILLER_79_1652 ();
 sg13g2_decap_8 FILLER_79_1659 ();
 sg13g2_decap_8 FILLER_79_1666 ();
 sg13g2_decap_8 FILLER_79_1673 ();
 sg13g2_decap_8 FILLER_79_1680 ();
 sg13g2_decap_8 FILLER_79_1687 ();
 sg13g2_decap_8 FILLER_79_1694 ();
 sg13g2_decap_8 FILLER_79_1701 ();
 sg13g2_decap_8 FILLER_79_1708 ();
 sg13g2_decap_8 FILLER_79_1715 ();
 sg13g2_decap_8 FILLER_79_1722 ();
 sg13g2_decap_8 FILLER_79_1729 ();
 sg13g2_decap_8 FILLER_79_1736 ();
 sg13g2_decap_8 FILLER_79_1743 ();
 sg13g2_decap_8 FILLER_79_1750 ();
 sg13g2_decap_8 FILLER_79_1757 ();
 sg13g2_decap_4 FILLER_79_1764 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_fill_1 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_103 ();
 sg13g2_fill_2 FILLER_80_142 ();
 sg13g2_fill_1 FILLER_80_183 ();
 sg13g2_fill_2 FILLER_80_201 ();
 sg13g2_fill_2 FILLER_80_219 ();
 sg13g2_fill_1 FILLER_80_314 ();
 sg13g2_fill_2 FILLER_80_321 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_4 FILLER_80_384 ();
 sg13g2_fill_1 FILLER_80_422 ();
 sg13g2_fill_2 FILLER_80_438 ();
 sg13g2_fill_2 FILLER_80_456 ();
 sg13g2_decap_4 FILLER_80_477 ();
 sg13g2_fill_2 FILLER_80_490 ();
 sg13g2_decap_8 FILLER_80_502 ();
 sg13g2_decap_8 FILLER_80_509 ();
 sg13g2_decap_8 FILLER_80_516 ();
 sg13g2_decap_8 FILLER_80_523 ();
 sg13g2_fill_1 FILLER_80_530 ();
 sg13g2_decap_8 FILLER_80_540 ();
 sg13g2_decap_8 FILLER_80_547 ();
 sg13g2_decap_8 FILLER_80_554 ();
 sg13g2_decap_8 FILLER_80_561 ();
 sg13g2_decap_8 FILLER_80_583 ();
 sg13g2_fill_2 FILLER_80_590 ();
 sg13g2_fill_1 FILLER_80_592 ();
 sg13g2_decap_4 FILLER_80_598 ();
 sg13g2_fill_2 FILLER_80_602 ();
 sg13g2_decap_4 FILLER_80_612 ();
 sg13g2_fill_1 FILLER_80_616 ();
 sg13g2_decap_8 FILLER_80_637 ();
 sg13g2_decap_4 FILLER_80_644 ();
 sg13g2_fill_2 FILLER_80_648 ();
 sg13g2_decap_8 FILLER_80_668 ();
 sg13g2_decap_8 FILLER_80_675 ();
 sg13g2_fill_1 FILLER_80_682 ();
 sg13g2_decap_8 FILLER_80_693 ();
 sg13g2_decap_4 FILLER_80_700 ();
 sg13g2_fill_1 FILLER_80_704 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_728 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_fill_2 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_752 ();
 sg13g2_decap_8 FILLER_80_759 ();
 sg13g2_fill_2 FILLER_80_774 ();
 sg13g2_fill_1 FILLER_80_776 ();
 sg13g2_decap_8 FILLER_80_790 ();
 sg13g2_decap_4 FILLER_80_797 ();
 sg13g2_fill_1 FILLER_80_801 ();
 sg13g2_decap_8 FILLER_80_820 ();
 sg13g2_decap_8 FILLER_80_827 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_decap_8 FILLER_80_861 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_decap_8 FILLER_80_875 ();
 sg13g2_decap_8 FILLER_80_882 ();
 sg13g2_decap_8 FILLER_80_889 ();
 sg13g2_decap_8 FILLER_80_896 ();
 sg13g2_fill_2 FILLER_80_903 ();
 sg13g2_fill_2 FILLER_80_962 ();
 sg13g2_fill_1 FILLER_80_972 ();
 sg13g2_fill_1 FILLER_80_1009 ();
 sg13g2_fill_1 FILLER_80_1019 ();
 sg13g2_decap_8 FILLER_80_1061 ();
 sg13g2_decap_8 FILLER_80_1068 ();
 sg13g2_decap_8 FILLER_80_1075 ();
 sg13g2_decap_8 FILLER_80_1082 ();
 sg13g2_decap_8 FILLER_80_1089 ();
 sg13g2_decap_8 FILLER_80_1096 ();
 sg13g2_decap_8 FILLER_80_1103 ();
 sg13g2_decap_8 FILLER_80_1110 ();
 sg13g2_decap_8 FILLER_80_1117 ();
 sg13g2_decap_8 FILLER_80_1124 ();
 sg13g2_decap_8 FILLER_80_1131 ();
 sg13g2_decap_8 FILLER_80_1138 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_decap_8 FILLER_80_1152 ();
 sg13g2_decap_8 FILLER_80_1159 ();
 sg13g2_decap_8 FILLER_80_1166 ();
 sg13g2_decap_8 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1180 ();
 sg13g2_decap_8 FILLER_80_1187 ();
 sg13g2_decap_8 FILLER_80_1194 ();
 sg13g2_decap_8 FILLER_80_1201 ();
 sg13g2_decap_8 FILLER_80_1208 ();
 sg13g2_decap_8 FILLER_80_1215 ();
 sg13g2_decap_8 FILLER_80_1222 ();
 sg13g2_decap_8 FILLER_80_1229 ();
 sg13g2_decap_8 FILLER_80_1236 ();
 sg13g2_decap_8 FILLER_80_1243 ();
 sg13g2_decap_8 FILLER_80_1250 ();
 sg13g2_decap_8 FILLER_80_1257 ();
 sg13g2_decap_8 FILLER_80_1264 ();
 sg13g2_decap_8 FILLER_80_1271 ();
 sg13g2_decap_8 FILLER_80_1278 ();
 sg13g2_decap_8 FILLER_80_1285 ();
 sg13g2_decap_8 FILLER_80_1292 ();
 sg13g2_decap_8 FILLER_80_1299 ();
 sg13g2_decap_8 FILLER_80_1306 ();
 sg13g2_decap_8 FILLER_80_1313 ();
 sg13g2_decap_8 FILLER_80_1320 ();
 sg13g2_decap_8 FILLER_80_1327 ();
 sg13g2_decap_8 FILLER_80_1334 ();
 sg13g2_decap_8 FILLER_80_1341 ();
 sg13g2_decap_8 FILLER_80_1348 ();
 sg13g2_decap_8 FILLER_80_1355 ();
 sg13g2_decap_8 FILLER_80_1362 ();
 sg13g2_decap_8 FILLER_80_1369 ();
 sg13g2_decap_8 FILLER_80_1376 ();
 sg13g2_decap_8 FILLER_80_1383 ();
 sg13g2_decap_8 FILLER_80_1390 ();
 sg13g2_decap_8 FILLER_80_1397 ();
 sg13g2_decap_8 FILLER_80_1404 ();
 sg13g2_decap_8 FILLER_80_1411 ();
 sg13g2_decap_8 FILLER_80_1418 ();
 sg13g2_decap_8 FILLER_80_1425 ();
 sg13g2_decap_8 FILLER_80_1432 ();
 sg13g2_decap_8 FILLER_80_1439 ();
 sg13g2_decap_8 FILLER_80_1446 ();
 sg13g2_decap_8 FILLER_80_1453 ();
 sg13g2_decap_8 FILLER_80_1460 ();
 sg13g2_decap_8 FILLER_80_1467 ();
 sg13g2_decap_8 FILLER_80_1474 ();
 sg13g2_decap_8 FILLER_80_1481 ();
 sg13g2_decap_8 FILLER_80_1488 ();
 sg13g2_decap_8 FILLER_80_1495 ();
 sg13g2_decap_8 FILLER_80_1502 ();
 sg13g2_decap_8 FILLER_80_1509 ();
 sg13g2_decap_8 FILLER_80_1516 ();
 sg13g2_decap_8 FILLER_80_1523 ();
 sg13g2_decap_8 FILLER_80_1530 ();
 sg13g2_decap_8 FILLER_80_1537 ();
 sg13g2_decap_8 FILLER_80_1544 ();
 sg13g2_decap_8 FILLER_80_1551 ();
 sg13g2_decap_8 FILLER_80_1558 ();
 sg13g2_decap_8 FILLER_80_1565 ();
 sg13g2_decap_8 FILLER_80_1572 ();
 sg13g2_decap_8 FILLER_80_1579 ();
 sg13g2_decap_8 FILLER_80_1586 ();
 sg13g2_decap_8 FILLER_80_1593 ();
 sg13g2_decap_8 FILLER_80_1600 ();
 sg13g2_decap_8 FILLER_80_1607 ();
 sg13g2_decap_8 FILLER_80_1614 ();
 sg13g2_decap_8 FILLER_80_1621 ();
 sg13g2_decap_8 FILLER_80_1628 ();
 sg13g2_decap_8 FILLER_80_1635 ();
 sg13g2_decap_8 FILLER_80_1642 ();
 sg13g2_decap_8 FILLER_80_1649 ();
 sg13g2_decap_8 FILLER_80_1656 ();
 sg13g2_decap_8 FILLER_80_1663 ();
 sg13g2_decap_8 FILLER_80_1670 ();
 sg13g2_decap_8 FILLER_80_1677 ();
 sg13g2_decap_8 FILLER_80_1684 ();
 sg13g2_decap_8 FILLER_80_1691 ();
 sg13g2_decap_8 FILLER_80_1698 ();
 sg13g2_decap_8 FILLER_80_1705 ();
 sg13g2_decap_8 FILLER_80_1712 ();
 sg13g2_decap_8 FILLER_80_1719 ();
 sg13g2_decap_8 FILLER_80_1726 ();
 sg13g2_decap_8 FILLER_80_1733 ();
 sg13g2_decap_8 FILLER_80_1740 ();
 sg13g2_decap_8 FILLER_80_1747 ();
 sg13g2_decap_8 FILLER_80_1754 ();
 sg13g2_decap_8 FILLER_80_1761 ();
 assign uo_out[6] = net12;
 assign uo_out[7] = net13;
endmodule

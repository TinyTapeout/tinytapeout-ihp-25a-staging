module tt_um_hack_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire clk_regs;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire \cpu.alu_instance.a_i[0] ;
 wire \cpu.alu_instance.a_i[10] ;
 wire \cpu.alu_instance.a_i[11] ;
 wire \cpu.alu_instance.a_i[12] ;
 wire \cpu.alu_instance.a_i[13] ;
 wire \cpu.alu_instance.a_i[14] ;
 wire \cpu.alu_instance.a_i[15] ;
 wire \cpu.alu_instance.a_i[1] ;
 wire \cpu.alu_instance.a_i[2] ;
 wire \cpu.alu_instance.a_i[3] ;
 wire \cpu.alu_instance.a_i[4] ;
 wire \cpu.alu_instance.a_i[5] ;
 wire \cpu.alu_instance.a_i[6] ;
 wire \cpu.alu_instance.a_i[7] ;
 wire \cpu.alu_instance.a_i[8] ;
 wire \cpu.alu_instance.a_i[9] ;
 wire \cpu.alu_instance.f_i ;
 wire \cpu.alu_instance.na_i ;
 wire \cpu.alu_instance.nb_i ;
 wire \cpu.alu_instance.no_i ;
 wire \cpu.alu_instance.za_i ;
 wire \cpu.alu_instance.zb_i ;
 wire \cpu.debug_out_o ;
 wire \cpu.fsm_instance.instruction_i[0] ;
 wire \cpu.fsm_instance.instruction_i[12] ;
 wire \cpu.fsm_instance.instruction_i[13] ;
 wire \cpu.fsm_instance.instruction_i[14] ;
 wire \cpu.fsm_instance.instruction_i[15] ;
 wire \cpu.fsm_instance.instruction_i[1] ;
 wire \cpu.fsm_instance.instruction_i[2] ;
 wire \cpu.fsm_instance.instruction_i[3] ;
 wire \cpu.fsm_instance.instruction_i[4] ;
 wire \cpu.fsm_instance.instruction_i[5] ;
 wire \cpu.fsm_instance.state_s[0] ;
 wire \cpu.fsm_instance.state_s[1] ;
 wire \cpu.inM_s[0] ;
 wire \cpu.inM_s[10] ;
 wire \cpu.inM_s[11] ;
 wire \cpu.inM_s[12] ;
 wire \cpu.inM_s[13] ;
 wire \cpu.inM_s[14] ;
 wire \cpu.inM_s[15] ;
 wire \cpu.inM_s[1] ;
 wire \cpu.inM_s[2] ;
 wire \cpu.inM_s[3] ;
 wire \cpu.inM_s[4] ;
 wire \cpu.inM_s[5] ;
 wire \cpu.inM_s[6] ;
 wire \cpu.inM_s[7] ;
 wire \cpu.inM_s[8] ;
 wire \cpu.inM_s[9] ;
 wire \cpu.mem_csb_o ;
 wire \cpu.mem_out_o ;
 wire \cpu.mem_sclk_o ;
 wire \cpu.pc_s[0] ;
 wire \cpu.pc_s[10] ;
 wire \cpu.pc_s[11] ;
 wire \cpu.pc_s[12] ;
 wire \cpu.pc_s[13] ;
 wire \cpu.pc_s[14] ;
 wire \cpu.pc_s[15] ;
 wire \cpu.pc_s[1] ;
 wire \cpu.pc_s[2] ;
 wire \cpu.pc_s[3] ;
 wire \cpu.pc_s[4] ;
 wire \cpu.pc_s[5] ;
 wire \cpu.pc_s[6] ;
 wire \cpu.pc_s[7] ;
 wire \cpu.pc_s[8] ;
 wire \cpu.pc_s[9] ;
 wire \cpu.regA_s[0] ;
 wire \cpu.regA_s[10] ;
 wire \cpu.regA_s[11] ;
 wire \cpu.regA_s[12] ;
 wire \cpu.regA_s[13] ;
 wire \cpu.regA_s[14] ;
 wire \cpu.regA_s[15] ;
 wire \cpu.regA_s[1] ;
 wire \cpu.regA_s[2] ;
 wire \cpu.regA_s[3] ;
 wire \cpu.regA_s[4] ;
 wire \cpu.regA_s[5] ;
 wire \cpu.regA_s[6] ;
 wire \cpu.regA_s[7] ;
 wire \cpu.regA_s[8] ;
 wire \cpu.regA_s[9] ;
 wire \cpu.spi_debug_instance.counter_s[0] ;
 wire \cpu.spi_debug_instance.counter_s[1] ;
 wire \cpu.spi_debug_instance.counter_s[2] ;
 wire \cpu.spi_debug_instance.counter_s[3] ;
 wire \cpu.spi_debug_instance.counter_s[4] ;
 wire \cpu.spi_debug_instance.in_s[0] ;
 wire \cpu.spi_debug_instance.in_s[1] ;
 wire \cpu.spi_mem_instance.count_s[0] ;
 wire \cpu.spi_mem_instance.count_s[1] ;
 wire \cpu.spi_mem_instance.count_s[2] ;
 wire \cpu.spi_mem_instance.count_s[3] ;
 wire \cpu.spi_mem_instance.count_s[4] ;
 wire \cpu.spi_mem_instance.count_s[5] ;
 wire \cpu.spi_mem_instance.next_state_s[0] ;
 wire \cpu.spi_mem_instance.next_state_s[1] ;
 wire \cpu.spi_mem_instance.next_state_s[2] ;
 wire \cpu.spi_mem_instance.state_s[0] ;
 wire \cpu.spi_mem_instance.state_s[1] ;
 wire \cpu.spi_mem_instance.state_s[2] ;
 wire net23;
 wire net24;
 wire net7;
 wire net25;
 wire net8;
 wire net9;
 wire net26;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net27;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire delaynet_0_clk;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;

 sg13g2_inv_1 _0733_ (.Y(_0115_),
    .A(\cpu.spi_mem_instance.count_s[5] ));
 sg13g2_inv_2 _0734_ (.Y(_0116_),
    .A(net141));
 sg13g2_inv_1 _0735_ (.Y(_0117_),
    .A(\cpu.spi_debug_instance.counter_s[1] ));
 sg13g2_inv_2 _0736_ (.Y(_0118_),
    .A(\cpu.spi_debug_instance.counter_s[0] ));
 sg13g2_inv_1 _0737_ (.Y(_0119_),
    .A(net82));
 sg13g2_inv_4 _0738_ (.A(net306),
    .Y(_0120_));
 sg13g2_inv_1 _0739_ (.Y(_0121_),
    .A(net44));
 sg13g2_inv_1 _0740_ (.Y(_0122_),
    .A(\cpu.alu_instance.zb_i ));
 sg13g2_inv_1 _0741_ (.Y(_0123_),
    .A(net311));
 sg13g2_inv_1 _0742_ (.Y(_0124_),
    .A(\cpu.inM_s[14] ));
 sg13g2_inv_1 _0743_ (.Y(_0125_),
    .A(net39));
 sg13g2_inv_1 _0744_ (.Y(_0126_),
    .A(\cpu.inM_s[12] ));
 sg13g2_inv_4 _0745_ (.A(net291),
    .Y(_0127_));
 sg13g2_inv_1 _0746_ (.Y(_0128_),
    .A(net59));
 sg13g2_inv_1 _0747_ (.Y(_0129_),
    .A(\cpu.fsm_instance.instruction_i[1] ));
 sg13g2_inv_1 _0748_ (.Y(_0130_),
    .A(net139));
 sg13g2_inv_1 _0749_ (.Y(_0131_),
    .A(net140));
 sg13g2_inv_1 _0750_ (.Y(_0132_),
    .A(net124));
 sg13g2_inv_1 _0751_ (.Y(_0133_),
    .A(net112));
 sg13g2_inv_1 _0752_ (.Y(_0134_),
    .A(\cpu.pc_s[14] ));
 sg13g2_inv_1 _1370__3 (.Y(net28),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _0754_ (.Y(_0009_),
    .A(net5));
 sg13g2_nor2b_2 _0755_ (.A(net95),
    .B_N(net33),
    .Y(_0135_));
 sg13g2_nand2_2 _0756_ (.Y(_0136_),
    .A(net82),
    .B(_0135_));
 sg13g2_nand2_1 _0757_ (.Y(_0137_),
    .A(\cpu.spi_mem_instance.state_s[1] ),
    .B(net33));
 sg13g2_nor2_1 _0758_ (.A(net82),
    .B(net34),
    .Y(_0138_));
 sg13g2_o21ai_1 _0759_ (.B1(_0136_),
    .Y(_0139_),
    .A1(\cpu.spi_mem_instance.state_s[0] ),
    .A2(_0137_));
 sg13g2_inv_2 _0760_ (.Y(\cpu.mem_csb_o ),
    .A(_0139_));
 sg13g2_nor2_1 _0761_ (.A(\cpu.spi_mem_instance.count_s[2] ),
    .B(net271),
    .Y(_0140_));
 sg13g2_nor2_1 _0762_ (.A(net275),
    .B(\cpu.mem_csb_o ),
    .Y(_0141_));
 sg13g2_nor3_1 _0763_ (.A(net270),
    .B(net275),
    .C(\cpu.mem_csb_o ),
    .Y(_0142_));
 sg13g2_nand2_1 _0764_ (.Y(_0143_),
    .A(_0116_),
    .B(_0142_));
 sg13g2_nor3_2 _0765_ (.A(net98),
    .B(\cpu.spi_mem_instance.count_s[2] ),
    .C(net270),
    .Y(_0144_));
 sg13g2_nand2_2 _0766_ (.Y(_0145_),
    .A(_0141_),
    .B(_0144_));
 sg13g2_nor3_1 _0767_ (.A(net107),
    .B(net128),
    .C(_0145_),
    .Y(_0146_));
 sg13g2_or3_1 _0768_ (.A(net107),
    .B(\cpu.spi_mem_instance.count_s[4] ),
    .C(_0145_),
    .X(_0147_));
 sg13g2_o21ai_1 _0769_ (.B1(net107),
    .Y(_0148_),
    .A1(\cpu.spi_mem_instance.count_s[4] ),
    .A2(_0145_));
 sg13g2_nand2_1 _0770_ (.Y(_0113_),
    .A(_0147_),
    .B(net108));
 sg13g2_xor2_1 _0771_ (.B(_0145_),
    .A(net128),
    .X(_0149_));
 sg13g2_nor2_1 _0772_ (.A(_0146_),
    .B(_0149_),
    .Y(_0112_));
 sg13g2_nand2_1 _0773_ (.Y(_0150_),
    .A(net98),
    .B(_0143_));
 sg13g2_a21oi_1 _0774_ (.A1(_0145_),
    .A2(_0150_),
    .Y(_0111_),
    .B1(_0146_));
 sg13g2_xnor2_1 _0775_ (.Y(_0110_),
    .A(_0116_),
    .B(_0142_));
 sg13g2_xor2_1 _0776_ (.B(net119),
    .A(net270),
    .X(_0109_));
 sg13g2_nand2_1 _0777_ (.Y(_0151_),
    .A(net275),
    .B(\cpu.mem_csb_o ));
 sg13g2_nand2_1 _0778_ (.Y(_0152_),
    .A(net36),
    .B(_0139_));
 sg13g2_nand3_1 _0779_ (.B(_0151_),
    .C(_0152_),
    .A(_0147_),
    .Y(_0108_));
 sg13g2_nor2_1 _0780_ (.A(\cpu.spi_debug_instance.counter_s[4] ),
    .B(\cpu.spi_debug_instance.counter_s[3] ),
    .Y(_0153_));
 sg13g2_nand2_2 _0781_ (.Y(_0154_),
    .A(_0117_),
    .B(_0118_));
 sg13g2_or2_1 _0782_ (.X(_0155_),
    .B(_0154_),
    .A(net3));
 sg13g2_nor2_1 _0783_ (.A(\cpu.spi_debug_instance.counter_s[2] ),
    .B(_0155_),
    .Y(_0156_));
 sg13g2_inv_1 _0784_ (.Y(_0157_),
    .A(_0156_));
 sg13g2_nor3_1 _0785_ (.A(\cpu.spi_debug_instance.counter_s[4] ),
    .B(net276),
    .C(\cpu.spi_debug_instance.counter_s[2] ),
    .Y(_0158_));
 sg13g2_nand2_1 _0786_ (.Y(_0159_),
    .A(_0153_),
    .B(_0156_));
 sg13g2_o21ai_1 _0787_ (.B1(\cpu.spi_debug_instance.counter_s[4] ),
    .Y(_0160_),
    .A1(net276),
    .A2(_0157_));
 sg13g2_nand2_1 _0788_ (.Y(_0056_),
    .A(_0159_),
    .B(_0160_));
 sg13g2_a21oi_1 _0789_ (.A1(\cpu.spi_debug_instance.counter_s[4] ),
    .A2(_0156_),
    .Y(_0161_),
    .B1(net276));
 sg13g2_a21oi_1 _0790_ (.A1(net276),
    .A2(_0156_),
    .Y(_0055_),
    .B1(_0161_));
 sg13g2_nand2_1 _0791_ (.Y(_0162_),
    .A(\cpu.spi_debug_instance.counter_s[2] ),
    .B(_0155_));
 sg13g2_o21ai_1 _0792_ (.B1(_0162_),
    .Y(_0054_),
    .A1(_0153_),
    .A2(_0157_));
 sg13g2_o21ai_1 _0793_ (.B1(\cpu.spi_debug_instance.counter_s[1] ),
    .Y(_0163_),
    .A1(net3),
    .A2(\cpu.spi_debug_instance.counter_s[0] ));
 sg13g2_o21ai_1 _0794_ (.B1(_0163_),
    .Y(_0053_),
    .A1(_0155_),
    .A2(_0158_));
 sg13g2_nor2b_1 _0795_ (.A(net3),
    .B_N(_0008_),
    .Y(_0164_));
 sg13g2_a21oi_1 _0796_ (.A1(net3),
    .A2(\cpu.spi_debug_instance.counter_s[0] ),
    .Y(_0165_),
    .B1(_0164_));
 sg13g2_nand2_1 _0797_ (.Y(_0052_),
    .A(_0159_),
    .B(_0165_));
 sg13g2_nand2b_1 _0798_ (.Y(_0166_),
    .B(_0135_),
    .A_N(net317));
 sg13g2_nand3_1 _0799_ (.B(_0147_),
    .C(_0166_),
    .A(net83),
    .Y(\cpu.spi_mem_instance.next_state_s[0] ));
 sg13g2_nor4_1 _0800_ (.A(\cpu.spi_mem_instance.count_s[5] ),
    .B(\cpu.spi_mem_instance.count_s[4] ),
    .C(net272),
    .D(_0136_),
    .Y(_0167_));
 sg13g2_nand4_1 _0801_ (.B(net313),
    .C(_0119_),
    .A(net317),
    .Y(_0168_),
    .D(_0135_));
 sg13g2_a21oi_1 _0802_ (.A1(_0144_),
    .A2(_0167_),
    .Y(_0169_),
    .B1(_0138_));
 sg13g2_nand2_1 _0803_ (.Y(\cpu.spi_mem_instance.next_state_s[1] ),
    .A(_0168_),
    .B(_0169_));
 sg13g2_nor2b_2 _0804_ (.A(net313),
    .B_N(net317),
    .Y(_0170_));
 sg13g2_nand2b_2 _0805_ (.Y(_0171_),
    .B(net317),
    .A_N(net313));
 sg13g2_nor3_1 _0806_ (.A(_0119_),
    .B(net34),
    .C(_0171_),
    .Y(\cpu.spi_mem_instance.next_state_s[2] ));
 sg13g2_nor2b_1 _0807_ (.A(net299),
    .B_N(\cpu.alu_instance.a_i[14] ),
    .Y(_0172_));
 sg13g2_xnor2_1 _0808_ (.Y(_0173_),
    .A(net298),
    .B(_0172_));
 sg13g2_a21oi_1 _0809_ (.A1(net302),
    .A2(_0124_),
    .Y(_0174_),
    .B1(\cpu.alu_instance.zb_i ));
 sg13g2_o21ai_1 _0810_ (.B1(_0174_),
    .Y(_0175_),
    .A1(net302),
    .A2(\cpu.regA_s[14] ));
 sg13g2_xnor2_1 _0811_ (.Y(_0176_),
    .A(net285),
    .B(_0175_));
 sg13g2_nand2_1 _0812_ (.Y(_0177_),
    .A(_0173_),
    .B(_0176_));
 sg13g2_nor2_1 _0813_ (.A(net291),
    .B(_0177_),
    .Y(_0178_));
 sg13g2_nor2b_1 _0814_ (.A(net301),
    .B_N(\cpu.alu_instance.a_i[1] ),
    .Y(_0179_));
 sg13g2_xnor2_1 _0815_ (.Y(_0180_),
    .A(net297),
    .B(_0179_));
 sg13g2_mux2_1 _0816_ (.A0(\cpu.regA_s[1] ),
    .A1(\cpu.inM_s[1] ),
    .S(net304),
    .X(_0181_));
 sg13g2_a21o_1 _0817_ (.A2(_0181_),
    .A1(net287),
    .B1(net283),
    .X(_0182_));
 sg13g2_nand3_1 _0818_ (.B(net283),
    .C(_0181_),
    .A(net287),
    .Y(_0183_));
 sg13g2_and3_1 _0819_ (.X(_0184_),
    .A(_0180_),
    .B(_0182_),
    .C(_0183_));
 sg13g2_nand3_1 _0820_ (.B(_0182_),
    .C(_0183_),
    .A(_0180_),
    .Y(_0185_));
 sg13g2_nor2b_1 _0821_ (.A(net300),
    .B_N(\cpu.alu_instance.a_i[0] ),
    .Y(_0186_));
 sg13g2_xnor2_1 _0822_ (.Y(_0187_),
    .A(_0004_),
    .B(_0186_));
 sg13g2_mux2_1 _0823_ (.A0(\cpu.regA_s[0] ),
    .A1(\cpu.inM_s[0] ),
    .S(net305),
    .X(_0188_));
 sg13g2_a21o_1 _0824_ (.A2(_0188_),
    .A1(net288),
    .B1(net283),
    .X(_0189_));
 sg13g2_nand3_1 _0825_ (.B(net283),
    .C(_0188_),
    .A(net288),
    .Y(_0190_));
 sg13g2_nand3_1 _0826_ (.B(_0189_),
    .C(_0190_),
    .A(_0187_),
    .Y(_0191_));
 sg13g2_a21oi_1 _0827_ (.A1(_0182_),
    .A2(_0183_),
    .Y(_0192_),
    .B1(_0180_));
 sg13g2_nor2_1 _0828_ (.A(_0184_),
    .B(_0192_),
    .Y(_0193_));
 sg13g2_o21ai_1 _0829_ (.B1(_0185_),
    .Y(_0194_),
    .A1(_0191_),
    .A2(_0192_));
 sg13g2_nor2b_1 _0830_ (.A(net301),
    .B_N(\cpu.alu_instance.a_i[2] ),
    .Y(_0195_));
 sg13g2_xnor2_1 _0831_ (.Y(_0196_),
    .A(net297),
    .B(_0195_));
 sg13g2_mux2_1 _0832_ (.A0(\cpu.regA_s[2] ),
    .A1(\cpu.inM_s[2] ),
    .S(net304),
    .X(_0197_));
 sg13g2_a21o_1 _0833_ (.A2(_0197_),
    .A1(net286),
    .B1(net284),
    .X(_0198_));
 sg13g2_nand3_1 _0834_ (.B(net284),
    .C(_0197_),
    .A(net286),
    .Y(_0199_));
 sg13g2_and3_1 _0835_ (.X(_0200_),
    .A(_0196_),
    .B(_0198_),
    .C(_0199_));
 sg13g2_a21oi_1 _0836_ (.A1(_0198_),
    .A2(_0199_),
    .Y(_0201_),
    .B1(_0196_));
 sg13g2_nor2_1 _0837_ (.A(_0200_),
    .B(_0201_),
    .Y(_0202_));
 sg13g2_nand2b_1 _0838_ (.Y(_0203_),
    .B(\cpu.alu_instance.a_i[3] ),
    .A_N(net300));
 sg13g2_xnor2_1 _0839_ (.Y(_0204_),
    .A(net297),
    .B(_0203_));
 sg13g2_mux2_1 _0840_ (.A0(\cpu.regA_s[3] ),
    .A1(\cpu.inM_s[3] ),
    .S(net305),
    .X(_0205_));
 sg13g2_a21o_1 _0841_ (.A2(_0205_),
    .A1(net286),
    .B1(net311),
    .X(_0206_));
 sg13g2_nand3_1 _0842_ (.B(net311),
    .C(_0205_),
    .A(net286),
    .Y(_0207_));
 sg13g2_a21oi_1 _0843_ (.A1(net286),
    .A2(_0205_),
    .Y(_0208_),
    .B1(net284));
 sg13g2_and3_1 _0844_ (.X(_0209_),
    .A(net286),
    .B(net284),
    .C(_0205_));
 sg13g2_nor3_1 _0845_ (.A(_0204_),
    .B(_0208_),
    .C(_0209_),
    .Y(_0210_));
 sg13g2_and3_1 _0846_ (.X(_0211_),
    .A(_0204_),
    .B(_0206_),
    .C(_0207_));
 sg13g2_o21ai_1 _0847_ (.B1(_0204_),
    .Y(_0212_),
    .A1(_0208_),
    .A2(_0209_));
 sg13g2_nor4_1 _0848_ (.A(_0200_),
    .B(_0201_),
    .C(_0210_),
    .D(_0211_),
    .Y(_0213_));
 sg13g2_a221oi_1 _0849_ (.B2(_0194_),
    .C1(_0210_),
    .B1(_0213_),
    .A1(_0200_),
    .Y(_0214_),
    .A2(_0212_));
 sg13g2_nand2b_1 _0850_ (.Y(_0215_),
    .B(\cpu.alu_instance.a_i[6] ),
    .A_N(net300));
 sg13g2_xnor2_1 _0851_ (.Y(_0216_),
    .A(net297),
    .B(_0215_));
 sg13g2_mux2_1 _0852_ (.A0(\cpu.regA_s[6] ),
    .A1(\cpu.inM_s[6] ),
    .S(net304),
    .X(_0217_));
 sg13g2_a21o_1 _0853_ (.A2(_0217_),
    .A1(net289),
    .B1(net311),
    .X(_0218_));
 sg13g2_nand3_1 _0854_ (.B(net311),
    .C(_0217_),
    .A(net288),
    .Y(_0219_));
 sg13g2_a21oi_2 _0855_ (.B1(_0216_),
    .Y(_0220_),
    .A2(_0219_),
    .A1(_0218_));
 sg13g2_and3_1 _0856_ (.X(_0221_),
    .A(_0216_),
    .B(_0218_),
    .C(_0219_));
 sg13g2_nor2_1 _0857_ (.A(_0220_),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_nand2b_1 _0858_ (.Y(_0223_),
    .B(\cpu.alu_instance.a_i[7] ),
    .A_N(net300));
 sg13g2_xnor2_1 _0859_ (.Y(_0224_),
    .A(net297),
    .B(_0223_));
 sg13g2_mux2_1 _0860_ (.A0(\cpu.regA_s[7] ),
    .A1(\cpu.inM_s[7] ),
    .S(net304),
    .X(_0225_));
 sg13g2_a21o_1 _0861_ (.A2(_0225_),
    .A1(net288),
    .B1(net311),
    .X(_0226_));
 sg13g2_nand3_1 _0862_ (.B(net311),
    .C(_0225_),
    .A(net288),
    .Y(_0227_));
 sg13g2_a21oi_1 _0863_ (.A1(net288),
    .A2(_0225_),
    .Y(_0228_),
    .B1(net283));
 sg13g2_and3_1 _0864_ (.X(_0229_),
    .A(net288),
    .B(net283),
    .C(_0225_));
 sg13g2_nor3_1 _0865_ (.A(_0224_),
    .B(_0228_),
    .C(_0229_),
    .Y(_0230_));
 sg13g2_and3_1 _0866_ (.X(_0231_),
    .A(_0224_),
    .B(_0226_),
    .C(_0227_));
 sg13g2_o21ai_1 _0867_ (.B1(_0224_),
    .Y(_0232_),
    .A1(_0228_),
    .A2(_0229_));
 sg13g2_nor2_1 _0868_ (.A(_0230_),
    .B(_0231_),
    .Y(_0233_));
 sg13g2_nor3_1 _0869_ (.A(_0220_),
    .B(_0221_),
    .C(_0231_),
    .Y(_0234_));
 sg13g2_nor2b_1 _0870_ (.A(net300),
    .B_N(\cpu.alu_instance.a_i[5] ),
    .Y(_0235_));
 sg13g2_xnor2_1 _0871_ (.Y(_0236_),
    .A(net297),
    .B(_0235_));
 sg13g2_mux2_1 _0872_ (.A0(\cpu.regA_s[5] ),
    .A1(\cpu.inM_s[5] ),
    .S(net304),
    .X(_0237_));
 sg13g2_a21o_1 _0873_ (.A2(_0237_),
    .A1(net287),
    .B1(net283),
    .X(_0238_));
 sg13g2_nand3_1 _0874_ (.B(net283),
    .C(_0237_),
    .A(net287),
    .Y(_0239_));
 sg13g2_and3_1 _0875_ (.X(_0240_),
    .A(_0236_),
    .B(_0238_),
    .C(_0239_));
 sg13g2_nand3_1 _0876_ (.B(_0238_),
    .C(_0239_),
    .A(_0236_),
    .Y(_0241_));
 sg13g2_a21oi_1 _0877_ (.A1(_0238_),
    .A2(_0239_),
    .Y(_0242_),
    .B1(_0236_));
 sg13g2_nor2_2 _0878_ (.A(_0240_),
    .B(_0242_),
    .Y(_0243_));
 sg13g2_nor2b_1 _0879_ (.A(net300),
    .B_N(\cpu.alu_instance.a_i[4] ),
    .Y(_0244_));
 sg13g2_xnor2_1 _0880_ (.Y(_0245_),
    .A(net297),
    .B(_0244_));
 sg13g2_mux2_1 _0881_ (.A0(\cpu.regA_s[4] ),
    .A1(\cpu.inM_s[4] ),
    .S(net304),
    .X(_0246_));
 sg13g2_a21oi_1 _0882_ (.A1(net286),
    .A2(_0246_),
    .Y(_0247_),
    .B1(net312));
 sg13g2_and3_1 _0883_ (.X(_0248_),
    .A(net286),
    .B(net311),
    .C(_0246_));
 sg13g2_nor2_1 _0884_ (.A(_0247_),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_o21ai_1 _0885_ (.B1(_0245_),
    .Y(_0250_),
    .A1(_0247_),
    .A2(_0248_));
 sg13g2_xnor2_1 _0886_ (.Y(_0251_),
    .A(_0245_),
    .B(_0249_));
 sg13g2_inv_1 _0887_ (.Y(_0252_),
    .A(_0251_));
 sg13g2_nand4_1 _0888_ (.B(_0233_),
    .C(_0243_),
    .A(_0222_),
    .Y(_0253_),
    .D(_0251_));
 sg13g2_a21oi_1 _0889_ (.A1(_0241_),
    .A2(_0250_),
    .Y(_0254_),
    .B1(_0242_));
 sg13g2_a221oi_1 _0890_ (.B2(_0254_),
    .C1(_0230_),
    .B1(_0234_),
    .A1(_0220_),
    .Y(_0255_),
    .A2(_0232_));
 sg13g2_o21ai_1 _0891_ (.B1(_0255_),
    .Y(_0256_),
    .A1(_0214_),
    .A2(_0253_));
 sg13g2_nor2b_1 _0892_ (.A(net300),
    .B_N(\cpu.alu_instance.a_i[8] ),
    .Y(_0257_));
 sg13g2_xnor2_1 _0893_ (.Y(_0258_),
    .A(net297),
    .B(_0257_));
 sg13g2_mux2_1 _0894_ (.A0(\cpu.regA_s[8] ),
    .A1(\cpu.inM_s[8] ),
    .S(net304),
    .X(_0259_));
 sg13g2_a21oi_1 _0895_ (.A1(net289),
    .A2(_0259_),
    .Y(_0260_),
    .B1(net312));
 sg13g2_and3_1 _0896_ (.X(_0261_),
    .A(net289),
    .B(net312),
    .C(_0259_));
 sg13g2_nor2_1 _0897_ (.A(_0260_),
    .B(_0261_),
    .Y(_0262_));
 sg13g2_o21ai_1 _0898_ (.B1(_0258_),
    .Y(_0263_),
    .A1(_0260_),
    .A2(_0261_));
 sg13g2_xnor2_1 _0899_ (.Y(_0264_),
    .A(_0258_),
    .B(_0262_));
 sg13g2_nand2_1 _0900_ (.Y(_0265_),
    .A(_0256_),
    .B(_0264_));
 sg13g2_nor2b_1 _0901_ (.A(net299),
    .B_N(\cpu.alu_instance.a_i[10] ),
    .Y(_0266_));
 sg13g2_xnor2_1 _0902_ (.Y(_0267_),
    .A(net298),
    .B(_0266_));
 sg13g2_nor2b_1 _0903_ (.A(\cpu.inM_s[10] ),
    .B_N(net303),
    .Y(_0268_));
 sg13g2_nor2_1 _0904_ (.A(net303),
    .B(\cpu.regA_s[10] ),
    .Y(_0269_));
 sg13g2_nor3_1 _0905_ (.A(\cpu.alu_instance.zb_i ),
    .B(_0268_),
    .C(_0269_),
    .Y(_0270_));
 sg13g2_xnor2_1 _0906_ (.Y(_0271_),
    .A(net312),
    .B(_0270_));
 sg13g2_nand2_1 _0907_ (.Y(_0272_),
    .A(_0267_),
    .B(_0271_));
 sg13g2_xor2_1 _0908_ (.B(_0271_),
    .A(_0267_),
    .X(_0273_));
 sg13g2_inv_1 _0909_ (.Y(_0274_),
    .A(_0273_));
 sg13g2_nor2b_1 _0910_ (.A(net299),
    .B_N(\cpu.alu_instance.a_i[11] ),
    .Y(_0275_));
 sg13g2_xnor2_1 _0911_ (.Y(_0276_),
    .A(net298),
    .B(_0275_));
 sg13g2_inv_1 _0912_ (.Y(_0277_),
    .A(_0276_));
 sg13g2_nor2b_1 _0913_ (.A(\cpu.inM_s[11] ),
    .B_N(net305),
    .Y(_0278_));
 sg13g2_nor2_1 _0914_ (.A(net303),
    .B(\cpu.regA_s[11] ),
    .Y(_0279_));
 sg13g2_nor3_1 _0915_ (.A(\cpu.alu_instance.zb_i ),
    .B(_0278_),
    .C(_0279_),
    .Y(_0280_));
 sg13g2_xnor2_1 _0916_ (.Y(_0281_),
    .A(net285),
    .B(_0280_));
 sg13g2_nor2_1 _0917_ (.A(_0277_),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_and2_1 _0918_ (.A(_0277_),
    .B(_0281_),
    .X(_0283_));
 sg13g2_xnor2_1 _0919_ (.Y(_0284_),
    .A(_0276_),
    .B(_0281_));
 sg13g2_nor2b_1 _0920_ (.A(net300),
    .B_N(\cpu.alu_instance.a_i[9] ),
    .Y(_0285_));
 sg13g2_xnor2_1 _0921_ (.Y(_0286_),
    .A(net298),
    .B(_0285_));
 sg13g2_mux2_1 _0922_ (.A0(\cpu.regA_s[9] ),
    .A1(\cpu.inM_s[9] ),
    .S(net304),
    .X(_0287_));
 sg13g2_a21o_1 _0923_ (.A2(_0287_),
    .A1(net290),
    .B1(net285),
    .X(_0288_));
 sg13g2_nand3_1 _0924_ (.B(net285),
    .C(_0287_),
    .A(net290),
    .Y(_0289_));
 sg13g2_and2_1 _0925_ (.A(_0288_),
    .B(_0289_),
    .X(_0290_));
 sg13g2_and2_1 _0926_ (.A(_0286_),
    .B(_0290_),
    .X(_0291_));
 sg13g2_nand3_1 _0927_ (.B(_0288_),
    .C(_0289_),
    .A(_0286_),
    .Y(_0292_));
 sg13g2_a21oi_1 _0928_ (.A1(_0288_),
    .A2(_0289_),
    .Y(_0293_),
    .B1(_0286_));
 sg13g2_xnor2_1 _0929_ (.Y(_0294_),
    .A(_0286_),
    .B(_0290_));
 sg13g2_inv_1 _0930_ (.Y(_0295_),
    .A(_0294_));
 sg13g2_and4_1 _0931_ (.A(_0264_),
    .B(_0273_),
    .C(_0284_),
    .D(_0295_),
    .X(_0296_));
 sg13g2_nor2_1 _0932_ (.A(_0263_),
    .B(_0294_),
    .Y(_0297_));
 sg13g2_nor2_1 _0933_ (.A(_0291_),
    .B(_0297_),
    .Y(_0298_));
 sg13g2_o21ai_1 _0934_ (.B1(_0292_),
    .Y(_0299_),
    .A1(_0263_),
    .A2(_0293_));
 sg13g2_nand3_1 _0935_ (.B(_0284_),
    .C(_0299_),
    .A(_0273_),
    .Y(_0300_));
 sg13g2_or2_1 _0936_ (.X(_0301_),
    .B(_0283_),
    .A(_0272_));
 sg13g2_nand3b_1 _0937_ (.B(_0300_),
    .C(_0301_),
    .Y(_0302_),
    .A_N(_0282_));
 sg13g2_a21oi_2 _0938_ (.B1(_0302_),
    .Y(_0303_),
    .A2(_0296_),
    .A1(_0256_));
 sg13g2_nor2b_1 _0939_ (.A(net301),
    .B_N(\cpu.alu_instance.a_i[12] ),
    .Y(_0304_));
 sg13g2_xnor2_1 _0940_ (.Y(_0305_),
    .A(net298),
    .B(_0304_));
 sg13g2_a21oi_1 _0941_ (.A1(net302),
    .A2(_0126_),
    .Y(_0306_),
    .B1(\cpu.alu_instance.zb_i ));
 sg13g2_o21ai_1 _0942_ (.B1(_0306_),
    .Y(_0307_),
    .A1(net305),
    .A2(\cpu.regA_s[12] ));
 sg13g2_xnor2_1 _0943_ (.Y(_0308_),
    .A(net285),
    .B(_0307_));
 sg13g2_nand2_1 _0944_ (.Y(_0309_),
    .A(_0305_),
    .B(_0308_));
 sg13g2_xor2_1 _0945_ (.B(_0308_),
    .A(_0305_),
    .X(_0310_));
 sg13g2_inv_1 _0946_ (.Y(_0311_),
    .A(_0310_));
 sg13g2_nand2b_1 _0947_ (.Y(_0312_),
    .B(_0310_),
    .A_N(_0303_));
 sg13g2_nor2b_1 _0948_ (.A(net299),
    .B_N(\cpu.alu_instance.a_i[13] ),
    .Y(_0313_));
 sg13g2_xnor2_1 _0949_ (.Y(_0314_),
    .A(net298),
    .B(_0313_));
 sg13g2_a21oi_1 _0950_ (.A1(net302),
    .A2(_0125_),
    .Y(_0315_),
    .B1(\cpu.alu_instance.zb_i ));
 sg13g2_o21ai_1 _0951_ (.B1(_0315_),
    .Y(_0316_),
    .A1(net302),
    .A2(\cpu.regA_s[13] ));
 sg13g2_xnor2_1 _0952_ (.Y(_0317_),
    .A(net285),
    .B(_0316_));
 sg13g2_nand2_1 _0953_ (.Y(_0318_),
    .A(_0314_),
    .B(_0317_));
 sg13g2_xnor2_1 _0954_ (.Y(_0319_),
    .A(_0314_),
    .B(_0317_));
 sg13g2_nor3_2 _0955_ (.A(_0303_),
    .B(_0311_),
    .C(_0319_),
    .Y(_0320_));
 sg13g2_or2_1 _0956_ (.X(_0321_),
    .B(_0319_),
    .A(_0309_));
 sg13g2_nand2_1 _0957_ (.Y(_0322_),
    .A(_0318_),
    .B(_0321_));
 sg13g2_xor2_1 _0958_ (.B(_0176_),
    .A(_0173_),
    .X(_0323_));
 sg13g2_nor3_1 _0959_ (.A(_0320_),
    .B(_0322_),
    .C(_0323_),
    .Y(_0324_));
 sg13g2_o21ai_1 _0960_ (.B1(_0323_),
    .Y(_0325_),
    .A1(_0320_),
    .A2(_0322_));
 sg13g2_nor2b_1 _0961_ (.A(_0324_),
    .B_N(_0325_),
    .Y(_0326_));
 sg13g2_a21oi_1 _0962_ (.A1(net291),
    .A2(_0326_),
    .Y(_0327_),
    .B1(_0178_));
 sg13g2_xnor2_1 _0963_ (.Y(_0328_),
    .A(net295),
    .B(_0327_));
 sg13g2_nand3_1 _0964_ (.B(_0177_),
    .C(_0325_),
    .A(net291),
    .Y(_0329_));
 sg13g2_a21oi_1 _0965_ (.A1(_0121_),
    .A2(net303),
    .Y(_0330_),
    .B1(\cpu.alu_instance.zb_i ));
 sg13g2_o21ai_1 _0966_ (.B1(_0330_),
    .Y(_0331_),
    .A1(\cpu.regA_s[15] ),
    .A2(net303));
 sg13g2_xnor2_1 _0967_ (.Y(_0332_),
    .A(net285),
    .B(_0331_));
 sg13g2_nand2b_1 _0968_ (.Y(_0333_),
    .B(\cpu.alu_instance.a_i[15] ),
    .A_N(net299));
 sg13g2_xnor2_1 _0969_ (.Y(_0334_),
    .A(net298),
    .B(_0333_));
 sg13g2_a21oi_1 _0970_ (.A1(net291),
    .A2(_0334_),
    .Y(_0335_),
    .B1(_0332_));
 sg13g2_a21o_1 _0971_ (.A2(_0334_),
    .A1(_0332_),
    .B1(_0335_),
    .X(_0336_));
 sg13g2_xnor2_1 _0972_ (.Y(_0337_),
    .A(net295),
    .B(_0336_));
 sg13g2_xnor2_1 _0973_ (.Y(_0338_),
    .A(_0329_),
    .B(_0337_));
 sg13g2_nor2_1 _0974_ (.A(net291),
    .B(_0318_),
    .Y(_0339_));
 sg13g2_nand3_1 _0975_ (.B(_0312_),
    .C(_0319_),
    .A(_0309_),
    .Y(_0340_));
 sg13g2_nand2_1 _0976_ (.Y(_0341_),
    .A(net291),
    .B(_0321_));
 sg13g2_nor2_1 _0977_ (.A(_0320_),
    .B(_0341_),
    .Y(_0342_));
 sg13g2_a21oi_1 _0978_ (.A1(_0340_),
    .A2(_0342_),
    .Y(_0343_),
    .B1(_0339_));
 sg13g2_xnor2_1 _0979_ (.Y(_0344_),
    .A(net295),
    .B(_0343_));
 sg13g2_nor2_1 _0980_ (.A(net291),
    .B(_0309_),
    .Y(_0345_));
 sg13g2_a21oi_1 _0981_ (.A1(_0303_),
    .A2(_0311_),
    .Y(_0346_),
    .B1(_0127_));
 sg13g2_a21oi_1 _0982_ (.A1(_0312_),
    .A2(_0346_),
    .Y(_0347_),
    .B1(_0345_));
 sg13g2_xnor2_1 _0983_ (.Y(_0348_),
    .A(net295),
    .B(_0347_));
 sg13g2_nand3_1 _0984_ (.B(_0267_),
    .C(_0271_),
    .A(_0127_),
    .Y(_0349_));
 sg13g2_nand3_1 _0985_ (.B(_0264_),
    .C(_0295_),
    .A(_0256_),
    .Y(_0350_));
 sg13g2_a21oi_1 _0986_ (.A1(_0298_),
    .A2(_0350_),
    .Y(_0351_),
    .B1(_0274_));
 sg13g2_nand2b_1 _0987_ (.Y(_0352_),
    .B(net292),
    .A_N(_0351_));
 sg13g2_and3_1 _0988_ (.X(_0353_),
    .A(_0274_),
    .B(_0298_),
    .C(_0350_));
 sg13g2_o21ai_1 _0989_ (.B1(_0349_),
    .Y(_0354_),
    .A1(_0352_),
    .A2(_0353_));
 sg13g2_xnor2_1 _0990_ (.Y(_0355_),
    .A(net295),
    .B(_0354_));
 sg13g2_nand3b_1 _0991_ (.B(net292),
    .C(_0272_),
    .Y(_0356_),
    .A_N(_0351_));
 sg13g2_a21oi_1 _0992_ (.A1(net292),
    .A2(_0283_),
    .Y(_0357_),
    .B1(_0282_));
 sg13g2_xnor2_1 _0993_ (.Y(_0358_),
    .A(net295),
    .B(_0357_));
 sg13g2_xnor2_1 _0994_ (.Y(_0359_),
    .A(_0356_),
    .B(_0358_));
 sg13g2_nand3_1 _0995_ (.B(_0265_),
    .C(_0294_),
    .A(_0263_),
    .Y(_0360_));
 sg13g2_o21ai_1 _0996_ (.B1(net294),
    .Y(_0361_),
    .A1(_0263_),
    .A2(_0294_));
 sg13g2_nor2b_1 _0997_ (.A(_0361_),
    .B_N(_0350_),
    .Y(_0362_));
 sg13g2_a22oi_1 _0998_ (.Y(_0363_),
    .B1(_0360_),
    .B2(_0362_),
    .A2(_0291_),
    .A1(_0127_));
 sg13g2_xnor2_1 _0999_ (.Y(_0364_),
    .A(net295),
    .B(_0363_));
 sg13g2_xnor2_1 _1000_ (.Y(_0365_),
    .A(_0256_),
    .B(_0264_));
 sg13g2_mux2_1 _1001_ (.A0(_0263_),
    .A1(_0365_),
    .S(net292),
    .X(_0366_));
 sg13g2_xnor2_1 _1002_ (.Y(_0367_),
    .A(net295),
    .B(_0366_));
 sg13g2_nor2_1 _1003_ (.A(_0116_),
    .B(_0338_),
    .Y(_0368_));
 sg13g2_o21ai_1 _1004_ (.B1(net272),
    .Y(_0369_),
    .A1(\cpu.spi_mem_instance.count_s[2] ),
    .A2(_0359_));
 sg13g2_o21ai_1 _1005_ (.B1(net270),
    .Y(_0370_),
    .A1(_0368_),
    .A2(_0369_));
 sg13g2_a21oi_1 _1006_ (.A1(_0116_),
    .A2(_0355_),
    .Y(_0371_),
    .B1(net272));
 sg13g2_o21ai_1 _1007_ (.B1(_0371_),
    .Y(_0372_),
    .A1(_0116_),
    .A2(_0328_));
 sg13g2_nand2b_1 _1008_ (.Y(_0373_),
    .B(_0372_),
    .A_N(_0370_));
 sg13g2_mux4_1 _1009_ (.S0(_0116_),
    .A0(_0348_),
    .A1(_0367_),
    .A2(_0344_),
    .A3(_0364_),
    .S1(net272),
    .X(_0374_));
 sg13g2_o21ai_1 _1010_ (.B1(_0373_),
    .Y(_0375_),
    .A1(net270),
    .A2(_0374_));
 sg13g2_or2_1 _1011_ (.X(_0376_),
    .B(_0220_),
    .A(net293));
 sg13g2_nor2_1 _1012_ (.A(_0214_),
    .B(_0252_),
    .Y(_0377_));
 sg13g2_a21o_1 _1013_ (.A2(_0377_),
    .A1(_0243_),
    .B1(_0254_),
    .X(_0378_));
 sg13g2_xor2_1 _1014_ (.B(_0378_),
    .A(_0222_),
    .X(_0379_));
 sg13g2_o21ai_1 _1015_ (.B1(_0376_),
    .Y(_0380_),
    .A1(_0127_),
    .A2(_0379_));
 sg13g2_xnor2_1 _1016_ (.Y(_0381_),
    .A(net296),
    .B(_0380_));
 sg13g2_nand2b_1 _1017_ (.Y(_0382_),
    .B(net293),
    .A_N(_0220_));
 sg13g2_a21oi_1 _1018_ (.A1(_0222_),
    .A2(_0378_),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_a21oi_1 _1019_ (.A1(net293),
    .A2(_0231_),
    .Y(_0384_),
    .B1(_0230_));
 sg13g2_xnor2_1 _1020_ (.Y(_0385_),
    .A(net296),
    .B(_0384_));
 sg13g2_xnor2_1 _1021_ (.Y(_0386_),
    .A(_0383_),
    .B(_0385_));
 sg13g2_and2_1 _1022_ (.A(_0127_),
    .B(_0241_),
    .X(_0387_));
 sg13g2_o21ai_1 _1023_ (.B1(_0250_),
    .Y(_0388_),
    .A1(_0214_),
    .A2(_0252_));
 sg13g2_xnor2_1 _1024_ (.Y(_0389_),
    .A(_0243_),
    .B(_0388_));
 sg13g2_a21oi_1 _1025_ (.A1(net294),
    .A2(_0389_),
    .Y(_0390_),
    .B1(_0387_));
 sg13g2_xnor2_1 _1026_ (.Y(_0391_),
    .A(net296),
    .B(_0390_));
 sg13g2_nand2_1 _1027_ (.Y(_0392_),
    .A(_0214_),
    .B(_0252_));
 sg13g2_nand3b_1 _1028_ (.B(_0392_),
    .C(net293),
    .Y(_0393_),
    .A_N(_0377_));
 sg13g2_o21ai_1 _1029_ (.B1(_0393_),
    .Y(_0394_),
    .A1(net293),
    .A2(_0250_));
 sg13g2_xnor2_1 _1030_ (.Y(_0395_),
    .A(net296),
    .B(_0394_));
 sg13g2_o21ai_1 _1031_ (.B1(net271),
    .Y(_0396_),
    .A1(net273),
    .A2(_0381_));
 sg13g2_a21o_1 _1032_ (.A2(_0386_),
    .A1(net273),
    .B1(_0396_),
    .X(_0397_));
 sg13g2_nand2b_1 _1033_ (.Y(_0398_),
    .B(_0395_),
    .A_N(net273));
 sg13g2_a21oi_1 _1034_ (.A1(net273),
    .A2(_0391_),
    .Y(_0399_),
    .B1(net271));
 sg13g2_a21oi_1 _1035_ (.A1(_0398_),
    .A2(_0399_),
    .Y(_0400_),
    .B1(_0116_));
 sg13g2_a21oi_1 _1036_ (.A1(_0194_),
    .A2(_0202_),
    .Y(_0401_),
    .B1(_0127_));
 sg13g2_or2_1 _1037_ (.X(_0402_),
    .B(_0202_),
    .A(_0194_));
 sg13g2_a22oi_1 _1038_ (.Y(_0403_),
    .B1(_0401_),
    .B2(_0402_),
    .A2(_0200_),
    .A1(_0127_));
 sg13g2_xnor2_1 _1039_ (.Y(_0404_),
    .A(net296),
    .B(_0403_));
 sg13g2_nand2b_1 _1040_ (.Y(_0405_),
    .B(_0404_),
    .A_N(net273));
 sg13g2_nor2b_1 _1041_ (.A(\cpu.spi_mem_instance.count_s[2] ),
    .B_N(net271),
    .Y(_0406_));
 sg13g2_nand2b_1 _1042_ (.Y(_0407_),
    .B(_0401_),
    .A_N(_0200_));
 sg13g2_a21oi_1 _1043_ (.A1(net294),
    .A2(_0211_),
    .Y(_0408_),
    .B1(_0210_));
 sg13g2_xnor2_1 _1044_ (.Y(_0409_),
    .A(net296),
    .B(_0408_));
 sg13g2_xnor2_1 _1045_ (.Y(_0410_),
    .A(_0407_),
    .B(_0409_));
 sg13g2_nand2_1 _1046_ (.Y(_0411_),
    .A(net273),
    .B(_0410_));
 sg13g2_nand3_1 _1047_ (.B(_0406_),
    .C(_0411_),
    .A(_0405_),
    .Y(_0412_));
 sg13g2_xnor2_1 _1048_ (.Y(_0413_),
    .A(_0191_),
    .B(_0193_));
 sg13g2_nor2_1 _1049_ (.A(net293),
    .B(_0185_),
    .Y(_0414_));
 sg13g2_a21oi_1 _1050_ (.A1(net293),
    .A2(_0413_),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_xnor2_1 _1051_ (.Y(_0416_),
    .A(net296),
    .B(_0415_));
 sg13g2_nand2_1 _1052_ (.Y(_0417_),
    .A(net273),
    .B(_0416_));
 sg13g2_a21oi_1 _1053_ (.A1(_0189_),
    .A2(_0190_),
    .Y(_0418_),
    .B1(_0187_));
 sg13g2_nand2b_1 _1054_ (.Y(_0419_),
    .B(net293),
    .A_N(_0418_));
 sg13g2_xnor2_1 _1055_ (.Y(_0420_),
    .A(net296),
    .B(_0191_));
 sg13g2_xnor2_1 _1056_ (.Y(_0421_),
    .A(_0419_),
    .B(_0420_));
 sg13g2_nand2b_1 _1057_ (.Y(_0422_),
    .B(_0421_),
    .A_N(net273));
 sg13g2_nand3_1 _1058_ (.B(_0417_),
    .C(_0422_),
    .A(_0140_),
    .Y(_0423_));
 sg13g2_nand3_1 _1059_ (.B(_0412_),
    .C(_0423_),
    .A(\cpu.spi_mem_instance.count_s[3] ),
    .Y(_0424_));
 sg13g2_a21oi_1 _1060_ (.A1(_0397_),
    .A2(_0400_),
    .Y(_0425_),
    .B1(_0424_));
 sg13g2_nor3_1 _1061_ (.A(\cpu.spi_mem_instance.count_s[5] ),
    .B(\cpu.spi_mem_instance.count_s[4] ),
    .C(_0425_),
    .Y(_0426_));
 sg13g2_o21ai_1 _1062_ (.B1(_0426_),
    .Y(_0427_),
    .A1(\cpu.spi_mem_instance.count_s[3] ),
    .A2(_0375_));
 sg13g2_nand2_1 _1063_ (.Y(_0428_),
    .A(\cpu.fsm_instance.state_s[0] ),
    .B(_0007_));
 sg13g2_nand4_1 _1064_ (.B(_0006_),
    .C(_0144_),
    .A(\cpu.spi_mem_instance.count_s[5] ),
    .Y(_0429_),
    .D(_0428_));
 sg13g2_mux4_1 _1065_ (.S0(net274),
    .A0(\cpu.pc_s[4] ),
    .A1(\cpu.pc_s[5] ),
    .A2(\cpu.regA_s[4] ),
    .A3(\cpu.regA_s[5] ),
    .S1(net315),
    .X(_0430_));
 sg13g2_nor2_1 _1066_ (.A(net271),
    .B(_0430_),
    .Y(_0431_));
 sg13g2_nor2b_1 _1067_ (.A(\cpu.regA_s[6] ),
    .B_N(net315),
    .Y(_0432_));
 sg13g2_nor2_1 _1068_ (.A(net316),
    .B(\cpu.pc_s[6] ),
    .Y(_0433_));
 sg13g2_nor3_1 _1069_ (.A(net274),
    .B(_0432_),
    .C(_0433_),
    .Y(_0434_));
 sg13g2_nor2b_1 _1070_ (.A(\cpu.regA_s[7] ),
    .B_N(net315),
    .Y(_0435_));
 sg13g2_o21ai_1 _1071_ (.B1(net274),
    .Y(_0436_),
    .A1(net315),
    .A2(\cpu.pc_s[7] ));
 sg13g2_o21ai_1 _1072_ (.B1(net270),
    .Y(_0437_),
    .A1(_0435_),
    .A2(_0436_));
 sg13g2_o21ai_1 _1073_ (.B1(\cpu.spi_mem_instance.count_s[2] ),
    .Y(_0438_),
    .A1(_0434_),
    .A2(_0437_));
 sg13g2_mux4_1 _1074_ (.S0(net274),
    .A0(\cpu.pc_s[0] ),
    .A1(\cpu.pc_s[1] ),
    .A2(\cpu.regA_s[0] ),
    .A3(\cpu.regA_s[1] ),
    .S1(net315),
    .X(_0439_));
 sg13g2_mux4_1 _1075_ (.S0(net274),
    .A0(\cpu.pc_s[2] ),
    .A1(\cpu.pc_s[3] ),
    .A2(\cpu.regA_s[2] ),
    .A3(\cpu.regA_s[3] ),
    .S1(net315),
    .X(_0440_));
 sg13g2_a221oi_1 _1076_ (.B2(_0406_),
    .C1(\cpu.spi_mem_instance.count_s[3] ),
    .B1(_0440_),
    .A1(_0140_),
    .Y(_0441_),
    .A2(_0439_));
 sg13g2_o21ai_1 _1077_ (.B1(_0441_),
    .Y(_0442_),
    .A1(_0431_),
    .A2(_0438_));
 sg13g2_mux4_1 _1078_ (.S0(net272),
    .A0(\cpu.pc_s[12] ),
    .A1(\cpu.pc_s[13] ),
    .A2(\cpu.regA_s[12] ),
    .A3(\cpu.regA_s[13] ),
    .S1(net313),
    .X(_0443_));
 sg13g2_nor2b_1 _1079_ (.A(\cpu.regA_s[14] ),
    .B_N(net314),
    .Y(_0444_));
 sg13g2_nor2_1 _1080_ (.A(net314),
    .B(\cpu.pc_s[14] ),
    .Y(_0445_));
 sg13g2_nor3_1 _1081_ (.A(net272),
    .B(_0444_),
    .C(_0445_),
    .Y(_0446_));
 sg13g2_nor2b_1 _1082_ (.A(\cpu.regA_s[15] ),
    .B_N(net314),
    .Y(_0447_));
 sg13g2_o21ai_1 _1083_ (.B1(net272),
    .Y(_0448_),
    .A1(net314),
    .A2(\cpu.pc_s[15] ));
 sg13g2_o21ai_1 _1084_ (.B1(net270),
    .Y(_0449_),
    .A1(_0447_),
    .A2(_0448_));
 sg13g2_o21ai_1 _1085_ (.B1(\cpu.spi_mem_instance.count_s[2] ),
    .Y(_0450_),
    .A1(_0446_),
    .A2(_0449_));
 sg13g2_inv_1 _1086_ (.Y(_0451_),
    .A(_0450_));
 sg13g2_o21ai_1 _1087_ (.B1(_0451_),
    .Y(_0452_),
    .A1(net270),
    .A2(_0443_));
 sg13g2_mux4_1 _1088_ (.S0(net274),
    .A0(\cpu.pc_s[8] ),
    .A1(\cpu.pc_s[9] ),
    .A2(\cpu.regA_s[8] ),
    .A3(\cpu.regA_s[9] ),
    .S1(net315),
    .X(_0453_));
 sg13g2_mux4_1 _1089_ (.S0(net272),
    .A0(\cpu.pc_s[10] ),
    .A1(\cpu.pc_s[11] ),
    .A2(\cpu.regA_s[10] ),
    .A3(\cpu.regA_s[11] ),
    .S1(net316),
    .X(_0454_));
 sg13g2_a22oi_1 _1090_ (.Y(_0455_),
    .B1(_0454_),
    .B2(_0406_),
    .A2(_0453_),
    .A1(_0140_));
 sg13g2_nand3_1 _1091_ (.B(_0452_),
    .C(_0455_),
    .A(\cpu.spi_mem_instance.count_s[3] ),
    .Y(_0456_));
 sg13g2_nand4_1 _1092_ (.B(\cpu.spi_mem_instance.count_s[4] ),
    .C(_0442_),
    .A(_0115_),
    .Y(_0457_),
    .D(_0456_));
 sg13g2_nand3_1 _1093_ (.B(_0429_),
    .C(_0457_),
    .A(_0427_),
    .Y(\cpu.mem_out_o ));
 sg13g2_nor2b_1 _1094_ (.A(\cpu.spi_debug_instance.in_s[1] ),
    .B_N(\cpu.spi_debug_instance.in_s[0] ),
    .Y(_0458_));
 sg13g2_nor2_1 _1095_ (.A(\cpu.spi_debug_instance.in_s[0] ),
    .B(\cpu.spi_debug_instance.in_s[1] ),
    .Y(_0459_));
 sg13g2_nor2b_1 _1096_ (.A(\cpu.spi_debug_instance.in_s[0] ),
    .B_N(\cpu.spi_debug_instance.in_s[1] ),
    .Y(_0460_));
 sg13g2_a21oi_1 _1097_ (.A1(\cpu.alu_instance.a_i[6] ),
    .A2(net279),
    .Y(_0461_),
    .B1(\cpu.spi_debug_instance.counter_s[0] ));
 sg13g2_a22oi_1 _1098_ (.Y(_0462_),
    .B1(net278),
    .B2(\cpu.pc_s[6] ),
    .A2(net281),
    .A1(\cpu.regA_s[6] ));
 sg13g2_a21oi_1 _1099_ (.A1(\cpu.pc_s[7] ),
    .A2(net277),
    .Y(_0463_),
    .B1(_0118_));
 sg13g2_a22oi_1 _1100_ (.Y(_0464_),
    .B1(net279),
    .B2(\cpu.alu_instance.a_i[7] ),
    .A2(_0458_),
    .A1(\cpu.regA_s[7] ));
 sg13g2_a221oi_1 _1101_ (.B2(_0464_),
    .C1(_0117_),
    .B1(_0463_),
    .A1(_0461_),
    .Y(_0465_),
    .A2(_0462_));
 sg13g2_nand2_1 _1102_ (.Y(_0466_),
    .A(_0117_),
    .B(\cpu.spi_debug_instance.counter_s[0] ));
 sg13g2_nand2_1 _1103_ (.Y(_0467_),
    .A(\cpu.alu_instance.a_i[5] ),
    .B(net279));
 sg13g2_a22oi_1 _1104_ (.Y(_0468_),
    .B1(net277),
    .B2(\cpu.pc_s[5] ),
    .A2(net281),
    .A1(\cpu.regA_s[5] ));
 sg13g2_a21oi_1 _1105_ (.A1(_0467_),
    .A2(_0468_),
    .Y(_0469_),
    .B1(_0466_));
 sg13g2_nand2_1 _1106_ (.Y(_0470_),
    .A(\cpu.alu_instance.a_i[4] ),
    .B(net279));
 sg13g2_a22oi_1 _1107_ (.Y(_0471_),
    .B1(net277),
    .B2(\cpu.pc_s[4] ),
    .A2(net281),
    .A1(\cpu.regA_s[4] ));
 sg13g2_a21oi_1 _1108_ (.A1(_0470_),
    .A2(_0471_),
    .Y(_0472_),
    .B1(_0154_));
 sg13g2_nor4_1 _1109_ (.A(net276),
    .B(_0465_),
    .C(_0469_),
    .D(_0472_),
    .Y(_0473_));
 sg13g2_a21oi_1 _1110_ (.A1(\cpu.pc_s[14] ),
    .A2(net278),
    .Y(_0474_),
    .B1(\cpu.spi_debug_instance.counter_s[0] ));
 sg13g2_a22oi_1 _1111_ (.Y(_0475_),
    .B1(net280),
    .B2(\cpu.alu_instance.a_i[14] ),
    .A2(net282),
    .A1(\cpu.regA_s[14] ));
 sg13g2_a21oi_1 _1112_ (.A1(\cpu.alu_instance.a_i[15] ),
    .A2(net280),
    .Y(_0476_),
    .B1(_0118_));
 sg13g2_a22oi_1 _1113_ (.Y(_0477_),
    .B1(net278),
    .B2(\cpu.pc_s[15] ),
    .A2(net282),
    .A1(\cpu.regA_s[15] ));
 sg13g2_a22oi_1 _1114_ (.Y(_0478_),
    .B1(_0476_),
    .B2(_0477_),
    .A2(_0475_),
    .A1(_0474_));
 sg13g2_and2_1 _1115_ (.A(\cpu.regA_s[12] ),
    .B(net282),
    .X(_0479_));
 sg13g2_a221oi_1 _1116_ (.B2(\cpu.pc_s[12] ),
    .C1(_0479_),
    .B1(net278),
    .A1(\cpu.alu_instance.a_i[12] ),
    .Y(_0480_),
    .A2(net280));
 sg13g2_nand2_1 _1117_ (.Y(_0481_),
    .A(\cpu.regA_s[13] ),
    .B(net282));
 sg13g2_a22oi_1 _1118_ (.Y(_0482_),
    .B1(net278),
    .B2(\cpu.pc_s[13] ),
    .A2(net280),
    .A1(\cpu.alu_instance.a_i[13] ));
 sg13g2_a21oi_1 _1119_ (.A1(_0481_),
    .A2(_0482_),
    .Y(_0483_),
    .B1(_0466_));
 sg13g2_o21ai_1 _1120_ (.B1(net276),
    .Y(_0484_),
    .A1(_0154_),
    .A2(_0480_));
 sg13g2_a21o_1 _1121_ (.A2(_0478_),
    .A1(\cpu.spi_debug_instance.counter_s[1] ),
    .B1(_0484_),
    .X(_0485_));
 sg13g2_o21ai_1 _1122_ (.B1(\cpu.spi_debug_instance.counter_s[2] ),
    .Y(_0486_),
    .A1(_0483_),
    .A2(_0485_));
 sg13g2_a22oi_1 _1123_ (.Y(_0487_),
    .B1(net277),
    .B2(\cpu.pc_s[3] ),
    .A2(net282),
    .A1(\cpu.regA_s[3] ));
 sg13g2_a21oi_1 _1124_ (.A1(\cpu.alu_instance.a_i[3] ),
    .A2(net279),
    .Y(_0488_),
    .B1(_0118_));
 sg13g2_a22oi_1 _1125_ (.Y(_0489_),
    .B1(net279),
    .B2(\cpu.alu_instance.a_i[2] ),
    .A2(net281),
    .A1(\cpu.regA_s[2] ));
 sg13g2_a21oi_1 _1126_ (.A1(\cpu.pc_s[2] ),
    .A2(net277),
    .Y(_0490_),
    .B1(\cpu.spi_debug_instance.counter_s[0] ));
 sg13g2_and2_1 _1127_ (.A(\cpu.spi_debug_instance.in_s[0] ),
    .B(\cpu.spi_debug_instance.in_s[1] ),
    .X(_0491_));
 sg13g2_nand2_1 _1128_ (.Y(_0492_),
    .A(\cpu.alu_instance.a_i[0] ),
    .B(net280));
 sg13g2_nand2_1 _1129_ (.Y(_0493_),
    .A(\cpu.fsm_instance.state_s[0] ),
    .B(_0491_));
 sg13g2_a21oi_1 _1130_ (.A1(\cpu.regA_s[11] ),
    .A2(net282),
    .Y(_0494_),
    .B1(_0118_));
 sg13g2_a22oi_1 _1131_ (.Y(_0495_),
    .B1(net278),
    .B2(\cpu.pc_s[11] ),
    .A2(net280),
    .A1(\cpu.alu_instance.a_i[11] ));
 sg13g2_a21oi_1 _1132_ (.A1(\cpu.alu_instance.a_i[10] ),
    .A2(net280),
    .Y(_0496_),
    .B1(\cpu.spi_debug_instance.counter_s[0] ));
 sg13g2_a22oi_1 _1133_ (.Y(_0497_),
    .B1(net278),
    .B2(\cpu.pc_s[10] ),
    .A2(net282),
    .A1(\cpu.regA_s[10] ));
 sg13g2_a22oi_1 _1134_ (.Y(_0498_),
    .B1(_0496_),
    .B2(_0497_),
    .A2(_0495_),
    .A1(_0494_));
 sg13g2_nand2_1 _1135_ (.Y(_0499_),
    .A(\cpu.regA_s[8] ),
    .B(net281));
 sg13g2_a22oi_1 _1136_ (.Y(_0500_),
    .B1(net277),
    .B2(\cpu.pc_s[8] ),
    .A2(net279),
    .A1(\cpu.alu_instance.a_i[8] ));
 sg13g2_a21o_1 _1137_ (.A2(_0500_),
    .A1(_0499_),
    .B1(_0154_),
    .X(_0501_));
 sg13g2_and2_1 _1138_ (.A(\cpu.pc_s[9] ),
    .B(net277),
    .X(_0502_));
 sg13g2_a221oi_1 _1139_ (.B2(\cpu.alu_instance.a_i[9] ),
    .C1(_0502_),
    .B1(net279),
    .A1(\cpu.regA_s[9] ),
    .Y(_0503_),
    .A2(net281));
 sg13g2_a22oi_1 _1140_ (.Y(_0504_),
    .B1(net277),
    .B2(\cpu.pc_s[0] ),
    .A2(net281),
    .A1(\cpu.regA_s[0] ));
 sg13g2_nand4_1 _1141_ (.B(_0492_),
    .C(_0493_),
    .A(_0118_),
    .Y(_0505_),
    .D(_0504_));
 sg13g2_a22oi_1 _1142_ (.Y(_0506_),
    .B1(_0460_),
    .B2(\cpu.pc_s[1] ),
    .A2(_0459_),
    .A1(\cpu.alu_instance.a_i[1] ));
 sg13g2_a221oi_1 _1143_ (.B2(net315),
    .C1(_0118_),
    .B1(_0491_),
    .A1(\cpu.regA_s[1] ),
    .Y(_0507_),
    .A2(net281));
 sg13g2_a21oi_1 _1144_ (.A1(_0506_),
    .A2(_0507_),
    .Y(_0508_),
    .B1(\cpu.spi_debug_instance.counter_s[1] ));
 sg13g2_a221oi_1 _1145_ (.B2(_0490_),
    .C1(_0117_),
    .B1(_0489_),
    .A1(_0487_),
    .Y(_0509_),
    .A2(_0488_));
 sg13g2_a21o_1 _1146_ (.A2(_0508_),
    .A1(_0505_),
    .B1(_0509_),
    .X(_0510_));
 sg13g2_o21ai_1 _1147_ (.B1(net276),
    .Y(_0511_),
    .A1(_0466_),
    .A2(_0503_));
 sg13g2_a21oi_1 _1148_ (.A1(\cpu.spi_debug_instance.counter_s[1] ),
    .A2(_0498_),
    .Y(_0512_),
    .B1(_0511_));
 sg13g2_a21oi_1 _1149_ (.A1(_0501_),
    .A2(_0512_),
    .Y(_0513_),
    .B1(\cpu.spi_debug_instance.counter_s[2] ));
 sg13g2_o21ai_1 _1150_ (.B1(_0513_),
    .Y(_0514_),
    .A1(net276),
    .A2(_0510_));
 sg13g2_o21ai_1 _1151_ (.B1(_0514_),
    .Y(\cpu.debug_out_o ),
    .A1(_0473_),
    .A2(_0486_));
 sg13g2_nand2_1 _1152_ (.Y(\cpu.mem_sclk_o ),
    .A(net27),
    .B(_0139_));
 sg13g2_and3_1 _1153_ (.X(_0515_),
    .A(net307),
    .B(\cpu.fsm_instance.instruction_i[4] ),
    .C(_0170_));
 sg13g2_nor2_1 _1154_ (.A(net64),
    .B(net268),
    .Y(_0516_));
 sg13g2_a21oi_1 _1155_ (.A1(_0421_),
    .A2(net268),
    .Y(_0020_),
    .B1(_0516_));
 sg13g2_nor2_1 _1156_ (.A(net57),
    .B(net268),
    .Y(_0517_));
 sg13g2_a21oi_1 _1157_ (.A1(_0416_),
    .A2(net269),
    .Y(_0021_),
    .B1(_0517_));
 sg13g2_nor2_1 _1158_ (.A(net84),
    .B(net268),
    .Y(_0518_));
 sg13g2_a21oi_1 _1159_ (.A1(_0404_),
    .A2(net268),
    .Y(_0022_),
    .B1(_0518_));
 sg13g2_nor2_1 _1160_ (.A(net91),
    .B(net268),
    .Y(_0519_));
 sg13g2_a21oi_1 _1161_ (.A1(_0410_),
    .A2(net268),
    .Y(_0023_),
    .B1(_0519_));
 sg13g2_mux2_1 _1162_ (.A0(net78),
    .A1(_0395_),
    .S(net268),
    .X(_0024_));
 sg13g2_mux2_1 _1163_ (.A0(net56),
    .A1(_0391_),
    .S(net269),
    .X(_0025_));
 sg13g2_nor2_1 _1164_ (.A(net77),
    .B(net269),
    .Y(_0520_));
 sg13g2_a21oi_1 _1165_ (.A1(_0381_),
    .A2(net269),
    .Y(_0026_),
    .B1(_0520_));
 sg13g2_mux2_1 _1166_ (.A0(net88),
    .A1(_0386_),
    .S(net269),
    .X(_0027_));
 sg13g2_nor2_1 _1167_ (.A(net52),
    .B(net267),
    .Y(_0521_));
 sg13g2_a21oi_1 _1168_ (.A1(_0367_),
    .A2(net267),
    .Y(_0028_),
    .B1(_0521_));
 sg13g2_nor2_1 _1169_ (.A(net55),
    .B(net267),
    .Y(_0522_));
 sg13g2_a21oi_1 _1170_ (.A1(_0364_),
    .A2(net267),
    .Y(_0029_),
    .B1(_0522_));
 sg13g2_mux2_1 _1171_ (.A0(net89),
    .A1(_0355_),
    .S(net266),
    .X(_0030_));
 sg13g2_nor2_1 _1172_ (.A(net86),
    .B(net267),
    .Y(_0523_));
 sg13g2_a21oi_1 _1173_ (.A1(_0359_),
    .A2(net267),
    .Y(_0031_),
    .B1(_0523_));
 sg13g2_nor2_1 _1174_ (.A(net87),
    .B(net267),
    .Y(_0524_));
 sg13g2_a21oi_1 _1175_ (.A1(_0348_),
    .A2(net266),
    .Y(_0032_),
    .B1(_0524_));
 sg13g2_nor2_1 _1176_ (.A(net69),
    .B(net266),
    .Y(_0525_));
 sg13g2_a21oi_1 _1177_ (.A1(_0344_),
    .A2(net266),
    .Y(_0033_),
    .B1(_0525_));
 sg13g2_nor2_1 _1178_ (.A(net90),
    .B(net266),
    .Y(_0526_));
 sg13g2_a21oi_1 _1179_ (.A1(_0328_),
    .A2(net266),
    .Y(_0034_),
    .B1(_0526_));
 sg13g2_nor2_1 _1180_ (.A(net65),
    .B(net266),
    .Y(_0527_));
 sg13g2_a21oi_1 _1181_ (.A1(_0338_),
    .A2(net266),
    .Y(_0035_),
    .B1(_0527_));
 sg13g2_nand2_1 _1182_ (.Y(_0528_),
    .A(net66),
    .B(_0170_));
 sg13g2_o21ai_1 _1183_ (.B1(_0170_),
    .Y(_0529_),
    .A1(_0120_),
    .A2(\cpu.fsm_instance.instruction_i[5] ));
 sg13g2_o21ai_1 _1184_ (.B1(_0528_),
    .Y(_0530_),
    .A1(net307),
    .A2(_0171_));
 sg13g2_o21ai_1 _1185_ (.B1(net262),
    .Y(_0531_),
    .A1(net306),
    .A2(\cpu.fsm_instance.instruction_i[0] ));
 sg13g2_a21oi_1 _1186_ (.A1(net308),
    .A2(_0421_),
    .Y(_0532_),
    .B1(_0531_));
 sg13g2_a21o_1 _1187_ (.A2(net264),
    .A1(net110),
    .B1(_0532_),
    .X(_0036_));
 sg13g2_o21ai_1 _1188_ (.B1(net262),
    .Y(_0533_),
    .A1(net310),
    .A2(\cpu.fsm_instance.instruction_i[1] ));
 sg13g2_a21oi_1 _1189_ (.A1(net309),
    .A2(_0416_),
    .Y(_0534_),
    .B1(_0533_));
 sg13g2_a21o_1 _1190_ (.A2(net264),
    .A1(net131),
    .B1(_0534_),
    .X(_0037_));
 sg13g2_o21ai_1 _1191_ (.B1(net262),
    .Y(_0535_),
    .A1(net310),
    .A2(net59));
 sg13g2_a21oi_1 _1192_ (.A1(net309),
    .A2(_0404_),
    .Y(_0536_),
    .B1(_0535_));
 sg13g2_a21o_1 _1193_ (.A2(net264),
    .A1(net118),
    .B1(_0536_),
    .X(_0038_));
 sg13g2_o21ai_1 _1194_ (.B1(net262),
    .Y(_0537_),
    .A1(net307),
    .A2(\cpu.fsm_instance.instruction_i[3] ));
 sg13g2_a21oi_1 _1195_ (.A1(net309),
    .A2(_0410_),
    .Y(_0538_),
    .B1(_0537_));
 sg13g2_a21o_1 _1196_ (.A2(_0529_),
    .A1(net125),
    .B1(_0538_),
    .X(_0039_));
 sg13g2_nand2_1 _1197_ (.Y(_0539_),
    .A(net103),
    .B(_0529_));
 sg13g2_or2_1 _1198_ (.X(_0540_),
    .B(net94),
    .A(net307));
 sg13g2_o21ai_1 _1199_ (.B1(_0540_),
    .Y(_0541_),
    .A1(_0120_),
    .A2(_0395_));
 sg13g2_o21ai_1 _1200_ (.B1(net104),
    .Y(_0040_),
    .A1(net264),
    .A2(_0541_));
 sg13g2_nand2_1 _1201_ (.Y(_0542_),
    .A(net97),
    .B(net264));
 sg13g2_nor2_1 _1202_ (.A(_0120_),
    .B(_0391_),
    .Y(_0543_));
 sg13g2_o21ai_1 _1203_ (.B1(_0542_),
    .Y(_0041_),
    .A1(_0528_),
    .A2(_0543_));
 sg13g2_o21ai_1 _1204_ (.B1(net263),
    .Y(_0544_),
    .A1(net307),
    .A2(net41));
 sg13g2_a21oi_1 _1205_ (.A1(net309),
    .A2(_0381_),
    .Y(_0545_),
    .B1(_0544_));
 sg13g2_a21o_1 _1206_ (.A2(_0529_),
    .A1(net120),
    .B1(_0545_),
    .X(_0042_));
 sg13g2_nand2_1 _1207_ (.Y(_0546_),
    .A(net102),
    .B(net264));
 sg13g2_nor2_1 _1208_ (.A(_0120_),
    .B(_0386_),
    .Y(_0547_));
 sg13g2_o21ai_1 _1209_ (.B1(net263),
    .Y(_0548_),
    .A1(net308),
    .A2(net292));
 sg13g2_o21ai_1 _1210_ (.B1(_0546_),
    .Y(_0043_),
    .A1(_0547_),
    .A2(_0548_));
 sg13g2_o21ai_1 _1211_ (.B1(net263),
    .Y(_0549_),
    .A1(net308),
    .A2(net48));
 sg13g2_a21oi_1 _1212_ (.A1(net308),
    .A2(_0367_),
    .Y(_0550_),
    .B1(_0549_));
 sg13g2_a21o_1 _1213_ (.A2(net264),
    .A1(net127),
    .B1(_0550_),
    .X(_0044_));
 sg13g2_o21ai_1 _1214_ (.B1(net263),
    .Y(_0551_),
    .A1(net308),
    .A2(\cpu.alu_instance.zb_i ));
 sg13g2_a21oi_1 _1215_ (.A1(net308),
    .A2(_0364_),
    .Y(_0552_),
    .B1(_0551_));
 sg13g2_a21o_1 _1216_ (.A2(net264),
    .A1(net116),
    .B1(_0552_),
    .X(_0045_));
 sg13g2_nand2_1 _1217_ (.Y(_0553_),
    .A(net96),
    .B(net265));
 sg13g2_nor2_1 _1218_ (.A(_0120_),
    .B(_0355_),
    .Y(_0554_));
 sg13g2_o21ai_1 _1219_ (.B1(net262),
    .Y(_0555_),
    .A1(net307),
    .A2(net70));
 sg13g2_o21ai_1 _1220_ (.B1(_0553_),
    .Y(_0046_),
    .A1(_0554_),
    .A2(_0555_));
 sg13g2_o21ai_1 _1221_ (.B1(net263),
    .Y(_0556_),
    .A1(net308),
    .A2(net299));
 sg13g2_a21oi_1 _1222_ (.A1(net308),
    .A2(_0359_),
    .Y(_0557_),
    .B1(_0556_));
 sg13g2_a21o_1 _1223_ (.A2(net265),
    .A1(net105),
    .B1(_0557_),
    .X(_0047_));
 sg13g2_o21ai_1 _1224_ (.B1(net262),
    .Y(_0558_),
    .A1(net306),
    .A2(net303));
 sg13g2_a21oi_1 _1225_ (.A1(net306),
    .A2(_0348_),
    .Y(_0559_),
    .B1(_0558_));
 sg13g2_a21o_1 _1226_ (.A2(net265),
    .A1(net121),
    .B1(_0559_),
    .X(_0048_));
 sg13g2_o21ai_1 _1227_ (.B1(net262),
    .Y(_0560_),
    .A1(net306),
    .A2(net58));
 sg13g2_a21oi_1 _1228_ (.A1(net306),
    .A2(_0344_),
    .Y(_0561_),
    .B1(_0560_));
 sg13g2_a21o_1 _1229_ (.A2(net265),
    .A1(net134),
    .B1(_0561_),
    .X(_0049_));
 sg13g2_o21ai_1 _1230_ (.B1(net262),
    .Y(_0562_),
    .A1(net306),
    .A2(net38));
 sg13g2_a21oi_1 _1231_ (.A1(net306),
    .A2(_0328_),
    .Y(_0563_),
    .B1(_0562_));
 sg13g2_a21o_1 _1232_ (.A2(net265),
    .A1(net117),
    .B1(_0563_),
    .X(_0050_));
 sg13g2_nor3_1 _1233_ (.A(net50),
    .B(_0338_),
    .C(net265),
    .Y(_0564_));
 sg13g2_a21o_1 _1234_ (.A2(net265),
    .A1(\cpu.regA_s[15] ),
    .B1(_0564_),
    .X(_0051_));
 sg13g2_nor3_1 _1235_ (.A(net1),
    .B(_0135_),
    .C(_0138_),
    .Y(_0565_));
 sg13g2_nor3_2 _1236_ (.A(net1),
    .B(_0139_),
    .C(_0171_),
    .Y(_0566_));
 sg13g2_nand3b_1 _1237_ (.B(\cpu.mem_csb_o ),
    .C(_0170_),
    .Y(_0567_),
    .A_N(net1));
 sg13g2_nand2b_1 _1238_ (.Y(_0568_),
    .B(net252),
    .A_N(_0565_));
 sg13g2_nor2_1 _1239_ (.A(net317),
    .B(_0565_),
    .Y(_0569_));
 sg13g2_a21oi_1 _1240_ (.A1(net307),
    .A2(net302),
    .Y(_0570_),
    .B1(net317));
 sg13g2_nor2_1 _1241_ (.A(net313),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_a21oi_1 _1242_ (.A1(_0568_),
    .A2(_0571_),
    .Y(_0057_),
    .B1(_0569_));
 sg13g2_nor2b_1 _1243_ (.A(net317),
    .B_N(net313),
    .Y(_0572_));
 sg13g2_nor2_1 _1244_ (.A(net303),
    .B(\cpu.fsm_instance.instruction_i[3] ),
    .Y(_0573_));
 sg13g2_nor4_1 _1245_ (.A(net317),
    .B(net313),
    .C(_0120_),
    .D(_0573_),
    .Y(_0574_));
 sg13g2_a21o_1 _1246_ (.A2(_0572_),
    .A1(net76),
    .B1(_0574_),
    .X(_0575_));
 sg13g2_mux2_1 _1247_ (.A0(net313),
    .A1(_0575_),
    .S(_0568_),
    .X(_0058_));
 sg13g2_nand4_1 _1248_ (.B(_0410_),
    .C(_0416_),
    .A(_0404_),
    .Y(_0576_),
    .D(_0421_));
 sg13g2_nor4_1 _1249_ (.A(_0386_),
    .B(_0391_),
    .C(_0395_),
    .D(_0576_),
    .Y(_0577_));
 sg13g2_and4_1 _1250_ (.A(_0344_),
    .B(_0348_),
    .C(_0367_),
    .D(_0577_),
    .X(_0578_));
 sg13g2_nand3_1 _1251_ (.B(_0364_),
    .C(_0381_),
    .A(_0359_),
    .Y(_0579_));
 sg13g2_nor2_1 _1252_ (.A(_0355_),
    .B(_0579_),
    .Y(_0580_));
 sg13g2_nand4_1 _1253_ (.B(_0338_),
    .C(_0578_),
    .A(_0328_),
    .Y(_0581_),
    .D(_0580_));
 sg13g2_nand2_1 _1254_ (.Y(_0582_),
    .A(\cpu.fsm_instance.instruction_i[0] ),
    .B(_0338_));
 sg13g2_or2_1 _1255_ (.X(_0583_),
    .B(_0338_),
    .A(_0128_));
 sg13g2_mux2_1 _1256_ (.A0(_0129_),
    .A1(_0582_),
    .S(_0581_),
    .X(_0584_));
 sg13g2_nand2b_1 _1257_ (.Y(_0585_),
    .B(_0170_),
    .A_N(net50));
 sg13g2_a21oi_2 _1258_ (.B1(_0585_),
    .Y(_0586_),
    .A2(_0584_),
    .A1(_0583_));
 sg13g2_nand2_2 _1259_ (.Y(_0587_),
    .A(_0566_),
    .B(net251));
 sg13g2_mux2_1 _1260_ (.A0(\cpu.regA_s[0] ),
    .A1(net92),
    .S(_0587_),
    .X(_0059_));
 sg13g2_mux2_1 _1261_ (.A0(_0005_),
    .A1(\cpu.regA_s[1] ),
    .S(net251),
    .X(_0588_));
 sg13g2_mux2_1 _1262_ (.A0(net100),
    .A1(_0588_),
    .S(_0566_),
    .X(_0060_));
 sg13g2_nand2_1 _1263_ (.Y(_0589_),
    .A(\cpu.pc_s[1] ),
    .B(\cpu.pc_s[2] ));
 sg13g2_nor2_2 _1264_ (.A(_0567_),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_a21oi_1 _1265_ (.A1(net100),
    .A2(_0566_),
    .Y(_0591_),
    .B1(net129));
 sg13g2_nor2_1 _1266_ (.A(_0590_),
    .B(_0591_),
    .Y(_0592_));
 sg13g2_mux2_1 _1267_ (.A0(net118),
    .A1(_0592_),
    .S(_0587_),
    .X(_0061_));
 sg13g2_xor2_1 _1268_ (.B(_0590_),
    .A(\cpu.pc_s[3] ),
    .X(_0593_));
 sg13g2_mux2_1 _1269_ (.A0(net125),
    .A1(_0593_),
    .S(_0587_),
    .X(_0062_));
 sg13g2_nand3_1 _1270_ (.B(\cpu.pc_s[4] ),
    .C(_0590_),
    .A(\cpu.pc_s[3] ),
    .Y(_0594_));
 sg13g2_a21o_1 _1271_ (.A2(_0590_),
    .A1(\cpu.pc_s[3] ),
    .B1(\cpu.pc_s[4] ),
    .X(_0595_));
 sg13g2_and2_1 _1272_ (.A(_0594_),
    .B(_0595_),
    .X(_0596_));
 sg13g2_mux2_1 _1273_ (.A0(net103),
    .A1(_0596_),
    .S(net250),
    .X(_0063_));
 sg13g2_nand3_1 _1274_ (.B(\cpu.pc_s[4] ),
    .C(\cpu.pc_s[5] ),
    .A(\cpu.pc_s[3] ),
    .Y(_0597_));
 sg13g2_nor2_2 _1275_ (.A(_0589_),
    .B(_0597_),
    .Y(_0598_));
 sg13g2_xnor2_1 _1276_ (.Y(_0599_),
    .A(net130),
    .B(_0594_));
 sg13g2_mux2_1 _1277_ (.A0(net97),
    .A1(_0599_),
    .S(net250),
    .X(_0064_));
 sg13g2_xnor2_1 _1278_ (.Y(_0600_),
    .A(_0130_),
    .B(_0598_));
 sg13g2_nand2b_1 _1279_ (.Y(_0601_),
    .B(_0600_),
    .A_N(_0586_));
 sg13g2_a21oi_1 _1280_ (.A1(net120),
    .A2(net251),
    .Y(_0602_),
    .B1(_0567_));
 sg13g2_a22oi_1 _1281_ (.Y(_0065_),
    .B1(_0601_),
    .B2(_0602_),
    .A2(net252),
    .A1(_0130_));
 sg13g2_nand3_1 _1282_ (.B(_0566_),
    .C(_0598_),
    .A(\cpu.pc_s[6] ),
    .Y(_0603_));
 sg13g2_xnor2_1 _1283_ (.Y(_0604_),
    .A(net136),
    .B(_0603_));
 sg13g2_mux2_1 _1284_ (.A0(net102),
    .A1(net137),
    .S(net250),
    .X(_0066_));
 sg13g2_nand3_1 _1285_ (.B(\cpu.pc_s[7] ),
    .C(_0598_),
    .A(\cpu.pc_s[6] ),
    .Y(_0605_));
 sg13g2_nor2_1 _1286_ (.A(_0131_),
    .B(_0605_),
    .Y(_0606_));
 sg13g2_xnor2_1 _1287_ (.Y(_0607_),
    .A(net140),
    .B(_0605_));
 sg13g2_nand2b_1 _1288_ (.Y(_0608_),
    .B(_0607_),
    .A_N(net251));
 sg13g2_a21oi_1 _1289_ (.A1(net127),
    .A2(_0586_),
    .Y(_0609_),
    .B1(net252));
 sg13g2_a22oi_1 _1290_ (.Y(_0067_),
    .B1(_0608_),
    .B2(_0609_),
    .A2(net252),
    .A1(_0131_));
 sg13g2_nor3_2 _1291_ (.A(_0131_),
    .B(_0132_),
    .C(_0605_),
    .Y(_0610_));
 sg13g2_nor2_1 _1292_ (.A(net124),
    .B(_0606_),
    .Y(_0611_));
 sg13g2_or3_1 _1293_ (.A(net251),
    .B(_0610_),
    .C(_0611_),
    .X(_0612_));
 sg13g2_a21oi_1 _1294_ (.A1(net116),
    .A2(net251),
    .Y(_0613_),
    .B1(net252));
 sg13g2_a22oi_1 _1295_ (.Y(_0068_),
    .B1(_0612_),
    .B2(_0613_),
    .A2(net252),
    .A1(_0132_));
 sg13g2_a21oi_1 _1296_ (.A1(_0566_),
    .A2(_0610_),
    .Y(_0614_),
    .B1(net114));
 sg13g2_and3_1 _1297_ (.X(_0615_),
    .A(\cpu.pc_s[10] ),
    .B(_0566_),
    .C(_0610_));
 sg13g2_nor2_1 _1298_ (.A(_0614_),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_mux2_1 _1299_ (.A0(net96),
    .A1(_0616_),
    .S(net250),
    .X(_0069_));
 sg13g2_nand3_1 _1300_ (.B(\cpu.pc_s[11] ),
    .C(_0610_),
    .A(\cpu.pc_s[10] ),
    .Y(_0617_));
 sg13g2_xor2_1 _1301_ (.B(_0615_),
    .A(\cpu.pc_s[11] ),
    .X(_0618_));
 sg13g2_mux2_1 _1302_ (.A0(net105),
    .A1(_0618_),
    .S(net250),
    .X(_0070_));
 sg13g2_xnor2_1 _1303_ (.Y(_0619_),
    .A(net112),
    .B(_0617_));
 sg13g2_nand2b_1 _1304_ (.Y(_0620_),
    .B(_0619_),
    .A_N(net251));
 sg13g2_a21oi_1 _1305_ (.A1(\cpu.regA_s[12] ),
    .A2(net251),
    .Y(_0621_),
    .B1(net252));
 sg13g2_a22oi_1 _1306_ (.Y(_0071_),
    .B1(_0620_),
    .B2(_0621_),
    .A2(net252),
    .A1(_0133_));
 sg13g2_nand3_1 _1307_ (.B(\cpu.pc_s[12] ),
    .C(_0615_),
    .A(\cpu.pc_s[11] ),
    .Y(_0622_));
 sg13g2_xnor2_1 _1308_ (.Y(_0623_),
    .A(\cpu.pc_s[13] ),
    .B(_0622_));
 sg13g2_mux2_1 _1309_ (.A0(net134),
    .A1(_0623_),
    .S(net250),
    .X(_0072_));
 sg13g2_nand4_1 _1310_ (.B(\cpu.pc_s[12] ),
    .C(\cpu.pc_s[13] ),
    .A(\cpu.pc_s[11] ),
    .Y(_0624_),
    .D(_0615_));
 sg13g2_nor2_1 _1311_ (.A(_0134_),
    .B(_0624_),
    .Y(_0625_));
 sg13g2_xnor2_1 _1312_ (.Y(_0626_),
    .A(net133),
    .B(_0624_));
 sg13g2_mux2_1 _1313_ (.A0(net117),
    .A1(_0626_),
    .S(net250),
    .X(_0073_));
 sg13g2_xor2_1 _1314_ (.B(_0625_),
    .A(\cpu.pc_s[15] ),
    .X(_0627_));
 sg13g2_mux2_1 _1315_ (.A0(net122),
    .A1(_0627_),
    .S(net250),
    .X(_0074_));
 sg13g2_nor2b_1 _1316_ (.A(_0136_),
    .B_N(_0572_),
    .Y(_0628_));
 sg13g2_mux2_1 _1317_ (.A0(net80),
    .A1(net2),
    .S(net260),
    .X(_0075_));
 sg13g2_nor2b_1 _1318_ (.A(net3),
    .B_N(\cpu.spi_debug_instance.counter_s[4] ),
    .Y(_0629_));
 sg13g2_mux2_1 _1319_ (.A0(\cpu.spi_debug_instance.in_s[0] ),
    .A1(net4),
    .S(_0629_),
    .X(_0076_));
 sg13g2_mux2_1 _1320_ (.A0(\cpu.spi_debug_instance.in_s[1] ),
    .A1(\cpu.spi_debug_instance.in_s[0] ),
    .S(_0629_),
    .X(_0077_));
 sg13g2_nor2_1 _1321_ (.A(net39),
    .B(net258),
    .Y(_0630_));
 sg13g2_a21oi_1 _1322_ (.A1(_0126_),
    .A2(net258),
    .Y(_0078_),
    .B1(_0630_));
 sg13g2_nor2_1 _1323_ (.A(net44),
    .B(net258),
    .Y(_0631_));
 sg13g2_a21oi_1 _1324_ (.A1(_0124_),
    .A2(net258),
    .Y(_0079_),
    .B1(_0631_));
 sg13g2_nand2_1 _1325_ (.Y(_0632_),
    .A(net42),
    .B(net259));
 sg13g2_o21ai_1 _1326_ (.B1(_0632_),
    .Y(_0080_),
    .A1(_0126_),
    .A2(net258));
 sg13g2_nor2_1 _1327_ (.A(net47),
    .B(net260),
    .Y(_0633_));
 sg13g2_a21oi_1 _1328_ (.A1(_0121_),
    .A2(net260),
    .Y(_0081_),
    .B1(_0633_));
 sg13g2_mux2_1 _1329_ (.A0(net79),
    .A1(net47),
    .S(net261),
    .X(_0082_));
 sg13g2_mux2_1 _1330_ (.A0(net72),
    .A1(\cpu.inM_s[1] ),
    .S(net260),
    .X(_0083_));
 sg13g2_mux2_1 _1331_ (.A0(net42),
    .A1(net63),
    .S(net258),
    .X(_0084_));
 sg13g2_mux2_1 _1332_ (.A0(net81),
    .A1(net72),
    .S(net260),
    .X(_0085_));
 sg13g2_mux2_1 _1333_ (.A0(net67),
    .A1(\cpu.inM_s[3] ),
    .S(net260),
    .X(_0086_));
 sg13g2_mux2_1 _1334_ (.A0(net75),
    .A1(net67),
    .S(net260),
    .X(_0087_));
 sg13g2_mux2_1 _1335_ (.A0(net63),
    .A1(net74),
    .S(net259),
    .X(_0088_));
 sg13g2_mux2_1 _1336_ (.A0(net85),
    .A1(net75),
    .S(net261),
    .X(_0089_));
 sg13g2_mux2_1 _1337_ (.A0(net53),
    .A1(\cpu.inM_s[6] ),
    .S(net260),
    .X(_0090_));
 sg13g2_nor2_1 _1338_ (.A(net46),
    .B(net258),
    .Y(_0634_));
 sg13g2_a21oi_1 _1339_ (.A1(_0125_),
    .A2(net258),
    .Y(_0091_),
    .B1(_0634_));
 sg13g2_nor2_1 _1340_ (.A(_0136_),
    .B(_0572_),
    .Y(_0635_));
 sg13g2_mux2_1 _1341_ (.A0(net48),
    .A1(net2),
    .S(net254),
    .X(_0092_));
 sg13g2_mux2_1 _1342_ (.A0(net74),
    .A1(net80),
    .S(net259),
    .X(_0093_));
 sg13g2_mux2_1 _1343_ (.A0(net58),
    .A1(net302),
    .S(net253),
    .X(_0094_));
 sg13g2_nand2_1 _1344_ (.Y(_0636_),
    .A(net38),
    .B(net253));
 sg13g2_o21ai_1 _1345_ (.B1(_0636_),
    .Y(_0095_),
    .A1(_0120_),
    .A2(net255));
 sg13g2_mux2_1 _1346_ (.A0(net302),
    .A1(net299),
    .S(net253),
    .X(_0096_));
 sg13g2_nor2_1 _1347_ (.A(net61),
    .B(net255),
    .Y(_0637_));
 sg13g2_a21oi_1 _1348_ (.A1(_0120_),
    .A2(net255),
    .Y(_0097_),
    .B1(_0637_));
 sg13g2_nand2_1 _1349_ (.Y(_0638_),
    .A(net61),
    .B(net255));
 sg13g2_o21ai_1 _1350_ (.B1(_0638_),
    .Y(_0098_),
    .A1(_0129_),
    .A2(net256));
 sg13g2_nor2_1 _1351_ (.A(net59),
    .B(net256),
    .Y(_0639_));
 sg13g2_a21oi_1 _1352_ (.A1(_0129_),
    .A2(net256),
    .Y(_0099_),
    .B1(_0639_));
 sg13g2_mux2_1 _1353_ (.A0(net299),
    .A1(net70),
    .S(net253),
    .X(_0100_));
 sg13g2_nor2_1 _1354_ (.A(net76),
    .B(net256),
    .Y(_0640_));
 sg13g2_a21oi_1 _1355_ (.A1(_0128_),
    .A2(net255),
    .Y(_0101_),
    .B1(_0640_));
 sg13g2_mux2_1 _1356_ (.A0(net94),
    .A1(net76),
    .S(net255),
    .X(_0102_));
 sg13g2_mux2_1 _1357_ (.A0(net66),
    .A1(net94),
    .S(net255),
    .X(_0103_));
 sg13g2_nor2_1 _1358_ (.A(net70),
    .B(net254),
    .Y(_0641_));
 sg13g2_a21oi_1 _1359_ (.A1(net290),
    .A2(net254),
    .Y(_0104_),
    .B1(_0641_));
 sg13g2_mux2_1 _1360_ (.A0(net41),
    .A1(net66),
    .S(net255),
    .X(_0105_));
 sg13g2_nand2_1 _1361_ (.Y(_0642_),
    .A(net41),
    .B(net253));
 sg13g2_o21ai_1 _1362_ (.B1(_0642_),
    .Y(_0106_),
    .A1(_0127_),
    .A2(net254));
 sg13g2_mux2_1 _1363_ (.A0(net38),
    .A1(net58),
    .S(net253),
    .X(_0107_));
 sg13g2_nand2_1 _1364_ (.Y(_0643_),
    .A(net48),
    .B(net253));
 sg13g2_o21ai_1 _1365_ (.B1(_0643_),
    .Y(_0114_),
    .A1(net290),
    .A2(net253));
 sg13g2_inv_1 _1366_ (.Y(_0010_),
    .A(net5));
 sg13g2_inv_1 _1367_ (.Y(_0011_),
    .A(net5));
 sg13g2_inv_1 _1368_ (.Y(_0012_),
    .A(net5));
 sg13g2_inv_1 _1369_ (.Y(_0013_),
    .A(net5));
 sg13g2_inv_1 _1371__4 (.Y(net29),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _1372__5 (.Y(net30),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _1373__6 (.Y(net31),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _1374__7 (.Y(net32),
    .A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbp_1 _1375_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net331),
    .D(_0020_),
    .Q_N(_0729_),
    .Q(\cpu.alu_instance.a_i[0] ));
 sg13g2_dfrbp_1 _1376_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net332),
    .D(_0021_),
    .Q_N(_0728_),
    .Q(\cpu.alu_instance.a_i[1] ));
 sg13g2_dfrbp_1 _1377_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net331),
    .D(_0022_),
    .Q_N(_0727_),
    .Q(\cpu.alu_instance.a_i[2] ));
 sg13g2_dfrbp_1 _1378_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net331),
    .D(_0023_),
    .Q_N(_0726_),
    .Q(\cpu.alu_instance.a_i[3] ));
 sg13g2_dfrbp_1 _1379_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net331),
    .D(_0024_),
    .Q_N(_0725_),
    .Q(\cpu.alu_instance.a_i[4] ));
 sg13g2_dfrbp_1 _1380_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net333),
    .D(_0025_),
    .Q_N(_0724_),
    .Q(\cpu.alu_instance.a_i[5] ));
 sg13g2_dfrbp_1 _1381_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net327),
    .D(_0026_),
    .Q_N(_0723_),
    .Q(\cpu.alu_instance.a_i[6] ));
 sg13g2_dfrbp_1 _1382_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net327),
    .D(_0027_),
    .Q_N(_0722_),
    .Q(\cpu.alu_instance.a_i[7] ));
 sg13g2_dfrbp_1 _1383_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net327),
    .D(_0028_),
    .Q_N(_0721_),
    .Q(\cpu.alu_instance.a_i[8] ));
 sg13g2_dfrbp_1 _1384_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net327),
    .D(_0029_),
    .Q_N(_0720_),
    .Q(\cpu.alu_instance.a_i[9] ));
 sg13g2_dfrbp_1 _1385_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net320),
    .D(_0030_),
    .Q_N(_0719_),
    .Q(\cpu.alu_instance.a_i[10] ));
 sg13g2_dfrbp_1 _1386_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net325),
    .D(_0031_),
    .Q_N(_0718_),
    .Q(\cpu.alu_instance.a_i[11] ));
 sg13g2_dfrbp_1 _1387_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net321),
    .D(_0032_),
    .Q_N(_0717_),
    .Q(\cpu.alu_instance.a_i[12] ));
 sg13g2_dfrbp_1 _1388_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net321),
    .D(_0033_),
    .Q_N(_0716_),
    .Q(\cpu.alu_instance.a_i[13] ));
 sg13g2_dfrbp_1 _1389_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net322),
    .D(_0034_),
    .Q_N(_0715_),
    .Q(\cpu.alu_instance.a_i[14] ));
 sg13g2_dfrbp_1 _1390_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net325),
    .D(_0035_),
    .Q_N(_0714_),
    .Q(\cpu.alu_instance.a_i[15] ));
 sg13g2_dfrbp_1 _1391_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net326),
    .D(net111),
    .Q_N(_0713_),
    .Q(\cpu.regA_s[0] ));
 sg13g2_dfrbp_1 _1392_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net326),
    .D(net132),
    .Q_N(_0712_),
    .Q(\cpu.regA_s[1] ));
 sg13g2_dfrbp_1 _1393_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net330),
    .D(_0038_),
    .Q_N(_0711_),
    .Q(\cpu.regA_s[2] ));
 sg13g2_dfrbp_1 _1394_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net331),
    .D(_0039_),
    .Q_N(_0710_),
    .Q(\cpu.regA_s[3] ));
 sg13g2_dfrbp_1 _1395_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net330),
    .D(_0040_),
    .Q_N(_0709_),
    .Q(\cpu.regA_s[4] ));
 sg13g2_dfrbp_1 _1396_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net330),
    .D(_0041_),
    .Q_N(_0708_),
    .Q(\cpu.regA_s[5] ));
 sg13g2_dfrbp_1 _1397_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net327),
    .D(_0042_),
    .Q_N(_0707_),
    .Q(\cpu.regA_s[6] ));
 sg13g2_dfrbp_1 _1398_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net326),
    .D(_0043_),
    .Q_N(_0706_),
    .Q(\cpu.regA_s[7] ));
 sg13g2_dfrbp_1 _1399_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net326),
    .D(_0044_),
    .Q_N(_0705_),
    .Q(\cpu.regA_s[8] ));
 sg13g2_dfrbp_1 _1400_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net326),
    .D(_0045_),
    .Q_N(_0704_),
    .Q(\cpu.regA_s[9] ));
 sg13g2_dfrbp_1 _1401_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net320),
    .D(_0046_),
    .Q_N(_0703_),
    .Q(\cpu.regA_s[10] ));
 sg13g2_dfrbp_1 _1402_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net320),
    .D(_0047_),
    .Q_N(_0702_),
    .Q(\cpu.regA_s[11] ));
 sg13g2_dfrbp_1 _1403_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net320),
    .D(_0048_),
    .Q_N(_0701_),
    .Q(\cpu.regA_s[12] ));
 sg13g2_dfrbp_1 _1404_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net318),
    .D(_0049_),
    .Q_N(_0700_),
    .Q(\cpu.regA_s[13] ));
 sg13g2_dfrbp_1 _1405_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net319),
    .D(_0050_),
    .Q_N(_0699_),
    .Q(\cpu.regA_s[14] ));
 sg13g2_dfrbp_1 _1406_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net319),
    .D(net51),
    .Q_N(_0698_),
    .Q(\cpu.regA_s[15] ));
 sg13g2_dfrbp_1 _1407_ (.CLK(_0009_),
    .RESET_B(net329),
    .D(_0052_),
    .Q_N(_0008_),
    .Q(\cpu.spi_debug_instance.counter_s[0] ));
 sg13g2_dfrbp_1 _1408_ (.CLK(_0010_),
    .RESET_B(net329),
    .D(_0053_),
    .Q_N(_0697_),
    .Q(\cpu.spi_debug_instance.counter_s[1] ));
 sg13g2_dfrbp_1 _1409_ (.CLK(_0011_),
    .RESET_B(net330),
    .D(_0054_),
    .Q_N(_0696_),
    .Q(\cpu.spi_debug_instance.counter_s[2] ));
 sg13g2_dfrbp_1 _1410_ (.CLK(_0012_),
    .RESET_B(net329),
    .D(_0055_),
    .Q_N(_0695_),
    .Q(\cpu.spi_debug_instance.counter_s[3] ));
 sg13g2_dfrbp_1 _1411_ (.CLK(_0013_),
    .RESET_B(net329),
    .D(_0056_),
    .Q_N(_0694_),
    .Q(\cpu.spi_debug_instance.counter_s[4] ));
 sg13g2_dfrbp_1 _1412_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net322),
    .D(_0057_),
    .Q_N(_0693_),
    .Q(\cpu.fsm_instance.state_s[0] ));
 sg13g2_dfrbp_1 _1413_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net323),
    .D(_0058_),
    .Q_N(_0692_),
    .Q(\cpu.fsm_instance.state_s[1] ));
 sg13g2_dfrbp_1 _1414_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net331),
    .D(net93),
    .Q_N(_0691_),
    .Q(\cpu.pc_s[0] ));
 sg13g2_dfrbp_1 _1415_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net332),
    .D(net101),
    .Q_N(_0005_),
    .Q(\cpu.pc_s[1] ));
 sg13g2_dfrbp_1 _1416_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net332),
    .D(_0061_),
    .Q_N(_0690_),
    .Q(\cpu.pc_s[2] ));
 sg13g2_dfrbp_1 _1417_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net332),
    .D(net126),
    .Q_N(_0689_),
    .Q(\cpu.pc_s[3] ));
 sg13g2_dfrbp_1 _1418_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net331),
    .D(_0063_),
    .Q_N(_0688_),
    .Q(\cpu.pc_s[4] ));
 sg13g2_dfrbp_1 _1419_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net331),
    .D(_0064_),
    .Q_N(_0687_),
    .Q(\cpu.pc_s[5] ));
 sg13g2_dfrbp_1 _1420_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net332),
    .D(_0065_),
    .Q_N(_0686_),
    .Q(\cpu.pc_s[6] ));
 sg13g2_dfrbp_1 _1421_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net332),
    .D(_0066_),
    .Q_N(_0685_),
    .Q(\cpu.pc_s[7] ));
 sg13g2_dfrbp_1 _1422_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net329),
    .D(_0067_),
    .Q_N(_0684_),
    .Q(\cpu.pc_s[8] ));
 sg13g2_dfrbp_1 _1423_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net329),
    .D(_0068_),
    .Q_N(_0683_),
    .Q(\cpu.pc_s[9] ));
 sg13g2_dfrbp_1 _1424_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net324),
    .D(_0069_),
    .Q_N(_0682_),
    .Q(\cpu.pc_s[10] ));
 sg13g2_dfrbp_1 _1425_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net324),
    .D(net106),
    .Q_N(_0681_),
    .Q(\cpu.pc_s[11] ));
 sg13g2_dfrbp_1 _1426_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net324),
    .D(net113),
    .Q_N(_0680_),
    .Q(\cpu.pc_s[12] ));
 sg13g2_dfrbp_1 _1427_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net324),
    .D(net135),
    .Q_N(_0679_),
    .Q(\cpu.pc_s[13] ));
 sg13g2_dfrbp_1 _1428_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net322),
    .D(_0073_),
    .Q_N(_0678_),
    .Q(\cpu.pc_s[14] ));
 sg13g2_dfrbp_1 _1429_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net322),
    .D(net123),
    .Q_N(_0677_),
    .Q(\cpu.pc_s[15] ));
 sg13g2_dfrbp_1 _1430_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net326),
    .D(_0075_),
    .Q_N(_0676_),
    .Q(\cpu.inM_s[8] ));
 sg13g2_dfrbp_1 _1431_ (.CLK(net5),
    .RESET_B(net329),
    .D(_0076_),
    .Q_N(_0675_),
    .Q(\cpu.spi_debug_instance.in_s[0] ));
 sg13g2_dfrbp_1 _1432_ (.CLK(net5),
    .RESET_B(net329),
    .D(_0077_),
    .Q_N(_0730_),
    .Q(\cpu.spi_debug_instance.in_s[1] ));
 sg13g2_dfrbp_1 _1433_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net323),
    .D(\cpu.spi_mem_instance.next_state_s[0] ),
    .Q_N(_0731_),
    .Q(\cpu.spi_mem_instance.state_s[0] ));
 sg13g2_dfrbp_1 _1434_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net323),
    .D(\cpu.spi_mem_instance.next_state_s[1] ),
    .Q_N(_0732_),
    .Q(\cpu.spi_mem_instance.state_s[1] ));
 sg13g2_dfrbp_1 _1435_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net323),
    .D(net35),
    .Q_N(_0000_),
    .Q(\cpu.spi_mem_instance.state_s[2] ));
 sg13g2_dfrbp_1 _1436_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net318),
    .D(net40),
    .Q_N(_0674_),
    .Q(\cpu.inM_s[13] ));
 sg13g2_dfrbp_1 _1437_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net318),
    .D(net45),
    .Q_N(_0673_),
    .Q(\cpu.inM_s[15] ));
 sg13g2_dfrbp_1 _1438_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net318),
    .D(net43),
    .Q_N(_0672_),
    .Q(\cpu.inM_s[12] ));
 sg13g2_dfrbp_1 _1439_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net326),
    .D(_0081_),
    .Q_N(_0671_),
    .Q(\cpu.inM_s[0] ));
 sg13g2_dfrbp_1 _1440_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net328),
    .D(_0082_),
    .Q_N(_0670_),
    .Q(\cpu.inM_s[1] ));
 sg13g2_dfrbp_1 _1441_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net328),
    .D(net73),
    .Q_N(_0669_),
    .Q(\cpu.inM_s[2] ));
 sg13g2_dfrbp_1 _1442_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net320),
    .D(_0084_),
    .Q_N(_0668_),
    .Q(\cpu.inM_s[11] ));
 sg13g2_dfrbp_1 _1443_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net328),
    .D(_0085_),
    .Q_N(_0667_),
    .Q(\cpu.inM_s[3] ));
 sg13g2_dfrbp_1 _1444_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net328),
    .D(net68),
    .Q_N(_0666_),
    .Q(\cpu.inM_s[4] ));
 sg13g2_dfrbp_1 _1445_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net328),
    .D(_0087_),
    .Q_N(_0665_),
    .Q(\cpu.inM_s[5] ));
 sg13g2_dfrbp_1 _1446_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net320),
    .D(_0088_),
    .Q_N(_0664_),
    .Q(\cpu.inM_s[10] ));
 sg13g2_dfrbp_1 _1447_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net333),
    .D(_0089_),
    .Q_N(_0663_),
    .Q(\cpu.inM_s[6] ));
 sg13g2_dfrbp_1 _1448_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net328),
    .D(net54),
    .Q_N(_0662_),
    .Q(\cpu.inM_s[7] ));
 sg13g2_dfrbp_1 _1449_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net318),
    .D(_0091_),
    .Q_N(_0661_),
    .Q(\cpu.inM_s[14] ));
 sg13g2_dfrbp_1 _1450_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net320),
    .D(_0092_),
    .Q_N(_0003_),
    .Q(\cpu.alu_instance.nb_i ));
 sg13g2_dfrbp_1 _1451_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net326),
    .D(_0093_),
    .Q_N(_0660_),
    .Q(\cpu.inM_s[9] ));
 sg13g2_dfrbp_1 _1452_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net318),
    .D(_0094_),
    .Q_N(_0659_),
    .Q(\cpu.fsm_instance.instruction_i[13] ));
 sg13g2_dfrbp_1 _1453_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net319),
    .D(_0095_),
    .Q_N(_0001_),
    .Q(\cpu.fsm_instance.instruction_i[15] ));
 sg13g2_dfrbp_1 _1454_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net318),
    .D(_0096_),
    .Q_N(_0658_),
    .Q(\cpu.fsm_instance.instruction_i[12] ));
 sg13g2_dfrbp_1 _1455_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net321),
    .D(_0097_),
    .Q_N(_0657_),
    .Q(\cpu.fsm_instance.instruction_i[0] ));
 sg13g2_dfrbp_1 _1456_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net321),
    .D(net62),
    .Q_N(_0656_),
    .Q(\cpu.fsm_instance.instruction_i[1] ));
 sg13g2_dfrbp_1 _1457_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net322),
    .D(net60),
    .Q_N(_0655_),
    .Q(\cpu.fsm_instance.instruction_i[2] ));
 sg13g2_dfrbp_1 _1458_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net318),
    .D(_0100_),
    .Q_N(_0654_),
    .Q(\cpu.alu_instance.za_i ));
 sg13g2_dfrbp_1 _1459_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net322),
    .D(_0101_),
    .Q_N(_0653_),
    .Q(\cpu.fsm_instance.instruction_i[3] ));
 sg13g2_dfrbp_1 _1460_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net322),
    .D(_0102_),
    .Q_N(_0652_),
    .Q(\cpu.fsm_instance.instruction_i[4] ));
 sg13g2_dfrbp_1 _1461_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net319),
    .D(_0103_),
    .Q_N(_0651_),
    .Q(\cpu.fsm_instance.instruction_i[5] ));
 sg13g2_dfrbp_1 _1462_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net319),
    .D(net71),
    .Q_N(_0004_),
    .Q(\cpu.alu_instance.na_i ));
 sg13g2_dfrbp_1 _1463_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net321),
    .D(_0105_),
    .Q_N(_0002_),
    .Q(\cpu.alu_instance.no_i ));
 sg13g2_dfrbp_1 _1464_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net319),
    .D(_0106_),
    .Q_N(_0650_),
    .Q(\cpu.alu_instance.f_i ));
 sg13g2_dfrbp_1 _1465_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net319),
    .D(_0107_),
    .Q_N(_0649_),
    .Q(\cpu.fsm_instance.instruction_i[14] ));
 sg13g2_dfrbp_1 _1466_ (.CLK(net26),
    .RESET_B(net323),
    .D(net37),
    .Q_N(_0007_),
    .Q(\cpu.spi_mem_instance.count_s[0] ));
 sg13g2_dfrbp_1 _1467_ (.CLK(net28),
    .RESET_B(net322),
    .D(_0109_),
    .Q_N(_0648_),
    .Q(\cpu.spi_mem_instance.count_s[1] ));
 sg13g2_dfrbp_1 _1468_ (.CLK(net29),
    .RESET_B(net324),
    .D(net142),
    .Q_N(_0647_),
    .Q(\cpu.spi_mem_instance.count_s[2] ));
 sg13g2_dfrbp_1 _1469_ (.CLK(net30),
    .RESET_B(net324),
    .D(net99),
    .Q_N(_0646_),
    .Q(\cpu.spi_mem_instance.count_s[3] ));
 sg13g2_dfrbp_1 _1470_ (.CLK(net31),
    .RESET_B(net323),
    .D(_0112_),
    .Q_N(_0006_),
    .Q(\cpu.spi_mem_instance.count_s[4] ));
 sg13g2_dfrbp_1 _1471_ (.CLK(net32),
    .RESET_B(net323),
    .D(net109),
    .Q_N(_0645_),
    .Q(\cpu.spi_mem_instance.count_s[5] ));
 sg13g2_dfrbp_1 _1472_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net320),
    .D(net49),
    .Q_N(_0644_),
    .Q(\cpu.alu_instance.zb_i ));
 sg13g2_tiehi tt_um_hack_cpu_23 (.L_HI(net23));
 sg13g2_tiehi tt_um_hack_cpu_24 (.L_HI(net24));
 sg13g2_tiehi tt_um_hack_cpu_25 (.L_HI(net25));
 sg13g2_inv_1 _0753__1 (.Y(net26),
    .A(clknet_1_1__leaf_clk));
 sg13g2_tielo tt_um_hack_cpu_7 (.L_LO(net7));
 sg13g2_tielo tt_um_hack_cpu_8 (.L_LO(net8));
 sg13g2_tielo tt_um_hack_cpu_9 (.L_LO(net9));
 sg13g2_tielo tt_um_hack_cpu_10 (.L_LO(net10));
 sg13g2_tielo tt_um_hack_cpu_11 (.L_LO(net11));
 sg13g2_tielo tt_um_hack_cpu_12 (.L_LO(net12));
 sg13g2_tielo tt_um_hack_cpu_13 (.L_LO(net13));
 sg13g2_tielo tt_um_hack_cpu_14 (.L_LO(net14));
 sg13g2_tielo tt_um_hack_cpu_15 (.L_LO(net15));
 sg13g2_tielo tt_um_hack_cpu_16 (.L_LO(net16));
 sg13g2_tielo tt_um_hack_cpu_17 (.L_LO(net17));
 sg13g2_tielo tt_um_hack_cpu_18 (.L_LO(net18));
 sg13g2_tielo tt_um_hack_cpu_19 (.L_LO(net19));
 sg13g2_tielo tt_um_hack_cpu_20 (.L_LO(net20));
 sg13g2_tielo tt_um_hack_cpu_21 (.L_LO(net21));
 sg13g2_tiehi tt_um_hack_cpu_22 (.L_HI(net22));
 sg13g2_buf_1 _1493_ (.A(\cpu.mem_csb_o ),
    .X(uio_out[0]));
 sg13g2_buf_1 _1494_ (.A(\cpu.mem_out_o ),
    .X(uio_out[1]));
 sg13g2_buf_1 _1495_ (.A(\cpu.mem_sclk_o ),
    .X(uio_out[3]));
 sg13g2_buf_1 _1496_ (.A(\cpu.debug_out_o ),
    .X(uio_out[6]));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(_0587_));
 sg13g2_buf_2 fanout251 (.A(_0586_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_0567_),
    .X(net252));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(net257));
 sg13g2_buf_2 fanout254 (.A(net257),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(net257),
    .X(net255));
 sg13g2_buf_1 fanout256 (.A(net257),
    .X(net256));
 sg13g2_buf_1 fanout257 (.A(_0635_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net259),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(net261),
    .X(net259));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(net261));
 sg13g2_buf_2 fanout261 (.A(_0628_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(net263),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_0530_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(net265),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_0529_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(net267),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_0515_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(net269),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_0515_),
    .X(net269));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(net138));
 sg13g2_buf_2 fanout271 (.A(\cpu.spi_mem_instance.count_s[1] ),
    .X(net271));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(net275));
 sg13g2_buf_2 fanout273 (.A(net275),
    .X(net273));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(net275));
 sg13g2_buf_2 fanout275 (.A(\cpu.spi_mem_instance.count_s[0] ),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(\cpu.spi_debug_instance.counter_s[3] ),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(net278),
    .X(net277));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(_0460_));
 sg13g2_buf_2 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_0459_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(net282),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_0458_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(net285),
    .X(net283));
 sg13g2_buf_1 fanout284 (.A(_0123_),
    .X(net284));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_0123_));
 sg13g2_buf_2 fanout286 (.A(net289),
    .X(net286));
 sg13g2_buf_1 fanout287 (.A(net288),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_1 fanout289 (.A(net290),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_0122_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(\cpu.alu_instance.f_i ),
    .X(net291));
 sg13g2_buf_1 fanout292 (.A(\cpu.alu_instance.f_i ),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(net294),
    .X(net293));
 sg13g2_buf_1 fanout294 (.A(\cpu.alu_instance.f_i ),
    .X(net294));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(_0002_));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(_0002_));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(net298));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(_0004_));
 sg13g2_buf_2 fanout299 (.A(net301),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(net301),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(\cpu.alu_instance.za_i ),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(net303),
    .X(net302));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(net305));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(net305));
 sg13g2_buf_2 fanout305 (.A(\cpu.fsm_instance.instruction_i[12] ),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(net307),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(net310),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(net309),
    .X(net308));
 sg13g2_buf_1 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_1 fanout310 (.A(\cpu.fsm_instance.instruction_i[15] ),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(net312),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_0003_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(net316),
    .X(net313));
 sg13g2_buf_1 fanout314 (.A(net316),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(net316),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(\cpu.fsm_instance.state_s[1] ),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(net115),
    .X(net317));
 sg13g2_buf_4 fanout318 (.X(net318),
    .A(net319));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(net321));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(net321));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(net325));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(net324));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(net324));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(net325));
 sg13g2_buf_2 fanout325 (.A(rst_n),
    .X(net325));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(net328));
 sg13g2_buf_2 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(net333));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(net330));
 sg13g2_buf_2 fanout330 (.A(net333),
    .X(net330));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(net332));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(net333));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(uio_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[5]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(uio_in[7]),
    .X(net5));
 sg13g2_tielo tt_um_hack_cpu_6 (.L_LO(net6));
 sg13g2_inv_1 _0753__2 (.Y(net27),
    .A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_4_1_0_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_4_5_0_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_4_6_0_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_4_7_0_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_4_9_0_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_4_10_0_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_4_11_0_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_4_13_0_clk_regs));
 sg13g2_inv_1 clkload10 (.A(clknet_4_14_0_clk_regs));
 sg13g2_inv_1 clkload11 (.A(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0000_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0137_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold3 (.A(\cpu.spi_mem_instance.next_state_s[2] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0007_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0108_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold6 (.A(\cpu.fsm_instance.instruction_i[14] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cpu.inM_s[13] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0078_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold9 (.A(\cpu.alu_instance.no_i ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cpu.inM_s[11] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0080_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cpu.inM_s[15] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0079_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cpu.inM_s[14] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold15 (.A(\cpu.inM_s[0] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cpu.alu_instance.nb_i ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0114_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0001_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0051_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold20 (.A(\cpu.alu_instance.a_i[8] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold21 (.A(\cpu.inM_s[7] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0090_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold23 (.A(\cpu.alu_instance.a_i[9] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cpu.alu_instance.a_i[5] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold25 (.A(\cpu.alu_instance.a_i[1] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold26 (.A(\cpu.fsm_instance.instruction_i[13] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold27 (.A(\cpu.fsm_instance.instruction_i[2] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0099_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cpu.fsm_instance.instruction_i[0] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0098_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cpu.inM_s[10] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold32 (.A(\cpu.alu_instance.a_i[0] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold33 (.A(\cpu.alu_instance.a_i[15] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cpu.fsm_instance.instruction_i[5] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cpu.inM_s[4] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0086_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold37 (.A(\cpu.alu_instance.a_i[13] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold38 (.A(\cpu.alu_instance.na_i ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0104_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cpu.inM_s[2] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0083_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold42 (.A(\cpu.inM_s[9] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cpu.inM_s[5] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold44 (.A(\cpu.fsm_instance.instruction_i[3] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold45 (.A(\cpu.alu_instance.a_i[6] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold46 (.A(\cpu.alu_instance.a_i[4] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cpu.inM_s[1] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cpu.inM_s[8] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold49 (.A(\cpu.inM_s[3] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cpu.spi_mem_instance.state_s[0] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0136_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cpu.alu_instance.a_i[2] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold53 (.A(\cpu.inM_s[6] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cpu.alu_instance.a_i[11] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cpu.alu_instance.a_i[12] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cpu.alu_instance.a_i[7] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold57 (.A(\cpu.alu_instance.a_i[10] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cpu.alu_instance.a_i[14] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cpu.alu_instance.a_i[3] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold60 (.A(\cpu.pc_s[0] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0059_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold62 (.A(\cpu.fsm_instance.instruction_i[4] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cpu.spi_mem_instance.state_s[1] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold64 (.A(\cpu.regA_s[10] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cpu.regA_s[5] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold66 (.A(\cpu.spi_mem_instance.count_s[3] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0111_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cpu.pc_s[1] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0060_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold70 (.A(\cpu.regA_s[7] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cpu.regA_s[4] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0539_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cpu.regA_s[11] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0070_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cpu.spi_mem_instance.count_s[5] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0148_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0113_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cpu.regA_s[0] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0036_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cpu.pc_s[12] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0071_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cpu.pc_s[10] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cpu.fsm_instance.state_s[0] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cpu.regA_s[9] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold85 (.A(\cpu.regA_s[14] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold86 (.A(\cpu.regA_s[2] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0141_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold88 (.A(\cpu.regA_s[6] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cpu.regA_s[12] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cpu.regA_s[15] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0074_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cpu.pc_s[9] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cpu.regA_s[3] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0062_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cpu.regA_s[8] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold96 (.A(\cpu.spi_mem_instance.count_s[4] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cpu.pc_s[2] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cpu.pc_s[5] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold99 (.A(\cpu.regA_s[1] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0037_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cpu.pc_s[14] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cpu.regA_s[13] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0072_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cpu.pc_s[7] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0604_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cpu.spi_mem_instance.count_s[1] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cpu.pc_s[6] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cpu.pc_s[8] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cpu.spi_mem_instance.count_s[2] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0110_),
    .X(net142));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_4 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_151 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_180 ();
 sg13g2_decap_4 FILLER_9_187 ();
 sg13g2_fill_1 FILLER_9_191 ();
 sg13g2_decap_8 FILLER_9_218 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_decap_8 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_239 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_260 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_281 ();
 sg13g2_decap_8 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_295 ();
 sg13g2_decap_8 FILLER_9_302 ();
 sg13g2_decap_8 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_316 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_337 ();
 sg13g2_decap_8 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_351 ();
 sg13g2_fill_1 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_4 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_185 ();
 sg13g2_fill_1 FILLER_10_187 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_234 ();
 sg13g2_decap_8 FILLER_10_241 ();
 sg13g2_decap_8 FILLER_10_248 ();
 sg13g2_decap_8 FILLER_10_255 ();
 sg13g2_decap_8 FILLER_10_262 ();
 sg13g2_decap_8 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_fill_2 FILLER_10_290 ();
 sg13g2_fill_1 FILLER_10_292 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_fill_2 FILLER_10_330 ();
 sg13g2_decap_4 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_fill_1 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_146 ();
 sg13g2_fill_1 FILLER_11_192 ();
 sg13g2_decap_4 FILLER_11_202 ();
 sg13g2_fill_2 FILLER_11_206 ();
 sg13g2_decap_4 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_233 ();
 sg13g2_fill_1 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_fill_2 FILLER_11_327 ();
 sg13g2_fill_1 FILLER_11_329 ();
 sg13g2_decap_4 FILLER_11_356 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_4 FILLER_12_91 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_decap_4 FILLER_12_132 ();
 sg13g2_fill_2 FILLER_12_136 ();
 sg13g2_fill_2 FILLER_12_156 ();
 sg13g2_decap_8 FILLER_12_167 ();
 sg13g2_decap_4 FILLER_12_174 ();
 sg13g2_fill_2 FILLER_12_191 ();
 sg13g2_fill_2 FILLER_12_203 ();
 sg13g2_decap_4 FILLER_12_241 ();
 sg13g2_fill_2 FILLER_12_245 ();
 sg13g2_fill_2 FILLER_12_275 ();
 sg13g2_fill_2 FILLER_12_303 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_fill_2 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_148 ();
 sg13g2_fill_1 FILLER_13_154 ();
 sg13g2_fill_2 FILLER_13_195 ();
 sg13g2_fill_1 FILLER_13_197 ();
 sg13g2_decap_8 FILLER_13_213 ();
 sg13g2_decap_4 FILLER_13_220 ();
 sg13g2_fill_2 FILLER_13_224 ();
 sg13g2_fill_2 FILLER_13_231 ();
 sg13g2_fill_1 FILLER_13_269 ();
 sg13g2_fill_2 FILLER_13_294 ();
 sg13g2_fill_1 FILLER_13_296 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_4 FILLER_13_322 ();
 sg13g2_fill_2 FILLER_13_326 ();
 sg13g2_decap_4 FILLER_13_338 ();
 sg13g2_fill_1 FILLER_13_342 ();
 sg13g2_fill_2 FILLER_13_353 ();
 sg13g2_fill_1 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_fill_1 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_4 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_90 ();
 sg13g2_decap_8 FILLER_14_97 ();
 sg13g2_decap_4 FILLER_14_104 ();
 sg13g2_fill_2 FILLER_14_108 ();
 sg13g2_decap_4 FILLER_14_145 ();
 sg13g2_fill_2 FILLER_14_170 ();
 sg13g2_decap_4 FILLER_14_180 ();
 sg13g2_fill_2 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_fill_1 FILLER_14_196 ();
 sg13g2_decap_4 FILLER_14_218 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_fill_2 FILLER_14_252 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_320 ();
 sg13g2_fill_2 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_fill_2 FILLER_14_360 ();
 sg13g2_fill_1 FILLER_14_372 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_63 ();
 sg13g2_fill_1 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_167 ();
 sg13g2_fill_1 FILLER_15_169 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_fill_2 FILLER_15_204 ();
 sg13g2_fill_1 FILLER_15_206 ();
 sg13g2_fill_1 FILLER_15_257 ();
 sg13g2_fill_1 FILLER_15_266 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_fill_1 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_fill_1 FILLER_15_304 ();
 sg13g2_fill_2 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_312 ();
 sg13g2_decap_4 FILLER_15_325 ();
 sg13g2_fill_2 FILLER_15_329 ();
 sg13g2_fill_2 FILLER_15_372 ();
 sg13g2_fill_2 FILLER_15_383 ();
 sg13g2_fill_1 FILLER_15_385 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_4 FILLER_16_42 ();
 sg13g2_fill_2 FILLER_16_46 ();
 sg13g2_fill_2 FILLER_16_74 ();
 sg13g2_fill_2 FILLER_16_159 ();
 sg13g2_fill_2 FILLER_16_183 ();
 sg13g2_fill_1 FILLER_16_195 ();
 sg13g2_fill_2 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_214 ();
 sg13g2_fill_1 FILLER_16_219 ();
 sg13g2_fill_2 FILLER_16_225 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_fill_2 FILLER_16_322 ();
 sg13g2_fill_1 FILLER_16_353 ();
 sg13g2_fill_2 FILLER_16_366 ();
 sg13g2_fill_2 FILLER_16_380 ();
 sg13g2_fill_1 FILLER_16_382 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_4 FILLER_17_49 ();
 sg13g2_fill_2 FILLER_17_73 ();
 sg13g2_fill_1 FILLER_17_82 ();
 sg13g2_fill_2 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_99 ();
 sg13g2_fill_2 FILLER_17_149 ();
 sg13g2_fill_1 FILLER_17_151 ();
 sg13g2_fill_1 FILLER_17_157 ();
 sg13g2_fill_2 FILLER_17_175 ();
 sg13g2_fill_2 FILLER_17_190 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_204 ();
 sg13g2_decap_4 FILLER_17_210 ();
 sg13g2_fill_2 FILLER_17_237 ();
 sg13g2_fill_1 FILLER_17_239 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_269 ();
 sg13g2_fill_2 FILLER_17_286 ();
 sg13g2_fill_2 FILLER_17_366 ();
 sg13g2_fill_1 FILLER_17_368 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_39 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_fill_2 FILLER_18_114 ();
 sg13g2_fill_1 FILLER_18_116 ();
 sg13g2_fill_1 FILLER_18_157 ();
 sg13g2_decap_4 FILLER_18_162 ();
 sg13g2_fill_2 FILLER_18_166 ();
 sg13g2_decap_8 FILLER_18_187 ();
 sg13g2_decap_8 FILLER_18_202 ();
 sg13g2_decap_4 FILLER_18_209 ();
 sg13g2_fill_1 FILLER_18_213 ();
 sg13g2_decap_4 FILLER_18_222 ();
 sg13g2_decap_4 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_240 ();
 sg13g2_fill_2 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_299 ();
 sg13g2_fill_1 FILLER_18_301 ();
 sg13g2_fill_2 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_321 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_2 FILLER_18_346 ();
 sg13g2_fill_2 FILLER_18_381 ();
 sg13g2_fill_1 FILLER_18_383 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_42 ();
 sg13g2_fill_1 FILLER_19_44 ();
 sg13g2_fill_2 FILLER_19_53 ();
 sg13g2_fill_1 FILLER_19_103 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_146 ();
 sg13g2_fill_2 FILLER_19_164 ();
 sg13g2_fill_1 FILLER_19_173 ();
 sg13g2_fill_1 FILLER_19_209 ();
 sg13g2_fill_2 FILLER_19_225 ();
 sg13g2_decap_4 FILLER_19_239 ();
 sg13g2_decap_4 FILLER_19_310 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_fill_2 FILLER_19_338 ();
 sg13g2_fill_1 FILLER_19_340 ();
 sg13g2_fill_2 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_fill_2 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_87 ();
 sg13g2_decap_8 FILLER_20_124 ();
 sg13g2_decap_8 FILLER_20_131 ();
 sg13g2_decap_4 FILLER_20_138 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_decap_8 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_155 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_175 ();
 sg13g2_fill_1 FILLER_20_177 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_decap_8 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_197 ();
 sg13g2_decap_4 FILLER_20_224 ();
 sg13g2_fill_2 FILLER_20_228 ();
 sg13g2_fill_1 FILLER_20_235 ();
 sg13g2_fill_2 FILLER_20_253 ();
 sg13g2_fill_1 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_fill_1 FILLER_20_334 ();
 sg13g2_decap_4 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_fill_2 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_4 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_53 ();
 sg13g2_fill_2 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_104 ();
 sg13g2_decap_8 FILLER_21_111 ();
 sg13g2_fill_1 FILLER_21_118 ();
 sg13g2_fill_1 FILLER_21_129 ();
 sg13g2_fill_1 FILLER_21_138 ();
 sg13g2_fill_1 FILLER_21_157 ();
 sg13g2_fill_1 FILLER_21_167 ();
 sg13g2_fill_2 FILLER_21_173 ();
 sg13g2_fill_1 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_199 ();
 sg13g2_fill_1 FILLER_21_201 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_fill_2 FILLER_21_326 ();
 sg13g2_fill_1 FILLER_21_328 ();
 sg13g2_fill_2 FILLER_21_337 ();
 sg13g2_fill_1 FILLER_21_339 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_4 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_25 ();
 sg13g2_fill_2 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_95 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_127 ();
 sg13g2_decap_4 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_138 ();
 sg13g2_decap_8 FILLER_22_148 ();
 sg13g2_fill_1 FILLER_22_155 ();
 sg13g2_fill_2 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_decap_4 FILLER_22_222 ();
 sg13g2_fill_2 FILLER_22_226 ();
 sg13g2_fill_1 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_265 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_4 FILLER_22_334 ();
 sg13g2_fill_1 FILLER_22_338 ();
 sg13g2_fill_1 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_2 FILLER_22_377 ();
 sg13g2_fill_1 FILLER_22_379 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_62 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_fill_2 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_175 ();
 sg13g2_fill_2 FILLER_23_189 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_305 ();
 sg13g2_fill_1 FILLER_23_307 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_decap_4 FILLER_23_336 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_fill_2 FILLER_24_104 ();
 sg13g2_fill_1 FILLER_24_122 ();
 sg13g2_decap_4 FILLER_24_153 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_fill_2 FILLER_24_363 ();
 sg13g2_fill_1 FILLER_24_365 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_fill_2 FILLER_25_67 ();
 sg13g2_fill_1 FILLER_25_69 ();
 sg13g2_fill_2 FILLER_25_79 ();
 sg13g2_fill_1 FILLER_25_81 ();
 sg13g2_fill_2 FILLER_25_106 ();
 sg13g2_decap_8 FILLER_25_113 ();
 sg13g2_decap_4 FILLER_25_134 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_decap_4 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_fill_2 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_decap_4 FILLER_25_229 ();
 sg13g2_decap_8 FILLER_25_237 ();
 sg13g2_decap_8 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_251 ();
 sg13g2_fill_2 FILLER_25_300 ();
 sg13g2_fill_1 FILLER_25_307 ();
 sg13g2_decap_4 FILLER_25_312 ();
 sg13g2_fill_1 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_353 ();
 sg13g2_fill_2 FILLER_25_385 ();
 sg13g2_fill_1 FILLER_25_387 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_46 ();
 sg13g2_fill_2 FILLER_26_74 ();
 sg13g2_fill_2 FILLER_26_104 ();
 sg13g2_fill_1 FILLER_26_132 ();
 sg13g2_fill_2 FILLER_26_176 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_fill_1 FILLER_26_217 ();
 sg13g2_fill_2 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_373 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_148 ();
 sg13g2_fill_2 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_209 ();
 sg13g2_decap_4 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_218 ();
 sg13g2_fill_1 FILLER_27_229 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_decap_8 FILLER_27_256 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_decap_4 FILLER_27_269 ();
 sg13g2_decap_8 FILLER_27_317 ();
 sg13g2_fill_1 FILLER_27_324 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_4 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_65 ();
 sg13g2_fill_1 FILLER_28_103 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_fill_2 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_199 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_fill_2 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_decap_4 FILLER_28_283 ();
 sg13g2_fill_1 FILLER_28_287 ();
 sg13g2_decap_4 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_fill_2 FILLER_28_324 ();
 sg13g2_fill_2 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_181 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_fill_1 FILLER_29_258 ();
 sg13g2_decap_8 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_302 ();
 sg13g2_fill_1 FILLER_29_313 ();
 sg13g2_decap_4 FILLER_29_338 ();
 sg13g2_fill_1 FILLER_29_342 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_46 ();
 sg13g2_fill_2 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_90 ();
 sg13g2_fill_1 FILLER_30_101 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_191 ();
 sg13g2_decap_4 FILLER_30_238 ();
 sg13g2_fill_1 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_257 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_fill_2 FILLER_31_91 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_104 ();
 sg13g2_fill_2 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_192 ();
 sg13g2_decap_4 FILLER_31_199 ();
 sg13g2_fill_2 FILLER_31_203 ();
 sg13g2_decap_4 FILLER_31_223 ();
 sg13g2_fill_2 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_258 ();
 sg13g2_fill_1 FILLER_31_263 ();
 sg13g2_decap_4 FILLER_31_269 ();
 sg13g2_decap_4 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_298 ();
 sg13g2_fill_2 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_316 ();
 sg13g2_fill_1 FILLER_31_320 ();
 sg13g2_fill_2 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_53 ();
 sg13g2_fill_2 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_92 ();
 sg13g2_fill_2 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_111 ();
 sg13g2_fill_1 FILLER_32_121 ();
 sg13g2_decap_4 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_decap_4 FILLER_32_175 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_decap_4 FILLER_32_185 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_decap_4 FILLER_32_208 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_4 FILLER_32_241 ();
 sg13g2_fill_1 FILLER_32_245 ();
 sg13g2_decap_4 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_274 ();
 sg13g2_fill_1 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_320 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_380 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_70 ();
 sg13g2_fill_2 FILLER_33_109 ();
 sg13g2_decap_4 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_163 ();
 sg13g2_fill_2 FILLER_33_172 ();
 sg13g2_fill_2 FILLER_33_184 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_219 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_decap_8 FILLER_33_257 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_317 ();
 sg13g2_decap_8 FILLER_33_324 ();
 sg13g2_fill_2 FILLER_33_356 ();
 sg13g2_fill_1 FILLER_33_367 ();
 sg13g2_fill_2 FILLER_33_378 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_fill_1 FILLER_34_56 ();
 sg13g2_fill_1 FILLER_34_170 ();
 sg13g2_fill_2 FILLER_34_177 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_fill_1 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_decap_4 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_295 ();
 sg13g2_decap_4 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_310 ();
 sg13g2_fill_1 FILLER_34_312 ();
 sg13g2_decap_4 FILLER_34_326 ();
 sg13g2_fill_2 FILLER_34_330 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_decap_4 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_86 ();
 sg13g2_fill_2 FILLER_35_96 ();
 sg13g2_fill_1 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_103 ();
 sg13g2_decap_4 FILLER_35_110 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_fill_1 FILLER_35_123 ();
 sg13g2_fill_1 FILLER_35_129 ();
 sg13g2_fill_2 FILLER_35_144 ();
 sg13g2_decap_8 FILLER_35_155 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_decap_4 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_234 ();
 sg13g2_decap_4 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_2 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_128 ();
 sg13g2_decap_8 FILLER_36_132 ();
 sg13g2_decap_8 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_146 ();
 sg13g2_decap_8 FILLER_36_153 ();
 sg13g2_decap_8 FILLER_36_160 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_decap_8 FILLER_36_178 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_193 ();
 sg13g2_fill_2 FILLER_36_200 ();
 sg13g2_decap_8 FILLER_36_211 ();
 sg13g2_decap_8 FILLER_36_218 ();
 sg13g2_decap_8 FILLER_36_225 ();
 sg13g2_decap_8 FILLER_36_232 ();
 sg13g2_decap_8 FILLER_36_239 ();
 sg13g2_decap_8 FILLER_36_246 ();
 sg13g2_decap_4 FILLER_36_253 ();
 sg13g2_decap_8 FILLER_36_292 ();
 sg13g2_decap_4 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_fill_2 FILLER_36_318 ();
 sg13g2_fill_2 FILLER_36_325 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_362 ();
 sg13g2_decap_8 FILLER_36_369 ();
 sg13g2_decap_8 FILLER_36_376 ();
 sg13g2_decap_8 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_4 FILLER_37_252 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_276 ();
 sg13g2_decap_8 FILLER_37_283 ();
 sg13g2_fill_2 FILLER_37_290 ();
 sg13g2_fill_2 FILLER_37_295 ();
 sg13g2_fill_1 FILLER_37_304 ();
 sg13g2_fill_1 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_131 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_155 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_decap_8 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_171 ();
 sg13g2_decap_4 FILLER_38_178 ();
 sg13g2_fill_2 FILLER_38_182 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_decap_4 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_decap_4 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_253 ();
 sg13g2_decap_4 FILLER_38_260 ();
 sg13g2_decap_4 FILLER_38_268 ();
 sg13g2_decap_8 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_283 ();
 sg13g2_fill_1 FILLER_38_285 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_decap_4 FILLER_38_323 ();
 sg13g2_fill_2 FILLER_38_327 ();
 sg13g2_decap_8 FILLER_38_355 ();
 sg13g2_decap_4 FILLER_38_362 ();
 sg13g2_fill_2 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net22;
 assign uio_oe[1] = net23;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net24;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net25;
 assign uio_oe[7] = net9;
 assign uio_out[2] = net10;
 assign uio_out[4] = net11;
 assign uio_out[5] = net12;
 assign uio_out[7] = net13;
 assign uo_out[0] = net14;
 assign uo_out[1] = net15;
 assign uo_out[2] = net16;
 assign uo_out[3] = net17;
 assign uo_out[4] = net18;
 assign uo_out[5] = net19;
 assign uo_out[6] = net20;
 assign uo_out[7] = net21;
endmodule

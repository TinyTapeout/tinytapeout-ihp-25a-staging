module tt_um_10_vga_crossyroad (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire net20;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire clknet_0_clk;
 wire \game1.hsync ;
 wire \game1.move_h ;
 wire \game1.move_v ;
 wire \game1.obstacle1_x[1] ;
 wire \game1.obstacle1_x[2] ;
 wire \game1.obstacle1_x[3] ;
 wire \game1.obstacle1_x[4] ;
 wire \game1.obstacle1_x[5] ;
 wire \game1.obstacle1_x[6] ;
 wire \game1.obstacle1_x[7] ;
 wire \game1.obstacle1_x[8] ;
 wire \game1.obstacle1_x[9] ;
 wire \game1.obstacle1_y[1] ;
 wire \game1.obstacle1_y[2] ;
 wire \game1.obstacle1_y[3] ;
 wire \game1.obstacle1_y[4] ;
 wire \game1.obstacle1_y[5] ;
 wire \game1.obstacle1_y[6] ;
 wire \game1.obstacle1_y[7] ;
 wire \game1.obstacle1_y[8] ;
 wire \game1.obstacle1_y[9] ;
 wire \game1.obstacle2_x[1] ;
 wire \game1.obstacle2_x[2] ;
 wire \game1.obstacle2_x[3] ;
 wire \game1.obstacle2_x[4] ;
 wire \game1.obstacle2_x[5] ;
 wire \game1.obstacle2_x[6] ;
 wire \game1.obstacle2_x[7] ;
 wire \game1.obstacle2_x[8] ;
 wire \game1.obstacle2_x[9] ;
 wire \game1.obstacle2_y[1] ;
 wire \game1.obstacle2_y[2] ;
 wire \game1.obstacle2_y[3] ;
 wire \game1.obstacle2_y[4] ;
 wire \game1.obstacle2_y[5] ;
 wire \game1.obstacle2_y[6] ;
 wire \game1.obstacle2_y[7] ;
 wire \game1.obstacle2_y[8] ;
 wire \game1.obstacle2_y[9] ;
 wire \game1.obstacle3_x[1] ;
 wire \game1.obstacle3_x[2] ;
 wire \game1.obstacle3_x[3] ;
 wire \game1.obstacle3_x[4] ;
 wire \game1.obstacle3_x[5] ;
 wire \game1.obstacle3_x[6] ;
 wire \game1.obstacle3_x[7] ;
 wire \game1.obstacle3_x[8] ;
 wire \game1.obstacle3_x[9] ;
 wire \game1.obstacle3_y[1] ;
 wire \game1.obstacle3_y[2] ;
 wire \game1.obstacle3_y[3] ;
 wire \game1.obstacle3_y[4] ;
 wire \game1.obstacle3_y[5] ;
 wire \game1.obstacle3_y[6] ;
 wire \game1.obstacle3_y[7] ;
 wire \game1.obstacle3_y[8] ;
 wire \game1.obstacle3_y[9] ;
 wire \game1.pixel_x[0] ;
 wire \game1.pixel_x[1] ;
 wire \game1.pixel_x[2] ;
 wire \game1.pixel_x[3] ;
 wire \game1.pixel_x[4] ;
 wire \game1.pixel_x[5] ;
 wire \game1.pixel_x[6] ;
 wire \game1.pixel_x[7] ;
 wire \game1.pixel_x[8] ;
 wire \game1.pixel_x[9] ;
 wire \game1.pixel_y[0] ;
 wire \game1.pixel_y[1] ;
 wire \game1.pixel_y[2] ;
 wire \game1.pixel_y[3] ;
 wire \game1.pixel_y[4] ;
 wire \game1.pixel_y[5] ;
 wire \game1.pixel_y[6] ;
 wire \game1.pixel_y[7] ;
 wire \game1.pixel_y[8] ;
 wire \game1.pixel_y[9] ;
 wire \game1.score[0] ;
 wire \game1.score[1] ;
 wire \game1.score[2] ;
 wire \game1.score[3] ;
 wire \game1.score[4] ;
 wire \game1.score[5] ;
 wire \game1.score[6] ;
 wire \game1.score_inst.o_score_rgb[0] ;
 wire \game1.scroll1_h_inst.ctr[0] ;
 wire \game1.scroll1_h_inst.ctr[10] ;
 wire \game1.scroll1_h_inst.ctr[11] ;
 wire \game1.scroll1_h_inst.ctr[12] ;
 wire \game1.scroll1_h_inst.ctr[13] ;
 wire \game1.scroll1_h_inst.ctr[14] ;
 wire \game1.scroll1_h_inst.ctr[15] ;
 wire \game1.scroll1_h_inst.ctr[16] ;
 wire \game1.scroll1_h_inst.ctr[17] ;
 wire \game1.scroll1_h_inst.ctr[1] ;
 wire \game1.scroll1_h_inst.ctr[2] ;
 wire \game1.scroll1_h_inst.ctr[3] ;
 wire \game1.scroll1_h_inst.ctr[4] ;
 wire \game1.scroll1_h_inst.ctr[5] ;
 wire \game1.scroll1_h_inst.ctr[6] ;
 wire \game1.scroll1_h_inst.ctr[7] ;
 wire \game1.scroll1_h_inst.ctr[8] ;
 wire \game1.scroll1_h_inst.ctr[9] ;
 wire \game1.scroll1_v_inst.ctr[0] ;
 wire \game1.scroll1_v_inst.ctr[10] ;
 wire \game1.scroll1_v_inst.ctr[11] ;
 wire \game1.scroll1_v_inst.ctr[12] ;
 wire \game1.scroll1_v_inst.ctr[13] ;
 wire \game1.scroll1_v_inst.ctr[14] ;
 wire \game1.scroll1_v_inst.ctr[15] ;
 wire \game1.scroll1_v_inst.ctr[16] ;
 wire \game1.scroll1_v_inst.ctr[17] ;
 wire \game1.scroll1_v_inst.ctr[1] ;
 wire \game1.scroll1_v_inst.ctr[2] ;
 wire \game1.scroll1_v_inst.ctr[3] ;
 wire \game1.scroll1_v_inst.ctr[4] ;
 wire \game1.scroll1_v_inst.ctr[5] ;
 wire \game1.scroll1_v_inst.ctr[6] ;
 wire \game1.scroll1_v_inst.ctr[7] ;
 wire \game1.scroll1_v_inst.ctr[8] ;
 wire \game1.scroll1_v_inst.ctr[9] ;
 wire \game1.scroll1_v_inst.score_ctr[0] ;
 wire \game1.scroll1_v_inst.score_ctr[1] ;
 wire \game1.scroll1_v_inst.score_ctr[2] ;
 wire \game1.scroll1_v_inst.score_ctr[3] ;
 wire \game1.scroll1_v_inst.score_ctr[4] ;
 wire \game1.scroll1_v_inst.score_ctr[5] ;
 wire \game1.scroll1_v_inst.score_ctr[6] ;
 wire \game1.vga_inst.vsync ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;

 sg13g2_inv_1 _1349_ (.Y(_0500_),
    .A(net387));
 sg13g2_inv_2 _1350_ (.Y(_0501_),
    .A(net2));
 sg13g2_inv_1 _1351_ (.Y(_0502_),
    .A(\game1.scroll1_v_inst.ctr[5] ));
 sg13g2_inv_1 _1352_ (.Y(_0503_),
    .A(\game1.score[4] ));
 sg13g2_inv_1 _1353_ (.Y(_0504_),
    .A(\game1.score[3] ));
 sg13g2_inv_1 _1354_ (.Y(_0505_),
    .A(\game1.obstacle2_y[9] ));
 sg13g2_inv_1 _1355_ (.Y(_0506_),
    .A(net165));
 sg13g2_inv_1 _1356_ (.Y(_0507_),
    .A(\game1.obstacle2_y[8] ));
 sg13g2_inv_1 _1357_ (.Y(_0508_),
    .A(\game1.obstacle2_y[7] ));
 sg13g2_inv_1 _1358_ (.Y(_0509_),
    .A(\game1.obstacle2_y[6] ));
 sg13g2_inv_1 _1359_ (.Y(_0510_),
    .A(\game1.obstacle2_y[5] ));
 sg13g2_inv_1 _1360_ (.Y(_0511_),
    .A(\game1.obstacle2_y[4] ));
 sg13g2_inv_1 _1361_ (.Y(_0512_),
    .A(net183));
 sg13g2_inv_1 _1362_ (.Y(_0513_),
    .A(\game1.obstacle1_x[8] ));
 sg13g2_inv_1 _1363_ (.Y(_0514_),
    .A(\game1.obstacle1_x[6] ));
 sg13g2_inv_1 _1364_ (.Y(_0515_),
    .A(\game1.obstacle1_x[4] ));
 sg13g2_inv_1 _1365_ (.Y(_0516_),
    .A(\game1.obstacle2_x[9] ));
 sg13g2_inv_2 _1366_ (.Y(_0517_),
    .A(net257));
 sg13g2_inv_1 _1367_ (.Y(_0518_),
    .A(\game1.obstacle2_x[8] ));
 sg13g2_inv_2 _1368_ (.Y(_0519_),
    .A(net415));
 sg13g2_inv_1 _1369_ (.Y(_0520_),
    .A(\game1.obstacle2_x[3] ));
 sg13g2_inv_1 _1370_ (.Y(_0521_),
    .A(\game1.obstacle2_x[1] ));
 sg13g2_inv_1 _1371_ (.Y(_0522_),
    .A(net286));
 sg13g2_inv_1 _1372_ (.Y(_0523_),
    .A(net317));
 sg13g2_inv_1 _1373_ (.Y(_0524_),
    .A(\game1.obstacle1_y[7] ));
 sg13g2_inv_1 _1374_ (.Y(_0525_),
    .A(\game1.obstacle1_y[6] ));
 sg13g2_inv_1 _1375_ (.Y(_0526_),
    .A(net310));
 sg13g2_inv_1 _1376_ (.Y(_0527_),
    .A(net287));
 sg13g2_inv_1 _1377_ (.Y(_0528_),
    .A(net348));
 sg13g2_inv_1 _1378_ (.Y(_0529_),
    .A(\game1.obstacle3_x[9] ));
 sg13g2_inv_1 _1379_ (.Y(_0530_),
    .A(\game1.obstacle3_x[8] ));
 sg13g2_inv_1 _1380_ (.Y(_0531_),
    .A(\game1.obstacle3_x[7] ));
 sg13g2_inv_1 _1381_ (.Y(_0532_),
    .A(net426));
 sg13g2_inv_1 _1382_ (.Y(_0533_),
    .A(net402));
 sg13g2_inv_1 _1383_ (.Y(_0534_),
    .A(net398));
 sg13g2_inv_1 _1384_ (.Y(_0535_),
    .A(net185));
 sg13g2_inv_1 _1385_ (.Y(_0536_),
    .A(\game1.obstacle3_y[8] ));
 sg13g2_inv_1 _1386_ (.Y(_0537_),
    .A(\game1.obstacle3_y[7] ));
 sg13g2_inv_1 _1387_ (.Y(_0538_),
    .A(\game1.obstacle3_y[6] ));
 sg13g2_inv_1 _1388_ (.Y(_0539_),
    .A(\game1.obstacle3_y[5] ));
 sg13g2_inv_1 _1389_ (.Y(_0540_),
    .A(\game1.obstacle3_y[4] ));
 sg13g2_inv_1 _1390_ (.Y(_0541_),
    .A(net1));
 sg13g2_inv_1 _1391_ (.Y(_0542_),
    .A(\game1.pixel_x[1] ));
 sg13g2_inv_2 _1392_ (.Y(_0543_),
    .A(net265));
 sg13g2_inv_2 _1393_ (.Y(_0544_),
    .A(net267));
 sg13g2_inv_2 _1394_ (.Y(_0545_),
    .A(net269));
 sg13g2_inv_4 _1395_ (.A(net271),
    .Y(_0546_));
 sg13g2_inv_1 _1396_ (.Y(_0547_),
    .A(net261));
 sg13g2_inv_2 _1397_ (.Y(_0548_),
    .A(\game1.pixel_x[8] ));
 sg13g2_inv_1 _1398_ (.Y(_0549_),
    .A(_0021_));
 sg13g2_inv_1 _1399_ (.Y(_0550_),
    .A(net250));
 sg13g2_inv_4 _1400_ (.A(net247),
    .Y(_0551_));
 sg13g2_inv_2 _1401_ (.Y(_0552_),
    .A(net249));
 sg13g2_inv_2 _1402_ (.Y(_0553_),
    .A(net239));
 sg13g2_inv_2 _1403_ (.Y(_0554_),
    .A(net241));
 sg13g2_inv_2 _1404_ (.Y(_0555_),
    .A(net243));
 sg13g2_inv_2 _1405_ (.Y(_0556_),
    .A(net245));
 sg13g2_inv_2 _1406_ (.Y(_0557_),
    .A(net237));
 sg13g2_inv_2 _1407_ (.Y(_0558_),
    .A(net238));
 sg13g2_inv_1 _1408_ (.Y(_0559_),
    .A(net388));
 sg13g2_inv_1 _1409_ (.Y(_0560_),
    .A(_0006_));
 sg13g2_inv_1 _1410_ (.Y(_0561_),
    .A(net355));
 sg13g2_inv_1 _1411_ (.Y(_0562_),
    .A(net405));
 sg13g2_inv_1 _1412_ (.Y(_0563_),
    .A(_0009_));
 sg13g2_inv_1 _1413_ (.Y(_0564_),
    .A(\game1.score_inst.o_score_rgb[0] ));
 sg13g2_nand2_1 _1414_ (.Y(_0565_),
    .A(net261),
    .B(net263));
 sg13g2_nand3_1 _1415_ (.B(_0545_),
    .C(_0546_),
    .A(_0544_),
    .Y(_0566_));
 sg13g2_nand3_1 _1416_ (.B(net261),
    .C(_0566_),
    .A(net264),
    .Y(_0567_));
 sg13g2_nand2_1 _1417_ (.Y(_0568_),
    .A(net269),
    .B(net272));
 sg13g2_nand2_2 _1418_ (.Y(_0569_),
    .A(net267),
    .B(net269));
 sg13g2_nand4_1 _1419_ (.B(net267),
    .C(net268),
    .A(net264),
    .Y(_0570_),
    .D(net271));
 sg13g2_nor2_1 _1420_ (.A(net234),
    .B(net263),
    .Y(_0571_));
 sg13g2_a21oi_1 _1421_ (.A1(_0570_),
    .A2(_0571_),
    .Y(_0572_),
    .B1(net423));
 sg13g2_a21oi_2 _1422_ (.B1(_0572_),
    .Y(_0000_),
    .A2(_0567_),
    .A1(_0565_));
 sg13g2_nand2_2 _1423_ (.Y(_0573_),
    .A(net240),
    .B(net242));
 sg13g2_nor2_1 _1424_ (.A(_0030_),
    .B(_0573_),
    .Y(_0574_));
 sg13g2_nand2_1 _1425_ (.Y(_0575_),
    .A(net244),
    .B(_0556_));
 sg13g2_and2_2 _1426_ (.A(net250),
    .B(\game1.pixel_y[0] ),
    .X(_0576_));
 sg13g2_nor2_1 _1427_ (.A(net248),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_nor2_2 _1428_ (.A(_0551_),
    .B(_0552_),
    .Y(_0578_));
 sg13g2_o21ai_1 _1429_ (.B1(net246),
    .Y(_0579_),
    .A1(net248),
    .A2(_0576_));
 sg13g2_nand2b_1 _1430_ (.Y(_0580_),
    .B(_0579_),
    .A_N(_0575_));
 sg13g2_nor2_2 _1431_ (.A(_0550_),
    .B(\game1.pixel_y[0] ),
    .Y(_0581_));
 sg13g2_nand2_1 _1432_ (.Y(_0582_),
    .A(net246),
    .B(_0581_));
 sg13g2_nor4_1 _1433_ (.A(net248),
    .B(_0573_),
    .C(_0575_),
    .D(_0582_),
    .Y(_0583_));
 sg13g2_a21oi_1 _1434_ (.A1(_0574_),
    .A2(_0580_),
    .Y(_0584_),
    .B1(_0583_));
 sg13g2_nor2_1 _1435_ (.A(net245),
    .B(_0578_),
    .Y(_0585_));
 sg13g2_nor2_1 _1436_ (.A(_0555_),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_nand2_1 _1437_ (.Y(_0587_),
    .A(_0557_),
    .B(net281));
 sg13g2_nor2_1 _1438_ (.A(_0573_),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_nor4_2 _1439_ (.A(_0573_),
    .B(_0584_),
    .C(_0586_),
    .Y(_0001_),
    .D(_0587_));
 sg13g2_nor3_1 _1440_ (.A(net246),
    .B(net248),
    .C(net245),
    .Y(_0589_));
 sg13g2_nor2_1 _1441_ (.A(net250),
    .B(\game1.pixel_y[0] ),
    .Y(_0590_));
 sg13g2_or2_1 _1442_ (.X(_0591_),
    .B(\game1.pixel_y[0] ),
    .A(net251));
 sg13g2_nor4_1 _1443_ (.A(net246),
    .B(net248),
    .C(_0575_),
    .D(_0591_),
    .Y(_0592_));
 sg13g2_nor2_2 _1444_ (.A(net265),
    .B(\game1.pixel_x[8] ),
    .Y(_0593_));
 sg13g2_or2_1 _1445_ (.X(_0594_),
    .B(\game1.pixel_x[8] ),
    .A(net265));
 sg13g2_o21ai_1 _1446_ (.B1(_0557_),
    .Y(_0595_),
    .A1(_0018_),
    .A2(_0593_));
 sg13g2_a22oi_1 _1447_ (.Y(_0596_),
    .B1(_0588_),
    .B2(_0592_),
    .A2(_0574_),
    .A1(net238));
 sg13g2_nand2b_2 _1448_ (.Y(_0597_),
    .B(_0596_),
    .A_N(_0595_));
 sg13g2_o21ai_1 _1449_ (.B1(\game1.obstacle3_y[3] ),
    .Y(_0598_),
    .A1(\game1.obstacle3_y[2] ),
    .A2(net279));
 sg13g2_nor2_1 _1450_ (.A(_0540_),
    .B(_0598_),
    .Y(_0599_));
 sg13g2_nand2_1 _1451_ (.Y(_0600_),
    .A(\game1.obstacle3_y[5] ),
    .B(_0599_));
 sg13g2_nand2_1 _1452_ (.Y(_0601_),
    .A(\game1.obstacle3_y[8] ),
    .B(\game1.obstacle3_y[7] ));
 sg13g2_a21o_1 _1453_ (.A2(_0600_),
    .A1(_0538_),
    .B1(_0601_),
    .X(_0602_));
 sg13g2_nor2_1 _1454_ (.A(_0014_),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_xnor2_1 _1455_ (.Y(_0604_),
    .A(_0535_),
    .B(_0602_));
 sg13g2_nand2_1 _1456_ (.Y(_0605_),
    .A(net237),
    .B(_0604_));
 sg13g2_nor3_1 _1457_ (.A(_0540_),
    .B(_0013_),
    .C(_0598_),
    .Y(_0606_));
 sg13g2_xnor2_1 _1458_ (.Y(_0607_),
    .A(\game1.obstacle3_y[6] ),
    .B(_0606_));
 sg13g2_inv_1 _1459_ (.Y(_0608_),
    .A(_0607_));
 sg13g2_xor2_1 _1460_ (.B(_0599_),
    .A(_0013_),
    .X(_0609_));
 sg13g2_nand2_1 _1461_ (.Y(_0610_),
    .A(net243),
    .B(_0609_));
 sg13g2_xnor2_1 _1462_ (.Y(_0611_),
    .A(\game1.obstacle3_y[4] ),
    .B(_0598_));
 sg13g2_nor2_1 _1463_ (.A(_0031_),
    .B(_0611_),
    .Y(_0612_));
 sg13g2_or3_1 _1464_ (.A(\game1.obstacle3_y[3] ),
    .B(\game1.obstacle3_y[2] ),
    .C(\game1.obstacle3_y[1] ),
    .X(_0613_));
 sg13g2_nand2_1 _1465_ (.Y(_0614_),
    .A(_0598_),
    .B(_0613_));
 sg13g2_nor2_1 _1466_ (.A(net247),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_xor2_1 _1467_ (.B(net279),
    .A(\game1.obstacle3_y[2] ),
    .X(_0616_));
 sg13g2_xnor2_1 _1468_ (.Y(_0617_),
    .A(_0032_),
    .B(_0616_));
 sg13g2_o21ai_1 _1469_ (.B1(_0617_),
    .Y(_0618_),
    .A1(net279),
    .A2(net250));
 sg13g2_a22oi_1 _1470_ (.Y(_0619_),
    .B1(_0616_),
    .B2(net249),
    .A2(_0614_),
    .A1(net247));
 sg13g2_a21oi_1 _1471_ (.A1(_0618_),
    .A2(_0619_),
    .Y(_0620_),
    .B1(_0615_));
 sg13g2_and2_1 _1472_ (.A(_0031_),
    .B(_0611_),
    .X(_0621_));
 sg13g2_xnor2_1 _1473_ (.Y(_0622_),
    .A(_0030_),
    .B(_0609_));
 sg13g2_o21ai_1 _1474_ (.B1(_0622_),
    .Y(_0623_),
    .A1(_0612_),
    .A2(_0620_));
 sg13g2_o21ai_1 _1475_ (.B1(_0610_),
    .Y(_0624_),
    .A1(_0621_),
    .A2(_0623_));
 sg13g2_xor2_1 _1476_ (.B(_0607_),
    .A(_0029_),
    .X(_0625_));
 sg13g2_a22oi_1 _1477_ (.Y(_0626_),
    .B1(_0624_),
    .B2(_0625_),
    .A2(_0608_),
    .A1(net241));
 sg13g2_o21ai_1 _1478_ (.B1(_0012_),
    .Y(_0627_),
    .A1(\game1.obstacle3_y[6] ),
    .A2(_0600_));
 sg13g2_nand2_1 _1479_ (.Y(_0628_),
    .A(\game1.obstacle3_y[7] ),
    .B(_0627_));
 sg13g2_xnor2_1 _1480_ (.Y(_0629_),
    .A(_0537_),
    .B(_0627_));
 sg13g2_a21oi_1 _1481_ (.A1(_0553_),
    .A2(_0629_),
    .Y(_0630_),
    .B1(_0626_));
 sg13g2_xor2_1 _1482_ (.B(_0628_),
    .A(_0015_),
    .X(_0631_));
 sg13g2_nand2b_1 _1483_ (.Y(_0632_),
    .B(net239),
    .A_N(_0629_));
 sg13g2_o21ai_1 _1484_ (.B1(_0632_),
    .Y(_0633_),
    .A1(_0025_),
    .A2(_0631_));
 sg13g2_xor2_1 _1485_ (.B(_0604_),
    .A(_0024_),
    .X(_0634_));
 sg13g2_a21oi_1 _1486_ (.A1(_0025_),
    .A2(_0631_),
    .Y(_0635_),
    .B1(_0634_));
 sg13g2_o21ai_1 _1487_ (.B1(_0635_),
    .Y(_0636_),
    .A1(_0630_),
    .A2(_0633_));
 sg13g2_a21oi_1 _1488_ (.A1(_0605_),
    .A2(_0636_),
    .Y(_0637_),
    .B1(_0603_));
 sg13g2_nor3_2 _1489_ (.A(net402),
    .B(\game1.obstacle3_x[4] ),
    .C(\game1.obstacle3_x[3] ),
    .Y(_0638_));
 sg13g2_nand2_2 _1490_ (.Y(_0639_),
    .A(_0532_),
    .B(_0638_));
 sg13g2_and3_1 _1491_ (.X(_0640_),
    .A(\game1.obstacle3_x[8] ),
    .B(\game1.obstacle3_x[7] ),
    .C(_0639_));
 sg13g2_xor2_1 _1492_ (.B(_0640_),
    .A(_0016_),
    .X(_0641_));
 sg13g2_xnor2_1 _1493_ (.Y(_0642_),
    .A(\game1.obstacle3_x[7] ),
    .B(_0639_));
 sg13g2_xnor2_1 _1494_ (.Y(_0643_),
    .A(\game1.obstacle3_x[6] ),
    .B(_0638_));
 sg13g2_nand2_1 _1495_ (.Y(_0644_),
    .A(net267),
    .B(_0643_));
 sg13g2_o21ai_1 _1496_ (.B1(\game1.obstacle3_x[5] ),
    .Y(_0645_),
    .A1(\game1.obstacle3_x[4] ),
    .A2(net278));
 sg13g2_nor2b_1 _1497_ (.A(_0638_),
    .B_N(_0645_),
    .Y(_0646_));
 sg13g2_nor2b_1 _1498_ (.A(net276),
    .B_N(\game1.obstacle3_x[2] ),
    .Y(_0647_));
 sg13g2_nand2b_1 _1499_ (.Y(_0648_),
    .B(net276),
    .A_N(\game1.obstacle3_x[2] ));
 sg13g2_nor2b_1 _1500_ (.A(\game1.pixel_x[1] ),
    .B_N(\game1.obstacle3_x[1] ),
    .Y(_0649_));
 sg13g2_o21ai_1 _1501_ (.B1(_0648_),
    .Y(_0650_),
    .A1(_0647_),
    .A2(_0649_));
 sg13g2_o21ai_1 _1502_ (.B1(net278),
    .Y(_0651_),
    .A1(net275),
    .A2(_0650_));
 sg13g2_xnor2_1 _1503_ (.Y(_0652_),
    .A(\game1.obstacle3_x[4] ),
    .B(net278));
 sg13g2_nor2_1 _1504_ (.A(net270),
    .B(_0652_),
    .Y(_0653_));
 sg13g2_a21oi_1 _1505_ (.A1(net275),
    .A2(_0650_),
    .Y(_0654_),
    .B1(_0653_));
 sg13g2_xnor2_1 _1506_ (.Y(_0655_),
    .A(_0021_),
    .B(_0646_));
 sg13g2_a22oi_1 _1507_ (.Y(_0656_),
    .B1(_0654_),
    .B2(_0651_),
    .A2(_0652_),
    .A1(net270));
 sg13g2_a22oi_1 _1508_ (.Y(_0657_),
    .B1(_0655_),
    .B2(_0656_),
    .A2(_0646_),
    .A1(net268));
 sg13g2_xor2_1 _1509_ (.B(_0643_),
    .A(_0020_),
    .X(_0658_));
 sg13g2_o21ai_1 _1510_ (.B1(_0644_),
    .Y(_0659_),
    .A1(_0657_),
    .A2(_0658_));
 sg13g2_o21ai_1 _1511_ (.B1(_0659_),
    .Y(_0660_),
    .A1(net264),
    .A2(_0642_));
 sg13g2_a21oi_1 _1512_ (.A1(\game1.obstacle3_x[7] ),
    .A2(_0639_),
    .Y(_0661_),
    .B1(\game1.obstacle3_x[8] ));
 sg13g2_nor2_1 _1513_ (.A(_0640_),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_nor2_1 _1514_ (.A(_0019_),
    .B(_0662_),
    .Y(_0663_));
 sg13g2_a21oi_1 _1515_ (.A1(net264),
    .A2(_0642_),
    .Y(_0664_),
    .B1(_0663_));
 sg13g2_xor2_1 _1516_ (.B(_0641_),
    .A(_0018_),
    .X(_0665_));
 sg13g2_a221oi_1 _1517_ (.B2(_0660_),
    .C1(_0665_),
    .B1(_0664_),
    .A1(_0019_),
    .Y(_0666_),
    .A2(_0662_));
 sg13g2_a21oi_1 _1518_ (.A1(net261),
    .A2(_0641_),
    .Y(_0667_),
    .B1(_0666_));
 sg13g2_a21oi_2 _1519_ (.B1(_0667_),
    .Y(_0668_),
    .A2(_0640_),
    .A1(\game1.obstacle3_x[9] ));
 sg13g2_nand2b_1 _1520_ (.Y(_0669_),
    .B(net278),
    .A_N(net275));
 sg13g2_nor2b_1 _1521_ (.A(net278),
    .B_N(net275),
    .Y(_0670_));
 sg13g2_a221oi_1 _1522_ (.B2(_0669_),
    .C1(_0670_),
    .B1(_0650_),
    .A1(_0534_),
    .Y(_0671_),
    .A2(net271));
 sg13g2_a221oi_1 _1523_ (.B2(\game1.obstacle3_x[4] ),
    .C1(_0671_),
    .B1(_0546_),
    .A1(\game1.obstacle3_x[5] ),
    .Y(_0672_),
    .A2(_0545_));
 sg13g2_a221oi_1 _1524_ (.B2(_0533_),
    .C1(_0672_),
    .B1(net268),
    .A1(_0532_),
    .Y(_0673_),
    .A2(net267));
 sg13g2_a221oi_1 _1525_ (.B2(\game1.obstacle3_x[6] ),
    .C1(_0673_),
    .B1(_0544_),
    .A1(\game1.obstacle3_x[7] ),
    .Y(_0674_),
    .A2(_0543_));
 sg13g2_a221oi_1 _1526_ (.B2(_0530_),
    .C1(_0674_),
    .B1(net263),
    .A1(_0531_),
    .Y(_0675_),
    .A2(net264));
 sg13g2_a221oi_1 _1527_ (.B2(\game1.obstacle3_x[8] ),
    .C1(_0675_),
    .B1(_0548_),
    .A1(\game1.obstacle3_x[9] ),
    .Y(_0676_),
    .A2(net234));
 sg13g2_a21oi_2 _1528_ (.B1(_0676_),
    .Y(_0677_),
    .A2(net261),
    .A1(_0529_));
 sg13g2_nor2b_1 _1529_ (.A(net250),
    .B_N(net279),
    .Y(_0678_));
 sg13g2_o21ai_1 _1530_ (.B1(_0678_),
    .Y(_0679_),
    .A1(\game1.obstacle3_y[2] ),
    .A2(_0552_));
 sg13g2_a22oi_1 _1531_ (.Y(_0680_),
    .B1(_0552_),
    .B2(\game1.obstacle3_y[2] ),
    .A2(_0551_),
    .A1(\game1.obstacle3_y[3] ));
 sg13g2_nor2_1 _1532_ (.A(\game1.obstacle3_y[3] ),
    .B(_0551_),
    .Y(_0681_));
 sg13g2_a221oi_1 _1533_ (.B2(_0680_),
    .C1(_0681_),
    .B1(_0679_),
    .A1(_0540_),
    .Y(_0682_),
    .A2(net245));
 sg13g2_a221oi_1 _1534_ (.B2(\game1.obstacle3_y[4] ),
    .C1(_0682_),
    .B1(_0556_),
    .A1(\game1.obstacle3_y[5] ),
    .Y(_0683_),
    .A2(_0555_));
 sg13g2_a221oi_1 _1535_ (.B2(_0539_),
    .C1(_0683_),
    .B1(net243),
    .A1(_0538_),
    .Y(_0684_),
    .A2(net241));
 sg13g2_a221oi_1 _1536_ (.B2(\game1.obstacle3_y[6] ),
    .C1(_0684_),
    .B1(_0554_),
    .A1(\game1.obstacle3_y[7] ),
    .Y(_0685_),
    .A2(_0553_));
 sg13g2_a221oi_1 _1537_ (.B2(_0536_),
    .C1(_0685_),
    .B1(net238),
    .A1(_0537_),
    .Y(_0686_),
    .A2(net239));
 sg13g2_a221oi_1 _1538_ (.B2(\game1.obstacle3_y[8] ),
    .C1(_0686_),
    .B1(_0558_),
    .A1(\game1.obstacle3_y[9] ),
    .Y(_0687_),
    .A2(_0557_));
 sg13g2_a21oi_1 _1539_ (.A1(_0535_),
    .A2(net237),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_nor4_2 _1540_ (.A(_0637_),
    .B(_0668_),
    .C(_0677_),
    .Y(_0689_),
    .D(_0688_));
 sg13g2_o21ai_1 _1541_ (.B1(\game1.obstacle2_y[3] ),
    .Y(_0690_),
    .A1(\game1.obstacle2_y[2] ),
    .A2(net256));
 sg13g2_nor2_1 _1542_ (.A(_0511_),
    .B(_0690_),
    .Y(_0691_));
 sg13g2_nand2_1 _1543_ (.Y(_0692_),
    .A(\game1.obstacle2_y[5] ),
    .B(_0691_));
 sg13g2_o21ai_1 _1544_ (.B1(_0035_),
    .Y(_0693_),
    .A1(\game1.obstacle2_y[6] ),
    .A2(_0692_));
 sg13g2_nand2_1 _1545_ (.Y(_0694_),
    .A(\game1.obstacle2_y[7] ),
    .B(_0693_));
 sg13g2_xor2_1 _1546_ (.B(_0694_),
    .A(_0034_),
    .X(_0695_));
 sg13g2_xnor2_1 _1547_ (.Y(_0696_),
    .A(\game1.obstacle2_y[7] ),
    .B(_0693_));
 sg13g2_nor3_1 _1548_ (.A(_0511_),
    .B(_0036_),
    .C(_0690_),
    .Y(_0697_));
 sg13g2_xor2_1 _1549_ (.B(_0691_),
    .A(_0036_),
    .X(_0698_));
 sg13g2_xnor2_1 _1550_ (.Y(_0699_),
    .A(\game1.obstacle2_y[4] ),
    .B(_0690_));
 sg13g2_xor2_1 _1551_ (.B(net256),
    .A(\game1.obstacle2_y[2] ),
    .X(_0700_));
 sg13g2_or2_1 _1552_ (.X(_0701_),
    .B(net250),
    .A(net256));
 sg13g2_xnor2_1 _1553_ (.Y(_0702_),
    .A(_0032_),
    .B(_0700_));
 sg13g2_or3_1 _1554_ (.A(\game1.obstacle2_y[3] ),
    .B(\game1.obstacle2_y[2] ),
    .C(net256),
    .X(_0703_));
 sg13g2_and2_1 _1555_ (.A(_0690_),
    .B(_0703_),
    .X(_0704_));
 sg13g2_nor2_1 _1556_ (.A(_0551_),
    .B(_0704_),
    .Y(_0705_));
 sg13g2_a221oi_1 _1557_ (.B2(_0702_),
    .C1(_0705_),
    .B1(_0701_),
    .A1(net249),
    .Y(_0706_),
    .A2(_0700_));
 sg13g2_a22oi_1 _1558_ (.Y(_0707_),
    .B1(_0704_),
    .B2(_0551_),
    .A2(_0699_),
    .A1(_0031_));
 sg13g2_nand2b_1 _1559_ (.Y(_0708_),
    .B(_0707_),
    .A_N(_0706_));
 sg13g2_o21ai_1 _1560_ (.B1(_0708_),
    .Y(_0709_),
    .A1(_0031_),
    .A2(_0699_));
 sg13g2_xnor2_1 _1561_ (.Y(_0710_),
    .A(_0030_),
    .B(_0698_));
 sg13g2_a22oi_1 _1562_ (.Y(_0711_),
    .B1(_0709_),
    .B2(_0710_),
    .A2(_0698_),
    .A1(net243));
 sg13g2_xnor2_1 _1563_ (.Y(_0712_),
    .A(\game1.obstacle2_y[6] ),
    .B(_0697_));
 sg13g2_xnor2_1 _1564_ (.Y(_0713_),
    .A(_0029_),
    .B(_0712_));
 sg13g2_nor2_1 _1565_ (.A(_0554_),
    .B(_0712_),
    .Y(_0714_));
 sg13g2_a21oi_1 _1566_ (.A1(net239),
    .A2(_0696_),
    .Y(_0715_),
    .B1(_0714_));
 sg13g2_o21ai_1 _1567_ (.B1(_0715_),
    .Y(_0716_),
    .A1(_0711_),
    .A2(_0713_));
 sg13g2_o21ai_1 _1568_ (.B1(_0716_),
    .Y(_0717_),
    .A1(net239),
    .A2(_0696_));
 sg13g2_o21ai_1 _1569_ (.B1(_0717_),
    .Y(_0718_),
    .A1(_0025_),
    .A2(_0695_));
 sg13g2_nand2_1 _1570_ (.Y(_0719_),
    .A(_0025_),
    .B(_0695_));
 sg13g2_a21oi_1 _1571_ (.A1(\game1.obstacle2_y[5] ),
    .A2(_0691_),
    .Y(_0720_),
    .B1(\game1.obstacle2_y[6] ));
 sg13g2_nand2_1 _1572_ (.Y(_0721_),
    .A(\game1.obstacle2_y[8] ),
    .B(\game1.obstacle2_y[7] ));
 sg13g2_or3_1 _1573_ (.A(_0505_),
    .B(_0720_),
    .C(_0721_),
    .X(_0722_));
 sg13g2_o21ai_1 _1574_ (.B1(_0505_),
    .Y(_0723_),
    .A1(_0720_),
    .A2(_0721_));
 sg13g2_a21o_1 _1575_ (.A2(_0723_),
    .A1(_0722_),
    .B1(_0024_),
    .X(_0724_));
 sg13g2_nand3_1 _1576_ (.B(_0722_),
    .C(_0723_),
    .A(_0024_),
    .Y(_0725_));
 sg13g2_and4_1 _1577_ (.A(_0719_),
    .B(_0722_),
    .C(_0724_),
    .D(_0725_),
    .X(_0726_));
 sg13g2_or2_1 _1578_ (.X(_0727_),
    .B(\game1.obstacle2_x[3] ),
    .A(\game1.obstacle2_x[4] ));
 sg13g2_nor3_2 _1579_ (.A(\game1.obstacle2_x[5] ),
    .B(\game1.obstacle2_x[4] ),
    .C(\game1.obstacle2_x[3] ),
    .Y(_0728_));
 sg13g2_nand2_2 _1580_ (.Y(_0729_),
    .A(_0519_),
    .B(_0728_));
 sg13g2_nand3_1 _1581_ (.B(\game1.obstacle2_x[7] ),
    .C(_0729_),
    .A(\game1.obstacle2_x[8] ),
    .Y(_0730_));
 sg13g2_inv_1 _1582_ (.Y(_0731_),
    .A(_0730_));
 sg13g2_xor2_1 _1583_ (.B(_0730_),
    .A(_0033_),
    .X(_0732_));
 sg13g2_nor2_1 _1584_ (.A(net234),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_xor2_1 _1585_ (.B(_0729_),
    .A(net260),
    .X(_0734_));
 sg13g2_nand2_1 _1586_ (.Y(_0735_),
    .A(_0543_),
    .B(_0734_));
 sg13g2_xnor2_1 _1587_ (.Y(_0736_),
    .A(\game1.obstacle2_x[6] ),
    .B(_0728_));
 sg13g2_nand2_1 _1588_ (.Y(_0737_),
    .A(net267),
    .B(_0736_));
 sg13g2_xor2_1 _1589_ (.B(_0727_),
    .A(\game1.obstacle2_x[5] ),
    .X(_0738_));
 sg13g2_nand2b_1 _1590_ (.Y(_0739_),
    .B(net276),
    .A_N(\game1.obstacle2_x[2] ));
 sg13g2_nand3_1 _1591_ (.B(_0542_),
    .C(_0739_),
    .A(\game1.obstacle2_x[1] ),
    .Y(_0740_));
 sg13g2_nand2b_1 _1592_ (.Y(_0741_),
    .B(\game1.obstacle2_x[2] ),
    .A_N(net276));
 sg13g2_o21ai_1 _1593_ (.B1(_0741_),
    .Y(_0742_),
    .A1(\game1.obstacle2_x[3] ),
    .A2(net275));
 sg13g2_nand2b_1 _1594_ (.Y(_0743_),
    .B(_0740_),
    .A_N(_0742_));
 sg13g2_xnor2_1 _1595_ (.Y(_0744_),
    .A(\game1.obstacle2_x[4] ),
    .B(\game1.obstacle2_x[3] ));
 sg13g2_nor2_1 _1596_ (.A(net270),
    .B(_0744_),
    .Y(_0745_));
 sg13g2_a21oi_1 _1597_ (.A1(\game1.obstacle2_x[3] ),
    .A2(net275),
    .Y(_0746_),
    .B1(_0745_));
 sg13g2_xnor2_1 _1598_ (.Y(_0747_),
    .A(_0549_),
    .B(_0738_));
 sg13g2_a221oi_1 _1599_ (.B2(_0743_),
    .C1(_0747_),
    .B1(_0746_),
    .A1(net270),
    .Y(_0748_),
    .A2(_0744_));
 sg13g2_a21oi_1 _1600_ (.A1(net268),
    .A2(_0738_),
    .Y(_0749_),
    .B1(_0748_));
 sg13g2_xor2_1 _1601_ (.B(_0736_),
    .A(_0020_),
    .X(_0750_));
 sg13g2_o21ai_1 _1602_ (.B1(_0737_),
    .Y(_0751_),
    .A1(_0749_),
    .A2(_0750_));
 sg13g2_a21oi_1 _1603_ (.A1(net260),
    .A2(_0729_),
    .Y(_0752_),
    .B1(\game1.obstacle2_x[8] ));
 sg13g2_nor2_1 _1604_ (.A(_0731_),
    .B(_0752_),
    .Y(_0753_));
 sg13g2_nand2b_1 _1605_ (.Y(_0754_),
    .B(net264),
    .A_N(_0734_));
 sg13g2_o21ai_1 _1606_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0019_),
    .A2(_0753_));
 sg13g2_a21o_1 _1607_ (.A2(_0751_),
    .A1(_0735_),
    .B1(_0755_),
    .X(_0756_));
 sg13g2_xnor2_1 _1608_ (.Y(_0757_),
    .A(_0018_),
    .B(_0732_));
 sg13g2_a21oi_1 _1609_ (.A1(_0019_),
    .A2(_0753_),
    .Y(_0758_),
    .B1(_0757_));
 sg13g2_a21oi_1 _1610_ (.A1(_0756_),
    .A2(_0758_),
    .Y(_0759_),
    .B1(_0733_));
 sg13g2_a21oi_1 _1611_ (.A1(\game1.obstacle2_x[9] ),
    .A2(_0731_),
    .Y(_0760_),
    .B1(_0759_));
 sg13g2_a22oi_1 _1612_ (.Y(_0761_),
    .B1(_0548_),
    .B2(\game1.obstacle2_x[8] ),
    .A2(net234),
    .A1(\game1.obstacle2_x[9] ));
 sg13g2_nand2_1 _1613_ (.Y(_0762_),
    .A(\game1.obstacle2_x[5] ),
    .B(_0545_));
 sg13g2_o21ai_1 _1614_ (.B1(_0762_),
    .Y(_0763_),
    .A1(_0519_),
    .A2(net267));
 sg13g2_nand2_1 _1615_ (.Y(_0764_),
    .A(net260),
    .B(_0543_));
 sg13g2_nor2_1 _1616_ (.A(\game1.obstacle2_x[5] ),
    .B(_0545_),
    .Y(_0765_));
 sg13g2_nor2_1 _1617_ (.A(\game1.obstacle2_x[4] ),
    .B(_0546_),
    .Y(_0766_));
 sg13g2_nor2_1 _1618_ (.A(_0765_),
    .B(_0766_),
    .Y(_0767_));
 sg13g2_nor2b_1 _1619_ (.A(net271),
    .B_N(\game1.obstacle2_x[4] ),
    .Y(_0768_));
 sg13g2_nor2b_1 _1620_ (.A(\game1.obstacle2_x[3] ),
    .B_N(net275),
    .Y(_0769_));
 sg13g2_o21ai_1 _1621_ (.B1(_0739_),
    .Y(_0770_),
    .A1(\game1.obstacle2_x[1] ),
    .A2(_0542_));
 sg13g2_nor2_1 _1622_ (.A(\game1.pixel_x[0] ),
    .B(_0770_),
    .Y(_0771_));
 sg13g2_o21ai_1 _1623_ (.B1(_0741_),
    .Y(_0772_),
    .A1(_0520_),
    .A2(net275));
 sg13g2_nor2_1 _1624_ (.A(_0771_),
    .B(_0772_),
    .Y(_0773_));
 sg13g2_a21oi_1 _1625_ (.A1(_0740_),
    .A2(_0773_),
    .Y(_0774_),
    .B1(_0769_));
 sg13g2_o21ai_1 _1626_ (.B1(_0767_),
    .Y(_0775_),
    .A1(_0768_),
    .A2(_0774_));
 sg13g2_nor4_1 _1627_ (.A(_0765_),
    .B(_0766_),
    .C(_0770_),
    .D(_0772_),
    .Y(_0776_));
 sg13g2_or2_1 _1628_ (.X(_0777_),
    .B(_0769_),
    .A(_0768_));
 sg13g2_o21ai_1 _1629_ (.B1(_0764_),
    .Y(_0778_),
    .A1(\game1.obstacle2_x[8] ),
    .A2(_0548_));
 sg13g2_nand2b_1 _1630_ (.Y(_0779_),
    .B(net264),
    .A_N(net260));
 sg13g2_o21ai_1 _1631_ (.B1(_0779_),
    .Y(_0780_),
    .A1(\game1.obstacle2_x[6] ),
    .A2(_0544_));
 sg13g2_o21ai_1 _1632_ (.B1(_0040_),
    .Y(_0781_),
    .A1(_0521_),
    .A2(\game1.pixel_x[1] ));
 sg13g2_nor4_1 _1633_ (.A(_0777_),
    .B(_0778_),
    .C(_0780_),
    .D(_0781_),
    .Y(_0782_));
 sg13g2_a22oi_1 _1634_ (.Y(_0783_),
    .B1(_0776_),
    .B2(_0782_),
    .A2(_0775_),
    .A1(_0764_));
 sg13g2_a22oi_1 _1635_ (.Y(_0784_),
    .B1(_0764_),
    .B2(_0780_),
    .A2(net263),
    .A1(_0518_));
 sg13g2_o21ai_1 _1636_ (.B1(_0784_),
    .Y(_0785_),
    .A1(_0763_),
    .A2(_0783_));
 sg13g2_a22oi_1 _1637_ (.Y(_0786_),
    .B1(_0761_),
    .B2(_0785_),
    .A2(net261),
    .A1(_0516_));
 sg13g2_nand2b_1 _1638_ (.Y(_0787_),
    .B(net247),
    .A_N(\game1.obstacle2_y[3] ));
 sg13g2_a22oi_1 _1639_ (.Y(_0788_),
    .B1(_0552_),
    .B2(\game1.obstacle2_y[2] ),
    .A2(_0550_),
    .A1(net256));
 sg13g2_o21ai_1 _1640_ (.B1(_0787_),
    .Y(_0789_),
    .A1(\game1.obstacle2_y[2] ),
    .A2(_0552_));
 sg13g2_nor2_1 _1641_ (.A(_0788_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_a221oi_1 _1642_ (.B2(\game1.obstacle2_y[4] ),
    .C1(_0790_),
    .B1(_0556_),
    .A1(\game1.obstacle2_y[3] ),
    .Y(_0791_),
    .A2(_0551_));
 sg13g2_a221oi_1 _1643_ (.B2(_0511_),
    .C1(_0791_),
    .B1(net245),
    .A1(_0510_),
    .Y(_0792_),
    .A2(net243));
 sg13g2_a221oi_1 _1644_ (.B2(\game1.obstacle2_y[5] ),
    .C1(_0792_),
    .B1(_0555_),
    .A1(\game1.obstacle2_y[6] ),
    .Y(_0793_),
    .A2(_0554_));
 sg13g2_a221oi_1 _1645_ (.B2(_0509_),
    .C1(_0793_),
    .B1(net241),
    .A1(_0508_),
    .Y(_0794_),
    .A2(net239));
 sg13g2_a221oi_1 _1646_ (.B2(\game1.obstacle2_y[8] ),
    .C1(_0794_),
    .B1(_0558_),
    .A1(\game1.obstacle2_y[7] ),
    .Y(_0795_),
    .A2(_0553_));
 sg13g2_a221oi_1 _1647_ (.B2(_0507_),
    .C1(_0795_),
    .B1(net238),
    .A1(_0505_),
    .Y(_0796_),
    .A2(net237));
 sg13g2_nand2_1 _1648_ (.Y(_0797_),
    .A(\game1.obstacle2_y[9] ),
    .B(_0557_));
 sg13g2_o21ai_1 _1649_ (.B1(_0797_),
    .Y(_0798_),
    .A1(_0557_),
    .A2(_0723_));
 sg13g2_or4_1 _1650_ (.A(_0760_),
    .B(_0786_),
    .C(_0796_),
    .D(_0798_),
    .X(_0799_));
 sg13g2_a21oi_2 _1651_ (.B1(_0799_),
    .Y(_0800_),
    .A2(_0726_),
    .A1(_0718_));
 sg13g2_o21ai_1 _1652_ (.B1(\game1.obstacle1_y[3] ),
    .Y(_0801_),
    .A1(\game1.obstacle1_y[2] ),
    .A2(net277));
 sg13g2_nor2_1 _1653_ (.A(_0527_),
    .B(_0801_),
    .Y(_0802_));
 sg13g2_nand2_1 _1654_ (.Y(_0803_),
    .A(\game1.obstacle1_y[5] ),
    .B(_0802_));
 sg13g2_nand2_1 _1655_ (.Y(_0804_),
    .A(_0525_),
    .B(_0803_));
 sg13g2_nand3_1 _1656_ (.B(\game1.obstacle1_y[7] ),
    .C(_0804_),
    .A(\game1.obstacle1_y[8] ),
    .Y(_0805_));
 sg13g2_xnor2_1 _1657_ (.Y(_0806_),
    .A(_0522_),
    .B(_0805_));
 sg13g2_and2_1 _1658_ (.A(net237),
    .B(_0806_),
    .X(_0807_));
 sg13g2_o21ai_1 _1659_ (.B1(_0027_),
    .Y(_0808_),
    .A1(\game1.obstacle1_y[6] ),
    .A2(_0803_));
 sg13g2_nand2_1 _1660_ (.Y(_0809_),
    .A(\game1.obstacle1_y[7] ),
    .B(_0808_));
 sg13g2_xnor2_1 _1661_ (.Y(_0810_),
    .A(\game1.obstacle1_y[7] ),
    .B(_0808_));
 sg13g2_nor3_1 _1662_ (.A(_0527_),
    .B(_0028_),
    .C(_0801_),
    .Y(_0811_));
 sg13g2_xnor2_1 _1663_ (.Y(_0812_),
    .A(\game1.obstacle1_y[6] ),
    .B(_0811_));
 sg13g2_nand2b_1 _1664_ (.Y(_0813_),
    .B(net241),
    .A_N(_0812_));
 sg13g2_xnor2_1 _1665_ (.Y(_0814_),
    .A(\game1.obstacle1_y[4] ),
    .B(_0801_));
 sg13g2_or3_1 _1666_ (.A(\game1.obstacle1_y[3] ),
    .B(\game1.obstacle1_y[2] ),
    .C(net277),
    .X(_0815_));
 sg13g2_nand2_1 _1667_ (.Y(_0816_),
    .A(_0801_),
    .B(_0815_));
 sg13g2_nor2_1 _1668_ (.A(net247),
    .B(_0816_),
    .Y(_0817_));
 sg13g2_xor2_1 _1669_ (.B(net277),
    .A(\game1.obstacle1_y[2] ),
    .X(_0818_));
 sg13g2_xnor2_1 _1670_ (.Y(_0819_),
    .A(_0032_),
    .B(_0818_));
 sg13g2_o21ai_1 _1671_ (.B1(_0819_),
    .Y(_0820_),
    .A1(net277),
    .A2(net250));
 sg13g2_a22oi_1 _1672_ (.Y(_0821_),
    .B1(_0818_),
    .B2(net249),
    .A2(_0816_),
    .A1(net246));
 sg13g2_a21o_1 _1673_ (.A2(_0821_),
    .A1(_0820_),
    .B1(_0817_),
    .X(_0822_));
 sg13g2_o21ai_1 _1674_ (.B1(_0822_),
    .Y(_0823_),
    .A1(_0031_),
    .A2(_0814_));
 sg13g2_xor2_1 _1675_ (.B(_0802_),
    .A(_0028_),
    .X(_0824_));
 sg13g2_xor2_1 _1676_ (.B(_0824_),
    .A(_0030_),
    .X(_0825_));
 sg13g2_a21oi_1 _1677_ (.A1(_0031_),
    .A2(_0814_),
    .Y(_0826_),
    .B1(_0825_));
 sg13g2_a22oi_1 _1678_ (.Y(_0827_),
    .B1(_0826_),
    .B2(_0823_),
    .A2(_0824_),
    .A1(net244));
 sg13g2_xnor2_1 _1679_ (.Y(_0828_),
    .A(_0029_),
    .B(_0812_));
 sg13g2_o21ai_1 _1680_ (.B1(_0813_),
    .Y(_0829_),
    .A1(_0827_),
    .A2(_0828_));
 sg13g2_o21ai_1 _1681_ (.B1(_0829_),
    .Y(_0830_),
    .A1(net240),
    .A2(_0810_));
 sg13g2_xor2_1 _1682_ (.B(_0809_),
    .A(_0026_),
    .X(_0831_));
 sg13g2_nor2_1 _1683_ (.A(_0025_),
    .B(_0831_),
    .Y(_0832_));
 sg13g2_a21oi_1 _1684_ (.A1(net240),
    .A2(_0810_),
    .Y(_0833_),
    .B1(_0832_));
 sg13g2_xor2_1 _1685_ (.B(_0806_),
    .A(_0024_),
    .X(_0834_));
 sg13g2_a221oi_1 _1686_ (.B2(_0830_),
    .C1(_0834_),
    .B1(_0833_),
    .A1(_0025_),
    .Y(_0835_),
    .A2(_0831_));
 sg13g2_or2_1 _1687_ (.X(_0836_),
    .B(_0805_),
    .A(_0023_));
 sg13g2_o21ai_1 _1688_ (.B1(_0836_),
    .Y(_0837_),
    .A1(_0807_),
    .A2(_0835_));
 sg13g2_nand2_1 _1689_ (.Y(_0838_),
    .A(net259),
    .B(_0543_));
 sg13g2_nor2b_1 _1690_ (.A(net276),
    .B_N(\game1.obstacle1_x[2] ),
    .Y(_0839_));
 sg13g2_nand2b_1 _1691_ (.Y(_0840_),
    .B(net276),
    .A_N(\game1.obstacle1_x[2] ));
 sg13g2_nor2b_1 _1692_ (.A(\game1.pixel_x[1] ),
    .B_N(\game1.obstacle1_x[1] ),
    .Y(_0841_));
 sg13g2_o21ai_1 _1693_ (.B1(_0840_),
    .Y(_0842_),
    .A1(_0839_),
    .A2(_0841_));
 sg13g2_nor2_1 _1694_ (.A(net274),
    .B(_0842_),
    .Y(_0843_));
 sg13g2_a22oi_1 _1695_ (.Y(_0844_),
    .B1(_0842_),
    .B2(net274),
    .A2(net271),
    .A1(_0515_));
 sg13g2_o21ai_1 _1696_ (.B1(_0844_),
    .Y(_0845_),
    .A1(\game1.obstacle1_x[3] ),
    .A2(_0843_));
 sg13g2_nor2_1 _1697_ (.A(\game1.obstacle1_x[5] ),
    .B(_0545_),
    .Y(_0846_));
 sg13g2_nor2_1 _1698_ (.A(_0514_),
    .B(net266),
    .Y(_0847_));
 sg13g2_a22oi_1 _1699_ (.Y(_0848_),
    .B1(_0546_),
    .B2(\game1.obstacle1_x[4] ),
    .A2(_0545_),
    .A1(\game1.obstacle1_x[5] ));
 sg13g2_nand2b_1 _1700_ (.Y(_0849_),
    .B(net265),
    .A_N(net259));
 sg13g2_a221oi_1 _1701_ (.B2(_0848_),
    .C1(_0846_),
    .B1(_0845_),
    .A1(_0514_),
    .Y(_0850_),
    .A2(net266));
 sg13g2_o21ai_1 _1702_ (.B1(_0849_),
    .Y(_0851_),
    .A1(_0847_),
    .A2(_0850_));
 sg13g2_a22oi_1 _1703_ (.Y(_0852_),
    .B1(_0838_),
    .B2(_0851_),
    .A2(net263),
    .A1(_0513_));
 sg13g2_a221oi_1 _1704_ (.B2(\game1.obstacle1_x[8] ),
    .C1(_0852_),
    .B1(_0548_),
    .A1(\game1.obstacle1_x[9] ),
    .Y(_0853_),
    .A2(_0547_));
 sg13g2_a21oi_1 _1705_ (.A1(_0512_),
    .A2(net262),
    .Y(_0854_),
    .B1(_0853_));
 sg13g2_nor3_2 _1706_ (.A(\game1.obstacle1_x[5] ),
    .B(\game1.obstacle1_x[4] ),
    .C(\game1.obstacle1_x[3] ),
    .Y(_0855_));
 sg13g2_and2_1 _1707_ (.A(_0514_),
    .B(_0855_),
    .X(_0856_));
 sg13g2_nor2b_1 _1708_ (.A(_0856_),
    .B_N(net259),
    .Y(_0857_));
 sg13g2_and2_1 _1709_ (.A(\game1.obstacle1_x[8] ),
    .B(_0857_),
    .X(_0858_));
 sg13g2_xor2_1 _1710_ (.B(_0858_),
    .A(_0017_),
    .X(_0859_));
 sg13g2_xnor2_1 _1711_ (.Y(_0860_),
    .A(_0513_),
    .B(_0857_));
 sg13g2_nor2_1 _1712_ (.A(_0019_),
    .B(_0860_),
    .Y(_0861_));
 sg13g2_xnor2_1 _1713_ (.Y(_0862_),
    .A(net259),
    .B(_0856_));
 sg13g2_inv_1 _1714_ (.Y(_0863_),
    .A(_0862_));
 sg13g2_nand2_1 _1715_ (.Y(_0864_),
    .A(_0543_),
    .B(_0862_));
 sg13g2_o21ai_1 _1716_ (.B1(\game1.obstacle1_x[5] ),
    .Y(_0865_),
    .A1(\game1.obstacle1_x[4] ),
    .A2(\game1.obstacle1_x[3] ));
 sg13g2_nor2b_1 _1717_ (.A(_0855_),
    .B_N(_0865_),
    .Y(_0866_));
 sg13g2_o21ai_1 _1718_ (.B1(\game1.obstacle1_x[3] ),
    .Y(_0867_),
    .A1(net274),
    .A2(_0842_));
 sg13g2_xnor2_1 _1719_ (.Y(_0868_),
    .A(\game1.obstacle1_x[4] ),
    .B(\game1.obstacle1_x[3] ));
 sg13g2_nor2_1 _1720_ (.A(net270),
    .B(_0868_),
    .Y(_0869_));
 sg13g2_a21oi_1 _1721_ (.A1(net274),
    .A2(_0842_),
    .Y(_0870_),
    .B1(_0869_));
 sg13g2_a22oi_1 _1722_ (.Y(_0871_),
    .B1(_0870_),
    .B2(_0867_),
    .A2(_0868_),
    .A1(net270));
 sg13g2_xnor2_1 _1723_ (.Y(_0872_),
    .A(_0021_),
    .B(_0866_));
 sg13g2_a22oi_1 _1724_ (.Y(_0873_),
    .B1(_0871_),
    .B2(_0872_),
    .A2(_0866_),
    .A1(net268));
 sg13g2_xnor2_1 _1725_ (.Y(_0874_),
    .A(\game1.obstacle1_x[6] ),
    .B(_0855_));
 sg13g2_xor2_1 _1726_ (.B(_0874_),
    .A(_0020_),
    .X(_0875_));
 sg13g2_a22oi_1 _1727_ (.Y(_0876_),
    .B1(_0874_),
    .B2(net266),
    .A2(_0863_),
    .A1(net264));
 sg13g2_o21ai_1 _1728_ (.B1(_0876_),
    .Y(_0877_),
    .A1(_0873_),
    .A2(_0875_));
 sg13g2_a21o_1 _1729_ (.A2(_0877_),
    .A1(_0864_),
    .B1(_0861_),
    .X(_0878_));
 sg13g2_xor2_1 _1730_ (.B(_0859_),
    .A(_0018_),
    .X(_0879_));
 sg13g2_a21oi_1 _1731_ (.A1(_0019_),
    .A2(_0860_),
    .Y(_0880_),
    .B1(_0879_));
 sg13g2_a22oi_1 _1732_ (.Y(_0881_),
    .B1(_0878_),
    .B2(_0880_),
    .A2(_0859_),
    .A1(net262));
 sg13g2_a21oi_1 _1733_ (.A1(\game1.obstacle1_x[9] ),
    .A2(_0858_),
    .Y(_0882_),
    .B1(_0881_));
 sg13g2_nand2b_1 _1734_ (.Y(_0883_),
    .B(\game1.obstacle1_y[2] ),
    .A_N(net249));
 sg13g2_nand2b_1 _1735_ (.Y(_0884_),
    .B(net248),
    .A_N(\game1.obstacle1_y[2] ));
 sg13g2_nand3b_1 _1736_ (.B(_0884_),
    .C(net277),
    .Y(_0885_),
    .A_N(net250));
 sg13g2_a22oi_1 _1737_ (.Y(_0886_),
    .B1(_0883_),
    .B2(_0885_),
    .A2(net246),
    .A1(_0528_));
 sg13g2_a221oi_1 _1738_ (.B2(\game1.obstacle1_y[4] ),
    .C1(_0886_),
    .B1(_0556_),
    .A1(\game1.obstacle1_y[3] ),
    .Y(_0887_),
    .A2(_0551_));
 sg13g2_a221oi_1 _1739_ (.B2(_0527_),
    .C1(_0887_),
    .B1(net245),
    .A1(_0526_),
    .Y(_0888_),
    .A2(net244));
 sg13g2_a221oi_1 _1740_ (.B2(\game1.obstacle1_y[5] ),
    .C1(_0888_),
    .B1(_0555_),
    .A1(\game1.obstacle1_y[6] ),
    .Y(_0889_),
    .A2(_0554_));
 sg13g2_a221oi_1 _1741_ (.B2(_0525_),
    .C1(_0889_),
    .B1(net241),
    .A1(_0524_),
    .Y(_0890_),
    .A2(net240));
 sg13g2_a221oi_1 _1742_ (.B2(\game1.obstacle1_y[8] ),
    .C1(_0890_),
    .B1(_0558_),
    .A1(\game1.obstacle1_y[7] ),
    .Y(_0891_),
    .A2(_0553_));
 sg13g2_a221oi_1 _1743_ (.B2(_0523_),
    .C1(_0891_),
    .B1(net238),
    .A1(_0522_),
    .Y(_0892_),
    .A2(\game1.pixel_y[9] ));
 sg13g2_nor2_1 _1744_ (.A(_0522_),
    .B(\game1.pixel_y[9] ),
    .Y(_0893_));
 sg13g2_nor4_1 _1745_ (.A(_0854_),
    .B(_0882_),
    .C(_0892_),
    .D(_0893_),
    .Y(_0894_));
 sg13g2_and2_1 _1746_ (.A(_0837_),
    .B(_0894_),
    .X(_0895_));
 sg13g2_nor3_2 _1747_ (.A(_0689_),
    .B(_0800_),
    .C(_0895_),
    .Y(_0896_));
 sg13g2_a21oi_2 _1748_ (.B1(_0597_),
    .Y(uo_out[6]),
    .A2(_0896_),
    .A1(_0564_));
 sg13g2_and2_2 _1749_ (.A(\game1.pixel_x[1] ),
    .B(net363),
    .X(_0897_));
 sg13g2_nor2_1 _1750_ (.A(net417),
    .B(net350),
    .Y(_0898_));
 sg13g2_nand2_1 _1751_ (.Y(_0899_),
    .A(\game1.pixel_x[2] ),
    .B(net272));
 sg13g2_nor2_1 _1752_ (.A(net241),
    .B(net243),
    .Y(_0900_));
 sg13g2_nand2_1 _1753_ (.Y(_0901_),
    .A(net263),
    .B(net240));
 sg13g2_nand2_1 _1754_ (.Y(_0902_),
    .A(_0555_),
    .B(_0585_));
 sg13g2_o21ai_1 _1755_ (.B1(_0902_),
    .Y(_0903_),
    .A1(net242),
    .A2(_0589_));
 sg13g2_nand2_1 _1756_ (.Y(_0904_),
    .A(net274),
    .B(net272));
 sg13g2_nor2b_1 _1757_ (.A(net269),
    .B_N(net272),
    .Y(_0905_));
 sg13g2_nand3_1 _1758_ (.B(_0898_),
    .C(_0905_),
    .A(net276),
    .Y(_0906_));
 sg13g2_o21ai_1 _1759_ (.B1(_0906_),
    .Y(_0907_),
    .A1(net266),
    .A2(_0897_));
 sg13g2_nand3b_1 _1760_ (.B(_0543_),
    .C(_0907_),
    .Y(_0908_),
    .A_N(net273));
 sg13g2_nor4_1 _1761_ (.A(net262),
    .B(_0587_),
    .C(_0900_),
    .D(_0901_),
    .Y(_0909_));
 sg13g2_nand2_1 _1762_ (.Y(_0910_),
    .A(_0543_),
    .B(_0544_));
 sg13g2_nor2_1 _1763_ (.A(net265),
    .B(net269),
    .Y(_0911_));
 sg13g2_nand4_1 _1764_ (.B(_0904_),
    .C(_0910_),
    .A(_0899_),
    .Y(_0912_),
    .D(_0911_));
 sg13g2_o21ai_1 _1765_ (.B1(_0912_),
    .Y(_0913_),
    .A1(_0568_),
    .A2(_0910_));
 sg13g2_nand4_1 _1766_ (.B(_0908_),
    .C(_0909_),
    .A(_0903_),
    .Y(_0914_),
    .D(_0913_));
 sg13g2_inv_1 _1767_ (.Y(_0915_),
    .A(_0914_));
 sg13g2_nand2_1 _1768_ (.Y(_0916_),
    .A(_0896_),
    .B(_0915_));
 sg13g2_a21oi_2 _1769_ (.B1(_0597_),
    .Y(uo_out[5]),
    .A2(_0916_),
    .A1(_0010_));
 sg13g2_nand2_1 _1770_ (.Y(_0917_),
    .A(_0896_),
    .B(_0914_));
 sg13g2_a21oi_2 _1771_ (.B1(_0597_),
    .Y(uo_out[4]),
    .A2(_0917_),
    .A1(_0010_));
 sg13g2_o21ai_1 _1772_ (.B1(net1),
    .Y(_0918_),
    .A1(_0896_),
    .A2(_0914_));
 sg13g2_inv_2 _1773_ (.Y(_0919_),
    .A(net226));
 sg13g2_nand3_1 _1774_ (.B(\game1.obstacle3_y[2] ),
    .C(net279),
    .A(net346),
    .Y(_0920_));
 sg13g2_or2_1 _1775_ (.X(_0921_),
    .B(_0920_),
    .A(_0540_));
 sg13g2_nand2_1 _1776_ (.Y(_0922_),
    .A(\game1.obstacle3_y[6] ),
    .B(\game1.obstacle3_y[5] ));
 sg13g2_nor2_1 _1777_ (.A(_0921_),
    .B(_0922_),
    .Y(_0923_));
 sg13g2_nor3_1 _1778_ (.A(_0011_),
    .B(_0921_),
    .C(_0922_),
    .Y(_0924_));
 sg13g2_xnor2_1 _1779_ (.Y(_0925_),
    .A(_0011_),
    .B(_0923_));
 sg13g2_nor2_1 _1780_ (.A(_0013_),
    .B(_0921_),
    .Y(_0926_));
 sg13g2_xor2_1 _1781_ (.B(_0921_),
    .A(_0013_),
    .X(_0927_));
 sg13g2_nor2_1 _1782_ (.A(_0012_),
    .B(_0015_),
    .Y(_0928_));
 sg13g2_xnor2_1 _1783_ (.Y(_0929_),
    .A(_0015_),
    .B(_0924_));
 sg13g2_nand3_1 _1784_ (.B(_0927_),
    .C(_0928_),
    .A(_0925_),
    .Y(_0930_));
 sg13g2_nand2b_1 _1785_ (.Y(_0931_),
    .B(_0923_),
    .A_N(_0601_));
 sg13g2_nor2_1 _1786_ (.A(\game1.obstacle3_y[9] ),
    .B(_0014_),
    .Y(_0932_));
 sg13g2_mux2_1 _1787_ (.A0(_0932_),
    .A1(_0014_),
    .S(_0931_),
    .X(_0933_));
 sg13g2_and3_2 _1788_ (.X(_0934_),
    .A(net165),
    .B(_0930_),
    .C(_0933_));
 sg13g2_nand2b_1 _1789_ (.Y(_0935_),
    .B(_0934_),
    .A_N(net279));
 sg13g2_nand2_1 _1790_ (.Y(_0936_),
    .A(net236),
    .B(net279));
 sg13g2_a21oi_1 _1791_ (.A1(_0935_),
    .A2(_0936_),
    .Y(_0041_),
    .B1(net225));
 sg13g2_a22oi_1 _1792_ (.Y(_0937_),
    .B1(_0616_),
    .B2(_0934_),
    .A2(net399),
    .A1(net236));
 sg13g2_nor2_1 _1793_ (.A(net225),
    .B(_0937_),
    .Y(_0042_));
 sg13g2_a21o_1 _1794_ (.A2(net279),
    .A1(\game1.obstacle3_y[2] ),
    .B1(\game1.obstacle3_y[3] ),
    .X(_0938_));
 sg13g2_and2_1 _1795_ (.A(_0920_),
    .B(_0938_),
    .X(_0939_));
 sg13g2_a22oi_1 _1796_ (.Y(_0940_),
    .B1(_0934_),
    .B2(_0939_),
    .A2(net346),
    .A1(net236));
 sg13g2_nor2_1 _1797_ (.A(net225),
    .B(net347),
    .Y(_0043_));
 sg13g2_xnor2_1 _1798_ (.Y(_0941_),
    .A(net354),
    .B(_0920_));
 sg13g2_a22oi_1 _1799_ (.Y(_0942_),
    .B1(_0934_),
    .B2(_0941_),
    .A2(net354),
    .A1(net236));
 sg13g2_nor2_1 _1800_ (.A(net225),
    .B(_0942_),
    .Y(_0044_));
 sg13g2_a22oi_1 _1801_ (.Y(_0943_),
    .B1(_0927_),
    .B2(_0934_),
    .A2(net315),
    .A1(net236));
 sg13g2_nor2_1 _1802_ (.A(net225),
    .B(net316),
    .Y(_0045_));
 sg13g2_xnor2_1 _1803_ (.Y(_0944_),
    .A(net368),
    .B(_0926_));
 sg13g2_a22oi_1 _1804_ (.Y(_0945_),
    .B1(_0934_),
    .B2(_0944_),
    .A2(\game1.obstacle3_y[6] ),
    .A1(net236));
 sg13g2_nand2_1 _1805_ (.Y(_0046_),
    .A(net220),
    .B(net369));
 sg13g2_a22oi_1 _1806_ (.Y(_0946_),
    .B1(_0925_),
    .B2(_0934_),
    .A2(net324),
    .A1(net236));
 sg13g2_nor2_1 _1807_ (.A(net225),
    .B(net325),
    .Y(_0047_));
 sg13g2_a22oi_1 _1808_ (.Y(_0947_),
    .B1(_0929_),
    .B2(_0934_),
    .A2(net329),
    .A1(net236));
 sg13g2_nand2_1 _1809_ (.Y(_0048_),
    .A(net220),
    .B(net330));
 sg13g2_nor3_1 _1810_ (.A(net165),
    .B(_0535_),
    .C(net225),
    .Y(_0049_));
 sg13g2_xnor2_1 _1811_ (.Y(_0948_),
    .A(net257),
    .B(net331));
 sg13g2_nor2_1 _1812_ (.A(net222),
    .B(net332),
    .Y(_0050_));
 sg13g2_o21ai_1 _1813_ (.B1(net300),
    .Y(_0949_),
    .A1(_0517_),
    .A2(\game1.obstacle3_x[1] ));
 sg13g2_nor2_1 _1814_ (.A(net300),
    .B(net331),
    .Y(_0950_));
 sg13g2_nand2_1 _1815_ (.Y(_0951_),
    .A(net257),
    .B(_0950_));
 sg13g2_a21oi_1 _1816_ (.A1(net301),
    .A2(_0951_),
    .Y(_0051_),
    .B1(net222));
 sg13g2_nor2_1 _1817_ (.A(net278),
    .B(_0951_),
    .Y(_0952_));
 sg13g2_xor2_1 _1818_ (.B(_0951_),
    .A(net278),
    .X(_0953_));
 sg13g2_nor2_1 _1819_ (.A(net223),
    .B(_0953_),
    .Y(_0052_));
 sg13g2_xnor2_1 _1820_ (.Y(_0954_),
    .A(net398),
    .B(_0952_));
 sg13g2_nand2_1 _1821_ (.Y(_0053_),
    .A(net220),
    .B(_0954_));
 sg13g2_nand3_1 _1822_ (.B(_0638_),
    .C(_0950_),
    .A(net257),
    .Y(_0955_));
 sg13g2_a21o_1 _1823_ (.A2(_0952_),
    .A1(_0534_),
    .B1(_0533_),
    .X(_0956_));
 sg13g2_a21oi_1 _1824_ (.A1(_0955_),
    .A2(_0956_),
    .Y(_0054_),
    .B1(net223));
 sg13g2_xnor2_1 _1825_ (.Y(_0957_),
    .A(_0532_),
    .B(_0955_));
 sg13g2_nor2_1 _1826_ (.A(net222),
    .B(net427),
    .Y(_0055_));
 sg13g2_nor2_1 _1827_ (.A(net300),
    .B(_0639_),
    .Y(_0958_));
 sg13g2_nor2_1 _1828_ (.A(\game1.obstacle3_x[8] ),
    .B(net278),
    .Y(_0959_));
 sg13g2_nand3_1 _1829_ (.B(_0638_),
    .C(_0950_),
    .A(_0532_),
    .Y(_0960_));
 sg13g2_nand2b_1 _1830_ (.Y(_0961_),
    .B(_0531_),
    .A_N(_0960_));
 sg13g2_nor2_1 _1831_ (.A(\game1.obstacle3_x[8] ),
    .B(_0961_),
    .Y(_0962_));
 sg13g2_xnor2_1 _1832_ (.Y(_0963_),
    .A(net385),
    .B(_0962_));
 sg13g2_nand4_1 _1833_ (.B(net385),
    .C(_0958_),
    .A(net331),
    .Y(_0964_),
    .D(_0959_));
 sg13g2_a21oi_1 _1834_ (.A1(\game1.obstacle3_x[7] ),
    .A2(_0960_),
    .Y(_0965_),
    .B1(_0517_));
 sg13g2_nand3_1 _1835_ (.B(_0964_),
    .C(_0965_),
    .A(_0961_),
    .Y(_0966_));
 sg13g2_o21ai_1 _1836_ (.B1(_0966_),
    .Y(_0967_),
    .A1(net257),
    .A2(net412));
 sg13g2_nand2_1 _1837_ (.Y(_0056_),
    .A(net220),
    .B(net413));
 sg13g2_nor2_1 _1838_ (.A(_0517_),
    .B(_0961_),
    .Y(_0968_));
 sg13g2_xnor2_1 _1839_ (.Y(_0969_),
    .A(net404),
    .B(_0968_));
 sg13g2_nand2_1 _1840_ (.Y(_0057_),
    .A(net220),
    .B(_0969_));
 sg13g2_nand4_1 _1841_ (.B(_0958_),
    .C(_0959_),
    .A(net331),
    .Y(_0970_),
    .D(_0965_));
 sg13g2_o21ai_1 _1842_ (.B1(_0970_),
    .Y(_0971_),
    .A1(net257),
    .A2(_0529_));
 sg13g2_a21oi_1 _1843_ (.A1(net257),
    .A2(_0963_),
    .Y(_0972_),
    .B1(_0971_));
 sg13g2_nor2_1 _1844_ (.A(net222),
    .B(net386),
    .Y(_0058_));
 sg13g2_nor2b_1 _1845_ (.A(\game1.scroll1_v_inst.ctr[8] ),
    .B_N(\game1.scroll1_v_inst.ctr[9] ),
    .Y(_0973_));
 sg13g2_nor2b_1 _1846_ (.A(\game1.scroll1_v_inst.ctr[6] ),
    .B_N(\game1.scroll1_v_inst.ctr[7] ),
    .Y(_0974_));
 sg13g2_a21o_1 _1847_ (.A2(_0974_),
    .A1(_0005_),
    .B1(_0004_),
    .X(_0975_));
 sg13g2_a21oi_1 _1848_ (.A1(_0973_),
    .A2(_0975_),
    .Y(_0976_),
    .B1(_0003_));
 sg13g2_nor4_1 _1849_ (.A(_0502_),
    .B(\game1.scroll1_v_inst.ctr[4] ),
    .C(\game1.scroll1_v_inst.ctr[3] ),
    .D(\game1.scroll1_v_inst.ctr[2] ),
    .Y(_0977_));
 sg13g2_nor2_1 _1850_ (.A(net191),
    .B(\game1.scroll1_v_inst.ctr[0] ),
    .Y(_0978_));
 sg13g2_and4_1 _1851_ (.A(_0973_),
    .B(_0974_),
    .C(_0977_),
    .D(_0978_),
    .X(_0979_));
 sg13g2_o21ai_1 _1852_ (.B1(\game1.scroll1_v_inst.ctr[10] ),
    .Y(_0980_),
    .A1(_0976_),
    .A2(_0979_));
 sg13g2_nor4_1 _1853_ (.A(\game1.scroll1_v_inst.ctr[14] ),
    .B(\game1.scroll1_v_inst.ctr[13] ),
    .C(\game1.scroll1_v_inst.ctr[12] ),
    .D(\game1.scroll1_v_inst.ctr[11] ),
    .Y(_0981_));
 sg13g2_nand2_1 _1854_ (.Y(_0982_),
    .A(\game1.scroll1_v_inst.ctr[16] ),
    .B(\game1.scroll1_v_inst.ctr[15] ));
 sg13g2_a21oi_1 _1855_ (.A1(_0980_),
    .A2(_0981_),
    .Y(_0983_),
    .B1(_0982_));
 sg13g2_nor2_1 _1856_ (.A(net177),
    .B(_0983_),
    .Y(_0984_));
 sg13g2_nor2_2 _1857_ (.A(_0501_),
    .B(_0984_),
    .Y(_0985_));
 sg13g2_or2_1 _1858_ (.X(_0986_),
    .B(_0985_),
    .A(net228));
 sg13g2_nor2_1 _1859_ (.A(net163),
    .B(net216),
    .Y(_0987_));
 sg13g2_nor2b_1 _1860_ (.A(net228),
    .B_N(_0985_),
    .Y(_0157_));
 sg13g2_nand3_1 _1861_ (.B(\game1.obstacle1_y[2] ),
    .C(net277),
    .A(\game1.obstacle1_y[3] ),
    .Y(_0988_));
 sg13g2_or2_1 _1862_ (.X(_0989_),
    .B(_0988_),
    .A(_0527_));
 sg13g2_or3_1 _1863_ (.A(_0525_),
    .B(_0526_),
    .C(_0989_),
    .X(_0990_));
 sg13g2_or2_1 _1864_ (.X(_0991_),
    .B(_0990_),
    .A(_0524_));
 sg13g2_xnor2_1 _1865_ (.Y(_0992_),
    .A(_0524_),
    .B(_0990_));
 sg13g2_nor2_1 _1866_ (.A(_0028_),
    .B(_0989_),
    .Y(_0993_));
 sg13g2_xnor2_1 _1867_ (.Y(_0994_),
    .A(_0028_),
    .B(_0989_));
 sg13g2_inv_1 _1868_ (.Y(_0995_),
    .A(_0994_));
 sg13g2_nor4_2 _1869_ (.A(_0027_),
    .B(_0026_),
    .C(_0992_),
    .Y(_0996_),
    .D(_0994_));
 sg13g2_or2_1 _1870_ (.X(_0997_),
    .B(_0991_),
    .A(_0523_));
 sg13g2_nand2_1 _1871_ (.Y(_0998_),
    .A(_0023_),
    .B(_0997_));
 sg13g2_xor2_1 _1872_ (.B(_0997_),
    .A(_0023_),
    .X(_0999_));
 sg13g2_or3_1 _1873_ (.A(net277),
    .B(_0996_),
    .C(_0999_),
    .X(_1000_));
 sg13g2_a21oi_1 _1874_ (.A1(net215),
    .A2(_1000_),
    .Y(_0059_),
    .B1(_0987_));
 sg13g2_nor2_1 _1875_ (.A(net364),
    .B(net216),
    .Y(_1001_));
 sg13g2_nor2_2 _1876_ (.A(_0996_),
    .B(_0998_),
    .Y(_1002_));
 sg13g2_nand2_1 _1877_ (.Y(_1003_),
    .A(_0818_),
    .B(_1002_));
 sg13g2_a21oi_1 _1878_ (.A1(net215),
    .A2(_1003_),
    .Y(_0060_),
    .B1(_1001_));
 sg13g2_a21o_1 _1879_ (.A2(net277),
    .A1(\game1.obstacle1_y[2] ),
    .B1(net348),
    .X(_1004_));
 sg13g2_nand4_1 _1880_ (.B(_0988_),
    .C(_1002_),
    .A(net215),
    .Y(_1005_),
    .D(_1004_));
 sg13g2_o21ai_1 _1881_ (.B1(_1005_),
    .Y(_0061_),
    .A1(_0528_),
    .A2(net216));
 sg13g2_nor2_1 _1882_ (.A(net287),
    .B(net216),
    .Y(_1006_));
 sg13g2_nand2_1 _1883_ (.Y(_1007_),
    .A(_0527_),
    .B(_0988_));
 sg13g2_nand3_1 _1884_ (.B(_1002_),
    .C(_1007_),
    .A(_0989_),
    .Y(_1008_));
 sg13g2_a21oi_1 _1885_ (.A1(_0157_),
    .A2(_1008_),
    .Y(_0062_),
    .B1(_1006_));
 sg13g2_nand3_1 _1886_ (.B(_0995_),
    .C(_1002_),
    .A(_0157_),
    .Y(_1009_));
 sg13g2_o21ai_1 _1887_ (.B1(_1009_),
    .Y(_0063_),
    .A1(_0526_),
    .A2(net216));
 sg13g2_xnor2_1 _1888_ (.Y(_1010_),
    .A(net370),
    .B(_0993_));
 sg13g2_nand3_1 _1889_ (.B(_1002_),
    .C(net371),
    .A(net215),
    .Y(_1011_));
 sg13g2_o21ai_1 _1890_ (.B1(net372),
    .Y(_0064_),
    .A1(_0525_),
    .A2(net216));
 sg13g2_nor2_1 _1891_ (.A(net333),
    .B(net219),
    .Y(_1012_));
 sg13g2_nand2b_1 _1892_ (.Y(_1013_),
    .B(_1002_),
    .A_N(_0992_));
 sg13g2_a21oi_1 _1893_ (.A1(net215),
    .A2(_1013_),
    .Y(_0065_),
    .B1(_1012_));
 sg13g2_xor2_1 _1894_ (.B(_0991_),
    .A(_0026_),
    .X(_1014_));
 sg13g2_nand3_1 _1895_ (.B(_1002_),
    .C(_1014_),
    .A(net215),
    .Y(_1015_));
 sg13g2_o21ai_1 _1896_ (.B1(_1015_),
    .Y(_0066_),
    .A1(_0523_),
    .A2(net219));
 sg13g2_nor2_1 _1897_ (.A(_0522_),
    .B(net216),
    .Y(_0067_));
 sg13g2_and2_2 _1898_ (.A(net273),
    .B(_0897_),
    .X(_1016_));
 sg13g2_and2_1 _1899_ (.A(net417),
    .B(net350),
    .X(_1017_));
 sg13g2_and2_1 _1900_ (.A(net350),
    .B(_1016_),
    .X(_1018_));
 sg13g2_nand2_2 _1901_ (.Y(_1019_),
    .A(net350),
    .B(_1016_));
 sg13g2_nor2_1 _1902_ (.A(_0565_),
    .B(_0910_),
    .Y(_1020_));
 sg13g2_nand3_1 _1903_ (.B(_1018_),
    .C(_1020_),
    .A(_0905_),
    .Y(_1021_));
 sg13g2_and2_1 _1904_ (.A(net1),
    .B(_1021_),
    .X(_1022_));
 sg13g2_nand2_1 _1905_ (.Y(_1023_),
    .A(net1),
    .B(_1021_));
 sg13g2_and2_1 _1906_ (.A(net152),
    .B(net232),
    .X(_0068_));
 sg13g2_nor3_1 _1907_ (.A(_0898_),
    .B(_1017_),
    .C(_1023_),
    .Y(_0069_));
 sg13g2_o21ai_1 _1908_ (.B1(net1),
    .Y(_1024_),
    .A1(net276),
    .A2(_1017_));
 sg13g2_a21oi_1 _1909_ (.A1(net350),
    .A2(_0897_),
    .Y(_0070_),
    .B1(_1024_));
 sg13g2_a21oi_1 _1910_ (.A1(net350),
    .A2(_0897_),
    .Y(_1025_),
    .B1(net273));
 sg13g2_nor3_1 _1911_ (.A(_0541_),
    .B(_1018_),
    .C(_1025_),
    .Y(_0071_));
 sg13g2_o21ai_1 _1912_ (.B1(net1),
    .Y(_1026_),
    .A1(_0546_),
    .A2(_1019_));
 sg13g2_a21oi_1 _1913_ (.A1(_0546_),
    .A2(_1019_),
    .Y(_0072_),
    .B1(_1026_));
 sg13g2_nor2_1 _1914_ (.A(net270),
    .B(_1019_),
    .Y(_1027_));
 sg13g2_o21ai_1 _1915_ (.B1(net232),
    .Y(_1028_),
    .A1(net268),
    .A2(_1027_));
 sg13g2_a21oi_1 _1916_ (.A1(net268),
    .A2(_1027_),
    .Y(_0073_),
    .B1(_1028_));
 sg13g2_nor2_1 _1917_ (.A(_0568_),
    .B(_1019_),
    .Y(_1029_));
 sg13g2_o21ai_1 _1918_ (.B1(net232),
    .Y(_1030_),
    .A1(net266),
    .A2(_1029_));
 sg13g2_a21oi_1 _1919_ (.A1(net266),
    .A2(_1029_),
    .Y(_0074_),
    .B1(_1030_));
 sg13g2_nor3_1 _1920_ (.A(_0020_),
    .B(_0568_),
    .C(_1019_),
    .Y(_1031_));
 sg13g2_o21ai_1 _1921_ (.B1(net232),
    .Y(_1032_),
    .A1(net265),
    .A2(_1031_));
 sg13g2_a21oi_1 _1922_ (.A1(net265),
    .A2(_1031_),
    .Y(_0075_),
    .B1(_1032_));
 sg13g2_nor2_1 _1923_ (.A(_0570_),
    .B(_1019_),
    .Y(_1033_));
 sg13g2_o21ai_1 _1924_ (.B1(net232),
    .Y(_1034_),
    .A1(net263),
    .A2(_1033_));
 sg13g2_a21oi_1 _1925_ (.A1(net263),
    .A2(_1033_),
    .Y(_0076_),
    .B1(_1034_));
 sg13g2_nor3_1 _1926_ (.A(_0019_),
    .B(_0570_),
    .C(_1019_),
    .Y(_1035_));
 sg13g2_o21ai_1 _1927_ (.B1(net232),
    .Y(_1036_),
    .A1(net261),
    .A2(_1035_));
 sg13g2_a21oi_1 _1928_ (.A1(net261),
    .A2(_1035_),
    .Y(_0077_),
    .B1(_1036_));
 sg13g2_xnor2_1 _1929_ (.Y(_1037_),
    .A(net257),
    .B(net359));
 sg13g2_nor2_1 _1930_ (.A(net222),
    .B(net360),
    .Y(_0078_));
 sg13g2_o21ai_1 _1931_ (.B1(net319),
    .Y(_1038_),
    .A1(_0517_),
    .A2(\game1.obstacle2_x[1] ));
 sg13g2_nor2_2 _1932_ (.A(net319),
    .B(net359),
    .Y(_1039_));
 sg13g2_nand2_2 _1933_ (.Y(_1040_),
    .A(net258),
    .B(_1039_));
 sg13g2_a21oi_1 _1934_ (.A1(net320),
    .A2(_1040_),
    .Y(_0079_),
    .B1(net222));
 sg13g2_xnor2_1 _1935_ (.Y(_1041_),
    .A(_0520_),
    .B(_1040_));
 sg13g2_nor2_1 _1936_ (.A(net222),
    .B(_1041_),
    .Y(_0080_));
 sg13g2_nand2_1 _1937_ (.Y(_1042_),
    .A(net361),
    .B(_1040_));
 sg13g2_nand3_1 _1938_ (.B(_0744_),
    .C(_1039_),
    .A(net258),
    .Y(_1043_));
 sg13g2_a21oi_1 _1939_ (.A1(_1042_),
    .A2(_1043_),
    .Y(_0081_),
    .B1(net223));
 sg13g2_nand3_1 _1940_ (.B(_0728_),
    .C(_1039_),
    .A(net258),
    .Y(_1044_));
 sg13g2_o21ai_1 _1941_ (.B1(net366),
    .Y(_1045_),
    .A1(_0727_),
    .A2(_1040_));
 sg13g2_a21oi_1 _1942_ (.A1(_1044_),
    .A2(_1045_),
    .Y(_0082_),
    .B1(net223));
 sg13g2_xnor2_1 _1943_ (.Y(_1046_),
    .A(_0519_),
    .B(_1044_));
 sg13g2_nor2_1 _1944_ (.A(net223),
    .B(_1046_),
    .Y(_0083_));
 sg13g2_nor4_1 _1945_ (.A(\game1.obstacle2_x[8] ),
    .B(\game1.obstacle2_x[3] ),
    .C(\game1.obstacle2_x[2] ),
    .D(_0521_),
    .Y(_1047_));
 sg13g2_nand2b_1 _1946_ (.Y(_1048_),
    .B(_1047_),
    .A_N(_0729_));
 sg13g2_nand3_1 _1947_ (.B(_0728_),
    .C(_1039_),
    .A(_0519_),
    .Y(_1049_));
 sg13g2_nor3_1 _1948_ (.A(\game1.obstacle2_x[8] ),
    .B(net260),
    .C(_1049_),
    .Y(_1050_));
 sg13g2_xnor2_1 _1949_ (.Y(_1051_),
    .A(_0033_),
    .B(_1050_));
 sg13g2_xnor2_1 _1950_ (.Y(_1052_),
    .A(net260),
    .B(_1049_));
 sg13g2_nor2_1 _1951_ (.A(_0517_),
    .B(_1052_),
    .Y(_1053_));
 sg13g2_o21ai_1 _1952_ (.B1(_1053_),
    .Y(_1054_),
    .A1(_1048_),
    .A2(_1051_));
 sg13g2_o21ai_1 _1953_ (.B1(_1054_),
    .Y(_1055_),
    .A1(net258),
    .A2(net260));
 sg13g2_nand2_1 _1954_ (.Y(_0084_),
    .A(net220),
    .B(net435));
 sg13g2_nor3_1 _1955_ (.A(net260),
    .B(_0729_),
    .C(_1040_),
    .Y(_1056_));
 sg13g2_xnor2_1 _1956_ (.Y(_1057_),
    .A(net391),
    .B(_1056_));
 sg13g2_nor2_1 _1957_ (.A(net222),
    .B(_1057_),
    .Y(_0085_));
 sg13g2_nor2_1 _1958_ (.A(net326),
    .B(net258),
    .Y(_1058_));
 sg13g2_o21ai_1 _1959_ (.B1(net258),
    .Y(_1059_),
    .A1(_1048_),
    .A2(_1052_));
 sg13g2_nor2_1 _1960_ (.A(_1051_),
    .B(_1059_),
    .Y(_1060_));
 sg13g2_o21ai_1 _1961_ (.B1(net220),
    .Y(_0086_),
    .A1(net327),
    .A2(_1060_));
 sg13g2_o21ai_1 _1962_ (.B1(\game1.scroll1_h_inst.ctr[7] ),
    .Y(_1061_),
    .A1(\game1.scroll1_h_inst.ctr[6] ),
    .A2(\game1.scroll1_h_inst.ctr[5] ));
 sg13g2_nand2b_1 _1963_ (.Y(_1062_),
    .B(_1061_),
    .A_N(\game1.scroll1_h_inst.ctr[8] ));
 sg13g2_nand3_1 _1964_ (.B(\game1.scroll1_h_inst.ctr[9] ),
    .C(_1062_),
    .A(\game1.scroll1_h_inst.ctr[10] ),
    .Y(_1063_));
 sg13g2_nor4_1 _1965_ (.A(\game1.scroll1_h_inst.ctr[14] ),
    .B(\game1.scroll1_h_inst.ctr[13] ),
    .C(\game1.scroll1_h_inst.ctr[12] ),
    .D(\game1.scroll1_h_inst.ctr[11] ),
    .Y(_1064_));
 sg13g2_nand2_1 _1966_ (.Y(_1065_),
    .A(\game1.scroll1_h_inst.ctr[15] ),
    .B(\game1.scroll1_h_inst.ctr[16] ));
 sg13g2_a21oi_1 _1967_ (.A1(_1063_),
    .A2(_1064_),
    .Y(_1066_),
    .B1(_1065_));
 sg13g2_nor2_1 _1968_ (.A(net433),
    .B(_1066_),
    .Y(_1067_));
 sg13g2_nor2_1 _1969_ (.A(net226),
    .B(_1067_),
    .Y(_0103_));
 sg13g2_nand2_1 _1970_ (.Y(_1068_),
    .A(net255),
    .B(net214));
 sg13g2_nor2b_2 _1971_ (.A(net226),
    .B_N(net231),
    .Y(_1069_));
 sg13g2_nand2_1 _1972_ (.Y(_1070_),
    .A(net221),
    .B(net231));
 sg13g2_and3_1 _1973_ (.X(_1071_),
    .A(net160),
    .B(\game1.scroll1_h_inst.ctr[1] ),
    .C(\game1.scroll1_h_inst.ctr[0] ));
 sg13g2_and2_1 _1974_ (.A(net175),
    .B(_1071_),
    .X(_1072_));
 sg13g2_and2_1 _1975_ (.A(net167),
    .B(_1072_),
    .X(_1073_));
 sg13g2_and2_1 _1976_ (.A(net188),
    .B(_1073_),
    .X(_1074_));
 sg13g2_and2_1 _1977_ (.A(net195),
    .B(_1074_),
    .X(_1075_));
 sg13g2_and2_1 _1978_ (.A(net193),
    .B(_1075_),
    .X(_1076_));
 sg13g2_and2_1 _1979_ (.A(net178),
    .B(_1076_),
    .X(_1077_));
 sg13g2_xnor2_1 _1980_ (.Y(_1078_),
    .A(net339),
    .B(_1077_));
 sg13g2_o21ai_1 _1981_ (.B1(_1068_),
    .Y(_0087_),
    .A1(net213),
    .A2(_1078_));
 sg13g2_nand2_1 _1982_ (.Y(_1079_),
    .A(net208),
    .B(net214));
 sg13g2_a21oi_1 _1983_ (.A1(\game1.scroll1_h_inst.ctr[9] ),
    .A2(_1077_),
    .Y(_1080_),
    .B1(net295));
 sg13g2_and3_1 _1984_ (.X(_1081_),
    .A(\game1.scroll1_h_inst.ctr[10] ),
    .B(\game1.scroll1_h_inst.ctr[9] ),
    .C(_1077_));
 sg13g2_or2_1 _1985_ (.X(_1082_),
    .B(_1081_),
    .A(net296));
 sg13g2_o21ai_1 _1986_ (.B1(_1079_),
    .Y(_0088_),
    .A1(net213),
    .A2(_1082_));
 sg13g2_nand2_1 _1987_ (.Y(_1083_),
    .A(net292),
    .B(net214));
 sg13g2_and2_1 _1988_ (.A(\game1.scroll1_h_inst.ctr[11] ),
    .B(_1081_),
    .X(_1084_));
 sg13g2_xnor2_1 _1989_ (.Y(_1085_),
    .A(\game1.scroll1_h_inst.ctr[11] ),
    .B(_1081_));
 sg13g2_o21ai_1 _1990_ (.B1(_1083_),
    .Y(_0089_),
    .A1(net213),
    .A2(_1085_));
 sg13g2_nand2_1 _1991_ (.Y(_1086_),
    .A(net254),
    .B(net214));
 sg13g2_xnor2_1 _1992_ (.Y(_1087_),
    .A(net340),
    .B(_1084_));
 sg13g2_o21ai_1 _1993_ (.B1(_1086_),
    .Y(_0090_),
    .A1(net213),
    .A2(net341));
 sg13g2_nand2_1 _1994_ (.Y(_1088_),
    .A(net253),
    .B(net214));
 sg13g2_nand3_1 _1995_ (.B(net340),
    .C(_1084_),
    .A(net393),
    .Y(_1089_));
 sg13g2_a21o_1 _1996_ (.A2(_1084_),
    .A1(net340),
    .B1(net393),
    .X(_1090_));
 sg13g2_nand2_1 _1997_ (.Y(_1091_),
    .A(_1089_),
    .B(_1090_));
 sg13g2_o21ai_1 _1998_ (.B1(_1088_),
    .Y(_0091_),
    .A1(net213),
    .A2(_1091_));
 sg13g2_nand2_1 _1999_ (.Y(_1092_),
    .A(net252),
    .B(net214));
 sg13g2_nor2_1 _2000_ (.A(_0559_),
    .B(_1089_),
    .Y(_1093_));
 sg13g2_xnor2_1 _2001_ (.Y(_1094_),
    .A(_0559_),
    .B(_1089_));
 sg13g2_o21ai_1 _2002_ (.B1(_1092_),
    .Y(_0092_),
    .A1(net213),
    .A2(net389));
 sg13g2_and2_1 _2003_ (.A(net313),
    .B(net214),
    .X(_1095_));
 sg13g2_nand2_1 _2004_ (.Y(_1096_),
    .A(\game1.scroll1_h_inst.ctr[15] ),
    .B(_1093_));
 sg13g2_xor2_1 _2005_ (.B(_1093_),
    .A(net400),
    .X(_1097_));
 sg13g2_a21o_1 _2006_ (.A2(_1097_),
    .A1(_1069_),
    .B1(_1095_),
    .X(_0093_));
 sg13g2_nor2b_1 _2007_ (.A(net231),
    .B_N(net283),
    .Y(_1098_));
 sg13g2_nand2_1 _2008_ (.Y(_1099_),
    .A(\game1.obstacle1_x[2] ),
    .B(\game1.obstacle1_x[1] ));
 sg13g2_nand4_1 _2009_ (.B(\game1.obstacle1_x[5] ),
    .C(\game1.obstacle1_x[4] ),
    .A(\game1.obstacle1_x[6] ),
    .Y(_1100_),
    .D(\game1.obstacle1_x[3] ));
 sg13g2_nor2_2 _2010_ (.A(_1099_),
    .B(_1100_),
    .Y(_1101_));
 sg13g2_o21ai_1 _2011_ (.B1(\game1.obstacle1_x[7] ),
    .Y(_1102_),
    .A1(_1099_),
    .A2(_1100_));
 sg13g2_nand3_1 _2012_ (.B(\game1.obstacle1_x[7] ),
    .C(_1101_),
    .A(\game1.obstacle1_x[8] ),
    .Y(_1103_));
 sg13g2_a21o_1 _2013_ (.A2(_1101_),
    .A1(net259),
    .B1(\game1.obstacle1_x[8] ),
    .X(_1104_));
 sg13g2_nand2_1 _2014_ (.Y(_1105_),
    .A(_1103_),
    .B(_1104_));
 sg13g2_xnor2_1 _2015_ (.Y(_1106_),
    .A(_0512_),
    .B(_1103_));
 sg13g2_a21oi_1 _2016_ (.A1(_1102_),
    .A2(_1105_),
    .Y(_1107_),
    .B1(_1106_));
 sg13g2_nor2_1 _2017_ (.A(net231),
    .B(_1107_),
    .Y(_1108_));
 sg13g2_nor2_1 _2018_ (.A(net283),
    .B(_1108_),
    .Y(_1109_));
 sg13g2_nor3_1 _2019_ (.A(net227),
    .B(_1098_),
    .C(_1109_),
    .Y(_0094_));
 sg13g2_nor2_1 _2020_ (.A(_0017_),
    .B(_1103_),
    .Y(_1110_));
 sg13g2_nand2b_1 _2021_ (.Y(_1111_),
    .B(_1101_),
    .A_N(net259));
 sg13g2_nor3_1 _2022_ (.A(_0512_),
    .B(\game1.obstacle1_x[8] ),
    .C(_1111_),
    .Y(_1112_));
 sg13g2_nor3_1 _2023_ (.A(_1107_),
    .B(_1110_),
    .C(_1112_),
    .Y(_1113_));
 sg13g2_or2_2 _2024_ (.X(_1114_),
    .B(_1113_),
    .A(net231));
 sg13g2_nor2_1 _2025_ (.A(net231),
    .B(_1099_),
    .Y(_1115_));
 sg13g2_xor2_1 _2026_ (.B(_1098_),
    .A(net424),
    .X(_1116_));
 sg13g2_a21o_1 _2027_ (.A2(_1116_),
    .A1(_1114_),
    .B1(net227),
    .X(_0095_));
 sg13g2_and2_1 _2028_ (.A(\game1.obstacle1_x[3] ),
    .B(_1115_),
    .X(_1117_));
 sg13g2_o21ai_1 _2029_ (.B1(_1114_),
    .Y(_1118_),
    .A1(net430),
    .A2(_1115_));
 sg13g2_o21ai_1 _2030_ (.B1(net221),
    .Y(_0096_),
    .A1(_1117_),
    .A2(_1118_));
 sg13g2_and2_1 _2031_ (.A(\game1.obstacle1_x[4] ),
    .B(_1117_),
    .X(_1119_));
 sg13g2_o21ai_1 _2032_ (.B1(_1114_),
    .Y(_1120_),
    .A1(net431),
    .A2(_1117_));
 sg13g2_o21ai_1 _2033_ (.B1(net221),
    .Y(_0097_),
    .A1(_1119_),
    .A2(_1120_));
 sg13g2_nor2_1 _2034_ (.A(net414),
    .B(_1119_),
    .Y(_1121_));
 sg13g2_nand2_1 _2035_ (.Y(_1122_),
    .A(\game1.obstacle1_x[5] ),
    .B(_1119_));
 sg13g2_nand2_1 _2036_ (.Y(_1123_),
    .A(_1114_),
    .B(_1122_));
 sg13g2_o21ai_1 _2037_ (.B1(net221),
    .Y(_0098_),
    .A1(_1121_),
    .A2(_1123_));
 sg13g2_xnor2_1 _2038_ (.Y(_1124_),
    .A(net425),
    .B(_1122_));
 sg13g2_a21o_1 _2039_ (.A2(_1124_),
    .A1(_1114_),
    .B1(net227),
    .X(_0099_));
 sg13g2_nand2_1 _2040_ (.Y(_1125_),
    .A(net259),
    .B(_1069_));
 sg13g2_xnor2_1 _2041_ (.Y(_1126_),
    .A(net259),
    .B(_1101_));
 sg13g2_nand2_1 _2042_ (.Y(_1127_),
    .A(_0103_),
    .B(_1113_));
 sg13g2_o21ai_1 _2043_ (.B1(_1125_),
    .Y(_0100_),
    .A1(_1126_),
    .A2(_1127_));
 sg13g2_nand2_1 _2044_ (.Y(_1128_),
    .A(net432),
    .B(net231));
 sg13g2_o21ai_1 _2045_ (.B1(_1128_),
    .Y(_1129_),
    .A1(net231),
    .A2(_1105_));
 sg13g2_a21o_1 _2046_ (.A2(_1129_),
    .A1(_1114_),
    .B1(net227),
    .X(_0101_));
 sg13g2_nand2_1 _2047_ (.Y(_0168_),
    .A(net183),
    .B(_1069_));
 sg13g2_o21ai_1 _2048_ (.B1(_0168_),
    .Y(_0102_),
    .A1(_1106_),
    .A2(_1127_));
 sg13g2_nand3_1 _2049_ (.B(\game1.obstacle2_y[2] ),
    .C(\game1.obstacle2_y[1] ),
    .A(\game1.obstacle2_y[3] ),
    .Y(_0169_));
 sg13g2_or2_2 _2050_ (.X(_0170_),
    .B(_0169_),
    .A(_0511_));
 sg13g2_nand2_1 _2051_ (.Y(_0171_),
    .A(\game1.obstacle2_y[6] ),
    .B(\game1.obstacle2_y[5] ));
 sg13g2_nor2_1 _2052_ (.A(_0170_),
    .B(_0171_),
    .Y(_0172_));
 sg13g2_nand2_1 _2053_ (.Y(_0173_),
    .A(\game1.obstacle2_y[7] ),
    .B(_0172_));
 sg13g2_xnor2_1 _2054_ (.Y(_0174_),
    .A(_0508_),
    .B(_0172_));
 sg13g2_nor2_1 _2055_ (.A(_0036_),
    .B(_0170_),
    .Y(_0175_));
 sg13g2_xor2_1 _2056_ (.B(_0170_),
    .A(_0036_),
    .X(_0176_));
 sg13g2_nor2_1 _2057_ (.A(_0035_),
    .B(_0034_),
    .Y(_0177_));
 sg13g2_and3_1 _2058_ (.X(_0178_),
    .A(_0174_),
    .B(_0176_),
    .C(_0177_));
 sg13g2_nor3_1 _2059_ (.A(_0721_),
    .B(_0170_),
    .C(_0171_),
    .Y(_0179_));
 sg13g2_nor4_2 _2060_ (.A(\game1.obstacle2_y[9] ),
    .B(net235),
    .C(_0178_),
    .Y(_0180_),
    .D(_0179_));
 sg13g2_nand2b_1 _2061_ (.Y(_0181_),
    .B(_0180_),
    .A_N(net256));
 sg13g2_nand2_1 _2062_ (.Y(_0182_),
    .A(net235),
    .B(net256));
 sg13g2_a21oi_1 _2063_ (.A1(_0181_),
    .A2(_0182_),
    .Y(_0104_),
    .B1(net224));
 sg13g2_a22oi_1 _2064_ (.Y(_0183_),
    .B1(_0700_),
    .B2(_0180_),
    .A2(net378),
    .A1(net235));
 sg13g2_nor2_1 _2065_ (.A(net230),
    .B(net379),
    .Y(_0105_));
 sg13g2_a21o_1 _2066_ (.A2(net256),
    .A1(\game1.obstacle2_y[2] ),
    .B1(\game1.obstacle2_y[3] ),
    .X(_0184_));
 sg13g2_and2_1 _2067_ (.A(_0169_),
    .B(_0184_),
    .X(_0185_));
 sg13g2_a22oi_1 _2068_ (.Y(_0186_),
    .B1(_0180_),
    .B2(_0185_),
    .A2(net352),
    .A1(net235));
 sg13g2_nor2_1 _2069_ (.A(net224),
    .B(net353),
    .Y(_0106_));
 sg13g2_xnor2_1 _2070_ (.Y(_0187_),
    .A(net337),
    .B(_0169_));
 sg13g2_a22oi_1 _2071_ (.Y(_0188_),
    .B1(_0180_),
    .B2(_0187_),
    .A2(net337),
    .A1(net235));
 sg13g2_nor2_1 _2072_ (.A(net224),
    .B(net338),
    .Y(_0107_));
 sg13g2_a22oi_1 _2073_ (.Y(_0189_),
    .B1(_0176_),
    .B2(_0180_),
    .A2(net335),
    .A1(net235));
 sg13g2_nor2_1 _2074_ (.A(net224),
    .B(net336),
    .Y(_0108_));
 sg13g2_xnor2_1 _2075_ (.Y(_0190_),
    .A(net343),
    .B(_0175_));
 sg13g2_a22oi_1 _2076_ (.Y(_0191_),
    .B1(_0180_),
    .B2(net344),
    .A2(\game1.obstacle2_y[6] ),
    .A1(_0506_));
 sg13g2_nor2_1 _2077_ (.A(net224),
    .B(net345),
    .Y(_0109_));
 sg13g2_a22oi_1 _2078_ (.Y(_0192_),
    .B1(_0174_),
    .B2(_0180_),
    .A2(net376),
    .A1(net235));
 sg13g2_nor2_1 _2079_ (.A(net224),
    .B(net377),
    .Y(_0110_));
 sg13g2_xor2_1 _2080_ (.B(_0173_),
    .A(_0034_),
    .X(_0193_));
 sg13g2_a22oi_1 _2081_ (.Y(_0194_),
    .B1(_0180_),
    .B2(_0193_),
    .A2(net303),
    .A1(net235));
 sg13g2_nor2_1 _2082_ (.A(net224),
    .B(net304),
    .Y(_0111_));
 sg13g2_nor3_1 _2083_ (.A(_0505_),
    .B(net165),
    .C(net224),
    .Y(_0112_));
 sg13g2_and2_2 _2084_ (.A(\game1.score[6] ),
    .B(\game1.score[5] ),
    .X(_0195_));
 sg13g2_nand3b_1 _2085_ (.B(net252),
    .C(\game1.score[6] ),
    .Y(_0196_),
    .A_N(net253));
 sg13g2_nor2_1 _2086_ (.A(net252),
    .B(net253),
    .Y(_0197_));
 sg13g2_o21ai_1 _2087_ (.B1(\game1.score[6] ),
    .Y(_0198_),
    .A1(net252),
    .A2(\game1.score[4] ));
 sg13g2_a22oi_1 _2088_ (.Y(_0199_),
    .B1(_0198_),
    .B2(_0561_),
    .A2(_0195_),
    .A1(_0503_));
 sg13g2_and2_1 _2089_ (.A(\game1.score[6] ),
    .B(_0197_),
    .X(_0200_));
 sg13g2_nand2_1 _2090_ (.Y(_0201_),
    .A(\game1.score[6] ),
    .B(_0197_));
 sg13g2_a22oi_1 _2091_ (.Y(_0202_),
    .B1(_0198_),
    .B2(_0560_),
    .A2(_0195_),
    .A1(net253));
 sg13g2_or2_1 _2092_ (.X(_0203_),
    .B(_0202_),
    .A(_0199_));
 sg13g2_nand2_1 _2093_ (.Y(_0204_),
    .A(net252),
    .B(_0196_));
 sg13g2_nand2b_1 _2094_ (.Y(_0205_),
    .B(net253),
    .A_N(\game1.score[6] ));
 sg13g2_nand4_1 _2095_ (.B(net254),
    .C(_0196_),
    .A(net252),
    .Y(_0206_),
    .D(_0205_));
 sg13g2_o21ai_1 _2096_ (.B1(_0206_),
    .Y(_0207_),
    .A1(_0199_),
    .A2(_0202_));
 sg13g2_nand2b_1 _2097_ (.Y(_0208_),
    .B(_0201_),
    .A_N(_0207_));
 sg13g2_o21ai_1 _2098_ (.B1(_0504_),
    .Y(_0209_),
    .A1(_0200_),
    .A2(_0207_));
 sg13g2_xor2_1 _2099_ (.B(_0209_),
    .A(_0199_),
    .X(_0210_));
 sg13g2_nand4_1 _2100_ (.B(_0201_),
    .C(_0203_),
    .A(net254),
    .Y(_0211_),
    .D(_0206_));
 sg13g2_and2_1 _2101_ (.A(_0209_),
    .B(_0211_),
    .X(_0212_));
 sg13g2_nand3_1 _2102_ (.B(_0209_),
    .C(_0211_),
    .A(_0008_),
    .Y(_0213_));
 sg13g2_nand3_1 _2103_ (.B(_0196_),
    .C(_0205_),
    .A(_0504_),
    .Y(_0214_));
 sg13g2_xnor2_1 _2104_ (.Y(_0215_),
    .A(_0202_),
    .B(_0214_));
 sg13g2_o21ai_1 _2105_ (.B1(_0215_),
    .Y(_0216_),
    .A1(_0200_),
    .A2(_0207_));
 sg13g2_nor3_1 _2106_ (.A(_0200_),
    .B(_0204_),
    .C(_0207_),
    .Y(_0217_));
 sg13g2_a21oi_1 _2107_ (.A1(_0208_),
    .A2(_0215_),
    .Y(_0218_),
    .B1(_0217_));
 sg13g2_nand3_1 _2108_ (.B(_0213_),
    .C(_0218_),
    .A(_0210_),
    .Y(_0219_));
 sg13g2_nor2_1 _2109_ (.A(_0201_),
    .B(_0203_),
    .Y(_0220_));
 sg13g2_o21ai_1 _2110_ (.B1(_0216_),
    .Y(_0221_),
    .A1(_0202_),
    .A2(_0208_));
 sg13g2_nor2_2 _2111_ (.A(_0220_),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_or2_1 _2112_ (.X(_0223_),
    .B(_0221_),
    .A(_0220_));
 sg13g2_nand2_1 _2113_ (.Y(_0224_),
    .A(_0219_),
    .B(_0222_));
 sg13g2_a21o_1 _2114_ (.A2(_0222_),
    .A1(_0219_),
    .B1(_0008_),
    .X(_0225_));
 sg13g2_nand3_1 _2115_ (.B(_0219_),
    .C(_0222_),
    .A(_0008_),
    .Y(_0226_));
 sg13g2_nand2_1 _2116_ (.Y(_0227_),
    .A(_0225_),
    .B(_0226_));
 sg13g2_and2_1 _2117_ (.A(_0225_),
    .B(_0226_),
    .X(_0228_));
 sg13g2_a21o_1 _2118_ (.A2(_0226_),
    .A1(_0225_),
    .B1(\game1.score[1] ),
    .X(_0229_));
 sg13g2_a21oi_1 _2119_ (.A1(_0219_),
    .A2(_0222_),
    .Y(_0230_),
    .B1(\game1.score[2] ));
 sg13g2_xnor2_1 _2120_ (.Y(_0231_),
    .A(_0212_),
    .B(_0230_));
 sg13g2_nand2b_1 _2121_ (.Y(_0232_),
    .B(_0221_),
    .A_N(_0213_));
 sg13g2_nand3b_1 _2122_ (.B(_0223_),
    .C(_0232_),
    .Y(_0233_),
    .A_N(_0210_));
 sg13g2_or2_1 _2123_ (.X(_0234_),
    .B(_0221_),
    .A(_0218_));
 sg13g2_a21oi_1 _2124_ (.A1(_0210_),
    .A2(_0219_),
    .Y(_0235_),
    .B1(_0220_));
 sg13g2_nand3_1 _2125_ (.B(_0234_),
    .C(_0235_),
    .A(_0233_),
    .Y(_0236_));
 sg13g2_a21oi_1 _2126_ (.A1(_0229_),
    .A2(_0236_),
    .Y(_0237_),
    .B1(_0231_));
 sg13g2_a21o_1 _2127_ (.A2(_0231_),
    .A1(_0229_),
    .B1(_0237_),
    .X(_0238_));
 sg13g2_a21oi_2 _2128_ (.B1(_0236_),
    .Y(_0239_),
    .A2(_0231_),
    .A1(_0229_));
 sg13g2_a21o_2 _2129_ (.A2(_0231_),
    .A1(_0229_),
    .B1(_0236_),
    .X(_0240_));
 sg13g2_a21oi_1 _2130_ (.A1(_0009_),
    .A2(_0240_),
    .Y(_0241_),
    .B1(_0228_));
 sg13g2_o21ai_1 _2131_ (.B1(_0227_),
    .Y(_0242_),
    .A1(_0563_),
    .A2(_0239_));
 sg13g2_nor3_1 _2132_ (.A(_0563_),
    .B(_0227_),
    .C(_0239_),
    .Y(_0243_));
 sg13g2_nand3_1 _2133_ (.B(_0228_),
    .C(_0240_),
    .A(_0009_),
    .Y(_0244_));
 sg13g2_o21ai_1 _2134_ (.B1(_0238_),
    .Y(_0245_),
    .A1(_0241_),
    .A2(_0243_));
 sg13g2_xnor2_1 _2135_ (.Y(_0246_),
    .A(_0563_),
    .B(_0239_));
 sg13g2_or2_1 _2136_ (.X(_0247_),
    .B(_0246_),
    .A(_0039_));
 sg13g2_nor2_1 _2137_ (.A(_0245_),
    .B(_0247_),
    .Y(_0248_));
 sg13g2_nor2_1 _2138_ (.A(net255),
    .B(_0246_),
    .Y(_0249_));
 sg13g2_a21oi_1 _2139_ (.A1(net255),
    .A2(_0039_),
    .Y(_0250_),
    .B1(_0246_));
 sg13g2_a21oi_1 _2140_ (.A1(_0242_),
    .A2(_0244_),
    .Y(_0251_),
    .B1(_0238_));
 sg13g2_and2_1 _2141_ (.A(_0250_),
    .B(_0251_),
    .X(_0252_));
 sg13g2_nand2_1 _2142_ (.Y(_0253_),
    .A(net255),
    .B(_0246_));
 sg13g2_and2_1 _2143_ (.A(_0039_),
    .B(_0246_),
    .X(_0254_));
 sg13g2_a21o_1 _2144_ (.A2(_0246_),
    .A1(net255),
    .B1(_0254_),
    .X(_0255_));
 sg13g2_nand3_1 _2145_ (.B(_0242_),
    .C(_0244_),
    .A(_0238_),
    .Y(_0256_));
 sg13g2_nor2_1 _2146_ (.A(_0253_),
    .B(_0256_),
    .Y(_0257_));
 sg13g2_nor2_1 _2147_ (.A(_0245_),
    .B(_0253_),
    .Y(_0258_));
 sg13g2_and2_1 _2148_ (.A(_0238_),
    .B(_0254_),
    .X(_0259_));
 sg13g2_nand2b_1 _2149_ (.Y(_0260_),
    .B(_0256_),
    .A_N(_0251_));
 sg13g2_a221oi_1 _2150_ (.B2(_0250_),
    .C1(_0248_),
    .B1(_0260_),
    .A1(_0238_),
    .Y(_0261_),
    .A2(_0255_));
 sg13g2_nand2_2 _2151_ (.Y(_0262_),
    .A(net262),
    .B(_0593_));
 sg13g2_nor2_1 _2152_ (.A(_0569_),
    .B(_0594_),
    .Y(_0263_));
 sg13g2_nand4_1 _2153_ (.B(net268),
    .C(_0022_),
    .A(net266),
    .Y(_0264_),
    .D(_0593_));
 sg13g2_nand4_1 _2154_ (.B(net266),
    .C(_0897_),
    .A(net273),
    .Y(_0265_),
    .D(_0905_));
 sg13g2_nor2_1 _2155_ (.A(\game1.pixel_x[1] ),
    .B(\game1.pixel_x[2] ),
    .Y(_0266_));
 sg13g2_nor3_1 _2156_ (.A(_0569_),
    .B(_0594_),
    .C(_0266_),
    .Y(_0267_));
 sg13g2_nor2b_1 _2157_ (.A(net271),
    .B_N(net273),
    .Y(_0268_));
 sg13g2_a221oi_1 _2158_ (.B2(_0268_),
    .C1(_0262_),
    .B1(_0267_),
    .A1(_0264_),
    .Y(_0269_),
    .A2(_0265_));
 sg13g2_and2_1 _2159_ (.A(net271),
    .B(_0269_),
    .X(_0270_));
 sg13g2_xnor2_1 _2160_ (.Y(_0271_),
    .A(net270),
    .B(_0269_));
 sg13g2_xor2_1 _2161_ (.B(_0269_),
    .A(_0022_),
    .X(_0272_));
 sg13g2_a21oi_1 _2162_ (.A1(net273),
    .A2(_0271_),
    .Y(_0273_),
    .B1(_0270_));
 sg13g2_a21o_1 _2163_ (.A2(_0271_),
    .A1(net273),
    .B1(_0270_),
    .X(_0274_));
 sg13g2_nor2b_1 _2164_ (.A(_0270_),
    .B_N(_0266_),
    .Y(_0275_));
 sg13g2_nor3_2 _2165_ (.A(_0569_),
    .B(_0273_),
    .C(_0275_),
    .Y(_0276_));
 sg13g2_o21ai_1 _2166_ (.B1(_0593_),
    .Y(_0277_),
    .A1(_0569_),
    .A2(_0273_));
 sg13g2_a21o_1 _2167_ (.A2(_0272_),
    .A1(_1016_),
    .B1(net271),
    .X(_0278_));
 sg13g2_a21oi_1 _2168_ (.A1(_0549_),
    .A2(_0278_),
    .Y(_0279_),
    .B1(_0269_));
 sg13g2_a21o_1 _2169_ (.A2(_0278_),
    .A1(_0549_),
    .B1(_0269_),
    .X(_0280_));
 sg13g2_nand3_1 _2170_ (.B(_1016_),
    .C(_0272_),
    .A(_0021_),
    .Y(_0281_));
 sg13g2_and2_1 _2171_ (.A(_0545_),
    .B(_0269_),
    .X(_0282_));
 sg13g2_a21oi_1 _2172_ (.A1(_0281_),
    .A2(_0282_),
    .Y(_0283_),
    .B1(_0020_));
 sg13g2_a21o_1 _2173_ (.A2(_0282_),
    .A1(_0281_),
    .B1(_0020_),
    .X(_0284_));
 sg13g2_nor4_2 _2174_ (.A(_0262_),
    .B(_0276_),
    .C(_0279_),
    .Y(_0285_),
    .D(_0284_));
 sg13g2_nor2_1 _2175_ (.A(net237),
    .B(net238),
    .Y(_0286_));
 sg13g2_nor2_1 _2176_ (.A(net240),
    .B(net242),
    .Y(_0287_));
 sg13g2_nor3_1 _2177_ (.A(net240),
    .B(net242),
    .C(net244),
    .Y(_0288_));
 sg13g2_and2_1 _2178_ (.A(_0286_),
    .B(_0288_),
    .X(_0289_));
 sg13g2_nand2_1 _2179_ (.Y(_0290_),
    .A(_0551_),
    .B(_0577_));
 sg13g2_nand2_1 _2180_ (.Y(_0291_),
    .A(_0581_),
    .B(_0288_));
 sg13g2_inv_1 _2181_ (.Y(_0292_),
    .A(_0291_));
 sg13g2_o21ai_1 _2182_ (.B1(\game1.pixel_y[4] ),
    .Y(_0293_),
    .A1(_0290_),
    .A2(_0292_));
 sg13g2_and2_1 _2183_ (.A(_0289_),
    .B(_0293_),
    .X(_0294_));
 sg13g2_nand2_1 _2184_ (.Y(_0295_),
    .A(_0578_),
    .B(_0581_));
 sg13g2_nand2_1 _2185_ (.Y(_0296_),
    .A(_0576_),
    .B(_0578_));
 sg13g2_nand3_1 _2186_ (.B(_0576_),
    .C(_0578_),
    .A(\game1.pixel_y[4] ),
    .Y(_0297_));
 sg13g2_xnor2_1 _2187_ (.Y(_0298_),
    .A(_0556_),
    .B(_0296_));
 sg13g2_nand2_1 _2188_ (.Y(_0299_),
    .A(_0295_),
    .B(_0298_));
 sg13g2_and3_1 _2189_ (.X(_0300_),
    .A(_0285_),
    .B(_0294_),
    .C(_0299_));
 sg13g2_a21oi_2 _2190_ (.B1(_0594_),
    .Y(_0301_),
    .A2(_0283_),
    .A1(_0280_));
 sg13g2_nor2_1 _2191_ (.A(net273),
    .B(_0272_),
    .Y(_0302_));
 sg13g2_nor2b_1 _2192_ (.A(_0569_),
    .B_N(_0897_),
    .Y(_0303_));
 sg13g2_a221oi_1 _2193_ (.B2(_0303_),
    .C1(_0594_),
    .B1(_0302_),
    .A1(_0263_),
    .Y(_0304_),
    .A2(_0274_));
 sg13g2_a21o_1 _2194_ (.A2(_0286_),
    .A1(net251),
    .B1(_0290_),
    .X(_0305_));
 sg13g2_and2_1 _2195_ (.A(_0556_),
    .B(_0288_),
    .X(_0306_));
 sg13g2_inv_1 _2196_ (.Y(_0307_),
    .A(_0306_));
 sg13g2_a21oi_1 _2197_ (.A1(net251),
    .A2(net248),
    .Y(_0308_),
    .B1(net246));
 sg13g2_nand3_1 _2198_ (.B(_0306_),
    .C(_0308_),
    .A(_0286_),
    .Y(_0309_));
 sg13g2_nor2b_1 _2199_ (.A(_0309_),
    .B_N(_0305_),
    .Y(_0310_));
 sg13g2_inv_1 _2200_ (.Y(_0311_),
    .A(_0310_));
 sg13g2_nand2_1 _2201_ (.Y(_0312_),
    .A(_0304_),
    .B(_0310_));
 sg13g2_nor3_2 _2202_ (.A(net234),
    .B(_0301_),
    .C(_0312_),
    .Y(_0313_));
 sg13g2_or3_1 _2203_ (.A(net234),
    .B(_0301_),
    .C(_0312_),
    .X(_0314_));
 sg13g2_nand3_1 _2204_ (.B(_0295_),
    .C(_0297_),
    .A(_0289_),
    .Y(_0315_));
 sg13g2_nand2_1 _2205_ (.Y(_0316_),
    .A(_0577_),
    .B(_0291_));
 sg13g2_nand3_1 _2206_ (.B(net245),
    .C(_0316_),
    .A(net246),
    .Y(_0317_));
 sg13g2_nor2_1 _2207_ (.A(_0315_),
    .B(_0317_),
    .Y(_0318_));
 sg13g2_and2_1 _2208_ (.A(_0285_),
    .B(_0318_),
    .X(_0319_));
 sg13g2_nand2_1 _2209_ (.Y(_0320_),
    .A(_0285_),
    .B(_0318_));
 sg13g2_o21ai_1 _2210_ (.B1(_0294_),
    .Y(_0321_),
    .A1(_0305_),
    .A2(_0307_));
 sg13g2_or3_1 _2211_ (.A(_0262_),
    .B(_0276_),
    .C(_0304_),
    .X(_0322_));
 sg13g2_nor2_2 _2212_ (.A(_0321_),
    .B(_0322_),
    .Y(_0323_));
 sg13g2_or2_1 _2213_ (.X(_0324_),
    .B(_0315_),
    .A(_0293_));
 sg13g2_or4_1 _2214_ (.A(_0262_),
    .B(_0276_),
    .C(_0304_),
    .D(_0324_),
    .X(_0325_));
 sg13g2_nor2b_1 _2215_ (.A(_0323_),
    .B_N(_0325_),
    .Y(_0326_));
 sg13g2_a21o_1 _2216_ (.A2(_0302_),
    .A1(_0267_),
    .B1(_0277_),
    .X(_0327_));
 sg13g2_nor3_1 _2217_ (.A(net234),
    .B(_0301_),
    .C(_0327_),
    .Y(_0328_));
 sg13g2_nor4_2 _2218_ (.A(net234),
    .B(_0301_),
    .C(_0321_),
    .Y(_0329_),
    .D(_0327_));
 sg13g2_nor2_1 _2219_ (.A(_0300_),
    .B(_0329_),
    .Y(_0330_));
 sg13g2_nand2_1 _2220_ (.Y(_0331_),
    .A(_0326_),
    .B(_0330_));
 sg13g2_nand2_1 _2221_ (.Y(_0332_),
    .A(_0289_),
    .B(_0317_));
 sg13g2_nor2b_1 _2222_ (.A(_0332_),
    .B_N(_0309_),
    .Y(_0333_));
 sg13g2_nand4_1 _2223_ (.B(_0304_),
    .C(_0327_),
    .A(net262),
    .Y(_0334_),
    .D(_0333_));
 sg13g2_o21ai_1 _2224_ (.B1(_0325_),
    .Y(_0335_),
    .A1(_0311_),
    .A2(_0322_));
 sg13g2_or4_1 _2225_ (.A(_0300_),
    .B(_0313_),
    .C(_0329_),
    .D(_0335_),
    .X(_0336_));
 sg13g2_nor2_1 _2226_ (.A(_0294_),
    .B(_0332_),
    .Y(_0337_));
 sg13g2_and2_1 _2227_ (.A(_0328_),
    .B(_0337_),
    .X(_0338_));
 sg13g2_a21oi_2 _2228_ (.B1(_0319_),
    .Y(_0339_),
    .A2(_0337_),
    .A1(_0328_));
 sg13g2_nor3_1 _2229_ (.A(net255),
    .B(_0246_),
    .C(_0339_),
    .Y(_0340_));
 sg13g2_or3_1 _2230_ (.A(_0323_),
    .B(_0336_),
    .C(_0340_),
    .X(_0341_));
 sg13g2_nand2b_1 _2231_ (.Y(_0342_),
    .B(_0320_),
    .A_N(_0300_));
 sg13g2_nor4_2 _2232_ (.A(_0313_),
    .B(_0323_),
    .C(_0338_),
    .Y(_0343_),
    .D(_0342_));
 sg13g2_inv_1 _2233_ (.Y(_0344_),
    .A(_0343_));
 sg13g2_a21oi_1 _2234_ (.A1(_0242_),
    .A2(_0244_),
    .Y(_0345_),
    .B1(_0343_));
 sg13g2_nor2_1 _2235_ (.A(_0319_),
    .B(_0336_),
    .Y(_0346_));
 sg13g2_nor3_1 _2236_ (.A(_0247_),
    .B(_0256_),
    .C(_0346_),
    .Y(_0347_));
 sg13g2_a221oi_1 _2237_ (.B2(_0259_),
    .C1(_0347_),
    .B1(_0345_),
    .A1(_0252_),
    .Y(_0348_),
    .A2(_0341_));
 sg13g2_nand2_2 _2238_ (.Y(_0349_),
    .A(_0314_),
    .B(_0326_));
 sg13g2_nand3_1 _2239_ (.B(_0320_),
    .C(_0334_),
    .A(_0314_),
    .Y(_0350_));
 sg13g2_a22oi_1 _2240_ (.Y(_0351_),
    .B1(_0350_),
    .B2(_0248_),
    .A2(_0349_),
    .A1(_0257_));
 sg13g2_nand2b_1 _2241_ (.Y(_0352_),
    .B(_0339_),
    .A_N(_0336_));
 sg13g2_a22oi_1 _2242_ (.Y(_0353_),
    .B1(_0352_),
    .B2(_0254_),
    .A2(_0331_),
    .A1(_0249_));
 sg13g2_or2_1 _2243_ (.X(_0354_),
    .B(_0353_),
    .A(_0256_));
 sg13g2_or2_1 _2244_ (.X(_0355_),
    .B(_0349_),
    .A(_0342_));
 sg13g2_nand2_1 _2245_ (.Y(_0356_),
    .A(_0258_),
    .B(_0355_));
 sg13g2_nand4_1 _2246_ (.B(_0351_),
    .C(_0354_),
    .A(_0348_),
    .Y(_0357_),
    .D(_0356_));
 sg13g2_nor2b_1 _2247_ (.A(_0329_),
    .B_N(_0339_),
    .Y(_0358_));
 sg13g2_nor2b_1 _2248_ (.A(_0349_),
    .B_N(_0358_),
    .Y(_0359_));
 sg13g2_nand2b_1 _2249_ (.Y(_0360_),
    .B(_0358_),
    .A_N(_0349_));
 sg13g2_nand2_1 _2250_ (.Y(_0361_),
    .A(_0546_),
    .B(_1016_));
 sg13g2_nor2_1 _2251_ (.A(_0569_),
    .B(_0262_),
    .Y(_0362_));
 sg13g2_o21ai_1 _2252_ (.B1(_0362_),
    .Y(_0363_),
    .A1(_0904_),
    .A2(_0266_));
 sg13g2_a221oi_1 _2253_ (.B2(net420),
    .C1(_0363_),
    .B1(_0361_),
    .A1(_0261_),
    .Y(_0364_),
    .A2(_0359_));
 sg13g2_o21ai_1 _2254_ (.B1(_0364_),
    .Y(_0365_),
    .A1(_0261_),
    .A2(_0357_));
 sg13g2_or2_1 _2255_ (.X(_0366_),
    .B(_0224_),
    .A(_0198_));
 sg13g2_nor2b_1 _2256_ (.A(_0366_),
    .B_N(_0207_),
    .Y(_0367_));
 sg13g2_a21oi_1 _2257_ (.A1(_0198_),
    .A2(_0224_),
    .Y(_0368_),
    .B1(_0367_));
 sg13g2_a21o_1 _2258_ (.A2(_0224_),
    .A1(_0198_),
    .B1(_0367_),
    .X(_0369_));
 sg13g2_and2_1 _2259_ (.A(_0208_),
    .B(_0366_),
    .X(_0370_));
 sg13g2_nand2_1 _2260_ (.Y(_0371_),
    .A(_0331_),
    .B(_0368_));
 sg13g2_or2_1 _2261_ (.X(_0372_),
    .B(_0366_),
    .A(_0207_));
 sg13g2_mux4_1 _2262_ (.S0(_0240_),
    .A0(_0344_),
    .A1(_0355_),
    .A2(_0360_),
    .A3(_0350_),
    .S1(_0368_),
    .X(_0373_));
 sg13g2_nand2b_1 _2263_ (.Y(_0374_),
    .B(_0373_),
    .A_N(_0370_));
 sg13g2_a21oi_1 _2264_ (.A1(_0349_),
    .A2(_0369_),
    .Y(_0375_),
    .B1(_0239_));
 sg13g2_o21ai_1 _2265_ (.B1(_0375_),
    .Y(_0376_),
    .A1(_0346_),
    .A2(_0369_));
 sg13g2_nand2_1 _2266_ (.Y(_0377_),
    .A(_0352_),
    .B(_0369_));
 sg13g2_nand3_1 _2267_ (.B(_0371_),
    .C(_0377_),
    .A(_0239_),
    .Y(_0378_));
 sg13g2_nand3_1 _2268_ (.B(_0376_),
    .C(_0378_),
    .A(_0370_),
    .Y(_0379_));
 sg13g2_nand3_1 _2269_ (.B(_0374_),
    .C(_0379_),
    .A(_0372_),
    .Y(_0380_));
 sg13g2_nor2_1 _2270_ (.A(_0240_),
    .B(_0339_),
    .Y(_0381_));
 sg13g2_or4_1 _2271_ (.A(_0323_),
    .B(_0336_),
    .C(_0372_),
    .D(_0381_),
    .X(_0382_));
 sg13g2_nand3_1 _2272_ (.B(_0380_),
    .C(_0382_),
    .A(_0269_),
    .Y(_0383_));
 sg13g2_or2_1 _2273_ (.X(_0384_),
    .B(_0592_),
    .A(_0030_));
 sg13g2_nand4_1 _2274_ (.B(_0286_),
    .C(_0287_),
    .A(net221),
    .Y(_0385_),
    .D(_0384_));
 sg13g2_a21oi_1 _2275_ (.A1(_0365_),
    .A2(_0383_),
    .Y(_0113_),
    .B1(_0385_));
 sg13g2_nand2b_1 _2276_ (.Y(_0386_),
    .B(\game1.scroll1_v_inst.score_ctr[1] ),
    .A_N(\game1.scroll1_v_inst.score_ctr[0] ));
 sg13g2_or3_1 _2277_ (.A(\game1.scroll1_v_inst.score_ctr[5] ),
    .B(\game1.scroll1_v_inst.score_ctr[4] ),
    .C(\game1.scroll1_v_inst.score_ctr[3] ),
    .X(_0387_));
 sg13g2_nor4_2 _2278_ (.A(_0500_),
    .B(_0002_),
    .C(_0386_),
    .Y(_0388_),
    .D(_0387_));
 sg13g2_nand2_2 _2279_ (.Y(_0389_),
    .A(net2),
    .B(_0388_));
 sg13g2_inv_1 _2280_ (.Y(_0390_),
    .A(_0389_));
 sg13g2_nand2_1 _2281_ (.Y(_0391_),
    .A(net208),
    .B(net308));
 sg13g2_nor3_1 _2282_ (.A(net253),
    .B(net254),
    .C(\game1.score[2] ),
    .Y(_0392_));
 sg13g2_nand2_1 _2283_ (.Y(_0393_),
    .A(_0391_),
    .B(_0392_));
 sg13g2_a21oi_2 _2284_ (.B1(_0389_),
    .Y(_0394_),
    .A2(_0393_),
    .A1(_0195_));
 sg13g2_nor2b_1 _2285_ (.A(net186),
    .B_N(_0394_),
    .Y(_0395_));
 sg13g2_nor2_1 _2286_ (.A(net255),
    .B(_0394_),
    .Y(_0396_));
 sg13g2_nor3_1 _2287_ (.A(net227),
    .B(_0395_),
    .C(_0396_),
    .Y(_0114_));
 sg13g2_a21oi_1 _2288_ (.A1(\game1.score[0] ),
    .A2(_0394_),
    .Y(_0397_),
    .B1(net208));
 sg13g2_nor3_2 _2289_ (.A(_0195_),
    .B(_0389_),
    .C(_0391_),
    .Y(_0398_));
 sg13g2_nor3_1 _2290_ (.A(net226),
    .B(net209),
    .C(_0398_),
    .Y(_0115_));
 sg13g2_and4_1 _2291_ (.A(net292),
    .B(net208),
    .C(net255),
    .D(_0394_),
    .X(_0399_));
 sg13g2_nor2_1 _2292_ (.A(net292),
    .B(net309),
    .Y(_0400_));
 sg13g2_nor3_1 _2293_ (.A(net226),
    .B(_0399_),
    .C(_0400_),
    .Y(_0116_));
 sg13g2_and2_1 _2294_ (.A(_0562_),
    .B(_0398_),
    .X(_0401_));
 sg13g2_xnor2_1 _2295_ (.Y(_0402_),
    .A(net254),
    .B(_0401_));
 sg13g2_nor2_1 _2296_ (.A(net229),
    .B(net406),
    .Y(_0117_));
 sg13g2_and3_1 _2297_ (.X(_0403_),
    .A(net253),
    .B(net254),
    .C(_0399_));
 sg13g2_a21oi_1 _2298_ (.A1(net254),
    .A2(_0399_),
    .Y(_0404_),
    .B1(net253));
 sg13g2_nor3_1 _2299_ (.A(net226),
    .B(_0403_),
    .C(net396),
    .Y(_0118_));
 sg13g2_nand3_1 _2300_ (.B(_0561_),
    .C(_0399_),
    .A(net254),
    .Y(_0405_));
 sg13g2_xnor2_1 _2301_ (.Y(_0406_),
    .A(net252),
    .B(_0405_));
 sg13g2_nor2b_1 _2302_ (.A(net226),
    .B_N(net356),
    .Y(_0119_));
 sg13g2_a21oi_1 _2303_ (.A1(net252),
    .A2(_0403_),
    .Y(_0407_),
    .B1(net313));
 sg13g2_nor2_1 _2304_ (.A(net226),
    .B(net314),
    .Y(_0120_));
 sg13g2_and2_1 _2305_ (.A(net149),
    .B(_1069_),
    .X(_0121_));
 sg13g2_xnor2_1 _2306_ (.Y(_0408_),
    .A(\game1.scroll1_h_inst.ctr[1] ),
    .B(net211));
 sg13g2_nor2_1 _2307_ (.A(net212),
    .B(net280),
    .Y(_0122_));
 sg13g2_a21oi_1 _2308_ (.A1(\game1.scroll1_h_inst.ctr[1] ),
    .A2(\game1.scroll1_h_inst.ctr[0] ),
    .Y(_0409_),
    .B1(net160));
 sg13g2_nor3_1 _2309_ (.A(net212),
    .B(_1071_),
    .C(net161),
    .Y(_0123_));
 sg13g2_nor2_1 _2310_ (.A(net175),
    .B(_1071_),
    .Y(_0410_));
 sg13g2_nor3_1 _2311_ (.A(net212),
    .B(_1072_),
    .C(net176),
    .Y(_0124_));
 sg13g2_nor2_1 _2312_ (.A(net167),
    .B(_1072_),
    .Y(_0411_));
 sg13g2_nor3_1 _2313_ (.A(net212),
    .B(_1073_),
    .C(net168),
    .Y(_0125_));
 sg13g2_nor2_1 _2314_ (.A(net188),
    .B(_1073_),
    .Y(_0412_));
 sg13g2_nor3_1 _2315_ (.A(net212),
    .B(_1074_),
    .C(_0412_),
    .Y(_0126_));
 sg13g2_nor2_1 _2316_ (.A(net195),
    .B(_1074_),
    .Y(_0413_));
 sg13g2_nor3_1 _2317_ (.A(net212),
    .B(_1075_),
    .C(_0413_),
    .Y(_0127_));
 sg13g2_nor2_1 _2318_ (.A(net193),
    .B(_1075_),
    .Y(_0414_));
 sg13g2_nor3_1 _2319_ (.A(net212),
    .B(_1076_),
    .C(net194),
    .Y(_0128_));
 sg13g2_nor2_1 _2320_ (.A(net178),
    .B(_1076_),
    .Y(_0415_));
 sg13g2_nor3_1 _2321_ (.A(net212),
    .B(_1077_),
    .C(net179),
    .Y(_0129_));
 sg13g2_xor2_1 _2322_ (.B(_1096_),
    .A(net289),
    .X(_0416_));
 sg13g2_nor2_1 _2323_ (.A(net213),
    .B(net290),
    .Y(_0130_));
 sg13g2_nor3_2 _2324_ (.A(net177),
    .B(_0501_),
    .C(_0983_),
    .Y(_0417_));
 sg13g2_nand2b_1 _2325_ (.Y(_0418_),
    .B(_0417_),
    .A_N(net202));
 sg13g2_nand2_1 _2326_ (.Y(_0419_),
    .A(_0501_),
    .B(net202));
 sg13g2_a21oi_1 _2327_ (.A1(_0418_),
    .A2(_0419_),
    .Y(_0132_),
    .B1(net228));
 sg13g2_and2_1 _2328_ (.A(net191),
    .B(\game1.scroll1_v_inst.ctr[0] ),
    .X(_0420_));
 sg13g2_nor2_1 _2329_ (.A(_0978_),
    .B(_0420_),
    .Y(_0421_));
 sg13g2_a22oi_1 _2330_ (.Y(_0422_),
    .B1(_0417_),
    .B2(_0421_),
    .A2(net191),
    .A1(_0501_));
 sg13g2_nor2_1 _2331_ (.A(net228),
    .B(net192),
    .Y(_0133_));
 sg13g2_and3_1 _2332_ (.X(_0423_),
    .A(net2),
    .B(net173),
    .C(_0420_));
 sg13g2_a21oi_1 _2333_ (.A1(net2),
    .A2(_0420_),
    .Y(_0424_),
    .B1(net173));
 sg13g2_nor3_1 _2334_ (.A(net218),
    .B(_0423_),
    .C(net174),
    .Y(_0134_));
 sg13g2_xnor2_1 _2335_ (.Y(_0425_),
    .A(net294),
    .B(_0423_));
 sg13g2_nor2_1 _2336_ (.A(net216),
    .B(_0425_),
    .Y(_0135_));
 sg13g2_and4_1 _2337_ (.A(\game1.scroll1_v_inst.ctr[4] ),
    .B(\game1.scroll1_v_inst.ctr[3] ),
    .C(\game1.scroll1_v_inst.ctr[2] ),
    .D(_0420_),
    .X(_0426_));
 sg13g2_and2_1 _2338_ (.A(net2),
    .B(_0426_),
    .X(_0427_));
 sg13g2_a21oi_1 _2339_ (.A1(\game1.scroll1_v_inst.ctr[3] ),
    .A2(_0423_),
    .Y(_0428_),
    .B1(net156));
 sg13g2_nor3_1 _2340_ (.A(net218),
    .B(_0427_),
    .C(net157),
    .Y(_0136_));
 sg13g2_xnor2_1 _2341_ (.Y(_0429_),
    .A(net297),
    .B(_0426_));
 sg13g2_a22oi_1 _2342_ (.Y(_0430_),
    .B1(_0417_),
    .B2(_0429_),
    .A2(\game1.scroll1_v_inst.ctr[5] ),
    .A1(_0501_));
 sg13g2_nor2_1 _2343_ (.A(net228),
    .B(net298),
    .Y(_0137_));
 sg13g2_and3_1 _2344_ (.X(_0431_),
    .A(net180),
    .B(\game1.scroll1_v_inst.ctr[5] ),
    .C(_0427_));
 sg13g2_a21oi_1 _2345_ (.A1(\game1.scroll1_v_inst.ctr[5] ),
    .A2(_0427_),
    .Y(_0432_),
    .B1(net180));
 sg13g2_nor3_1 _2346_ (.A(net218),
    .B(_0431_),
    .C(net181),
    .Y(_0138_));
 sg13g2_nand3_1 _2347_ (.B(\game1.scroll1_v_inst.ctr[5] ),
    .C(_0426_),
    .A(net180),
    .Y(_0433_));
 sg13g2_xor2_1 _2348_ (.B(_0433_),
    .A(net305),
    .X(_0434_));
 sg13g2_a22oi_1 _2349_ (.Y(_0435_),
    .B1(_0417_),
    .B2(net306),
    .A2(\game1.scroll1_v_inst.ctr[7] ),
    .A1(_0501_));
 sg13g2_nor2_1 _2350_ (.A(net228),
    .B(net307),
    .Y(_0139_));
 sg13g2_a21oi_1 _2351_ (.A1(\game1.scroll1_v_inst.ctr[7] ),
    .A2(_0431_),
    .Y(_0436_),
    .B1(net357));
 sg13g2_nand2_1 _2352_ (.Y(_0437_),
    .A(\game1.scroll1_v_inst.ctr[8] ),
    .B(\game1.scroll1_v_inst.ctr[7] ));
 sg13g2_nor2_1 _2353_ (.A(_0433_),
    .B(_0437_),
    .Y(_0438_));
 sg13g2_a21o_1 _2354_ (.A2(_0438_),
    .A1(net2),
    .B1(net358),
    .X(_0439_));
 sg13g2_nor2_1 _2355_ (.A(net217),
    .B(_0439_),
    .Y(_0140_));
 sg13g2_xnor2_1 _2356_ (.Y(_0440_),
    .A(_0003_),
    .B(_0438_));
 sg13g2_a22oi_1 _2357_ (.Y(_0441_),
    .B1(_0417_),
    .B2(_0440_),
    .A2(net284),
    .A1(_0501_));
 sg13g2_nor2_1 _2358_ (.A(net228),
    .B(net285),
    .Y(_0141_));
 sg13g2_nand4_1 _2359_ (.B(\game1.scroll1_v_inst.ctr[8] ),
    .C(\game1.scroll1_v_inst.ctr[7] ),
    .A(net284),
    .Y(_0442_),
    .D(_0431_));
 sg13g2_and4_1 _2360_ (.A(\game1.scroll1_v_inst.ctr[9] ),
    .B(\game1.scroll1_v_inst.ctr[8] ),
    .C(\game1.scroll1_v_inst.ctr[7] ),
    .D(_0431_),
    .X(_0443_));
 sg13g2_xor2_1 _2361_ (.B(_0442_),
    .A(net322),
    .X(_0444_));
 sg13g2_nor2_1 _2362_ (.A(net217),
    .B(net323),
    .Y(_0142_));
 sg13g2_a21oi_1 _2363_ (.A1(\game1.scroll1_v_inst.ctr[10] ),
    .A2(_0443_),
    .Y(_0445_),
    .B1(net170));
 sg13g2_and3_1 _2364_ (.X(_0446_),
    .A(net170),
    .B(\game1.scroll1_v_inst.ctr[10] ),
    .C(_0443_));
 sg13g2_nor3_1 _2365_ (.A(net217),
    .B(net171),
    .C(_0446_),
    .Y(_0143_));
 sg13g2_nor2_1 _2366_ (.A(net205),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_and2_1 _2367_ (.A(net205),
    .B(_0446_),
    .X(_0448_));
 sg13g2_nor3_1 _2368_ (.A(net217),
    .B(net206),
    .C(_0448_),
    .Y(_0144_));
 sg13g2_nor2_1 _2369_ (.A(net207),
    .B(_0448_),
    .Y(_0449_));
 sg13g2_and2_1 _2370_ (.A(net207),
    .B(_0448_),
    .X(_0450_));
 sg13g2_nor3_1 _2371_ (.A(net217),
    .B(_0449_),
    .C(_0450_),
    .Y(_0145_));
 sg13g2_nor2_1 _2372_ (.A(net199),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_and2_1 _2373_ (.A(net199),
    .B(_0450_),
    .X(_0452_));
 sg13g2_nor3_1 _2374_ (.A(net217),
    .B(net200),
    .C(_0452_),
    .Y(_0146_));
 sg13g2_nor2_1 _2375_ (.A(net196),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_and2_1 _2376_ (.A(net196),
    .B(_0452_),
    .X(_0454_));
 sg13g2_nor3_1 _2377_ (.A(net217),
    .B(net197),
    .C(_0454_),
    .Y(_0147_));
 sg13g2_xnor2_1 _2378_ (.Y(_0455_),
    .A(net189),
    .B(_0454_));
 sg13g2_nor2_1 _2379_ (.A(net217),
    .B(net190),
    .Y(_0148_));
 sg13g2_and3_1 _2380_ (.X(_0149_),
    .A(net177),
    .B(_0501_),
    .C(net221));
 sg13g2_a21o_1 _2381_ (.A2(_0985_),
    .A1(net291),
    .B1(_0390_),
    .X(_0456_));
 sg13g2_nor2_1 _2382_ (.A(net291),
    .B(_0985_),
    .Y(_0457_));
 sg13g2_nor3_1 _2383_ (.A(net229),
    .B(_0456_),
    .C(_0457_),
    .Y(_0150_));
 sg13g2_xnor2_1 _2384_ (.Y(_0458_),
    .A(net312),
    .B(_0456_));
 sg13g2_nor2_1 _2385_ (.A(net228),
    .B(_0458_),
    .Y(_0151_));
 sg13g2_nand3_1 _2386_ (.B(net291),
    .C(_0985_),
    .A(net312),
    .Y(_0459_));
 sg13g2_and2_1 _2387_ (.A(_0500_),
    .B(_0459_),
    .X(_0460_));
 sg13g2_nor2_1 _2388_ (.A(_0500_),
    .B(_0459_),
    .Y(_0461_));
 sg13g2_nor4_1 _2389_ (.A(net229),
    .B(_0390_),
    .C(_0460_),
    .D(_0461_),
    .Y(_0152_));
 sg13g2_and2_1 _2390_ (.A(net203),
    .B(_0461_),
    .X(_0462_));
 sg13g2_nor2_1 _2391_ (.A(net203),
    .B(_0461_),
    .Y(_0463_));
 sg13g2_nor3_1 _2392_ (.A(net229),
    .B(_0462_),
    .C(net204),
    .Y(_0153_));
 sg13g2_xnor2_1 _2393_ (.Y(_0464_),
    .A(net299),
    .B(_0462_));
 sg13g2_nor2_1 _2394_ (.A(net229),
    .B(_0464_),
    .Y(_0154_));
 sg13g2_a21oi_1 _2395_ (.A1(\game1.scroll1_v_inst.score_ctr[4] ),
    .A2(_0462_),
    .Y(_0465_),
    .B1(net153));
 sg13g2_and3_1 _2396_ (.X(_0466_),
    .A(\game1.scroll1_v_inst.score_ctr[5] ),
    .B(\game1.scroll1_v_inst.score_ctr[4] ),
    .C(\game1.scroll1_v_inst.score_ctr[3] ));
 sg13g2_nand4_1 _2397_ (.B(\game1.scroll1_v_inst.score_ctr[1] ),
    .C(\game1.scroll1_v_inst.score_ctr[0] ),
    .A(\game1.scroll1_v_inst.score_ctr[2] ),
    .Y(_0467_),
    .D(_0466_));
 sg13g2_nand2_1 _2398_ (.Y(_0468_),
    .A(net220),
    .B(_0467_));
 sg13g2_a21oi_1 _2399_ (.A1(net218),
    .A2(_0468_),
    .Y(_0155_),
    .B1(net154));
 sg13g2_xor2_1 _2400_ (.B(_0467_),
    .A(_0002_),
    .X(_0469_));
 sg13g2_nand3b_1 _2401_ (.B(_0469_),
    .C(net215),
    .Y(_0470_),
    .A_N(_0388_));
 sg13g2_nand2_1 _2402_ (.Y(_0471_),
    .A(net158),
    .B(_0389_));
 sg13g2_o21ai_1 _2403_ (.B1(_0470_),
    .Y(_0156_),
    .A1(net218),
    .A2(_0471_));
 sg13g2_nor2_1 _2404_ (.A(net238),
    .B(_0591_),
    .Y(_0472_));
 sg13g2_nand4_1 _2405_ (.B(_0578_),
    .C(_0306_),
    .A(\game1.pixel_y[9] ),
    .Y(_0473_),
    .D(_0472_));
 sg13g2_nand2_1 _2406_ (.Y(_0474_),
    .A(net1),
    .B(_0473_));
 sg13g2_or2_2 _2407_ (.X(_0475_),
    .B(_0474_),
    .A(_1021_));
 sg13g2_inv_1 _2408_ (.Y(_0476_),
    .A(_0475_));
 sg13g2_a22oi_1 _2409_ (.Y(_0477_),
    .B1(_0476_),
    .B2(net150),
    .A2(net233),
    .A1(\game1.pixel_y[0] ));
 sg13g2_inv_1 _2410_ (.Y(_0158_),
    .A(net151));
 sg13g2_nor3_1 _2411_ (.A(_0576_),
    .B(_0590_),
    .C(_0475_),
    .Y(_0478_));
 sg13g2_a21o_1 _2412_ (.A2(net233),
    .A1(net251),
    .B1(_0478_),
    .X(_0159_));
 sg13g2_nand2_1 _2413_ (.Y(_0479_),
    .A(_0576_),
    .B(_1023_));
 sg13g2_o21ai_1 _2414_ (.B1(net1),
    .Y(_0480_),
    .A1(_1021_),
    .A2(_0473_));
 sg13g2_xor2_1 _2415_ (.B(_0479_),
    .A(net248),
    .X(_0481_));
 sg13g2_nor2_1 _2416_ (.A(_0480_),
    .B(_0481_),
    .Y(_0160_));
 sg13g2_nand2_1 _2417_ (.Y(_0482_),
    .A(net247),
    .B(net233));
 sg13g2_nor2b_1 _2418_ (.A(_0032_),
    .B_N(_0576_),
    .Y(_0483_));
 sg13g2_xnor2_1 _2419_ (.Y(_0484_),
    .A(net247),
    .B(_0483_));
 sg13g2_o21ai_1 _2420_ (.B1(_0482_),
    .Y(_0161_),
    .A1(_0475_),
    .A2(_0484_));
 sg13g2_nand2_1 _2421_ (.Y(_0485_),
    .A(net245),
    .B(net233));
 sg13g2_o21ai_1 _2422_ (.B1(_0485_),
    .Y(_0162_),
    .A1(_0298_),
    .A2(_0475_));
 sg13g2_nand2_1 _2423_ (.Y(_0486_),
    .A(net243),
    .B(net233));
 sg13g2_nor2_1 _2424_ (.A(_0031_),
    .B(_0296_),
    .Y(_0487_));
 sg13g2_xnor2_1 _2425_ (.Y(_0488_),
    .A(net243),
    .B(_0487_));
 sg13g2_o21ai_1 _2426_ (.B1(_0486_),
    .Y(_0163_),
    .A1(_0475_),
    .A2(_0488_));
 sg13g2_or2_1 _2427_ (.X(_0489_),
    .B(_0297_),
    .A(_0555_));
 sg13g2_nor2_1 _2428_ (.A(net233),
    .B(_0489_),
    .Y(_0490_));
 sg13g2_xnor2_1 _2429_ (.Y(_0491_),
    .A(net241),
    .B(_0490_));
 sg13g2_nor2_1 _2430_ (.A(_0480_),
    .B(_0491_),
    .Y(_0164_));
 sg13g2_nand2_1 _2431_ (.Y(_0492_),
    .A(net239),
    .B(net232));
 sg13g2_nor2_1 _2432_ (.A(_0029_),
    .B(_0489_),
    .Y(_0493_));
 sg13g2_xnor2_1 _2433_ (.Y(_0494_),
    .A(net239),
    .B(_0493_));
 sg13g2_o21ai_1 _2434_ (.B1(_0492_),
    .Y(_0165_),
    .A1(_0475_),
    .A2(_0494_));
 sg13g2_nor3_1 _2435_ (.A(_0573_),
    .B(net232),
    .C(_0489_),
    .Y(_0495_));
 sg13g2_xnor2_1 _2436_ (.Y(_0496_),
    .A(net238),
    .B(_0495_));
 sg13g2_nor2_1 _2437_ (.A(_0480_),
    .B(_0496_),
    .Y(_0166_));
 sg13g2_nor3_1 _2438_ (.A(_0025_),
    .B(_0573_),
    .C(_0489_),
    .Y(_0497_));
 sg13g2_o21ai_1 _2439_ (.B1(_0476_),
    .Y(_0498_),
    .A1(net237),
    .A2(_0497_));
 sg13g2_a21o_1 _2440_ (.A2(_0497_),
    .A1(net237),
    .B1(_0498_),
    .X(_0499_));
 sg13g2_o21ai_1 _2441_ (.B1(_0499_),
    .Y(_0167_),
    .A1(_0557_),
    .A2(_1023_));
 sg13g2_dfrbp_1 _2442_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net135),
    .D(_0041_),
    .Q_N(_1218_),
    .Q(\game1.obstacle3_y[1] ));
 sg13g2_dfrbp_1 _2443_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net142),
    .D(_0042_),
    .Q_N(_1217_),
    .Q(\game1.obstacle3_y[2] ));
 sg13g2_dfrbp_1 _2444_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net140),
    .D(_0043_),
    .Q_N(_1216_),
    .Q(\game1.obstacle3_y[3] ));
 sg13g2_dfrbp_1 _2445_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net138),
    .D(_0044_),
    .Q_N(_1215_),
    .Q(\game1.obstacle3_y[4] ));
 sg13g2_dfrbp_1 _2446_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net134),
    .D(_0045_),
    .Q_N(_0013_),
    .Q(\game1.obstacle3_y[5] ));
 sg13g2_dfrbp_1 _2447_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net132),
    .D(_0046_),
    .Q_N(_0012_),
    .Q(\game1.obstacle3_y[6] ));
 sg13g2_dfrbp_1 _2448_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net130),
    .D(_0047_),
    .Q_N(_0011_),
    .Q(\game1.obstacle3_y[7] ));
 sg13g2_dfrbp_1 _2449_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net128),
    .D(_0048_),
    .Q_N(_0015_),
    .Q(\game1.obstacle3_y[8] ));
 sg13g2_dfrbp_1 _2450_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net126),
    .D(_0049_),
    .Q_N(_0014_),
    .Q(\game1.obstacle3_y[9] ));
 sg13g2_dfrbp_1 _2451_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net124),
    .D(_0050_),
    .Q_N(_1214_),
    .Q(\game1.obstacle3_x[1] ));
 sg13g2_dfrbp_1 _2452_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net122),
    .D(net302),
    .Q_N(_1213_),
    .Q(\game1.obstacle3_x[2] ));
 sg13g2_dfrbp_1 _2453_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net120),
    .D(_0052_),
    .Q_N(_1212_),
    .Q(\game1.obstacle3_x[3] ));
 sg13g2_dfrbp_1 _2454_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net118),
    .D(_0053_),
    .Q_N(_1211_),
    .Q(\game1.obstacle3_x[4] ));
 sg13g2_dfrbp_1 _2455_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net116),
    .D(net403),
    .Q_N(_1210_),
    .Q(\game1.obstacle3_x[5] ));
 sg13g2_dfrbp_1 _2456_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net114),
    .D(_0055_),
    .Q_N(_1209_),
    .Q(\game1.obstacle3_x[6] ));
 sg13g2_dfrbp_1 _2457_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net112),
    .D(_0056_),
    .Q_N(_1208_),
    .Q(\game1.obstacle3_x[7] ));
 sg13g2_dfrbp_1 _2458_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net110),
    .D(_0057_),
    .Q_N(_1207_),
    .Q(\game1.obstacle3_x[8] ));
 sg13g2_dfrbp_1 _2459_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net108),
    .D(_0058_),
    .Q_N(_0016_),
    .Q(\game1.obstacle3_x[9] ));
 sg13g2_dfrbp_1 _2460_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net106),
    .D(net164),
    .Q_N(_1206_),
    .Q(\game1.obstacle1_y[1] ));
 sg13g2_dfrbp_1 _2461_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net104),
    .D(net365),
    .Q_N(_1205_),
    .Q(\game1.obstacle1_y[2] ));
 sg13g2_dfrbp_1 _2462_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net102),
    .D(net349),
    .Q_N(_1204_),
    .Q(\game1.obstacle1_y[3] ));
 sg13g2_dfrbp_1 _2463_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net100),
    .D(net288),
    .Q_N(_1203_),
    .Q(\game1.obstacle1_y[4] ));
 sg13g2_dfrbp_1 _2464_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net98),
    .D(net311),
    .Q_N(_0028_),
    .Q(\game1.obstacle1_y[5] ));
 sg13g2_dfrbp_1 _2465_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net96),
    .D(net373),
    .Q_N(_0027_),
    .Q(\game1.obstacle1_y[6] ));
 sg13g2_dfrbp_1 _2466_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net94),
    .D(net334),
    .Q_N(_1202_),
    .Q(\game1.obstacle1_y[7] ));
 sg13g2_dfrbp_1 _2467_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net92),
    .D(net318),
    .Q_N(_0026_),
    .Q(\game1.obstacle1_y[8] ));
 sg13g2_dfrbp_1 _2468_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net90),
    .D(_0067_),
    .Q_N(_0023_),
    .Q(\game1.obstacle1_y[9] ));
 sg13g2_dfrbp_1 _2469_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net88),
    .D(_0068_),
    .Q_N(_0040_),
    .Q(\game1.pixel_x[0] ));
 sg13g2_dfrbp_1 _2470_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net87),
    .D(_0069_),
    .Q_N(_1201_),
    .Q(\game1.pixel_x[1] ));
 sg13g2_dfrbp_1 _2471_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net86),
    .D(net351),
    .Q_N(_1200_),
    .Q(\game1.pixel_x[2] ));
 sg13g2_dfrbp_1 _2472_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net85),
    .D(_0071_),
    .Q_N(_1199_),
    .Q(\game1.pixel_x[3] ));
 sg13g2_dfrbp_1 _2473_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net84),
    .D(_0072_),
    .Q_N(_0022_),
    .Q(\game1.pixel_x[4] ));
 sg13g2_dfrbp_1 _2474_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net83),
    .D(_0073_),
    .Q_N(_0021_),
    .Q(\game1.pixel_x[5] ));
 sg13g2_dfrbp_1 _2475_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net82),
    .D(_0074_),
    .Q_N(_0020_),
    .Q(\game1.pixel_x[6] ));
 sg13g2_dfrbp_1 _2476_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net81),
    .D(_0075_),
    .Q_N(_1198_),
    .Q(\game1.pixel_x[7] ));
 sg13g2_dfrbp_1 _2477_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net80),
    .D(_0076_),
    .Q_N(_0019_),
    .Q(\game1.pixel_x[8] ));
 sg13g2_dfrbp_1 _2478_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net79),
    .D(net375),
    .Q_N(_0018_),
    .Q(\game1.pixel_x[9] ));
 sg13g2_dfrbp_1 _2479_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net78),
    .D(_0078_),
    .Q_N(_1197_),
    .Q(\game1.obstacle2_x[1] ));
 sg13g2_dfrbp_1 _2480_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net76),
    .D(net321),
    .Q_N(_1196_),
    .Q(\game1.obstacle2_x[2] ));
 sg13g2_dfrbp_1 _2481_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net74),
    .D(_0080_),
    .Q_N(_1195_),
    .Q(\game1.obstacle2_x[3] ));
 sg13g2_dfrbp_1 _2482_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net72),
    .D(net362),
    .Q_N(_1194_),
    .Q(\game1.obstacle2_x[4] ));
 sg13g2_dfrbp_1 _2483_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net70),
    .D(net367),
    .Q_N(_1193_),
    .Q(\game1.obstacle2_x[5] ));
 sg13g2_dfrbp_1 _2484_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net68),
    .D(_0083_),
    .Q_N(_1192_),
    .Q(\game1.obstacle2_x[6] ));
 sg13g2_dfrbp_1 _2485_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net66),
    .D(_0084_),
    .Q_N(_1191_),
    .Q(\game1.obstacle2_x[7] ));
 sg13g2_dfrbp_1 _2486_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net64),
    .D(_0085_),
    .Q_N(_1190_),
    .Q(\game1.obstacle2_x[8] ));
 sg13g2_dfrbp_1 _2487_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net62),
    .D(net328),
    .Q_N(_0033_),
    .Q(\game1.obstacle2_x[9] ));
 sg13g2_dfrbp_1 _2488_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net60),
    .D(_0087_),
    .Q_N(_1189_),
    .Q(\game1.scroll1_h_inst.ctr[9] ));
 sg13g2_dfrbp_1 _2489_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net59),
    .D(_0088_),
    .Q_N(_1188_),
    .Q(\game1.scroll1_h_inst.ctr[10] ));
 sg13g2_dfrbp_1 _2490_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net58),
    .D(net293),
    .Q_N(_1187_),
    .Q(\game1.scroll1_h_inst.ctr[11] ));
 sg13g2_dfrbp_1 _2491_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net57),
    .D(net342),
    .Q_N(_1186_),
    .Q(\game1.scroll1_h_inst.ctr[12] ));
 sg13g2_dfrbp_1 _2492_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net56),
    .D(net394),
    .Q_N(_1185_),
    .Q(\game1.scroll1_h_inst.ctr[13] ));
 sg13g2_dfrbp_1 _2493_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net55),
    .D(net390),
    .Q_N(_1184_),
    .Q(\game1.scroll1_h_inst.ctr[14] ));
 sg13g2_dfrbp_1 _2494_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net54),
    .D(_0093_),
    .Q_N(_1183_),
    .Q(\game1.scroll1_h_inst.ctr[15] ));
 sg13g2_dfrbp_1 _2495_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net53),
    .D(_0094_),
    .Q_N(_1182_),
    .Q(\game1.obstacle1_x[1] ));
 sg13g2_dfrbp_1 _2496_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net51),
    .D(_0095_),
    .Q_N(_1181_),
    .Q(\game1.obstacle1_x[2] ));
 sg13g2_dfrbp_1 _2497_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net49),
    .D(_0096_),
    .Q_N(_1180_),
    .Q(\game1.obstacle1_x[3] ));
 sg13g2_dfrbp_1 _2498_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net47),
    .D(_0097_),
    .Q_N(_1179_),
    .Q(\game1.obstacle1_x[4] ));
 sg13g2_dfrbp_1 _2499_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net45),
    .D(_0098_),
    .Q_N(_1178_),
    .Q(\game1.obstacle1_x[5] ));
 sg13g2_dfrbp_1 _2500_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net43),
    .D(_0099_),
    .Q_N(_1177_),
    .Q(\game1.obstacle1_x[6] ));
 sg13g2_dfrbp_1 _2501_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net41),
    .D(net422),
    .Q_N(_1176_),
    .Q(\game1.obstacle1_x[7] ));
 sg13g2_dfrbp_1 _2502_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net39),
    .D(_0101_),
    .Q_N(_1175_),
    .Q(\game1.obstacle1_x[8] ));
 sg13g2_dfrbp_1 _2503_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net37),
    .D(net184),
    .Q_N(_0017_),
    .Q(\game1.obstacle1_x[9] ));
 sg13g2_dfrbp_1 _2504_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net35),
    .D(net214),
    .Q_N(_1174_),
    .Q(\game1.move_h ));
 sg13g2_dfrbp_1 _2505_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net34),
    .D(net419),
    .Q_N(_1173_),
    .Q(\game1.obstacle2_y[1] ));
 sg13g2_dfrbp_1 _2506_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net32),
    .D(_0105_),
    .Q_N(_1172_),
    .Q(\game1.obstacle2_y[2] ));
 sg13g2_dfrbp_1 _2507_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net30),
    .D(_0106_),
    .Q_N(_1171_),
    .Q(\game1.obstacle2_y[3] ));
 sg13g2_dfrbp_1 _2508_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net28),
    .D(_0107_),
    .Q_N(_1170_),
    .Q(\game1.obstacle2_y[4] ));
 sg13g2_dfrbp_1 _2509_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net26),
    .D(_0108_),
    .Q_N(_0036_),
    .Q(\game1.obstacle2_y[5] ));
 sg13g2_dfrbp_1 _2510_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net24),
    .D(_0109_),
    .Q_N(_0035_),
    .Q(\game1.obstacle2_y[6] ));
 sg13g2_dfrbp_1 _2511_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net22),
    .D(_0110_),
    .Q_N(_1169_),
    .Q(\game1.obstacle2_y[7] ));
 sg13g2_dfrbp_1 _2512_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net20),
    .D(_0111_),
    .Q_N(_0034_),
    .Q(\game1.obstacle2_y[8] ));
 sg13g2_dfrbp_1 _2513_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net147),
    .D(net166),
    .Q_N(_1168_),
    .Q(\game1.obstacle2_y[9] ));
 sg13g2_dfrbp_1 _2514_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net145),
    .D(_0113_),
    .Q_N(_0010_),
    .Q(\game1.score_inst.o_score_rgb[0] ));
 sg13g2_dfrbp_1 _2515_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net144),
    .D(net187),
    .Q_N(_0039_),
    .Q(\game1.score[0] ));
 sg13g2_dfrbp_1 _2516_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net141),
    .D(net210),
    .Q_N(_0009_),
    .Q(\game1.score[1] ));
 sg13g2_dfrbp_1 _2517_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net137),
    .D(_0116_),
    .Q_N(_0008_),
    .Q(\game1.score[2] ));
 sg13g2_dfrbp_1 _2518_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net131),
    .D(_0117_),
    .Q_N(_1167_),
    .Q(\game1.score[3] ));
 sg13g2_dfrbp_1 _2519_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net127),
    .D(_0118_),
    .Q_N(_0007_),
    .Q(\game1.score[4] ));
 sg13g2_dfrbp_1 _2520_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net123),
    .D(_0119_),
    .Q_N(_0006_),
    .Q(\game1.score[5] ));
 sg13g2_dfrbp_1 _2521_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net119),
    .D(_0120_),
    .Q_N(_1166_),
    .Q(\game1.score[6] ));
 sg13g2_dfrbp_1 _2522_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net115),
    .D(_0121_),
    .Q_N(_0038_),
    .Q(\game1.scroll1_h_inst.ctr[0] ));
 sg13g2_dfrbp_1 _2523_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net113),
    .D(_0122_),
    .Q_N(_1165_),
    .Q(\game1.scroll1_h_inst.ctr[1] ));
 sg13g2_dfrbp_1 _2524_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net111),
    .D(net162),
    .Q_N(_1164_),
    .Q(\game1.scroll1_h_inst.ctr[2] ));
 sg13g2_dfrbp_1 _2525_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net109),
    .D(_0124_),
    .Q_N(_1163_),
    .Q(\game1.scroll1_h_inst.ctr[3] ));
 sg13g2_dfrbp_1 _2526_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net107),
    .D(net169),
    .Q_N(_1162_),
    .Q(\game1.scroll1_h_inst.ctr[4] ));
 sg13g2_dfrbp_1 _2527_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net105),
    .D(_0126_),
    .Q_N(_1161_),
    .Q(\game1.scroll1_h_inst.ctr[5] ));
 sg13g2_dfrbp_1 _2528_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net103),
    .D(_0127_),
    .Q_N(_1160_),
    .Q(\game1.scroll1_h_inst.ctr[6] ));
 sg13g2_dfrbp_1 _2529_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net101),
    .D(_0128_),
    .Q_N(_1159_),
    .Q(\game1.scroll1_h_inst.ctr[7] ));
 sg13g2_dfrbp_1 _2530_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net99),
    .D(_0129_),
    .Q_N(_1158_),
    .Q(\game1.scroll1_h_inst.ctr[8] ));
 sg13g2_dfrbp_1 _2531_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net97),
    .D(_0130_),
    .Q_N(_1157_),
    .Q(\game1.scroll1_h_inst.ctr[16] ));
 sg13g2_dfrbp_1 _2532_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net95),
    .D(net19),
    .Q_N(_1156_),
    .Q(\game1.scroll1_h_inst.ctr[17] ));
 sg13g2_dfrbp_1 _2533_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net93),
    .D(_0132_),
    .Q_N(_1155_),
    .Q(\game1.scroll1_v_inst.ctr[0] ));
 sg13g2_dfrbp_1 _2534_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net89),
    .D(_0133_),
    .Q_N(_1154_),
    .Q(\game1.scroll1_v_inst.ctr[1] ));
 sg13g2_dfrbp_1 _2535_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net75),
    .D(_0134_),
    .Q_N(_1153_),
    .Q(\game1.scroll1_v_inst.ctr[2] ));
 sg13g2_dfrbp_1 _2536_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net71),
    .D(_0135_),
    .Q_N(_1152_),
    .Q(\game1.scroll1_v_inst.ctr[3] ));
 sg13g2_dfrbp_1 _2537_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net67),
    .D(_0136_),
    .Q_N(_1151_),
    .Q(\game1.scroll1_v_inst.ctr[4] ));
 sg13g2_dfrbp_1 _2538_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net63),
    .D(_0137_),
    .Q_N(_0005_),
    .Q(\game1.scroll1_v_inst.ctr[5] ));
 sg13g2_dfrbp_1 _2539_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net52),
    .D(net182),
    .Q_N(_1150_),
    .Q(\game1.scroll1_v_inst.ctr[6] ));
 sg13g2_dfrbp_1 _2540_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net48),
    .D(_0139_),
    .Q_N(_0004_),
    .Q(\game1.scroll1_v_inst.ctr[7] ));
 sg13g2_dfrbp_1 _2541_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net44),
    .D(_0140_),
    .Q_N(_1149_),
    .Q(\game1.scroll1_v_inst.ctr[8] ));
 sg13g2_dfrbp_1 _2542_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net40),
    .D(_0141_),
    .Q_N(_0003_),
    .Q(\game1.scroll1_v_inst.ctr[9] ));
 sg13g2_dfrbp_1 _2543_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net36),
    .D(_0142_),
    .Q_N(_1148_),
    .Q(\game1.scroll1_v_inst.ctr[10] ));
 sg13g2_dfrbp_1 _2544_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net31),
    .D(net172),
    .Q_N(_1147_),
    .Q(\game1.scroll1_v_inst.ctr[11] ));
 sg13g2_dfrbp_1 _2545_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net27),
    .D(_0144_),
    .Q_N(_1146_),
    .Q(\game1.scroll1_v_inst.ctr[12] ));
 sg13g2_dfrbp_1 _2546_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net23),
    .D(_0145_),
    .Q_N(_1145_),
    .Q(\game1.scroll1_v_inst.ctr[13] ));
 sg13g2_dfrbp_1 _2547_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net148),
    .D(net201),
    .Q_N(_1144_),
    .Q(\game1.scroll1_v_inst.ctr[14] ));
 sg13g2_dfrbp_1 _2548_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net143),
    .D(net198),
    .Q_N(_1143_),
    .Q(\game1.scroll1_v_inst.ctr[15] ));
 sg13g2_dfrbp_1 _2549_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net133),
    .D(_0148_),
    .Q_N(_1142_),
    .Q(\game1.scroll1_v_inst.ctr[16] ));
 sg13g2_dfrbp_1 _2550_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net125),
    .D(_0149_),
    .Q_N(_1141_),
    .Q(\game1.scroll1_v_inst.ctr[17] ));
 sg13g2_dfrbp_1 _2551_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net117),
    .D(_0150_),
    .Q_N(_1140_),
    .Q(\game1.scroll1_v_inst.score_ctr[0] ));
 sg13g2_dfrbp_1 _2552_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net77),
    .D(_0151_),
    .Q_N(_1139_),
    .Q(\game1.scroll1_v_inst.score_ctr[1] ));
 sg13g2_dfrbp_1 _2553_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net69),
    .D(_0152_),
    .Q_N(_1138_),
    .Q(\game1.scroll1_v_inst.score_ctr[2] ));
 sg13g2_dfrbp_1 _2554_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net61),
    .D(_0153_),
    .Q_N(_1137_),
    .Q(\game1.scroll1_v_inst.score_ctr[3] ));
 sg13g2_dfrbp_1 _2555_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net46),
    .D(_0154_),
    .Q_N(_1136_),
    .Q(\game1.scroll1_v_inst.score_ctr[4] ));
 sg13g2_dfrbp_1 _2556_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net38),
    .D(net155),
    .Q_N(_1135_),
    .Q(\game1.scroll1_v_inst.score_ctr[5] ));
 sg13g2_dfrbp_1 _2557_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net136),
    .D(net159),
    .Q_N(_0002_),
    .Q(\game1.scroll1_v_inst.score_ctr[6] ));
 sg13g2_dfrbp_1 _2558_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net73),
    .D(_0000_),
    .Q_N(_1219_),
    .Q(\game1.hsync ));
 sg13g2_dfrbp_1 _2559_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net29),
    .D(net282),
    .Q_N(_1134_),
    .Q(\game1.vga_inst.vsync ));
 sg13g2_dfrbp_1 _2560_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net21),
    .D(net215),
    .Q_N(_1133_),
    .Q(\game1.move_v ));
 sg13g2_dfrbp_1 _2561_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net146),
    .D(_0158_),
    .Q_N(_0037_),
    .Q(\game1.pixel_y[0] ));
 sg13g2_dfrbp_1 _2562_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net129),
    .D(net408),
    .Q_N(_1132_),
    .Q(\game1.pixel_y[1] ));
 sg13g2_dfrbp_1 _2563_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net91),
    .D(_0160_),
    .Q_N(_0032_),
    .Q(\game1.pixel_y[2] ));
 sg13g2_dfrbp_1 _2564_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net65),
    .D(net383),
    .Q_N(_1131_),
    .Q(\game1.pixel_y[3] ));
 sg13g2_dfrbp_1 _2565_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net42),
    .D(_0162_),
    .Q_N(_0031_),
    .Q(\game1.pixel_y[4] ));
 sg13g2_dfrbp_1 _2566_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net25),
    .D(net381),
    .Q_N(_0030_),
    .Q(\game1.pixel_y[5] ));
 sg13g2_dfrbp_1 _2567_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net121),
    .D(_0164_),
    .Q_N(_0029_),
    .Q(\game1.pixel_y[6] ));
 sg13g2_dfrbp_1 _2568_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net50),
    .D(net410),
    .Q_N(_1130_),
    .Q(\game1.pixel_y[7] ));
 sg13g2_dfrbp_1 _2569_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net139),
    .D(_0166_),
    .Q_N(_0025_),
    .Q(\game1.pixel_y[8] ));
 sg13g2_dfrbp_1 _2570_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net33),
    .D(_0167_),
    .Q_N(_0024_),
    .Q(\game1.pixel_y[9] ));
 sg13g2_tiehi _2560__21 (.L_HI(net21));
 sg13g2_tiehi _2511__22 (.L_HI(net22));
 sg13g2_tiehi _2546__23 (.L_HI(net23));
 sg13g2_tiehi _2510__24 (.L_HI(net24));
 sg13g2_tiehi _2566__25 (.L_HI(net25));
 sg13g2_tiehi _2509__26 (.L_HI(net26));
 sg13g2_tiehi _2545__27 (.L_HI(net27));
 sg13g2_tiehi _2508__28 (.L_HI(net28));
 sg13g2_tiehi _2559__29 (.L_HI(net29));
 sg13g2_tiehi _2507__30 (.L_HI(net30));
 sg13g2_tiehi _2544__31 (.L_HI(net31));
 sg13g2_tiehi _2506__32 (.L_HI(net32));
 sg13g2_tiehi _2570__33 (.L_HI(net33));
 sg13g2_tiehi _2505__34 (.L_HI(net34));
 sg13g2_tiehi _2504__35 (.L_HI(net35));
 sg13g2_tiehi _2543__36 (.L_HI(net36));
 sg13g2_tiehi _2503__37 (.L_HI(net37));
 sg13g2_tiehi _2556__38 (.L_HI(net38));
 sg13g2_tiehi _2502__39 (.L_HI(net39));
 sg13g2_tiehi _2542__40 (.L_HI(net40));
 sg13g2_tiehi _2501__41 (.L_HI(net41));
 sg13g2_tiehi _2565__42 (.L_HI(net42));
 sg13g2_tiehi _2500__43 (.L_HI(net43));
 sg13g2_tiehi _2541__44 (.L_HI(net44));
 sg13g2_tiehi _2499__45 (.L_HI(net45));
 sg13g2_tiehi _2555__46 (.L_HI(net46));
 sg13g2_tiehi _2498__47 (.L_HI(net47));
 sg13g2_tiehi _2540__48 (.L_HI(net48));
 sg13g2_tiehi _2497__49 (.L_HI(net49));
 sg13g2_tiehi _2568__50 (.L_HI(net50));
 sg13g2_tiehi _2496__51 (.L_HI(net51));
 sg13g2_tiehi _2539__52 (.L_HI(net52));
 sg13g2_tiehi _2495__53 (.L_HI(net53));
 sg13g2_tiehi _2494__54 (.L_HI(net54));
 sg13g2_tiehi _2493__55 (.L_HI(net55));
 sg13g2_tiehi _2492__56 (.L_HI(net56));
 sg13g2_tiehi _2491__57 (.L_HI(net57));
 sg13g2_tiehi _2490__58 (.L_HI(net58));
 sg13g2_tiehi _2489__59 (.L_HI(net59));
 sg13g2_tiehi _2488__60 (.L_HI(net60));
 sg13g2_tiehi _2554__61 (.L_HI(net61));
 sg13g2_tiehi _2487__62 (.L_HI(net62));
 sg13g2_tiehi _2538__63 (.L_HI(net63));
 sg13g2_tiehi _2486__64 (.L_HI(net64));
 sg13g2_tiehi _2564__65 (.L_HI(net65));
 sg13g2_tiehi _2485__66 (.L_HI(net66));
 sg13g2_tiehi _2537__67 (.L_HI(net67));
 sg13g2_tiehi _2484__68 (.L_HI(net68));
 sg13g2_tiehi _2553__69 (.L_HI(net69));
 sg13g2_tiehi _2483__70 (.L_HI(net70));
 sg13g2_tiehi _2536__71 (.L_HI(net71));
 sg13g2_tiehi _2482__72 (.L_HI(net72));
 sg13g2_tiehi _2558__73 (.L_HI(net73));
 sg13g2_tiehi _2481__74 (.L_HI(net74));
 sg13g2_tiehi _2535__75 (.L_HI(net75));
 sg13g2_tiehi _2480__76 (.L_HI(net76));
 sg13g2_tiehi _2552__77 (.L_HI(net77));
 sg13g2_tiehi _2479__78 (.L_HI(net78));
 sg13g2_tiehi _2478__79 (.L_HI(net79));
 sg13g2_tiehi _2477__80 (.L_HI(net80));
 sg13g2_tiehi _2476__81 (.L_HI(net81));
 sg13g2_tiehi _2475__82 (.L_HI(net82));
 sg13g2_tiehi _2474__83 (.L_HI(net83));
 sg13g2_tiehi _2473__84 (.L_HI(net84));
 sg13g2_tiehi _2472__85 (.L_HI(net85));
 sg13g2_tiehi _2471__86 (.L_HI(net86));
 sg13g2_tiehi _2470__87 (.L_HI(net87));
 sg13g2_tiehi _2469__88 (.L_HI(net88));
 sg13g2_tiehi _2534__89 (.L_HI(net89));
 sg13g2_tiehi _2468__90 (.L_HI(net90));
 sg13g2_tiehi _2563__91 (.L_HI(net91));
 sg13g2_tiehi _2467__92 (.L_HI(net92));
 sg13g2_tiehi _2533__93 (.L_HI(net93));
 sg13g2_tiehi _2466__94 (.L_HI(net94));
 sg13g2_tiehi _2532__95 (.L_HI(net95));
 sg13g2_tiehi _2465__96 (.L_HI(net96));
 sg13g2_tiehi _2531__97 (.L_HI(net97));
 sg13g2_tiehi _2464__98 (.L_HI(net98));
 sg13g2_tiehi _2530__99 (.L_HI(net99));
 sg13g2_tiehi _2463__100 (.L_HI(net100));
 sg13g2_tiehi _2529__101 (.L_HI(net101));
 sg13g2_tiehi _2462__102 (.L_HI(net102));
 sg13g2_tiehi _2528__103 (.L_HI(net103));
 sg13g2_tiehi _2461__104 (.L_HI(net104));
 sg13g2_tiehi _2527__105 (.L_HI(net105));
 sg13g2_tiehi _2460__106 (.L_HI(net106));
 sg13g2_tiehi _2526__107 (.L_HI(net107));
 sg13g2_tiehi _2459__108 (.L_HI(net108));
 sg13g2_tiehi _2525__109 (.L_HI(net109));
 sg13g2_tiehi _2458__110 (.L_HI(net110));
 sg13g2_tiehi _2524__111 (.L_HI(net111));
 sg13g2_tiehi _2457__112 (.L_HI(net112));
 sg13g2_tiehi _2523__113 (.L_HI(net113));
 sg13g2_tiehi _2456__114 (.L_HI(net114));
 sg13g2_tiehi _2522__115 (.L_HI(net115));
 sg13g2_tiehi _2455__116 (.L_HI(net116));
 sg13g2_tiehi _2551__117 (.L_HI(net117));
 sg13g2_tiehi _2454__118 (.L_HI(net118));
 sg13g2_tiehi _2521__119 (.L_HI(net119));
 sg13g2_tiehi _2453__120 (.L_HI(net120));
 sg13g2_tiehi _2567__121 (.L_HI(net121));
 sg13g2_tiehi _2452__122 (.L_HI(net122));
 sg13g2_tiehi _2520__123 (.L_HI(net123));
 sg13g2_tiehi _2451__124 (.L_HI(net124));
 sg13g2_tiehi _2550__125 (.L_HI(net125));
 sg13g2_tiehi _2450__126 (.L_HI(net126));
 sg13g2_tiehi _2519__127 (.L_HI(net127));
 sg13g2_tiehi _2449__128 (.L_HI(net128));
 sg13g2_tiehi _2562__129 (.L_HI(net129));
 sg13g2_tiehi _2448__130 (.L_HI(net130));
 sg13g2_tiehi _2518__131 (.L_HI(net131));
 sg13g2_tiehi _2447__132 (.L_HI(net132));
 sg13g2_tiehi _2549__133 (.L_HI(net133));
 sg13g2_tiehi _2446__134 (.L_HI(net134));
 sg13g2_tiehi _2442__135 (.L_HI(net135));
 sg13g2_tiehi _2557__136 (.L_HI(net136));
 sg13g2_tiehi _2517__137 (.L_HI(net137));
 sg13g2_tiehi _2445__138 (.L_HI(net138));
 sg13g2_tiehi _2569__139 (.L_HI(net139));
 sg13g2_tiehi _2444__140 (.L_HI(net140));
 sg13g2_tiehi _2516__141 (.L_HI(net141));
 sg13g2_tiehi _2443__142 (.L_HI(net142));
 sg13g2_tiehi _2548__143 (.L_HI(net143));
 sg13g2_tiehi _2515__144 (.L_HI(net144));
 sg13g2_tiehi _2514__145 (.L_HI(net145));
 sg13g2_tiehi _2561__146 (.L_HI(net146));
 sg13g2_tiehi _2513__147 (.L_HI(net147));
 sg13g2_tiehi _2547__148 (.L_HI(net148));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_10_vga_crossyroad_4 (.L_LO(net4));
 sg13g2_tielo tt_um_10_vga_crossyroad_5 (.L_LO(net5));
 sg13g2_tielo tt_um_10_vga_crossyroad_6 (.L_LO(net6));
 sg13g2_tielo tt_um_10_vga_crossyroad_7 (.L_LO(net7));
 sg13g2_tielo tt_um_10_vga_crossyroad_8 (.L_LO(net8));
 sg13g2_tielo tt_um_10_vga_crossyroad_9 (.L_LO(net9));
 sg13g2_tielo tt_um_10_vga_crossyroad_10 (.L_LO(net10));
 sg13g2_tielo tt_um_10_vga_crossyroad_11 (.L_LO(net11));
 sg13g2_tielo tt_um_10_vga_crossyroad_12 (.L_LO(net12));
 sg13g2_tielo tt_um_10_vga_crossyroad_13 (.L_LO(net13));
 sg13g2_tielo tt_um_10_vga_crossyroad_14 (.L_LO(net14));
 sg13g2_tielo tt_um_10_vga_crossyroad_15 (.L_LO(net15));
 sg13g2_tielo tt_um_10_vga_crossyroad_16 (.L_LO(net16));
 sg13g2_tielo tt_um_10_vga_crossyroad_17 (.L_LO(net17));
 sg13g2_tielo tt_um_10_vga_crossyroad_18 (.L_LO(net18));
 sg13g2_tielo _2532__19 (.L_LO(net19));
 sg13g2_tiehi _2512__20 (.L_HI(net20));
 sg13g2_buf_1 _2717_ (.A(uo_out[4]),
    .X(uo_out[0]));
 sg13g2_buf_1 _2718_ (.A(uo_out[5]),
    .X(uo_out[1]));
 sg13g2_buf_1 _2719_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_1 _2720_ (.A(\game1.vga_inst.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2721_ (.A(\game1.hsync ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout212 (.A(_1070_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_1070_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_0103_),
    .X(net214));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(_0157_));
 sg13g2_buf_2 fanout216 (.A(net219),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(net218),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(net219),
    .X(net218));
 sg13g2_buf_1 fanout219 (.A(_0986_),
    .X(net219));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(_0919_));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(_0919_));
 sg13g2_buf_2 fanout222 (.A(net223),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(net230),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(net225),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(net230),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(net227),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(net230),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(net229),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(net230),
    .X(net229));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(_0918_));
 sg13g2_buf_2 fanout231 (.A(_1067_),
    .X(net231));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(_1022_));
 sg13g2_buf_2 fanout233 (.A(_1022_),
    .X(net233));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(_0547_));
 sg13g2_buf_2 fanout235 (.A(_0506_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_0506_),
    .X(net236));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(\game1.pixel_y[9] ));
 sg13g2_buf_4 fanout238 (.X(net238),
    .A(net281));
 sg13g2_buf_2 fanout239 (.A(net409),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(net409),
    .X(net240));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(net397));
 sg13g2_buf_1 fanout242 (.A(net397),
    .X(net242));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(net380));
 sg13g2_buf_1 fanout244 (.A(\game1.pixel_y[5] ),
    .X(net244));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(net401));
 sg13g2_buf_2 fanout246 (.A(net247),
    .X(net246));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(net382));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(net249));
 sg13g2_buf_2 fanout249 (.A(\game1.pixel_y[2] ),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(\game1.pixel_y[1] ),
    .X(net250));
 sg13g2_buf_1 fanout251 (.A(net407),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(\game1.score[5] ),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(net395),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(\game1.score[3] ),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(net308),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(net418),
    .X(net256));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(\game1.move_h ));
 sg13g2_buf_2 fanout258 (.A(net434),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(net421),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(\game1.obstacle2_x[7] ),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(net374));
 sg13g2_buf_2 fanout262 (.A(\game1.pixel_x[9] ),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(net428));
 sg13g2_buf_2 fanout264 (.A(net392),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(net392),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(net267),
    .X(net266));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(\game1.pixel_x[6] ));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(net384));
 sg13g2_buf_2 fanout269 (.A(\game1.pixel_x[5] ),
    .X(net269));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(_0022_));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(net416));
 sg13g2_buf_1 fanout272 (.A(\game1.pixel_x[4] ),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(\game1.pixel_x[3] ),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(\game1.pixel_x[3] ),
    .X(net275));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(\game1.pixel_x[2] ));
 sg13g2_buf_2 fanout277 (.A(\game1.obstacle1_y[1] ),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(net429),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(net411),
    .X(net279));
 sg13g2_buf_4 input1 (.X(net1),
    .A(rst_n));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_tielo tt_um_10_vga_crossyroad_3 (.L_LO(net3));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0038_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0037_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0477_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0040_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold5 (.A(\game1.scroll1_v_inst.score_ctr[5] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0465_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0155_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold8 (.A(\game1.scroll1_v_inst.ctr[4] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0428_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold10 (.A(\game1.scroll1_v_inst.score_ctr[6] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0156_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold12 (.A(\game1.scroll1_h_inst.ctr[2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0409_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0123_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold15 (.A(\game1.obstacle1_y[1] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0059_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold17 (.A(\game1.move_v ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0112_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold19 (.A(\game1.scroll1_h_inst.ctr[4] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0411_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0125_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold22 (.A(\game1.scroll1_v_inst.ctr[11] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0445_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0143_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold25 (.A(\game1.scroll1_v_inst.ctr[2] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0424_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold27 (.A(\game1.scroll1_h_inst.ctr[3] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0410_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold29 (.A(\game1.scroll1_v_inst.ctr[17] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold30 (.A(\game1.scroll1_h_inst.ctr[8] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0415_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold32 (.A(\game1.scroll1_v_inst.ctr[6] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0432_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0138_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold35 (.A(\game1.obstacle1_x[9] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0102_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold37 (.A(\game1.obstacle3_y[9] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0039_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0114_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold40 (.A(\game1.scroll1_h_inst.ctr[5] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold41 (.A(\game1.scroll1_v_inst.ctr[16] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0455_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold43 (.A(\game1.scroll1_v_inst.ctr[1] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0422_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold45 (.A(\game1.scroll1_h_inst.ctr[7] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0414_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold47 (.A(\game1.scroll1_h_inst.ctr[6] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold48 (.A(\game1.scroll1_v_inst.ctr[15] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0453_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0147_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold51 (.A(\game1.scroll1_v_inst.ctr[14] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0451_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0146_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold54 (.A(\game1.scroll1_v_inst.ctr[0] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold55 (.A(\game1.scroll1_v_inst.score_ctr[3] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0463_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold57 (.A(\game1.scroll1_v_inst.ctr[12] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0447_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold59 (.A(\game1.scroll1_v_inst.ctr[13] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold60 (.A(\game1.score[1] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0397_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0115_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold63 (.A(\game1.scroll1_h_inst.ctr[0] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0408_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold65 (.A(\game1.pixel_y[8] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0001_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold67 (.A(\game1.obstacle1_x[1] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold68 (.A(\game1.scroll1_v_inst.ctr[9] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0441_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold70 (.A(\game1.obstacle1_y[9] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold71 (.A(\game1.obstacle1_y[4] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0062_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold73 (.A(\game1.scroll1_h_inst.ctr[16] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0416_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold75 (.A(\game1.scroll1_v_inst.score_ctr[0] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold76 (.A(\game1.score[2] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0089_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold78 (.A(\game1.scroll1_v_inst.ctr[3] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold79 (.A(\game1.scroll1_h_inst.ctr[10] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold80 (.A(_1080_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0005_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0430_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold83 (.A(\game1.scroll1_v_inst.score_ctr[4] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold84 (.A(\game1.obstacle3_x[2] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0949_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0051_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold87 (.A(\game1.obstacle2_y[8] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0194_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0004_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0434_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0435_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold92 (.A(\game1.score[0] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0398_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold94 (.A(\game1.obstacle1_y[5] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0063_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold96 (.A(\game1.scroll1_v_inst.score_ctr[1] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold97 (.A(\game1.score[6] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0407_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold99 (.A(\game1.obstacle3_y[5] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0943_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold101 (.A(\game1.obstacle1_y[8] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0066_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold103 (.A(\game1.obstacle2_x[2] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold104 (.A(_1038_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0079_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold106 (.A(\game1.scroll1_v_inst.ctr[10] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0444_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold108 (.A(\game1.obstacle3_y[7] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0946_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold110 (.A(\game1.obstacle2_x[9] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold111 (.A(_1058_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0086_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold113 (.A(\game1.obstacle3_y[8] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0947_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold115 (.A(\game1.obstacle3_x[1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0948_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold117 (.A(\game1.obstacle1_y[7] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0065_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold119 (.A(\game1.obstacle2_y[5] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0189_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold121 (.A(\game1.obstacle2_y[4] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0188_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold123 (.A(\game1.scroll1_h_inst.ctr[9] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold124 (.A(\game1.scroll1_h_inst.ctr[12] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold125 (.A(_1087_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0090_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0035_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0190_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0191_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold130 (.A(\game1.obstacle3_y[3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0940_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold132 (.A(\game1.obstacle1_y[3] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0061_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold134 (.A(\game1.pixel_x[0] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0070_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold136 (.A(\game1.obstacle2_y[3] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0186_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold138 (.A(\game1.obstacle3_y[4] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0007_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0406_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold141 (.A(\game1.scroll1_v_inst.ctr[8] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0436_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold143 (.A(\game1.obstacle2_x[1] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold144 (.A(_1037_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold145 (.A(\game1.obstacle2_x[4] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0081_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold147 (.A(\game1.pixel_x[2] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold148 (.A(\game1.obstacle1_y[2] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0060_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold150 (.A(\game1.obstacle2_x[5] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0082_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0012_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0945_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0027_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold155 (.A(_1010_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold156 (.A(_1011_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0064_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold158 (.A(\game1.pixel_x[9] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0077_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold160 (.A(\game1.obstacle2_y[7] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0192_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold162 (.A(\game1.obstacle2_y[2] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0183_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold164 (.A(\game1.pixel_y[5] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0163_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold166 (.A(\game1.pixel_y[3] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0161_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold168 (.A(\game1.pixel_x[5] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0016_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0972_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold171 (.A(\game1.scroll1_v_inst.score_ctr[2] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold172 (.A(\game1.scroll1_h_inst.ctr[14] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold173 (.A(_1094_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0092_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold175 (.A(\game1.obstacle2_x[8] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold176 (.A(\game1.pixel_x[7] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold177 (.A(\game1.scroll1_h_inst.ctr[13] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0091_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold179 (.A(\game1.score[4] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0404_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold181 (.A(\game1.pixel_y[6] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold182 (.A(\game1.obstacle3_x[4] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold183 (.A(\game1.obstacle3_y[2] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold184 (.A(\game1.scroll1_h_inst.ctr[15] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold185 (.A(\game1.pixel_y[4] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold186 (.A(\game1.obstacle3_x[5] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0054_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold188 (.A(\game1.obstacle3_x[8] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0008_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0402_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold191 (.A(\game1.pixel_y[1] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0159_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold193 (.A(\game1.pixel_y[7] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0165_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold195 (.A(\game1.obstacle3_y[1] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold196 (.A(\game1.obstacle3_x[7] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0967_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold198 (.A(\game1.obstacle1_x[5] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold199 (.A(\game1.obstacle2_x[6] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold200 (.A(\game1.pixel_x[4] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold201 (.A(\game1.pixel_x[1] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold202 (.A(\game1.obstacle2_y[1] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0104_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0022_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold205 (.A(\game1.obstacle1_x[7] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0100_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0018_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold208 (.A(\game1.obstacle1_x[2] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold209 (.A(\game1.obstacle1_x[6] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold210 (.A(\game1.obstacle3_x[6] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0957_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold212 (.A(\game1.pixel_x[8] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold213 (.A(\game1.obstacle3_x[3] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold214 (.A(\game1.obstacle1_x[3] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold215 (.A(\game1.obstacle1_x[4] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold216 (.A(\game1.obstacle1_x[8] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold217 (.A(\game1.scroll1_h_inst.ctr[17] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold218 (.A(\game1.move_h ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold219 (.A(_1055_),
    .X(net435));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_4 FILLER_0_329 ();
 sg13g2_fill_1 FILLER_0_333 ();
 sg13g2_decap_4 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_4 FILLER_1_301 ();
 sg13g2_fill_2 FILLER_1_305 ();
 sg13g2_fill_2 FILLER_1_311 ();
 sg13g2_fill_1 FILLER_1_313 ();
 sg13g2_fill_2 FILLER_1_332 ();
 sg13g2_fill_2 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_fill_2 FILLER_2_294 ();
 sg13g2_fill_1 FILLER_2_329 ();
 sg13g2_fill_1 FILLER_2_356 ();
 sg13g2_fill_2 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_137 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_4 FILLER_3_207 ();
 sg13g2_fill_1 FILLER_3_211 ();
 sg13g2_decap_4 FILLER_3_238 ();
 sg13g2_fill_1 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_247 ();
 sg13g2_decap_8 FILLER_3_267 ();
 sg13g2_fill_2 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_276 ();
 sg13g2_fill_2 FILLER_3_303 ();
 sg13g2_fill_1 FILLER_3_305 ();
 sg13g2_fill_1 FILLER_3_338 ();
 sg13g2_fill_2 FILLER_3_357 ();
 sg13g2_fill_1 FILLER_3_359 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_4 FILLER_4_49 ();
 sg13g2_fill_1 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_80 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_fill_2 FILLER_4_109 ();
 sg13g2_fill_1 FILLER_4_111 ();
 sg13g2_decap_8 FILLER_4_115 ();
 sg13g2_decap_8 FILLER_4_122 ();
 sg13g2_decap_8 FILLER_4_129 ();
 sg13g2_decap_8 FILLER_4_136 ();
 sg13g2_decap_8 FILLER_4_143 ();
 sg13g2_decap_8 FILLER_4_150 ();
 sg13g2_decap_8 FILLER_4_157 ();
 sg13g2_decap_8 FILLER_4_164 ();
 sg13g2_decap_8 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_178 ();
 sg13g2_fill_2 FILLER_4_185 ();
 sg13g2_decap_8 FILLER_4_213 ();
 sg13g2_fill_2 FILLER_4_246 ();
 sg13g2_decap_4 FILLER_4_283 ();
 sg13g2_fill_1 FILLER_4_287 ();
 sg13g2_fill_2 FILLER_4_318 ();
 sg13g2_fill_1 FILLER_4_320 ();
 sg13g2_fill_2 FILLER_4_367 ();
 sg13g2_fill_1 FILLER_4_369 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_4 FILLER_5_14 ();
 sg13g2_fill_1 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_27 ();
 sg13g2_decap_4 FILLER_5_42 ();
 sg13g2_fill_1 FILLER_5_46 ();
 sg13g2_fill_2 FILLER_5_122 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_fill_1 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_145 ();
 sg13g2_decap_8 FILLER_5_152 ();
 sg13g2_decap_8 FILLER_5_159 ();
 sg13g2_decap_8 FILLER_5_166 ();
 sg13g2_decap_8 FILLER_5_173 ();
 sg13g2_decap_8 FILLER_5_180 ();
 sg13g2_decap_8 FILLER_5_187 ();
 sg13g2_decap_8 FILLER_5_194 ();
 sg13g2_fill_2 FILLER_5_201 ();
 sg13g2_fill_1 FILLER_5_253 ();
 sg13g2_fill_2 FILLER_5_290 ();
 sg13g2_fill_2 FILLER_5_310 ();
 sg13g2_fill_2 FILLER_5_361 ();
 sg13g2_fill_1 FILLER_5_363 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_33 ();
 sg13g2_fill_2 FILLER_6_93 ();
 sg13g2_fill_1 FILLER_6_102 ();
 sg13g2_decap_8 FILLER_6_156 ();
 sg13g2_decap_8 FILLER_6_163 ();
 sg13g2_decap_8 FILLER_6_170 ();
 sg13g2_decap_8 FILLER_6_177 ();
 sg13g2_decap_8 FILLER_6_184 ();
 sg13g2_fill_2 FILLER_6_191 ();
 sg13g2_fill_1 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_207 ();
 sg13g2_fill_2 FILLER_6_218 ();
 sg13g2_fill_2 FILLER_6_229 ();
 sg13g2_fill_1 FILLER_6_231 ();
 sg13g2_fill_2 FILLER_6_247 ();
 sg13g2_fill_1 FILLER_6_254 ();
 sg13g2_decap_4 FILLER_6_283 ();
 sg13g2_fill_1 FILLER_6_366 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_72 ();
 sg13g2_fill_1 FILLER_7_103 ();
 sg13g2_fill_2 FILLER_7_112 ();
 sg13g2_decap_4 FILLER_7_127 ();
 sg13g2_fill_2 FILLER_7_152 ();
 sg13g2_fill_1 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_fill_1 FILLER_7_168 ();
 sg13g2_fill_1 FILLER_7_189 ();
 sg13g2_decap_4 FILLER_7_213 ();
 sg13g2_fill_1 FILLER_7_217 ();
 sg13g2_fill_2 FILLER_7_223 ();
 sg13g2_decap_8 FILLER_7_237 ();
 sg13g2_fill_1 FILLER_7_244 ();
 sg13g2_decap_4 FILLER_7_260 ();
 sg13g2_fill_1 FILLER_7_264 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_9 ();
 sg13g2_decap_4 FILLER_8_115 ();
 sg13g2_decap_4 FILLER_8_124 ();
 sg13g2_fill_2 FILLER_8_133 ();
 sg13g2_fill_1 FILLER_8_151 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_fill_1 FILLER_8_193 ();
 sg13g2_fill_1 FILLER_8_208 ();
 sg13g2_fill_1 FILLER_8_232 ();
 sg13g2_fill_2 FILLER_8_239 ();
 sg13g2_fill_1 FILLER_8_309 ();
 sg13g2_fill_1 FILLER_8_329 ();
 sg13g2_fill_1 FILLER_8_334 ();
 sg13g2_fill_1 FILLER_8_360 ();
 sg13g2_fill_2 FILLER_9_26 ();
 sg13g2_decap_4 FILLER_9_109 ();
 sg13g2_fill_2 FILLER_9_113 ();
 sg13g2_decap_8 FILLER_9_145 ();
 sg13g2_decap_8 FILLER_9_152 ();
 sg13g2_fill_2 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_176 ();
 sg13g2_decap_4 FILLER_9_183 ();
 sg13g2_decap_4 FILLER_9_192 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_fill_2 FILLER_9_217 ();
 sg13g2_fill_1 FILLER_9_219 ();
 sg13g2_decap_8 FILLER_9_237 ();
 sg13g2_decap_8 FILLER_9_244 ();
 sg13g2_fill_2 FILLER_9_267 ();
 sg13g2_fill_1 FILLER_9_269 ();
 sg13g2_fill_1 FILLER_9_284 ();
 sg13g2_fill_2 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_11 ();
 sg13g2_fill_2 FILLER_10_20 ();
 sg13g2_fill_1 FILLER_10_26 ();
 sg13g2_fill_1 FILLER_10_48 ();
 sg13g2_fill_2 FILLER_10_62 ();
 sg13g2_fill_2 FILLER_10_76 ();
 sg13g2_fill_2 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_116 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_decap_4 FILLER_10_131 ();
 sg13g2_fill_2 FILLER_10_135 ();
 sg13g2_fill_1 FILLER_10_146 ();
 sg13g2_decap_4 FILLER_10_151 ();
 sg13g2_fill_1 FILLER_10_165 ();
 sg13g2_fill_2 FILLER_10_218 ();
 sg13g2_fill_1 FILLER_10_220 ();
 sg13g2_decap_8 FILLER_10_239 ();
 sg13g2_decap_4 FILLER_10_246 ();
 sg13g2_fill_1 FILLER_10_250 ();
 sg13g2_fill_2 FILLER_10_272 ();
 sg13g2_fill_1 FILLER_10_287 ();
 sg13g2_fill_2 FILLER_10_307 ();
 sg13g2_fill_1 FILLER_10_309 ();
 sg13g2_fill_2 FILLER_10_317 ();
 sg13g2_fill_2 FILLER_10_326 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_50 ();
 sg13g2_fill_2 FILLER_11_60 ();
 sg13g2_fill_1 FILLER_11_93 ();
 sg13g2_fill_1 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_114 ();
 sg13g2_fill_2 FILLER_11_129 ();
 sg13g2_decap_8 FILLER_11_181 ();
 sg13g2_decap_4 FILLER_11_198 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_fill_2 FILLER_11_218 ();
 sg13g2_fill_1 FILLER_11_220 ();
 sg13g2_fill_2 FILLER_11_248 ();
 sg13g2_fill_1 FILLER_11_250 ();
 sg13g2_fill_2 FILLER_11_282 ();
 sg13g2_fill_2 FILLER_11_341 ();
 sg13g2_fill_1 FILLER_11_378 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_83 ();
 sg13g2_fill_2 FILLER_12_90 ();
 sg13g2_fill_2 FILLER_12_124 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_132 ();
 sg13g2_fill_2 FILLER_12_137 ();
 sg13g2_decap_4 FILLER_12_143 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_fill_2 FILLER_12_162 ();
 sg13g2_fill_1 FILLER_12_164 ();
 sg13g2_fill_1 FILLER_12_218 ();
 sg13g2_fill_1 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_244 ();
 sg13g2_decap_4 FILLER_12_254 ();
 sg13g2_fill_2 FILLER_12_263 ();
 sg13g2_fill_1 FILLER_12_274 ();
 sg13g2_fill_2 FILLER_12_294 ();
 sg13g2_fill_2 FILLER_12_305 ();
 sg13g2_fill_1 FILLER_12_307 ();
 sg13g2_fill_2 FILLER_12_321 ();
 sg13g2_fill_1 FILLER_12_327 ();
 sg13g2_fill_1 FILLER_12_337 ();
 sg13g2_fill_1 FILLER_12_346 ();
 sg13g2_fill_1 FILLER_12_361 ();
 sg13g2_fill_2 FILLER_12_391 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_4 ();
 sg13g2_fill_1 FILLER_13_102 ();
 sg13g2_decap_4 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_120 ();
 sg13g2_fill_1 FILLER_13_154 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_188 ();
 sg13g2_decap_4 FILLER_13_195 ();
 sg13g2_fill_2 FILLER_13_199 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_207 ();
 sg13g2_decap_4 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_319 ();
 sg13g2_fill_2 FILLER_13_325 ();
 sg13g2_fill_1 FILLER_13_327 ();
 sg13g2_fill_2 FILLER_13_359 ();
 sg13g2_fill_1 FILLER_13_361 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_2 FILLER_14_75 ();
 sg13g2_fill_1 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_fill_2 FILLER_14_133 ();
 sg13g2_fill_1 FILLER_14_135 ();
 sg13g2_fill_2 FILLER_14_160 ();
 sg13g2_fill_2 FILLER_14_181 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_fill_1 FILLER_14_260 ();
 sg13g2_decap_4 FILLER_14_265 ();
 sg13g2_fill_2 FILLER_14_269 ();
 sg13g2_fill_1 FILLER_14_306 ();
 sg13g2_fill_1 FILLER_14_321 ();
 sg13g2_fill_2 FILLER_14_339 ();
 sg13g2_fill_1 FILLER_14_341 ();
 sg13g2_fill_2 FILLER_14_351 ();
 sg13g2_fill_1 FILLER_14_353 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_51 ();
 sg13g2_fill_2 FILLER_15_72 ();
 sg13g2_decap_4 FILLER_15_95 ();
 sg13g2_decap_4 FILLER_15_103 ();
 sg13g2_fill_2 FILLER_15_107 ();
 sg13g2_decap_8 FILLER_15_118 ();
 sg13g2_fill_2 FILLER_15_125 ();
 sg13g2_fill_2 FILLER_15_150 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_1 FILLER_15_171 ();
 sg13g2_fill_1 FILLER_15_183 ();
 sg13g2_decap_4 FILLER_15_192 ();
 sg13g2_decap_8 FILLER_15_205 ();
 sg13g2_fill_2 FILLER_15_212 ();
 sg13g2_fill_1 FILLER_15_214 ();
 sg13g2_fill_1 FILLER_15_229 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_4 FILLER_15_273 ();
 sg13g2_fill_2 FILLER_15_285 ();
 sg13g2_decap_8 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_298 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_11 ();
 sg13g2_fill_1 FILLER_16_39 ();
 sg13g2_fill_2 FILLER_16_60 ();
 sg13g2_fill_1 FILLER_16_62 ();
 sg13g2_fill_1 FILLER_16_76 ();
 sg13g2_fill_2 FILLER_16_89 ();
 sg13g2_fill_1 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_120 ();
 sg13g2_fill_1 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_205 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_fill_2 FILLER_16_224 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_232 ();
 sg13g2_fill_1 FILLER_16_234 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_271 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_decap_8 FILLER_16_297 ();
 sg13g2_decap_4 FILLER_16_304 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_fill_2 FILLER_16_377 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_2 FILLER_17_29 ();
 sg13g2_fill_1 FILLER_17_31 ();
 sg13g2_fill_2 FILLER_17_55 ();
 sg13g2_decap_4 FILLER_17_81 ();
 sg13g2_fill_2 FILLER_17_85 ();
 sg13g2_decap_8 FILLER_17_96 ();
 sg13g2_fill_2 FILLER_17_117 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_2 FILLER_17_155 ();
 sg13g2_fill_1 FILLER_17_157 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_fill_2 FILLER_17_185 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_fill_1 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_248 ();
 sg13g2_fill_2 FILLER_17_270 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_357 ();
 sg13g2_fill_2 FILLER_17_367 ();
 sg13g2_fill_2 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_11 ();
 sg13g2_fill_1 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_38 ();
 sg13g2_fill_2 FILLER_18_57 ();
 sg13g2_fill_2 FILLER_18_69 ();
 sg13g2_fill_1 FILLER_18_79 ();
 sg13g2_fill_2 FILLER_18_88 ();
 sg13g2_fill_2 FILLER_18_111 ();
 sg13g2_fill_1 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_4 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_247 ();
 sg13g2_fill_2 FILLER_18_254 ();
 sg13g2_fill_1 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_fill_1 FILLER_18_295 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_4 FILLER_18_308 ();
 sg13g2_fill_1 FILLER_18_312 ();
 sg13g2_decap_4 FILLER_18_336 ();
 sg13g2_fill_1 FILLER_18_348 ();
 sg13g2_fill_2 FILLER_18_359 ();
 sg13g2_fill_2 FILLER_18_369 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_18_388 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_100 ();
 sg13g2_decap_4 FILLER_19_115 ();
 sg13g2_fill_1 FILLER_19_119 ();
 sg13g2_fill_1 FILLER_19_138 ();
 sg13g2_decap_4 FILLER_19_233 ();
 sg13g2_fill_1 FILLER_19_237 ();
 sg13g2_decap_4 FILLER_19_291 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_decap_4 FILLER_19_306 ();
 sg13g2_fill_2 FILLER_19_314 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_fill_2 FILLER_19_345 ();
 sg13g2_fill_1 FILLER_19_347 ();
 sg13g2_fill_1 FILLER_19_391 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_45 ();
 sg13g2_fill_1 FILLER_20_51 ();
 sg13g2_fill_1 FILLER_20_99 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_decap_8 FILLER_20_181 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_fill_1 FILLER_20_194 ();
 sg13g2_fill_2 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_225 ();
 sg13g2_decap_8 FILLER_20_232 ();
 sg13g2_decap_4 FILLER_20_251 ();
 sg13g2_fill_1 FILLER_20_255 ();
 sg13g2_decap_4 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_fill_1 FILLER_20_275 ();
 sg13g2_decap_4 FILLER_20_296 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_fill_2 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_4 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_82 ();
 sg13g2_fill_1 FILLER_21_99 ();
 sg13g2_fill_2 FILLER_21_104 ();
 sg13g2_fill_1 FILLER_21_106 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_fill_2 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_decap_4 FILLER_21_133 ();
 sg13g2_fill_2 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_fill_2 FILLER_21_157 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_227 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_287 ();
 sg13g2_decap_4 FILLER_21_312 ();
 sg13g2_fill_1 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_4 FILLER_21_345 ();
 sg13g2_fill_1 FILLER_21_349 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_47 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_decap_4 FILLER_22_81 ();
 sg13g2_fill_2 FILLER_22_85 ();
 sg13g2_fill_2 FILLER_22_176 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_fill_1 FILLER_22_217 ();
 sg13g2_decap_4 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_227 ();
 sg13g2_fill_1 FILLER_22_234 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_fill_2 FILLER_22_272 ();
 sg13g2_fill_2 FILLER_22_278 ();
 sg13g2_decap_8 FILLER_22_297 ();
 sg13g2_decap_4 FILLER_22_304 ();
 sg13g2_fill_1 FILLER_22_308 ();
 sg13g2_fill_2 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_11 ();
 sg13g2_fill_1 FILLER_23_17 ();
 sg13g2_fill_2 FILLER_23_37 ();
 sg13g2_fill_1 FILLER_23_39 ();
 sg13g2_decap_4 FILLER_23_60 ();
 sg13g2_fill_1 FILLER_23_73 ();
 sg13g2_decap_8 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_90 ();
 sg13g2_decap_8 FILLER_23_95 ();
 sg13g2_decap_4 FILLER_23_102 ();
 sg13g2_fill_2 FILLER_23_106 ();
 sg13g2_fill_2 FILLER_23_121 ();
 sg13g2_fill_1 FILLER_23_123 ();
 sg13g2_fill_1 FILLER_23_137 ();
 sg13g2_fill_1 FILLER_23_157 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_174 ();
 sg13g2_decap_4 FILLER_23_179 ();
 sg13g2_fill_2 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_230 ();
 sg13g2_decap_4 FILLER_23_248 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_267 ();
 sg13g2_decap_8 FILLER_23_282 ();
 sg13g2_decap_4 FILLER_23_289 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_fill_2 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_fill_1 FILLER_23_351 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_57 ();
 sg13g2_fill_1 FILLER_24_66 ();
 sg13g2_fill_2 FILLER_24_75 ();
 sg13g2_fill_1 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_88 ();
 sg13g2_decap_4 FILLER_24_124 ();
 sg13g2_fill_1 FILLER_24_164 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_decap_8 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_268 ();
 sg13g2_fill_2 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_346 ();
 sg13g2_fill_2 FILLER_24_355 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_11 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_80 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_decap_4 FILLER_25_125 ();
 sg13g2_fill_2 FILLER_25_129 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_fill_1 FILLER_25_190 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_decap_4 FILLER_25_222 ();
 sg13g2_decap_4 FILLER_25_230 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_decap_4 FILLER_25_247 ();
 sg13g2_fill_1 FILLER_25_251 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_decap_4 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_273 ();
 sg13g2_fill_2 FILLER_25_279 ();
 sg13g2_fill_2 FILLER_25_292 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_fill_1 FILLER_25_309 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_346 ();
 sg13g2_fill_1 FILLER_25_364 ();
 sg13g2_fill_2 FILLER_25_381 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_27 ();
 sg13g2_fill_1 FILLER_26_74 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_4 FILLER_26_109 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_174 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_decap_4 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_decap_4 FILLER_26_235 ();
 sg13g2_fill_2 FILLER_26_257 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_15 ();
 sg13g2_fill_2 FILLER_27_77 ();
 sg13g2_decap_4 FILLER_27_96 ();
 sg13g2_fill_2 FILLER_27_100 ();
 sg13g2_decap_4 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_fill_2 FILLER_27_149 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_160 ();
 sg13g2_decap_8 FILLER_27_216 ();
 sg13g2_fill_2 FILLER_27_233 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_fill_2 FILLER_27_264 ();
 sg13g2_fill_1 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_367 ();
 sg13g2_fill_1 FILLER_27_377 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_28_26 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_decap_4 FILLER_28_108 ();
 sg13g2_fill_2 FILLER_28_117 ();
 sg13g2_decap_4 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_fill_1 FILLER_28_169 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_decap_8 FILLER_28_212 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_decap_4 FILLER_28_239 ();
 sg13g2_fill_2 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_328 ();
 sg13g2_fill_2 FILLER_28_381 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_64 ();
 sg13g2_fill_2 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_78 ();
 sg13g2_fill_2 FILLER_29_88 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_2 FILLER_29_122 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_decap_8 FILLER_29_135 ();
 sg13g2_decap_4 FILLER_29_142 ();
 sg13g2_decap_8 FILLER_29_183 ();
 sg13g2_decap_8 FILLER_29_190 ();
 sg13g2_fill_2 FILLER_29_197 ();
 sg13g2_decap_8 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_fill_2 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_323 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_fill_1 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_29_357 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_38 ();
 sg13g2_fill_1 FILLER_30_40 ();
 sg13g2_decap_4 FILLER_30_79 ();
 sg13g2_fill_2 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_107 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_fill_1 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_228 ();
 sg13g2_fill_2 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_289 ();
 sg13g2_fill_1 FILLER_30_291 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_355 ();
 sg13g2_fill_2 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_33 ();
 sg13g2_fill_2 FILLER_31_59 ();
 sg13g2_fill_2 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_103 ();
 sg13g2_fill_1 FILLER_31_114 ();
 sg13g2_decap_8 FILLER_31_125 ();
 sg13g2_fill_1 FILLER_31_132 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_fill_1 FILLER_31_210 ();
 sg13g2_decap_4 FILLER_31_216 ();
 sg13g2_decap_4 FILLER_31_241 ();
 sg13g2_decap_4 FILLER_31_248 ();
 sg13g2_fill_2 FILLER_31_334 ();
 sg13g2_fill_1 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_367 ();
 sg13g2_fill_2 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_109 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_160 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_decap_4 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_259 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_fill_1 FILLER_32_370 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_30 ();
 sg13g2_fill_2 FILLER_33_41 ();
 sg13g2_fill_2 FILLER_33_71 ();
 sg13g2_fill_1 FILLER_33_82 ();
 sg13g2_decap_8 FILLER_33_107 ();
 sg13g2_fill_2 FILLER_33_114 ();
 sg13g2_fill_1 FILLER_33_130 ();
 sg13g2_decap_4 FILLER_33_135 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_4 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_2 FILLER_33_195 ();
 sg13g2_fill_1 FILLER_33_197 ();
 sg13g2_fill_2 FILLER_33_212 ();
 sg13g2_fill_1 FILLER_33_214 ();
 sg13g2_fill_2 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_fill_2 FILLER_33_385 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_73 ();
 sg13g2_fill_2 FILLER_34_104 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_decap_8 FILLER_34_129 ();
 sg13g2_decap_8 FILLER_34_136 ();
 sg13g2_decap_4 FILLER_34_143 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_fill_1 FILLER_34_208 ();
 sg13g2_decap_8 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_fill_2 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_366 ();
 sg13g2_fill_1 FILLER_34_368 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_decap_4 FILLER_35_138 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_decap_4 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_fill_1 FILLER_35_179 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_296 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_fill_2 FILLER_35_397 ();
 sg13g2_fill_1 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_40 ();
 sg13g2_fill_1 FILLER_36_101 ();
 sg13g2_fill_2 FILLER_36_111 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_decap_8 FILLER_36_132 ();
 sg13g2_fill_1 FILLER_36_139 ();
 sg13g2_fill_2 FILLER_36_180 ();
 sg13g2_fill_1 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_205 ();
 sg13g2_fill_2 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_fill_2 FILLER_36_267 ();
 sg13g2_fill_1 FILLER_36_278 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_132 ();
 sg13g2_fill_1 FILLER_37_134 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_fill_2 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_200 ();
 sg13g2_fill_1 FILLER_37_214 ();
 sg13g2_fill_1 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_313 ();
 sg13g2_fill_2 FILLER_37_369 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_23 ();
 sg13g2_fill_1 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_2 FILLER_38_149 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_187 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_240 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_265 ();
 sg13g2_fill_2 FILLER_38_275 ();
 sg13g2_fill_1 FILLER_38_277 ();
 sg13g2_fill_1 FILLER_38_321 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
endmodule

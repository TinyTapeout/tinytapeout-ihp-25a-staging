module tt_um_levenshtein (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire \arbiter.cyc ;
 wire \arbiter.gnt ;
 wire \arbiter.wbm_ack_i ;
 wire \arbiter.wbm_dat_i[0] ;
 wire \arbiter.wbm_dat_i[1] ;
 wire \arbiter.wbm_dat_i[2] ;
 wire \arbiter.wbm_dat_i[3] ;
 wire \arbiter.wbm_dat_i[4] ;
 wire \arbiter.wbm_dat_i[5] ;
 wire \arbiter.wbm_dat_i[6] ;
 wire \arbiter.wbm_dat_i[7] ;
 wire \arbiter.wbs0_adr_i[0] ;
 wire \arbiter.wbs0_adr_i[10] ;
 wire \arbiter.wbs0_adr_i[11] ;
 wire \arbiter.wbs0_adr_i[12] ;
 wire \arbiter.wbs0_adr_i[13] ;
 wire \arbiter.wbs0_adr_i[14] ;
 wire \arbiter.wbs0_adr_i[15] ;
 wire \arbiter.wbs0_adr_i[16] ;
 wire \arbiter.wbs0_adr_i[17] ;
 wire \arbiter.wbs0_adr_i[18] ;
 wire \arbiter.wbs0_adr_i[19] ;
 wire \arbiter.wbs0_adr_i[1] ;
 wire \arbiter.wbs0_adr_i[20] ;
 wire \arbiter.wbs0_adr_i[21] ;
 wire \arbiter.wbs0_adr_i[22] ;
 wire \arbiter.wbs0_adr_i[2] ;
 wire \arbiter.wbs0_adr_i[3] ;
 wire \arbiter.wbs0_adr_i[4] ;
 wire \arbiter.wbs0_adr_i[5] ;
 wire \arbiter.wbs0_adr_i[6] ;
 wire \arbiter.wbs0_adr_i[7] ;
 wire \arbiter.wbs0_adr_i[8] ;
 wire \arbiter.wbs0_adr_i[9] ;
 wire \arbiter.wbs0_dat_i[0] ;
 wire \arbiter.wbs0_dat_i[1] ;
 wire \arbiter.wbs0_dat_i[2] ;
 wire \arbiter.wbs0_dat_i[3] ;
 wire \arbiter.wbs0_dat_i[4] ;
 wire \arbiter.wbs0_dat_i[5] ;
 wire \arbiter.wbs0_dat_i[6] ;
 wire \arbiter.wbs0_dat_i[7] ;
 wire \arbiter.wbs0_we_i ;
 wire \arbiter.wbs1_cyc_i ;
 wire ctrl_slave_ack;
 wire \intercon.wbs_cyc_i ;
 wire \levenshtein_ctrl.best_distance[0] ;
 wire \levenshtein_ctrl.best_distance[1] ;
 wire \levenshtein_ctrl.best_distance[2] ;
 wire \levenshtein_ctrl.best_distance[3] ;
 wire \levenshtein_ctrl.best_distance[4] ;
 wire \levenshtein_ctrl.best_distance[5] ;
 wire \levenshtein_ctrl.best_distance[6] ;
 wire \levenshtein_ctrl.best_distance[7] ;
 wire \levenshtein_ctrl.best_idx[0] ;
 wire \levenshtein_ctrl.best_idx[10] ;
 wire \levenshtein_ctrl.best_idx[11] ;
 wire \levenshtein_ctrl.best_idx[12] ;
 wire \levenshtein_ctrl.best_idx[13] ;
 wire \levenshtein_ctrl.best_idx[14] ;
 wire \levenshtein_ctrl.best_idx[15] ;
 wire \levenshtein_ctrl.best_idx[1] ;
 wire \levenshtein_ctrl.best_idx[2] ;
 wire \levenshtein_ctrl.best_idx[3] ;
 wire \levenshtein_ctrl.best_idx[4] ;
 wire \levenshtein_ctrl.best_idx[5] ;
 wire \levenshtein_ctrl.best_idx[6] ;
 wire \levenshtein_ctrl.best_idx[7] ;
 wire \levenshtein_ctrl.best_idx[8] ;
 wire \levenshtein_ctrl.best_idx[9] ;
 wire \levenshtein_ctrl.d[0] ;
 wire \levenshtein_ctrl.d[1] ;
 wire \levenshtein_ctrl.d[2] ;
 wire \levenshtein_ctrl.d[3] ;
 wire \levenshtein_ctrl.d[4] ;
 wire \levenshtein_ctrl.d[5] ;
 wire \levenshtein_ctrl.d[6] ;
 wire \levenshtein_ctrl.d[7] ;
 wire \levenshtein_ctrl.dict_address[0] ;
 wire \levenshtein_ctrl.dict_address[10] ;
 wire \levenshtein_ctrl.dict_address[11] ;
 wire \levenshtein_ctrl.dict_address[12] ;
 wire \levenshtein_ctrl.dict_address[13] ;
 wire \levenshtein_ctrl.dict_address[14] ;
 wire \levenshtein_ctrl.dict_address[15] ;
 wire \levenshtein_ctrl.dict_address[16] ;
 wire \levenshtein_ctrl.dict_address[17] ;
 wire \levenshtein_ctrl.dict_address[18] ;
 wire \levenshtein_ctrl.dict_address[19] ;
 wire \levenshtein_ctrl.dict_address[1] ;
 wire \levenshtein_ctrl.dict_address[20] ;
 wire \levenshtein_ctrl.dict_address[2] ;
 wire \levenshtein_ctrl.dict_address[3] ;
 wire \levenshtein_ctrl.dict_address[4] ;
 wire \levenshtein_ctrl.dict_address[5] ;
 wire \levenshtein_ctrl.dict_address[6] ;
 wire \levenshtein_ctrl.dict_address[7] ;
 wire \levenshtein_ctrl.dict_address[8] ;
 wire \levenshtein_ctrl.dict_address[9] ;
 wire \levenshtein_ctrl.enabled ;
 wire \levenshtein_ctrl.idx[0] ;
 wire \levenshtein_ctrl.idx[10] ;
 wire \levenshtein_ctrl.idx[11] ;
 wire \levenshtein_ctrl.idx[12] ;
 wire \levenshtein_ctrl.idx[13] ;
 wire \levenshtein_ctrl.idx[14] ;
 wire \levenshtein_ctrl.idx[15] ;
 wire \levenshtein_ctrl.idx[1] ;
 wire \levenshtein_ctrl.idx[2] ;
 wire \levenshtein_ctrl.idx[3] ;
 wire \levenshtein_ctrl.idx[4] ;
 wire \levenshtein_ctrl.idx[5] ;
 wire \levenshtein_ctrl.idx[6] ;
 wire \levenshtein_ctrl.idx[7] ;
 wire \levenshtein_ctrl.idx[8] ;
 wire \levenshtein_ctrl.idx[9] ;
 wire \levenshtein_ctrl.next_symbol[0] ;
 wire \levenshtein_ctrl.next_symbol[1] ;
 wire \levenshtein_ctrl.next_symbol[2] ;
 wire \levenshtein_ctrl.next_symbol[3] ;
 wire \levenshtein_ctrl.next_symbol[4] ;
 wire \levenshtein_ctrl.next_symbol[5] ;
 wire \levenshtein_ctrl.next_symbol[6] ;
 wire \levenshtein_ctrl.next_symbol[7] ;
 wire \levenshtein_ctrl.pm[0] ;
 wire \levenshtein_ctrl.pm[10] ;
 wire \levenshtein_ctrl.pm[11] ;
 wire \levenshtein_ctrl.pm[12] ;
 wire \levenshtein_ctrl.pm[13] ;
 wire \levenshtein_ctrl.pm[14] ;
 wire \levenshtein_ctrl.pm[15] ;
 wire \levenshtein_ctrl.pm[1] ;
 wire \levenshtein_ctrl.pm[2] ;
 wire \levenshtein_ctrl.pm[3] ;
 wire \levenshtein_ctrl.pm[4] ;
 wire \levenshtein_ctrl.pm[5] ;
 wire \levenshtein_ctrl.pm[6] ;
 wire \levenshtein_ctrl.pm[7] ;
 wire \levenshtein_ctrl.pm[8] ;
 wire \levenshtein_ctrl.pm[9] ;
 wire \levenshtein_ctrl.sram_config[0] ;
 wire \levenshtein_ctrl.sram_config[1] ;
 wire \levenshtein_ctrl.state[0] ;
 wire \levenshtein_ctrl.state[1] ;
 wire \levenshtein_ctrl.state[2] ;
 wire \levenshtein_ctrl.state[3] ;
 wire \levenshtein_ctrl.state[4] ;
 wire \levenshtein_ctrl.state[5] ;
 wire \levenshtein_ctrl.state[6] ;
 wire \levenshtein_ctrl.state[7] ;
 wire \levenshtein_ctrl.symbol[0] ;
 wire \levenshtein_ctrl.symbol[1] ;
 wire \levenshtein_ctrl.symbol[2] ;
 wire \levenshtein_ctrl.symbol[3] ;
 wire \levenshtein_ctrl.symbol[4] ;
 wire \levenshtein_ctrl.symbol[5] ;
 wire \levenshtein_ctrl.symbol[6] ;
 wire \levenshtein_ctrl.symbol[7] ;
 wire \levenshtein_ctrl.symbol_idx[0] ;
 wire \levenshtein_ctrl.symbol_idx[1] ;
 wire \levenshtein_ctrl.symbols[10] ;
 wire \levenshtein_ctrl.symbols[11] ;
 wire \levenshtein_ctrl.symbols[12] ;
 wire \levenshtein_ctrl.symbols[13] ;
 wire \levenshtein_ctrl.symbols[14] ;
 wire \levenshtein_ctrl.symbols[15] ;
 wire \levenshtein_ctrl.symbols[16] ;
 wire \levenshtein_ctrl.symbols[17] ;
 wire \levenshtein_ctrl.symbols[18] ;
 wire \levenshtein_ctrl.symbols[19] ;
 wire \levenshtein_ctrl.symbols[20] ;
 wire \levenshtein_ctrl.symbols[21] ;
 wire \levenshtein_ctrl.symbols[22] ;
 wire \levenshtein_ctrl.symbols[23] ;
 wire \levenshtein_ctrl.symbols[8] ;
 wire \levenshtein_ctrl.symbols[9] ;
 wire \levenshtein_ctrl.vn[0] ;
 wire \levenshtein_ctrl.vn[10] ;
 wire \levenshtein_ctrl.vn[11] ;
 wire \levenshtein_ctrl.vn[12] ;
 wire \levenshtein_ctrl.vn[13] ;
 wire \levenshtein_ctrl.vn[14] ;
 wire \levenshtein_ctrl.vn[15] ;
 wire \levenshtein_ctrl.vn[1] ;
 wire \levenshtein_ctrl.vn[2] ;
 wire \levenshtein_ctrl.vn[3] ;
 wire \levenshtein_ctrl.vn[4] ;
 wire \levenshtein_ctrl.vn[5] ;
 wire \levenshtein_ctrl.vn[6] ;
 wire \levenshtein_ctrl.vn[7] ;
 wire \levenshtein_ctrl.vn[8] ;
 wire \levenshtein_ctrl.vn[9] ;
 wire \levenshtein_ctrl.vp[0] ;
 wire \levenshtein_ctrl.vp[10] ;
 wire \levenshtein_ctrl.vp[11] ;
 wire \levenshtein_ctrl.vp[12] ;
 wire \levenshtein_ctrl.vp[13] ;
 wire \levenshtein_ctrl.vp[14] ;
 wire \levenshtein_ctrl.vp[15] ;
 wire \levenshtein_ctrl.vp[1] ;
 wire \levenshtein_ctrl.vp[2] ;
 wire \levenshtein_ctrl.vp[3] ;
 wire \levenshtein_ctrl.vp[4] ;
 wire \levenshtein_ctrl.vp[5] ;
 wire \levenshtein_ctrl.vp[6] ;
 wire \levenshtein_ctrl.vp[7] ;
 wire \levenshtein_ctrl.vp[8] ;
 wire \levenshtein_ctrl.vp[9] ;
 wire \levenshtein_ctrl.word_length_reg[0] ;
 wire \levenshtein_ctrl.word_length_reg[1] ;
 wire \levenshtein_ctrl.word_length_reg[2] ;
 wire \levenshtein_ctrl.word_length_reg[3] ;
 wire \spi.counter[0] ;
 wire \spi.counter[1] ;
 wire \spi.counter[2] ;
 wire \spi.counter[3] ;
 wire \spi.counter[4] ;
 wire \spi.last_sck ;
 wire \spi.miso ;
 wire \spi.mosi ;
 wire \spi.mosi_sync[0] ;
 wire \spi.sck ;
 wire \spi.sck_sync[0] ;
 wire \spi.ss_n ;
 wire \spi.ss_n_sync[0] ;
 wire \spi.state[0] ;
 wire \spi.state[2] ;
 wire \spi_ctrl.bit_counter[0] ;
 wire \spi_ctrl.bit_counter[1] ;
 wire \spi_ctrl.bit_counter[2] ;
 wire \spi_ctrl.bit_counter[3] ;
 wire \spi_ctrl.bit_counter[4] ;
 wire \spi_ctrl.cs2_n ;
 wire \spi_ctrl.cs3_n ;
 wire \spi_ctrl.cs_n ;
 wire \spi_ctrl.sck ;
 wire \spi_ctrl.ss_n ;
 wire net258;
 wire net259;
 wire net260;
 wire clknet_leaf_0_clk;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;

 sg13g2_inv_1 _1744_ (.Y(_0929_),
    .A(net404));
 sg13g2_inv_1 _1745_ (.Y(_0930_),
    .A(net634));
 sg13g2_inv_1 _1746_ (.Y(_0931_),
    .A(net606));
 sg13g2_inv_2 _1747_ (.Y(_0932_),
    .A(net408));
 sg13g2_inv_1 _1748_ (.Y(_0933_),
    .A(net418));
 sg13g2_inv_1 _1749_ (.Y(_0934_),
    .A(net540));
 sg13g2_inv_1 _1750_ (.Y(_0935_),
    .A(net641));
 sg13g2_inv_1 _1751_ (.Y(_0936_),
    .A(net678));
 sg13g2_inv_2 _1752_ (.Y(_0937_),
    .A(\arbiter.wbs0_we_i ));
 sg13g2_inv_1 _1753_ (.Y(_0938_),
    .A(net515));
 sg13g2_inv_1 _1754_ (.Y(_0939_),
    .A(\levenshtein_ctrl.d[0] ));
 sg13g2_inv_1 _1755_ (.Y(_0940_),
    .A(net692));
 sg13g2_inv_1 _1756_ (.Y(_0941_),
    .A(\levenshtein_ctrl.d[1] ));
 sg13g2_inv_1 _1757_ (.Y(_0942_),
    .A(net701));
 sg13g2_inv_1 _1758_ (.Y(_0943_),
    .A(\levenshtein_ctrl.d[2] ));
 sg13g2_inv_1 _1759_ (.Y(_0944_),
    .A(net709));
 sg13g2_inv_2 _1760_ (.Y(_0945_),
    .A(\levenshtein_ctrl.d[3] ));
 sg13g2_inv_1 _1761_ (.Y(_0946_),
    .A(net578));
 sg13g2_inv_2 _1762_ (.Y(_0947_),
    .A(\levenshtein_ctrl.d[4] ));
 sg13g2_inv_1 _1763_ (.Y(_0948_),
    .A(net538));
 sg13g2_inv_1 _1764_ (.Y(_0949_),
    .A(\levenshtein_ctrl.d[5] ));
 sg13g2_inv_1 _1765_ (.Y(_0950_),
    .A(net541));
 sg13g2_inv_1 _1766_ (.Y(_0951_),
    .A(\levenshtein_ctrl.d[6] ));
 sg13g2_inv_1 _1767_ (.Y(_0952_),
    .A(net568));
 sg13g2_inv_1 _1768_ (.Y(_0953_),
    .A(\levenshtein_ctrl.d[7] ));
 sg13g2_inv_1 _1769_ (.Y(_0954_),
    .A(\levenshtein_ctrl.state[4] ));
 sg13g2_inv_2 _1770_ (.Y(_0955_),
    .A(\levenshtein_ctrl.state[6] ));
 sg13g2_inv_1 _1771_ (.Y(_0956_),
    .A(net314));
 sg13g2_inv_1 _1772_ (.Y(_0957_),
    .A(net559));
 sg13g2_inv_1 _1773_ (.Y(_0958_),
    .A(net582));
 sg13g2_inv_1 _1774_ (.Y(_0959_),
    .A(net320));
 sg13g2_inv_1 _1775_ (.Y(_0960_),
    .A(net322));
 sg13g2_inv_1 _1776_ (.Y(_0961_),
    .A(net478));
 sg13g2_inv_1 _1777_ (.Y(_0962_),
    .A(net439));
 sg13g2_inv_4 _1778_ (.A(net661),
    .Y(_0963_));
 sg13g2_inv_1 _1779_ (.Y(_0964_),
    .A(_0066_));
 sg13g2_inv_1 _1780_ (.Y(_0965_),
    .A(\levenshtein_ctrl.dict_address[6] ));
 sg13g2_inv_1 _1781_ (.Y(_0966_),
    .A(\levenshtein_ctrl.dict_address[7] ));
 sg13g2_inv_1 _1782_ (.Y(_0967_),
    .A(_0018_));
 sg13g2_inv_1 _1783_ (.Y(_0968_),
    .A(\arbiter.wbs0_adr_i[10] ));
 sg13g2_inv_1 _1784_ (.Y(_0969_),
    .A(net502));
 sg13g2_inv_1 _1785_ (.Y(_0970_),
    .A(\levenshtein_ctrl.dict_address[13] ));
 sg13g2_inv_2 _1786_ (.Y(_0971_),
    .A(net413));
 sg13g2_inv_2 _1787_ (.Y(_0972_),
    .A(net434));
 sg13g2_inv_1 _1788_ (.Y(_0973_),
    .A(net283));
 sg13g2_inv_1 _1789_ (.Y(_0974_),
    .A(\levenshtein_ctrl.vp[2] ));
 sg13g2_inv_1 _1790_ (.Y(_0975_),
    .A(\levenshtein_ctrl.vp[4] ));
 sg13g2_inv_1 _1791_ (.Y(_0976_),
    .A(\levenshtein_ctrl.vp[5] ));
 sg13g2_inv_1 _1792_ (.Y(_0977_),
    .A(net308));
 sg13g2_inv_1 _1793_ (.Y(_0978_),
    .A(\levenshtein_ctrl.vp[6] ));
 sg13g2_inv_1 _1794_ (.Y(_0979_),
    .A(\levenshtein_ctrl.vp[7] ));
 sg13g2_inv_1 _1795_ (.Y(_0980_),
    .A(\levenshtein_ctrl.vp[9] ));
 sg13g2_inv_1 _1796_ (.Y(_0981_),
    .A(\levenshtein_ctrl.vn[11] ));
 sg13g2_inv_1 _1797_ (.Y(_0982_),
    .A(\levenshtein_ctrl.vn[12] ));
 sg13g2_inv_1 _1798_ (.Y(_0983_),
    .A(\levenshtein_ctrl.vn[13] ));
 sg13g2_inv_1 _1799_ (.Y(_0984_),
    .A(\levenshtein_ctrl.vp[14] ));
 sg13g2_inv_1 _1800_ (.Y(_0985_),
    .A(net438));
 sg13g2_inv_1 _1801_ (.Y(_0986_),
    .A(\levenshtein_ctrl.idx[0] ));
 sg13g2_inv_1 _1802_ (.Y(_0987_),
    .A(net520));
 sg13g2_nor2b_1 _1803_ (.A(\spi_ctrl.ss_n ),
    .B_N(\levenshtein_ctrl.sram_config[1] ),
    .Y(_0988_));
 sg13g2_nor2b_1 _1804_ (.A(\spi_ctrl.ss_n ),
    .B_N(\levenshtein_ctrl.sram_config[0] ),
    .Y(_0989_));
 sg13g2_nand2_1 _1805_ (.Y(\spi_ctrl.cs3_n ),
    .A(\levenshtein_ctrl.sram_config[0] ),
    .B(_0988_));
 sg13g2_nand2b_1 _1806_ (.Y(\spi_ctrl.cs2_n ),
    .B(_0988_),
    .A_N(\levenshtein_ctrl.sram_config[0] ));
 sg13g2_nand2b_1 _1807_ (.Y(\spi_ctrl.cs_n ),
    .B(_0989_),
    .A_N(\levenshtein_ctrl.sram_config[1] ));
 sg13g2_and2_1 _1808_ (.A(\levenshtein_ctrl.enabled ),
    .B(net437),
    .X(_0990_));
 sg13g2_nand2_2 _1809_ (.Y(_0991_),
    .A(net416),
    .B(net435));
 sg13g2_nor4_1 _1810_ (.A(\arbiter.wbs0_adr_i[20] ),
    .B(\arbiter.wbs0_adr_i[5] ),
    .C(\arbiter.wbs0_adr_i[9] ),
    .D(\arbiter.wbs0_adr_i[13] ),
    .Y(_0992_));
 sg13g2_nor4_1 _1811_ (.A(\arbiter.wbs0_adr_i[4] ),
    .B(\arbiter.wbs0_adr_i[8] ),
    .C(\arbiter.wbs0_adr_i[12] ),
    .D(\arbiter.wbs0_adr_i[16] ),
    .Y(_0993_));
 sg13g2_and2_1 _1812_ (.A(_0992_),
    .B(_0993_),
    .X(_0994_));
 sg13g2_nor4_1 _1813_ (.A(\arbiter.wbs0_adr_i[7] ),
    .B(\arbiter.wbs0_adr_i[11] ),
    .C(\arbiter.wbs0_adr_i[15] ),
    .D(\arbiter.wbs0_adr_i[19] ),
    .Y(_0995_));
 sg13g2_nor4_1 _1814_ (.A(\arbiter.wbs0_adr_i[14] ),
    .B(\arbiter.wbs0_adr_i[18] ),
    .C(\arbiter.wbs0_adr_i[22] ),
    .D(\arbiter.wbs0_adr_i[3] ),
    .Y(_0996_));
 sg13g2_nor4_1 _1815_ (.A(\arbiter.wbs0_adr_i[17] ),
    .B(\arbiter.wbs0_adr_i[21] ),
    .C(\arbiter.wbs0_adr_i[6] ),
    .D(\arbiter.wbs0_adr_i[10] ),
    .Y(_0997_));
 sg13g2_and3_1 _1816_ (.X(_0998_),
    .A(_0995_),
    .B(_0996_),
    .C(_0997_));
 sg13g2_and2_1 _1817_ (.A(_0994_),
    .B(_0998_),
    .X(_0999_));
 sg13g2_nand2_1 _1818_ (.Y(_1000_),
    .A(_0994_),
    .B(_0998_));
 sg13g2_nor3_2 _1819_ (.A(net727),
    .B(net733),
    .C(_1000_),
    .Y(_1001_));
 sg13g2_and2_1 _1820_ (.A(net436),
    .B(_1001_),
    .X(_0086_));
 sg13g2_nor2_1 _1821_ (.A(\arbiter.wbs0_adr_i[0] ),
    .B(\arbiter.wbs0_adr_i[1] ),
    .Y(_1002_));
 sg13g2_nand2_2 _1822_ (.Y(_1003_),
    .A(_0018_),
    .B(_1002_));
 sg13g2_inv_1 _1823_ (.Y(_1004_),
    .A(_1003_));
 sg13g2_nor2_1 _1824_ (.A(\levenshtein_ctrl.enabled ),
    .B(net431),
    .Y(_1005_));
 sg13g2_nand2b_1 _1825_ (.Y(_1006_),
    .B(net435),
    .A_N(net416));
 sg13g2_a21oi_1 _1826_ (.A1(_1003_),
    .A2(_1005_),
    .Y(_1007_),
    .B1(_0937_));
 sg13g2_nand2_1 _1827_ (.Y(_1008_),
    .A(\arbiter.wbs0_we_i ),
    .B(_1001_));
 sg13g2_inv_1 _1828_ (.Y(_1009_),
    .A(_1008_));
 sg13g2_a22oi_1 _1829_ (.Y(_1010_),
    .B1(_0086_),
    .B2(_0056_),
    .A2(_1001_),
    .A1(\arbiter.wbs0_we_i ));
 sg13g2_or2_1 _1830_ (.X(_1011_),
    .B(_1010_),
    .A(_1007_));
 sg13g2_o21ai_1 _1831_ (.B1(_1011_),
    .Y(_1012_),
    .A1(net396),
    .A2(_0086_));
 sg13g2_nor2_2 _1832_ (.A(net431),
    .B(_0056_),
    .Y(_1013_));
 sg13g2_nand2b_1 _1833_ (.Y(_1014_),
    .B(net436),
    .A_N(_0056_));
 sg13g2_nor2b_1 _1834_ (.A(\arbiter.gnt ),
    .B_N(\arbiter.wbm_ack_i ),
    .Y(_1015_));
 sg13g2_a21oi_1 _1835_ (.A1(\arbiter.wbs1_cyc_i ),
    .A2(net394),
    .Y(_1016_),
    .B1(_1014_));
 sg13g2_o21ai_1 _1836_ (.B1(\levenshtein_ctrl.state[3] ),
    .Y(_1017_),
    .A1(_1012_),
    .A2(_1016_));
 sg13g2_nor2_1 _1837_ (.A(\levenshtein_ctrl.next_symbol[1] ),
    .B(\levenshtein_ctrl.next_symbol[4] ),
    .Y(_1018_));
 sg13g2_nor3_1 _1838_ (.A(\levenshtein_ctrl.next_symbol[5] ),
    .B(\levenshtein_ctrl.next_symbol[6] ),
    .C(\levenshtein_ctrl.next_symbol[7] ),
    .Y(_1019_));
 sg13g2_and2_1 _1839_ (.A(_1018_),
    .B(_1019_),
    .X(_1020_));
 sg13g2_nor2_1 _1840_ (.A(\levenshtein_ctrl.next_symbol[2] ),
    .B(\levenshtein_ctrl.next_symbol[3] ),
    .Y(_1021_));
 sg13g2_nand3_1 _1841_ (.B(_1020_),
    .C(_1021_),
    .A(\levenshtein_ctrl.next_symbol[0] ),
    .Y(_1022_));
 sg13g2_nor3_1 _1842_ (.A(\levenshtein_ctrl.next_symbol[0] ),
    .B(\levenshtein_ctrl.next_symbol[2] ),
    .C(\levenshtein_ctrl.next_symbol[3] ),
    .Y(_1023_));
 sg13g2_and2_2 _1843_ (.A(_1020_),
    .B(_1023_),
    .X(_1024_));
 sg13g2_nand3_1 _1844_ (.B(_1013_),
    .C(_1022_),
    .A(net570),
    .Y(_1025_));
 sg13g2_o21ai_1 _1845_ (.B1(_1017_),
    .Y(_0003_),
    .A1(_1024_),
    .A2(net571));
 sg13g2_and4_2 _1846_ (.A(net423),
    .B(_1018_),
    .C(_1019_),
    .D(_1023_),
    .X(_1026_));
 sg13g2_nand2_2 _1847_ (.Y(_1027_),
    .A(net423),
    .B(_1024_));
 sg13g2_nor2_1 _1848_ (.A(_0991_),
    .B(_1027_),
    .Y(_1028_));
 sg13g2_nor2_1 _1849_ (.A(\levenshtein_ctrl.symbol_idx[0] ),
    .B(net617),
    .Y(_1029_));
 sg13g2_nand2_1 _1850_ (.Y(_1030_),
    .A(net422),
    .B(_1013_));
 sg13g2_nand3_1 _1851_ (.B(_1013_),
    .C(_1029_),
    .A(net422),
    .Y(_1031_));
 sg13g2_o21ai_1 _1852_ (.B1(net425),
    .Y(_1032_),
    .A1(_0991_),
    .A2(_1016_));
 sg13g2_and2_1 _1853_ (.A(net416),
    .B(net423),
    .X(_1033_));
 sg13g2_nand2_1 _1854_ (.Y(_1034_),
    .A(net416),
    .B(net423));
 sg13g2_nand2_2 _1855_ (.Y(_1035_),
    .A(net423),
    .B(net397));
 sg13g2_and3_2 _1856_ (.X(_1036_),
    .A(net423),
    .B(net397),
    .C(_1024_));
 sg13g2_nand3_1 _1857_ (.B(net617),
    .C(_1036_),
    .A(\levenshtein_ctrl.symbol_idx[0] ),
    .Y(_1037_));
 sg13g2_nand3_1 _1858_ (.B(_1032_),
    .C(_1037_),
    .A(_1031_),
    .Y(_1038_));
 sg13g2_nor3_1 _1859_ (.A(net431),
    .B(_1003_),
    .C(_1008_),
    .Y(_1039_));
 sg13g2_nand3_1 _1860_ (.B(_1001_),
    .C(_1004_),
    .A(\arbiter.wbs0_we_i ),
    .Y(_1040_));
 sg13g2_a21o_1 _1861_ (.A2(_1039_),
    .A1(net711),
    .B1(_1038_),
    .X(_0000_));
 sg13g2_and2_1 _1862_ (.A(net396),
    .B(net394),
    .X(_1041_));
 sg13g2_nand2_2 _1863_ (.Y(_1042_),
    .A(net396),
    .B(net394));
 sg13g2_nand2b_1 _1864_ (.Y(_1043_),
    .B(net416),
    .A_N(net394));
 sg13g2_nand2b_2 _1865_ (.Y(_1044_),
    .B(_1043_),
    .A_N(_1012_));
 sg13g2_a22oi_1 _1866_ (.Y(_1045_),
    .B1(_1044_),
    .B2(net683),
    .A2(_1041_),
    .A1(net667));
 sg13g2_inv_1 _1867_ (.Y(_0002_),
    .A(_1045_));
 sg13g2_a22oi_1 _1868_ (.Y(_1046_),
    .B1(_1041_),
    .B2(net703),
    .A2(_1012_),
    .A1(net422));
 sg13g2_inv_1 _1869_ (.Y(_0005_),
    .A(_1046_));
 sg13g2_a22oi_1 _1870_ (.Y(_1047_),
    .B1(_1044_),
    .B2(net674),
    .A2(_1041_),
    .A1(\levenshtein_ctrl.state[2] ));
 sg13g2_inv_1 _1871_ (.Y(_0006_),
    .A(net675));
 sg13g2_and3_1 _1872_ (.X(_1048_),
    .A(\arbiter.wbs1_cyc_i ),
    .B(_1013_),
    .C(net394));
 sg13g2_a22oi_1 _1873_ (.Y(_1049_),
    .B1(_1048_),
    .B2(net425),
    .A2(_1044_),
    .A1(net667));
 sg13g2_inv_1 _1874_ (.Y(_0004_),
    .A(net668));
 sg13g2_a21oi_1 _1875_ (.A1(\levenshtein_ctrl.symbol_idx[0] ),
    .A2(\levenshtein_ctrl.symbol_idx[1] ),
    .Y(_1050_),
    .B1(_0991_));
 sg13g2_a21oi_1 _1876_ (.A1(_1024_),
    .A2(_1050_),
    .Y(_1051_),
    .B1(_1012_));
 sg13g2_o21ai_1 _1877_ (.B1(_1051_),
    .Y(_1052_),
    .A1(_1014_),
    .A2(_1022_));
 sg13g2_nand2_1 _1878_ (.Y(_1053_),
    .A(\levenshtein_ctrl.state[6] ),
    .B(_1015_));
 sg13g2_nor2_2 _1879_ (.A(_0955_),
    .B(_1042_),
    .Y(_1054_));
 sg13g2_a21oi_1 _1880_ (.A1(net570),
    .A2(_1052_),
    .Y(_1055_),
    .B1(_1054_));
 sg13g2_o21ai_1 _1881_ (.B1(_1055_),
    .Y(_0001_),
    .A1(_1029_),
    .A2(net689));
 sg13g2_nand2b_1 _1882_ (.Y(_1056_),
    .B(net437),
    .A_N(\spi.ss_n ));
 sg13g2_nor2b_2 _1883_ (.A(\spi.last_sck ),
    .B_N(net264),
    .Y(_1057_));
 sg13g2_nand2b_2 _1884_ (.Y(_1058_),
    .B(net264),
    .A_N(\spi.last_sck ));
 sg13g2_and3_1 _1885_ (.X(_1059_),
    .A(net299),
    .B(\spi.counter[0] ),
    .C(_1057_));
 sg13g2_and2_1 _1886_ (.A(net317),
    .B(_1059_),
    .X(_1060_));
 sg13g2_and2_1 _1887_ (.A(net450),
    .B(_1060_),
    .X(_1061_));
 sg13g2_and2_1 _1888_ (.A(net483),
    .B(_1061_),
    .X(_1062_));
 sg13g2_nand2_1 _1889_ (.Y(_1063_),
    .A(\spi.state[0] ),
    .B(_1062_));
 sg13g2_a21o_1 _1890_ (.A2(\arbiter.wbm_ack_i ),
    .A1(net404),
    .B1(net370),
    .X(_1064_));
 sg13g2_o21ai_1 _1891_ (.B1(_1064_),
    .Y(_1065_),
    .A1(ctrl_slave_ack),
    .A2(_1000_));
 sg13g2_nand2_1 _1892_ (.Y(_1066_),
    .A(net671),
    .B(_1065_));
 sg13g2_a21oi_1 _1893_ (.A1(_1063_),
    .A2(_1066_),
    .Y(_0009_),
    .B1(net393));
 sg13g2_nand2b_1 _1894_ (.Y(_1067_),
    .B(net694),
    .A_N(_1062_));
 sg13g2_nand2b_1 _1895_ (.Y(_0008_),
    .B(_1067_),
    .A_N(net393));
 sg13g2_a22oi_1 _1896_ (.Y(_1068_),
    .B1(_1048_),
    .B2(net715),
    .A2(_1044_),
    .A1(net703));
 sg13g2_inv_1 _1897_ (.Y(_0007_),
    .A(net716));
 sg13g2_nor2_1 _1898_ (.A(net292),
    .B(_1058_),
    .Y(_1069_));
 sg13g2_nor2_1 _1899_ (.A(\spi.counter[0] ),
    .B(_1057_),
    .Y(_1070_));
 sg13g2_nor3_1 _1900_ (.A(_1056_),
    .B(net293),
    .C(_1070_),
    .Y(_0068_));
 sg13g2_a21oi_1 _1901_ (.A1(\spi.counter[0] ),
    .A2(_1057_),
    .Y(_1071_),
    .B1(net299));
 sg13g2_nor3_1 _1902_ (.A(_1056_),
    .B(_1059_),
    .C(net300),
    .Y(_0069_));
 sg13g2_nor2_1 _1903_ (.A(net317),
    .B(_1059_),
    .Y(_1072_));
 sg13g2_nor3_1 _1904_ (.A(_1056_),
    .B(_1060_),
    .C(net318),
    .Y(_0070_));
 sg13g2_nor2_1 _1905_ (.A(net450),
    .B(_1060_),
    .Y(_1073_));
 sg13g2_nor3_1 _1906_ (.A(net393),
    .B(_1061_),
    .C(_1073_),
    .Y(_0071_));
 sg13g2_nor2_1 _1907_ (.A(net483),
    .B(_1061_),
    .Y(_1074_));
 sg13g2_nor3_1 _1908_ (.A(net393),
    .B(_1062_),
    .C(_1074_),
    .Y(_0072_));
 sg13g2_nor2_1 _1909_ (.A(net416),
    .B(_1040_),
    .Y(_1075_));
 sg13g2_or2_1 _1910_ (.X(_1076_),
    .B(_1040_),
    .A(net416));
 sg13g2_nand3_1 _1911_ (.B(_1034_),
    .C(net344),
    .A(\levenshtein_ctrl.symbol_idx[0] ),
    .Y(_1077_));
 sg13g2_nand2_1 _1912_ (.Y(_1078_),
    .A(net704),
    .B(_1033_));
 sg13g2_nand3_1 _1913_ (.B(_1077_),
    .C(_1078_),
    .A(net435),
    .Y(_1079_));
 sg13g2_o21ai_1 _1914_ (.B1(net705),
    .Y(_1080_),
    .A1(\levenshtein_ctrl.symbol_idx[0] ),
    .A2(net435));
 sg13g2_inv_1 _1915_ (.Y(_0073_),
    .A(net706));
 sg13g2_nand3_1 _1916_ (.B(\levenshtein_ctrl.symbol_idx[0] ),
    .C(net397),
    .A(net423),
    .Y(_1081_));
 sg13g2_nor2_2 _1917_ (.A(net431),
    .B(net346),
    .Y(_1082_));
 sg13g2_nand4_1 _1918_ (.B(_1001_),
    .C(_1004_),
    .A(\arbiter.wbs0_we_i ),
    .Y(_1083_),
    .D(_1005_));
 sg13g2_nand2_1 _1919_ (.Y(_1084_),
    .A(net617),
    .B(net359));
 sg13g2_xor2_1 _1920_ (.B(_1084_),
    .A(_1081_),
    .X(_0074_));
 sg13g2_nor2_1 _1921_ (.A(\spi.state[0] ),
    .B(\spi.state[2] ),
    .Y(_1085_));
 sg13g2_nor4_1 _1922_ (.A(\arbiter.wbs0_adr_i[0] ),
    .B(\spi.state[0] ),
    .C(\spi.state[2] ),
    .D(_1058_),
    .Y(_1086_));
 sg13g2_a21oi_1 _1923_ (.A1(_1057_),
    .A2(_1085_),
    .Y(_1087_),
    .B1(net287));
 sg13g2_nor3_1 _1924_ (.A(net393),
    .B(_1086_),
    .C(net288),
    .Y(_0075_));
 sg13g2_or2_1 _1925_ (.X(_1088_),
    .B(\spi.state[0] ),
    .A(net641));
 sg13g2_a22oi_1 _1926_ (.Y(_1089_),
    .B1(_1088_),
    .B2(_1063_),
    .A2(_1065_),
    .A1(_0935_));
 sg13g2_nor2_1 _1927_ (.A(\intercon.wbs_cyc_i ),
    .B(_1089_),
    .Y(_1090_));
 sg13g2_or2_1 _1928_ (.X(_1091_),
    .B(_1090_),
    .A(net393));
 sg13g2_a21oi_1 _1929_ (.A1(_0935_),
    .A2(_1089_),
    .Y(_0076_),
    .B1(_1091_));
 sg13g2_nor2_1 _1930_ (.A(net727),
    .B(net370),
    .Y(_1092_));
 sg13g2_and4_1 _1931_ (.A(net399),
    .B(\arbiter.cyc ),
    .C(\arbiter.wbs1_cyc_i ),
    .D(net436),
    .X(_1093_));
 sg13g2_and3_1 _1932_ (.X(_1094_),
    .A(net404),
    .B(net718),
    .C(net436));
 sg13g2_a21oi_1 _1933_ (.A1(_1092_),
    .A2(_1094_),
    .Y(_1095_),
    .B1(_1093_));
 sg13g2_nor2_2 _1934_ (.A(net417),
    .B(net420),
    .Y(_1096_));
 sg13g2_or2_2 _1935_ (.X(_1097_),
    .B(net420),
    .A(net417));
 sg13g2_nor2_1 _1936_ (.A(net406),
    .B(_1097_),
    .Y(_1098_));
 sg13g2_nor3_2 _1937_ (.A(net405),
    .B(\spi_ctrl.bit_counter[3] ),
    .C(_1097_),
    .Y(_1099_));
 sg13g2_nor2_2 _1938_ (.A(net399),
    .B(_0937_),
    .Y(_1100_));
 sg13g2_nand2_2 _1939_ (.Y(_1101_),
    .A(net404),
    .B(\arbiter.wbs0_we_i ));
 sg13g2_nand3_1 _1940_ (.B(_1099_),
    .C(_1100_),
    .A(net634),
    .Y(_1102_));
 sg13g2_nor2b_1 _1941_ (.A(\spi_ctrl.bit_counter[3] ),
    .B_N(net405),
    .Y(_1103_));
 sg13g2_and2_2 _1942_ (.A(\spi_ctrl.bit_counter[1] ),
    .B(net420),
    .X(_1104_));
 sg13g2_nand2_1 _1943_ (.Y(_1105_),
    .A(net417),
    .B(net420));
 sg13g2_nor3_1 _1944_ (.A(_0066_),
    .B(_1100_),
    .C(_1105_),
    .Y(_1106_));
 sg13g2_a21oi_1 _1945_ (.A1(_1103_),
    .A2(_1106_),
    .Y(_1107_),
    .B1(net351));
 sg13g2_nand2_1 _1946_ (.Y(_1108_),
    .A(_1102_),
    .B(_1107_));
 sg13g2_nor2b_1 _1947_ (.A(\levenshtein_ctrl.state[3] ),
    .B_N(_0061_),
    .Y(_1109_));
 sg13g2_nor3_2 _1948_ (.A(\levenshtein_ctrl.state[4] ),
    .B(\levenshtein_ctrl.state[2] ),
    .C(\levenshtein_ctrl.state[6] ),
    .Y(_1110_));
 sg13g2_or3_1 _1949_ (.A(\levenshtein_ctrl.state[4] ),
    .B(\levenshtein_ctrl.state[2] ),
    .C(\levenshtein_ctrl.state[6] ),
    .X(_1111_));
 sg13g2_nor2_1 _1950_ (.A(net425),
    .B(_1111_),
    .Y(_1112_));
 sg13g2_o21ai_1 _1951_ (.B1(_0061_),
    .Y(_1113_),
    .A1(_0955_),
    .A2(\levenshtein_ctrl.state[3] ));
 sg13g2_a22oi_1 _1952_ (.Y(_1114_),
    .B1(_1113_),
    .B2(_0010_),
    .A2(_1112_),
    .A1(_1109_));
 sg13g2_nand2_1 _1953_ (.Y(_1115_),
    .A(net399),
    .B(_1114_));
 sg13g2_nor2_2 _1954_ (.A(net417),
    .B(_0933_),
    .Y(_1116_));
 sg13g2_and4_1 _1955_ (.A(\spi_ctrl.bit_counter[4] ),
    .B(_1101_),
    .C(_1103_),
    .D(_1116_),
    .X(_1117_));
 sg13g2_nand4_1 _1956_ (.B(_0931_),
    .C(_1114_),
    .A(net400),
    .Y(_1118_),
    .D(_1117_));
 sg13g2_nand3_1 _1957_ (.B(_1107_),
    .C(_1118_),
    .A(_1102_),
    .Y(_1119_));
 sg13g2_mux2_1 _1958_ (.A0(net398),
    .A1(_0934_),
    .S(net407),
    .X(_1120_));
 sg13g2_nor2_1 _1959_ (.A(_1119_),
    .B(_1120_),
    .Y(_0077_));
 sg13g2_nor2_2 _1960_ (.A(_1096_),
    .B(_1104_),
    .Y(_1121_));
 sg13g2_nor3_1 _1961_ (.A(_0932_),
    .B(_1096_),
    .C(_1104_),
    .Y(_1122_));
 sg13g2_a21oi_1 _1962_ (.A1(_0932_),
    .A2(net417),
    .Y(_1123_),
    .B1(_1122_));
 sg13g2_nor2_1 _1963_ (.A(_1119_),
    .B(_1123_),
    .Y(_0078_));
 sg13g2_and2_2 _1964_ (.A(net405),
    .B(_1104_),
    .X(_1124_));
 sg13g2_nand2_1 _1965_ (.Y(_1125_),
    .A(net407),
    .B(_1124_));
 sg13g2_nand2_1 _1966_ (.Y(_1126_),
    .A(net405),
    .B(\spi_ctrl.bit_counter[3] ));
 sg13g2_nand2_1 _1967_ (.Y(_1127_),
    .A(\spi_ctrl.bit_counter[3] ),
    .B(_1124_));
 sg13g2_xor2_1 _1968_ (.B(_1125_),
    .A(net736),
    .X(_1128_));
 sg13g2_nor2_1 _1969_ (.A(_1119_),
    .B(_1128_),
    .Y(_0079_));
 sg13g2_nand2_2 _1970_ (.Y(_1129_),
    .A(_0066_),
    .B(_1099_));
 sg13g2_nor3_1 _1971_ (.A(\spi_ctrl.bit_counter[4] ),
    .B(_1101_),
    .C(_1127_),
    .Y(_1130_));
 sg13g2_o21ai_1 _1972_ (.B1(net408),
    .Y(_1131_),
    .A1(_1117_),
    .A2(_1130_));
 sg13g2_inv_1 _1973_ (.Y(_1132_),
    .A(_1131_));
 sg13g2_a22oi_1 _1974_ (.Y(_1133_),
    .B1(_1132_),
    .B2(_1115_),
    .A2(_1129_),
    .A1(net729));
 sg13g2_nand2b_1 _1975_ (.Y(_0080_),
    .B(net730),
    .A_N(net351));
 sg13g2_nor2_1 _1976_ (.A(_1100_),
    .B(_1129_),
    .Y(_1134_));
 sg13g2_a21oi_1 _1977_ (.A1(net749),
    .A2(_1129_),
    .Y(_1135_),
    .B1(_1134_));
 sg13g2_nand2b_1 _1978_ (.Y(_1136_),
    .B(_0932_),
    .A_N(_1135_));
 sg13g2_nor2_1 _1979_ (.A(\spi_ctrl.bit_counter[3] ),
    .B(_1124_),
    .Y(_1137_));
 sg13g2_o21ai_1 _1980_ (.B1(_0964_),
    .Y(_1138_),
    .A1(\spi_ctrl.bit_counter[4] ),
    .A2(_1126_));
 sg13g2_o21ai_1 _1981_ (.B1(_1138_),
    .Y(_1139_),
    .A1(_1096_),
    .A2(_1126_));
 sg13g2_a21oi_2 _1982_ (.B1(_1139_),
    .Y(_1140_),
    .A2(_1137_),
    .A1(_0930_));
 sg13g2_xnor2_1 _1983_ (.Y(_1141_),
    .A(net405),
    .B(_1104_));
 sg13g2_nor2_2 _1984_ (.A(_1098_),
    .B(_1124_),
    .Y(_1142_));
 sg13g2_inv_1 _1985_ (.Y(_1143_),
    .A(_1142_));
 sg13g2_a21oi_2 _1986_ (.B1(_1143_),
    .Y(_1144_),
    .A2(_1121_),
    .A1(net406));
 sg13g2_nor2_2 _1987_ (.A(\levenshtein_ctrl.state[7] ),
    .B(\levenshtein_ctrl.state[3] ),
    .Y(_1145_));
 sg13g2_or2_1 _1988_ (.X(_1146_),
    .B(\levenshtein_ctrl.state[3] ),
    .A(\levenshtein_ctrl.state[7] ));
 sg13g2_a21oi_1 _1989_ (.A1(net424),
    .A2(\levenshtein_ctrl.dict_address[6] ),
    .Y(_1147_),
    .B1(net389));
 sg13g2_nand2_1 _1990_ (.Y(_1148_),
    .A(net417),
    .B(net398));
 sg13g2_a21oi_1 _1991_ (.A1(net424),
    .A2(\levenshtein_ctrl.dict_address[10] ),
    .Y(_1149_),
    .B1(net389));
 sg13g2_a21oi_2 _1992_ (.B1(_1148_),
    .Y(_1150_),
    .A2(_0012_),
    .A1(net402));
 sg13g2_a21oi_1 _1993_ (.A1(_0048_),
    .A2(net391),
    .Y(_1151_),
    .B1(net385));
 sg13g2_nor2b_1 _1994_ (.A(_1147_),
    .B_N(_1151_),
    .Y(_1152_));
 sg13g2_o21ai_1 _1995_ (.B1(net399),
    .Y(_1153_),
    .A1(_0021_),
    .A2(_1145_));
 sg13g2_o21ai_1 _1996_ (.B1(_1150_),
    .Y(_1154_),
    .A1(_1152_),
    .A2(_1153_));
 sg13g2_a21oi_1 _1997_ (.A1(_0045_),
    .A2(net389),
    .Y(_1155_),
    .B1(_1149_));
 sg13g2_a21oi_1 _1998_ (.A1(_1109_),
    .A2(_1155_),
    .Y(_1156_),
    .B1(net401));
 sg13g2_o21ai_1 _1999_ (.B1(_1116_),
    .Y(_1157_),
    .A1(net400),
    .A2(\arbiter.wbs0_adr_i[12] ));
 sg13g2_o21ai_1 _2000_ (.B1(_1154_),
    .Y(_1158_),
    .A1(_1156_),
    .A2(_1157_));
 sg13g2_a21oi_1 _2001_ (.A1(net424),
    .A2(\levenshtein_ctrl.dict_address[2] ),
    .Y(_1159_),
    .B1(net390));
 sg13g2_a21oi_1 _2002_ (.A1(_0052_),
    .A2(net390),
    .Y(_1160_),
    .B1(_1159_));
 sg13g2_a21oi_1 _2003_ (.A1(_0025_),
    .A2(_1146_),
    .Y(_1161_),
    .B1(net398));
 sg13g2_o21ai_1 _2004_ (.B1(_1161_),
    .Y(_1162_),
    .A1(_1146_),
    .A2(_1160_));
 sg13g2_o21ai_1 _2005_ (.B1(_0064_),
    .Y(_1163_),
    .A1(_0954_),
    .A2(\levenshtein_ctrl.state[2] ));
 sg13g2_a21oi_1 _2006_ (.A1(_0062_),
    .A2(_1163_),
    .Y(_1164_),
    .B1(\levenshtein_ctrl.state[7] ));
 sg13g2_o21ai_1 _2007_ (.B1(net399),
    .Y(_1165_),
    .A1(net421),
    .A2(_1164_));
 sg13g2_nor2b_1 _2008_ (.A(_1165_),
    .B_N(_1162_),
    .Y(_1166_));
 sg13g2_o21ai_1 _2009_ (.B1(net403),
    .Y(_1167_),
    .A1(net398),
    .A2(_0016_));
 sg13g2_a21oi_1 _2010_ (.A1(net398),
    .A2(\arbiter.wbs0_adr_i[0] ),
    .Y(_1168_),
    .B1(_1167_));
 sg13g2_nor3_1 _2011_ (.A(_1121_),
    .B(_1166_),
    .C(_1168_),
    .Y(_1169_));
 sg13g2_o21ai_1 _2012_ (.B1(_1144_),
    .Y(_1170_),
    .A1(_1158_),
    .A2(_1169_));
 sg13g2_o21ai_1 _2013_ (.B1(_1109_),
    .Y(_1171_),
    .A1(net424),
    .A2(net388));
 sg13g2_nor2_2 _2014_ (.A(net403),
    .B(_1171_),
    .Y(_1172_));
 sg13g2_nand2_1 _2015_ (.Y(_1173_),
    .A(_0037_),
    .B(net387));
 sg13g2_o21ai_1 _2016_ (.B1(_1173_),
    .Y(_1174_),
    .A1(\levenshtein_ctrl.dict_address[18] ),
    .A2(net386));
 sg13g2_a21oi_1 _2017_ (.A1(_0041_),
    .A2(net387),
    .Y(_1175_),
    .B1(net418));
 sg13g2_o21ai_1 _2018_ (.B1(_1175_),
    .Y(_1176_),
    .A1(\levenshtein_ctrl.dict_address[14] ),
    .A2(net387));
 sg13g2_o21ai_1 _2019_ (.B1(_1176_),
    .Y(_1177_),
    .A1(net398),
    .A2(_1174_));
 sg13g2_mux2_1 _2020_ (.A0(\arbiter.wbs0_adr_i[16] ),
    .A1(\arbiter.wbs0_adr_i[20] ),
    .S(net419),
    .X(_1178_));
 sg13g2_a22oi_1 _2021_ (.Y(_1179_),
    .B1(_1178_),
    .B2(net402),
    .A2(_1177_),
    .A1(_1172_));
 sg13g2_o21ai_1 _2022_ (.B1(_1170_),
    .Y(_1180_),
    .A1(_1142_),
    .A2(_1179_));
 sg13g2_nand4_1 _2023_ (.B(\spi_ctrl.bit_counter[3] ),
    .C(_0066_),
    .A(net406),
    .Y(_1181_),
    .D(_1116_));
 sg13g2_nor3_1 _2024_ (.A(_0964_),
    .B(_1126_),
    .C(_1148_),
    .Y(_1182_));
 sg13g2_nand2_1 _2025_ (.Y(_1183_),
    .A(\arbiter.wbs0_dat_i[0] ),
    .B(net367));
 sg13g2_a21oi_1 _2026_ (.A1(_1181_),
    .A2(_1183_),
    .Y(_1184_),
    .B1(_1101_));
 sg13g2_nor2_1 _2027_ (.A(\spi_ctrl.bit_counter[4] ),
    .B(_1148_),
    .Y(_1185_));
 sg13g2_a22oi_1 _2028_ (.Y(_1186_),
    .B1(_1185_),
    .B2(_1103_),
    .A2(_1137_),
    .A1(_0066_));
 sg13g2_nand2b_1 _2029_ (.Y(_1187_),
    .B(_1186_),
    .A_N(_1135_));
 sg13g2_nand2_1 _2030_ (.Y(_1188_),
    .A(_1100_),
    .B(_1141_));
 sg13g2_o21ai_1 _2031_ (.B1(_1101_),
    .Y(_1189_),
    .A1(net405),
    .A2(net420));
 sg13g2_nand3_1 _2032_ (.B(_1188_),
    .C(_1189_),
    .A(_1121_),
    .Y(_1190_));
 sg13g2_o21ai_1 _2033_ (.B1(_1188_),
    .Y(_1191_),
    .A1(_0934_),
    .A2(_1141_));
 sg13g2_nand2b_1 _2034_ (.Y(_1192_),
    .B(_1191_),
    .A_N(_1121_));
 sg13g2_nand4_1 _2035_ (.B(_1137_),
    .C(_1190_),
    .A(_0066_),
    .Y(_1193_),
    .D(_1192_));
 sg13g2_a21oi_1 _2036_ (.A1(_1187_),
    .A2(_1193_),
    .Y(_1194_),
    .B1(_1140_));
 sg13g2_a21o_1 _2037_ (.A2(_1180_),
    .A1(_1140_),
    .B1(_1194_),
    .X(_1195_));
 sg13g2_nor2_1 _2038_ (.A(\arbiter.wbs0_dat_i[4] ),
    .B(_1181_),
    .Y(_1196_));
 sg13g2_a21oi_1 _2039_ (.A1(\arbiter.wbs0_dat_i[0] ),
    .A2(net367),
    .Y(_1197_),
    .B1(_1101_));
 sg13g2_o21ai_1 _2040_ (.B1(_1197_),
    .Y(_1198_),
    .A1(net367),
    .A2(_1196_));
 sg13g2_and2_1 _2041_ (.A(net407),
    .B(_1198_),
    .X(_1199_));
 sg13g2_o21ai_1 _2042_ (.B1(_1199_),
    .Y(_1200_),
    .A1(_1184_),
    .A2(_1195_));
 sg13g2_a21oi_1 _2043_ (.A1(_1136_),
    .A2(_1200_),
    .Y(_0081_),
    .B1(net351));
 sg13g2_nor2_1 _2044_ (.A(net718),
    .B(net431),
    .Y(_1201_));
 sg13g2_o21ai_1 _2045_ (.B1(_1201_),
    .Y(_1202_),
    .A1(\arbiter.wbs1_cyc_i ),
    .A2(_1092_));
 sg13g2_nand2_1 _2046_ (.Y(_0082_),
    .A(net352),
    .B(net719));
 sg13g2_nor3_2 _2047_ (.A(_0936_),
    .B(\arbiter.wbs0_adr_i[1] ),
    .C(_0967_),
    .Y(_1203_));
 sg13g2_nand3_1 _2048_ (.B(_1009_),
    .C(_1203_),
    .A(net436),
    .Y(_1204_));
 sg13g2_mux2_1 _2049_ (.A0(\arbiter.wbs0_dat_i[0] ),
    .A1(net686),
    .S(_1204_),
    .X(_0083_));
 sg13g2_mux2_1 _2050_ (.A0(\arbiter.wbs0_dat_i[1] ),
    .A1(net619),
    .S(_1204_),
    .X(_0084_));
 sg13g2_o21ai_1 _2051_ (.B1(_1053_),
    .Y(_1205_),
    .A1(\arbiter.wbs1_cyc_i ),
    .A2(net425));
 sg13g2_nand2_1 _2052_ (.Y(_1206_),
    .A(\levenshtein_ctrl.state[3] ),
    .B(net695));
 sg13g2_a221oi_1 _2053_ (.B2(_1206_),
    .C1(_0991_),
    .B1(_1205_),
    .A1(\levenshtein_ctrl.state[7] ),
    .Y(_1207_),
    .A2(net394));
 sg13g2_a21o_1 _2054_ (.A2(net395),
    .A1(\arbiter.wbs1_cyc_i ),
    .B1(_1207_),
    .X(_0085_));
 sg13g2_nor2_1 _2055_ (.A(net396),
    .B(_1039_),
    .Y(_1208_));
 sg13g2_nor2_1 _2056_ (.A(net725),
    .B(_1040_),
    .Y(_1209_));
 sg13g2_nor2_1 _2057_ (.A(_1022_),
    .B(_1034_),
    .Y(_1210_));
 sg13g2_nor3_1 _2058_ (.A(_1208_),
    .B(_1209_),
    .C(_1210_),
    .Y(_0087_));
 sg13g2_nor2b_1 _2059_ (.A(\arbiter.wbs0_adr_i[0] ),
    .B_N(\arbiter.wbs0_adr_i[1] ),
    .Y(_1211_));
 sg13g2_and2_1 _2060_ (.A(_0018_),
    .B(_1211_),
    .X(_1212_));
 sg13g2_nand3_1 _2061_ (.B(_1009_),
    .C(_1212_),
    .A(net436),
    .Y(_1213_));
 sg13g2_mux2_1 _2062_ (.A0(net725),
    .A1(\levenshtein_ctrl.word_length_reg[0] ),
    .S(_1213_),
    .X(_0088_));
 sg13g2_mux2_1 _2063_ (.A0(net662),
    .A1(net414),
    .S(_1213_),
    .X(_0089_));
 sg13g2_nor2_1 _2064_ (.A(net628),
    .B(_1213_),
    .Y(_1214_));
 sg13g2_a21oi_1 _2065_ (.A1(_0971_),
    .A2(_1213_),
    .Y(_0090_),
    .B1(_1214_));
 sg13g2_mux2_1 _2066_ (.A0(net650),
    .A1(net411),
    .S(_1213_),
    .X(_0091_));
 sg13g2_nor2b_1 _2067_ (.A(_1054_),
    .B_N(\levenshtein_ctrl.dict_address[0] ),
    .Y(_1215_));
 sg13g2_a21oi_1 _2068_ (.A1(net297),
    .A2(_1054_),
    .Y(_1216_),
    .B1(_1215_));
 sg13g2_nor2_1 _2069_ (.A(_1082_),
    .B(net298),
    .Y(_0092_));
 sg13g2_a22oi_1 _2070_ (.Y(_1217_),
    .B1(net359),
    .B2(net512),
    .A2(_1054_),
    .A1(\levenshtein_ctrl.dict_address[0] ));
 sg13g2_nand2_1 _2071_ (.Y(_1218_),
    .A(\levenshtein_ctrl.dict_address[0] ),
    .B(net512));
 sg13g2_nand3_1 _2072_ (.B(net512),
    .C(_1054_),
    .A(\levenshtein_ctrl.dict_address[0] ),
    .Y(_1219_));
 sg13g2_nor2b_1 _2073_ (.A(net513),
    .B_N(_1219_),
    .Y(_0093_));
 sg13g2_nand2_1 _2074_ (.Y(_1220_),
    .A(net527),
    .B(net358));
 sg13g2_xor2_1 _2075_ (.B(_1220_),
    .A(_1219_),
    .X(_0094_));
 sg13g2_nor2_1 _2076_ (.A(net455),
    .B(_1219_),
    .Y(_1221_));
 sg13g2_nand2_1 _2077_ (.Y(_1222_),
    .A(\levenshtein_ctrl.dict_address[3] ),
    .B(net358));
 sg13g2_xnor2_1 _2078_ (.Y(_0095_),
    .A(net456),
    .B(_1222_));
 sg13g2_nand2_1 _2079_ (.Y(_1223_),
    .A(net527),
    .B(\levenshtein_ctrl.dict_address[3] ));
 sg13g2_nor4_2 _2080_ (.A(_0955_),
    .B(_1042_),
    .C(_1218_),
    .Y(_1224_),
    .D(_1223_));
 sg13g2_nand2_1 _2081_ (.Y(_1225_),
    .A(net510),
    .B(net358));
 sg13g2_xnor2_1 _2082_ (.Y(_0096_),
    .A(_1224_),
    .B(_1225_));
 sg13g2_nor2b_1 _2083_ (.A(net500),
    .B_N(_1224_),
    .Y(_1226_));
 sg13g2_nand2_1 _2084_ (.Y(_1227_),
    .A(\levenshtein_ctrl.dict_address[5] ),
    .B(net358));
 sg13g2_xnor2_1 _2085_ (.Y(_0097_),
    .A(_1226_),
    .B(_1227_));
 sg13g2_nand2_1 _2086_ (.Y(_1228_),
    .A(net583),
    .B(net358));
 sg13g2_nand3_1 _2087_ (.B(\levenshtein_ctrl.dict_address[5] ),
    .C(_1224_),
    .A(net510),
    .Y(_1229_));
 sg13g2_xor2_1 _2088_ (.B(_1229_),
    .A(_1228_),
    .X(_0098_));
 sg13g2_nand2_1 _2089_ (.Y(_1230_),
    .A(\levenshtein_ctrl.dict_address[7] ),
    .B(net358));
 sg13g2_nor2_1 _2090_ (.A(net621),
    .B(_1229_),
    .Y(_1231_));
 sg13g2_xnor2_1 _2091_ (.Y(_0099_),
    .A(_1230_),
    .B(net622));
 sg13g2_nor3_2 _2092_ (.A(_0965_),
    .B(_0966_),
    .C(_1229_),
    .Y(_1232_));
 sg13g2_nor3_1 _2093_ (.A(net466),
    .B(_1082_),
    .C(_1232_),
    .Y(_1233_));
 sg13g2_a21oi_1 _2094_ (.A1(net466),
    .A2(_1232_),
    .Y(_0100_),
    .B1(_1233_));
 sg13g2_nand2_1 _2095_ (.Y(_1234_),
    .A(\levenshtein_ctrl.dict_address[9] ),
    .B(net356));
 sg13g2_nor2b_1 _2096_ (.A(net495),
    .B_N(_1232_),
    .Y(_1235_));
 sg13g2_xnor2_1 _2097_ (.Y(_0101_),
    .A(_1234_),
    .B(net496));
 sg13g2_nand2_1 _2098_ (.Y(_1236_),
    .A(net624),
    .B(net356));
 sg13g2_and3_1 _2099_ (.X(_1237_),
    .A(net466),
    .B(\levenshtein_ctrl.dict_address[9] ),
    .C(_1232_));
 sg13g2_xnor2_1 _2100_ (.Y(_0102_),
    .A(_1236_),
    .B(_1237_));
 sg13g2_nand2_1 _2101_ (.Y(_1238_),
    .A(\levenshtein_ctrl.dict_address[11] ),
    .B(net356));
 sg13g2_nand2b_1 _2102_ (.Y(_1239_),
    .B(_1237_),
    .A_N(net461));
 sg13g2_xor2_1 _2103_ (.B(net462),
    .A(_1238_),
    .X(_0103_));
 sg13g2_nand2_1 _2104_ (.Y(_1240_),
    .A(net656),
    .B(net356));
 sg13g2_nand3_1 _2105_ (.B(\levenshtein_ctrl.dict_address[11] ),
    .C(_1237_),
    .A(net624),
    .Y(_1241_));
 sg13g2_xor2_1 _2106_ (.B(_1241_),
    .A(_1240_),
    .X(_0104_));
 sg13g2_nand2_1 _2107_ (.Y(_1242_),
    .A(\levenshtein_ctrl.dict_address[13] ),
    .B(net356));
 sg13g2_nor2_1 _2108_ (.A(net543),
    .B(_1241_),
    .Y(_1243_));
 sg13g2_xnor2_1 _2109_ (.Y(_0105_),
    .A(_1242_),
    .B(net544));
 sg13g2_nand2_1 _2110_ (.Y(_1244_),
    .A(net608),
    .B(net357));
 sg13g2_nor3_2 _2111_ (.A(_0970_),
    .B(_1240_),
    .C(_1241_),
    .Y(_1245_));
 sg13g2_and2_1 _2112_ (.A(\levenshtein_ctrl.dict_address[14] ),
    .B(_1245_),
    .X(_1246_));
 sg13g2_xnor2_1 _2113_ (.Y(_0106_),
    .A(_1244_),
    .B(_1245_));
 sg13g2_nand2_1 _2114_ (.Y(_1247_),
    .A(\levenshtein_ctrl.dict_address[15] ),
    .B(net357));
 sg13g2_nor2b_1 _2115_ (.A(net447),
    .B_N(_1245_),
    .Y(_1248_));
 sg13g2_xnor2_1 _2116_ (.Y(_0107_),
    .A(_1247_),
    .B(net448));
 sg13g2_nand2_1 _2117_ (.Y(_1249_),
    .A(net593),
    .B(net357));
 sg13g2_nand2_1 _2118_ (.Y(_1250_),
    .A(\levenshtein_ctrl.dict_address[15] ),
    .B(_1246_));
 sg13g2_xor2_1 _2119_ (.B(_1250_),
    .A(_1249_),
    .X(_0108_));
 sg13g2_nand2_1 _2120_ (.Y(_1251_),
    .A(\levenshtein_ctrl.dict_address[17] ),
    .B(net356));
 sg13g2_nor2_1 _2121_ (.A(net535),
    .B(_1250_),
    .Y(_1252_));
 sg13g2_xnor2_1 _2122_ (.Y(_0109_),
    .A(_1251_),
    .B(net536));
 sg13g2_nand2_1 _2123_ (.Y(_1253_),
    .A(net563),
    .B(net356));
 sg13g2_nand4_1 _2124_ (.B(\levenshtein_ctrl.dict_address[16] ),
    .C(\levenshtein_ctrl.dict_address[17] ),
    .A(\levenshtein_ctrl.dict_address[15] ),
    .Y(_1254_),
    .D(_1246_));
 sg13g2_xor2_1 _2125_ (.B(_1254_),
    .A(_1253_),
    .X(_0110_));
 sg13g2_nand2_1 _2126_ (.Y(_1255_),
    .A(\levenshtein_ctrl.dict_address[19] ),
    .B(net356));
 sg13g2_nor2_1 _2127_ (.A(net546),
    .B(_1254_),
    .Y(_1256_));
 sg13g2_xnor2_1 _2128_ (.Y(_0111_),
    .A(_1255_),
    .B(net547));
 sg13g2_nand2_1 _2129_ (.Y(_1257_),
    .A(net553),
    .B(net357));
 sg13g2_nand2_1 _2130_ (.Y(_1258_),
    .A(\levenshtein_ctrl.dict_address[18] ),
    .B(\levenshtein_ctrl.dict_address[19] ));
 sg13g2_nor2_1 _2131_ (.A(_1254_),
    .B(_1258_),
    .Y(_1259_));
 sg13g2_xnor2_1 _2132_ (.Y(_0112_),
    .A(_1257_),
    .B(_1259_));
 sg13g2_and3_2 _2133_ (.X(_1260_),
    .A(\levenshtein_ctrl.state[7] ),
    .B(_1013_),
    .C(net394));
 sg13g2_mux2_1 _2134_ (.A0(net646),
    .A1(\arbiter.wbm_dat_i[0] ),
    .S(net384),
    .X(_0113_));
 sg13g2_mux2_1 _2135_ (.A0(net517),
    .A1(net761),
    .S(net384),
    .X(_0114_));
 sg13g2_mux2_1 _2136_ (.A0(net645),
    .A1(\arbiter.wbm_dat_i[2] ),
    .S(net384),
    .X(_0115_));
 sg13g2_nor2_1 _2137_ (.A(net508),
    .B(net384),
    .Y(_1261_));
 sg13g2_a21oi_1 _2138_ (.A1(_0963_),
    .A2(net384),
    .Y(_0116_),
    .B1(_1261_));
 sg13g2_mux2_1 _2139_ (.A0(net717),
    .A1(\arbiter.wbm_dat_i[4] ),
    .S(_1260_),
    .X(_0117_));
 sg13g2_mux2_1 _2140_ (.A0(net615),
    .A1(\arbiter.wbm_dat_i[5] ),
    .S(net384),
    .X(_0118_));
 sg13g2_mux2_1 _2141_ (.A0(net680),
    .A1(\arbiter.wbm_dat_i[6] ),
    .S(net384),
    .X(_0119_));
 sg13g2_mux2_1 _2142_ (.A0(net643),
    .A1(\arbiter.wbm_dat_i[7] ),
    .S(net384),
    .X(_0120_));
 sg13g2_nand2_1 _2143_ (.Y(_1262_),
    .A(net431),
    .B(\levenshtein_ctrl.vp[0] ));
 sg13g2_nand2_1 _2144_ (.Y(_1263_),
    .A(net416),
    .B(_1026_));
 sg13g2_and3_1 _2145_ (.X(_1264_),
    .A(_0034_),
    .B(net346),
    .C(_1263_));
 sg13g2_a21oi_1 _2146_ (.A1(net436),
    .A2(net468),
    .Y(_1265_),
    .B1(net395));
 sg13g2_o21ai_1 _2147_ (.B1(_1262_),
    .Y(_0121_),
    .A1(_1264_),
    .A2(_1265_));
 sg13g2_nor2_1 _2148_ (.A(\levenshtein_ctrl.vp[1] ),
    .B(net348),
    .Y(_1266_));
 sg13g2_nor2_2 _2149_ (.A(net415),
    .B(\levenshtein_ctrl.word_length_reg[0] ),
    .Y(_1267_));
 sg13g2_or2_2 _2150_ (.X(_1268_),
    .B(\levenshtein_ctrl.word_length_reg[0] ),
    .A(net414));
 sg13g2_nor2_2 _2151_ (.A(net412),
    .B(net410),
    .Y(_1269_));
 sg13g2_or2_2 _2152_ (.X(_1270_),
    .B(net410),
    .A(net413));
 sg13g2_nor2_1 _2153_ (.A(net412),
    .B(_1268_),
    .Y(_1271_));
 sg13g2_nor2_2 _2154_ (.A(_1268_),
    .B(_1270_),
    .Y(_1272_));
 sg13g2_a21oi_1 _2155_ (.A1(net348),
    .A2(_1272_),
    .Y(_1273_),
    .B1(_1266_));
 sg13g2_nand2b_1 _2156_ (.Y(_1274_),
    .B(_1026_),
    .A_N(_1272_));
 sg13g2_a21oi_1 _2157_ (.A1(_1027_),
    .A2(_1273_),
    .Y(_1275_),
    .B1(net688));
 sg13g2_a21o_1 _2158_ (.A2(\levenshtein_ctrl.pm[0] ),
    .A1(\levenshtein_ctrl.vp[0] ),
    .B1(\levenshtein_ctrl.pm[1] ),
    .X(_1276_));
 sg13g2_nand2b_2 _2159_ (.Y(_1277_),
    .B(_0973_),
    .A_N(_1276_));
 sg13g2_o21ai_1 _2160_ (.B1(_0032_),
    .Y(_1278_),
    .A1(\levenshtein_ctrl.vp[0] ),
    .A2(\levenshtein_ctrl.pm[0] ));
 sg13g2_nor2_1 _2161_ (.A(_1277_),
    .B(_1278_),
    .Y(_1279_));
 sg13g2_nand2b_1 _2162_ (.Y(_1280_),
    .B(_0032_),
    .A_N(\levenshtein_ctrl.pm[0] ));
 sg13g2_a21oi_1 _2163_ (.A1(\levenshtein_ctrl.vp[0] ),
    .A2(_1280_),
    .Y(_1281_),
    .B1(_1279_));
 sg13g2_a221oi_1 _2164_ (.B2(net422),
    .C1(_0991_),
    .B1(_1281_),
    .A1(_1274_),
    .Y(_1282_),
    .A2(_1275_));
 sg13g2_a221oi_1 _2165_ (.B2(_1273_),
    .C1(_1282_),
    .B1(net395),
    .A1(net430),
    .Y(_1283_),
    .A2(net747));
 sg13g2_inv_1 _2166_ (.Y(_0122_),
    .A(_1283_));
 sg13g2_nor2_2 _2167_ (.A(net422),
    .B(_0991_),
    .Y(_1284_));
 sg13g2_nand2b_2 _2168_ (.Y(_1285_),
    .B(net397),
    .A_N(net422));
 sg13g2_a21oi_2 _2169_ (.B1(net395),
    .Y(_1286_),
    .A2(_1284_),
    .A1(_1027_));
 sg13g2_o21ai_1 _2170_ (.B1(_1006_),
    .Y(_1287_),
    .A1(_1026_),
    .A2(_1285_));
 sg13g2_nor2_1 _2171_ (.A(net414),
    .B(_1270_),
    .Y(_1288_));
 sg13g2_a21oi_1 _2172_ (.A1(net348),
    .A2(_1288_),
    .Y(_1289_),
    .B1(_1286_));
 sg13g2_o21ai_1 _2173_ (.B1(_1289_),
    .Y(_1290_),
    .A1(net734),
    .A2(net348));
 sg13g2_and2_1 _2174_ (.A(net422),
    .B(net396),
    .X(_1291_));
 sg13g2_nand2_2 _2175_ (.Y(_1292_),
    .A(net422),
    .B(net396));
 sg13g2_nand2_1 _2176_ (.Y(_1293_),
    .A(\levenshtein_ctrl.vp[1] ),
    .B(_1277_));
 sg13g2_a21oi_2 _2177_ (.B1(\levenshtein_ctrl.pm[2] ),
    .Y(_1294_),
    .A2(_1276_),
    .A1(\levenshtein_ctrl.vp[1] ));
 sg13g2_nand2b_2 _2178_ (.Y(_1295_),
    .B(_1294_),
    .A_N(net441));
 sg13g2_o21ai_1 _2179_ (.B1(_0973_),
    .Y(_1296_),
    .A1(\levenshtein_ctrl.vp[1] ),
    .A2(_1276_));
 sg13g2_o21ai_1 _2180_ (.B1(_1293_),
    .Y(_1297_),
    .A1(_1295_),
    .A2(_1296_));
 sg13g2_nor2_1 _2181_ (.A(_1027_),
    .B(_1285_),
    .Y(_1298_));
 sg13g2_nand2b_1 _2182_ (.Y(_1299_),
    .B(net350),
    .A_N(_1288_));
 sg13g2_a22oi_1 _2183_ (.Y(_1300_),
    .B1(net383),
    .B2(_1297_),
    .A2(net734),
    .A1(net431));
 sg13g2_nand3_1 _2184_ (.B(_1299_),
    .C(_1300_),
    .A(_1290_),
    .Y(_0123_));
 sg13g2_nand2_2 _2185_ (.Y(_1301_),
    .A(net415),
    .B(\levenshtein_ctrl.word_length_reg[0] ));
 sg13g2_nand2_1 _2186_ (.Y(_1302_),
    .A(_0971_),
    .B(_1301_));
 sg13g2_nand2_1 _2187_ (.Y(_1303_),
    .A(_1269_),
    .B(_1301_));
 sg13g2_nor2_1 _2188_ (.A(net345),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_o21ai_1 _2189_ (.B1(net366),
    .Y(_1305_),
    .A1(net745),
    .A2(net348));
 sg13g2_or2_2 _2190_ (.X(_1306_),
    .B(\levenshtein_ctrl.pm[3] ),
    .A(\levenshtein_ctrl.vp[2] ));
 sg13g2_or2_1 _2191_ (.X(_1307_),
    .B(\levenshtein_ctrl.pm[3] ),
    .A(\levenshtein_ctrl.pm[2] ));
 sg13g2_a21o_2 _2192_ (.A2(_1276_),
    .A1(\levenshtein_ctrl.vp[1] ),
    .B1(_1307_),
    .X(_1308_));
 sg13g2_a21oi_1 _2193_ (.A1(_1306_),
    .A2(_1308_),
    .Y(_1309_),
    .B1(net676));
 sg13g2_a21o_1 _2194_ (.A2(_1308_),
    .A1(_1306_),
    .B1(\levenshtein_ctrl.vn[3] ),
    .X(_1310_));
 sg13g2_a21oi_2 _2195_ (.B1(net441),
    .Y(_1311_),
    .A2(_1294_),
    .A1(_0974_));
 sg13g2_a22oi_1 _2196_ (.Y(_1312_),
    .B1(_1309_),
    .B2(_1311_),
    .A2(_1295_),
    .A1(\levenshtein_ctrl.vp[2] ));
 sg13g2_nor2_1 _2197_ (.A(net378),
    .B(_1312_),
    .Y(_1313_));
 sg13g2_a221oi_1 _2198_ (.B2(_1303_),
    .C1(_1313_),
    .B1(net350),
    .A1(_0972_),
    .Y(_1314_),
    .A2(net745));
 sg13g2_o21ai_1 _2199_ (.B1(_1314_),
    .Y(_0124_),
    .A1(_1304_),
    .A2(_1305_));
 sg13g2_a21oi_1 _2200_ (.A1(net348),
    .A2(_1269_),
    .Y(_1315_),
    .B1(_1286_));
 sg13g2_o21ai_1 _2201_ (.B1(_1315_),
    .Y(_1316_),
    .A1(net750),
    .A2(net348));
 sg13g2_and3_1 _2202_ (.X(_1317_),
    .A(\levenshtein_ctrl.vp[3] ),
    .B(_1306_),
    .C(_1308_));
 sg13g2_nor3_2 _2203_ (.A(\levenshtein_ctrl.pm[4] ),
    .B(\levenshtein_ctrl.vn[4] ),
    .C(_1317_),
    .Y(_0293_));
 sg13g2_a21oi_1 _2204_ (.A1(_1306_),
    .A2(_1308_),
    .Y(_0294_),
    .B1(\levenshtein_ctrl.vp[3] ));
 sg13g2_nor2_1 _2205_ (.A(net757),
    .B(_0294_),
    .Y(_0295_));
 sg13g2_a22oi_1 _2206_ (.Y(_0296_),
    .B1(_0293_),
    .B2(_0295_),
    .A2(_1310_),
    .A1(\levenshtein_ctrl.vp[3] ));
 sg13g2_a22oi_1 _2207_ (.Y(_0297_),
    .B1(_1270_),
    .B2(net350),
    .A2(\levenshtein_ctrl.vp[4] ),
    .A1(net430));
 sg13g2_o21ai_1 _2208_ (.B1(_0297_),
    .Y(_0298_),
    .A1(net378),
    .A2(_0296_));
 sg13g2_nand2b_1 _2209_ (.Y(_0125_),
    .B(_1316_),
    .A_N(_0298_));
 sg13g2_o21ai_1 _2210_ (.B1(net436),
    .Y(_0299_),
    .A1(net348),
    .A2(_1286_));
 sg13g2_nand2_1 _2211_ (.Y(_0300_),
    .A(net728),
    .B(net336));
 sg13g2_nor2_1 _2212_ (.A(_0975_),
    .B(_0293_),
    .Y(_0301_));
 sg13g2_o21ai_1 _2213_ (.B1(\levenshtein_ctrl.vp[4] ),
    .Y(_0302_),
    .A1(\levenshtein_ctrl.pm[4] ),
    .A2(_1317_));
 sg13g2_nand3b_1 _2214_ (.B(_0977_),
    .C(_0302_),
    .Y(_0303_),
    .A_N(\levenshtein_ctrl.pm[5] ));
 sg13g2_nor3_1 _2215_ (.A(\levenshtein_ctrl.vp[4] ),
    .B(\levenshtein_ctrl.pm[4] ),
    .C(_1317_),
    .Y(_0304_));
 sg13g2_nor2_1 _2216_ (.A(\levenshtein_ctrl.vn[4] ),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_nor2b_1 _2217_ (.A(_0303_),
    .B_N(_0305_),
    .Y(_0306_));
 sg13g2_o21ai_1 _2218_ (.B1(net382),
    .Y(_0307_),
    .A1(_0301_),
    .A2(_0306_));
 sg13g2_nor2_2 _2219_ (.A(_0971_),
    .B(net410),
    .Y(_0308_));
 sg13g2_nand2_1 _2220_ (.Y(_0309_),
    .A(_1267_),
    .B(_0308_));
 sg13g2_a21oi_1 _2221_ (.A1(_1267_),
    .A2(_0308_),
    .Y(_0310_),
    .B1(_1269_));
 sg13g2_o21ai_1 _2222_ (.B1(_0310_),
    .Y(_0311_),
    .A1(_1082_),
    .A2(net350));
 sg13g2_nand3_1 _2223_ (.B(_0307_),
    .C(_0311_),
    .A(_0300_),
    .Y(_0126_));
 sg13g2_nand2_1 _2224_ (.Y(_0312_),
    .A(\levenshtein_ctrl.vp[5] ),
    .B(_0303_));
 sg13g2_or2_1 _2225_ (.X(_0313_),
    .B(\levenshtein_ctrl.pm[5] ),
    .A(\levenshtein_ctrl.pm[4] ));
 sg13g2_a21oi_1 _2226_ (.A1(\levenshtein_ctrl.vp[4] ),
    .A2(\levenshtein_ctrl.pm[4] ),
    .Y(_0314_),
    .B1(\levenshtein_ctrl.pm[5] ));
 sg13g2_nand2b_1 _2227_ (.Y(_0315_),
    .B(\levenshtein_ctrl.vp[5] ),
    .A_N(_0314_));
 sg13g2_nand2_1 _2228_ (.Y(_0316_),
    .A(\levenshtein_ctrl.vp[4] ),
    .B(\levenshtein_ctrl.vp[5] ));
 sg13g2_nor2_1 _2229_ (.A(_0313_),
    .B(_0316_),
    .Y(_0317_));
 sg13g2_nand4_1 _2230_ (.B(_1306_),
    .C(_1308_),
    .A(\levenshtein_ctrl.vp[3] ),
    .Y(_0318_),
    .D(_0317_));
 sg13g2_nor2_1 _2231_ (.A(\levenshtein_ctrl.pm[6] ),
    .B(\levenshtein_ctrl.vn[6] ),
    .Y(_0319_));
 sg13g2_nand3_1 _2232_ (.B(_0318_),
    .C(_0319_),
    .A(_0315_),
    .Y(_0320_));
 sg13g2_o21ai_1 _2233_ (.B1(_0977_),
    .Y(_0321_),
    .A1(\levenshtein_ctrl.vp[5] ),
    .A2(_0303_));
 sg13g2_o21ai_1 _2234_ (.B1(_0312_),
    .Y(_0322_),
    .A1(_0320_),
    .A2(_0321_));
 sg13g2_nand2_1 _2235_ (.Y(_0323_),
    .A(net382),
    .B(_0322_));
 sg13g2_nand2b_2 _2236_ (.Y(_0324_),
    .B(\levenshtein_ctrl.word_length_reg[0] ),
    .A_N(net415));
 sg13g2_nor3_2 _2237_ (.A(_0971_),
    .B(net410),
    .C(_0324_),
    .Y(_0325_));
 sg13g2_o21ai_1 _2238_ (.B1(_0323_),
    .Y(_0326_),
    .A1(_0311_),
    .A2(_0325_));
 sg13g2_a21o_1 _2239_ (.A2(net336),
    .A1(net713),
    .B1(_0326_),
    .X(_0127_));
 sg13g2_a21o_1 _2240_ (.A2(\levenshtein_ctrl.pm[6] ),
    .A1(\levenshtein_ctrl.vp[6] ),
    .B1(\levenshtein_ctrl.pm[7] ),
    .X(_0327_));
 sg13g2_nand2b_1 _2241_ (.Y(_0328_),
    .B(\levenshtein_ctrl.vp[6] ),
    .A_N(\levenshtein_ctrl.pm[6] ));
 sg13g2_a21oi_1 _2242_ (.A1(_0315_),
    .A2(_0318_),
    .Y(_0329_),
    .B1(_0328_));
 sg13g2_nor3_2 _2243_ (.A(net698),
    .B(_0327_),
    .C(_0329_),
    .Y(_0330_));
 sg13g2_nand4_1 _2244_ (.B(_0315_),
    .C(_0318_),
    .A(_0978_),
    .Y(_0331_),
    .D(_0319_));
 sg13g2_nor2b_2 _2245_ (.A(net452),
    .B_N(_0331_),
    .Y(_0332_));
 sg13g2_a22oi_1 _2246_ (.Y(_0333_),
    .B1(_0330_),
    .B2(_0332_),
    .A2(_0320_),
    .A1(net713));
 sg13g2_nand3_1 _2247_ (.B(net412),
    .C(\levenshtein_ctrl.word_length_reg[0] ),
    .A(net414),
    .Y(_0334_));
 sg13g2_nand2b_1 _2248_ (.Y(_0335_),
    .B(_0334_),
    .A_N(net410));
 sg13g2_o21ai_1 _2249_ (.B1(net366),
    .Y(_0336_),
    .A1(net345),
    .A2(_0335_));
 sg13g2_a21oi_1 _2250_ (.A1(_0979_),
    .A2(net345),
    .Y(_0337_),
    .B1(_0336_));
 sg13g2_a221oi_1 _2251_ (.B2(_0335_),
    .C1(_0337_),
    .B1(net350),
    .A1(net430),
    .Y(_0338_),
    .A2(net735));
 sg13g2_o21ai_1 _2252_ (.B1(_0338_),
    .Y(_0128_),
    .A1(_1292_),
    .A2(_0333_));
 sg13g2_nand2b_1 _2253_ (.Y(_0339_),
    .B(\levenshtein_ctrl.vp[7] ),
    .A_N(_0330_));
 sg13g2_nand3b_1 _2254_ (.B(\levenshtein_ctrl.vp[7] ),
    .C(\levenshtein_ctrl.vp[6] ),
    .Y(_0340_),
    .A_N(\levenshtein_ctrl.pm[6] ));
 sg13g2_nor4_1 _2255_ (.A(\levenshtein_ctrl.pm[7] ),
    .B(_0313_),
    .C(_0316_),
    .D(_0340_),
    .Y(_0341_));
 sg13g2_nand4_1 _2256_ (.B(_1306_),
    .C(_1308_),
    .A(\levenshtein_ctrl.vp[3] ),
    .Y(_0342_),
    .D(_0341_));
 sg13g2_nor4_1 _2257_ (.A(_0976_),
    .B(\levenshtein_ctrl.pm[7] ),
    .C(_0314_),
    .D(_0340_),
    .Y(_0343_));
 sg13g2_a21oi_2 _2258_ (.B1(_0343_),
    .Y(_0344_),
    .A2(_0327_),
    .A1(\levenshtein_ctrl.vp[7] ));
 sg13g2_nor2_1 _2259_ (.A(\levenshtein_ctrl.pm[8] ),
    .B(\levenshtein_ctrl.vn[8] ),
    .Y(_0345_));
 sg13g2_nand3_1 _2260_ (.B(_0344_),
    .C(_0345_),
    .A(_0342_),
    .Y(_0346_));
 sg13g2_nor3_1 _2261_ (.A(\levenshtein_ctrl.vp[7] ),
    .B(_0327_),
    .C(_0329_),
    .Y(_0347_));
 sg13g2_nor2_1 _2262_ (.A(\levenshtein_ctrl.vn[7] ),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_nand2b_1 _2263_ (.Y(_0349_),
    .B(_0348_),
    .A_N(_0346_));
 sg13g2_a21oi_1 _2264_ (.A1(_0339_),
    .A2(_0349_),
    .Y(_0350_),
    .B1(net378));
 sg13g2_nor2_1 _2265_ (.A(net739),
    .B(net349),
    .Y(_0351_));
 sg13g2_o21ai_1 _2266_ (.B1(_1287_),
    .Y(_0352_),
    .A1(net410),
    .A2(net345));
 sg13g2_and2_1 _2267_ (.A(net409),
    .B(net350),
    .X(_0353_));
 sg13g2_a221oi_1 _2268_ (.B2(net411),
    .C1(_0350_),
    .B1(_1298_),
    .A1(net430),
    .Y(_0354_),
    .A2(net739));
 sg13g2_o21ai_1 _2269_ (.B1(_0354_),
    .Y(_0129_),
    .A1(_0351_),
    .A2(_0352_));
 sg13g2_a21oi_1 _2270_ (.A1(\levenshtein_ctrl.vp[8] ),
    .A2(\levenshtein_ctrl.pm[8] ),
    .Y(_0355_),
    .B1(\levenshtein_ctrl.pm[9] ));
 sg13g2_a21o_1 _2271_ (.A2(\levenshtein_ctrl.pm[8] ),
    .A1(\levenshtein_ctrl.vp[8] ),
    .B1(\levenshtein_ctrl.pm[9] ),
    .X(_0356_));
 sg13g2_nand2b_1 _2272_ (.Y(_0357_),
    .B(\levenshtein_ctrl.vp[8] ),
    .A_N(\levenshtein_ctrl.pm[8] ));
 sg13g2_a21oi_2 _2273_ (.B1(_0357_),
    .Y(_0358_),
    .A2(_0344_),
    .A1(_0342_));
 sg13g2_a21o_1 _2274_ (.A2(_0344_),
    .A1(_0342_),
    .B1(_0357_),
    .X(_0359_));
 sg13g2_nor3_2 _2275_ (.A(\levenshtein_ctrl.vn[9] ),
    .B(_0356_),
    .C(_0358_),
    .Y(_0360_));
 sg13g2_nor2_1 _2276_ (.A(\levenshtein_ctrl.vp[8] ),
    .B(_0346_),
    .Y(_0361_));
 sg13g2_nor2_1 _2277_ (.A(net481),
    .B(_0361_),
    .Y(_0362_));
 sg13g2_a22oi_1 _2278_ (.Y(_0363_),
    .B1(_0360_),
    .B2(_0362_),
    .A2(_0346_),
    .A1(net758));
 sg13g2_nor2_1 _2279_ (.A(net378),
    .B(net759),
    .Y(_0364_));
 sg13g2_o21ai_1 _2280_ (.B1(net409),
    .Y(_0365_),
    .A1(net412),
    .A2(_1268_));
 sg13g2_a21oi_1 _2281_ (.A1(net349),
    .A2(_1287_),
    .Y(_0366_),
    .B1(net350));
 sg13g2_nand2_1 _2282_ (.Y(_0367_),
    .A(\levenshtein_ctrl.vp[9] ),
    .B(_1287_));
 sg13g2_a21oi_1 _2283_ (.A1(net349),
    .A2(_0365_),
    .Y(_0368_),
    .B1(_0367_));
 sg13g2_a21oi_1 _2284_ (.A1(net430),
    .A2(\levenshtein_ctrl.vp[9] ),
    .Y(_0369_),
    .B1(_0368_));
 sg13g2_o21ai_1 _2285_ (.B1(_0369_),
    .Y(_0370_),
    .A1(_0365_),
    .A2(_0366_));
 sg13g2_or2_1 _2286_ (.X(_0130_),
    .B(_0370_),
    .A(_0364_));
 sg13g2_nor2_1 _2287_ (.A(_0980_),
    .B(_0360_),
    .Y(_0371_));
 sg13g2_a21oi_2 _2288_ (.B1(_0980_),
    .Y(_0372_),
    .A2(_0359_),
    .A1(_0355_));
 sg13g2_o21ai_1 _2289_ (.B1(\levenshtein_ctrl.vp[9] ),
    .Y(_0373_),
    .A1(_0356_),
    .A2(_0358_));
 sg13g2_nor3_2 _2290_ (.A(net658),
    .B(net565),
    .C(_0372_),
    .Y(_0374_));
 sg13g2_nor3_1 _2291_ (.A(\levenshtein_ctrl.vp[9] ),
    .B(_0356_),
    .C(_0358_),
    .Y(_0375_));
 sg13g2_nor2_2 _2292_ (.A(net654),
    .B(_0375_),
    .Y(_0376_));
 sg13g2_a21oi_1 _2293_ (.A1(_0374_),
    .A2(_0376_),
    .Y(_0377_),
    .B1(_0371_));
 sg13g2_nor2_1 _2294_ (.A(net412),
    .B(_0324_),
    .Y(_0378_));
 sg13g2_nor3_1 _2295_ (.A(_0365_),
    .B(_0366_),
    .C(_0378_),
    .Y(_0379_));
 sg13g2_a21oi_1 _2296_ (.A1(net723),
    .A2(net336),
    .Y(_0380_),
    .B1(_0379_));
 sg13g2_o21ai_1 _2297_ (.B1(_0380_),
    .Y(_0131_),
    .A1(net379),
    .A2(_0377_));
 sg13g2_nor2b_1 _2298_ (.A(_0374_),
    .B_N(net723),
    .Y(_0381_));
 sg13g2_nor2_1 _2299_ (.A(\levenshtein_ctrl.vp[10] ),
    .B(net760),
    .Y(_0382_));
 sg13g2_nor2_1 _2300_ (.A(\levenshtein_ctrl.pm[10] ),
    .B(\levenshtein_ctrl.pm[11] ),
    .Y(_0383_));
 sg13g2_a21oi_2 _2301_ (.B1(_0382_),
    .Y(_0384_),
    .A2(_0383_),
    .A1(_0373_));
 sg13g2_nor2_1 _2302_ (.A(net551),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_nor3_1 _2303_ (.A(\levenshtein_ctrl.vp[10] ),
    .B(\levenshtein_ctrl.pm[10] ),
    .C(_0372_),
    .Y(_0386_));
 sg13g2_or2_1 _2304_ (.X(_0387_),
    .B(_0386_),
    .A(\levenshtein_ctrl.vn[10] ));
 sg13g2_inv_1 _2305_ (.Y(_0388_),
    .A(_0387_));
 sg13g2_a21oi_1 _2306_ (.A1(_0385_),
    .A2(_0388_),
    .Y(_0389_),
    .B1(_0381_));
 sg13g2_o21ai_1 _2307_ (.B1(net366),
    .Y(_0390_),
    .A1(\levenshtein_ctrl.vp[11] ),
    .A2(net349));
 sg13g2_a21oi_1 _2308_ (.A1(net409),
    .A2(_1302_),
    .Y(_0391_),
    .B1(net345));
 sg13g2_nor2_1 _2309_ (.A(_0390_),
    .B(_0391_),
    .Y(_0392_));
 sg13g2_a221oi_1 _2310_ (.B2(_0353_),
    .C1(_0392_),
    .B1(_1302_),
    .A1(net430),
    .Y(_0393_),
    .A2(net737));
 sg13g2_o21ai_1 _2311_ (.B1(_0393_),
    .Y(_0132_),
    .A1(net379),
    .A2(_0389_));
 sg13g2_o21ai_1 _2312_ (.B1(\levenshtein_ctrl.vp[11] ),
    .Y(_0394_),
    .A1(\levenshtein_ctrl.vn[11] ),
    .A2(_0384_));
 sg13g2_nand4_1 _2313_ (.B(\levenshtein_ctrl.vp[10] ),
    .C(\levenshtein_ctrl.vp[11] ),
    .A(\levenshtein_ctrl.vp[9] ),
    .Y(_0395_),
    .D(_0383_));
 sg13g2_or3_1 _2314_ (.A(\levenshtein_ctrl.pm[9] ),
    .B(_0357_),
    .C(_0395_),
    .X(_0396_));
 sg13g2_a21oi_2 _2315_ (.B1(_0396_),
    .Y(_0397_),
    .A2(_0344_),
    .A1(_0342_));
 sg13g2_o21ai_1 _2316_ (.B1(\levenshtein_ctrl.vp[11] ),
    .Y(_0398_),
    .A1(\levenshtein_ctrl.vp[10] ),
    .A2(\levenshtein_ctrl.pm[11] ));
 sg13g2_or2_1 _2317_ (.X(_0399_),
    .B(_0398_),
    .A(_0383_));
 sg13g2_o21ai_1 _2318_ (.B1(_0399_),
    .Y(_0400_),
    .A1(_0355_),
    .A2(_0395_));
 sg13g2_or4_2 _2319_ (.A(\levenshtein_ctrl.pm[12] ),
    .B(\levenshtein_ctrl.vn[12] ),
    .C(_0397_),
    .D(_0400_),
    .X(_0401_));
 sg13g2_o21ai_1 _2320_ (.B1(_0981_),
    .Y(_0402_),
    .A1(\levenshtein_ctrl.vp[11] ),
    .A2(_0384_));
 sg13g2_o21ai_1 _2321_ (.B1(_0394_),
    .Y(_0403_),
    .A1(_0401_),
    .A2(_0402_));
 sg13g2_and2_2 _2322_ (.A(net412),
    .B(net409),
    .X(_0404_));
 sg13g2_nand2_1 _2323_ (.Y(_0405_),
    .A(net412),
    .B(net409));
 sg13g2_nand3_1 _2324_ (.B(net366),
    .C(_0404_),
    .A(net347),
    .Y(_0406_));
 sg13g2_nand2_1 _2325_ (.Y(_0407_),
    .A(net412),
    .B(_0353_));
 sg13g2_inv_1 _2326_ (.Y(_0408_),
    .A(_0407_));
 sg13g2_nand2_1 _2327_ (.Y(_0409_),
    .A(net429),
    .B(\levenshtein_ctrl.vp[12] ));
 sg13g2_nand3_1 _2328_ (.B(net345),
    .C(net366),
    .A(\levenshtein_ctrl.vp[12] ),
    .Y(_0410_));
 sg13g2_nand4_1 _2329_ (.B(_0407_),
    .C(_0409_),
    .A(_0406_),
    .Y(_0411_),
    .D(_0410_));
 sg13g2_a21o_1 _2330_ (.A2(_0403_),
    .A1(net380),
    .B1(_0411_),
    .X(_0133_));
 sg13g2_a21o_1 _2331_ (.A2(\levenshtein_ctrl.pm[12] ),
    .A1(\levenshtein_ctrl.vp[12] ),
    .B1(\levenshtein_ctrl.pm[13] ),
    .X(_0412_));
 sg13g2_o21ai_1 _2332_ (.B1(\levenshtein_ctrl.vp[12] ),
    .Y(_0413_),
    .A1(_0397_),
    .A2(_0400_));
 sg13g2_nand2b_1 _2333_ (.Y(_0414_),
    .B(_0413_),
    .A_N(_0412_));
 sg13g2_nor2_1 _2334_ (.A(net614),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_or2_1 _2335_ (.X(_0416_),
    .B(_0401_),
    .A(\levenshtein_ctrl.vp[12] ));
 sg13g2_and2_1 _2336_ (.A(_0982_),
    .B(_0416_),
    .X(_0417_));
 sg13g2_a22oi_1 _2337_ (.Y(_0418_),
    .B1(_0415_),
    .B2(_0417_),
    .A2(_0401_),
    .A1(net742));
 sg13g2_o21ai_1 _2338_ (.B1(net366),
    .Y(_0419_),
    .A1(\levenshtein_ctrl.vp[13] ),
    .A2(net347));
 sg13g2_a21oi_1 _2339_ (.A1(_1268_),
    .A2(_0404_),
    .Y(_0420_),
    .B1(net344));
 sg13g2_nor2_1 _2340_ (.A(_0419_),
    .B(_0420_),
    .Y(_0421_));
 sg13g2_a221oi_1 _2341_ (.B2(_0408_),
    .C1(_0421_),
    .B1(_1268_),
    .A1(net430),
    .Y(_0422_),
    .A2(\levenshtein_ctrl.vp[13] ));
 sg13g2_o21ai_1 _2342_ (.B1(_0422_),
    .Y(_0134_),
    .A1(net379),
    .A2(net743));
 sg13g2_o21ai_1 _2343_ (.B1(\levenshtein_ctrl.vp[13] ),
    .Y(_0423_),
    .A1(\levenshtein_ctrl.vn[13] ),
    .A2(_0414_));
 sg13g2_nand3b_1 _2344_ (.B(\levenshtein_ctrl.vp[13] ),
    .C(\levenshtein_ctrl.vp[12] ),
    .Y(_0424_),
    .A_N(\levenshtein_ctrl.pm[12] ));
 sg13g2_nor2_1 _2345_ (.A(\levenshtein_ctrl.pm[13] ),
    .B(_0424_),
    .Y(_0425_));
 sg13g2_o21ai_1 _2346_ (.B1(_0425_),
    .Y(_0426_),
    .A1(_0397_),
    .A2(_0400_));
 sg13g2_a21oi_1 _2347_ (.A1(\levenshtein_ctrl.vp[13] ),
    .A2(_0412_),
    .Y(_0427_),
    .B1(\levenshtein_ctrl.pm[14] ));
 sg13g2_nand3_1 _2348_ (.B(_0426_),
    .C(_0427_),
    .A(_0985_),
    .Y(_0428_));
 sg13g2_o21ai_1 _2349_ (.B1(_0983_),
    .Y(_0429_),
    .A1(\levenshtein_ctrl.vp[13] ),
    .A2(_0414_));
 sg13g2_o21ai_1 _2350_ (.B1(_0423_),
    .Y(_0430_),
    .A1(_0428_),
    .A2(_0429_));
 sg13g2_nand2_1 _2351_ (.Y(_0431_),
    .A(net380),
    .B(_0430_));
 sg13g2_nand4_1 _2352_ (.B(net347),
    .C(net366),
    .A(net414),
    .Y(_0432_),
    .D(_0404_));
 sg13g2_a22oi_1 _2353_ (.Y(_0433_),
    .B1(_0408_),
    .B2(net414),
    .A2(net741),
    .A1(net429));
 sg13g2_nand3_1 _2354_ (.B(net345),
    .C(net366),
    .A(net741),
    .Y(_0434_));
 sg13g2_nand4_1 _2355_ (.B(_0432_),
    .C(_0433_),
    .A(_0431_),
    .Y(_0135_),
    .D(_0434_));
 sg13g2_nand2_1 _2356_ (.Y(_0435_),
    .A(net741),
    .B(_0428_));
 sg13g2_a21oi_1 _2357_ (.A1(_0426_),
    .A2(_0427_),
    .Y(_0436_),
    .B1(_0984_));
 sg13g2_xnor2_1 _2358_ (.Y(_0437_),
    .A(\levenshtein_ctrl.vp[15] ),
    .B(_0033_));
 sg13g2_xnor2_1 _2359_ (.Y(_0438_),
    .A(_0436_),
    .B(_0437_));
 sg13g2_nor2b_1 _2360_ (.A(\levenshtein_ctrl.pm[15] ),
    .B_N(_0031_),
    .Y(_0439_));
 sg13g2_nand2_1 _2361_ (.Y(_0440_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_nand3_1 _2362_ (.B(_0426_),
    .C(_0427_),
    .A(_0984_),
    .Y(_0441_));
 sg13g2_nand2_2 _2363_ (.Y(_0442_),
    .A(_0985_),
    .B(_0441_));
 sg13g2_o21ai_1 _2364_ (.B1(_0435_),
    .Y(_0443_),
    .A1(_0440_),
    .A2(_0442_));
 sg13g2_nor2_2 _2365_ (.A(_1301_),
    .B(_0405_),
    .Y(_0444_));
 sg13g2_inv_1 _2366_ (.Y(_0445_),
    .A(_0444_));
 sg13g2_a22oi_1 _2367_ (.Y(_0446_),
    .B1(net350),
    .B2(_0444_),
    .A2(net746),
    .A1(net429));
 sg13g2_nor2_1 _2368_ (.A(net344),
    .B(_0445_),
    .Y(_0447_));
 sg13g2_a21oi_1 _2369_ (.A1(net746),
    .A2(net344),
    .Y(_0448_),
    .B1(_0447_));
 sg13g2_o21ai_1 _2370_ (.B1(_0446_),
    .Y(_0449_),
    .A1(_1286_),
    .A2(_0448_));
 sg13g2_a21o_1 _2371_ (.A2(_0443_),
    .A1(net381),
    .B1(_0449_),
    .X(_0136_));
 sg13g2_a22oi_1 _2372_ (.Y(_0450_),
    .B1(net335),
    .B2(net269),
    .A2(net382),
    .A1(_1280_));
 sg13g2_inv_1 _2373_ (.Y(_0137_),
    .A(net270));
 sg13g2_nand2_1 _2374_ (.Y(_0451_),
    .A(net283),
    .B(net335));
 sg13g2_nand3_1 _2375_ (.B(_1278_),
    .C(net382),
    .A(_1277_),
    .Y(_0452_));
 sg13g2_nand2_1 _2376_ (.Y(_0138_),
    .A(_0451_),
    .B(_0452_));
 sg13g2_nand2_1 _2377_ (.Y(_0453_),
    .A(net441),
    .B(net335));
 sg13g2_nand3_1 _2378_ (.B(_1295_),
    .C(_1296_),
    .A(net382),
    .Y(_0454_));
 sg13g2_nand2_1 _2379_ (.Y(_0139_),
    .A(_0453_),
    .B(_0454_));
 sg13g2_nor3_1 _2380_ (.A(net378),
    .B(_1309_),
    .C(_1311_),
    .Y(_0455_));
 sg13g2_a21o_1 _2381_ (.A2(net335),
    .A1(net676),
    .B1(_0455_),
    .X(_0140_));
 sg13g2_nor3_1 _2382_ (.A(net378),
    .B(_0293_),
    .C(_0295_),
    .Y(_0456_));
 sg13g2_a21o_1 _2383_ (.A2(net335),
    .A1(net581),
    .B1(_0456_),
    .X(_0141_));
 sg13g2_nand2_1 _2384_ (.Y(_0457_),
    .A(net308),
    .B(net335));
 sg13g2_nand2_1 _2385_ (.Y(_0458_),
    .A(net382),
    .B(_0303_));
 sg13g2_o21ai_1 _2386_ (.B1(_0457_),
    .Y(_0142_),
    .A1(_0305_),
    .A2(_0458_));
 sg13g2_nand2_1 _2387_ (.Y(_0459_),
    .A(net452),
    .B(net335));
 sg13g2_nand3_1 _2388_ (.B(_0320_),
    .C(_0321_),
    .A(net382),
    .Y(_0460_));
 sg13g2_nand2_1 _2389_ (.Y(_0143_),
    .A(_0459_),
    .B(_0460_));
 sg13g2_nor3_1 _2390_ (.A(net378),
    .B(_0330_),
    .C(_0332_),
    .Y(_0461_));
 sg13g2_a21o_1 _2391_ (.A2(net335),
    .A1(net698),
    .B1(_0461_),
    .X(_0144_));
 sg13g2_nand2_1 _2392_ (.Y(_0462_),
    .A(net481),
    .B(net336));
 sg13g2_nand2_1 _2393_ (.Y(_0463_),
    .A(net382),
    .B(_0346_));
 sg13g2_o21ai_1 _2394_ (.B1(_0462_),
    .Y(_0145_),
    .A1(_0348_),
    .A2(_0463_));
 sg13g2_nor3_1 _2395_ (.A(net378),
    .B(_0360_),
    .C(_0362_),
    .Y(_0464_));
 sg13g2_a21o_1 _2396_ (.A2(net336),
    .A1(net654),
    .B1(_0464_),
    .X(_0146_));
 sg13g2_nor3_1 _2397_ (.A(net379),
    .B(_0374_),
    .C(_0376_),
    .Y(_0465_));
 sg13g2_a21o_1 _2398_ (.A2(net334),
    .A1(net565),
    .B1(_0465_),
    .X(_0147_));
 sg13g2_a22oi_1 _2399_ (.Y(_0466_),
    .B1(_0387_),
    .B2(net381),
    .A2(net334),
    .A1(net551));
 sg13g2_nor2_1 _2400_ (.A(_0385_),
    .B(net552),
    .Y(_0148_));
 sg13g2_nand2_1 _2401_ (.Y(_0467_),
    .A(net324),
    .B(_0299_));
 sg13g2_nand3_1 _2402_ (.B(_0401_),
    .C(_0402_),
    .A(net380),
    .Y(_0468_));
 sg13g2_nand2_1 _2403_ (.Y(_0149_),
    .A(_0467_),
    .B(_0468_));
 sg13g2_nor3_1 _2404_ (.A(net379),
    .B(_0415_),
    .C(_0417_),
    .Y(_0469_));
 sg13g2_a21o_1 _2405_ (.A2(net334),
    .A1(net614),
    .B1(_0469_),
    .X(_0150_));
 sg13g2_and2_1 _2406_ (.A(net380),
    .B(_0428_),
    .X(_0470_));
 sg13g2_a22oi_1 _2407_ (.Y(_0471_),
    .B1(_0429_),
    .B2(_0470_),
    .A2(net334),
    .A1(net438));
 sg13g2_inv_1 _2408_ (.Y(_0151_),
    .A(_0471_));
 sg13g2_nand2_1 _2409_ (.Y(_0472_),
    .A(net285),
    .B(net334));
 sg13g2_nand3_1 _2410_ (.B(_0440_),
    .C(_0442_),
    .A(net380),
    .Y(_0473_));
 sg13g2_nand2_1 _2411_ (.Y(_0152_),
    .A(_0472_),
    .B(_0473_));
 sg13g2_nand2b_1 _2412_ (.Y(_0474_),
    .B(_0444_),
    .A_N(_0033_));
 sg13g2_a21oi_1 _2413_ (.A1(_0438_),
    .A2(_0439_),
    .Y(_0475_),
    .B1(_0474_));
 sg13g2_nand2_1 _2414_ (.Y(_0476_),
    .A(_0971_),
    .B(net409));
 sg13g2_nor2_1 _2415_ (.A(_1301_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_nor2b_1 _2416_ (.A(_0394_),
    .B_N(_0477_),
    .Y(_0478_));
 sg13g2_nor2b_2 _2417_ (.A(\levenshtein_ctrl.word_length_reg[0] ),
    .B_N(net414),
    .Y(_0479_));
 sg13g2_and2_1 _2418_ (.A(_0404_),
    .B(_0479_),
    .X(_0480_));
 sg13g2_nand3_1 _2419_ (.B(_0428_),
    .C(_0480_),
    .A(\levenshtein_ctrl.vp[14] ),
    .Y(_0481_));
 sg13g2_nor2_1 _2420_ (.A(_0324_),
    .B(_0476_),
    .Y(_0482_));
 sg13g2_inv_1 _2421_ (.Y(_0483_),
    .A(_0482_));
 sg13g2_nand2_1 _2422_ (.Y(_0484_),
    .A(_0371_),
    .B(_0482_));
 sg13g2_nand4_1 _2423_ (.B(_0308_),
    .C(_0320_),
    .A(\levenshtein_ctrl.vp[6] ),
    .Y(_0485_),
    .D(_0479_));
 sg13g2_nor3_1 _2424_ (.A(_0975_),
    .B(_0293_),
    .C(_0309_),
    .Y(_0486_));
 sg13g2_nor2_1 _2425_ (.A(_1270_),
    .B(_1301_),
    .Y(_0487_));
 sg13g2_nand3_1 _2426_ (.B(_1310_),
    .C(_0487_),
    .A(\levenshtein_ctrl.vp[3] ),
    .Y(_0488_));
 sg13g2_nand2_1 _2427_ (.Y(_0489_),
    .A(_1269_),
    .B(_0479_));
 sg13g2_nand4_1 _2428_ (.B(_1269_),
    .C(_1295_),
    .A(\levenshtein_ctrl.vp[2] ),
    .Y(_0490_),
    .D(_0479_));
 sg13g2_nand3_1 _2429_ (.B(_1272_),
    .C(_1280_),
    .A(\levenshtein_ctrl.vp[0] ),
    .Y(_0491_));
 sg13g2_nor2_1 _2430_ (.A(_1270_),
    .B(_0324_),
    .Y(_0492_));
 sg13g2_nand3_1 _2431_ (.B(_1277_),
    .C(_0492_),
    .A(\levenshtein_ctrl.vp[1] ),
    .Y(_0493_));
 sg13g2_nand4_1 _2432_ (.B(_0490_),
    .C(_0491_),
    .A(_0488_),
    .Y(_0494_),
    .D(_0493_));
 sg13g2_nand3_1 _2433_ (.B(_0303_),
    .C(_0325_),
    .A(\levenshtein_ctrl.vp[5] ),
    .Y(_0495_));
 sg13g2_nand2_1 _2434_ (.Y(_0496_),
    .A(net409),
    .B(_1271_));
 sg13g2_and4_1 _2435_ (.A(net410),
    .B(\levenshtein_ctrl.vp[8] ),
    .C(_1271_),
    .D(_0346_),
    .X(_0497_));
 sg13g2_nor3_1 _2436_ (.A(_0486_),
    .B(_0494_),
    .C(_0497_),
    .Y(_0498_));
 sg13g2_nor2_1 _2437_ (.A(net409),
    .B(_0334_),
    .Y(_0499_));
 sg13g2_nand2b_1 _2438_ (.Y(_0500_),
    .B(_0499_),
    .A_N(_0339_));
 sg13g2_nand2_1 _2439_ (.Y(_0501_),
    .A(_1267_),
    .B(_0404_));
 sg13g2_nand4_1 _2440_ (.B(_1267_),
    .C(_0401_),
    .A(\levenshtein_ctrl.vp[12] ),
    .Y(_0502_),
    .D(_0404_));
 sg13g2_and4_1 _2441_ (.A(_0485_),
    .B(_0495_),
    .C(_0498_),
    .D(_0502_),
    .X(_0503_));
 sg13g2_nand4_1 _2442_ (.B(_0484_),
    .C(_0500_),
    .A(_0481_),
    .Y(_0504_),
    .D(_0503_));
 sg13g2_nor2b_1 _2443_ (.A(_0476_),
    .B_N(_0479_),
    .Y(_0505_));
 sg13g2_nand3b_1 _2444_ (.B(_0505_),
    .C(\levenshtein_ctrl.vp[10] ),
    .Y(_0506_),
    .A_N(_0374_));
 sg13g2_nor2_1 _2445_ (.A(_0324_),
    .B(_0405_),
    .Y(_0507_));
 sg13g2_inv_1 _2446_ (.Y(_0508_),
    .A(_0507_));
 sg13g2_o21ai_1 _2447_ (.B1(_0506_),
    .Y(_0509_),
    .A1(_0423_),
    .A2(_0508_));
 sg13g2_nor4_2 _2448_ (.A(_0475_),
    .B(_0478_),
    .C(_0504_),
    .Y(_0510_),
    .D(_0509_));
 sg13g2_or4_2 _2449_ (.A(_0475_),
    .B(_0478_),
    .C(_0504_),
    .D(_0509_),
    .X(_0511_));
 sg13g2_nand3b_1 _2450_ (.B(_0438_),
    .C(_0439_),
    .Y(_0512_),
    .A_N(\levenshtein_ctrl.vp[15] ));
 sg13g2_nand2_1 _2451_ (.Y(_0513_),
    .A(_0031_),
    .B(_0512_));
 sg13g2_a21oi_2 _2452_ (.B1(_0445_),
    .Y(_0514_),
    .A2(_0512_),
    .A1(_0031_));
 sg13g2_nand2_1 _2453_ (.Y(_0515_),
    .A(_0429_),
    .B(_0507_));
 sg13g2_a22oi_1 _2454_ (.Y(_0516_),
    .B1(_0505_),
    .B2(_0387_),
    .A2(_0480_),
    .A1(_0442_));
 sg13g2_nand2_1 _2455_ (.Y(_0517_),
    .A(_0402_),
    .B(_0477_));
 sg13g2_o21ai_1 _2456_ (.B1(_0487_),
    .Y(_0518_),
    .A1(\levenshtein_ctrl.vn[3] ),
    .A2(_0294_));
 sg13g2_a22oi_1 _2457_ (.Y(_0519_),
    .B1(_1296_),
    .B2(_0492_),
    .A2(_1278_),
    .A1(_1272_));
 sg13g2_o21ai_1 _2458_ (.B1(_0519_),
    .Y(_0520_),
    .A1(_1311_),
    .A2(_0489_));
 sg13g2_nor2b_1 _2459_ (.A(_0520_),
    .B_N(_0518_),
    .Y(_0521_));
 sg13g2_o21ai_1 _2460_ (.B1(_0521_),
    .Y(_0522_),
    .A1(_0305_),
    .A2(_0309_));
 sg13g2_a21o_1 _2461_ (.A2(_0325_),
    .A1(_0321_),
    .B1(_0522_),
    .X(_0523_));
 sg13g2_nand3b_1 _2462_ (.B(_0479_),
    .C(_0308_),
    .Y(_0524_),
    .A_N(_0332_));
 sg13g2_o21ai_1 _2463_ (.B1(_0524_),
    .Y(_0525_),
    .A1(_0362_),
    .A2(_0496_));
 sg13g2_o21ai_1 _2464_ (.B1(_0499_),
    .Y(_0526_),
    .A1(\levenshtein_ctrl.vn[7] ),
    .A2(_0347_));
 sg13g2_o21ai_1 _2465_ (.B1(_0526_),
    .Y(_0527_),
    .A1(_0376_),
    .A2(_0483_));
 sg13g2_a21oi_2 _2466_ (.B1(_0501_),
    .Y(_0528_),
    .A2(_0416_),
    .A1(_0982_));
 sg13g2_nor4_2 _2467_ (.A(_0523_),
    .B(_0525_),
    .C(_0527_),
    .Y(_0529_),
    .D(_0528_));
 sg13g2_nand4_1 _2468_ (.B(_0516_),
    .C(_0517_),
    .A(_0515_),
    .Y(_0530_),
    .D(_0529_));
 sg13g2_nor2_2 _2469_ (.A(_0514_),
    .B(_0530_),
    .Y(_0531_));
 sg13g2_or2_2 _2470_ (.X(_0532_),
    .B(_0530_),
    .A(_0514_));
 sg13g2_a21oi_1 _2471_ (.A1(_0510_),
    .A2(_0531_),
    .Y(_0533_),
    .B1(net267));
 sg13g2_nor2_2 _2472_ (.A(_1026_),
    .B(net347),
    .Y(_0534_));
 sg13g2_nand2_1 _2473_ (.Y(_0535_),
    .A(_1027_),
    .B(net344));
 sg13g2_nor2_1 _2474_ (.A(_0055_),
    .B(_0534_),
    .Y(_0536_));
 sg13g2_a21oi_1 _2475_ (.A1(_0939_),
    .A2(_0534_),
    .Y(_0537_),
    .B1(_0536_));
 sg13g2_nor4_1 _2476_ (.A(_0511_),
    .B(_0514_),
    .C(_0530_),
    .D(_0537_),
    .Y(_0538_));
 sg13g2_nand2b_1 _2477_ (.Y(_0539_),
    .B(net381),
    .A_N(_0538_));
 sg13g2_o21ai_1 _2478_ (.B1(net395),
    .Y(_0540_),
    .A1(_0055_),
    .A2(_1040_));
 sg13g2_a21oi_1 _2479_ (.A1(_0939_),
    .A2(net344),
    .Y(_0541_),
    .B1(_0540_));
 sg13g2_a221oi_1 _2480_ (.B2(_0537_),
    .C1(_0541_),
    .B1(_1284_),
    .A1(\levenshtein_ctrl.d[0] ),
    .Y(_0542_),
    .A2(net429));
 sg13g2_o21ai_1 _2481_ (.B1(_0542_),
    .Y(_0153_),
    .A1(_0533_),
    .A2(_0539_));
 sg13g2_xor2_1 _2482_ (.B(\levenshtein_ctrl.word_length_reg[0] ),
    .A(net414),
    .X(_0543_));
 sg13g2_nor2_1 _2483_ (.A(_0534_),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_a21oi_1 _2484_ (.A1(_0941_),
    .A2(_0534_),
    .Y(_0545_),
    .B1(_0544_));
 sg13g2_nand2_1 _2485_ (.Y(_0546_),
    .A(_0510_),
    .B(_0545_));
 sg13g2_xnor2_1 _2486_ (.Y(_0547_),
    .A(\levenshtein_ctrl.d[0] ),
    .B(\levenshtein_ctrl.d[1] ));
 sg13g2_a221oi_1 _2487_ (.B2(_0511_),
    .C1(_0530_),
    .B1(_0547_),
    .A1(_0444_),
    .Y(_0548_),
    .A2(_0513_));
 sg13g2_a221oi_1 _2488_ (.B2(_0546_),
    .C1(net379),
    .B1(_0548_),
    .A1(_0532_),
    .Y(_0549_),
    .A2(_0547_));
 sg13g2_o21ai_1 _2489_ (.B1(net395),
    .Y(_0550_),
    .A1(\levenshtein_ctrl.d[1] ),
    .A2(net347));
 sg13g2_nor2_1 _2490_ (.A(net344),
    .B(_0543_),
    .Y(_0551_));
 sg13g2_a22oi_1 _2491_ (.Y(_0552_),
    .B1(_1284_),
    .B2(_0545_),
    .A2(net429),
    .A1(\levenshtein_ctrl.d[1] ));
 sg13g2_o21ai_1 _2492_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_0550_),
    .A2(_0551_));
 sg13g2_or2_1 _2493_ (.X(_0154_),
    .B(_0553_),
    .A(_0549_));
 sg13g2_nand2_1 _2494_ (.Y(_0554_),
    .A(_1302_),
    .B(_0334_));
 sg13g2_nand2_1 _2495_ (.Y(_0555_),
    .A(\levenshtein_ctrl.d[2] ),
    .B(_0534_));
 sg13g2_o21ai_1 _2496_ (.B1(_0555_),
    .Y(_0556_),
    .A1(_0534_),
    .A2(_0554_));
 sg13g2_nor3_2 _2497_ (.A(\levenshtein_ctrl.d[0] ),
    .B(\levenshtein_ctrl.d[1] ),
    .C(\levenshtein_ctrl.d[2] ),
    .Y(_0557_));
 sg13g2_o21ai_1 _2498_ (.B1(\levenshtein_ctrl.d[2] ),
    .Y(_0558_),
    .A1(\levenshtein_ctrl.d[0] ),
    .A2(\levenshtein_ctrl.d[1] ));
 sg13g2_nand2b_1 _2499_ (.Y(_0559_),
    .B(_0558_),
    .A_N(_0557_));
 sg13g2_mux2_1 _2500_ (.A0(_0556_),
    .A1(_0559_),
    .S(_0511_),
    .X(_0560_));
 sg13g2_nor2_1 _2501_ (.A(_0532_),
    .B(_0560_),
    .Y(_0561_));
 sg13g2_nand3_1 _2502_ (.B(\levenshtein_ctrl.d[1] ),
    .C(\levenshtein_ctrl.d[2] ),
    .A(\levenshtein_ctrl.d[0] ),
    .Y(_0562_));
 sg13g2_o21ai_1 _2503_ (.B1(_0943_),
    .Y(_0563_),
    .A1(_0939_),
    .A2(_0941_));
 sg13g2_and2_1 _2504_ (.A(_0562_),
    .B(_0563_),
    .X(_0564_));
 sg13g2_o21ai_1 _2505_ (.B1(net381),
    .Y(_0565_),
    .A1(_0531_),
    .A2(_0564_));
 sg13g2_o21ai_1 _2506_ (.B1(net395),
    .Y(_0566_),
    .A1(\levenshtein_ctrl.d[2] ),
    .A2(net347));
 sg13g2_a21oi_1 _2507_ (.A1(net347),
    .A2(_0554_),
    .Y(_0567_),
    .B1(_0566_));
 sg13g2_a221oi_1 _2508_ (.B2(_0556_),
    .C1(_0567_),
    .B1(_1284_),
    .A1(net752),
    .Y(_0568_),
    .A2(net429));
 sg13g2_o21ai_1 _2509_ (.B1(_0568_),
    .Y(_0155_),
    .A1(_0561_),
    .A2(_0565_));
 sg13g2_xor2_1 _2510_ (.B(_0334_),
    .A(net411),
    .X(_0569_));
 sg13g2_nor2_1 _2511_ (.A(_0534_),
    .B(_0569_),
    .Y(_0570_));
 sg13g2_a21oi_1 _2512_ (.A1(\levenshtein_ctrl.d[3] ),
    .A2(_0534_),
    .Y(_0571_),
    .B1(_0570_));
 sg13g2_inv_1 _2513_ (.Y(_0572_),
    .A(_0571_));
 sg13g2_nor2_1 _2514_ (.A(_0511_),
    .B(_0571_),
    .Y(_0573_));
 sg13g2_and2_1 _2515_ (.A(_0945_),
    .B(_0557_),
    .X(_0574_));
 sg13g2_xnor2_1 _2516_ (.Y(_0575_),
    .A(\levenshtein_ctrl.d[3] ),
    .B(_0557_));
 sg13g2_nor2_1 _2517_ (.A(_0510_),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_nor3_1 _2518_ (.A(_0532_),
    .B(_0573_),
    .C(_0576_),
    .Y(_0577_));
 sg13g2_nor2_2 _2519_ (.A(_0945_),
    .B(_0562_),
    .Y(_0578_));
 sg13g2_xnor2_1 _2520_ (.Y(_0579_),
    .A(\levenshtein_ctrl.d[3] ),
    .B(_0562_));
 sg13g2_o21ai_1 _2521_ (.B1(net381),
    .Y(_0580_),
    .A1(_0531_),
    .A2(_0579_));
 sg13g2_a221oi_1 _2522_ (.B2(_0569_),
    .C1(_1006_),
    .B1(net347),
    .A1(_0945_),
    .Y(_0581_),
    .A2(_1040_));
 sg13g2_a221oi_1 _2523_ (.B2(_0572_),
    .C1(_0581_),
    .B1(_1284_),
    .A1(\levenshtein_ctrl.d[3] ),
    .Y(_0582_),
    .A2(net429));
 sg13g2_o21ai_1 _2524_ (.B1(_0582_),
    .Y(_0156_),
    .A1(_0577_),
    .A2(_0580_));
 sg13g2_and2_1 _2525_ (.A(_0947_),
    .B(_0574_),
    .X(_0583_));
 sg13g2_nor2_1 _2526_ (.A(_0947_),
    .B(_0574_),
    .Y(_0584_));
 sg13g2_or3_1 _2527_ (.A(_0510_),
    .B(_0583_),
    .C(_0584_),
    .X(_0585_));
 sg13g2_a21o_1 _2528_ (.A2(net344),
    .A1(\levenshtein_ctrl.d[4] ),
    .B1(_0447_),
    .X(_0586_));
 sg13g2_mux2_1 _2529_ (.A0(_0947_),
    .A1(_0445_),
    .S(_0535_),
    .X(_0587_));
 sg13g2_a221oi_1 _2530_ (.B2(_0510_),
    .C1(_0530_),
    .B1(_0587_),
    .A1(_0444_),
    .Y(_0588_),
    .A2(_0513_));
 sg13g2_xnor2_1 _2531_ (.Y(_0589_),
    .A(_0947_),
    .B(_0578_));
 sg13g2_a22oi_1 _2532_ (.Y(_0590_),
    .B1(_0589_),
    .B2(_0532_),
    .A2(_0588_),
    .A1(_0585_));
 sg13g2_nor2_1 _2533_ (.A(_1285_),
    .B(_0587_),
    .Y(_0591_));
 sg13g2_a221oi_1 _2534_ (.B2(_0586_),
    .C1(_0591_),
    .B1(net395),
    .A1(net748),
    .Y(_0592_),
    .A2(net429));
 sg13g2_o21ai_1 _2535_ (.B1(_0592_),
    .Y(_0157_),
    .A1(net379),
    .A2(_0590_));
 sg13g2_nand2_1 _2536_ (.Y(_0593_),
    .A(net638),
    .B(net334));
 sg13g2_nor2_1 _2537_ (.A(_0511_),
    .B(_0535_),
    .Y(_0594_));
 sg13g2_and2_1 _2538_ (.A(_0949_),
    .B(_0583_),
    .X(_0595_));
 sg13g2_xnor2_1 _2539_ (.Y(_0596_),
    .A(_0949_),
    .B(_0583_));
 sg13g2_a221oi_1 _2540_ (.B2(_0511_),
    .C1(_0532_),
    .B1(_0596_),
    .A1(net638),
    .Y(_0597_),
    .A2(_0594_));
 sg13g2_nand3_1 _2541_ (.B(\levenshtein_ctrl.d[5] ),
    .C(_0578_),
    .A(\levenshtein_ctrl.d[4] ),
    .Y(_0598_));
 sg13g2_a21o_1 _2542_ (.A2(_0578_),
    .A1(\levenshtein_ctrl.d[4] ),
    .B1(\levenshtein_ctrl.d[5] ),
    .X(_0599_));
 sg13g2_and2_1 _2543_ (.A(_0598_),
    .B(_0599_),
    .X(_0600_));
 sg13g2_o21ai_1 _2544_ (.B1(net380),
    .Y(_0601_),
    .A1(_0531_),
    .A2(_0600_));
 sg13g2_o21ai_1 _2545_ (.B1(_0593_),
    .Y(_0158_),
    .A1(_0597_),
    .A2(_0601_));
 sg13g2_nand2_1 _2546_ (.Y(_0602_),
    .A(net647),
    .B(net334));
 sg13g2_and2_1 _2547_ (.A(_0951_),
    .B(_0595_),
    .X(_0603_));
 sg13g2_xnor2_1 _2548_ (.Y(_0604_),
    .A(_0951_),
    .B(_0595_));
 sg13g2_a221oi_1 _2549_ (.B2(_0511_),
    .C1(_0532_),
    .B1(_0604_),
    .A1(net647),
    .Y(_0605_),
    .A2(_0594_));
 sg13g2_or2_1 _2550_ (.X(_0606_),
    .B(_0598_),
    .A(_0951_));
 sg13g2_xnor2_1 _2551_ (.Y(_0607_),
    .A(\levenshtein_ctrl.d[6] ),
    .B(_0598_));
 sg13g2_o21ai_1 _2552_ (.B1(net380),
    .Y(_0608_),
    .A1(_0531_),
    .A2(_0607_));
 sg13g2_o21ai_1 _2553_ (.B1(_0602_),
    .Y(_0159_),
    .A1(_0605_),
    .A2(_0608_));
 sg13g2_nand2_1 _2554_ (.Y(_0609_),
    .A(net576),
    .B(net334));
 sg13g2_xnor2_1 _2555_ (.Y(_0610_),
    .A(_0953_),
    .B(_0603_));
 sg13g2_a221oi_1 _2556_ (.B2(_0511_),
    .C1(_0532_),
    .B1(_0610_),
    .A1(net576),
    .Y(_0611_),
    .A2(_0594_));
 sg13g2_xnor2_1 _2557_ (.Y(_0612_),
    .A(\levenshtein_ctrl.d[7] ),
    .B(_0606_));
 sg13g2_o21ai_1 _2558_ (.B1(net380),
    .Y(_0613_),
    .A1(_0531_),
    .A2(_0612_));
 sg13g2_o21ai_1 _2559_ (.B1(_0609_),
    .Y(_0160_),
    .A1(_0611_),
    .A2(_0613_));
 sg13g2_nor3_1 _2560_ (.A(_0986_),
    .B(_1028_),
    .C(_1082_),
    .Y(_0614_));
 sg13g2_a21o_1 _2561_ (.A2(_1036_),
    .A1(net265),
    .B1(_0614_),
    .X(_0161_));
 sg13g2_a22oi_1 _2562_ (.Y(_0615_),
    .B1(net355),
    .B2(net590),
    .A2(_1036_),
    .A1(\levenshtein_ctrl.idx[0] ));
 sg13g2_and4_1 _2563_ (.A(\levenshtein_ctrl.idx[0] ),
    .B(\levenshtein_ctrl.idx[1] ),
    .C(net397),
    .D(_1026_),
    .X(_0616_));
 sg13g2_and3_1 _2564_ (.X(_0617_),
    .A(\levenshtein_ctrl.idx[0] ),
    .B(net590),
    .C(_1036_));
 sg13g2_nor2_1 _2565_ (.A(net591),
    .B(_0617_),
    .Y(_0162_));
 sg13g2_a21oi_1 _2566_ (.A1(net493),
    .A2(net355),
    .Y(_0618_),
    .B1(_0617_));
 sg13g2_a21oi_1 _2567_ (.A1(net493),
    .A2(_0617_),
    .Y(_0163_),
    .B1(_0618_));
 sg13g2_a22oi_1 _2568_ (.Y(_0619_),
    .B1(_0617_),
    .B2(net493),
    .A2(net355),
    .A1(net522));
 sg13g2_nand3_1 _2569_ (.B(net522),
    .C(_0616_),
    .A(net493),
    .Y(_0620_));
 sg13g2_nor2b_1 _2570_ (.A(net523),
    .B_N(_0620_),
    .Y(_0164_));
 sg13g2_nand2_1 _2571_ (.Y(_0621_),
    .A(net520),
    .B(net353));
 sg13g2_nor2_1 _2572_ (.A(_0987_),
    .B(_0620_),
    .Y(_0622_));
 sg13g2_xor2_1 _2573_ (.B(_0621_),
    .A(_0620_),
    .X(_0165_));
 sg13g2_nand2_1 _2574_ (.Y(_0623_),
    .A(net595),
    .B(net353));
 sg13g2_nor3_1 _2575_ (.A(_0987_),
    .B(_0620_),
    .C(_0623_),
    .Y(_0624_));
 sg13g2_xnor2_1 _2576_ (.Y(_0166_),
    .A(_0622_),
    .B(_0623_));
 sg13g2_a21oi_1 _2577_ (.A1(net555),
    .A2(net353),
    .Y(_0625_),
    .B1(_0624_));
 sg13g2_and4_1 _2578_ (.A(\levenshtein_ctrl.idx[5] ),
    .B(net555),
    .C(net353),
    .D(_0622_),
    .X(_0626_));
 sg13g2_nor2_1 _2579_ (.A(net556),
    .B(_0626_),
    .Y(_0167_));
 sg13g2_nand2_1 _2580_ (.Y(_0627_),
    .A(net518),
    .B(net353));
 sg13g2_and2_1 _2581_ (.A(net518),
    .B(_0626_),
    .X(_0628_));
 sg13g2_xnor2_1 _2582_ (.Y(_0168_),
    .A(_0626_),
    .B(_0627_));
 sg13g2_nand2_1 _2583_ (.Y(_0629_),
    .A(net573),
    .B(net353));
 sg13g2_xnor2_1 _2584_ (.Y(_0169_),
    .A(_0628_),
    .B(_0629_));
 sg13g2_and2_1 _2585_ (.A(\levenshtein_ctrl.idx[9] ),
    .B(net354),
    .X(_0630_));
 sg13g2_a21oi_1 _2586_ (.A1(net573),
    .A2(_0628_),
    .Y(_0631_),
    .B1(_0630_));
 sg13g2_nand3_1 _2587_ (.B(\levenshtein_ctrl.idx[9] ),
    .C(_0628_),
    .A(net573),
    .Y(_0632_));
 sg13g2_nor2b_1 _2588_ (.A(net574),
    .B_N(_0632_),
    .Y(_0170_));
 sg13g2_nand2_1 _2589_ (.Y(_0633_),
    .A(net529),
    .B(net354));
 sg13g2_nor2_1 _2590_ (.A(_0632_),
    .B(_0633_),
    .Y(_0634_));
 sg13g2_xor2_1 _2591_ (.B(_0633_),
    .A(_0632_),
    .X(_0171_));
 sg13g2_a21oi_1 _2592_ (.A1(net684),
    .A2(net354),
    .Y(_0635_),
    .B1(_0634_));
 sg13g2_and2_1 _2593_ (.A(net684),
    .B(_0634_),
    .X(_0636_));
 sg13g2_nor2_1 _2594_ (.A(net685),
    .B(_0636_),
    .Y(_0172_));
 sg13g2_a21oi_1 _2595_ (.A1(net669),
    .A2(net353),
    .Y(_0637_),
    .B1(_0636_));
 sg13g2_nand2_1 _2596_ (.Y(_0638_),
    .A(net669),
    .B(_0636_));
 sg13g2_nor2b_1 _2597_ (.A(net670),
    .B_N(_0638_),
    .Y(_0173_));
 sg13g2_nand2_1 _2598_ (.Y(_0639_),
    .A(net600),
    .B(net353));
 sg13g2_nand4_1 _2599_ (.B(net669),
    .C(net600),
    .A(net684),
    .Y(_0640_),
    .D(_0634_));
 sg13g2_xor2_1 _2600_ (.B(_0639_),
    .A(_0638_),
    .X(_0174_));
 sg13g2_nand2_1 _2601_ (.Y(_0641_),
    .A(net707),
    .B(net354));
 sg13g2_nand4_1 _2602_ (.B(\levenshtein_ctrl.idx[13] ),
    .C(\levenshtein_ctrl.idx[14] ),
    .A(\levenshtein_ctrl.idx[12] ),
    .Y(_0642_),
    .D(_0636_));
 sg13g2_mux2_1 _2603_ (.A0(net707),
    .A1(_0641_),
    .S(_0640_),
    .X(_0643_));
 sg13g2_inv_1 _2604_ (.Y(_0175_),
    .A(_0643_));
 sg13g2_nand2_1 _2605_ (.Y(_0644_),
    .A(net498),
    .B(net354));
 sg13g2_xor2_1 _2606_ (.B(_0644_),
    .A(_0642_),
    .X(_0176_));
 sg13g2_nand2_1 _2607_ (.Y(_0645_),
    .A(net428),
    .B(net464));
 sg13g2_nand2_1 _2608_ (.Y(_0646_),
    .A(\levenshtein_ctrl.best_distance[2] ),
    .B(_0943_));
 sg13g2_a22oi_1 _2609_ (.Y(_0647_),
    .B1(\levenshtein_ctrl.best_distance[1] ),
    .B2(_0941_),
    .A2(_0939_),
    .A1(\levenshtein_ctrl.best_distance[0] ));
 sg13g2_a22oi_1 _2610_ (.Y(_0648_),
    .B1(_0942_),
    .B2(\levenshtein_ctrl.d[2] ),
    .A2(\levenshtein_ctrl.d[1] ),
    .A1(_0940_));
 sg13g2_nand2b_1 _2611_ (.Y(_0649_),
    .B(_0648_),
    .A_N(_0647_));
 sg13g2_a22oi_1 _2612_ (.Y(_0650_),
    .B1(_0646_),
    .B2(_0649_),
    .A2(\levenshtein_ctrl.d[3] ),
    .A1(_0944_));
 sg13g2_a221oi_1 _2613_ (.B2(_0947_),
    .C1(_0650_),
    .B1(\levenshtein_ctrl.best_distance[4] ),
    .A1(\levenshtein_ctrl.best_distance[3] ),
    .Y(_0651_),
    .A2(_0945_));
 sg13g2_a221oi_1 _2614_ (.B2(\levenshtein_ctrl.d[5] ),
    .C1(_0651_),
    .B1(_0948_),
    .A1(_0946_),
    .Y(_0652_),
    .A2(\levenshtein_ctrl.d[4] ));
 sg13g2_a221oi_1 _2615_ (.B2(_0951_),
    .C1(_0652_),
    .B1(\levenshtein_ctrl.best_distance[6] ),
    .A1(\levenshtein_ctrl.best_distance[5] ),
    .Y(_0653_),
    .A2(_0949_));
 sg13g2_a221oi_1 _2616_ (.B2(\levenshtein_ctrl.d[7] ),
    .C1(_0653_),
    .B1(_0952_),
    .A1(_0950_),
    .Y(_0654_),
    .A2(\levenshtein_ctrl.d[6] ));
 sg13g2_a21o_1 _2617_ (.A2(_0953_),
    .A1(\levenshtein_ctrl.best_distance[7] ),
    .B1(_0654_),
    .X(_0655_));
 sg13g2_nor2b_1 _2618_ (.A(_1263_),
    .B_N(_0655_),
    .Y(_0656_));
 sg13g2_nand2b_1 _2619_ (.Y(_0657_),
    .B(_0655_),
    .A_N(_1263_));
 sg13g2_a21oi_1 _2620_ (.A1(net464),
    .A2(net343),
    .Y(_0658_),
    .B1(net333));
 sg13g2_o21ai_1 _2621_ (.B1(net435),
    .Y(_0659_),
    .A1(\levenshtein_ctrl.idx[0] ),
    .A2(net330));
 sg13g2_o21ai_1 _2622_ (.B1(_0645_),
    .Y(_0177_),
    .A1(_0658_),
    .A2(_0659_));
 sg13g2_nand2_1 _2623_ (.Y(_0660_),
    .A(net532),
    .B(net428));
 sg13g2_a21oi_1 _2624_ (.A1(net532),
    .A2(net343),
    .Y(_0661_),
    .B1(net333));
 sg13g2_o21ai_1 _2625_ (.B1(net435),
    .Y(_0662_),
    .A1(\levenshtein_ctrl.idx[1] ),
    .A2(net330));
 sg13g2_o21ai_1 _2626_ (.B1(_0660_),
    .Y(_0178_),
    .A1(_0661_),
    .A2(_0662_));
 sg13g2_nand2_1 _2627_ (.Y(_0663_),
    .A(net302),
    .B(net426));
 sg13g2_a21oi_1 _2628_ (.A1(net302),
    .A2(net342),
    .Y(_0664_),
    .B1(net333));
 sg13g2_o21ai_1 _2629_ (.B1(net434),
    .Y(_0665_),
    .A1(\levenshtein_ctrl.idx[2] ),
    .A2(net330));
 sg13g2_o21ai_1 _2630_ (.B1(_0663_),
    .Y(_0179_),
    .A1(_0664_),
    .A2(_0665_));
 sg13g2_nand2_1 _2631_ (.Y(_0666_),
    .A(net560),
    .B(net428));
 sg13g2_a21oi_1 _2632_ (.A1(net560),
    .A2(net343),
    .Y(_0667_),
    .B1(net333));
 sg13g2_o21ai_1 _2633_ (.B1(net435),
    .Y(_0668_),
    .A1(net522),
    .A2(net330));
 sg13g2_o21ai_1 _2634_ (.B1(_0666_),
    .Y(_0180_),
    .A1(_0667_),
    .A2(_0668_));
 sg13g2_nand2_1 _2635_ (.Y(_0669_),
    .A(net310),
    .B(net426));
 sg13g2_a21oi_1 _2636_ (.A1(net310),
    .A2(net342),
    .Y(_0670_),
    .B1(net332));
 sg13g2_o21ai_1 _2637_ (.B1(net432),
    .Y(_0671_),
    .A1(\levenshtein_ctrl.idx[4] ),
    .A2(net329));
 sg13g2_o21ai_1 _2638_ (.B1(_0669_),
    .Y(_0181_),
    .A1(_0670_),
    .A2(_0671_));
 sg13g2_nand2_1 _2639_ (.Y(_0672_),
    .A(net475),
    .B(net426));
 sg13g2_a21oi_1 _2640_ (.A1(net475),
    .A2(net341),
    .Y(_0673_),
    .B1(net331));
 sg13g2_o21ai_1 _2641_ (.B1(net432),
    .Y(_0674_),
    .A1(\levenshtein_ctrl.idx[5] ),
    .A2(net329));
 sg13g2_o21ai_1 _2642_ (.B1(_0672_),
    .Y(_0182_),
    .A1(_0673_),
    .A2(_0674_));
 sg13g2_nand2_1 _2643_ (.Y(_0675_),
    .A(net306),
    .B(net426));
 sg13g2_a21oi_1 _2644_ (.A1(net306),
    .A2(net341),
    .Y(_0676_),
    .B1(net331));
 sg13g2_o21ai_1 _2645_ (.B1(net432),
    .Y(_0677_),
    .A1(\levenshtein_ctrl.idx[6] ),
    .A2(net328));
 sg13g2_o21ai_1 _2646_ (.B1(_0675_),
    .Y(_0183_),
    .A1(_0676_),
    .A2(_0677_));
 sg13g2_nand2_1 _2647_ (.Y(_0678_),
    .A(net304),
    .B(net426));
 sg13g2_a21oi_1 _2648_ (.A1(net304),
    .A2(net341),
    .Y(_0679_),
    .B1(net331));
 sg13g2_o21ai_1 _2649_ (.B1(net432),
    .Y(_0680_),
    .A1(\levenshtein_ctrl.idx[7] ),
    .A2(net328));
 sg13g2_o21ai_1 _2650_ (.B1(_0678_),
    .Y(_0184_),
    .A1(_0679_),
    .A2(_0680_));
 sg13g2_nand2_1 _2651_ (.Y(_0681_),
    .A(net580),
    .B(net426));
 sg13g2_a21oi_1 _2652_ (.A1(net580),
    .A2(net341),
    .Y(_0682_),
    .B1(net332));
 sg13g2_o21ai_1 _2653_ (.B1(net432),
    .Y(_0683_),
    .A1(net573),
    .A2(net328));
 sg13g2_o21ai_1 _2654_ (.B1(_0681_),
    .Y(_0185_),
    .A1(_0682_),
    .A2(_0683_));
 sg13g2_nand2_1 _2655_ (.Y(_0684_),
    .A(net699),
    .B(net426));
 sg13g2_a21oi_1 _2656_ (.A1(net699),
    .A2(net341),
    .Y(_0685_),
    .B1(net331));
 sg13g2_o21ai_1 _2657_ (.B1(net432),
    .Y(_0686_),
    .A1(\levenshtein_ctrl.idx[9] ),
    .A2(net328));
 sg13g2_o21ai_1 _2658_ (.B1(_0684_),
    .Y(_0186_),
    .A1(_0685_),
    .A2(_0686_));
 sg13g2_nand2_1 _2659_ (.Y(_0687_),
    .A(net644),
    .B(net426));
 sg13g2_a21oi_1 _2660_ (.A1(net644),
    .A2(net341),
    .Y(_0688_),
    .B1(net331));
 sg13g2_o21ai_1 _2661_ (.B1(net432),
    .Y(_0689_),
    .A1(net529),
    .A2(net328));
 sg13g2_o21ai_1 _2662_ (.B1(_0687_),
    .Y(_0187_),
    .A1(_0688_),
    .A2(_0689_));
 sg13g2_nand2_1 _2663_ (.Y(_0690_),
    .A(net714),
    .B(net427));
 sg13g2_a21oi_1 _2664_ (.A1(net714),
    .A2(net342),
    .Y(_0691_),
    .B1(net331));
 sg13g2_o21ai_1 _2665_ (.B1(net433),
    .Y(_0692_),
    .A1(net684),
    .A2(net329));
 sg13g2_o21ai_1 _2666_ (.B1(_0690_),
    .Y(_0188_),
    .A1(_0691_),
    .A2(_0692_));
 sg13g2_nand2_1 _2667_ (.Y(_0693_),
    .A(net525),
    .B(net427));
 sg13g2_a21oi_1 _2668_ (.A1(net525),
    .A2(net342),
    .Y(_0694_),
    .B1(net332));
 sg13g2_o21ai_1 _2669_ (.B1(net433),
    .Y(_0695_),
    .A1(\levenshtein_ctrl.idx[12] ),
    .A2(net329));
 sg13g2_o21ai_1 _2670_ (.B1(_0693_),
    .Y(_0189_),
    .A1(_0694_),
    .A2(_0695_));
 sg13g2_nand2_1 _2671_ (.Y(_0696_),
    .A(net471),
    .B(net427));
 sg13g2_a21oi_1 _2672_ (.A1(net471),
    .A2(net341),
    .Y(_0697_),
    .B1(net332));
 sg13g2_o21ai_1 _2673_ (.B1(net433),
    .Y(_0698_),
    .A1(\levenshtein_ctrl.idx[13] ),
    .A2(net328));
 sg13g2_o21ai_1 _2674_ (.B1(_0696_),
    .Y(_0190_),
    .A1(_0697_),
    .A2(_0698_));
 sg13g2_nand2_1 _2675_ (.Y(_0699_),
    .A(net491),
    .B(net427));
 sg13g2_a21oi_1 _2676_ (.A1(net491),
    .A2(net342),
    .Y(_0700_),
    .B1(net331));
 sg13g2_o21ai_1 _2677_ (.B1(net433),
    .Y(_0701_),
    .A1(\levenshtein_ctrl.idx[14] ),
    .A2(net328));
 sg13g2_o21ai_1 _2678_ (.B1(_0699_),
    .Y(_0191_),
    .A1(_0700_),
    .A2(_0701_));
 sg13g2_nand2_1 _2679_ (.Y(_0702_),
    .A(net473),
    .B(net427));
 sg13g2_a21oi_1 _2680_ (.A1(net473),
    .A2(net341),
    .Y(_0703_),
    .B1(net331));
 sg13g2_o21ai_1 _2681_ (.B1(net432),
    .Y(_0704_),
    .A1(\levenshtein_ctrl.idx[15] ),
    .A2(net328));
 sg13g2_o21ai_1 _2682_ (.B1(_0702_),
    .Y(_0192_),
    .A1(_0703_),
    .A2(_0704_));
 sg13g2_and4_2 _2683_ (.A(net435),
    .B(_1024_),
    .C(_1033_),
    .D(_0655_),
    .X(_0705_));
 sg13g2_nor2_2 _2684_ (.A(_1082_),
    .B(_0705_),
    .Y(_0706_));
 sg13g2_a22oi_1 _2685_ (.Y(_0193_),
    .B1(_0706_),
    .B2(_0938_),
    .A2(_0705_),
    .A1(_0939_));
 sg13g2_a22oi_1 _2686_ (.Y(_0194_),
    .B1(_0706_),
    .B2(_0940_),
    .A2(_0705_),
    .A1(_0941_));
 sg13g2_a22oi_1 _2687_ (.Y(_0195_),
    .B1(_0706_),
    .B2(_0942_),
    .A2(_0705_),
    .A1(_0943_));
 sg13g2_a22oi_1 _2688_ (.Y(_0196_),
    .B1(_0706_),
    .B2(_0944_),
    .A2(_0705_),
    .A1(_0945_));
 sg13g2_a22oi_1 _2689_ (.Y(_0197_),
    .B1(_0706_),
    .B2(_0946_),
    .A2(_0705_),
    .A1(_0947_));
 sg13g2_a22oi_1 _2690_ (.Y(_0198_),
    .B1(_0706_),
    .B2(_0948_),
    .A2(_0705_),
    .A1(_0949_));
 sg13g2_a22oi_1 _2691_ (.Y(_0199_),
    .B1(_0706_),
    .B2(_0950_),
    .A2(_0705_),
    .A1(_0951_));
 sg13g2_a22oi_1 _2692_ (.Y(_0200_),
    .B1(net355),
    .B2(_0952_),
    .A2(_1036_),
    .A1(_0953_));
 sg13g2_a21oi_1 _2693_ (.A1(\arbiter.wbs1_cyc_i ),
    .A2(net425),
    .Y(_0707_),
    .B1(net391));
 sg13g2_inv_1 _2694_ (.Y(_0708_),
    .A(_0707_));
 sg13g2_a22oi_1 _2695_ (.Y(_0709_),
    .B1(_1041_),
    .B2(_0708_),
    .A2(net396),
    .A1(\levenshtein_ctrl.state[1] ));
 sg13g2_mux2_1 _2696_ (.A0(net443),
    .A1(\levenshtein_ctrl.next_symbol[0] ),
    .S(net363),
    .X(_0201_));
 sg13g2_mux2_1 _2697_ (.A0(net451),
    .A1(net453),
    .S(net360),
    .X(_0202_));
 sg13g2_mux2_1 _2698_ (.A0(net316),
    .A1(net487),
    .S(net360),
    .X(_0203_));
 sg13g2_mux2_1 _2699_ (.A0(net445),
    .A1(\levenshtein_ctrl.next_symbol[3] ),
    .S(net364),
    .X(_0204_));
 sg13g2_mux2_1 _2700_ (.A0(net454),
    .A1(net458),
    .S(net365),
    .X(_0205_));
 sg13g2_mux2_1 _2701_ (.A0(net459),
    .A1(net490),
    .S(net362),
    .X(_0206_));
 sg13g2_mux2_1 _2702_ (.A0(net327),
    .A1(net480),
    .S(net361),
    .X(_0207_));
 sg13g2_mux2_1 _2703_ (.A0(net470),
    .A1(net484),
    .S(net362),
    .X(_0208_));
 sg13g2_mux2_1 _2704_ (.A0(net295),
    .A1(net443),
    .S(net363),
    .X(_0209_));
 sg13g2_mux2_1 _2705_ (.A0(net281),
    .A1(net451),
    .S(net360),
    .X(_0210_));
 sg13g2_mux2_1 _2706_ (.A0(net273),
    .A1(net316),
    .S(net360),
    .X(_0211_));
 sg13g2_mux2_1 _2707_ (.A0(net477),
    .A1(net445),
    .S(net364),
    .X(_0212_));
 sg13g2_mux2_1 _2708_ (.A0(net271),
    .A1(net454),
    .S(net361),
    .X(_0213_));
 sg13g2_mux2_1 _2709_ (.A0(net290),
    .A1(net459),
    .S(net362),
    .X(_0214_));
 sg13g2_mux2_1 _2710_ (.A0(net277),
    .A1(net327),
    .S(net361),
    .X(_0215_));
 sg13g2_mux2_1 _2711_ (.A0(net275),
    .A1(net470),
    .S(net362),
    .X(_0216_));
 sg13g2_nand2_1 _2712_ (.Y(_0710_),
    .A(net295),
    .B(net363));
 sg13g2_o21ai_1 _2713_ (.B1(_0710_),
    .Y(_0217_),
    .A1(_0956_),
    .A2(net363));
 sg13g2_nand2_1 _2714_ (.Y(_0711_),
    .A(net281),
    .B(net360));
 sg13g2_o21ai_1 _2715_ (.B1(_0711_),
    .Y(_0218_),
    .A1(_0957_),
    .A2(net360));
 sg13g2_nand2_1 _2716_ (.Y(_0712_),
    .A(net273),
    .B(net360));
 sg13g2_o21ai_1 _2717_ (.B1(_0712_),
    .Y(_0219_),
    .A1(_0958_),
    .A2(net360));
 sg13g2_mux2_1 _2718_ (.A0(net312),
    .A1(\levenshtein_ctrl.symbols[19] ),
    .S(net363),
    .X(_0220_));
 sg13g2_nand2_1 _2719_ (.Y(_0713_),
    .A(net271),
    .B(net361));
 sg13g2_o21ai_1 _2720_ (.B1(_0713_),
    .Y(_0221_),
    .A1(_0959_),
    .A2(net361));
 sg13g2_nand2_1 _2721_ (.Y(_0714_),
    .A(net290),
    .B(net364));
 sg13g2_o21ai_1 _2722_ (.B1(_0714_),
    .Y(_0222_),
    .A1(_0960_),
    .A2(net364));
 sg13g2_nand2_1 _2723_ (.Y(_0715_),
    .A(net277),
    .B(net361));
 sg13g2_o21ai_1 _2724_ (.B1(_0715_),
    .Y(_0223_),
    .A1(_0961_),
    .A2(net361));
 sg13g2_nand2_1 _2725_ (.Y(_0716_),
    .A(net275),
    .B(net364));
 sg13g2_o21ai_1 _2726_ (.B1(_0716_),
    .Y(_0224_),
    .A1(_0962_),
    .A2(net362));
 sg13g2_nor3_2 _2727_ (.A(net423),
    .B(_1042_),
    .C(_0707_),
    .Y(_0717_));
 sg13g2_nand2b_1 _2728_ (.Y(_0718_),
    .B(_0717_),
    .A_N(\arbiter.wbm_dat_i[0] ));
 sg13g2_o21ai_1 _2729_ (.B1(_0718_),
    .Y(_0719_),
    .A1(\levenshtein_ctrl.next_symbol[0] ),
    .A2(_1035_));
 sg13g2_a21oi_1 _2730_ (.A1(_0956_),
    .A2(net364),
    .Y(_0225_),
    .B1(_0719_));
 sg13g2_nand2b_1 _2731_ (.Y(_0720_),
    .B(_0717_),
    .A_N(\arbiter.wbm_dat_i[1] ));
 sg13g2_o21ai_1 _2732_ (.B1(_0720_),
    .Y(_0721_),
    .A1(net453),
    .A2(_1035_));
 sg13g2_a21oi_1 _2733_ (.A1(_0957_),
    .A2(net363),
    .Y(_0226_),
    .B1(_0721_));
 sg13g2_nand2b_1 _2734_ (.Y(_0722_),
    .B(_0717_),
    .A_N(\arbiter.wbm_dat_i[2] ));
 sg13g2_o21ai_1 _2735_ (.B1(_0722_),
    .Y(_0723_),
    .A1(net487),
    .A2(_1035_));
 sg13g2_a21oi_1 _2736_ (.A1(_0958_),
    .A2(net363),
    .Y(_0227_),
    .B1(_0723_));
 sg13g2_nand2b_1 _2737_ (.Y(_0724_),
    .B(net363),
    .A_N(net312));
 sg13g2_o21ai_1 _2738_ (.B1(_0724_),
    .Y(_0725_),
    .A1(net691),
    .A2(_1035_));
 sg13g2_a21oi_1 _2739_ (.A1(_0963_),
    .A2(_0717_),
    .Y(_0228_),
    .B1(_0725_));
 sg13g2_nand2b_1 _2740_ (.Y(_0726_),
    .B(_0717_),
    .A_N(\arbiter.wbm_dat_i[4] ));
 sg13g2_o21ai_1 _2741_ (.B1(_0726_),
    .Y(_0727_),
    .A1(\levenshtein_ctrl.next_symbol[4] ),
    .A2(_1035_));
 sg13g2_a21oi_1 _2742_ (.A1(_0959_),
    .A2(net365),
    .Y(_0229_),
    .B1(_0727_));
 sg13g2_nand2b_1 _2743_ (.Y(_0728_),
    .B(_0717_),
    .A_N(\arbiter.wbm_dat_i[5] ));
 sg13g2_o21ai_1 _2744_ (.B1(_0728_),
    .Y(_0729_),
    .A1(\levenshtein_ctrl.next_symbol[5] ),
    .A2(_1035_));
 sg13g2_a21oi_1 _2745_ (.A1(_0960_),
    .A2(net362),
    .Y(_0230_),
    .B1(_0729_));
 sg13g2_nand2b_1 _2746_ (.Y(_0730_),
    .B(_0717_),
    .A_N(\arbiter.wbm_dat_i[6] ));
 sg13g2_o21ai_1 _2747_ (.B1(_0730_),
    .Y(_0731_),
    .A1(\levenshtein_ctrl.next_symbol[6] ),
    .A2(_1035_));
 sg13g2_a21oi_1 _2748_ (.A1(_0961_),
    .A2(net362),
    .Y(_0231_),
    .B1(_0731_));
 sg13g2_nand2b_1 _2749_ (.Y(_0732_),
    .B(_0717_),
    .A_N(\arbiter.wbm_dat_i[7] ));
 sg13g2_o21ai_1 _2750_ (.B1(_0732_),
    .Y(_0733_),
    .A1(\levenshtein_ctrl.next_symbol[7] ),
    .A2(_1035_));
 sg13g2_a21oi_1 _2751_ (.A1(_0962_),
    .A2(net362),
    .Y(_0232_),
    .B1(_0733_));
 sg13g2_and4_1 _2752_ (.A(\arbiter.wbs1_cyc_i ),
    .B(\levenshtein_ctrl.state[3] ),
    .C(net396),
    .D(net394),
    .X(_0734_));
 sg13g2_mux2_1 _2753_ (.A0(net679),
    .A1(\arbiter.wbm_dat_i[0] ),
    .S(net377),
    .X(_0233_));
 sg13g2_mux2_1 _2754_ (.A0(net549),
    .A1(\arbiter.wbm_dat_i[1] ),
    .S(net377),
    .X(_0234_));
 sg13g2_mux2_1 _2755_ (.A0(net658),
    .A1(\arbiter.wbm_dat_i[2] ),
    .S(net377),
    .X(_0235_));
 sg13g2_nor2_1 _2756_ (.A(net585),
    .B(_0734_),
    .Y(_0735_));
 sg13g2_a21oi_1 _2757_ (.A1(_0963_),
    .A2(net377),
    .Y(_0236_),
    .B1(net586));
 sg13g2_mux2_1 _2758_ (.A0(net630),
    .A1(\arbiter.wbm_dat_i[4] ),
    .S(net377),
    .X(_0237_));
 sg13g2_mux2_1 _2759_ (.A0(net488),
    .A1(\arbiter.wbm_dat_i[5] ),
    .S(net377),
    .X(_0238_));
 sg13g2_mux2_1 _2760_ (.A0(net460),
    .A1(\arbiter.wbm_dat_i[6] ),
    .S(net377),
    .X(_0239_));
 sg13g2_mux2_1 _2761_ (.A0(net326),
    .A1(\arbiter.wbm_dat_i[7] ),
    .S(net377),
    .X(_0240_));
 sg13g2_a221oi_1 _2762_ (.B2(_1058_),
    .C1(net393),
    .B1(_1088_),
    .A1(_0935_),
    .Y(_0736_),
    .A2(_1065_));
 sg13g2_nor2_1 _2763_ (.A(net662),
    .B(net338),
    .Y(_0737_));
 sg13g2_nand2b_2 _2764_ (.Y(_0738_),
    .B(\spi.state[2] ),
    .A_N(\spi.state[0] ));
 sg13g2_and2_2 _2765_ (.A(\arbiter.wbs0_adr_i[2] ),
    .B(_1002_),
    .X(_0739_));
 sg13g2_and2_2 _2766_ (.A(_0967_),
    .B(_1211_),
    .X(_0740_));
 sg13g2_nor3_2 _2767_ (.A(_0936_),
    .B(\arbiter.wbs0_adr_i[1] ),
    .C(_0018_),
    .Y(_0741_));
 sg13g2_a22oi_1 _2768_ (.Y(_0742_),
    .B1(_0740_),
    .B2(\levenshtein_ctrl.best_distance[1] ),
    .A2(_1212_),
    .A1(net415));
 sg13g2_and3_1 _2769_ (.X(_0743_),
    .A(\arbiter.wbs0_adr_i[0] ),
    .B(\arbiter.wbs0_adr_i[1] ),
    .C(_0018_));
 sg13g2_a21oi_1 _2770_ (.A1(\levenshtein_ctrl.best_idx[9] ),
    .A2(_0739_),
    .Y(_0744_),
    .B1(_0743_));
 sg13g2_a22oi_1 _2771_ (.Y(_0745_),
    .B1(_0741_),
    .B2(\levenshtein_ctrl.best_idx[1] ),
    .A2(_1203_),
    .A1(\levenshtein_ctrl.sram_config[1] ));
 sg13g2_nand4_1 _2772_ (.B(_0742_),
    .C(_0744_),
    .A(net371),
    .Y(_0746_),
    .D(_0745_));
 sg13g2_nor2_2 _2773_ (.A(net641),
    .B(_1085_),
    .Y(_0747_));
 sg13g2_o21ai_1 _2774_ (.B1(_0747_),
    .Y(_0748_),
    .A1(\arbiter.wbm_dat_i[1] ),
    .A2(net368));
 sg13g2_inv_1 _2775_ (.Y(_0749_),
    .A(_0748_));
 sg13g2_a22oi_1 _2776_ (.Y(_0750_),
    .B1(_0746_),
    .B2(_0749_),
    .A2(_0738_),
    .A1(\arbiter.wbs0_dat_i[0] ));
 sg13g2_a21oi_1 _2777_ (.A1(net338),
    .A2(_0750_),
    .Y(_0241_),
    .B1(_0737_));
 sg13g2_nor2_1 _2778_ (.A(net628),
    .B(net338),
    .Y(_0751_));
 sg13g2_a22oi_1 _2779_ (.Y(_0752_),
    .B1(_0741_),
    .B2(\levenshtein_ctrl.best_idx[2] ),
    .A2(_0739_),
    .A1(\levenshtein_ctrl.best_idx[10] ));
 sg13g2_a221oi_1 _2780_ (.B2(\levenshtein_ctrl.best_distance[2] ),
    .C1(_0743_),
    .B1(_0740_),
    .A1(net413),
    .Y(_0753_),
    .A2(_1212_));
 sg13g2_nand3_1 _2781_ (.B(_0752_),
    .C(_0753_),
    .A(net371),
    .Y(_0754_));
 sg13g2_o21ai_1 _2782_ (.B1(_0747_),
    .Y(_0755_),
    .A1(\arbiter.wbm_dat_i[2] ),
    .A2(net368));
 sg13g2_inv_1 _2783_ (.Y(_0756_),
    .A(_0755_));
 sg13g2_a22oi_1 _2784_ (.Y(_0757_),
    .B1(_0754_),
    .B2(_0756_),
    .A2(_0738_),
    .A1(\arbiter.wbs0_dat_i[1] ));
 sg13g2_a21oi_1 _2785_ (.A1(net338),
    .A2(_0757_),
    .Y(_0242_),
    .B1(_0751_));
 sg13g2_nor2_1 _2786_ (.A(net650),
    .B(net338),
    .Y(_0758_));
 sg13g2_a22oi_1 _2787_ (.Y(_0759_),
    .B1(_0741_),
    .B2(\levenshtein_ctrl.best_idx[3] ),
    .A2(_1212_),
    .A1(net411));
 sg13g2_a221oi_1 _2788_ (.B2(\levenshtein_ctrl.best_distance[3] ),
    .C1(_0743_),
    .B1(_0740_),
    .A1(\levenshtein_ctrl.best_idx[11] ),
    .Y(_0760_),
    .A2(_0739_));
 sg13g2_nand3_1 _2789_ (.B(_0759_),
    .C(_0760_),
    .A(net371),
    .Y(_0761_));
 sg13g2_o21ai_1 _2790_ (.B1(_0747_),
    .Y(_0762_),
    .A1(net661),
    .A2(net369));
 sg13g2_inv_1 _2791_ (.Y(_0763_),
    .A(_0762_));
 sg13g2_a22oi_1 _2792_ (.Y(_0764_),
    .B1(_0761_),
    .B2(_0763_),
    .A2(_0738_),
    .A1(net628));
 sg13g2_a21oi_1 _2793_ (.A1(net338),
    .A2(_0764_),
    .Y(_0243_),
    .B1(_0758_));
 sg13g2_and2_1 _2794_ (.A(\levenshtein_ctrl.best_idx[12] ),
    .B(_0739_),
    .X(_0765_));
 sg13g2_a221oi_1 _2795_ (.B2(\levenshtein_ctrl.best_idx[4] ),
    .C1(_0765_),
    .B1(_0741_),
    .A1(\levenshtein_ctrl.best_distance[4] ),
    .Y(_0766_),
    .A2(_0740_));
 sg13g2_o21ai_1 _2796_ (.B1(_0747_),
    .Y(_0767_),
    .A1(\arbiter.wbm_dat_i[4] ),
    .A2(net368));
 sg13g2_a21oi_1 _2797_ (.A1(net370),
    .A2(_0766_),
    .Y(_0768_),
    .B1(_0767_));
 sg13g2_a21oi_1 _2798_ (.A1(\arbiter.wbs0_dat_i[3] ),
    .A2(_0738_),
    .Y(_0769_),
    .B1(_0768_));
 sg13g2_nor2_1 _2799_ (.A(net506),
    .B(net340),
    .Y(_0770_));
 sg13g2_a21oi_1 _2800_ (.A1(net338),
    .A2(_0769_),
    .Y(_0244_),
    .B1(_0770_));
 sg13g2_and2_1 _2801_ (.A(\levenshtein_ctrl.best_idx[13] ),
    .B(_0739_),
    .X(_0771_));
 sg13g2_a221oi_1 _2802_ (.B2(\levenshtein_ctrl.best_idx[5] ),
    .C1(_0771_),
    .B1(_0741_),
    .A1(\levenshtein_ctrl.best_distance[5] ),
    .Y(_0772_),
    .A2(_0740_));
 sg13g2_o21ai_1 _2803_ (.B1(_0747_),
    .Y(_0773_),
    .A1(\arbiter.wbm_dat_i[5] ),
    .A2(net368));
 sg13g2_a21oi_1 _2804_ (.A1(net369),
    .A2(_0772_),
    .Y(_0774_),
    .B1(_0773_));
 sg13g2_a21oi_1 _2805_ (.A1(net506),
    .A2(_0738_),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_nor2_1 _2806_ (.A(net534),
    .B(net339),
    .Y(_0776_));
 sg13g2_a21oi_1 _2807_ (.A1(net338),
    .A2(_0775_),
    .Y(_0245_),
    .B1(_0776_));
 sg13g2_and2_1 _2808_ (.A(\levenshtein_ctrl.best_idx[6] ),
    .B(_0741_),
    .X(_0777_));
 sg13g2_a221oi_1 _2809_ (.B2(\levenshtein_ctrl.best_distance[6] ),
    .C1(_0777_),
    .B1(_0740_),
    .A1(\levenshtein_ctrl.best_idx[14] ),
    .Y(_0778_),
    .A2(_0739_));
 sg13g2_o21ai_1 _2810_ (.B1(_0747_),
    .Y(_0779_),
    .A1(\arbiter.wbm_dat_i[6] ),
    .A2(net368));
 sg13g2_a21oi_1 _2811_ (.A1(net369),
    .A2(_0778_),
    .Y(_0780_),
    .B1(_0779_));
 sg13g2_a21oi_1 _2812_ (.A1(\arbiter.wbs0_dat_i[5] ),
    .A2(_0738_),
    .Y(_0781_),
    .B1(_0780_));
 sg13g2_nor2_1 _2813_ (.A(net485),
    .B(net339),
    .Y(_0782_));
 sg13g2_a21oi_1 _2814_ (.A1(net339),
    .A2(_0781_),
    .Y(_0246_),
    .B1(_0782_));
 sg13g2_and2_1 _2815_ (.A(\levenshtein_ctrl.best_idx[15] ),
    .B(_0739_),
    .X(_0783_));
 sg13g2_a221oi_1 _2816_ (.B2(\levenshtein_ctrl.best_idx[7] ),
    .C1(_0783_),
    .B1(_0741_),
    .A1(\levenshtein_ctrl.best_distance[7] ),
    .Y(_0784_),
    .A2(_0740_));
 sg13g2_o21ai_1 _2817_ (.B1(_0747_),
    .Y(_0785_),
    .A1(\arbiter.wbm_dat_i[7] ),
    .A2(net368));
 sg13g2_a21oi_1 _2818_ (.A1(net368),
    .A2(_0784_),
    .Y(_0786_),
    .B1(_0785_));
 sg13g2_a21oi_1 _2819_ (.A1(net485),
    .A2(_0738_),
    .Y(_0787_),
    .B1(_0786_));
 sg13g2_nor2_1 _2820_ (.A(net531),
    .B(net339),
    .Y(_0788_));
 sg13g2_a21oi_1 _2821_ (.A1(net340),
    .A2(_0787_),
    .Y(_0247_),
    .B1(_0788_));
 sg13g2_nor2_1 _2822_ (.A(net531),
    .B(net671),
    .Y(_0789_));
 sg13g2_nor2_1 _2823_ (.A(net678),
    .B(net339),
    .Y(_0790_));
 sg13g2_a21oi_1 _2824_ (.A1(net339),
    .A2(_0789_),
    .Y(_0248_),
    .B1(_0790_));
 sg13g2_nor2_1 _2825_ (.A(_1100_),
    .B(_1181_),
    .Y(_0791_));
 sg13g2_o21ai_1 _2826_ (.B1(net407),
    .Y(_0792_),
    .A1(_1130_),
    .A2(_0791_));
 sg13g2_nand2b_2 _2827_ (.Y(_0793_),
    .B(_0792_),
    .A_N(net352));
 sg13g2_nand2_2 _2828_ (.Y(_0794_),
    .A(net407),
    .B(_1140_));
 sg13g2_a21oi_1 _2829_ (.A1(_0066_),
    .A2(_1099_),
    .Y(_0795_),
    .B1(net596));
 sg13g2_a21oi_1 _2830_ (.A1(_0794_),
    .A2(net597),
    .Y(_0249_),
    .B1(_0793_));
 sg13g2_nand2_1 _2831_ (.Y(_0796_),
    .A(net558),
    .B(_1129_));
 sg13g2_a21oi_1 _2832_ (.A1(_0794_),
    .A2(_0796_),
    .Y(_0250_),
    .B1(_0793_));
 sg13g2_nand2_1 _2833_ (.Y(_0797_),
    .A(net627),
    .B(_1129_));
 sg13g2_a21oi_1 _2834_ (.A1(_0794_),
    .A2(_0797_),
    .Y(_0251_),
    .B1(_0793_));
 sg13g2_nand2_1 _2835_ (.Y(_0798_),
    .A(net613),
    .B(_1129_));
 sg13g2_a21oi_1 _2836_ (.A1(_0794_),
    .A2(_0798_),
    .Y(_0252_),
    .B1(_0793_));
 sg13g2_nor3_1 _2837_ (.A(net279),
    .B(net352),
    .C(_1131_),
    .Y(_0253_));
 sg13g2_a21oi_1 _2838_ (.A1(net425),
    .A2(\levenshtein_ctrl.dict_address[3] ),
    .Y(_0799_),
    .B1(net391));
 sg13g2_a21oi_1 _2839_ (.A1(_0051_),
    .A2(net391),
    .Y(_0800_),
    .B1(_0799_));
 sg13g2_nand2_1 _2840_ (.Y(_0801_),
    .A(_1145_),
    .B(_0800_));
 sg13g2_o21ai_1 _2841_ (.B1(_0801_),
    .Y(_0802_),
    .A1(_0024_),
    .A2(_1145_));
 sg13g2_a21oi_1 _2842_ (.A1(net402),
    .A2(_0015_),
    .Y(_0803_),
    .B1(_1105_));
 sg13g2_o21ai_1 _2843_ (.B1(_0803_),
    .Y(_0804_),
    .A1(net403),
    .A2(_0802_));
 sg13g2_nor2_1 _2844_ (.A(\levenshtein_ctrl.dict_address[11] ),
    .B(net388),
    .Y(_0805_));
 sg13g2_a21oi_1 _2845_ (.A1(_0044_),
    .A2(net388),
    .Y(_0806_),
    .B1(_0805_));
 sg13g2_a22oi_1 _2846_ (.Y(_0807_),
    .B1(_1172_),
    .B2(_0806_),
    .A2(\arbiter.wbs0_adr_i[13] ),
    .A1(net403));
 sg13g2_nor2_1 _2847_ (.A(net417),
    .B(_0807_),
    .Y(_0808_));
 sg13g2_o21ai_1 _2848_ (.B1(\levenshtein_ctrl.dict_address[7] ),
    .Y(_0809_),
    .A1(net424),
    .A2(net389));
 sg13g2_a21oi_1 _2849_ (.A1(_1145_),
    .A2(_0809_),
    .Y(_0810_),
    .B1(net401));
 sg13g2_a21oi_1 _2850_ (.A1(net403),
    .A2(\arbiter.wbs0_adr_i[9] ),
    .Y(_0811_),
    .B1(_0810_));
 sg13g2_a21oi_1 _2851_ (.A1(net417),
    .A2(_0811_),
    .Y(_0812_),
    .B1(net419));
 sg13g2_nor2_1 _2852_ (.A(_0808_),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_and2_1 _2853_ (.A(_0028_),
    .B(_1146_),
    .X(_0814_));
 sg13g2_nor3_1 _2854_ (.A(\levenshtein_ctrl.state[2] ),
    .B(\levenshtein_ctrl.state[6] ),
    .C(net385),
    .Y(_0815_));
 sg13g2_nor3_1 _2855_ (.A(net401),
    .B(_0814_),
    .C(_0815_),
    .Y(_0816_));
 sg13g2_o21ai_1 _2856_ (.B1(_1096_),
    .Y(_0817_),
    .A1(net399),
    .A2(_0019_));
 sg13g2_o21ai_1 _2857_ (.B1(_1144_),
    .Y(_0818_),
    .A1(_0816_),
    .A2(_0817_));
 sg13g2_a21oi_1 _2858_ (.A1(_0804_),
    .A2(_0813_),
    .Y(_0819_),
    .B1(_0818_));
 sg13g2_nand2_1 _2859_ (.Y(_0820_),
    .A(_0036_),
    .B(net386));
 sg13g2_o21ai_1 _2860_ (.B1(_0820_),
    .Y(_0821_),
    .A1(\levenshtein_ctrl.dict_address[19] ),
    .A2(net386));
 sg13g2_a21oi_1 _2861_ (.A1(_0040_),
    .A2(net387),
    .Y(_0822_),
    .B1(net418));
 sg13g2_o21ai_1 _2862_ (.B1(_0822_),
    .Y(_0823_),
    .A1(\levenshtein_ctrl.dict_address[15] ),
    .A2(net386));
 sg13g2_o21ai_1 _2863_ (.B1(_0823_),
    .Y(_0824_),
    .A1(net398),
    .A2(_0821_));
 sg13g2_mux2_1 _2864_ (.A0(\arbiter.wbs0_adr_i[17] ),
    .A1(\arbiter.wbs0_adr_i[21] ),
    .S(net419),
    .X(_0825_));
 sg13g2_a22oi_1 _2865_ (.Y(_0826_),
    .B1(_0825_),
    .B2(net402),
    .A2(_0824_),
    .A1(_1172_));
 sg13g2_nor2_1 _2866_ (.A(_1142_),
    .B(_0826_),
    .Y(_0827_));
 sg13g2_nor3_1 _2867_ (.A(_0794_),
    .B(_0819_),
    .C(_0827_),
    .Y(_0828_));
 sg13g2_nand2_2 _2868_ (.Y(_0829_),
    .A(net407),
    .B(_1100_));
 sg13g2_nor2_1 _2869_ (.A(net534),
    .B(_1181_),
    .Y(_0830_));
 sg13g2_a21oi_1 _2870_ (.A1(net662),
    .A2(net367),
    .Y(_0831_),
    .B1(_0829_));
 sg13g2_o21ai_1 _2871_ (.B1(_0831_),
    .Y(_0832_),
    .A1(net367),
    .A2(_0830_));
 sg13g2_nand4_1 _2872_ (.B(\spi_ctrl.bit_counter[3] ),
    .C(_0066_),
    .A(net405),
    .Y(_0833_),
    .D(_1121_));
 sg13g2_o21ai_1 _2873_ (.B1(_0794_),
    .Y(_0834_),
    .A1(_0829_),
    .A2(_0833_));
 sg13g2_o21ai_1 _2874_ (.B1(_0832_),
    .Y(_0835_),
    .A1(net732),
    .A2(_0834_));
 sg13g2_nor3_1 _2875_ (.A(net351),
    .B(_0828_),
    .C(_0835_),
    .Y(_0254_));
 sg13g2_a21oi_1 _2876_ (.A1(\levenshtein_ctrl.dict_address[8] ),
    .A2(net392),
    .Y(_0836_),
    .B1(net418));
 sg13g2_o21ai_1 _2877_ (.B1(_0836_),
    .Y(_0837_),
    .A1(_0047_),
    .A2(net392));
 sg13g2_o21ai_1 _2878_ (.B1(net418),
    .Y(_0838_),
    .A1(_0043_),
    .A2(net392));
 sg13g2_a21oi_1 _2879_ (.A1(\levenshtein_ctrl.dict_address[12] ),
    .A2(net392),
    .Y(_0839_),
    .B1(_0838_));
 sg13g2_nor2_1 _2880_ (.A(_1171_),
    .B(_0839_),
    .Y(_0840_));
 sg13g2_a21oi_1 _2881_ (.A1(_0837_),
    .A2(_0840_),
    .Y(_0841_),
    .B1(net401));
 sg13g2_o21ai_1 _2882_ (.B1(net402),
    .Y(_0842_),
    .A1(net419),
    .A2(_0968_));
 sg13g2_a21oi_1 _2883_ (.A1(net419),
    .A2(\arbiter.wbs0_adr_i[14] ),
    .Y(_0843_),
    .B1(_0842_));
 sg13g2_o21ai_1 _2884_ (.B1(_1121_),
    .Y(_0844_),
    .A1(_0841_),
    .A2(_0843_));
 sg13g2_a21oi_1 _2885_ (.A1(net424),
    .A2(\levenshtein_ctrl.dict_address[4] ),
    .Y(_0845_),
    .B1(net390));
 sg13g2_a21oi_1 _2886_ (.A1(_0050_),
    .A2(net390),
    .Y(_0846_),
    .B1(_0845_));
 sg13g2_nand2_1 _2887_ (.Y(_0847_),
    .A(_1145_),
    .B(_0846_));
 sg13g2_o21ai_1 _2888_ (.B1(_0847_),
    .Y(_0848_),
    .A1(_0023_),
    .A2(_1145_));
 sg13g2_o21ai_1 _2889_ (.B1(_1104_),
    .Y(_0849_),
    .A1(net400),
    .A2(_0014_));
 sg13g2_a21o_1 _2890_ (.A2(_0848_),
    .A1(net399),
    .B1(_0849_),
    .X(_0850_));
 sg13g2_a21oi_1 _2891_ (.A1(net425),
    .A2(\levenshtein_ctrl.dict_address[0] ),
    .Y(_0851_),
    .B1(net390));
 sg13g2_a21oi_1 _2892_ (.A1(_0054_),
    .A2(net391),
    .Y(_0852_),
    .B1(_0851_));
 sg13g2_a21oi_1 _2893_ (.A1(_0027_),
    .A2(net385),
    .Y(_0853_),
    .B1(net401));
 sg13g2_o21ai_1 _2894_ (.B1(_0853_),
    .Y(_0854_),
    .A1(net385),
    .A2(_0852_));
 sg13g2_a21oi_1 _2895_ (.A1(net404),
    .A2(_0967_),
    .Y(_0855_),
    .B1(_1097_));
 sg13g2_nand2_1 _2896_ (.Y(_0856_),
    .A(_0854_),
    .B(_0855_));
 sg13g2_nand4_1 _2897_ (.B(_0844_),
    .C(_0850_),
    .A(_1144_),
    .Y(_0857_),
    .D(_0856_));
 sg13g2_nand2_1 _2898_ (.Y(_0858_),
    .A(_0035_),
    .B(net386));
 sg13g2_o21ai_1 _2899_ (.B1(_0858_),
    .Y(_0859_),
    .A1(\levenshtein_ctrl.dict_address[20] ),
    .A2(net386));
 sg13g2_a21oi_1 _2900_ (.A1(_0039_),
    .A2(net386),
    .Y(_0860_),
    .B1(net418));
 sg13g2_o21ai_1 _2901_ (.B1(_0860_),
    .Y(_0861_),
    .A1(\levenshtein_ctrl.dict_address[16] ),
    .A2(net386));
 sg13g2_o21ai_1 _2902_ (.B1(_0861_),
    .Y(_0862_),
    .A1(net398),
    .A2(_0859_));
 sg13g2_mux2_1 _2903_ (.A0(\arbiter.wbs0_adr_i[18] ),
    .A1(\arbiter.wbs0_adr_i[22] ),
    .S(net419),
    .X(_0863_));
 sg13g2_a22oi_1 _2904_ (.Y(_0864_),
    .B1(_0863_),
    .B2(net402),
    .A2(_0862_),
    .A1(_1172_));
 sg13g2_o21ai_1 _2905_ (.B1(_0857_),
    .Y(_0865_),
    .A1(_1142_),
    .A2(_0864_));
 sg13g2_nor2_1 _2906_ (.A(_0794_),
    .B(_0865_),
    .Y(_0866_));
 sg13g2_nor2_1 _2907_ (.A(net485),
    .B(_1181_),
    .Y(_0867_));
 sg13g2_a21oi_1 _2908_ (.A1(net628),
    .A2(net367),
    .Y(_0868_),
    .B1(_0829_));
 sg13g2_o21ai_1 _2909_ (.B1(_0868_),
    .Y(_0869_),
    .A1(net367),
    .A2(_0867_));
 sg13g2_o21ai_1 _2910_ (.B1(_0869_),
    .Y(_0870_),
    .A1(net731),
    .A2(_0834_));
 sg13g2_nor3_1 _2911_ (.A(net351),
    .B(_0866_),
    .C(_0870_),
    .Y(_0255_));
 sg13g2_a21oi_1 _2912_ (.A1(\levenshtein_ctrl.dict_address[9] ),
    .A2(net392),
    .Y(_0871_),
    .B1(net418));
 sg13g2_o21ai_1 _2913_ (.B1(_0871_),
    .Y(_0872_),
    .A1(_0046_),
    .A2(net392));
 sg13g2_o21ai_1 _2914_ (.B1(net418),
    .Y(_0873_),
    .A1(_0042_),
    .A2(net392));
 sg13g2_a21oi_1 _2915_ (.A1(\levenshtein_ctrl.dict_address[13] ),
    .A2(net392),
    .Y(_0874_),
    .B1(_0873_));
 sg13g2_nor2_1 _2916_ (.A(_1171_),
    .B(_0874_),
    .Y(_0875_));
 sg13g2_a21oi_1 _2917_ (.A1(_0872_),
    .A2(_0875_),
    .Y(_0876_),
    .B1(net401));
 sg13g2_o21ai_1 _2918_ (.B1(net402),
    .Y(_0877_),
    .A1(net419),
    .A2(_0969_));
 sg13g2_a21oi_1 _2919_ (.A1(net419),
    .A2(\arbiter.wbs0_adr_i[15] ),
    .Y(_0878_),
    .B1(_0877_));
 sg13g2_o21ai_1 _2920_ (.B1(_1121_),
    .Y(_0879_),
    .A1(_0876_),
    .A2(_0878_));
 sg13g2_a21oi_1 _2921_ (.A1(net424),
    .A2(\levenshtein_ctrl.dict_address[5] ),
    .Y(_0880_),
    .B1(net390));
 sg13g2_a21oi_1 _2922_ (.A1(_0049_),
    .A2(net390),
    .Y(_0881_),
    .B1(_0880_));
 sg13g2_a21oi_1 _2923_ (.A1(_0022_),
    .A2(net385),
    .Y(_0882_),
    .B1(net401));
 sg13g2_o21ai_1 _2924_ (.B1(_0882_),
    .Y(_0883_),
    .A1(net385),
    .A2(_0881_));
 sg13g2_o21ai_1 _2925_ (.B1(_1104_),
    .Y(_0884_),
    .A1(net400),
    .A2(_0013_));
 sg13g2_nand2b_1 _2926_ (.Y(_0885_),
    .B(_0883_),
    .A_N(_0884_));
 sg13g2_a21oi_1 _2927_ (.A1(net424),
    .A2(\levenshtein_ctrl.dict_address[1] ),
    .Y(_0886_),
    .B1(net390));
 sg13g2_a21oi_1 _2928_ (.A1(_0053_),
    .A2(net391),
    .Y(_0887_),
    .B1(_0886_));
 sg13g2_a21oi_1 _2929_ (.A1(_0026_),
    .A2(net385),
    .Y(_0888_),
    .B1(net401));
 sg13g2_o21ai_1 _2930_ (.B1(_0888_),
    .Y(_0889_),
    .A1(net385),
    .A2(_0887_));
 sg13g2_o21ai_1 _2931_ (.B1(_1096_),
    .Y(_0890_),
    .A1(net399),
    .A2(_0017_));
 sg13g2_nand2b_1 _2932_ (.Y(_0891_),
    .B(_0889_),
    .A_N(_0890_));
 sg13g2_nand4_1 _2933_ (.B(_0879_),
    .C(_0885_),
    .A(_1144_),
    .Y(_0892_),
    .D(_0891_));
 sg13g2_nand2_1 _2934_ (.Y(_0893_),
    .A(\levenshtein_ctrl.dict_address[17] ),
    .B(_1110_));
 sg13g2_o21ai_1 _2935_ (.B1(_0893_),
    .Y(_0894_),
    .A1(_0038_),
    .A2(_1110_));
 sg13g2_a22oi_1 _2936_ (.Y(_0895_),
    .B1(_1172_),
    .B2(_0894_),
    .A2(\arbiter.wbs0_adr_i[19] ),
    .A1(net402));
 sg13g2_nand2b_1 _2937_ (.Y(_0896_),
    .B(_1098_),
    .A_N(_0895_));
 sg13g2_nand3_1 _2938_ (.B(_0892_),
    .C(_0896_),
    .A(_1140_),
    .Y(_0897_));
 sg13g2_nor2_1 _2939_ (.A(net531),
    .B(_1181_),
    .Y(_0898_));
 sg13g2_nor2_1 _2940_ (.A(_1182_),
    .B(_0898_),
    .Y(_0899_));
 sg13g2_nand2_1 _2941_ (.Y(_0900_),
    .A(net650),
    .B(net367));
 sg13g2_nand2_1 _2942_ (.Y(_0901_),
    .A(_1100_),
    .B(_0900_));
 sg13g2_o21ai_1 _2943_ (.B1(_0897_),
    .Y(_0902_),
    .A1(_0899_),
    .A2(_0901_));
 sg13g2_a21o_1 _2944_ (.A2(_0900_),
    .A1(_1181_),
    .B1(_0829_),
    .X(_0903_));
 sg13g2_a21oi_1 _2945_ (.A1(net408),
    .A2(_1140_),
    .Y(_0904_),
    .B1(net722));
 sg13g2_a221oi_1 _2946_ (.B2(_0904_),
    .C1(net351),
    .B1(_0903_),
    .A1(net407),
    .Y(_0256_),
    .A2(_0902_));
 sg13g2_mux2_1 _2947_ (.A0(_0931_),
    .A1(_0932_),
    .S(\spi_ctrl.ss_n ),
    .X(_0905_));
 sg13g2_nor2_1 _2948_ (.A(net351),
    .B(net607),
    .Y(_0257_));
 sg13g2_or2_1 _2949_ (.X(_0906_),
    .B(net351),
    .A(_0932_));
 sg13g2_mux2_1 _2950_ (.A0(net4),
    .A1(\arbiter.wbm_dat_i[0] ),
    .S(_0906_),
    .X(_0258_));
 sg13g2_mux2_1 _2951_ (.A0(net5),
    .A1(net756),
    .S(_0906_),
    .X(_0259_));
 sg13g2_mux2_1 _2952_ (.A0(net6),
    .A1(\arbiter.wbm_dat_i[2] ),
    .S(net337),
    .X(_0260_));
 sg13g2_nor2_1 _2953_ (.A(net7),
    .B(net337),
    .Y(_0907_));
 sg13g2_a21oi_1 _2954_ (.A1(_0963_),
    .A2(net337),
    .Y(_0261_),
    .B1(_0907_));
 sg13g2_mux2_1 _2955_ (.A0(\arbiter.wbm_dat_i[0] ),
    .A1(\arbiter.wbm_dat_i[4] ),
    .S(net337),
    .X(_0262_));
 sg13g2_mux2_1 _2956_ (.A0(\arbiter.wbm_dat_i[1] ),
    .A1(net754),
    .S(net337),
    .X(_0263_));
 sg13g2_mux2_1 _2957_ (.A0(\arbiter.wbm_dat_i[2] ),
    .A1(\arbiter.wbm_dat_i[6] ),
    .S(net337),
    .X(_0264_));
 sg13g2_nand2_1 _2958_ (.Y(_0908_),
    .A(net693),
    .B(net337));
 sg13g2_o21ai_1 _2959_ (.B1(_0908_),
    .Y(_0265_),
    .A1(_0963_),
    .A2(net337));
 sg13g2_nor3_1 _2960_ (.A(net660),
    .B(net393),
    .C(_1058_),
    .Y(_0909_));
 sg13g2_nor2_1 _2961_ (.A(net721),
    .B(net376),
    .Y(_0910_));
 sg13g2_a21oi_1 _2962_ (.A1(_0936_),
    .A2(net376),
    .Y(_0266_),
    .B1(_0910_));
 sg13g2_mux2_1 _2963_ (.A0(net588),
    .A1(\arbiter.wbs0_adr_i[1] ),
    .S(net376),
    .X(_0267_));
 sg13g2_mux2_1 _2964_ (.A0(net652),
    .A1(net588),
    .S(net376),
    .X(_0268_));
 sg13g2_mux2_1 _2965_ (.A0(net598),
    .A1(\arbiter.wbs0_adr_i[3] ),
    .S(net375),
    .X(_0269_));
 sg13g2_mux2_1 _2966_ (.A0(net561),
    .A1(\arbiter.wbs0_adr_i[4] ),
    .S(net375),
    .X(_0270_));
 sg13g2_mux2_1 _2967_ (.A0(net504),
    .A1(\arbiter.wbs0_adr_i[5] ),
    .S(net374),
    .X(_0271_));
 sg13g2_mux2_1 _2968_ (.A0(net524),
    .A1(net504),
    .S(net372),
    .X(_0272_));
 sg13g2_mux2_1 _2969_ (.A0(net567),
    .A1(net524),
    .S(net374),
    .X(_0273_));
 sg13g2_mux2_1 _2970_ (.A0(net636),
    .A1(net567),
    .S(net374),
    .X(_0274_));
 sg13g2_nand2_1 _2971_ (.Y(_0911_),
    .A(net636),
    .B(net372));
 sg13g2_o21ai_1 _2972_ (.B1(_0911_),
    .Y(_0275_),
    .A1(_0968_),
    .A2(net373));
 sg13g2_nor2_1 _2973_ (.A(net502),
    .B(net372),
    .Y(_0912_));
 sg13g2_a21oi_1 _2974_ (.A1(_0968_),
    .A2(net373),
    .Y(_0276_),
    .B1(_0912_));
 sg13g2_nor2_1 _2975_ (.A(net655),
    .B(net375),
    .Y(_0913_));
 sg13g2_a21oi_1 _2976_ (.A1(_0969_),
    .A2(net375),
    .Y(_0277_),
    .B1(_0913_));
 sg13g2_mux2_1 _2977_ (.A0(net659),
    .A1(net655),
    .S(net375),
    .X(_0278_));
 sg13g2_mux2_1 _2978_ (.A0(net639),
    .A1(\arbiter.wbs0_adr_i[13] ),
    .S(net375),
    .X(_0279_));
 sg13g2_mux2_1 _2979_ (.A0(net632),
    .A1(\arbiter.wbs0_adr_i[14] ),
    .S(net375),
    .X(_0280_));
 sg13g2_mux2_1 _2980_ (.A0(net604),
    .A1(\arbiter.wbs0_adr_i[15] ),
    .S(net372),
    .X(_0281_));
 sg13g2_mux2_1 _2981_ (.A0(net602),
    .A1(\arbiter.wbs0_adr_i[16] ),
    .S(net372),
    .X(_0282_));
 sg13g2_mux2_1 _2982_ (.A0(net626),
    .A1(net602),
    .S(net372),
    .X(_0283_));
 sg13g2_mux2_1 _2983_ (.A0(net677),
    .A1(net626),
    .S(net372),
    .X(_0284_));
 sg13g2_mux2_1 _2984_ (.A0(net697),
    .A1(net677),
    .S(net373),
    .X(_0285_));
 sg13g2_mux2_1 _2985_ (.A0(net681),
    .A1(\arbiter.wbs0_adr_i[20] ),
    .S(net373),
    .X(_0286_));
 sg13g2_mux2_1 _2986_ (.A0(net610),
    .A1(net681),
    .S(net372),
    .X(_0287_));
 sg13g2_nand2_1 _2987_ (.Y(_0914_),
    .A(net610),
    .B(net376));
 sg13g2_o21ai_1 _2988_ (.B1(net611),
    .Y(_0288_),
    .A1(_0937_),
    .A2(net376));
 sg13g2_a21oi_1 _2989_ (.A1(net407),
    .A2(_1104_),
    .Y(_0915_),
    .B1(net405));
 sg13g2_nor2_1 _2990_ (.A(_1108_),
    .B(_0915_),
    .Y(_0916_));
 sg13g2_and2_1 _2991_ (.A(_1125_),
    .B(_0916_),
    .X(_0289_));
 sg13g2_xnor2_1 _2992_ (.Y(_0917_),
    .A(_0964_),
    .B(_1127_));
 sg13g2_nor2_1 _2993_ (.A(_0932_),
    .B(_0917_),
    .Y(_0918_));
 sg13g2_a221oi_1 _2994_ (.B2(_0918_),
    .C1(_1108_),
    .B1(_1118_),
    .A1(_0930_),
    .Y(_0290_),
    .A2(_0932_));
 sg13g2_a21o_1 _2995_ (.A2(_1201_),
    .A1(_1092_),
    .B1(_1094_),
    .X(_0291_));
 sg13g2_nor2_1 _2996_ (.A(\arbiter.wbs0_dat_i[0] ),
    .B(net339),
    .Y(_0919_));
 sg13g2_nor2b_1 _2997_ (.A(_0055_),
    .B_N(_1212_),
    .Y(_0920_));
 sg13g2_a22oi_1 _2998_ (.Y(_0921_),
    .B1(_0741_),
    .B2(\levenshtein_ctrl.best_idx[0] ),
    .A2(_0739_),
    .A1(\levenshtein_ctrl.best_idx[8] ));
 sg13g2_o21ai_1 _2999_ (.B1(_0921_),
    .Y(_0922_),
    .A1(_0056_),
    .A2(_1003_));
 sg13g2_a22oi_1 _3000_ (.Y(_0923_),
    .B1(_0740_),
    .B2(\levenshtein_ctrl.best_distance[0] ),
    .A2(_1203_),
    .A1(\levenshtein_ctrl.sram_config[0] ));
 sg13g2_inv_1 _3001_ (.Y(_0924_),
    .A(_0923_));
 sg13g2_nor4_2 _3002_ (.A(_0743_),
    .B(_0920_),
    .C(_0922_),
    .Y(_0925_),
    .D(_0924_));
 sg13g2_o21ai_1 _3003_ (.B1(_0747_),
    .Y(_0926_),
    .A1(\arbiter.wbm_dat_i[0] ),
    .A2(net369));
 sg13g2_a21oi_1 _3004_ (.A1(net368),
    .A2(_0925_),
    .Y(_0927_),
    .B1(_0926_));
 sg13g2_a21oi_1 _3005_ (.A1(\spi.state[0] ),
    .A2(net664),
    .Y(_0928_),
    .B1(_0927_));
 sg13g2_a21oi_1 _3006_ (.A1(net339),
    .A2(net665),
    .Y(_0292_),
    .B1(_0919_));
 sg13g2_dfrbp_1 _3007_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net17),
    .D(net712),
    .Q_N(_1492_),
    .Q(\levenshtein_ctrl.state[0] ));
 sg13g2_dfrbp_1 _3008_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net18),
    .D(net690),
    .Q_N(_1493_),
    .Q(\levenshtein_ctrl.state[1] ));
 sg13g2_dfrbp_1 _3009_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net19),
    .D(_0002_),
    .Q_N(_1494_),
    .Q(\levenshtein_ctrl.state[2] ));
 sg13g2_dfrbp_1 _3010_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net20),
    .D(net572),
    .Q_N(_0062_),
    .Q(\levenshtein_ctrl.state[3] ));
 sg13g2_dfrbp_1 _3011_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net21),
    .D(_0004_),
    .Q_N(_1495_),
    .Q(\levenshtein_ctrl.state[4] ));
 sg13g2_dfrbp_1 _3012_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net22),
    .D(_0005_),
    .Q_N(_0063_),
    .Q(\levenshtein_ctrl.state[5] ));
 sg13g2_dfrbp_1 _3013_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net28),
    .D(_0006_),
    .Q_N(_0064_),
    .Q(\levenshtein_ctrl.state[6] ));
 sg13g2_dfrbp_1 _3014_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net16),
    .D(_0007_),
    .Q_N(_0061_),
    .Q(\levenshtein_ctrl.state[7] ));
 sg13g2_dfrbp_1 _3015_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net222),
    .D(net294),
    .Q_N(_0060_),
    .Q(\spi.counter[0] ));
 sg13g2_dfrbp_1 _3016_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net220),
    .D(net301),
    .Q_N(_1491_),
    .Q(\spi.counter[1] ));
 sg13g2_dfrbp_1 _3017_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net218),
    .D(net319),
    .Q_N(_1490_),
    .Q(\spi.counter[2] ));
 sg13g2_dfrbp_1 _3018_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net216),
    .D(_0071_),
    .Q_N(_1489_),
    .Q(\spi.counter[3] ));
 sg13g2_dfrbp_1 _3019_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net32),
    .D(_0072_),
    .Q_N(_1496_),
    .Q(\spi.counter[4] ));
 sg13g2_dfrbp_1 _3020_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net214),
    .D(net264),
    .Q_N(_1488_),
    .Q(\spi.last_sck ));
 sg13g2_dfrbp_1 _3021_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net212),
    .D(_0073_),
    .Q_N(_0059_),
    .Q(\levenshtein_ctrl.symbol_idx[0] ));
 sg13g2_dfrbp_1 _3022_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net211),
    .D(net618),
    .Q_N(_1487_),
    .Q(\levenshtein_ctrl.symbol_idx[1] ));
 sg13g2_dfrbp_1 _3023_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net33),
    .D(net289),
    .Q_N(_1497_),
    .Q(\spi.miso ));
 sg13g2_dfrbp_1 _3024_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net34),
    .D(net1),
    .Q_N(_1498_),
    .Q(\spi.ss_n_sync[0] ));
 sg13g2_dfrbp_1 _3025_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net35),
    .D(net263),
    .Q_N(_1499_),
    .Q(\spi.ss_n ));
 sg13g2_dfrbp_1 _3026_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net37),
    .D(net3),
    .Q_N(_1500_),
    .Q(\spi.mosi_sync[0] ));
 sg13g2_dfrbp_1 _3027_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net210),
    .D(net262),
    .Q_N(_1486_),
    .Q(\spi.mosi ));
 sg13g2_dfrbp_1 _3028_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net38),
    .D(net642),
    .Q_N(_0065_),
    .Q(\intercon.wbs_cyc_i ));
 sg13g2_dfrbp_1 _3029_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net253),
    .D(net2),
    .Q_N(_1501_),
    .Q(\spi.sck_sync[0] ));
 sg13g2_dfrbp_1 _3030_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net208),
    .D(net261),
    .Q_N(_1485_),
    .Q(\spi.sck ));
 sg13g2_dfrbp_1 _3031_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net206),
    .D(_0077_),
    .Q_N(_0058_),
    .Q(\spi_ctrl.bit_counter[0] ));
 sg13g2_dfrbp_1 _3032_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net204),
    .D(_0078_),
    .Q_N(_1484_),
    .Q(\spi_ctrl.bit_counter[1] ));
 sg13g2_dfrbp_1 _3033_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net202),
    .D(_0079_),
    .Q_N(_1483_),
    .Q(\spi_ctrl.bit_counter[3] ));
 sg13g2_dfrbp_1 _3034_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net200),
    .D(_0080_),
    .Q_N(_1482_),
    .Q(\spi_ctrl.ss_n ));
 sg13g2_dfrbp_1 _3035_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net199),
    .D(_0081_),
    .Q_N(_1481_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _3036_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net198),
    .D(net720),
    .Q_N(_1480_),
    .Q(\arbiter.cyc ));
 sg13g2_dfrbp_1 _3037_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net197),
    .D(net687),
    .Q_N(_1479_),
    .Q(\levenshtein_ctrl.sram_config[0] ));
 sg13g2_dfrbp_1 _3038_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net196),
    .D(net620),
    .Q_N(_1478_),
    .Q(\levenshtein_ctrl.sram_config[1] ));
 sg13g2_dfrbp_1 _3039_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net195),
    .D(net696),
    .Q_N(_0057_),
    .Q(\arbiter.wbs1_cyc_i ));
 sg13g2_dfrbp_1 _3040_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net193),
    .D(_0086_),
    .Q_N(_1477_),
    .Q(ctrl_slave_ack));
 sg13g2_dfrbp_1 _3041_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net192),
    .D(_0087_),
    .Q_N(_0056_),
    .Q(\levenshtein_ctrl.enabled ));
 sg13g2_dfrbp_1 _3042_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net191),
    .D(net726),
    .Q_N(_0055_),
    .Q(\levenshtein_ctrl.word_length_reg[0] ));
 sg13g2_dfrbp_1 _3043_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net190),
    .D(_0089_),
    .Q_N(_1476_),
    .Q(\levenshtein_ctrl.word_length_reg[1] ));
 sg13g2_dfrbp_1 _3044_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net189),
    .D(_0090_),
    .Q_N(_1475_),
    .Q(\levenshtein_ctrl.word_length_reg[2] ));
 sg13g2_dfrbp_1 _3045_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net188),
    .D(net651),
    .Q_N(_1474_),
    .Q(\levenshtein_ctrl.word_length_reg[3] ));
 sg13g2_dfrbp_1 _3046_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net187),
    .D(_0092_),
    .Q_N(_0054_),
    .Q(\levenshtein_ctrl.dict_address[0] ));
 sg13g2_dfrbp_1 _3047_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net186),
    .D(net514),
    .Q_N(_0053_),
    .Q(\levenshtein_ctrl.dict_address[1] ));
 sg13g2_dfrbp_1 _3048_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net185),
    .D(net528),
    .Q_N(_0052_),
    .Q(\levenshtein_ctrl.dict_address[2] ));
 sg13g2_dfrbp_1 _3049_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net184),
    .D(net457),
    .Q_N(_0051_),
    .Q(\levenshtein_ctrl.dict_address[3] ));
 sg13g2_dfrbp_1 _3050_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net183),
    .D(net511),
    .Q_N(_0050_),
    .Q(\levenshtein_ctrl.dict_address[4] ));
 sg13g2_dfrbp_1 _3051_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net182),
    .D(net501),
    .Q_N(_0049_),
    .Q(\levenshtein_ctrl.dict_address[5] ));
 sg13g2_dfrbp_1 _3052_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net181),
    .D(net584),
    .Q_N(_0048_),
    .Q(\levenshtein_ctrl.dict_address[6] ));
 sg13g2_dfrbp_1 _3053_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net180),
    .D(net623),
    .Q_N(_1473_),
    .Q(\levenshtein_ctrl.dict_address[7] ));
 sg13g2_dfrbp_1 _3054_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net179),
    .D(net467),
    .Q_N(_0047_),
    .Q(\levenshtein_ctrl.dict_address[8] ));
 sg13g2_dfrbp_1 _3055_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net178),
    .D(net497),
    .Q_N(_0046_),
    .Q(\levenshtein_ctrl.dict_address[9] ));
 sg13g2_dfrbp_1 _3056_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net177),
    .D(net625),
    .Q_N(_0045_),
    .Q(\levenshtein_ctrl.dict_address[10] ));
 sg13g2_dfrbp_1 _3057_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net176),
    .D(net463),
    .Q_N(_0044_),
    .Q(\levenshtein_ctrl.dict_address[11] ));
 sg13g2_dfrbp_1 _3058_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net175),
    .D(net657),
    .Q_N(_0043_),
    .Q(\levenshtein_ctrl.dict_address[12] ));
 sg13g2_dfrbp_1 _3059_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net174),
    .D(net545),
    .Q_N(_0042_),
    .Q(\levenshtein_ctrl.dict_address[13] ));
 sg13g2_dfrbp_1 _3060_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net173),
    .D(net609),
    .Q_N(_0041_),
    .Q(\levenshtein_ctrl.dict_address[14] ));
 sg13g2_dfrbp_1 _3061_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net172),
    .D(net449),
    .Q_N(_0040_),
    .Q(\levenshtein_ctrl.dict_address[15] ));
 sg13g2_dfrbp_1 _3062_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net171),
    .D(net594),
    .Q_N(_0039_),
    .Q(\levenshtein_ctrl.dict_address[16] ));
 sg13g2_dfrbp_1 _3063_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net170),
    .D(net537),
    .Q_N(_0038_),
    .Q(\levenshtein_ctrl.dict_address[17] ));
 sg13g2_dfrbp_1 _3064_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net169),
    .D(net564),
    .Q_N(_0037_),
    .Q(\levenshtein_ctrl.dict_address[18] ));
 sg13g2_dfrbp_1 _3065_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net168),
    .D(net548),
    .Q_N(_0036_),
    .Q(\levenshtein_ctrl.dict_address[19] ));
 sg13g2_dfrbp_1 _3066_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net167),
    .D(net554),
    .Q_N(_0035_),
    .Q(\levenshtein_ctrl.dict_address[20] ));
 sg13g2_dfrbp_1 _3067_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net166),
    .D(_0113_),
    .Q_N(_1472_),
    .Q(\levenshtein_ctrl.pm[0] ));
 sg13g2_dfrbp_1 _3068_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net165),
    .D(_0114_),
    .Q_N(_1471_),
    .Q(\levenshtein_ctrl.pm[1] ));
 sg13g2_dfrbp_1 _3069_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net164),
    .D(_0115_),
    .Q_N(_1470_),
    .Q(\levenshtein_ctrl.pm[2] ));
 sg13g2_dfrbp_1 _3070_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net163),
    .D(net509),
    .Q_N(_1469_),
    .Q(\levenshtein_ctrl.pm[3] ));
 sg13g2_dfrbp_1 _3071_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net162),
    .D(_0117_),
    .Q_N(_1468_),
    .Q(\levenshtein_ctrl.pm[4] ));
 sg13g2_dfrbp_1 _3072_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net161),
    .D(net616),
    .Q_N(_1467_),
    .Q(\levenshtein_ctrl.pm[5] ));
 sg13g2_dfrbp_1 _3073_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net160),
    .D(_0119_),
    .Q_N(_1466_),
    .Q(\levenshtein_ctrl.pm[6] ));
 sg13g2_dfrbp_1 _3074_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net159),
    .D(_0120_),
    .Q_N(_1465_),
    .Q(\levenshtein_ctrl.pm[7] ));
 sg13g2_dfrbp_1 _3075_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net158),
    .D(net469),
    .Q_N(_0034_),
    .Q(\levenshtein_ctrl.vp[0] ));
 sg13g2_dfrbp_1 _3076_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net157),
    .D(_0122_),
    .Q_N(_1464_),
    .Q(\levenshtein_ctrl.vp[1] ));
 sg13g2_dfrbp_1 _3077_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net156),
    .D(_0123_),
    .Q_N(_1463_),
    .Q(\levenshtein_ctrl.vp[2] ));
 sg13g2_dfrbp_1 _3078_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net155),
    .D(_0124_),
    .Q_N(_1462_),
    .Q(\levenshtein_ctrl.vp[3] ));
 sg13g2_dfrbp_1 _3079_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net154),
    .D(net751),
    .Q_N(_1461_),
    .Q(\levenshtein_ctrl.vp[4] ));
 sg13g2_dfrbp_1 _3080_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net153),
    .D(_0126_),
    .Q_N(_1460_),
    .Q(\levenshtein_ctrl.vp[5] ));
 sg13g2_dfrbp_1 _3081_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net152),
    .D(_0127_),
    .Q_N(_1459_),
    .Q(\levenshtein_ctrl.vp[6] ));
 sg13g2_dfrbp_1 _3082_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net151),
    .D(_0128_),
    .Q_N(_1458_),
    .Q(\levenshtein_ctrl.vp[7] ));
 sg13g2_dfrbp_1 _3083_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net150),
    .D(net740),
    .Q_N(_1457_),
    .Q(\levenshtein_ctrl.vp[8] ));
 sg13g2_dfrbp_1 _3084_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net149),
    .D(_0130_),
    .Q_N(_1456_),
    .Q(\levenshtein_ctrl.vp[9] ));
 sg13g2_dfrbp_1 _3085_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net148),
    .D(net724),
    .Q_N(_1455_),
    .Q(\levenshtein_ctrl.vp[10] ));
 sg13g2_dfrbp_1 _3086_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net147),
    .D(net738),
    .Q_N(_1454_),
    .Q(\levenshtein_ctrl.vp[11] ));
 sg13g2_dfrbp_1 _3087_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net146),
    .D(_0133_),
    .Q_N(_1453_),
    .Q(\levenshtein_ctrl.vp[12] ));
 sg13g2_dfrbp_1 _3088_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net145),
    .D(net744),
    .Q_N(_1452_),
    .Q(\levenshtein_ctrl.vp[13] ));
 sg13g2_dfrbp_1 _3089_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net144),
    .D(_0135_),
    .Q_N(_1451_),
    .Q(\levenshtein_ctrl.vp[14] ));
 sg13g2_dfrbp_1 _3090_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net143),
    .D(_0136_),
    .Q_N(_0033_),
    .Q(\levenshtein_ctrl.vp[15] ));
 sg13g2_dfrbp_1 _3091_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net142),
    .D(_0137_),
    .Q_N(_0032_),
    .Q(\levenshtein_ctrl.vn[0] ));
 sg13g2_dfrbp_1 _3092_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net141),
    .D(net284),
    .Q_N(_1450_),
    .Q(\levenshtein_ctrl.vn[1] ));
 sg13g2_dfrbp_1 _3093_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net140),
    .D(net442),
    .Q_N(_1449_),
    .Q(\levenshtein_ctrl.vn[2] ));
 sg13g2_dfrbp_1 _3094_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net139),
    .D(_0140_),
    .Q_N(_1448_),
    .Q(\levenshtein_ctrl.vn[3] ));
 sg13g2_dfrbp_1 _3095_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net138),
    .D(_0141_),
    .Q_N(_1447_),
    .Q(\levenshtein_ctrl.vn[4] ));
 sg13g2_dfrbp_1 _3096_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net137),
    .D(net309),
    .Q_N(_1446_),
    .Q(\levenshtein_ctrl.vn[5] ));
 sg13g2_dfrbp_1 _3097_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net136),
    .D(_0143_),
    .Q_N(_1445_),
    .Q(\levenshtein_ctrl.vn[6] ));
 sg13g2_dfrbp_1 _3098_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net135),
    .D(_0144_),
    .Q_N(_1444_),
    .Q(\levenshtein_ctrl.vn[7] ));
 sg13g2_dfrbp_1 _3099_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net134),
    .D(net482),
    .Q_N(_1443_),
    .Q(\levenshtein_ctrl.vn[8] ));
 sg13g2_dfrbp_1 _3100_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net133),
    .D(_0146_),
    .Q_N(_1442_),
    .Q(\levenshtein_ctrl.vn[9] ));
 sg13g2_dfrbp_1 _3101_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net132),
    .D(net566),
    .Q_N(_1441_),
    .Q(\levenshtein_ctrl.vn[10] ));
 sg13g2_dfrbp_1 _3102_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net131),
    .D(_0148_),
    .Q_N(_1440_),
    .Q(\levenshtein_ctrl.vn[11] ));
 sg13g2_dfrbp_1 _3103_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net130),
    .D(net325),
    .Q_N(_1439_),
    .Q(\levenshtein_ctrl.vn[12] ));
 sg13g2_dfrbp_1 _3104_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net129),
    .D(_0150_),
    .Q_N(_1438_),
    .Q(\levenshtein_ctrl.vn[13] ));
 sg13g2_dfrbp_1 _3105_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net128),
    .D(_0151_),
    .Q_N(_1437_),
    .Q(\levenshtein_ctrl.vn[14] ));
 sg13g2_dfrbp_1 _3106_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net127),
    .D(net286),
    .Q_N(_0031_),
    .Q(\levenshtein_ctrl.vn[15] ));
 sg13g2_dfrbp_1 _3107_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net126),
    .D(net268),
    .Q_N(_0030_),
    .Q(\levenshtein_ctrl.d[0] ));
 sg13g2_dfrbp_1 _3108_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net125),
    .D(_0154_),
    .Q_N(_1436_),
    .Q(\levenshtein_ctrl.d[1] ));
 sg13g2_dfrbp_1 _3109_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net124),
    .D(_0155_),
    .Q_N(_1435_),
    .Q(\levenshtein_ctrl.d[2] ));
 sg13g2_dfrbp_1 _3110_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net123),
    .D(_0156_),
    .Q_N(_1434_),
    .Q(\levenshtein_ctrl.d[3] ));
 sg13g2_dfrbp_1 _3111_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net122),
    .D(_0157_),
    .Q_N(_1433_),
    .Q(\levenshtein_ctrl.d[4] ));
 sg13g2_dfrbp_1 _3112_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net121),
    .D(_0158_),
    .Q_N(_1432_),
    .Q(\levenshtein_ctrl.d[5] ));
 sg13g2_dfrbp_1 _3113_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net120),
    .D(net648),
    .Q_N(_1431_),
    .Q(\levenshtein_ctrl.d[6] ));
 sg13g2_dfrbp_1 _3114_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net119),
    .D(net577),
    .Q_N(_1430_),
    .Q(\levenshtein_ctrl.d[7] ));
 sg13g2_dfrbp_1 _3115_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net118),
    .D(net266),
    .Q_N(_0029_),
    .Q(\levenshtein_ctrl.idx[0] ));
 sg13g2_dfrbp_1 _3116_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net117),
    .D(net592),
    .Q_N(_1429_),
    .Q(\levenshtein_ctrl.idx[1] ));
 sg13g2_dfrbp_1 _3117_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net116),
    .D(net494),
    .Q_N(_1428_),
    .Q(\levenshtein_ctrl.idx[2] ));
 sg13g2_dfrbp_1 _3118_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net115),
    .D(_0164_),
    .Q_N(_1427_),
    .Q(\levenshtein_ctrl.idx[3] ));
 sg13g2_dfrbp_1 _3119_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net114),
    .D(net521),
    .Q_N(_1426_),
    .Q(\levenshtein_ctrl.idx[4] ));
 sg13g2_dfrbp_1 _3120_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net113),
    .D(_0166_),
    .Q_N(_1425_),
    .Q(\levenshtein_ctrl.idx[5] ));
 sg13g2_dfrbp_1 _3121_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net112),
    .D(net557),
    .Q_N(_1424_),
    .Q(\levenshtein_ctrl.idx[6] ));
 sg13g2_dfrbp_1 _3122_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net111),
    .D(net519),
    .Q_N(_1423_),
    .Q(\levenshtein_ctrl.idx[7] ));
 sg13g2_dfrbp_1 _3123_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net110),
    .D(_0169_),
    .Q_N(_1422_),
    .Q(\levenshtein_ctrl.idx[8] ));
 sg13g2_dfrbp_1 _3124_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net109),
    .D(net575),
    .Q_N(_1421_),
    .Q(\levenshtein_ctrl.idx[9] ));
 sg13g2_dfrbp_1 _3125_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net108),
    .D(net530),
    .Q_N(_1420_),
    .Q(\levenshtein_ctrl.idx[10] ));
 sg13g2_dfrbp_1 _3126_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net107),
    .D(_0172_),
    .Q_N(_1419_),
    .Q(\levenshtein_ctrl.idx[11] ));
 sg13g2_dfrbp_1 _3127_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net106),
    .D(_0173_),
    .Q_N(_1418_),
    .Q(\levenshtein_ctrl.idx[12] ));
 sg13g2_dfrbp_1 _3128_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net105),
    .D(net601),
    .Q_N(_1417_),
    .Q(\levenshtein_ctrl.idx[13] ));
 sg13g2_dfrbp_1 _3129_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net104),
    .D(_0175_),
    .Q_N(_1416_),
    .Q(\levenshtein_ctrl.idx[14] ));
 sg13g2_dfrbp_1 _3130_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net103),
    .D(net499),
    .Q_N(_1415_),
    .Q(\levenshtein_ctrl.idx[15] ));
 sg13g2_dfrbp_1 _3131_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net102),
    .D(net465),
    .Q_N(_1414_),
    .Q(\levenshtein_ctrl.best_idx[0] ));
 sg13g2_dfrbp_1 _3132_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net101),
    .D(net533),
    .Q_N(_1413_),
    .Q(\levenshtein_ctrl.best_idx[1] ));
 sg13g2_dfrbp_1 _3133_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net100),
    .D(net303),
    .Q_N(_1412_),
    .Q(\levenshtein_ctrl.best_idx[2] ));
 sg13g2_dfrbp_1 _3134_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net99),
    .D(_0180_),
    .Q_N(_1411_),
    .Q(\levenshtein_ctrl.best_idx[3] ));
 sg13g2_dfrbp_1 _3135_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net98),
    .D(net311),
    .Q_N(_1410_),
    .Q(\levenshtein_ctrl.best_idx[4] ));
 sg13g2_dfrbp_1 _3136_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net97),
    .D(net476),
    .Q_N(_1409_),
    .Q(\levenshtein_ctrl.best_idx[5] ));
 sg13g2_dfrbp_1 _3137_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net96),
    .D(net307),
    .Q_N(_1408_),
    .Q(\levenshtein_ctrl.best_idx[6] ));
 sg13g2_dfrbp_1 _3138_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net95),
    .D(net305),
    .Q_N(_1407_),
    .Q(\levenshtein_ctrl.best_idx[7] ));
 sg13g2_dfrbp_1 _3139_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net94),
    .D(_0185_),
    .Q_N(_1406_),
    .Q(\levenshtein_ctrl.best_idx[8] ));
 sg13g2_dfrbp_1 _3140_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net93),
    .D(net700),
    .Q_N(_1405_),
    .Q(\levenshtein_ctrl.best_idx[9] ));
 sg13g2_dfrbp_1 _3141_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net92),
    .D(_0187_),
    .Q_N(_1404_),
    .Q(\levenshtein_ctrl.best_idx[10] ));
 sg13g2_dfrbp_1 _3142_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net91),
    .D(_0188_),
    .Q_N(_1403_),
    .Q(\levenshtein_ctrl.best_idx[11] ));
 sg13g2_dfrbp_1 _3143_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net90),
    .D(net526),
    .Q_N(_1402_),
    .Q(\levenshtein_ctrl.best_idx[12] ));
 sg13g2_dfrbp_1 _3144_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net89),
    .D(net472),
    .Q_N(_1401_),
    .Q(\levenshtein_ctrl.best_idx[13] ));
 sg13g2_dfrbp_1 _3145_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net88),
    .D(net492),
    .Q_N(_1400_),
    .Q(\levenshtein_ctrl.best_idx[14] ));
 sg13g2_dfrbp_1 _3146_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net87),
    .D(net474),
    .Q_N(_1399_),
    .Q(\levenshtein_ctrl.best_idx[15] ));
 sg13g2_dfrbp_1 _3147_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net86),
    .D(net516),
    .Q_N(_1398_),
    .Q(\levenshtein_ctrl.best_distance[0] ));
 sg13g2_dfrbp_1 _3148_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net85),
    .D(_0194_),
    .Q_N(_1397_),
    .Q(\levenshtein_ctrl.best_distance[1] ));
 sg13g2_dfrbp_1 _3149_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net84),
    .D(net702),
    .Q_N(_1396_),
    .Q(\levenshtein_ctrl.best_distance[2] ));
 sg13g2_dfrbp_1 _3150_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net83),
    .D(net710),
    .Q_N(_1395_),
    .Q(\levenshtein_ctrl.best_distance[3] ));
 sg13g2_dfrbp_1 _3151_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net82),
    .D(net579),
    .Q_N(_1394_),
    .Q(\levenshtein_ctrl.best_distance[4] ));
 sg13g2_dfrbp_1 _3152_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net81),
    .D(net539),
    .Q_N(_1393_),
    .Q(\levenshtein_ctrl.best_distance[5] ));
 sg13g2_dfrbp_1 _3153_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net80),
    .D(net542),
    .Q_N(_1392_),
    .Q(\levenshtein_ctrl.best_distance[6] ));
 sg13g2_dfrbp_1 _3154_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net79),
    .D(net569),
    .Q_N(_1391_),
    .Q(\levenshtein_ctrl.best_distance[7] ));
 sg13g2_dfrbp_1 _3155_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net78),
    .D(net444),
    .Q_N(_1390_),
    .Q(\levenshtein_ctrl.next_symbol[0] ));
 sg13g2_dfrbp_1 _3156_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net77),
    .D(_0202_),
    .Q_N(_1389_),
    .Q(\levenshtein_ctrl.next_symbol[1] ));
 sg13g2_dfrbp_1 _3157_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net76),
    .D(_0203_),
    .Q_N(_1388_),
    .Q(\levenshtein_ctrl.next_symbol[2] ));
 sg13g2_dfrbp_1 _3158_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net75),
    .D(net446),
    .Q_N(_1387_),
    .Q(\levenshtein_ctrl.next_symbol[3] ));
 sg13g2_dfrbp_1 _3159_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net74),
    .D(_0205_),
    .Q_N(_1386_),
    .Q(\levenshtein_ctrl.next_symbol[4] ));
 sg13g2_dfrbp_1 _3160_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net73),
    .D(_0206_),
    .Q_N(_1385_),
    .Q(\levenshtein_ctrl.next_symbol[5] ));
 sg13g2_dfrbp_1 _3161_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net72),
    .D(_0207_),
    .Q_N(_1384_),
    .Q(\levenshtein_ctrl.next_symbol[6] ));
 sg13g2_dfrbp_1 _3162_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net71),
    .D(_0208_),
    .Q_N(_1383_),
    .Q(\levenshtein_ctrl.next_symbol[7] ));
 sg13g2_dfrbp_1 _3163_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net70),
    .D(_0209_),
    .Q_N(_1382_),
    .Q(\levenshtein_ctrl.symbols[8] ));
 sg13g2_dfrbp_1 _3164_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net69),
    .D(_0210_),
    .Q_N(_1381_),
    .Q(\levenshtein_ctrl.symbols[9] ));
 sg13g2_dfrbp_1 _3165_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net68),
    .D(_0211_),
    .Q_N(_1380_),
    .Q(\levenshtein_ctrl.symbols[10] ));
 sg13g2_dfrbp_1 _3166_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net67),
    .D(_0212_),
    .Q_N(_1379_),
    .Q(\levenshtein_ctrl.symbols[11] ));
 sg13g2_dfrbp_1 _3167_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net66),
    .D(_0213_),
    .Q_N(_1378_),
    .Q(\levenshtein_ctrl.symbols[12] ));
 sg13g2_dfrbp_1 _3168_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net65),
    .D(_0214_),
    .Q_N(_1377_),
    .Q(\levenshtein_ctrl.symbols[13] ));
 sg13g2_dfrbp_1 _3169_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net64),
    .D(_0215_),
    .Q_N(_1376_),
    .Q(\levenshtein_ctrl.symbols[14] ));
 sg13g2_dfrbp_1 _3170_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net63),
    .D(_0216_),
    .Q_N(_1375_),
    .Q(\levenshtein_ctrl.symbols[15] ));
 sg13g2_dfrbp_1 _3171_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net62),
    .D(net296),
    .Q_N(_1374_),
    .Q(\levenshtein_ctrl.symbols[16] ));
 sg13g2_dfrbp_1 _3172_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net61),
    .D(net282),
    .Q_N(_1373_),
    .Q(\levenshtein_ctrl.symbols[17] ));
 sg13g2_dfrbp_1 _3173_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net60),
    .D(net274),
    .Q_N(_1372_),
    .Q(\levenshtein_ctrl.symbols[18] ));
 sg13g2_dfrbp_1 _3174_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net59),
    .D(net313),
    .Q_N(_1371_),
    .Q(\levenshtein_ctrl.symbols[19] ));
 sg13g2_dfrbp_1 _3175_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net58),
    .D(net272),
    .Q_N(_1370_),
    .Q(\levenshtein_ctrl.symbols[20] ));
 sg13g2_dfrbp_1 _3176_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net57),
    .D(net291),
    .Q_N(_1369_),
    .Q(\levenshtein_ctrl.symbols[21] ));
 sg13g2_dfrbp_1 _3177_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net56),
    .D(net278),
    .Q_N(_1368_),
    .Q(\levenshtein_ctrl.symbols[22] ));
 sg13g2_dfrbp_1 _3178_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net55),
    .D(net276),
    .Q_N(_1367_),
    .Q(\levenshtein_ctrl.symbols[23] ));
 sg13g2_dfrbp_1 _3179_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net54),
    .D(net315),
    .Q_N(_0028_),
    .Q(\levenshtein_ctrl.symbol[0] ));
 sg13g2_dfrbp_1 _3180_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net53),
    .D(_0226_),
    .Q_N(_0027_),
    .Q(\levenshtein_ctrl.symbol[1] ));
 sg13g2_dfrbp_1 _3181_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net52),
    .D(_0227_),
    .Q_N(_0026_),
    .Q(\levenshtein_ctrl.symbol[2] ));
 sg13g2_dfrbp_1 _3182_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net51),
    .D(_0228_),
    .Q_N(_0025_),
    .Q(\levenshtein_ctrl.symbol[3] ));
 sg13g2_dfrbp_1 _3183_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net50),
    .D(net321),
    .Q_N(_0024_),
    .Q(\levenshtein_ctrl.symbol[4] ));
 sg13g2_dfrbp_1 _3184_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net49),
    .D(net323),
    .Q_N(_0023_),
    .Q(\levenshtein_ctrl.symbol[5] ));
 sg13g2_dfrbp_1 _3185_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net48),
    .D(net479),
    .Q_N(_0022_),
    .Q(\levenshtein_ctrl.symbol[6] ));
 sg13g2_dfrbp_1 _3186_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net47),
    .D(net440),
    .Q_N(_0021_),
    .Q(\levenshtein_ctrl.symbol[7] ));
 sg13g2_dfrbp_1 _3187_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net46),
    .D(_0233_),
    .Q_N(_1366_),
    .Q(\levenshtein_ctrl.pm[8] ));
 sg13g2_dfrbp_1 _3188_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net45),
    .D(net550),
    .Q_N(_1365_),
    .Q(\levenshtein_ctrl.pm[9] ));
 sg13g2_dfrbp_1 _3189_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net44),
    .D(_0235_),
    .Q_N(_1364_),
    .Q(\levenshtein_ctrl.pm[10] ));
 sg13g2_dfrbp_1 _3190_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net43),
    .D(net587),
    .Q_N(_1363_),
    .Q(\levenshtein_ctrl.pm[11] ));
 sg13g2_dfrbp_1 _3191_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net42),
    .D(net631),
    .Q_N(_1362_),
    .Q(\levenshtein_ctrl.pm[12] ));
 sg13g2_dfrbp_1 _3192_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net41),
    .D(net489),
    .Q_N(_1361_),
    .Q(\levenshtein_ctrl.pm[13] ));
 sg13g2_dfrbp_1 _3193_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net40),
    .D(_0239_),
    .Q_N(_1360_),
    .Q(\levenshtein_ctrl.pm[14] ));
 sg13g2_dfrbp_1 _3194_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net39),
    .D(_0240_),
    .Q_N(_1359_),
    .Q(\levenshtein_ctrl.pm[15] ));
 sg13g2_dfrbp_1 _3195_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net36),
    .D(net663),
    .Q_N(_1358_),
    .Q(\arbiter.wbs0_dat_i[1] ));
 sg13g2_dfrbp_1 _3196_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net31),
    .D(net629),
    .Q_N(_1357_),
    .Q(\arbiter.wbs0_dat_i[2] ));
 sg13g2_dfrbp_1 _3197_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net30),
    .D(_0243_),
    .Q_N(_1356_),
    .Q(\arbiter.wbs0_dat_i[3] ));
 sg13g2_dfrbp_1 _3198_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net29),
    .D(net507),
    .Q_N(_1355_),
    .Q(\arbiter.wbs0_dat_i[4] ));
 sg13g2_dfrbp_1 _3199_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net27),
    .D(_0245_),
    .Q_N(_1354_),
    .Q(\arbiter.wbs0_dat_i[5] ));
 sg13g2_dfrbp_1 _3200_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net26),
    .D(net486),
    .Q_N(_1353_),
    .Q(\arbiter.wbs0_dat_i[6] ));
 sg13g2_dfrbp_1 _3201_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net25),
    .D(_0247_),
    .Q_N(_1352_),
    .Q(\arbiter.wbs0_dat_i[7] ));
 sg13g2_dfrbp_1 _3202_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net24),
    .D(_0248_),
    .Q_N(_1351_),
    .Q(\arbiter.wbs0_adr_i[0] ));
 sg13g2_dfrbp_1 _3203_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net23),
    .D(_0249_),
    .Q_N(_1350_),
    .Q(uio_oe[1]));
 sg13g2_dfrbp_1 _3204_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net15),
    .D(_0250_),
    .Q_N(_1349_),
    .Q(uio_oe[2]));
 sg13g2_dfrbp_1 _3205_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net256),
    .D(_0251_),
    .Q_N(_1348_),
    .Q(uio_oe[4]));
 sg13g2_dfrbp_1 _3206_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net255),
    .D(_0252_),
    .Q_N(_1347_),
    .Q(uio_oe[5]));
 sg13g2_dfrbp_1 _3207_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net252),
    .D(net280),
    .Q_N(_1346_),
    .Q(\arbiter.wbm_ack_i ));
 sg13g2_dfrbp_1 _3208_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net251),
    .D(_0254_),
    .Q_N(_1345_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _3209_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net249),
    .D(_0255_),
    .Q_N(_1344_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _3210_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net247),
    .D(_0256_),
    .Q_N(_1343_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _3211_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net245),
    .D(_0257_),
    .Q_N(_0020_),
    .Q(\spi_ctrl.sck ));
 sg13g2_dfrbp_1 _3212_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net243),
    .D(_0258_),
    .Q_N(_1342_),
    .Q(\arbiter.wbm_dat_i[0] ));
 sg13g2_dfrbp_1 _3213_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net242),
    .D(_0259_),
    .Q_N(_1341_),
    .Q(\arbiter.wbm_dat_i[1] ));
 sg13g2_dfrbp_1 _3214_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net241),
    .D(_0260_),
    .Q_N(_1340_),
    .Q(\arbiter.wbm_dat_i[2] ));
 sg13g2_dfrbp_1 _3215_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net240),
    .D(_0261_),
    .Q_N(_1339_),
    .Q(\arbiter.wbm_dat_i[3] ));
 sg13g2_dfrbp_1 _3216_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net239),
    .D(_0262_),
    .Q_N(_1338_),
    .Q(\arbiter.wbm_dat_i[4] ));
 sg13g2_dfrbp_1 _3217_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net238),
    .D(net755),
    .Q_N(_1337_),
    .Q(\arbiter.wbm_dat_i[5] ));
 sg13g2_dfrbp_1 _3218_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net237),
    .D(_0264_),
    .Q_N(_1336_),
    .Q(\arbiter.wbm_dat_i[6] ));
 sg13g2_dfrbp_1 _3219_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net236),
    .D(_0265_),
    .Q_N(_1335_),
    .Q(\arbiter.wbm_dat_i[7] ));
 sg13g2_dfrbp_1 _3220_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net235),
    .D(_0266_),
    .Q_N(_0019_),
    .Q(\arbiter.wbs0_adr_i[1] ));
 sg13g2_dfrbp_1 _3221_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net234),
    .D(net589),
    .Q_N(_0018_),
    .Q(\arbiter.wbs0_adr_i[2] ));
 sg13g2_dfrbp_1 _3222_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net233),
    .D(net653),
    .Q_N(_0017_),
    .Q(\arbiter.wbs0_adr_i[3] ));
 sg13g2_dfrbp_1 _3223_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net232),
    .D(net599),
    .Q_N(_0016_),
    .Q(\arbiter.wbs0_adr_i[4] ));
 sg13g2_dfrbp_1 _3224_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net231),
    .D(net562),
    .Q_N(_0015_),
    .Q(\arbiter.wbs0_adr_i[5] ));
 sg13g2_dfrbp_1 _3225_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net230),
    .D(net505),
    .Q_N(_0014_),
    .Q(\arbiter.wbs0_adr_i[6] ));
 sg13g2_dfrbp_1 _3226_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net229),
    .D(_0272_),
    .Q_N(_0013_),
    .Q(\arbiter.wbs0_adr_i[7] ));
 sg13g2_dfrbp_1 _3227_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net228),
    .D(_0273_),
    .Q_N(_0012_),
    .Q(\arbiter.wbs0_adr_i[8] ));
 sg13g2_dfrbp_1 _3228_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net227),
    .D(_0274_),
    .Q_N(_1334_),
    .Q(\arbiter.wbs0_adr_i[9] ));
 sg13g2_dfrbp_1 _3229_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net226),
    .D(net637),
    .Q_N(_1333_),
    .Q(\arbiter.wbs0_adr_i[10] ));
 sg13g2_dfrbp_1 _3230_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net225),
    .D(net503),
    .Q_N(_1332_),
    .Q(\arbiter.wbs0_adr_i[11] ));
 sg13g2_dfrbp_1 _3231_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net224),
    .D(_0277_),
    .Q_N(_1331_),
    .Q(\arbiter.wbs0_adr_i[12] ));
 sg13g2_dfrbp_1 _3232_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net223),
    .D(_0278_),
    .Q_N(_1330_),
    .Q(\arbiter.wbs0_adr_i[13] ));
 sg13g2_dfrbp_1 _3233_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net221),
    .D(net640),
    .Q_N(_1329_),
    .Q(\arbiter.wbs0_adr_i[14] ));
 sg13g2_dfrbp_1 _3234_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net219),
    .D(net633),
    .Q_N(_1328_),
    .Q(\arbiter.wbs0_adr_i[15] ));
 sg13g2_dfrbp_1 _3235_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net217),
    .D(net605),
    .Q_N(_1327_),
    .Q(\arbiter.wbs0_adr_i[16] ));
 sg13g2_dfrbp_1 _3236_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net215),
    .D(net603),
    .Q_N(_1326_),
    .Q(\arbiter.wbs0_adr_i[17] ));
 sg13g2_dfrbp_1 _3237_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net213),
    .D(_0283_),
    .Q_N(_1325_),
    .Q(\arbiter.wbs0_adr_i[18] ));
 sg13g2_dfrbp_1 _3238_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net209),
    .D(_0284_),
    .Q_N(_1324_),
    .Q(\arbiter.wbs0_adr_i[19] ));
 sg13g2_dfrbp_1 _3239_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net207),
    .D(_0285_),
    .Q_N(_1323_),
    .Q(\arbiter.wbs0_adr_i[20] ));
 sg13g2_dfrbp_1 _3240_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net205),
    .D(net682),
    .Q_N(_1322_),
    .Q(\arbiter.wbs0_adr_i[21] ));
 sg13g2_dfrbp_1 _3241_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net203),
    .D(_0287_),
    .Q_N(_1321_),
    .Q(\arbiter.wbs0_adr_i[22] ));
 sg13g2_dfrbp_1 _3242_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net201),
    .D(net612),
    .Q_N(_1320_),
    .Q(\arbiter.wbs0_we_i ));
 sg13g2_dfrbp_1 _3243_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net194),
    .D(_0289_),
    .Q_N(_1319_),
    .Q(\spi_ctrl.bit_counter[2] ));
 sg13g2_dfrbp_1 _3244_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net254),
    .D(net635),
    .Q_N(_0066_),
    .Q(\spi_ctrl.bit_counter[4] ));
 sg13g2_dfrbp_1 _3245_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net250),
    .D(_0008_),
    .Q_N(_0067_),
    .Q(\spi.state[0] ));
 sg13g2_dfrbp_1 _3246_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net248),
    .D(net672),
    .Q_N(_0011_),
    .Q(\spi.state[2] ));
 sg13g2_dfrbp_1 _3247_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net244),
    .D(_0291_),
    .Q_N(_0010_),
    .Q(\arbiter.gnt ));
 sg13g2_dfrbp_1 _3248_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net246),
    .D(net666),
    .Q_N(_1318_),
    .Q(\arbiter.wbs0_dat_i[0] ));
 sg13g2_tiehi _3014__16 (.L_HI(net16));
 sg13g2_tiehi _3007__17 (.L_HI(net17));
 sg13g2_tiehi _3008__18 (.L_HI(net18));
 sg13g2_tiehi _3009__19 (.L_HI(net19));
 sg13g2_tiehi _3010__20 (.L_HI(net20));
 sg13g2_tiehi _3011__21 (.L_HI(net21));
 sg13g2_tiehi _3012__22 (.L_HI(net22));
 sg13g2_tiehi _3203__23 (.L_HI(net23));
 sg13g2_tiehi _3202__24 (.L_HI(net24));
 sg13g2_tiehi _3201__25 (.L_HI(net25));
 sg13g2_tiehi _3200__26 (.L_HI(net26));
 sg13g2_tiehi _3199__27 (.L_HI(net27));
 sg13g2_tiehi _3013__28 (.L_HI(net28));
 sg13g2_tiehi _3198__29 (.L_HI(net29));
 sg13g2_tiehi _3197__30 (.L_HI(net30));
 sg13g2_tiehi _3196__31 (.L_HI(net31));
 sg13g2_tiehi _3019__32 (.L_HI(net32));
 sg13g2_tiehi _3023__33 (.L_HI(net33));
 sg13g2_tiehi _3024__34 (.L_HI(net34));
 sg13g2_tiehi _3025__35 (.L_HI(net35));
 sg13g2_tiehi _3195__36 (.L_HI(net36));
 sg13g2_tiehi _3026__37 (.L_HI(net37));
 sg13g2_tiehi _3028__38 (.L_HI(net38));
 sg13g2_tiehi _3194__39 (.L_HI(net39));
 sg13g2_tiehi _3193__40 (.L_HI(net40));
 sg13g2_tiehi _3192__41 (.L_HI(net41));
 sg13g2_tiehi _3191__42 (.L_HI(net42));
 sg13g2_tiehi _3190__43 (.L_HI(net43));
 sg13g2_tiehi _3189__44 (.L_HI(net44));
 sg13g2_tiehi _3188__45 (.L_HI(net45));
 sg13g2_tiehi _3187__46 (.L_HI(net46));
 sg13g2_tiehi _3186__47 (.L_HI(net47));
 sg13g2_tiehi _3185__48 (.L_HI(net48));
 sg13g2_tiehi _3184__49 (.L_HI(net49));
 sg13g2_tiehi _3183__50 (.L_HI(net50));
 sg13g2_tiehi _3182__51 (.L_HI(net51));
 sg13g2_tiehi _3181__52 (.L_HI(net52));
 sg13g2_tiehi _3180__53 (.L_HI(net53));
 sg13g2_tiehi _3179__54 (.L_HI(net54));
 sg13g2_tiehi _3178__55 (.L_HI(net55));
 sg13g2_tiehi _3177__56 (.L_HI(net56));
 sg13g2_tiehi _3176__57 (.L_HI(net57));
 sg13g2_tiehi _3175__58 (.L_HI(net58));
 sg13g2_tiehi _3174__59 (.L_HI(net59));
 sg13g2_tiehi _3173__60 (.L_HI(net60));
 sg13g2_tiehi _3172__61 (.L_HI(net61));
 sg13g2_tiehi _3171__62 (.L_HI(net62));
 sg13g2_tiehi _3170__63 (.L_HI(net63));
 sg13g2_tiehi _3169__64 (.L_HI(net64));
 sg13g2_tiehi _3168__65 (.L_HI(net65));
 sg13g2_tiehi _3167__66 (.L_HI(net66));
 sg13g2_tiehi _3166__67 (.L_HI(net67));
 sg13g2_tiehi _3165__68 (.L_HI(net68));
 sg13g2_tiehi _3164__69 (.L_HI(net69));
 sg13g2_tiehi _3163__70 (.L_HI(net70));
 sg13g2_tiehi _3162__71 (.L_HI(net71));
 sg13g2_tiehi _3161__72 (.L_HI(net72));
 sg13g2_tiehi _3160__73 (.L_HI(net73));
 sg13g2_tiehi _3159__74 (.L_HI(net74));
 sg13g2_tiehi _3158__75 (.L_HI(net75));
 sg13g2_tiehi _3157__76 (.L_HI(net76));
 sg13g2_tiehi _3156__77 (.L_HI(net77));
 sg13g2_tiehi _3155__78 (.L_HI(net78));
 sg13g2_tiehi _3154__79 (.L_HI(net79));
 sg13g2_tiehi _3153__80 (.L_HI(net80));
 sg13g2_tiehi _3152__81 (.L_HI(net81));
 sg13g2_tiehi _3151__82 (.L_HI(net82));
 sg13g2_tiehi _3150__83 (.L_HI(net83));
 sg13g2_tiehi _3149__84 (.L_HI(net84));
 sg13g2_tiehi _3148__85 (.L_HI(net85));
 sg13g2_tiehi _3147__86 (.L_HI(net86));
 sg13g2_tiehi _3146__87 (.L_HI(net87));
 sg13g2_tiehi _3145__88 (.L_HI(net88));
 sg13g2_tiehi _3144__89 (.L_HI(net89));
 sg13g2_tiehi _3143__90 (.L_HI(net90));
 sg13g2_tiehi _3142__91 (.L_HI(net91));
 sg13g2_tiehi _3141__92 (.L_HI(net92));
 sg13g2_tiehi _3140__93 (.L_HI(net93));
 sg13g2_tiehi _3139__94 (.L_HI(net94));
 sg13g2_tiehi _3138__95 (.L_HI(net95));
 sg13g2_tiehi _3137__96 (.L_HI(net96));
 sg13g2_tiehi _3136__97 (.L_HI(net97));
 sg13g2_tiehi _3135__98 (.L_HI(net98));
 sg13g2_tiehi _3134__99 (.L_HI(net99));
 sg13g2_tiehi _3133__100 (.L_HI(net100));
 sg13g2_tiehi _3132__101 (.L_HI(net101));
 sg13g2_tiehi _3131__102 (.L_HI(net102));
 sg13g2_tiehi _3130__103 (.L_HI(net103));
 sg13g2_tiehi _3129__104 (.L_HI(net104));
 sg13g2_tiehi _3128__105 (.L_HI(net105));
 sg13g2_tiehi _3127__106 (.L_HI(net106));
 sg13g2_tiehi _3126__107 (.L_HI(net107));
 sg13g2_tiehi _3125__108 (.L_HI(net108));
 sg13g2_tiehi _3124__109 (.L_HI(net109));
 sg13g2_tiehi _3123__110 (.L_HI(net110));
 sg13g2_tiehi _3122__111 (.L_HI(net111));
 sg13g2_tiehi _3121__112 (.L_HI(net112));
 sg13g2_tiehi _3120__113 (.L_HI(net113));
 sg13g2_tiehi _3119__114 (.L_HI(net114));
 sg13g2_tiehi _3118__115 (.L_HI(net115));
 sg13g2_tiehi _3117__116 (.L_HI(net116));
 sg13g2_tiehi _3116__117 (.L_HI(net117));
 sg13g2_tiehi _3115__118 (.L_HI(net118));
 sg13g2_tiehi _3114__119 (.L_HI(net119));
 sg13g2_tiehi _3113__120 (.L_HI(net120));
 sg13g2_tiehi _3112__121 (.L_HI(net121));
 sg13g2_tiehi _3111__122 (.L_HI(net122));
 sg13g2_tiehi _3110__123 (.L_HI(net123));
 sg13g2_tiehi _3109__124 (.L_HI(net124));
 sg13g2_tiehi _3108__125 (.L_HI(net125));
 sg13g2_tiehi _3107__126 (.L_HI(net126));
 sg13g2_tiehi _3106__127 (.L_HI(net127));
 sg13g2_tiehi _3105__128 (.L_HI(net128));
 sg13g2_tiehi _3104__129 (.L_HI(net129));
 sg13g2_tiehi _3103__130 (.L_HI(net130));
 sg13g2_tiehi _3102__131 (.L_HI(net131));
 sg13g2_tiehi _3101__132 (.L_HI(net132));
 sg13g2_tiehi _3100__133 (.L_HI(net133));
 sg13g2_tiehi _3099__134 (.L_HI(net134));
 sg13g2_tiehi _3098__135 (.L_HI(net135));
 sg13g2_tiehi _3097__136 (.L_HI(net136));
 sg13g2_tiehi _3096__137 (.L_HI(net137));
 sg13g2_tiehi _3095__138 (.L_HI(net138));
 sg13g2_tiehi _3094__139 (.L_HI(net139));
 sg13g2_tiehi _3093__140 (.L_HI(net140));
 sg13g2_tiehi _3092__141 (.L_HI(net141));
 sg13g2_tiehi _3091__142 (.L_HI(net142));
 sg13g2_tiehi _3090__143 (.L_HI(net143));
 sg13g2_tiehi _3089__144 (.L_HI(net144));
 sg13g2_tiehi _3088__145 (.L_HI(net145));
 sg13g2_tiehi _3087__146 (.L_HI(net146));
 sg13g2_tiehi _3086__147 (.L_HI(net147));
 sg13g2_tiehi _3085__148 (.L_HI(net148));
 sg13g2_tiehi _3084__149 (.L_HI(net149));
 sg13g2_tiehi _3083__150 (.L_HI(net150));
 sg13g2_tiehi _3082__151 (.L_HI(net151));
 sg13g2_tiehi _3081__152 (.L_HI(net152));
 sg13g2_tiehi _3080__153 (.L_HI(net153));
 sg13g2_tiehi _3079__154 (.L_HI(net154));
 sg13g2_tiehi _3078__155 (.L_HI(net155));
 sg13g2_tiehi _3077__156 (.L_HI(net156));
 sg13g2_tiehi _3076__157 (.L_HI(net157));
 sg13g2_tiehi _3075__158 (.L_HI(net158));
 sg13g2_tiehi _3074__159 (.L_HI(net159));
 sg13g2_tiehi _3073__160 (.L_HI(net160));
 sg13g2_tiehi _3072__161 (.L_HI(net161));
 sg13g2_tiehi _3071__162 (.L_HI(net162));
 sg13g2_tiehi _3070__163 (.L_HI(net163));
 sg13g2_tiehi _3069__164 (.L_HI(net164));
 sg13g2_tiehi _3068__165 (.L_HI(net165));
 sg13g2_tiehi _3067__166 (.L_HI(net166));
 sg13g2_tiehi _3066__167 (.L_HI(net167));
 sg13g2_tiehi _3065__168 (.L_HI(net168));
 sg13g2_tiehi _3064__169 (.L_HI(net169));
 sg13g2_tiehi _3063__170 (.L_HI(net170));
 sg13g2_tiehi _3062__171 (.L_HI(net171));
 sg13g2_tiehi _3061__172 (.L_HI(net172));
 sg13g2_tiehi _3060__173 (.L_HI(net173));
 sg13g2_tiehi _3059__174 (.L_HI(net174));
 sg13g2_tiehi _3058__175 (.L_HI(net175));
 sg13g2_tiehi _3057__176 (.L_HI(net176));
 sg13g2_tiehi _3056__177 (.L_HI(net177));
 sg13g2_tiehi _3055__178 (.L_HI(net178));
 sg13g2_tiehi _3054__179 (.L_HI(net179));
 sg13g2_tiehi _3053__180 (.L_HI(net180));
 sg13g2_tiehi _3052__181 (.L_HI(net181));
 sg13g2_tiehi _3051__182 (.L_HI(net182));
 sg13g2_tiehi _3050__183 (.L_HI(net183));
 sg13g2_tiehi _3049__184 (.L_HI(net184));
 sg13g2_tiehi _3048__185 (.L_HI(net185));
 sg13g2_tiehi _3047__186 (.L_HI(net186));
 sg13g2_tiehi _3046__187 (.L_HI(net187));
 sg13g2_tiehi _3045__188 (.L_HI(net188));
 sg13g2_tiehi _3044__189 (.L_HI(net189));
 sg13g2_tiehi _3043__190 (.L_HI(net190));
 sg13g2_tiehi _3042__191 (.L_HI(net191));
 sg13g2_tiehi _3041__192 (.L_HI(net192));
 sg13g2_tiehi _3040__193 (.L_HI(net193));
 sg13g2_tiehi _3243__194 (.L_HI(net194));
 sg13g2_tiehi _3039__195 (.L_HI(net195));
 sg13g2_tiehi _3038__196 (.L_HI(net196));
 sg13g2_tiehi _3037__197 (.L_HI(net197));
 sg13g2_tiehi _3036__198 (.L_HI(net198));
 sg13g2_tiehi _3035__199 (.L_HI(net199));
 sg13g2_tiehi _3034__200 (.L_HI(net200));
 sg13g2_tiehi _3242__201 (.L_HI(net201));
 sg13g2_tiehi _3033__202 (.L_HI(net202));
 sg13g2_tiehi _3241__203 (.L_HI(net203));
 sg13g2_tiehi _3032__204 (.L_HI(net204));
 sg13g2_tiehi _3240__205 (.L_HI(net205));
 sg13g2_tiehi _3031__206 (.L_HI(net206));
 sg13g2_tiehi _3239__207 (.L_HI(net207));
 sg13g2_tiehi _3030__208 (.L_HI(net208));
 sg13g2_tiehi _3238__209 (.L_HI(net209));
 sg13g2_tiehi _3027__210 (.L_HI(net210));
 sg13g2_tiehi _3022__211 (.L_HI(net211));
 sg13g2_tiehi _3021__212 (.L_HI(net212));
 sg13g2_tiehi _3237__213 (.L_HI(net213));
 sg13g2_tiehi _3020__214 (.L_HI(net214));
 sg13g2_tiehi _3236__215 (.L_HI(net215));
 sg13g2_tiehi _3018__216 (.L_HI(net216));
 sg13g2_tiehi _3235__217 (.L_HI(net217));
 sg13g2_tiehi _3017__218 (.L_HI(net218));
 sg13g2_tiehi _3234__219 (.L_HI(net219));
 sg13g2_tiehi _3016__220 (.L_HI(net220));
 sg13g2_tiehi _3233__221 (.L_HI(net221));
 sg13g2_tiehi _3015__222 (.L_HI(net222));
 sg13g2_tiehi _3232__223 (.L_HI(net223));
 sg13g2_tiehi _3231__224 (.L_HI(net224));
 sg13g2_tiehi _3230__225 (.L_HI(net225));
 sg13g2_tiehi _3229__226 (.L_HI(net226));
 sg13g2_tiehi _3228__227 (.L_HI(net227));
 sg13g2_tiehi _3227__228 (.L_HI(net228));
 sg13g2_tiehi _3226__229 (.L_HI(net229));
 sg13g2_tiehi _3225__230 (.L_HI(net230));
 sg13g2_tiehi _3224__231 (.L_HI(net231));
 sg13g2_tiehi _3223__232 (.L_HI(net232));
 sg13g2_tiehi _3222__233 (.L_HI(net233));
 sg13g2_tiehi _3221__234 (.L_HI(net234));
 sg13g2_tiehi _3220__235 (.L_HI(net235));
 sg13g2_tiehi _3219__236 (.L_HI(net236));
 sg13g2_tiehi _3218__237 (.L_HI(net237));
 sg13g2_tiehi _3217__238 (.L_HI(net238));
 sg13g2_tiehi _3216__239 (.L_HI(net239));
 sg13g2_tiehi _3215__240 (.L_HI(net240));
 sg13g2_tiehi _3214__241 (.L_HI(net241));
 sg13g2_tiehi _3213__242 (.L_HI(net242));
 sg13g2_tiehi _3212__243 (.L_HI(net243));
 sg13g2_tiehi _3247__244 (.L_HI(net244));
 sg13g2_tiehi _3211__245 (.L_HI(net245));
 sg13g2_tiehi _3248__246 (.L_HI(net246));
 sg13g2_tiehi _3210__247 (.L_HI(net247));
 sg13g2_tiehi _3246__248 (.L_HI(net248));
 sg13g2_tiehi _3209__249 (.L_HI(net249));
 sg13g2_tiehi _3245__250 (.L_HI(net250));
 sg13g2_tiehi _3208__251 (.L_HI(net251));
 sg13g2_tiehi _3207__252 (.L_HI(net252));
 sg13g2_tiehi _3029__253 (.L_HI(net253));
 sg13g2_tiehi _3244__254 (.L_HI(net254));
 sg13g2_tiehi _3206__255 (.L_HI(net255));
 sg13g2_tiehi _3205__256 (.L_HI(net256));
 sg13g2_tiehi tt_um_levenshtein_257 (.L_HI(net257));
 sg13g2_tiehi tt_um_levenshtein_258 (.L_HI(net258));
 sg13g2_tiehi tt_um_levenshtein_259 (.L_HI(net259));
 sg13g2_tiehi tt_um_levenshtein_260 (.L_HI(net260));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_levenshtein_9 (.L_LO(net9));
 sg13g2_tielo tt_um_levenshtein_10 (.L_LO(net10));
 sg13g2_tielo tt_um_levenshtein_11 (.L_LO(net11));
 sg13g2_tielo tt_um_levenshtein_12 (.L_LO(net12));
 sg13g2_tielo tt_um_levenshtein_13 (.L_LO(net13));
 sg13g2_tielo tt_um_levenshtein_14 (.L_LO(net14));
 sg13g2_tiehi _3204__15 (.L_HI(net15));
 sg13g2_buf_2 _3502_ (.A(\spi_ctrl.cs_n ),
    .X(uio_out[0]));
 sg13g2_buf_1 _3503_ (.A(net408),
    .X(uio_out[3]));
 sg13g2_buf_2 _3504_ (.A(\spi_ctrl.cs2_n ),
    .X(uio_out[6]));
 sg13g2_buf_2 _3505_ (.A(\spi_ctrl.cs3_n ),
    .X(uio_out[7]));
 sg13g2_buf_1 _3506_ (.A(\spi.miso ),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout328 (.A(net329),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(net330),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_0657_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(net332),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_1 fanout333 (.A(_0656_),
    .X(net333));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(_0299_));
 sg13g2_buf_2 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_0299_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_0906_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(net340),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(net340),
    .X(net339));
 sg13g2_buf_1 fanout340 (.A(_0736_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(net342),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(net343),
    .X(net342));
 sg13g2_buf_1 fanout343 (.A(net346),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(net345),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(net346),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_1076_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(net349),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(net349),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_1075_),
    .X(net349));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(_1298_));
 sg13g2_buf_2 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_1095_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(net355),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(net355),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(net359),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(net358),
    .X(net356));
 sg13g2_buf_1 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(net359),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_1083_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(net361),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(net365),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(net364),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(net365),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_0709_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_1287_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_1182_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(net370),
    .X(net368));
 sg13g2_buf_1 fanout369 (.A(net370),
    .X(net369));
 sg13g2_buf_1 fanout370 (.A(net371),
    .X(net370));
 sg13g2_buf_1 fanout371 (.A(_0999_),
    .X(net371));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(net374));
 sg13g2_buf_2 fanout373 (.A(net374),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(net375),
    .X(net374));
 sg13g2_buf_4 fanout375 (.X(net375),
    .A(net376));
 sg13g2_buf_4 fanout376 (.X(net376),
    .A(_0909_));
 sg13g2_buf_4 fanout377 (.X(net377),
    .A(_0734_));
 sg13g2_buf_4 fanout378 (.X(net378),
    .A(net379));
 sg13g2_buf_4 fanout379 (.X(net379),
    .A(_1292_));
 sg13g2_buf_4 fanout380 (.X(net380),
    .A(net383));
 sg13g2_buf_2 fanout381 (.A(net383),
    .X(net381));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(net383));
 sg13g2_buf_2 fanout383 (.A(_1291_),
    .X(net383));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(_1260_));
 sg13g2_buf_2 fanout385 (.A(_1146_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(net387),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(net388),
    .X(net387));
 sg13g2_buf_1 fanout388 (.A(net389),
    .X(net388));
 sg13g2_buf_1 fanout389 (.A(_1111_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(net391),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_1111_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_1110_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_1056_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_1015_),
    .X(net394));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(_1005_));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(net397));
 sg13g2_buf_2 fanout397 (.A(_0990_),
    .X(net397));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(_0933_));
 sg13g2_buf_2 fanout399 (.A(_0929_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_0929_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(\arbiter.gnt ),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(net403),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(net404),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(\arbiter.gnt ),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(\spi_ctrl.bit_counter[2] ),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(net408),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(net708),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(net410),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(\levenshtein_ctrl.word_length_reg[3] ),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(net413),
    .X(net412));
 sg13g2_buf_1 fanout413 (.A(net649),
    .X(net413));
 sg13g2_buf_4 fanout414 (.X(net414),
    .A(net673));
 sg13g2_buf_2 fanout415 (.A(\levenshtein_ctrl.word_length_reg[1] ),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(\levenshtein_ctrl.enabled ),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(net753),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(net421),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(net421),
    .X(net419));
 sg13g2_buf_1 fanout420 (.A(net421),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(\spi_ctrl.bit_counter[0] ),
    .X(net421));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(net688));
 sg13g2_buf_4 fanout423 (.X(net423),
    .A(net570));
 sg13g2_buf_2 fanout424 (.A(net425),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(\levenshtein_ctrl.state[0] ),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(net428),
    .X(net426));
 sg13g2_buf_1 fanout427 (.A(net428),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_0972_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(net431));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(_0972_));
 sg13g2_buf_2 fanout432 (.A(net434),
    .X(net432));
 sg13g2_buf_1 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(net437),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(net437),
    .X(net435));
 sg13g2_buf_4 fanout436 (.X(net436),
    .A(net437));
 sg13g2_buf_2 fanout437 (.A(rst_n),
    .X(net437));
 sg13g2_buf_1 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[5]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[6]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[2]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[5]),
    .X(net7));
 sg13g2_tielo tt_um_levenshtein_8 (.L_LO(net8));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_leaf_24_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_12_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_22_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_18_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_19_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_20_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\spi.sck_sync[0] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold2 (.A(\spi.mosi_sync[0] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold3 (.A(\spi.ss_n_sync[0] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold4 (.A(\spi.sck ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0029_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0161_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0030_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0153_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold9 (.A(\levenshtein_ctrl.vn[0] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0450_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold11 (.A(\levenshtein_ctrl.symbols[20] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0221_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold13 (.A(\levenshtein_ctrl.symbols[18] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0219_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold15 (.A(\levenshtein_ctrl.symbols[23] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0224_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold17 (.A(\levenshtein_ctrl.symbols[22] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0223_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold19 (.A(\arbiter.wbm_ack_i ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0253_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold21 (.A(\levenshtein_ctrl.symbols[17] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0218_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold23 (.A(\levenshtein_ctrl.vn[1] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0138_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold25 (.A(\levenshtein_ctrl.vn[15] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0152_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold27 (.A(\spi.miso ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold28 (.A(_1087_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0075_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold30 (.A(\levenshtein_ctrl.symbols[21] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0222_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0060_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold33 (.A(_1069_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0068_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold35 (.A(\levenshtein_ctrl.symbols[16] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0217_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0054_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold38 (.A(_1216_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold39 (.A(\spi.counter[1] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold40 (.A(_1071_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0069_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold42 (.A(\levenshtein_ctrl.best_idx[2] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0179_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold44 (.A(\levenshtein_ctrl.best_idx[7] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0184_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold46 (.A(\levenshtein_ctrl.best_idx[6] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0183_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold48 (.A(\levenshtein_ctrl.vn[5] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0142_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold50 (.A(\levenshtein_ctrl.best_idx[4] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0181_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold52 (.A(\levenshtein_ctrl.symbol[3] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0220_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold54 (.A(\levenshtein_ctrl.symbol[0] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0225_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold56 (.A(\levenshtein_ctrl.symbols[10] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold57 (.A(\spi.counter[2] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold58 (.A(_1072_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0070_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold60 (.A(\levenshtein_ctrl.symbol[4] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0229_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold62 (.A(\levenshtein_ctrl.symbol[5] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0230_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold64 (.A(\levenshtein_ctrl.vn[12] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0149_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold66 (.A(\levenshtein_ctrl.pm[15] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold67 (.A(\levenshtein_ctrl.symbols[14] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold68 (.A(\levenshtein_ctrl.vn[14] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold69 (.A(\levenshtein_ctrl.symbol[7] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0232_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold71 (.A(\levenshtein_ctrl.vn[2] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0139_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold73 (.A(\levenshtein_ctrl.symbols[8] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0201_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold75 (.A(\levenshtein_ctrl.symbols[11] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0204_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0041_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold78 (.A(_1248_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0107_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold80 (.A(\spi.counter[3] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold81 (.A(\levenshtein_ctrl.symbols[9] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold82 (.A(\levenshtein_ctrl.vn[6] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold83 (.A(\levenshtein_ctrl.next_symbol[1] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold84 (.A(\levenshtein_ctrl.symbols[12] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0052_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold86 (.A(_1221_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0095_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold88 (.A(\levenshtein_ctrl.next_symbol[4] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold89 (.A(\levenshtein_ctrl.symbols[13] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold90 (.A(\levenshtein_ctrl.pm[14] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0045_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold92 (.A(_1239_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0103_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold94 (.A(\levenshtein_ctrl.best_idx[0] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0177_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold96 (.A(\levenshtein_ctrl.dict_address[8] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0100_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0063_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0121_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold100 (.A(\levenshtein_ctrl.symbols[15] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold101 (.A(\levenshtein_ctrl.best_idx[13] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0190_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold103 (.A(\levenshtein_ctrl.best_idx[15] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0192_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold105 (.A(\levenshtein_ctrl.best_idx[5] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0182_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold107 (.A(\levenshtein_ctrl.symbols[19] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold108 (.A(\levenshtein_ctrl.symbol[6] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0231_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold110 (.A(\levenshtein_ctrl.next_symbol[6] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold111 (.A(\levenshtein_ctrl.vn[8] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0145_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold113 (.A(\spi.counter[4] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold114 (.A(\levenshtein_ctrl.next_symbol[7] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold115 (.A(\arbiter.wbs0_dat_i[6] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0246_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold117 (.A(\levenshtein_ctrl.next_symbol[2] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold118 (.A(\levenshtein_ctrl.pm[13] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0238_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold120 (.A(\levenshtein_ctrl.next_symbol[5] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold121 (.A(\levenshtein_ctrl.best_idx[14] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0191_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold123 (.A(\levenshtein_ctrl.idx[2] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0163_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0047_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold126 (.A(_1235_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0101_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold128 (.A(\levenshtein_ctrl.idx[15] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0176_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0050_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0097_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold132 (.A(\arbiter.wbs0_adr_i[11] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0276_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold134 (.A(\arbiter.wbs0_adr_i[6] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0271_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold136 (.A(\arbiter.wbs0_dat_i[4] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0244_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold138 (.A(\levenshtein_ctrl.pm[3] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0116_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold140 (.A(\levenshtein_ctrl.dict_address[4] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0096_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold142 (.A(\levenshtein_ctrl.dict_address[1] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold143 (.A(_1217_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0093_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold145 (.A(\levenshtein_ctrl.best_distance[0] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0193_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold147 (.A(\levenshtein_ctrl.pm[1] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold148 (.A(\levenshtein_ctrl.idx[7] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0168_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold150 (.A(\levenshtein_ctrl.idx[4] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0165_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold152 (.A(\levenshtein_ctrl.idx[3] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0619_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold154 (.A(\arbiter.wbs0_adr_i[7] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold155 (.A(\levenshtein_ctrl.best_idx[12] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0189_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold157 (.A(\levenshtein_ctrl.dict_address[2] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0094_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold159 (.A(\levenshtein_ctrl.idx[10] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0171_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold161 (.A(\arbiter.wbs0_dat_i[7] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold162 (.A(\levenshtein_ctrl.best_idx[1] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0178_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold164 (.A(\arbiter.wbs0_dat_i[5] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0039_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold166 (.A(_1252_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0109_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold168 (.A(\levenshtein_ctrl.best_distance[5] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0198_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0058_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold171 (.A(\levenshtein_ctrl.best_distance[6] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0199_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0043_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold174 (.A(_1243_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0105_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0037_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold177 (.A(_1256_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0111_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold179 (.A(\levenshtein_ctrl.pm[9] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0234_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold181 (.A(\levenshtein_ctrl.vn[11] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0466_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold183 (.A(\levenshtein_ctrl.dict_address[20] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0112_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold185 (.A(\levenshtein_ctrl.idx[6] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0625_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0167_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold188 (.A(uio_oe[2]),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold189 (.A(\levenshtein_ctrl.symbol[1] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold190 (.A(\levenshtein_ctrl.best_idx[3] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold191 (.A(\arbiter.wbs0_adr_i[5] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0270_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold193 (.A(\levenshtein_ctrl.dict_address[18] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0110_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold195 (.A(\levenshtein_ctrl.vn[10] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0147_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold197 (.A(\arbiter.wbs0_adr_i[8] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold198 (.A(\levenshtein_ctrl.best_distance[7] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0200_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold200 (.A(\levenshtein_ctrl.state[1] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold201 (.A(_1025_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0003_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold203 (.A(\levenshtein_ctrl.idx[8] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0631_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0170_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold206 (.A(\levenshtein_ctrl.d[7] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0160_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold208 (.A(\levenshtein_ctrl.best_distance[4] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0197_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold210 (.A(\levenshtein_ctrl.best_idx[8] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold211 (.A(\levenshtein_ctrl.vn[4] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold212 (.A(\levenshtein_ctrl.symbol[2] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold213 (.A(\levenshtein_ctrl.dict_address[6] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0098_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold215 (.A(\levenshtein_ctrl.pm[11] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0735_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0236_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold218 (.A(\arbiter.wbs0_adr_i[2] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0267_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold220 (.A(\levenshtein_ctrl.idx[1] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0615_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0162_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold223 (.A(\levenshtein_ctrl.dict_address[16] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0108_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold225 (.A(\levenshtein_ctrl.idx[5] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold226 (.A(uio_oe[1]),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0795_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold228 (.A(\arbiter.wbs0_adr_i[4] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0269_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold230 (.A(\levenshtein_ctrl.idx[13] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0174_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold232 (.A(\arbiter.wbs0_adr_i[17] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0282_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold234 (.A(\arbiter.wbs0_adr_i[16] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0281_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0020_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0905_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold238 (.A(\levenshtein_ctrl.dict_address[14] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0106_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold240 (.A(\arbiter.wbs0_adr_i[22] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0914_),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0288_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold243 (.A(uio_oe[5]),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold244 (.A(\levenshtein_ctrl.vn[13] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold245 (.A(\levenshtein_ctrl.pm[5] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0118_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold247 (.A(\levenshtein_ctrl.symbol_idx[1] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0074_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold249 (.A(\levenshtein_ctrl.sram_config[1] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0084_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0048_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold252 (.A(_1231_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0099_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold254 (.A(\levenshtein_ctrl.dict_address[10] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0102_),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold256 (.A(\arbiter.wbs0_adr_i[18] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold257 (.A(uio_oe[4]),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold258 (.A(\arbiter.wbs0_dat_i[2] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0242_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold260 (.A(\levenshtein_ctrl.pm[12] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0237_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold262 (.A(\arbiter.wbs0_adr_i[15] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0280_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold264 (.A(\spi_ctrl.bit_counter[4] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0290_),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold266 (.A(\arbiter.wbs0_adr_i[9] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0275_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold268 (.A(\levenshtein_ctrl.d[5] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold269 (.A(\arbiter.wbs0_adr_i[14] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0279_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0011_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0076_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold273 (.A(\levenshtein_ctrl.pm[7] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold274 (.A(\levenshtein_ctrl.best_idx[10] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold275 (.A(\levenshtein_ctrl.pm[2] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold276 (.A(\levenshtein_ctrl.pm[0] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold277 (.A(\levenshtein_ctrl.d[6] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0159_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold279 (.A(\levenshtein_ctrl.word_length_reg[2] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold280 (.A(\arbiter.wbs0_dat_i[3] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0091_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold282 (.A(\arbiter.wbs0_adr_i[3] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0268_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold284 (.A(\levenshtein_ctrl.vn[9] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold285 (.A(\arbiter.wbs0_adr_i[12] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold286 (.A(\levenshtein_ctrl.dict_address[12] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0104_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold288 (.A(\levenshtein_ctrl.pm[10] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold289 (.A(\arbiter.wbs0_adr_i[13] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0067_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold291 (.A(\arbiter.wbm_dat_i[3] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold292 (.A(\arbiter.wbs0_dat_i[1] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0241_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold294 (.A(\spi.mosi ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0928_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0292_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold297 (.A(\levenshtein_ctrl.state[4] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold298 (.A(_1049_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold299 (.A(\levenshtein_ctrl.idx[12] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0637_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold301 (.A(\spi.state[2] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0009_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold303 (.A(\levenshtein_ctrl.word_length_reg[1] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold304 (.A(\levenshtein_ctrl.state[6] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold305 (.A(_1047_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold306 (.A(\levenshtein_ctrl.vn[3] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold307 (.A(\arbiter.wbs0_adr_i[19] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold308 (.A(\arbiter.wbs0_adr_i[0] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold309 (.A(\levenshtein_ctrl.pm[8] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold310 (.A(\levenshtein_ctrl.pm[6] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold311 (.A(\arbiter.wbs0_adr_i[21] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0286_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold313 (.A(\levenshtein_ctrl.state[2] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold314 (.A(\levenshtein_ctrl.idx[11] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0635_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold316 (.A(\levenshtein_ctrl.sram_config[0] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0083_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold318 (.A(\levenshtein_ctrl.state[5] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold319 (.A(_1030_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0001_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold321 (.A(\levenshtein_ctrl.next_symbol[3] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold322 (.A(\levenshtein_ctrl.best_distance[1] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold323 (.A(\arbiter.wbm_dat_i[7] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold324 (.A(\spi.state[0] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0057_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0085_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold327 (.A(\arbiter.wbs0_adr_i[20] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold328 (.A(\levenshtein_ctrl.vn[7] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold329 (.A(\levenshtein_ctrl.best_idx[9] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0186_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold331 (.A(\levenshtein_ctrl.best_distance[2] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0195_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold333 (.A(\levenshtein_ctrl.state[7] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0059_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold335 (.A(_1079_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold336 (.A(_1080_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold337 (.A(\levenshtein_ctrl.idx[14] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold338 (.A(\spi_ctrl.sck ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold339 (.A(\levenshtein_ctrl.best_distance[3] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0196_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0056_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0000_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold343 (.A(\levenshtein_ctrl.vp[6] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold344 (.A(\levenshtein_ctrl.best_idx[11] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold345 (.A(\levenshtein_ctrl.state[3] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold346 (.A(_1068_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold347 (.A(\levenshtein_ctrl.pm[4] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold348 (.A(\arbiter.cyc ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold349 (.A(_1202_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0082_),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold351 (.A(\arbiter.wbs0_adr_i[1] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold352 (.A(uio_out[5]),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold353 (.A(\levenshtein_ctrl.vp[10] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0131_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold355 (.A(\arbiter.wbs0_dat_i[0] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0088_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0065_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold358 (.A(\levenshtein_ctrl.vp[5] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold359 (.A(\spi_ctrl.ss_n ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold360 (.A(_1133_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold361 (.A(uio_out[4]),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold362 (.A(uio_out[2]),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold363 (.A(ctrl_slave_ack),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold364 (.A(\levenshtein_ctrl.vp[2] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold365 (.A(\levenshtein_ctrl.vp[7] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold366 (.A(\spi_ctrl.bit_counter[3] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold367 (.A(\levenshtein_ctrl.vp[11] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0132_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold369 (.A(\levenshtein_ctrl.vp[8] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0129_),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold371 (.A(\levenshtein_ctrl.vp[14] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold372 (.A(\levenshtein_ctrl.vp[12] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0418_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0134_),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold375 (.A(\levenshtein_ctrl.vp[3] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold376 (.A(\levenshtein_ctrl.vp[15] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold377 (.A(\levenshtein_ctrl.vp[1] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold378 (.A(\levenshtein_ctrl.d[4] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold379 (.A(uio_out[1]),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold380 (.A(\levenshtein_ctrl.vp[4] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0125_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold382 (.A(\levenshtein_ctrl.d[2] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold383 (.A(\spi_ctrl.bit_counter[1] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold384 (.A(\arbiter.wbm_dat_i[5] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0263_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold386 (.A(\arbiter.wbm_dat_i[1] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold387 (.A(\levenshtein_ctrl.vn[3] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold388 (.A(\levenshtein_ctrl.vp[8] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0363_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold390 (.A(\levenshtein_ctrl.pm[11] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold391 (.A(\arbiter.wbm_dat_i[1] ),
    .X(net761));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_fill_2 FILLER_7_182 ();
 sg13g2_fill_1 FILLER_7_184 ();
 sg13g2_decap_4 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_197 ();
 sg13g2_decap_4 FILLER_7_204 ();
 sg13g2_decap_4 FILLER_7_212 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_fill_2 FILLER_8_183 ();
 sg13g2_fill_1 FILLER_8_185 ();
 sg13g2_fill_2 FILLER_8_195 ();
 sg13g2_fill_1 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_163 ();
 sg13g2_decap_8 FILLER_9_244 ();
 sg13g2_decap_8 FILLER_9_251 ();
 sg13g2_decap_8 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_265 ();
 sg13g2_decap_8 FILLER_9_272 ();
 sg13g2_decap_8 FILLER_9_279 ();
 sg13g2_decap_8 FILLER_9_286 ();
 sg13g2_decap_8 FILLER_9_293 ();
 sg13g2_decap_8 FILLER_9_300 ();
 sg13g2_decap_8 FILLER_9_307 ();
 sg13g2_decap_8 FILLER_9_314 ();
 sg13g2_decap_8 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_156 ();
 sg13g2_decap_8 FILLER_10_258 ();
 sg13g2_decap_8 FILLER_10_265 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_decap_8 FILLER_10_279 ();
 sg13g2_decap_8 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_293 ();
 sg13g2_decap_8 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_decap_8 FILLER_10_314 ();
 sg13g2_decap_8 FILLER_10_321 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_261 ();
 sg13g2_decap_8 FILLER_11_268 ();
 sg13g2_decap_8 FILLER_11_275 ();
 sg13g2_decap_8 FILLER_11_282 ();
 sg13g2_decap_8 FILLER_11_289 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_fill_2 FILLER_12_168 ();
 sg13g2_fill_2 FILLER_12_220 ();
 sg13g2_fill_1 FILLER_12_222 ();
 sg13g2_decap_8 FILLER_12_272 ();
 sg13g2_decap_8 FILLER_12_279 ();
 sg13g2_decap_8 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_293 ();
 sg13g2_decap_8 FILLER_12_300 ();
 sg13g2_decap_8 FILLER_12_307 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_4 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_193 ();
 sg13g2_fill_2 FILLER_13_201 ();
 sg13g2_decap_8 FILLER_13_272 ();
 sg13g2_decap_8 FILLER_13_279 ();
 sg13g2_decap_8 FILLER_13_286 ();
 sg13g2_decap_8 FILLER_13_293 ();
 sg13g2_decap_8 FILLER_13_300 ();
 sg13g2_decap_8 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_314 ();
 sg13g2_decap_8 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_328 ();
 sg13g2_decap_8 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_139 ();
 sg13g2_fill_2 FILLER_14_146 ();
 sg13g2_fill_1 FILLER_14_148 ();
 sg13g2_decap_8 FILLER_14_153 ();
 sg13g2_decap_8 FILLER_14_160 ();
 sg13g2_fill_2 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_276 ();
 sg13g2_decap_8 FILLER_14_283 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_decap_8 FILLER_14_297 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_318 ();
 sg13g2_decap_8 FILLER_14_325 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_374 ();
 sg13g2_decap_8 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_14_388 ();
 sg13g2_decap_8 FILLER_14_395 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_4 FILLER_15_119 ();
 sg13g2_fill_2 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_2 FILLER_15_193 ();
 sg13g2_fill_1 FILLER_15_210 ();
 sg13g2_fill_2 FILLER_15_258 ();
 sg13g2_fill_1 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_278 ();
 sg13g2_decap_8 FILLER_15_285 ();
 sg13g2_decap_8 FILLER_15_292 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_fill_2 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_121 ();
 sg13g2_fill_2 FILLER_16_183 ();
 sg13g2_fill_1 FILLER_16_185 ();
 sg13g2_fill_2 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_224 ();
 sg13g2_fill_2 FILLER_16_240 ();
 sg13g2_fill_1 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_4 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_123 ();
 sg13g2_fill_2 FILLER_17_157 ();
 sg13g2_fill_2 FILLER_17_202 ();
 sg13g2_fill_2 FILLER_17_235 ();
 sg13g2_decap_8 FILLER_17_271 ();
 sg13g2_decap_8 FILLER_17_278 ();
 sg13g2_decap_8 FILLER_17_285 ();
 sg13g2_decap_8 FILLER_17_292 ();
 sg13g2_decap_8 FILLER_17_299 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_decap_8 FILLER_17_313 ();
 sg13g2_decap_8 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_327 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_4 FILLER_18_119 ();
 sg13g2_fill_2 FILLER_18_123 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_decap_8 FILLER_18_163 ();
 sg13g2_decap_4 FILLER_18_170 ();
 sg13g2_fill_1 FILLER_18_174 ();
 sg13g2_fill_2 FILLER_18_206 ();
 sg13g2_fill_2 FILLER_18_234 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_fill_1 FILLER_18_255 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_166 ();
 sg13g2_fill_2 FILLER_19_170 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_decap_4 FILLER_19_295 ();
 sg13g2_fill_1 FILLER_19_299 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_4 FILLER_20_105 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_237 ();
 sg13g2_fill_1 FILLER_20_261 ();
 sg13g2_fill_2 FILLER_20_281 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_93 ();
 sg13g2_fill_1 FILLER_21_144 ();
 sg13g2_fill_2 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_84 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_fill_2 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_fill_2 FILLER_22_328 ();
 sg13g2_fill_2 FILLER_22_335 ();
 sg13g2_fill_1 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_132 ();
 sg13g2_fill_1 FILLER_23_161 ();
 sg13g2_fill_1 FILLER_23_184 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_209 ();
 sg13g2_fill_1 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_254 ();
 sg13g2_decap_4 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_123 ();
 sg13g2_decap_4 FILLER_24_211 ();
 sg13g2_fill_1 FILLER_24_215 ();
 sg13g2_fill_2 FILLER_24_220 ();
 sg13g2_fill_2 FILLER_24_231 ();
 sg13g2_fill_1 FILLER_24_233 ();
 sg13g2_fill_2 FILLER_24_242 ();
 sg13g2_fill_1 FILLER_24_280 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_fill_2 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_fill_1 FILLER_25_138 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_230 ();
 sg13g2_decap_4 FILLER_25_246 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_decap_8 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_288 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_4 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_88 ();
 sg13g2_fill_1 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_185 ();
 sg13g2_decap_4 FILLER_26_209 ();
 sg13g2_fill_1 FILLER_26_213 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_fill_2 FILLER_26_282 ();
 sg13g2_decap_8 FILLER_26_293 ();
 sg13g2_decap_4 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_304 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_4 FILLER_26_323 ();
 sg13g2_fill_2 FILLER_26_327 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_4 FILLER_27_81 ();
 sg13g2_fill_1 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_184 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_202 ();
 sg13g2_fill_2 FILLER_27_209 ();
 sg13g2_fill_1 FILLER_27_211 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_fill_2 FILLER_27_289 ();
 sg13g2_fill_1 FILLER_27_305 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_70 ();
 sg13g2_fill_1 FILLER_28_72 ();
 sg13g2_fill_1 FILLER_28_131 ();
 sg13g2_decap_4 FILLER_28_186 ();
 sg13g2_fill_2 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_63 ();
 sg13g2_fill_1 FILLER_29_65 ();
 sg13g2_fill_2 FILLER_29_102 ();
 sg13g2_fill_2 FILLER_29_113 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_decap_4 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_1 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_178 ();
 sg13g2_decap_8 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_263 ();
 sg13g2_fill_2 FILLER_30_300 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_316 ();
 sg13g2_fill_2 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_178 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_196 ();
 sg13g2_fill_2 FILLER_31_214 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_fill_2 FILLER_31_291 ();
 sg13g2_decap_4 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_348 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_363 ();
 sg13g2_fill_1 FILLER_31_365 ();
 sg13g2_fill_1 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_4 FILLER_32_70 ();
 sg13g2_fill_2 FILLER_32_74 ();
 sg13g2_fill_2 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_4 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_fill_1 FILLER_33_114 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_187 ();
 sg13g2_fill_1 FILLER_33_189 ();
 sg13g2_fill_2 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_281 ();
 sg13g2_fill_1 FILLER_33_291 ();
 sg13g2_fill_2 FILLER_33_363 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_67 ();
 sg13g2_fill_2 FILLER_34_95 ();
 sg13g2_fill_1 FILLER_34_97 ();
 sg13g2_fill_2 FILLER_34_138 ();
 sg13g2_decap_4 FILLER_34_186 ();
 sg13g2_decap_4 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_280 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_4 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_67 ();
 sg13g2_fill_1 FILLER_35_130 ();
 sg13g2_fill_2 FILLER_35_175 ();
 sg13g2_fill_1 FILLER_35_177 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_4 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_fill_2 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_395 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_90 ();
 sg13g2_decap_8 FILLER_36_95 ();
 sg13g2_decap_8 FILLER_36_102 ();
 sg13g2_decap_4 FILLER_36_109 ();
 sg13g2_decap_8 FILLER_36_162 ();
 sg13g2_decap_4 FILLER_36_169 ();
 sg13g2_fill_1 FILLER_36_173 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_fill_2 FILLER_36_266 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_356 ();
 sg13g2_decap_8 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_fill_1 FILLER_37_108 ();
 sg13g2_fill_2 FILLER_37_163 ();
 sg13g2_fill_1 FILLER_37_165 ();
 sg13g2_fill_2 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_319 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_fill_2 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_91 ();
 sg13g2_fill_1 FILLER_38_93 ();
 sg13g2_fill_2 FILLER_38_204 ();
 sg13g2_fill_1 FILLER_38_206 ();
 sg13g2_fill_1 FILLER_38_282 ();
 sg13g2_fill_2 FILLER_38_376 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_fill_2 FILLER_39_117 ();
 sg13g2_fill_1 FILLER_39_119 ();
 sg13g2_fill_2 FILLER_39_129 ();
 sg13g2_fill_1 FILLER_39_131 ();
 sg13g2_fill_2 FILLER_39_178 ();
 sg13g2_fill_1 FILLER_39_180 ();
 sg13g2_fill_1 FILLER_39_190 ();
 sg13g2_fill_1 FILLER_39_219 ();
 sg13g2_fill_1 FILLER_39_306 ();
 sg13g2_fill_2 FILLER_39_311 ();
 sg13g2_fill_1 FILLER_39_313 ();
 sg13g2_fill_2 FILLER_39_352 ();
 sg13g2_fill_2 FILLER_39_363 ();
 sg13g2_decap_8 FILLER_39_395 ();
 sg13g2_decap_8 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_4 FILLER_40_77 ();
 sg13g2_fill_1 FILLER_40_81 ();
 sg13g2_fill_2 FILLER_40_112 ();
 sg13g2_fill_1 FILLER_40_114 ();
 sg13g2_fill_2 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_181 ();
 sg13g2_decap_4 FILLER_40_213 ();
 sg13g2_decap_4 FILLER_40_221 ();
 sg13g2_fill_1 FILLER_40_225 ();
 sg13g2_decap_4 FILLER_40_239 ();
 sg13g2_fill_2 FILLER_40_243 ();
 sg13g2_fill_1 FILLER_40_278 ();
 sg13g2_fill_2 FILLER_40_287 ();
 sg13g2_fill_1 FILLER_40_289 ();
 sg13g2_decap_8 FILLER_40_303 ();
 sg13g2_decap_8 FILLER_40_310 ();
 sg13g2_decap_8 FILLER_40_317 ();
 sg13g2_decap_8 FILLER_40_324 ();
 sg13g2_decap_4 FILLER_40_339 ();
 sg13g2_fill_1 FILLER_40_354 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_fill_1 FILLER_41_77 ();
 sg13g2_fill_2 FILLER_41_101 ();
 sg13g2_fill_2 FILLER_41_126 ();
 sg13g2_decap_4 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_214 ();
 sg13g2_decap_8 FILLER_41_221 ();
 sg13g2_fill_1 FILLER_41_228 ();
 sg13g2_fill_2 FILLER_41_234 ();
 sg13g2_fill_1 FILLER_41_236 ();
 sg13g2_decap_8 FILLER_41_248 ();
 sg13g2_fill_1 FILLER_41_255 ();
 sg13g2_decap_8 FILLER_41_260 ();
 sg13g2_fill_2 FILLER_41_283 ();
 sg13g2_decap_8 FILLER_41_290 ();
 sg13g2_decap_8 FILLER_41_297 ();
 sg13g2_decap_8 FILLER_41_304 ();
 sg13g2_decap_8 FILLER_41_311 ();
 sg13g2_decap_4 FILLER_41_318 ();
 sg13g2_fill_1 FILLER_41_331 ();
 sg13g2_fill_1 FILLER_41_362 ();
 sg13g2_fill_1 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_fill_2 FILLER_42_70 ();
 sg13g2_fill_1 FILLER_42_72 ();
 sg13g2_fill_2 FILLER_42_94 ();
 sg13g2_fill_2 FILLER_42_104 ();
 sg13g2_fill_1 FILLER_42_106 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_fill_1 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_166 ();
 sg13g2_fill_1 FILLER_42_173 ();
 sg13g2_fill_1 FILLER_42_249 ();
 sg13g2_decap_4 FILLER_42_259 ();
 sg13g2_decap_4 FILLER_42_267 ();
 sg13g2_fill_1 FILLER_42_271 ();
 sg13g2_decap_8 FILLER_42_277 ();
 sg13g2_decap_8 FILLER_42_284 ();
 sg13g2_decap_4 FILLER_42_291 ();
 sg13g2_fill_1 FILLER_42_295 ();
 sg13g2_fill_2 FILLER_42_312 ();
 sg13g2_fill_2 FILLER_42_367 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_fill_2 FILLER_43_103 ();
 sg13g2_fill_1 FILLER_43_105 ();
 sg13g2_fill_1 FILLER_43_155 ();
 sg13g2_fill_2 FILLER_43_159 ();
 sg13g2_fill_1 FILLER_43_161 ();
 sg13g2_fill_1 FILLER_43_166 ();
 sg13g2_decap_4 FILLER_43_171 ();
 sg13g2_fill_2 FILLER_43_175 ();
 sg13g2_fill_1 FILLER_43_182 ();
 sg13g2_decap_4 FILLER_43_235 ();
 sg13g2_fill_1 FILLER_43_239 ();
 sg13g2_fill_2 FILLER_43_248 ();
 sg13g2_decap_4 FILLER_43_255 ();
 sg13g2_fill_2 FILLER_43_271 ();
 sg13g2_fill_1 FILLER_43_273 ();
 sg13g2_fill_2 FILLER_43_289 ();
 sg13g2_fill_1 FILLER_43_321 ();
 sg13g2_fill_2 FILLER_43_365 ();
 sg13g2_decap_4 FILLER_43_386 ();
 sg13g2_fill_2 FILLER_43_390 ();
 sg13g2_decap_4 FILLER_43_405 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_4 FILLER_44_70 ();
 sg13g2_fill_2 FILLER_44_74 ();
 sg13g2_fill_2 FILLER_44_141 ();
 sg13g2_fill_1 FILLER_44_143 ();
 sg13g2_fill_2 FILLER_44_149 ();
 sg13g2_fill_2 FILLER_44_177 ();
 sg13g2_fill_1 FILLER_44_179 ();
 sg13g2_fill_2 FILLER_44_193 ();
 sg13g2_fill_1 FILLER_44_195 ();
 sg13g2_fill_2 FILLER_44_206 ();
 sg13g2_fill_1 FILLER_44_213 ();
 sg13g2_fill_1 FILLER_44_222 ();
 sg13g2_fill_2 FILLER_44_237 ();
 sg13g2_decap_8 FILLER_44_243 ();
 sg13g2_fill_1 FILLER_44_250 ();
 sg13g2_fill_2 FILLER_44_255 ();
 sg13g2_fill_2 FILLER_44_292 ();
 sg13g2_decap_8 FILLER_44_339 ();
 sg13g2_decap_4 FILLER_44_346 ();
 sg13g2_fill_2 FILLER_44_362 ();
 sg13g2_fill_1 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_fill_1 FILLER_45_77 ();
 sg13g2_fill_1 FILLER_45_93 ();
 sg13g2_fill_2 FILLER_45_137 ();
 sg13g2_fill_2 FILLER_45_144 ();
 sg13g2_decap_4 FILLER_45_191 ();
 sg13g2_decap_4 FILLER_45_215 ();
 sg13g2_fill_2 FILLER_45_219 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_fill_2 FILLER_45_342 ();
 sg13g2_fill_2 FILLER_45_363 ();
 sg13g2_decap_8 FILLER_45_401 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_4 FILLER_46_63 ();
 sg13g2_fill_1 FILLER_46_140 ();
 sg13g2_fill_1 FILLER_46_146 ();
 sg13g2_fill_2 FILLER_46_191 ();
 sg13g2_fill_1 FILLER_46_219 ();
 sg13g2_fill_2 FILLER_46_268 ();
 sg13g2_fill_1 FILLER_46_270 ();
 sg13g2_fill_1 FILLER_46_343 ();
 sg13g2_fill_1 FILLER_46_350 ();
 sg13g2_fill_2 FILLER_46_377 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_4 FILLER_47_56 ();
 sg13g2_fill_2 FILLER_47_60 ();
 sg13g2_fill_1 FILLER_47_66 ();
 sg13g2_fill_1 FILLER_47_135 ();
 sg13g2_fill_1 FILLER_47_173 ();
 sg13g2_fill_1 FILLER_47_201 ();
 sg13g2_fill_1 FILLER_47_213 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_fill_2 FILLER_47_263 ();
 sg13g2_fill_1 FILLER_47_265 ();
 sg13g2_fill_1 FILLER_47_275 ();
 sg13g2_fill_1 FILLER_47_302 ();
 sg13g2_fill_2 FILLER_47_336 ();
 sg13g2_fill_1 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_402 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_fill_1 FILLER_48_56 ();
 sg13g2_fill_2 FILLER_48_110 ();
 sg13g2_fill_1 FILLER_48_112 ();
 sg13g2_fill_1 FILLER_48_138 ();
 sg13g2_fill_1 FILLER_48_214 ();
 sg13g2_fill_2 FILLER_48_228 ();
 sg13g2_fill_1 FILLER_48_230 ();
 sg13g2_fill_2 FILLER_48_319 ();
 sg13g2_fill_1 FILLER_48_321 ();
 sg13g2_fill_1 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_4 FILLER_49_49 ();
 sg13g2_fill_2 FILLER_49_53 ();
 sg13g2_fill_2 FILLER_49_90 ();
 sg13g2_fill_1 FILLER_49_92 ();
 sg13g2_fill_1 FILLER_49_118 ();
 sg13g2_fill_1 FILLER_49_128 ();
 sg13g2_fill_1 FILLER_49_133 ();
 sg13g2_fill_2 FILLER_49_139 ();
 sg13g2_fill_1 FILLER_49_141 ();
 sg13g2_fill_1 FILLER_49_181 ();
 sg13g2_fill_2 FILLER_49_191 ();
 sg13g2_fill_1 FILLER_49_193 ();
 sg13g2_fill_1 FILLER_49_198 ();
 sg13g2_fill_1 FILLER_49_204 ();
 sg13g2_fill_1 FILLER_49_216 ();
 sg13g2_fill_2 FILLER_49_241 ();
 sg13g2_fill_1 FILLER_49_243 ();
 sg13g2_fill_1 FILLER_49_250 ();
 sg13g2_decap_4 FILLER_49_287 ();
 sg13g2_fill_2 FILLER_49_326 ();
 sg13g2_fill_2 FILLER_49_358 ();
 sg13g2_fill_2 FILLER_49_391 ();
 sg13g2_fill_1 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_398 ();
 sg13g2_decap_4 FILLER_49_405 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_4 FILLER_50_42 ();
 sg13g2_fill_1 FILLER_50_46 ();
 sg13g2_fill_1 FILLER_50_86 ();
 sg13g2_fill_1 FILLER_50_115 ();
 sg13g2_fill_1 FILLER_50_125 ();
 sg13g2_decap_8 FILLER_50_135 ();
 sg13g2_decap_8 FILLER_50_142 ();
 sg13g2_fill_2 FILLER_50_184 ();
 sg13g2_fill_1 FILLER_50_186 ();
 sg13g2_decap_8 FILLER_50_195 ();
 sg13g2_fill_2 FILLER_50_202 ();
 sg13g2_fill_1 FILLER_50_204 ();
 sg13g2_decap_8 FILLER_50_209 ();
 sg13g2_fill_2 FILLER_50_216 ();
 sg13g2_fill_1 FILLER_50_218 ();
 sg13g2_fill_1 FILLER_50_240 ();
 sg13g2_fill_1 FILLER_50_251 ();
 sg13g2_fill_2 FILLER_50_260 ();
 sg13g2_decap_8 FILLER_50_277 ();
 sg13g2_decap_4 FILLER_50_284 ();
 sg13g2_decap_8 FILLER_50_293 ();
 sg13g2_decap_8 FILLER_50_300 ();
 sg13g2_fill_2 FILLER_50_307 ();
 sg13g2_fill_1 FILLER_50_309 ();
 sg13g2_fill_2 FILLER_50_322 ();
 sg13g2_fill_2 FILLER_50_338 ();
 sg13g2_decap_4 FILLER_50_362 ();
 sg13g2_fill_2 FILLER_50_371 ();
 sg13g2_decap_8 FILLER_50_386 ();
 sg13g2_decap_8 FILLER_50_393 ();
 sg13g2_decap_8 FILLER_50_400 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_4 FILLER_51_35 ();
 sg13g2_fill_1 FILLER_51_39 ();
 sg13g2_fill_2 FILLER_51_83 ();
 sg13g2_fill_1 FILLER_51_85 ();
 sg13g2_fill_2 FILLER_51_110 ();
 sg13g2_fill_1 FILLER_51_112 ();
 sg13g2_fill_2 FILLER_51_128 ();
 sg13g2_fill_1 FILLER_51_155 ();
 sg13g2_decap_8 FILLER_51_183 ();
 sg13g2_decap_4 FILLER_51_190 ();
 sg13g2_fill_1 FILLER_51_194 ();
 sg13g2_fill_2 FILLER_51_256 ();
 sg13g2_fill_1 FILLER_51_258 ();
 sg13g2_fill_2 FILLER_51_303 ();
 sg13g2_fill_1 FILLER_51_305 ();
 sg13g2_decap_8 FILLER_51_321 ();
 sg13g2_fill_1 FILLER_51_328 ();
 sg13g2_fill_1 FILLER_51_341 ();
 sg13g2_fill_1 FILLER_51_345 ();
 sg13g2_fill_1 FILLER_51_351 ();
 sg13g2_fill_1 FILLER_51_371 ();
 sg13g2_fill_1 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_fill_1 FILLER_52_42 ();
 sg13g2_fill_1 FILLER_52_79 ();
 sg13g2_fill_1 FILLER_52_123 ();
 sg13g2_fill_2 FILLER_52_134 ();
 sg13g2_fill_1 FILLER_52_145 ();
 sg13g2_fill_1 FILLER_52_161 ();
 sg13g2_decap_4 FILLER_52_168 ();
 sg13g2_fill_2 FILLER_52_172 ();
 sg13g2_fill_1 FILLER_52_179 ();
 sg13g2_fill_2 FILLER_52_197 ();
 sg13g2_fill_2 FILLER_52_244 ();
 sg13g2_fill_2 FILLER_52_256 ();
 sg13g2_fill_1 FILLER_52_270 ();
 sg13g2_fill_2 FILLER_52_283 ();
 sg13g2_fill_1 FILLER_52_285 ();
 sg13g2_decap_4 FILLER_52_290 ();
 sg13g2_fill_1 FILLER_52_294 ();
 sg13g2_fill_2 FILLER_52_314 ();
 sg13g2_fill_2 FILLER_52_322 ();
 sg13g2_fill_1 FILLER_52_324 ();
 sg13g2_decap_4 FILLER_52_330 ();
 sg13g2_fill_1 FILLER_52_347 ();
 sg13g2_fill_1 FILLER_52_381 ();
 sg13g2_fill_1 FILLER_52_391 ();
 sg13g2_decap_4 FILLER_52_405 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_fill_2 FILLER_53_42 ();
 sg13g2_fill_1 FILLER_53_44 ();
 sg13g2_fill_2 FILLER_53_66 ();
 sg13g2_fill_1 FILLER_53_111 ();
 sg13g2_fill_1 FILLER_53_146 ();
 sg13g2_fill_2 FILLER_53_206 ();
 sg13g2_fill_1 FILLER_53_208 ();
 sg13g2_fill_2 FILLER_53_249 ();
 sg13g2_fill_1 FILLER_53_251 ();
 sg13g2_fill_1 FILLER_53_262 ();
 sg13g2_fill_1 FILLER_53_306 ();
 sg13g2_fill_2 FILLER_53_325 ();
 sg13g2_fill_1 FILLER_53_327 ();
 sg13g2_decap_4 FILLER_53_359 ();
 sg13g2_decap_8 FILLER_53_396 ();
 sg13g2_decap_4 FILLER_53_403 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_4 FILLER_54_42 ();
 sg13g2_fill_2 FILLER_54_67 ();
 sg13g2_fill_2 FILLER_54_105 ();
 sg13g2_fill_1 FILLER_54_120 ();
 sg13g2_fill_2 FILLER_54_135 ();
 sg13g2_fill_2 FILLER_54_142 ();
 sg13g2_fill_1 FILLER_54_144 ();
 sg13g2_fill_1 FILLER_54_159 ();
 sg13g2_fill_1 FILLER_54_187 ();
 sg13g2_fill_2 FILLER_54_197 ();
 sg13g2_fill_1 FILLER_54_199 ();
 sg13g2_fill_2 FILLER_54_229 ();
 sg13g2_fill_1 FILLER_54_231 ();
 sg13g2_decap_8 FILLER_54_235 ();
 sg13g2_fill_2 FILLER_54_242 ();
 sg13g2_fill_1 FILLER_54_244 ();
 sg13g2_fill_2 FILLER_54_280 ();
 sg13g2_fill_2 FILLER_54_321 ();
 sg13g2_fill_2 FILLER_54_329 ();
 sg13g2_fill_2 FILLER_54_366 ();
 sg13g2_fill_1 FILLER_54_368 ();
 sg13g2_decap_8 FILLER_54_395 ();
 sg13g2_decap_8 FILLER_54_402 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_fill_2 FILLER_55_42 ();
 sg13g2_fill_2 FILLER_55_88 ();
 sg13g2_fill_1 FILLER_55_90 ();
 sg13g2_decap_8 FILLER_55_100 ();
 sg13g2_decap_8 FILLER_55_107 ();
 sg13g2_fill_2 FILLER_55_124 ();
 sg13g2_decap_4 FILLER_55_155 ();
 sg13g2_fill_2 FILLER_55_159 ();
 sg13g2_fill_2 FILLER_55_187 ();
 sg13g2_fill_2 FILLER_55_205 ();
 sg13g2_decap_8 FILLER_55_215 ();
 sg13g2_decap_8 FILLER_55_222 ();
 sg13g2_fill_2 FILLER_55_229 ();
 sg13g2_fill_1 FILLER_55_231 ();
 sg13g2_fill_1 FILLER_55_262 ();
 sg13g2_fill_2 FILLER_55_354 ();
 sg13g2_fill_2 FILLER_55_361 ();
 sg13g2_fill_2 FILLER_55_377 ();
 sg13g2_fill_1 FILLER_55_379 ();
 sg13g2_decap_8 FILLER_55_397 ();
 sg13g2_decap_4 FILLER_55_404 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_fill_2 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_37 ();
 sg13g2_decap_8 FILLER_56_95 ();
 sg13g2_decap_8 FILLER_56_102 ();
 sg13g2_decap_8 FILLER_56_109 ();
 sg13g2_decap_8 FILLER_56_116 ();
 sg13g2_decap_8 FILLER_56_123 ();
 sg13g2_fill_2 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_132 ();
 sg13g2_fill_2 FILLER_56_137 ();
 sg13g2_fill_1 FILLER_56_139 ();
 sg13g2_decap_8 FILLER_56_150 ();
 sg13g2_fill_1 FILLER_56_160 ();
 sg13g2_fill_1 FILLER_56_170 ();
 sg13g2_decap_4 FILLER_56_223 ();
 sg13g2_fill_2 FILLER_56_253 ();
 sg13g2_decap_4 FILLER_56_300 ();
 sg13g2_fill_2 FILLER_56_304 ();
 sg13g2_fill_1 FILLER_56_315 ();
 sg13g2_fill_1 FILLER_56_326 ();
 sg13g2_fill_2 FILLER_56_342 ();
 sg13g2_fill_2 FILLER_56_351 ();
 sg13g2_decap_8 FILLER_56_358 ();
 sg13g2_decap_8 FILLER_56_370 ();
 sg13g2_decap_8 FILLER_56_377 ();
 sg13g2_decap_8 FILLER_56_384 ();
 sg13g2_decap_8 FILLER_56_391 ();
 sg13g2_decap_8 FILLER_56_398 ();
 sg13g2_decap_4 FILLER_56_405 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_fill_2 FILLER_57_35 ();
 sg13g2_fill_1 FILLER_57_37 ();
 sg13g2_fill_2 FILLER_57_69 ();
 sg13g2_fill_1 FILLER_57_106 ();
 sg13g2_fill_2 FILLER_57_144 ();
 sg13g2_fill_2 FILLER_57_151 ();
 sg13g2_fill_2 FILLER_57_169 ();
 sg13g2_fill_1 FILLER_57_171 ();
 sg13g2_fill_1 FILLER_57_186 ();
 sg13g2_fill_1 FILLER_57_200 ();
 sg13g2_decap_8 FILLER_57_285 ();
 sg13g2_fill_1 FILLER_57_292 ();
 sg13g2_decap_4 FILLER_57_298 ();
 sg13g2_decap_4 FILLER_57_307 ();
 sg13g2_fill_1 FILLER_57_311 ();
 sg13g2_fill_2 FILLER_57_316 ();
 sg13g2_fill_1 FILLER_57_318 ();
 sg13g2_fill_2 FILLER_57_333 ();
 sg13g2_fill_1 FILLER_57_335 ();
 sg13g2_fill_2 FILLER_57_360 ();
 sg13g2_fill_2 FILLER_57_376 ();
 sg13g2_decap_8 FILLER_57_391 ();
 sg13g2_decap_8 FILLER_57_398 ();
 sg13g2_decap_4 FILLER_57_405 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_fill_2 FILLER_58_42 ();
 sg13g2_fill_1 FILLER_58_44 ();
 sg13g2_fill_2 FILLER_58_130 ();
 sg13g2_fill_2 FILLER_58_152 ();
 sg13g2_fill_1 FILLER_58_154 ();
 sg13g2_fill_2 FILLER_58_169 ();
 sg13g2_fill_1 FILLER_58_171 ();
 sg13g2_decap_4 FILLER_58_180 ();
 sg13g2_fill_1 FILLER_58_207 ();
 sg13g2_decap_4 FILLER_58_217 ();
 sg13g2_fill_1 FILLER_58_221 ();
 sg13g2_fill_1 FILLER_58_240 ();
 sg13g2_fill_2 FILLER_58_246 ();
 sg13g2_decap_8 FILLER_58_278 ();
 sg13g2_fill_2 FILLER_58_285 ();
 sg13g2_fill_1 FILLER_58_292 ();
 sg13g2_decap_4 FILLER_58_325 ();
 sg13g2_fill_2 FILLER_58_339 ();
 sg13g2_fill_1 FILLER_58_341 ();
 sg13g2_decap_8 FILLER_58_393 ();
 sg13g2_decap_8 FILLER_58_400 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_fill_2 FILLER_59_106 ();
 sg13g2_fill_2 FILLER_59_160 ();
 sg13g2_fill_2 FILLER_59_194 ();
 sg13g2_decap_8 FILLER_59_222 ();
 sg13g2_fill_1 FILLER_59_239 ();
 sg13g2_fill_1 FILLER_59_370 ();
 sg13g2_decap_8 FILLER_59_397 ();
 sg13g2_decap_4 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_fill_1 FILLER_60_49 ();
 sg13g2_fill_1 FILLER_60_76 ();
 sg13g2_fill_1 FILLER_60_118 ();
 sg13g2_fill_1 FILLER_60_147 ();
 sg13g2_fill_1 FILLER_60_205 ();
 sg13g2_fill_1 FILLER_60_237 ();
 sg13g2_decap_4 FILLER_60_273 ();
 sg13g2_fill_2 FILLER_60_281 ();
 sg13g2_fill_1 FILLER_60_330 ();
 sg13g2_fill_2 FILLER_60_342 ();
 sg13g2_fill_1 FILLER_60_344 ();
 sg13g2_fill_1 FILLER_60_350 ();
 sg13g2_fill_2 FILLER_60_371 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_fill_1 FILLER_60_383 ();
 sg13g2_decap_8 FILLER_60_393 ();
 sg13g2_decap_8 FILLER_60_400 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_4 FILLER_61_42 ();
 sg13g2_fill_2 FILLER_61_62 ();
 sg13g2_fill_1 FILLER_61_64 ();
 sg13g2_fill_2 FILLER_61_79 ();
 sg13g2_fill_2 FILLER_61_100 ();
 sg13g2_fill_1 FILLER_61_102 ();
 sg13g2_fill_1 FILLER_61_112 ();
 sg13g2_fill_2 FILLER_61_129 ();
 sg13g2_fill_2 FILLER_61_149 ();
 sg13g2_fill_1 FILLER_61_155 ();
 sg13g2_fill_2 FILLER_61_160 ();
 sg13g2_fill_1 FILLER_61_167 ();
 sg13g2_fill_2 FILLER_61_276 ();
 sg13g2_fill_1 FILLER_61_278 ();
 sg13g2_fill_2 FILLER_61_292 ();
 sg13g2_fill_1 FILLER_61_318 ();
 sg13g2_fill_1 FILLER_61_336 ();
 sg13g2_fill_2 FILLER_61_352 ();
 sg13g2_fill_2 FILLER_61_380 ();
 sg13g2_decap_8 FILLER_61_389 ();
 sg13g2_decap_8 FILLER_61_396 ();
 sg13g2_decap_4 FILLER_61_403 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_4 FILLER_62_42 ();
 sg13g2_fill_2 FILLER_62_46 ();
 sg13g2_fill_2 FILLER_62_74 ();
 sg13g2_fill_2 FILLER_62_86 ();
 sg13g2_fill_1 FILLER_62_88 ();
 sg13g2_fill_2 FILLER_62_98 ();
 sg13g2_fill_2 FILLER_62_104 ();
 sg13g2_fill_2 FILLER_62_128 ();
 sg13g2_fill_1 FILLER_62_130 ();
 sg13g2_fill_2 FILLER_62_135 ();
 sg13g2_fill_1 FILLER_62_137 ();
 sg13g2_decap_8 FILLER_62_159 ();
 sg13g2_decap_8 FILLER_62_166 ();
 sg13g2_decap_8 FILLER_62_173 ();
 sg13g2_fill_2 FILLER_62_180 ();
 sg13g2_fill_2 FILLER_62_203 ();
 sg13g2_fill_2 FILLER_62_244 ();
 sg13g2_fill_1 FILLER_62_246 ();
 sg13g2_fill_2 FILLER_62_338 ();
 sg13g2_fill_1 FILLER_62_340 ();
 sg13g2_fill_2 FILLER_62_353 ();
 sg13g2_fill_2 FILLER_62_361 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_fill_1 FILLER_63_87 ();
 sg13g2_fill_2 FILLER_63_144 ();
 sg13g2_fill_2 FILLER_63_150 ();
 sg13g2_fill_1 FILLER_63_152 ();
 sg13g2_fill_1 FILLER_63_162 ();
 sg13g2_fill_2 FILLER_63_216 ();
 sg13g2_fill_1 FILLER_63_218 ();
 sg13g2_fill_2 FILLER_63_242 ();
 sg13g2_fill_1 FILLER_63_244 ();
 sg13g2_fill_1 FILLER_63_270 ();
 sg13g2_fill_1 FILLER_63_300 ();
 sg13g2_fill_2 FILLER_63_328 ();
 sg13g2_fill_1 FILLER_63_330 ();
 sg13g2_fill_2 FILLER_63_355 ();
 sg13g2_fill_1 FILLER_63_357 ();
 sg13g2_decap_8 FILLER_63_393 ();
 sg13g2_decap_8 FILLER_63_400 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_fill_1 FILLER_64_83 ();
 sg13g2_fill_2 FILLER_64_126 ();
 sg13g2_fill_2 FILLER_64_147 ();
 sg13g2_fill_1 FILLER_64_149 ();
 sg13g2_fill_1 FILLER_64_160 ();
 sg13g2_fill_2 FILLER_64_195 ();
 sg13g2_fill_1 FILLER_64_207 ();
 sg13g2_fill_2 FILLER_64_221 ();
 sg13g2_fill_1 FILLER_64_223 ();
 sg13g2_fill_2 FILLER_64_229 ();
 sg13g2_fill_1 FILLER_64_231 ();
 sg13g2_fill_2 FILLER_64_241 ();
 sg13g2_fill_1 FILLER_64_243 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_decap_4 FILLER_64_273 ();
 sg13g2_fill_1 FILLER_64_322 ();
 sg13g2_fill_1 FILLER_64_332 ();
 sg13g2_fill_2 FILLER_64_368 ();
 sg13g2_fill_1 FILLER_64_370 ();
 sg13g2_decap_8 FILLER_64_401 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_4 FILLER_65_35 ();
 sg13g2_fill_2 FILLER_65_39 ();
 sg13g2_fill_2 FILLER_65_80 ();
 sg13g2_fill_2 FILLER_65_97 ();
 sg13g2_fill_1 FILLER_65_99 ();
 sg13g2_fill_2 FILLER_65_127 ();
 sg13g2_fill_2 FILLER_65_137 ();
 sg13g2_fill_1 FILLER_65_151 ();
 sg13g2_fill_2 FILLER_65_186 ();
 sg13g2_fill_2 FILLER_65_202 ();
 sg13g2_fill_1 FILLER_65_204 ();
 sg13g2_fill_2 FILLER_65_235 ();
 sg13g2_fill_1 FILLER_65_237 ();
 sg13g2_decap_4 FILLER_65_278 ();
 sg13g2_fill_1 FILLER_65_282 ();
 sg13g2_fill_1 FILLER_65_300 ();
 sg13g2_fill_1 FILLER_65_314 ();
 sg13g2_fill_1 FILLER_65_346 ();
 sg13g2_decap_8 FILLER_65_390 ();
 sg13g2_decap_8 FILLER_65_397 ();
 sg13g2_decap_4 FILLER_65_404 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_4 FILLER_66_42 ();
 sg13g2_fill_2 FILLER_66_46 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_fill_1 FILLER_66_178 ();
 sg13g2_fill_1 FILLER_66_189 ();
 sg13g2_decap_4 FILLER_66_195 ();
 sg13g2_fill_1 FILLER_66_199 ();
 sg13g2_fill_1 FILLER_66_204 ();
 sg13g2_fill_2 FILLER_66_209 ();
 sg13g2_decap_8 FILLER_66_284 ();
 sg13g2_fill_2 FILLER_66_291 ();
 sg13g2_decap_8 FILLER_66_381 ();
 sg13g2_decap_8 FILLER_66_388 ();
 sg13g2_decap_8 FILLER_66_395 ();
 sg13g2_decap_8 FILLER_66_402 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_fill_2 FILLER_67_56 ();
 sg13g2_fill_1 FILLER_67_58 ();
 sg13g2_fill_1 FILLER_67_102 ();
 sg13g2_fill_1 FILLER_67_120 ();
 sg13g2_fill_2 FILLER_67_130 ();
 sg13g2_fill_1 FILLER_67_132 ();
 sg13g2_fill_2 FILLER_67_149 ();
 sg13g2_fill_2 FILLER_67_166 ();
 sg13g2_fill_1 FILLER_67_179 ();
 sg13g2_fill_2 FILLER_67_201 ();
 sg13g2_decap_4 FILLER_67_212 ();
 sg13g2_fill_2 FILLER_67_274 ();
 sg13g2_fill_1 FILLER_67_319 ();
 sg13g2_fill_1 FILLER_67_341 ();
 sg13g2_fill_1 FILLER_67_347 ();
 sg13g2_fill_1 FILLER_67_360 ();
 sg13g2_decap_8 FILLER_67_369 ();
 sg13g2_decap_8 FILLER_67_376 ();
 sg13g2_decap_8 FILLER_67_383 ();
 sg13g2_decap_8 FILLER_67_390 ();
 sg13g2_decap_8 FILLER_67_397 ();
 sg13g2_decap_4 FILLER_67_404 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_fill_1 FILLER_68_63 ();
 sg13g2_fill_1 FILLER_68_94 ();
 sg13g2_fill_1 FILLER_68_137 ();
 sg13g2_fill_1 FILLER_68_224 ();
 sg13g2_fill_1 FILLER_68_242 ();
 sg13g2_decap_8 FILLER_68_325 ();
 sg13g2_decap_4 FILLER_68_332 ();
 sg13g2_decap_8 FILLER_68_346 ();
 sg13g2_decap_4 FILLER_68_353 ();
 sg13g2_decap_8 FILLER_68_366 ();
 sg13g2_decap_8 FILLER_68_373 ();
 sg13g2_decap_8 FILLER_68_380 ();
 sg13g2_decap_8 FILLER_68_387 ();
 sg13g2_decap_8 FILLER_68_394 ();
 sg13g2_decap_8 FILLER_68_401 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_fill_2 FILLER_69_70 ();
 sg13g2_fill_2 FILLER_69_134 ();
 sg13g2_fill_1 FILLER_69_176 ();
 sg13g2_fill_2 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_209 ();
 sg13g2_fill_2 FILLER_69_215 ();
 sg13g2_fill_2 FILLER_69_229 ();
 sg13g2_fill_2 FILLER_69_263 ();
 sg13g2_fill_1 FILLER_69_265 ();
 sg13g2_fill_1 FILLER_69_279 ();
 sg13g2_fill_2 FILLER_69_320 ();
 sg13g2_decap_8 FILLER_69_374 ();
 sg13g2_decap_8 FILLER_69_381 ();
 sg13g2_decap_8 FILLER_69_388 ();
 sg13g2_decap_8 FILLER_69_395 ();
 sg13g2_decap_8 FILLER_69_402 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_fill_2 FILLER_70_70 ();
 sg13g2_fill_1 FILLER_70_72 ();
 sg13g2_fill_2 FILLER_70_159 ();
 sg13g2_fill_1 FILLER_70_192 ();
 sg13g2_fill_1 FILLER_70_255 ();
 sg13g2_fill_2 FILLER_70_266 ();
 sg13g2_fill_2 FILLER_70_277 ();
 sg13g2_fill_1 FILLER_70_279 ();
 sg13g2_fill_2 FILLER_70_297 ();
 sg13g2_fill_1 FILLER_70_299 ();
 sg13g2_fill_2 FILLER_70_358 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_decap_8 FILLER_70_371 ();
 sg13g2_decap_8 FILLER_70_378 ();
 sg13g2_decap_8 FILLER_70_385 ();
 sg13g2_decap_8 FILLER_70_392 ();
 sg13g2_decap_8 FILLER_70_399 ();
 sg13g2_fill_2 FILLER_70_406 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_fill_2 FILLER_71_63 ();
 sg13g2_fill_1 FILLER_71_65 ();
 sg13g2_fill_1 FILLER_71_124 ();
 sg13g2_fill_2 FILLER_71_151 ();
 sg13g2_fill_2 FILLER_71_172 ();
 sg13g2_fill_1 FILLER_71_200 ();
 sg13g2_fill_1 FILLER_71_234 ();
 sg13g2_fill_2 FILLER_71_261 ();
 sg13g2_fill_1 FILLER_71_289 ();
 sg13g2_decap_8 FILLER_71_299 ();
 sg13g2_decap_8 FILLER_71_306 ();
 sg13g2_decap_8 FILLER_71_313 ();
 sg13g2_fill_1 FILLER_71_320 ();
 sg13g2_decap_4 FILLER_71_325 ();
 sg13g2_fill_1 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_375 ();
 sg13g2_decap_8 FILLER_71_382 ();
 sg13g2_decap_8 FILLER_71_389 ();
 sg13g2_decap_8 FILLER_71_396 ();
 sg13g2_decap_4 FILLER_71_403 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_fill_2 FILLER_72_102 ();
 sg13g2_fill_1 FILLER_72_104 ();
 sg13g2_fill_2 FILLER_72_115 ();
 sg13g2_fill_1 FILLER_72_117 ();
 sg13g2_decap_4 FILLER_72_131 ();
 sg13g2_fill_1 FILLER_72_143 ();
 sg13g2_fill_2 FILLER_72_188 ();
 sg13g2_fill_2 FILLER_72_230 ();
 sg13g2_fill_2 FILLER_72_250 ();
 sg13g2_fill_1 FILLER_72_312 ();
 sg13g2_fill_2 FILLER_72_322 ();
 sg13g2_fill_1 FILLER_72_324 ();
 sg13g2_decap_8 FILLER_72_370 ();
 sg13g2_decap_8 FILLER_72_377 ();
 sg13g2_decap_8 FILLER_72_384 ();
 sg13g2_decap_8 FILLER_72_391 ();
 sg13g2_decap_8 FILLER_72_398 ();
 sg13g2_decap_4 FILLER_72_405 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_fill_2 FILLER_73_70 ();
 sg13g2_fill_1 FILLER_73_72 ();
 sg13g2_fill_1 FILLER_73_99 ();
 sg13g2_decap_4 FILLER_73_140 ();
 sg13g2_fill_2 FILLER_73_149 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_fill_2 FILLER_73_166 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_fill_2 FILLER_73_182 ();
 sg13g2_fill_1 FILLER_73_184 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_4 FILLER_73_196 ();
 sg13g2_fill_1 FILLER_73_200 ();
 sg13g2_decap_4 FILLER_73_205 ();
 sg13g2_fill_2 FILLER_73_209 ();
 sg13g2_fill_2 FILLER_73_223 ();
 sg13g2_fill_2 FILLER_73_254 ();
 sg13g2_fill_2 FILLER_73_270 ();
 sg13g2_fill_1 FILLER_73_272 ();
 sg13g2_decap_4 FILLER_73_309 ();
 sg13g2_decap_8 FILLER_73_357 ();
 sg13g2_decap_8 FILLER_73_364 ();
 sg13g2_decap_8 FILLER_73_371 ();
 sg13g2_decap_8 FILLER_73_378 ();
 sg13g2_decap_8 FILLER_73_385 ();
 sg13g2_decap_8 FILLER_73_392 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_fill_2 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_fill_2 FILLER_74_70 ();
 sg13g2_fill_2 FILLER_74_160 ();
 sg13g2_decap_4 FILLER_74_176 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_fill_2 FILLER_74_203 ();
 sg13g2_fill_1 FILLER_74_205 ();
 sg13g2_fill_2 FILLER_74_219 ();
 sg13g2_fill_2 FILLER_74_236 ();
 sg13g2_fill_2 FILLER_74_243 ();
 sg13g2_fill_1 FILLER_74_245 ();
 sg13g2_fill_2 FILLER_74_281 ();
 sg13g2_fill_1 FILLER_74_283 ();
 sg13g2_fill_2 FILLER_74_336 ();
 sg13g2_fill_1 FILLER_74_338 ();
 sg13g2_fill_2 FILLER_74_343 ();
 sg13g2_fill_1 FILLER_74_345 ();
 sg13g2_decap_8 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_357 ();
 sg13g2_decap_8 FILLER_74_364 ();
 sg13g2_decap_8 FILLER_74_371 ();
 sg13g2_decap_8 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_fill_1 FILLER_75_77 ();
 sg13g2_decap_4 FILLER_75_104 ();
 sg13g2_fill_2 FILLER_75_134 ();
 sg13g2_fill_2 FILLER_75_140 ();
 sg13g2_fill_2 FILLER_75_172 ();
 sg13g2_fill_2 FILLER_75_180 ();
 sg13g2_fill_1 FILLER_75_282 ();
 sg13g2_fill_1 FILLER_75_296 ();
 sg13g2_decap_8 FILLER_75_337 ();
 sg13g2_decap_8 FILLER_75_344 ();
 sg13g2_decap_8 FILLER_75_351 ();
 sg13g2_decap_8 FILLER_75_358 ();
 sg13g2_decap_8 FILLER_75_365 ();
 sg13g2_decap_8 FILLER_75_372 ();
 sg13g2_decap_8 FILLER_75_379 ();
 sg13g2_decap_8 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_fill_1 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_131 ();
 sg13g2_decap_4 FILLER_76_138 ();
 sg13g2_fill_2 FILLER_76_142 ();
 sg13g2_fill_2 FILLER_76_170 ();
 sg13g2_fill_1 FILLER_76_172 ();
 sg13g2_fill_2 FILLER_76_229 ();
 sg13g2_fill_2 FILLER_76_297 ();
 sg13g2_fill_1 FILLER_76_299 ();
 sg13g2_decap_8 FILLER_76_332 ();
 sg13g2_decap_8 FILLER_76_339 ();
 sg13g2_decap_8 FILLER_76_346 ();
 sg13g2_decap_8 FILLER_76_353 ();
 sg13g2_decap_8 FILLER_76_360 ();
 sg13g2_decap_8 FILLER_76_367 ();
 sg13g2_decap_8 FILLER_76_374 ();
 sg13g2_decap_8 FILLER_76_381 ();
 sg13g2_decap_8 FILLER_76_388 ();
 sg13g2_decap_8 FILLER_76_395 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_fill_1 FILLER_77_84 ();
 sg13g2_decap_4 FILLER_77_111 ();
 sg13g2_fill_2 FILLER_77_115 ();
 sg13g2_fill_1 FILLER_77_143 ();
 sg13g2_fill_1 FILLER_77_206 ();
 sg13g2_fill_2 FILLER_77_216 ();
 sg13g2_decap_8 FILLER_77_309 ();
 sg13g2_decap_8 FILLER_77_316 ();
 sg13g2_decap_8 FILLER_77_323 ();
 sg13g2_decap_8 FILLER_77_330 ();
 sg13g2_decap_8 FILLER_77_337 ();
 sg13g2_decap_8 FILLER_77_344 ();
 sg13g2_decap_8 FILLER_77_351 ();
 sg13g2_decap_8 FILLER_77_358 ();
 sg13g2_decap_8 FILLER_77_365 ();
 sg13g2_decap_8 FILLER_77_372 ();
 sg13g2_decap_8 FILLER_77_379 ();
 sg13g2_decap_8 FILLER_77_386 ();
 sg13g2_decap_8 FILLER_77_393 ();
 sg13g2_decap_8 FILLER_77_400 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_135 ();
 sg13g2_decap_4 FILLER_78_142 ();
 sg13g2_fill_1 FILLER_78_146 ();
 sg13g2_fill_1 FILLER_78_208 ();
 sg13g2_fill_1 FILLER_78_213 ();
 sg13g2_fill_1 FILLER_78_255 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_4 FILLER_79_84 ();
 sg13g2_fill_2 FILLER_79_88 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_fill_2 FILLER_79_161 ();
 sg13g2_fill_2 FILLER_79_173 ();
 sg13g2_fill_1 FILLER_79_175 ();
 sg13g2_fill_2 FILLER_79_181 ();
 sg13g2_fill_2 FILLER_79_192 ();
 sg13g2_fill_2 FILLER_79_224 ();
 sg13g2_fill_1 FILLER_79_252 ();
 sg13g2_fill_1 FILLER_79_262 ();
 sg13g2_fill_2 FILLER_79_289 ();
 sg13g2_fill_1 FILLER_79_291 ();
 sg13g2_decap_8 FILLER_79_310 ();
 sg13g2_decap_8 FILLER_79_317 ();
 sg13g2_decap_8 FILLER_79_324 ();
 sg13g2_decap_8 FILLER_79_331 ();
 sg13g2_decap_8 FILLER_79_338 ();
 sg13g2_decap_8 FILLER_79_345 ();
 sg13g2_decap_8 FILLER_79_352 ();
 sg13g2_decap_8 FILLER_79_359 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_decap_8 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_8 FILLER_80_68 ();
 sg13g2_decap_8 FILLER_80_75 ();
 sg13g2_decap_4 FILLER_80_82 ();
 sg13g2_fill_2 FILLER_80_86 ();
 sg13g2_fill_2 FILLER_80_92 ();
 sg13g2_fill_1 FILLER_80_94 ();
 sg13g2_decap_8 FILLER_80_121 ();
 sg13g2_decap_8 FILLER_80_128 ();
 sg13g2_decap_8 FILLER_80_135 ();
 sg13g2_decap_8 FILLER_80_142 ();
 sg13g2_decap_8 FILLER_80_149 ();
 sg13g2_decap_8 FILLER_80_156 ();
 sg13g2_decap_8 FILLER_80_163 ();
 sg13g2_decap_8 FILLER_80_170 ();
 sg13g2_fill_2 FILLER_80_193 ();
 sg13g2_fill_1 FILLER_80_195 ();
 sg13g2_fill_1 FILLER_80_212 ();
 sg13g2_fill_1 FILLER_80_230 ();
 sg13g2_decap_8 FILLER_80_308 ();
 sg13g2_decap_4 FILLER_80_315 ();
 sg13g2_fill_1 FILLER_80_319 ();
 sg13g2_decap_4 FILLER_80_324 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_8 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_347 ();
 sg13g2_decap_8 FILLER_80_354 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_decap_8 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_382 ();
 sg13g2_decap_8 FILLER_80_389 ();
 sg13g2_decap_8 FILLER_80_396 ();
 sg13g2_decap_4 FILLER_80_403 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net257;
 assign uio_oe[3] = net258;
 assign uio_oe[6] = net259;
 assign uio_oe[7] = net260;
 assign uo_out[0] = net8;
 assign uo_out[1] = net9;
 assign uo_out[2] = net10;
 assign uo_out[3] = net11;
 assign uo_out[4] = net12;
 assign uo_out[5] = net13;
 assign uo_out[6] = net14;
endmodule

module tt_um_tappu_tobias1012 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \ChiselTop.tappu.cpuState[0] ;
 wire \ChiselTop.tappu.cpuState[1] ;
 wire \ChiselTop.tappu.cpuState[2] ;
 wire \ChiselTop.tappu.cpuState[3] ;
 wire \ChiselTop.tappu.cpuState[5] ;
 wire \ChiselTop.tappu.instrStepReg[0] ;
 wire \ChiselTop.tappu.instrStepReg[1] ;
 wire \ChiselTop.tappu.instrStepReg[2] ;
 wire \ChiselTop.tappu.instrStepReg[4] ;
 wire \ChiselTop.tappu.instrStepReg[5] ;
 wire \ChiselTop.tappu.mem._GEN_198[1] ;
 wire \ChiselTop.tappu.mem._GEN_198[2] ;
 wire \ChiselTop.tappu.mem._GEN_198[3] ;
 wire \ChiselTop.tappu.mem._GEN_198[4] ;
 wire \ChiselTop.tappu.mem._GEN_198[5] ;
 wire \ChiselTop.tappu.mem.state ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[0] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[10] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[11] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[12] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[13] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[14] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[15] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[1] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[2] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[3] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[4] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[5] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[6] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[7] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[8] ;
 wire \ChiselTop.tappu.mem.tapeCounterReg[9] ;
 wire \ChiselTop.tappu.mem.tape[0][0] ;
 wire \ChiselTop.tappu.mem.tape[0][1] ;
 wire \ChiselTop.tappu.mem.tape[0][2] ;
 wire \ChiselTop.tappu.mem.tape[0][3] ;
 wire \ChiselTop.tappu.mem.tape[0][4] ;
 wire \ChiselTop.tappu.mem.tape[0][5] ;
 wire \ChiselTop.tappu.mem.tape[0][6] ;
 wire \ChiselTop.tappu.mem.tape[0][7] ;
 wire \ChiselTop.tappu.mem.tape[1][0] ;
 wire \ChiselTop.tappu.mem.tape[1][1] ;
 wire \ChiselTop.tappu.mem.tape[1][2] ;
 wire \ChiselTop.tappu.mem.tape[1][3] ;
 wire \ChiselTop.tappu.mem.tape[1][4] ;
 wire \ChiselTop.tappu.mem.tape[1][5] ;
 wire \ChiselTop.tappu.mem.tape[1][6] ;
 wire \ChiselTop.tappu.mem.tape[1][7] ;
 wire \ChiselTop.tappu.mem.tape[2][0] ;
 wire \ChiselTop.tappu.mem.tape[2][1] ;
 wire \ChiselTop.tappu.mem.tape[2][2] ;
 wire \ChiselTop.tappu.mem.tape[2][3] ;
 wire \ChiselTop.tappu.mem.tape[2][4] ;
 wire \ChiselTop.tappu.mem.tape[2][5] ;
 wire \ChiselTop.tappu.mem.tape[2][6] ;
 wire \ChiselTop.tappu.mem.tape[2][7] ;
 wire \ChiselTop.tappu.mem.tape_readData_addr[0] ;
 wire \ChiselTop.tappu.mem.tape_readData_addr[1] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire net19;
 wire net18;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire clknet_0_clk;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net1;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;

 sg13g2_inv_1 _0696_ (.Y(_0089_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[12] ));
 sg13g2_inv_1 _0697_ (.Y(_0090_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[11] ));
 sg13g2_inv_1 _0698_ (.Y(_0091_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[10] ));
 sg13g2_inv_1 _0699_ (.Y(_0092_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[8] ));
 sg13g2_inv_1 _0700_ (.Y(_0093_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[7] ));
 sg13g2_inv_1 _0701_ (.Y(_0094_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[4] ));
 sg13g2_inv_1 _0702_ (.Y(_0095_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[2] ));
 sg13g2_inv_1 _0703_ (.Y(_0096_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[0] ));
 sg13g2_inv_1 _0704_ (.Y(_0097_),
    .A(\ChiselTop.tappu.mem._GEN_198[4] ));
 sg13g2_inv_1 _0705_ (.Y(_0098_),
    .A(net135));
 sg13g2_inv_1 _0706_ (.Y(_0099_),
    .A(net138));
 sg13g2_inv_1 _0707_ (.Y(_0100_),
    .A(net133));
 sg13g2_inv_1 _0708_ (.Y(_0101_),
    .A(net123));
 sg13g2_inv_1 _0709_ (.Y(_0102_),
    .A(_0016_));
 sg13g2_inv_1 _0710_ (.Y(_0103_),
    .A(_0018_));
 sg13g2_inv_1 _0711_ (.Y(_0104_),
    .A(_0020_));
 sg13g2_inv_1 _0712_ (.Y(_0105_),
    .A(_0017_));
 sg13g2_inv_1 _0713_ (.Y(_0106_),
    .A(net202));
 sg13g2_inv_2 _0714_ (.Y(_0107_),
    .A(net181));
 sg13g2_nand2b_1 _0715_ (.Y(_0108_),
    .B(net132),
    .A_N(\ChiselTop.tappu.mem.tape[1][5] ));
 sg13g2_nor2_1 _0716_ (.A(net132),
    .B(\ChiselTop.tappu.mem.tape[0][5] ),
    .Y(_0109_));
 sg13g2_nor2_1 _0717_ (.A(net130),
    .B(_0109_),
    .Y(_0110_));
 sg13g2_a22oi_1 _0718_ (.Y(_0111_),
    .B1(_0108_),
    .B2(_0110_),
    .A2(net148),
    .A1(net130));
 sg13g2_inv_1 _0719_ (.Y(_0112_),
    .A(_0111_));
 sg13g2_nor2_1 _0720_ (.A(net123),
    .B(_0111_),
    .Y(_0113_));
 sg13g2_inv_1 _0721_ (.Y(_0114_),
    .A(_0113_));
 sg13g2_nand2b_1 _0722_ (.Y(_0115_),
    .B(net132),
    .A_N(\ChiselTop.tappu.mem.tape[1][7] ));
 sg13g2_nor2_1 _0723_ (.A(net132),
    .B(\ChiselTop.tappu.mem.tape[0][7] ),
    .Y(_0116_));
 sg13g2_nor2_1 _0724_ (.A(net130),
    .B(_0116_),
    .Y(_0117_));
 sg13g2_a22oi_1 _0725_ (.Y(_0118_),
    .B1(_0115_),
    .B2(_0117_),
    .A2(net106),
    .A1(net130));
 sg13g2_nor2_1 _0726_ (.A(net122),
    .B(_0118_),
    .Y(_0119_));
 sg13g2_inv_1 _0727_ (.Y(_0120_),
    .A(_0119_));
 sg13g2_nand2b_1 _0728_ (.Y(_0121_),
    .B(net132),
    .A_N(\ChiselTop.tappu.mem.tape[1][4] ));
 sg13g2_nor2_1 _0729_ (.A(net132),
    .B(\ChiselTop.tappu.mem.tape[0][4] ),
    .Y(_0122_));
 sg13g2_nor2_1 _0730_ (.A(net130),
    .B(_0122_),
    .Y(_0123_));
 sg13g2_a22oi_1 _0731_ (.Y(_0124_),
    .B1(_0121_),
    .B2(_0123_),
    .A2(\ChiselTop.tappu.mem.tape[2][4] ),
    .A1(net130));
 sg13g2_inv_1 _0732_ (.Y(_0125_),
    .A(_0124_));
 sg13g2_nand2_1 _0733_ (.Y(_0126_),
    .A(_0101_),
    .B(_0125_));
 sg13g2_nand2b_1 _0734_ (.Y(_0127_),
    .B(net132),
    .A_N(\ChiselTop.tappu.mem.tape[1][6] ));
 sg13g2_nor2_1 _0735_ (.A(net132),
    .B(\ChiselTop.tappu.mem.tape[0][6] ),
    .Y(_0128_));
 sg13g2_nor2_1 _0736_ (.A(net130),
    .B(_0128_),
    .Y(_0129_));
 sg13g2_a22oi_1 _0737_ (.Y(_0130_),
    .B1(_0127_),
    .B2(_0129_),
    .A2(\ChiselTop.tappu.mem.tape[2][6] ),
    .A1(net130));
 sg13g2_or2_1 _0738_ (.X(_0131_),
    .B(_0130_),
    .A(net122));
 sg13g2_and4_1 _0739_ (.A(_0114_),
    .B(_0120_),
    .C(_0126_),
    .D(_0131_),
    .X(_0132_));
 sg13g2_nand2b_1 _0740_ (.Y(_0133_),
    .B(net131),
    .A_N(\ChiselTop.tappu.mem.tape[1][0] ));
 sg13g2_nor2_1 _0741_ (.A(\ChiselTop.tappu.mem.tape[0][0] ),
    .B(net131),
    .Y(_0134_));
 sg13g2_nor2_1 _0742_ (.A(net129),
    .B(_0134_),
    .Y(_0135_));
 sg13g2_a22oi_1 _0743_ (.Y(_0136_),
    .B1(_0133_),
    .B2(_0135_),
    .A2(net129),
    .A1(\ChiselTop.tappu.mem.tape[2][0] ));
 sg13g2_inv_1 _0744_ (.Y(_0137_),
    .A(_0136_));
 sg13g2_nand2_1 _0745_ (.Y(_0138_),
    .A(_0101_),
    .B(_0137_));
 sg13g2_nand2b_1 _0746_ (.Y(_0139_),
    .B(net131),
    .A_N(\ChiselTop.tappu.mem.tape[1][1] ));
 sg13g2_nor2_1 _0747_ (.A(net131),
    .B(\ChiselTop.tappu.mem.tape[0][1] ),
    .Y(_0140_));
 sg13g2_nor2_1 _0748_ (.A(net129),
    .B(_0140_),
    .Y(_0141_));
 sg13g2_a22oi_1 _0749_ (.Y(_0142_),
    .B1(_0139_),
    .B2(_0141_),
    .A2(\ChiselTop.tappu.mem.tape[2][1] ),
    .A1(net129));
 sg13g2_or2_1 _0750_ (.X(_0143_),
    .B(_0142_),
    .A(net122));
 sg13g2_nand2b_1 _0751_ (.Y(_0144_),
    .B(net131),
    .A_N(\ChiselTop.tappu.mem.tape[1][3] ));
 sg13g2_nor2_1 _0752_ (.A(net131),
    .B(\ChiselTop.tappu.mem.tape[0][3] ),
    .Y(_0145_));
 sg13g2_nor2_1 _0753_ (.A(net129),
    .B(_0145_),
    .Y(_0146_));
 sg13g2_a22oi_1 _0754_ (.Y(_0147_),
    .B1(_0144_),
    .B2(_0146_),
    .A2(\ChiselTop.tappu.mem.tape[2][3] ),
    .A1(net129));
 sg13g2_or2_1 _0755_ (.X(_0148_),
    .B(_0147_),
    .A(net122));
 sg13g2_nand2b_1 _0756_ (.Y(_0149_),
    .B(net131),
    .A_N(\ChiselTop.tappu.mem.tape[1][2] ));
 sg13g2_nor2_1 _0757_ (.A(net131),
    .B(\ChiselTop.tappu.mem.tape[0][2] ),
    .Y(_0150_));
 sg13g2_nor2_1 _0758_ (.A(net129),
    .B(_0150_),
    .Y(_0151_));
 sg13g2_a22oi_1 _0759_ (.Y(_0152_),
    .B1(_0149_),
    .B2(_0151_),
    .A2(\ChiselTop.tappu.mem.tape[2][2] ),
    .A1(net129));
 sg13g2_inv_1 _0760_ (.Y(_0153_),
    .A(_0152_));
 sg13g2_nand2_1 _0761_ (.Y(_0154_),
    .A(_0101_),
    .B(_0153_));
 sg13g2_and2_1 _0762_ (.A(_0148_),
    .B(_0154_),
    .X(_0155_));
 sg13g2_and4_1 _0763_ (.A(_0132_),
    .B(_0138_),
    .C(_0143_),
    .D(_0155_),
    .X(_0156_));
 sg13g2_nor2b_2 _0764_ (.A(net138),
    .B_N(\ChiselTop.tappu.mem._GEN_198[1] ),
    .Y(_0157_));
 sg13g2_nand2b_2 _0765_ (.Y(_0158_),
    .B(\ChiselTop.tappu.mem._GEN_198[1] ),
    .A_N(\ChiselTop.tappu.mem._GEN_198[2] ));
 sg13g2_nor2b_1 _0766_ (.A(net135),
    .B_N(net133),
    .Y(_0159_));
 sg13g2_nand2b_1 _0767_ (.Y(_0160_),
    .B(net133),
    .A_N(net135));
 sg13g2_nand3b_1 _0768_ (.B(net133),
    .C(\ChiselTop.tappu.mem._GEN_198[4] ),
    .Y(_0161_),
    .A_N(net136));
 sg13g2_or2_1 _0769_ (.X(_0162_),
    .B(_0161_),
    .A(_0158_));
 sg13g2_nor2b_1 _0770_ (.A(net134),
    .B_N(\ChiselTop.tappu.mem._GEN_198[5] ),
    .Y(_0163_));
 sg13g2_nand2b_1 _0771_ (.Y(_0164_),
    .B(\ChiselTop.tappu.mem._GEN_198[5] ),
    .A_N(net134));
 sg13g2_or2_1 _0772_ (.X(_0165_),
    .B(\ChiselTop.tappu.mem._GEN_198[1] ),
    .A(\ChiselTop.tappu.mem._GEN_198[2] ));
 sg13g2_nand3b_1 _0773_ (.B(net136),
    .C(\ChiselTop.tappu.mem._GEN_198[5] ),
    .Y(_0166_),
    .A_N(net134));
 sg13g2_or2_1 _0774_ (.X(_0167_),
    .B(_0166_),
    .A(_0165_));
 sg13g2_nor2_1 _0775_ (.A(net135),
    .B(_0164_),
    .Y(_0168_));
 sg13g2_nand3_1 _0776_ (.B(_0157_),
    .C(_0163_),
    .A(_0098_),
    .Y(_0169_));
 sg13g2_nand3_1 _0777_ (.B(_0167_),
    .C(_0169_),
    .A(_0162_),
    .Y(_0170_));
 sg13g2_nor2b_1 _0778_ (.A(_0156_),
    .B_N(_0170_),
    .Y(_0171_));
 sg13g2_nand4_1 _0779_ (.B(net140),
    .C(\ChiselTop.tappu.cpuState[2] ),
    .A(net124),
    .Y(_0172_),
    .D(_0171_));
 sg13g2_nand3b_1 _0780_ (.B(_0172_),
    .C(net140),
    .Y(_0005_),
    .A_N(net88));
 sg13g2_nand2b_2 _0781_ (.Y(_0173_),
    .B(\ChiselTop.tappu.mem._GEN_198[2] ),
    .A_N(\ChiselTop.tappu.mem._GEN_198[1] ));
 sg13g2_and4_1 _0782_ (.A(net136),
    .B(net133),
    .C(_0158_),
    .D(_0173_),
    .X(_0174_));
 sg13g2_nand4_1 _0783_ (.B(net133),
    .C(_0158_),
    .A(net135),
    .Y(_0175_),
    .D(_0173_));
 sg13g2_nand2_1 _0784_ (.Y(_0176_),
    .A(_0097_),
    .B(_0159_));
 sg13g2_nand3_1 _0785_ (.B(_0157_),
    .C(_0159_),
    .A(_0097_),
    .Y(_0177_));
 sg13g2_o21ai_1 _0786_ (.B1(net124),
    .Y(_0178_),
    .A1(_0165_),
    .A2(_0166_));
 sg13g2_nor2b_1 _0787_ (.A(_0178_),
    .B_N(_0169_),
    .Y(_0179_));
 sg13g2_nand2b_1 _0788_ (.Y(_0180_),
    .B(_0169_),
    .A_N(_0178_));
 sg13g2_a221oi_1 _0789_ (.B2(_0177_),
    .C1(_0178_),
    .B1(_0175_),
    .A1(_0157_),
    .Y(_0181_),
    .A2(_0168_));
 sg13g2_a21o_1 _0790_ (.A2(_0170_),
    .A1(net124),
    .B1(_0181_),
    .X(_0182_));
 sg13g2_nor4_2 _0791_ (.A(\ChiselTop.tappu.mem._GEN_198[5] ),
    .B(_0097_),
    .C(net135),
    .Y(_0183_),
    .D(_0173_));
 sg13g2_nor3_1 _0792_ (.A(net135),
    .B(_0164_),
    .C(_0165_),
    .Y(_0184_));
 sg13g2_nor2_2 _0793_ (.A(_0183_),
    .B(_0184_),
    .Y(_0185_));
 sg13g2_nor3_2 _0794_ (.A(net136),
    .B(_0099_),
    .C(_0164_),
    .Y(_0186_));
 sg13g2_nand3_1 _0795_ (.B(net138),
    .C(_0163_),
    .A(_0098_),
    .Y(_0187_));
 sg13g2_nand4_1 _0796_ (.B(_0158_),
    .C(_0159_),
    .A(net134),
    .Y(_0188_),
    .D(_0173_));
 sg13g2_and4_2 _0797_ (.A(_0175_),
    .B(_0177_),
    .C(_0187_),
    .D(_0188_),
    .X(_0189_));
 sg13g2_nand2_1 _0798_ (.Y(_0190_),
    .A(_0185_),
    .B(_0189_));
 sg13g2_o21ai_1 _0799_ (.B1(net124),
    .Y(_0191_),
    .A1(_0170_),
    .A2(_0190_));
 sg13g2_o21ai_1 _0800_ (.B1(_0182_),
    .Y(_0192_),
    .A1(_0171_),
    .A2(_0191_));
 sg13g2_and3_1 _0801_ (.X(_0006_),
    .A(net140),
    .B(net96),
    .C(_0192_));
 sg13g2_nor2_1 _0802_ (.A(net127),
    .B(net94),
    .Y(_0193_));
 sg13g2_a21oi_1 _0803_ (.A1(net119),
    .A2(net127),
    .Y(_0007_),
    .B1(_0193_));
 sg13g2_mux2_1 _0804_ (.A0(net91),
    .A1(net121),
    .S(net127),
    .X(_0008_));
 sg13g2_and2_1 _0805_ (.A(net139),
    .B(net193),
    .X(_0004_));
 sg13g2_and2_1 _0806_ (.A(net140),
    .B(net87),
    .X(_0002_));
 sg13g2_and2_1 _0807_ (.A(net140),
    .B(net90),
    .X(_0003_));
 sg13g2_and2_2 _0808_ (.A(net124),
    .B(\ChiselTop.tappu.cpuState[0] ),
    .X(_0194_));
 sg13g2_nand2_2 _0809_ (.Y(_0195_),
    .A(net124),
    .B(net193));
 sg13g2_or3_1 _0810_ (.A(\ChiselTop.tappu.instrStepReg[0] ),
    .B(\ChiselTop.tappu.instrStepReg[1] ),
    .C(\ChiselTop.tappu.instrStepReg[2] ),
    .X(_0196_));
 sg13g2_or2_1 _0811_ (.X(_0197_),
    .B(_0196_),
    .A(\ChiselTop.tappu.instrStepReg[4] ));
 sg13g2_nor2b_1 _0812_ (.A(\ChiselTop.tappu.instrStepReg[0] ),
    .B_N(\ChiselTop.tappu.cpuState[0] ),
    .Y(_0198_));
 sg13g2_o21ai_1 _0813_ (.B1(\ChiselTop.tappu.cpuState[0] ),
    .Y(_0199_),
    .A1(\ChiselTop.tappu.instrStepReg[0] ),
    .A2(\ChiselTop.tappu.instrStepReg[1] ));
 sg13g2_and2_1 _0814_ (.A(\ChiselTop.tappu.cpuState[0] ),
    .B(_0196_),
    .X(_0200_));
 sg13g2_nand2_1 _0815_ (.Y(_0201_),
    .A(\ChiselTop.tappu.cpuState[0] ),
    .B(_0197_));
 sg13g2_o21ai_1 _0816_ (.B1(_0198_),
    .Y(_0202_),
    .A1(\ChiselTop.tappu.instrStepReg[5] ),
    .A2(_0197_));
 sg13g2_a21oi_1 _0817_ (.A1(_0194_),
    .A2(_0202_),
    .Y(_0203_),
    .B1(net172));
 sg13g2_nand2_1 _0818_ (.Y(_0204_),
    .A(\ChiselTop.tappu.mem._GEN_198[1] ),
    .B(_0202_));
 sg13g2_o21ai_1 _0819_ (.B1(net142),
    .Y(_0205_),
    .A1(_0195_),
    .A2(_0204_));
 sg13g2_nor2_1 _0820_ (.A(net173),
    .B(_0205_),
    .Y(_0028_));
 sg13g2_a21oi_1 _0821_ (.A1(\ChiselTop.tappu.instrStepReg[0] ),
    .A2(\ChiselTop.tappu.instrStepReg[1] ),
    .Y(_0206_),
    .B1(_0199_));
 sg13g2_nand2_1 _0822_ (.Y(_0207_),
    .A(net138),
    .B(_0206_));
 sg13g2_xnor2_1 _0823_ (.Y(_0208_),
    .A(net138),
    .B(_0206_));
 sg13g2_or2_1 _0824_ (.X(_0209_),
    .B(_0208_),
    .A(_0204_));
 sg13g2_xor2_1 _0825_ (.B(_0208_),
    .A(_0204_),
    .X(_0210_));
 sg13g2_o21ai_1 _0826_ (.B1(net142),
    .Y(_0211_),
    .A1(_0195_),
    .A2(_0210_));
 sg13g2_a21oi_1 _0827_ (.A1(_0099_),
    .A2(_0195_),
    .Y(_0029_),
    .B1(_0211_));
 sg13g2_o21ai_1 _0828_ (.B1(\ChiselTop.tappu.instrStepReg[2] ),
    .Y(_0212_),
    .A1(\ChiselTop.tappu.instrStepReg[0] ),
    .A2(\ChiselTop.tappu.instrStepReg[1] ));
 sg13g2_nand3_1 _0829_ (.B(_0200_),
    .C(_0212_),
    .A(net137),
    .Y(_0213_));
 sg13g2_a21o_1 _0830_ (.A2(_0212_),
    .A1(_0200_),
    .B1(net137),
    .X(_0214_));
 sg13g2_nand2_1 _0831_ (.Y(_0215_),
    .A(_0213_),
    .B(_0214_));
 sg13g2_nand3_1 _0832_ (.B(_0209_),
    .C(_0215_),
    .A(_0207_),
    .Y(_0216_));
 sg13g2_a21o_1 _0833_ (.A2(_0209_),
    .A1(_0207_),
    .B1(_0215_),
    .X(_0217_));
 sg13g2_a21oi_1 _0834_ (.A1(_0216_),
    .A2(_0217_),
    .Y(_0218_),
    .B1(_0195_));
 sg13g2_o21ai_1 _0835_ (.B1(net142),
    .Y(_0219_),
    .A1(net137),
    .A2(_0194_));
 sg13g2_nor2_1 _0836_ (.A(_0218_),
    .B(_0219_),
    .Y(_0030_));
 sg13g2_nor2_1 _0837_ (.A(\ChiselTop.tappu.instrStepReg[2] ),
    .B(_0199_),
    .Y(_0220_));
 sg13g2_xnor2_1 _0838_ (.Y(_0221_),
    .A(net134),
    .B(_0220_));
 sg13g2_and3_1 _0839_ (.X(_0222_),
    .A(_0213_),
    .B(_0217_),
    .C(_0221_));
 sg13g2_a21oi_1 _0840_ (.A1(_0213_),
    .A2(_0217_),
    .Y(_0223_),
    .B1(_0221_));
 sg13g2_o21ai_1 _0841_ (.B1(_0194_),
    .Y(_0224_),
    .A1(_0222_),
    .A2(_0223_));
 sg13g2_o21ai_1 _0842_ (.B1(net142),
    .Y(_0225_),
    .A1(net134),
    .A2(_0194_));
 sg13g2_nor2b_1 _0843_ (.A(_0225_),
    .B_N(_0224_),
    .Y(_0031_));
 sg13g2_a21oi_1 _0844_ (.A1(net134),
    .A2(_0220_),
    .Y(_0226_),
    .B1(_0223_));
 sg13g2_a21oi_1 _0845_ (.A1(\ChiselTop.tappu.instrStepReg[4] ),
    .A2(_0196_),
    .Y(_0227_),
    .B1(_0201_));
 sg13g2_xnor2_1 _0846_ (.Y(_0228_),
    .A(net133),
    .B(_0227_));
 sg13g2_o21ai_1 _0847_ (.B1(_0194_),
    .Y(_0229_),
    .A1(_0226_),
    .A2(_0228_));
 sg13g2_a21oi_1 _0848_ (.A1(_0226_),
    .A2(_0228_),
    .Y(_0230_),
    .B1(_0229_));
 sg13g2_o21ai_1 _0849_ (.B1(net142),
    .Y(_0231_),
    .A1(net178),
    .A2(_0194_));
 sg13g2_nor2_1 _0850_ (.A(_0230_),
    .B(_0231_),
    .Y(_0032_));
 sg13g2_nor4_2 _0851_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[13] ),
    .B(\ChiselTop.tappu.mem.tapeCounterReg[12] ),
    .C(\ChiselTop.tappu.mem.tapeCounterReg[11] ),
    .Y(_0232_),
    .D(\ChiselTop.tappu.mem.tapeCounterReg[10] ));
 sg13g2_nor4_1 _0852_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[15] ),
    .B(\ChiselTop.tappu.mem.tapeCounterReg[14] ),
    .C(\ChiselTop.tappu.mem.tapeCounterReg[9] ),
    .D(net120),
    .Y(_0233_));
 sg13g2_nand2_2 _0853_ (.Y(_0234_),
    .A(_0232_),
    .B(_0233_));
 sg13g2_nor4_1 _0854_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[7] ),
    .B(\ChiselTop.tappu.mem.tapeCounterReg[6] ),
    .C(\ChiselTop.tappu.mem.tapeCounterReg[5] ),
    .D(\ChiselTop.tappu.mem.tapeCounterReg[2] ),
    .Y(_0235_));
 sg13g2_nor2_1 _0855_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[4] ),
    .B(\ChiselTop.tappu.mem.tapeCounterReg[3] ),
    .Y(_0236_));
 sg13g2_nand2_1 _0856_ (.Y(_0237_),
    .A(net121),
    .B(\ChiselTop.tappu.mem.tapeCounterReg[0] ));
 sg13g2_nand4_1 _0857_ (.B(\ChiselTop.tappu.mem.tapeCounterReg[0] ),
    .C(_0235_),
    .A(net121),
    .Y(_0238_),
    .D(_0236_));
 sg13g2_nor2_1 _0858_ (.A(_0234_),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_o21ai_1 _0859_ (.B1(net123),
    .Y(_0240_),
    .A1(_0234_),
    .A2(_0238_));
 sg13g2_nand3b_1 _0860_ (.B(net133),
    .C(net136),
    .Y(_0241_),
    .A_N(net138));
 sg13g2_o21ai_1 _0861_ (.B1(_0241_),
    .Y(_0242_),
    .A1(_0158_),
    .A2(_0161_));
 sg13g2_nor3_1 _0862_ (.A(net134),
    .B(_0160_),
    .C(_0173_),
    .Y(_0243_));
 sg13g2_nor4_2 _0863_ (.A(_0183_),
    .B(_0186_),
    .C(_0242_),
    .Y(_0244_),
    .D(_0243_));
 sg13g2_nand2_2 _0864_ (.Y(_0245_),
    .A(_0179_),
    .B(_0244_));
 sg13g2_a21o_2 _0865_ (.A2(_0189_),
    .A1(_0185_),
    .B1(_0180_),
    .X(_0246_));
 sg13g2_nor2_1 _0866_ (.A(_0190_),
    .B(_0245_),
    .Y(_0247_));
 sg13g2_nand2b_2 _0867_ (.Y(_0248_),
    .B(_0246_),
    .A_N(_0245_));
 sg13g2_nor2b_1 _0868_ (.A(\ChiselTop.tappu.cpuState[3] ),
    .B_N(_0015_),
    .Y(_0249_));
 sg13g2_nor2b_2 _0869_ (.A(_0014_),
    .B_N(_0249_),
    .Y(_0250_));
 sg13g2_nand2b_2 _0870_ (.Y(_0251_),
    .B(_0249_),
    .A_N(_0014_));
 sg13g2_nand2_2 _0871_ (.Y(_0252_),
    .A(net128),
    .B(_0250_));
 sg13g2_nor2_2 _0872_ (.A(_0248_),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_or2_1 _0873_ (.X(_0254_),
    .B(_0252_),
    .A(_0248_));
 sg13g2_nand2_1 _0874_ (.Y(_0255_),
    .A(_0240_),
    .B(_0254_));
 sg13g2_nand3_1 _0875_ (.B(_0167_),
    .C(_0169_),
    .A(_0101_),
    .Y(_0256_));
 sg13g2_a21oi_2 _0876_ (.B1(_0256_),
    .Y(_0257_),
    .A2(_0189_),
    .A1(_0185_));
 sg13g2_a21o_1 _0877_ (.A2(_0189_),
    .A1(_0185_),
    .B1(_0256_),
    .X(_0258_));
 sg13g2_nor3_1 _0878_ (.A(_0182_),
    .B(_0245_),
    .C(_0258_),
    .Y(_0259_));
 sg13g2_and4_1 _0879_ (.A(_0179_),
    .B(_0190_),
    .C(_0250_),
    .D(_0259_),
    .X(_0260_));
 sg13g2_or2_1 _0880_ (.X(_0261_),
    .B(_0260_),
    .A(_0255_));
 sg13g2_nor2_1 _0881_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[1] ),
    .B(net119),
    .Y(_0262_));
 sg13g2_nand2_2 _0882_ (.Y(_0263_),
    .A(_0261_),
    .B(_0262_));
 sg13g2_nor3_1 _0883_ (.A(_0174_),
    .B(_0183_),
    .C(_0184_),
    .Y(_0264_));
 sg13g2_nand3_1 _0884_ (.B(_0013_),
    .C(_0157_),
    .A(net135),
    .Y(_0265_));
 sg13g2_nand2_1 _0885_ (.Y(_0266_),
    .A(_0176_),
    .B(_0265_));
 sg13g2_and3_1 _0886_ (.X(_0267_),
    .A(_0176_),
    .B(_0188_),
    .C(_0265_));
 sg13g2_a22oi_1 _0887_ (.Y(_0268_),
    .B1(_0264_),
    .B2(_0267_),
    .A2(_0168_),
    .A1(_0157_));
 sg13g2_nand2_1 _0888_ (.Y(_0269_),
    .A(_0167_),
    .B(_0187_));
 sg13g2_o21ai_1 _0889_ (.B1(_0101_),
    .Y(_0270_),
    .A1(_0268_),
    .A2(_0269_));
 sg13g2_and2_1 _0890_ (.A(\ChiselTop.tappu.cpuState[2] ),
    .B(_0249_),
    .X(_0271_));
 sg13g2_o21ai_1 _0891_ (.B1(_0271_),
    .Y(_0272_),
    .A1(_0247_),
    .A2(_0259_));
 sg13g2_or2_1 _0892_ (.X(_0273_),
    .B(_0272_),
    .A(_0270_));
 sg13g2_nand2_1 _0893_ (.Y(_0274_),
    .A(_0137_),
    .B(_0273_));
 sg13g2_nor3_1 _0894_ (.A(_0137_),
    .B(_0270_),
    .C(_0272_),
    .Y(_0275_));
 sg13g2_xnor2_1 _0895_ (.Y(_0276_),
    .A(_0136_),
    .B(_0273_));
 sg13g2_nor2_1 _0896_ (.A(_0161_),
    .B(_0165_),
    .Y(_0277_));
 sg13g2_nor3_1 _0897_ (.A(_0098_),
    .B(_0100_),
    .C(_0173_),
    .Y(_0278_));
 sg13g2_nand2_1 _0898_ (.Y(_0279_),
    .A(net138),
    .B(\ChiselTop.tappu.mem._GEN_198[1] ));
 sg13g2_nand2_1 _0899_ (.Y(_0280_),
    .A(_0266_),
    .B(_0279_));
 sg13g2_nor4_1 _0900_ (.A(net122),
    .B(_0170_),
    .C(_0277_),
    .D(_0278_),
    .Y(_0281_));
 sg13g2_nand4_1 _0901_ (.B(_0264_),
    .C(_0280_),
    .A(_0187_),
    .Y(_0282_),
    .D(_0281_));
 sg13g2_or2_1 _0902_ (.X(_0283_),
    .B(_0282_),
    .A(_0272_));
 sg13g2_nand2_1 _0903_ (.Y(_0284_),
    .A(_0112_),
    .B(_0283_));
 sg13g2_inv_1 _0904_ (.Y(_0285_),
    .A(_0284_));
 sg13g2_or2_1 _0905_ (.X(_0286_),
    .B(_0283_),
    .A(_0112_));
 sg13g2_and2_1 _0906_ (.A(_0284_),
    .B(_0286_),
    .X(_0287_));
 sg13g2_nand2_1 _0907_ (.Y(_0288_),
    .A(_0284_),
    .B(_0286_));
 sg13g2_or2_1 _0908_ (.X(_0289_),
    .B(_0279_),
    .A(_0160_));
 sg13g2_or4_1 _0909_ (.A(_0160_),
    .B(_0168_),
    .C(_0252_),
    .D(_0279_),
    .X(_0290_));
 sg13g2_a21oi_2 _0910_ (.B1(_0290_),
    .Y(_0291_),
    .A2(_0248_),
    .A1(net122));
 sg13g2_a21o_2 _0911_ (.A2(_0248_),
    .A1(net122),
    .B1(_0290_),
    .X(_0292_));
 sg13g2_xnor2_1 _0912_ (.Y(_0293_),
    .A(_0118_),
    .B(net118));
 sg13g2_inv_1 _0913_ (.Y(_0294_),
    .A(_0293_));
 sg13g2_nor2_1 _0914_ (.A(_0130_),
    .B(net118),
    .Y(_0295_));
 sg13g2_nand2b_1 _0915_ (.Y(_0296_),
    .B(_0291_),
    .A_N(_0130_));
 sg13g2_xnor2_1 _0916_ (.Y(_0297_),
    .A(_0130_),
    .B(_0292_));
 sg13g2_xnor2_1 _0917_ (.Y(_0298_),
    .A(_0130_),
    .B(_0291_));
 sg13g2_nor2_1 _0918_ (.A(_0293_),
    .B(_0298_),
    .Y(_0299_));
 sg13g2_nand2_1 _0919_ (.Y(_0300_),
    .A(_0248_),
    .B(_0258_));
 sg13g2_a221oi_1 _0920_ (.B2(_0244_),
    .C1(_0181_),
    .B1(_0179_),
    .A1(net124),
    .Y(_0301_),
    .A2(_0170_));
 sg13g2_nand2_1 _0921_ (.Y(_0302_),
    .A(_0257_),
    .B(_0301_));
 sg13g2_nand2b_1 _0922_ (.Y(_0303_),
    .B(_0289_),
    .A_N(_0278_));
 sg13g2_nand4_1 _0923_ (.B(_0300_),
    .C(_0302_),
    .A(_0271_),
    .Y(_0304_),
    .D(_0303_));
 sg13g2_nand2_1 _0924_ (.Y(_0305_),
    .A(_0125_),
    .B(_0304_));
 sg13g2_nor2_1 _0925_ (.A(_0125_),
    .B(_0304_),
    .Y(_0306_));
 sg13g2_xnor2_1 _0926_ (.Y(_0307_),
    .A(_0125_),
    .B(_0304_));
 sg13g2_inv_1 _0927_ (.Y(_0308_),
    .A(_0307_));
 sg13g2_nand3_1 _0928_ (.B(_0299_),
    .C(_0308_),
    .A(_0287_),
    .Y(_0309_));
 sg13g2_nand4_1 _0929_ (.B(_0167_),
    .C(_0169_),
    .A(_0162_),
    .Y(_0310_),
    .D(_0289_));
 sg13g2_a21oi_1 _0930_ (.A1(\ChiselTop.tappu.mem._GEN_198[1] ),
    .A2(_0186_),
    .Y(_0311_),
    .B1(net122));
 sg13g2_and2_1 _0931_ (.A(_0310_),
    .B(_0311_),
    .X(_0312_));
 sg13g2_inv_1 _0932_ (.Y(_0313_),
    .A(_0312_));
 sg13g2_nand4_1 _0933_ (.B(_0271_),
    .C(_0310_),
    .A(net138),
    .Y(_0314_),
    .D(_0311_));
 sg13g2_a221oi_1 _0934_ (.B2(_0246_),
    .C1(_0314_),
    .B1(_0301_),
    .A1(_0245_),
    .Y(_0315_),
    .A2(_0257_));
 sg13g2_nand2b_1 _0935_ (.Y(_0316_),
    .B(_0315_),
    .A_N(_0142_));
 sg13g2_or2_1 _0936_ (.X(_0317_),
    .B(_0315_),
    .A(_0142_));
 sg13g2_xnor2_1 _0937_ (.Y(_0318_),
    .A(_0142_),
    .B(_0315_));
 sg13g2_xor2_1 _0938_ (.B(_0315_),
    .A(_0142_),
    .X(_0319_));
 sg13g2_nor2_1 _0939_ (.A(_0275_),
    .B(_0318_),
    .Y(_0320_));
 sg13g2_nor2_1 _0940_ (.A(_0153_),
    .B(_0292_),
    .Y(_0321_));
 sg13g2_nor2_1 _0941_ (.A(_0152_),
    .B(net118),
    .Y(_0322_));
 sg13g2_xnor2_1 _0942_ (.Y(_0323_),
    .A(_0153_),
    .B(net118));
 sg13g2_nor2_1 _0943_ (.A(_0147_),
    .B(net118),
    .Y(_0324_));
 sg13g2_xnor2_1 _0944_ (.Y(_0325_),
    .A(_0147_),
    .B(net118));
 sg13g2_nor3_2 _0945_ (.A(_0321_),
    .B(_0322_),
    .C(_0325_),
    .Y(_0326_));
 sg13g2_nand2_1 _0946_ (.Y(_0327_),
    .A(_0274_),
    .B(_0326_));
 sg13g2_nor2_1 _0947_ (.A(_0309_),
    .B(_0327_),
    .Y(_0328_));
 sg13g2_o21ai_1 _0948_ (.B1(_0291_),
    .Y(_0329_),
    .A1(_0118_),
    .A2(_0130_));
 sg13g2_inv_1 _0949_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_nand2_1 _0950_ (.Y(_0331_),
    .A(_0284_),
    .B(_0306_));
 sg13g2_nand2_1 _0951_ (.Y(_0332_),
    .A(_0286_),
    .B(_0331_));
 sg13g2_a21oi_1 _0952_ (.A1(_0299_),
    .A2(_0332_),
    .Y(_0333_),
    .B1(_0330_));
 sg13g2_nand3_1 _0953_ (.B(_0317_),
    .C(_0326_),
    .A(_0274_),
    .Y(_0334_));
 sg13g2_o21ai_1 _0954_ (.B1(net118),
    .Y(_0335_),
    .A1(_0147_),
    .A2(_0152_));
 sg13g2_a21o_1 _0955_ (.A2(_0335_),
    .A1(_0334_),
    .B1(_0309_),
    .X(_0336_));
 sg13g2_a22oi_1 _0956_ (.Y(_0337_),
    .B1(_0333_),
    .B2(_0336_),
    .A2(_0328_),
    .A1(_0320_));
 sg13g2_nand2b_2 _0957_ (.Y(_0338_),
    .B(_0260_),
    .A_N(_0337_));
 sg13g2_a21oi_2 _0958_ (.B1(_0276_),
    .Y(_0339_),
    .A2(_0338_),
    .A1(_0254_));
 sg13g2_mux2_1 _0959_ (.A0(_0339_),
    .A1(net99),
    .S(_0263_),
    .X(_0033_));
 sg13g2_or4_1 _0960_ (.A(_0136_),
    .B(_0270_),
    .C(_0272_),
    .D(_0319_),
    .X(_0340_));
 sg13g2_o21ai_1 _0961_ (.B1(_0319_),
    .Y(_0341_),
    .A1(_0136_),
    .A2(_0273_));
 sg13g2_and2_1 _0962_ (.A(_0253_),
    .B(_0341_),
    .X(_0342_));
 sg13g2_and2_1 _0963_ (.A(_0275_),
    .B(_0318_),
    .X(_0343_));
 sg13g2_nor3_1 _0964_ (.A(_0320_),
    .B(_0338_),
    .C(_0343_),
    .Y(_0344_));
 sg13g2_a21o_1 _0965_ (.A2(_0342_),
    .A1(_0340_),
    .B1(_0344_),
    .X(_0345_));
 sg13g2_mux2_1 _0966_ (.A0(_0345_),
    .A1(net103),
    .S(_0263_),
    .X(_0034_));
 sg13g2_nand3_1 _0967_ (.B(_0323_),
    .C(_0340_),
    .A(_0316_),
    .Y(_0346_));
 sg13g2_a21oi_1 _0968_ (.A1(_0316_),
    .A2(_0340_),
    .Y(_0347_),
    .B1(_0323_));
 sg13g2_nand3b_1 _0969_ (.B(_0253_),
    .C(_0346_),
    .Y(_0348_),
    .A_N(_0347_));
 sg13g2_o21ai_1 _0970_ (.B1(_0317_),
    .Y(_0349_),
    .A1(_0275_),
    .A2(_0318_));
 sg13g2_xnor2_1 _0971_ (.Y(_0350_),
    .A(_0323_),
    .B(_0349_));
 sg13g2_o21ai_1 _0972_ (.B1(_0348_),
    .Y(_0351_),
    .A1(_0338_),
    .A2(_0350_));
 sg13g2_mux2_1 _0973_ (.A0(_0351_),
    .A1(net101),
    .S(_0263_),
    .X(_0035_));
 sg13g2_nor2_1 _0974_ (.A(_0152_),
    .B(_0292_),
    .Y(_0352_));
 sg13g2_or3_1 _0975_ (.A(_0325_),
    .B(_0347_),
    .C(_0352_),
    .X(_0353_));
 sg13g2_o21ai_1 _0976_ (.B1(_0325_),
    .Y(_0354_),
    .A1(_0347_),
    .A2(_0352_));
 sg13g2_nand3_1 _0977_ (.B(_0353_),
    .C(_0354_),
    .A(_0253_),
    .Y(_0355_));
 sg13g2_a21oi_1 _0978_ (.A1(_0323_),
    .A2(_0349_),
    .Y(_0356_),
    .B1(_0322_));
 sg13g2_xnor2_1 _0979_ (.Y(_0357_),
    .A(_0325_),
    .B(_0356_));
 sg13g2_o21ai_1 _0980_ (.B1(_0355_),
    .Y(_0358_),
    .A1(_0338_),
    .A2(_0357_));
 sg13g2_mux2_1 _0981_ (.A0(_0358_),
    .A1(net157),
    .S(_0263_),
    .X(_0036_));
 sg13g2_nand2b_1 _0982_ (.Y(_0359_),
    .B(net118),
    .A_N(_0147_));
 sg13g2_a21oi_1 _0983_ (.A1(_0354_),
    .A2(_0359_),
    .Y(_0360_),
    .B1(_0308_));
 sg13g2_nand3_1 _0984_ (.B(_0354_),
    .C(_0359_),
    .A(_0308_),
    .Y(_0361_));
 sg13g2_nand3b_1 _0985_ (.B(_0361_),
    .C(_0253_),
    .Y(_0362_),
    .A_N(_0360_));
 sg13g2_a221oi_1 _0986_ (.B2(_0349_),
    .C1(_0324_),
    .B1(_0326_),
    .A1(_0153_),
    .Y(_0363_),
    .A2(_0292_));
 sg13g2_xnor2_1 _0987_ (.Y(_0364_),
    .A(_0307_),
    .B(_0363_));
 sg13g2_o21ai_1 _0988_ (.B1(_0362_),
    .Y(_0365_),
    .A1(_0338_),
    .A2(_0364_));
 sg13g2_mux2_1 _0989_ (.A0(_0365_),
    .A1(net98),
    .S(_0263_),
    .X(_0037_));
 sg13g2_nor2_1 _0990_ (.A(_0124_),
    .B(_0304_),
    .Y(_0366_));
 sg13g2_o21ai_1 _0991_ (.B1(_0288_),
    .Y(_0367_),
    .A1(_0360_),
    .A2(_0366_));
 sg13g2_nor3_1 _0992_ (.A(_0288_),
    .B(_0360_),
    .C(_0366_),
    .Y(_0368_));
 sg13g2_nand3b_1 _0993_ (.B(_0253_),
    .C(_0367_),
    .Y(_0369_),
    .A_N(_0368_));
 sg13g2_o21ai_1 _0994_ (.B1(_0305_),
    .Y(_0370_),
    .A1(_0307_),
    .A2(_0363_));
 sg13g2_xnor2_1 _0995_ (.Y(_0371_),
    .A(_0287_),
    .B(_0370_));
 sg13g2_o21ai_1 _0996_ (.B1(_0369_),
    .Y(_0372_),
    .A1(_0338_),
    .A2(_0371_));
 sg13g2_mux2_1 _0997_ (.A0(_0372_),
    .A1(net97),
    .S(_0263_),
    .X(_0038_));
 sg13g2_nand2b_1 _0998_ (.Y(_0373_),
    .B(_0112_),
    .A_N(_0283_));
 sg13g2_a21o_1 _0999_ (.A2(_0373_),
    .A1(_0367_),
    .B1(_0297_),
    .X(_0374_));
 sg13g2_nand3_1 _1000_ (.B(_0367_),
    .C(_0373_),
    .A(_0297_),
    .Y(_0375_));
 sg13g2_nand3_1 _1001_ (.B(_0374_),
    .C(_0375_),
    .A(_0253_),
    .Y(_0376_));
 sg13g2_a21oi_1 _1002_ (.A1(_0287_),
    .A2(_0370_),
    .Y(_0377_),
    .B1(_0285_));
 sg13g2_nor2_1 _1003_ (.A(_0298_),
    .B(_0377_),
    .Y(_0378_));
 sg13g2_a21o_1 _1004_ (.A2(_0377_),
    .A1(_0298_),
    .B1(_0338_),
    .X(_0379_));
 sg13g2_o21ai_1 _1005_ (.B1(_0376_),
    .Y(_0380_),
    .A1(_0378_),
    .A2(_0379_));
 sg13g2_mux2_1 _1006_ (.A0(_0380_),
    .A1(net153),
    .S(_0263_),
    .X(_0039_));
 sg13g2_a21oi_1 _1007_ (.A1(_0296_),
    .A2(_0374_),
    .Y(_0381_),
    .B1(_0294_));
 sg13g2_nand3_1 _1008_ (.B(_0296_),
    .C(_0374_),
    .A(_0294_),
    .Y(_0382_));
 sg13g2_nand3b_1 _1009_ (.B(_0382_),
    .C(_0253_),
    .Y(_0383_),
    .A_N(_0381_));
 sg13g2_nor2_1 _1010_ (.A(_0295_),
    .B(_0378_),
    .Y(_0384_));
 sg13g2_nor2_1 _1011_ (.A(_0293_),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_a21o_1 _1012_ (.A2(_0384_),
    .A1(_0293_),
    .B1(_0338_),
    .X(_0386_));
 sg13g2_o21ai_1 _1013_ (.B1(_0383_),
    .Y(_0387_),
    .A1(_0385_),
    .A2(_0386_));
 sg13g2_mux2_1 _1014_ (.A0(_0387_),
    .A1(net104),
    .S(_0263_),
    .X(_0040_));
 sg13g2_nand3b_1 _1015_ (.B(net119),
    .C(_0261_),
    .Y(_0388_),
    .A_N(\ChiselTop.tappu.mem.tapeCounterReg[1] ));
 sg13g2_mux2_1 _1016_ (.A0(_0339_),
    .A1(net105),
    .S(_0388_),
    .X(_0041_));
 sg13g2_mux2_1 _1017_ (.A0(_0345_),
    .A1(net154),
    .S(_0388_),
    .X(_0042_));
 sg13g2_mux2_1 _1018_ (.A0(_0351_),
    .A1(net149),
    .S(_0388_),
    .X(_0043_));
 sg13g2_mux2_1 _1019_ (.A0(_0358_),
    .A1(net151),
    .S(_0388_),
    .X(_0044_));
 sg13g2_mux2_1 _1020_ (.A0(_0365_),
    .A1(net150),
    .S(_0388_),
    .X(_0045_));
 sg13g2_mux2_1 _1021_ (.A0(_0372_),
    .A1(net102),
    .S(_0388_),
    .X(_0046_));
 sg13g2_mux2_1 _1022_ (.A0(_0380_),
    .A1(net146),
    .S(_0388_),
    .X(_0047_));
 sg13g2_mux2_1 _1023_ (.A0(_0387_),
    .A1(net155),
    .S(_0388_),
    .X(_0048_));
 sg13g2_nor2b_1 _1024_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[0] ),
    .B_N(\ChiselTop.tappu.mem.tapeCounterReg[1] ),
    .Y(_0389_));
 sg13g2_nand2_2 _1025_ (.Y(_0390_),
    .A(_0261_),
    .B(_0389_));
 sg13g2_mux2_1 _1026_ (.A0(_0339_),
    .A1(net152),
    .S(_0390_),
    .X(_0049_));
 sg13g2_mux2_1 _1027_ (.A0(_0345_),
    .A1(net156),
    .S(_0390_),
    .X(_0050_));
 sg13g2_mux2_1 _1028_ (.A0(_0351_),
    .A1(net100),
    .S(_0390_),
    .X(_0051_));
 sg13g2_mux2_1 _1029_ (.A0(_0358_),
    .A1(net145),
    .S(_0390_),
    .X(_0052_));
 sg13g2_mux2_1 _1030_ (.A0(_0365_),
    .A1(net107),
    .S(_0390_),
    .X(_0053_));
 sg13g2_mux2_1 _1031_ (.A0(_0372_),
    .A1(net148),
    .S(_0390_),
    .X(_0054_));
 sg13g2_mux2_1 _1032_ (.A0(_0380_),
    .A1(net147),
    .S(_0390_),
    .X(_0055_));
 sg13g2_mux2_1 _1033_ (.A0(_0387_),
    .A1(net106),
    .S(_0390_),
    .X(_0056_));
 sg13g2_and2_1 _1034_ (.A(net141),
    .B(_0240_),
    .X(_0057_));
 sg13g2_and3_1 _1035_ (.X(_0391_),
    .A(_0181_),
    .B(_0245_),
    .C(_0257_));
 sg13g2_and2_1 _1036_ (.A(_0271_),
    .B(_0391_),
    .X(_0392_));
 sg13g2_o21ai_1 _1037_ (.B1(net143),
    .Y(_0393_),
    .A1(net158),
    .A2(net117));
 sg13g2_a21oi_1 _1038_ (.A1(_0138_),
    .A2(net117),
    .Y(_0058_),
    .B1(_0393_));
 sg13g2_o21ai_1 _1039_ (.B1(net143),
    .Y(_0394_),
    .A1(net161),
    .A2(net117));
 sg13g2_a21oi_1 _1040_ (.A1(_0143_),
    .A2(net117),
    .Y(_0059_),
    .B1(_0394_));
 sg13g2_o21ai_1 _1041_ (.B1(net143),
    .Y(_0395_),
    .A1(net162),
    .A2(net117));
 sg13g2_a21oi_1 _1042_ (.A1(_0154_),
    .A2(net117),
    .Y(_0060_),
    .B1(_0395_));
 sg13g2_o21ai_1 _1043_ (.B1(net143),
    .Y(_0396_),
    .A1(net167),
    .A2(net117));
 sg13g2_a21oi_1 _1044_ (.A1(_0148_),
    .A2(net117),
    .Y(_0061_),
    .B1(_0396_));
 sg13g2_o21ai_1 _1045_ (.B1(net143),
    .Y(_0397_),
    .A1(net159),
    .A2(net116));
 sg13g2_a21oi_1 _1046_ (.A1(_0126_),
    .A2(net116),
    .Y(_0062_),
    .B1(_0397_));
 sg13g2_o21ai_1 _1047_ (.B1(net142),
    .Y(_0398_),
    .A1(net163),
    .A2(net116));
 sg13g2_a21oi_1 _1048_ (.A1(_0114_),
    .A2(net116),
    .Y(_0063_),
    .B1(_0398_));
 sg13g2_o21ai_1 _1049_ (.B1(net142),
    .Y(_0399_),
    .A1(net165),
    .A2(net116));
 sg13g2_a21oi_1 _1050_ (.A1(_0131_),
    .A2(net116),
    .Y(_0064_),
    .B1(_0399_));
 sg13g2_o21ai_1 _1051_ (.B1(net142),
    .Y(_0400_),
    .A1(net166),
    .A2(net116));
 sg13g2_a21oi_1 _1052_ (.A1(_0120_),
    .A2(net116),
    .Y(_0065_),
    .B1(_0400_));
 sg13g2_o21ai_1 _1053_ (.B1(_0301_),
    .Y(_0401_),
    .A1(_0246_),
    .A2(_0257_));
 sg13g2_nor4_2 _1054_ (.A(_0251_),
    .B(_0270_),
    .C(_0391_),
    .Y(_0402_),
    .D(_0401_));
 sg13g2_nor3_2 _1055_ (.A(_0251_),
    .B(_0282_),
    .C(_0401_),
    .Y(_0403_));
 sg13g2_nor3_1 _1056_ (.A(net199),
    .B(net90),
    .C(net170),
    .Y(_0404_));
 sg13g2_nand3_1 _1057_ (.B(_0301_),
    .C(_0404_),
    .A(_0257_),
    .Y(_0405_));
 sg13g2_nor3_2 _1058_ (.A(net125),
    .B(_0251_),
    .C(_0313_),
    .Y(_0406_));
 sg13g2_nand3b_1 _1059_ (.B(_0250_),
    .C(_0312_),
    .Y(_0407_),
    .A_N(net124));
 sg13g2_nand2_1 _1060_ (.Y(_0408_),
    .A(_0405_),
    .B(_0407_));
 sg13g2_nor4_2 _1061_ (.A(net123),
    .B(_0402_),
    .C(_0403_),
    .Y(_0409_),
    .D(_0408_));
 sg13g2_or4_1 _1062_ (.A(net123),
    .B(net115),
    .C(_0403_),
    .D(_0408_),
    .X(_0410_));
 sg13g2_nand2_1 _1063_ (.Y(_0411_),
    .A(_0026_),
    .B(_0406_));
 sg13g2_nor2_1 _1064_ (.A(net119),
    .B(net115),
    .Y(_0412_));
 sg13g2_nor2_1 _1065_ (.A(_0026_),
    .B(_0406_),
    .Y(_0413_));
 sg13g2_nand3b_1 _1066_ (.B(_0236_),
    .C(_0025_),
    .Y(_0414_),
    .A_N(_0413_));
 sg13g2_a21oi_1 _1067_ (.A1(_0411_),
    .A2(_0412_),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_xnor2_1 _1068_ (.Y(_0416_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[5] ),
    .B(_0403_));
 sg13g2_a22oi_1 _1069_ (.Y(_0417_),
    .B1(_0415_),
    .B2(_0416_),
    .A2(_0403_),
    .A1(_0019_));
 sg13g2_nor2_1 _1070_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[7] ),
    .B(_0107_),
    .Y(_0418_));
 sg13g2_nor4_1 _1071_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[7] ),
    .B(_0107_),
    .C(_0234_),
    .D(_0417_),
    .Y(_0419_));
 sg13g2_and2_1 _1072_ (.A(_0416_),
    .B(_0418_),
    .X(_0420_));
 sg13g2_nor2_2 _1073_ (.A(_0405_),
    .B(_0419_),
    .Y(_0421_));
 sg13g2_and2_1 _1074_ (.A(net119),
    .B(net115),
    .X(_0422_));
 sg13g2_o21ai_1 _1075_ (.B1(_0421_),
    .Y(_0423_),
    .A1(_0412_),
    .A2(_0422_));
 sg13g2_nand2_1 _1076_ (.Y(_0424_),
    .A(_0102_),
    .B(net115));
 sg13g2_xnor2_1 _1077_ (.Y(_0425_),
    .A(_0102_),
    .B(net115));
 sg13g2_nor2_1 _1078_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[14] ),
    .B(\ChiselTop.tappu.mem.tapeCounterReg[13] ),
    .Y(_0426_));
 sg13g2_nand4_1 _1079_ (.B(\ChiselTop.tappu.mem.tapeCounterReg[10] ),
    .C(\ChiselTop.tappu.mem.tapeCounterReg[9] ),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[11] ),
    .Y(_0427_),
    .D(net120));
 sg13g2_nand2_1 _1080_ (.Y(_0428_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[6] ),
    .B(_0103_));
 sg13g2_nand2_1 _1081_ (.Y(_0429_),
    .A(net121),
    .B(_0406_));
 sg13g2_xor2_1 _1082_ (.B(_0407_),
    .A(net121),
    .X(_0430_));
 sg13g2_nand3b_1 _1083_ (.B(_0102_),
    .C(net115),
    .Y(_0431_),
    .A_N(_0430_));
 sg13g2_nand2_1 _1084_ (.Y(_0432_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[2] ),
    .B(_0104_));
 sg13g2_a21oi_2 _1085_ (.B1(_0432_),
    .Y(_0433_),
    .A2(_0431_),
    .A1(_0429_));
 sg13g2_nor2_1 _1086_ (.A(_0019_),
    .B(_0403_),
    .Y(_0434_));
 sg13g2_xnor2_1 _1087_ (.Y(_0435_),
    .A(_0019_),
    .B(_0403_));
 sg13g2_and2_1 _1088_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[4] ),
    .B(_0435_),
    .X(_0436_));
 sg13g2_a22oi_1 _1089_ (.Y(_0437_),
    .B1(_0433_),
    .B2(_0436_),
    .A2(_0403_),
    .A1(\ChiselTop.tappu.mem.tapeCounterReg[5] ));
 sg13g2_nor4_1 _1090_ (.A(_0089_),
    .B(_0427_),
    .C(_0428_),
    .D(_0437_),
    .Y(_0438_));
 sg13g2_a21oi_1 _1091_ (.A1(\ChiselTop.tappu.mem.tapeCounterReg[14] ),
    .A2(_0438_),
    .Y(_0439_),
    .B1(_0426_));
 sg13g2_nand3_1 _1092_ (.B(\ChiselTop.tappu.mem.tapeCounterReg[12] ),
    .C(_0105_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[13] ),
    .Y(_0440_));
 sg13g2_nor4_1 _1093_ (.A(_0427_),
    .B(_0428_),
    .C(_0437_),
    .D(_0440_),
    .Y(_0441_));
 sg13g2_xor2_1 _1094_ (.B(_0441_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[15] ),
    .X(_0442_));
 sg13g2_nor2b_1 _1095_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[13] ),
    .B_N(_0438_),
    .Y(_0443_));
 sg13g2_o21ai_1 _1096_ (.B1(_0106_),
    .Y(_0444_),
    .A1(_0428_),
    .A2(_0437_));
 sg13g2_nor3_1 _1097_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[10] ),
    .B(\ChiselTop.tappu.mem.tapeCounterReg[6] ),
    .C(_0103_),
    .Y(_0445_));
 sg13g2_a21o_1 _1098_ (.A2(_0445_),
    .A1(_0437_),
    .B1(_0106_),
    .X(_0446_));
 sg13g2_nor3_1 _1099_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[4] ),
    .B(_0433_),
    .C(_0435_),
    .Y(_0447_));
 sg13g2_a21o_1 _1100_ (.A2(_0436_),
    .A1(_0433_),
    .B1(_0447_),
    .X(_0448_));
 sg13g2_nand4_1 _1101_ (.B(_0020_),
    .C(_0429_),
    .A(_0095_),
    .Y(_0449_),
    .D(_0431_));
 sg13g2_nor2b_1 _1102_ (.A(_0433_),
    .B_N(_0449_),
    .Y(_0450_));
 sg13g2_nor2_1 _1103_ (.A(_0425_),
    .B(_0430_),
    .Y(_0451_));
 sg13g2_a21oi_1 _1104_ (.A1(net120),
    .A2(_0106_),
    .Y(_0452_),
    .B1(\ChiselTop.tappu.mem.tapeCounterReg[9] ));
 sg13g2_nand2_1 _1105_ (.Y(_0453_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[11] ),
    .B(_0021_));
 sg13g2_nand3_1 _1106_ (.B(net120),
    .C(_0453_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[9] ),
    .Y(_0454_));
 sg13g2_nor2_1 _1107_ (.A(_0091_),
    .B(_0022_),
    .Y(_0455_));
 sg13g2_a21oi_1 _1108_ (.A1(_0090_),
    .A2(_0021_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_a221oi_1 _1109_ (.B2(_0090_),
    .C1(_0456_),
    .B1(_0455_),
    .A1(\ChiselTop.tappu.mem.tapeCounterReg[10] ),
    .Y(_0457_),
    .A2(_0454_));
 sg13g2_o21ai_1 _1110_ (.B1(_0457_),
    .Y(_0458_),
    .A1(\ChiselTop.tappu.mem.tapeCounterReg[10] ),
    .A2(_0452_));
 sg13g2_nor3_1 _1111_ (.A(_0450_),
    .B(_0451_),
    .C(_0458_),
    .Y(_0459_));
 sg13g2_nand4_1 _1112_ (.B(_0446_),
    .C(_0448_),
    .A(_0444_),
    .Y(_0460_),
    .D(_0459_));
 sg13g2_nor4_1 _1113_ (.A(_0439_),
    .B(_0442_),
    .C(_0443_),
    .D(_0460_),
    .Y(_0461_));
 sg13g2_or4_1 _1114_ (.A(_0439_),
    .B(_0442_),
    .C(_0443_),
    .D(_0460_),
    .X(_0462_));
 sg13g2_nand3b_1 _1115_ (.B(_0461_),
    .C(_0405_),
    .Y(_0463_),
    .A_N(_0425_));
 sg13g2_nand3_1 _1116_ (.B(_0423_),
    .C(_0463_),
    .A(net126),
    .Y(_0464_));
 sg13g2_o21ai_1 _1117_ (.B1(_0464_),
    .Y(_0465_),
    .A1(net119),
    .A2(net126));
 sg13g2_o21ai_1 _1118_ (.B1(net141),
    .Y(_0466_),
    .A1(net192),
    .A2(net112));
 sg13g2_a21oi_1 _1119_ (.A1(net111),
    .A2(_0465_),
    .Y(_0066_),
    .B1(_0466_));
 sg13g2_xor2_1 _1120_ (.B(_0430_),
    .A(_0424_),
    .X(_0467_));
 sg13g2_o21ai_1 _1121_ (.B1(_0405_),
    .Y(_0468_),
    .A1(_0462_),
    .A2(_0467_));
 sg13g2_xor2_1 _1122_ (.B(_0407_),
    .A(_0026_),
    .X(_0469_));
 sg13g2_nand3_1 _1123_ (.B(net115),
    .C(_0469_),
    .A(net119),
    .Y(_0470_));
 sg13g2_a21oi_1 _1124_ (.A1(net119),
    .A2(net115),
    .Y(_0471_),
    .B1(_0469_));
 sg13g2_nand3b_1 _1125_ (.B(_0421_),
    .C(_0470_),
    .Y(_0472_),
    .A_N(_0471_));
 sg13g2_nand3_1 _1126_ (.B(_0468_),
    .C(_0472_),
    .A(net126),
    .Y(_0473_));
 sg13g2_or2_1 _1127_ (.X(_0474_),
    .B(_0389_),
    .A(_0262_));
 sg13g2_o21ai_1 _1128_ (.B1(_0473_),
    .Y(_0475_),
    .A1(net126),
    .A2(_0474_));
 sg13g2_o21ai_1 _1129_ (.B1(net141),
    .Y(_0476_),
    .A1(net121),
    .A2(net111));
 sg13g2_a21oi_1 _1130_ (.A1(net111),
    .A2(_0475_),
    .Y(_0067_),
    .B1(_0476_));
 sg13g2_nor2_2 _1131_ (.A(net126),
    .B(_0239_),
    .Y(_0477_));
 sg13g2_or2_2 _1132_ (.X(_0478_),
    .B(_0239_),
    .A(net126));
 sg13g2_nor2_1 _1133_ (.A(_0025_),
    .B(_0237_),
    .Y(_0479_));
 sg13g2_xor2_1 _1134_ (.B(_0237_),
    .A(_0025_),
    .X(_0480_));
 sg13g2_nor3_1 _1135_ (.A(_0025_),
    .B(_0413_),
    .C(_0471_),
    .Y(_0481_));
 sg13g2_o21ai_1 _1136_ (.B1(_0025_),
    .Y(_0482_),
    .A1(_0413_),
    .A2(_0471_));
 sg13g2_nor2b_1 _1137_ (.A(_0481_),
    .B_N(_0482_),
    .Y(_0483_));
 sg13g2_and2_1 _1138_ (.A(net126),
    .B(_0421_),
    .X(_0484_));
 sg13g2_a221oi_1 _1139_ (.B2(net109),
    .C1(net114),
    .B1(_0483_),
    .A1(_0477_),
    .Y(_0485_),
    .A2(_0480_));
 sg13g2_o21ai_1 _1140_ (.B1(net141),
    .Y(_0486_),
    .A1(net179),
    .A2(net112));
 sg13g2_nor2_1 _1141_ (.A(_0485_),
    .B(_0486_),
    .Y(_0068_));
 sg13g2_xnor2_1 _1142_ (.Y(_0487_),
    .A(_0020_),
    .B(_0479_));
 sg13g2_a21oi_1 _1143_ (.A1(_0095_),
    .A2(_0482_),
    .Y(_0488_),
    .B1(\ChiselTop.tappu.mem.tapeCounterReg[3] ));
 sg13g2_nand3_1 _1144_ (.B(_0095_),
    .C(_0482_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[3] ),
    .Y(_0489_));
 sg13g2_nor2b_1 _1145_ (.A(_0488_),
    .B_N(_0489_),
    .Y(_0490_));
 sg13g2_a221oi_1 _1146_ (.B2(net108),
    .C1(net113),
    .B1(_0490_),
    .A1(_0477_),
    .Y(_0491_),
    .A2(_0487_));
 sg13g2_o21ai_1 _1147_ (.B1(net140),
    .Y(_0492_),
    .A1(net174),
    .A2(net110));
 sg13g2_nor2_1 _1148_ (.A(_0491_),
    .B(_0492_),
    .Y(_0069_));
 sg13g2_or3_2 _1149_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[4] ),
    .B(_0104_),
    .C(_0488_),
    .X(_0493_));
 sg13g2_o21ai_1 _1150_ (.B1(\ChiselTop.tappu.mem.tapeCounterReg[4] ),
    .Y(_0494_),
    .A1(_0104_),
    .A2(_0488_));
 sg13g2_nand2_1 _1151_ (.Y(_0495_),
    .A(_0493_),
    .B(_0494_));
 sg13g2_nand2_1 _1152_ (.Y(_0496_),
    .A(_0421_),
    .B(_0495_));
 sg13g2_nand4_1 _1153_ (.B(\ChiselTop.tappu.mem.tapeCounterReg[2] ),
    .C(net121),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[3] ),
    .Y(_0497_),
    .D(\ChiselTop.tappu.mem.tapeCounterReg[0] ));
 sg13g2_nor2_1 _1154_ (.A(_0094_),
    .B(_0497_),
    .Y(_0498_));
 sg13g2_xnor2_1 _1155_ (.Y(_0499_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[4] ),
    .B(_0497_));
 sg13g2_o21ai_1 _1156_ (.B1(net111),
    .Y(_0500_),
    .A1(net125),
    .A2(_0499_));
 sg13g2_a21oi_1 _1157_ (.A1(net125),
    .A2(_0496_),
    .Y(_0501_),
    .B1(_0500_));
 sg13g2_a21oi_1 _1158_ (.A1(net187),
    .A2(net113),
    .Y(_0502_),
    .B1(_0501_));
 sg13g2_nor2b_1 _1159_ (.A(_0502_),
    .B_N(net140),
    .Y(_0070_));
 sg13g2_xnor2_1 _1160_ (.Y(_0503_),
    .A(_0019_),
    .B(_0498_));
 sg13g2_xor2_1 _1161_ (.B(_0493_),
    .A(_0416_),
    .X(_0504_));
 sg13g2_a221oi_1 _1162_ (.B2(net109),
    .C1(net114),
    .B1(_0504_),
    .A1(_0477_),
    .Y(_0505_),
    .A2(_0503_));
 sg13g2_o21ai_1 _1163_ (.B1(net141),
    .Y(_0506_),
    .A1(net171),
    .A2(net111));
 sg13g2_nor2_1 _1164_ (.A(_0505_),
    .B(_0506_),
    .Y(_0071_));
 sg13g2_and2_1 _1165_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[5] ),
    .B(_0498_),
    .X(_0507_));
 sg13g2_inv_1 _1166_ (.Y(_0508_),
    .A(_0507_));
 sg13g2_nand2_1 _1167_ (.Y(_0509_),
    .A(_0107_),
    .B(_0507_));
 sg13g2_a21oi_1 _1168_ (.A1(net181),
    .A2(_0508_),
    .Y(_0510_),
    .B1(_0478_));
 sg13g2_a21oi_1 _1169_ (.A1(_0509_),
    .A2(_0510_),
    .Y(_0511_),
    .B1(net114));
 sg13g2_a21oi_1 _1170_ (.A1(_0416_),
    .A2(_0493_),
    .Y(_0512_),
    .B1(_0434_));
 sg13g2_nand2_1 _1171_ (.Y(_0513_),
    .A(_0107_),
    .B(_0512_));
 sg13g2_nor2_1 _1172_ (.A(_0107_),
    .B(_0512_),
    .Y(_0514_));
 sg13g2_nand3b_1 _1173_ (.B(net109),
    .C(_0513_),
    .Y(_0515_),
    .A_N(_0514_));
 sg13g2_o21ai_1 _1174_ (.B1(net144),
    .Y(_0516_),
    .A1(\ChiselTop.tappu.mem.tapeCounterReg[6] ),
    .A2(net111));
 sg13g2_a21oi_1 _1175_ (.A1(_0511_),
    .A2(_0515_),
    .Y(_0072_),
    .B1(_0516_));
 sg13g2_nor2_1 _1176_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[6] ),
    .B(_0514_),
    .Y(_0517_));
 sg13g2_xnor2_1 _1177_ (.Y(_0518_),
    .A(_0093_),
    .B(_0517_));
 sg13g2_nand3_1 _1178_ (.B(_0107_),
    .C(_0507_),
    .A(_0103_),
    .Y(_0519_));
 sg13g2_a21oi_1 _1179_ (.A1(_0018_),
    .A2(_0509_),
    .Y(_0520_),
    .B1(_0478_));
 sg13g2_a221oi_1 _1180_ (.B2(_0520_),
    .C1(net114),
    .B1(_0519_),
    .A1(net109),
    .Y(_0521_),
    .A2(_0518_));
 sg13g2_o21ai_1 _1181_ (.B1(net144),
    .Y(_0522_),
    .A1(net190),
    .A2(net111));
 sg13g2_nor2_1 _1182_ (.A(_0521_),
    .B(_0522_),
    .Y(_0073_));
 sg13g2_nand3_1 _1183_ (.B(\ChiselTop.tappu.mem.tapeCounterReg[6] ),
    .C(_0507_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[7] ),
    .Y(_0523_));
 sg13g2_nor2_1 _1184_ (.A(_0092_),
    .B(_0523_),
    .Y(_0524_));
 sg13g2_xnor2_1 _1185_ (.Y(_0525_),
    .A(_0092_),
    .B(_0523_));
 sg13g2_o21ai_1 _1186_ (.B1(net111),
    .Y(_0526_),
    .A1(net125),
    .A2(_0525_));
 sg13g2_a22oi_1 _1187_ (.Y(_0527_),
    .B1(_0418_),
    .B2(_0434_),
    .A2(\ChiselTop.tappu.mem.tapeCounterReg[6] ),
    .A1(_0093_));
 sg13g2_nand2_1 _1188_ (.Y(_0528_),
    .A(_0018_),
    .B(_0527_));
 sg13g2_a21o_2 _1189_ (.A2(_0493_),
    .A1(_0420_),
    .B1(_0528_),
    .X(_0529_));
 sg13g2_xnor2_1 _1190_ (.Y(_0530_),
    .A(_0106_),
    .B(_0529_));
 sg13g2_a21oi_1 _1191_ (.A1(net109),
    .A2(_0530_),
    .Y(_0531_),
    .B1(_0526_));
 sg13g2_o21ai_1 _1192_ (.B1(net141),
    .Y(_0532_),
    .A1(net120),
    .A2(net110));
 sg13g2_nor2_1 _1193_ (.A(_0531_),
    .B(_0532_),
    .Y(_0074_));
 sg13g2_xnor2_1 _1194_ (.Y(_0533_),
    .A(net196),
    .B(_0524_));
 sg13g2_nor2_1 _1195_ (.A(net120),
    .B(_0529_),
    .Y(_0534_));
 sg13g2_xnor2_1 _1196_ (.Y(_0535_),
    .A(net196),
    .B(_0534_));
 sg13g2_a221oi_1 _1197_ (.B2(net108),
    .C1(net114),
    .B1(_0535_),
    .A1(_0477_),
    .Y(_0536_),
    .A2(_0533_));
 sg13g2_o21ai_1 _1198_ (.B1(net139),
    .Y(_0537_),
    .A1(\ChiselTop.tappu.mem.tapeCounterReg[9] ),
    .A2(net110));
 sg13g2_nor2_1 _1199_ (.A(_0536_),
    .B(_0537_),
    .Y(_0075_));
 sg13g2_nor3_2 _1200_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[9] ),
    .B(net120),
    .C(_0529_),
    .Y(_0538_));
 sg13g2_xnor2_1 _1201_ (.Y(_0539_),
    .A(_0022_),
    .B(_0538_));
 sg13g2_nand2_1 _1202_ (.Y(_0540_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[9] ),
    .B(_0524_));
 sg13g2_nor2_1 _1203_ (.A(_0022_),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_inv_1 _1204_ (.Y(_0542_),
    .A(_0541_));
 sg13g2_a21oi_1 _1205_ (.A1(_0022_),
    .A2(_0540_),
    .Y(_0543_),
    .B1(_0478_));
 sg13g2_a221oi_1 _1206_ (.B2(_0543_),
    .C1(net113),
    .B1(_0542_),
    .A1(net108),
    .Y(_0544_),
    .A2(_0539_));
 sg13g2_o21ai_1 _1207_ (.B1(net139),
    .Y(_0545_),
    .A1(net200),
    .A2(net110));
 sg13g2_nor2_1 _1208_ (.A(_0544_),
    .B(_0545_),
    .Y(_0076_));
 sg13g2_a21oi_1 _1209_ (.A1(_0009_),
    .A2(_0542_),
    .Y(_0546_),
    .B1(_0478_));
 sg13g2_nand2b_1 _1210_ (.Y(_0547_),
    .B(_0541_),
    .A_N(_0009_));
 sg13g2_nor4_2 _1211_ (.A(\ChiselTop.tappu.mem.tapeCounterReg[10] ),
    .B(\ChiselTop.tappu.mem.tapeCounterReg[9] ),
    .C(net120),
    .Y(_0548_),
    .D(_0529_));
 sg13g2_xnor2_1 _1212_ (.Y(_0549_),
    .A(_0009_),
    .B(_0548_));
 sg13g2_a221oi_1 _1213_ (.B2(net108),
    .C1(net113),
    .B1(_0549_),
    .A1(_0546_),
    .Y(_0550_),
    .A2(_0547_));
 sg13g2_o21ai_1 _1214_ (.B1(net139),
    .Y(_0551_),
    .A1(net185),
    .A2(net110));
 sg13g2_nor2_1 _1215_ (.A(_0550_),
    .B(_0551_),
    .Y(_0077_));
 sg13g2_and2_1 _1216_ (.A(_0090_),
    .B(_0548_),
    .X(_0552_));
 sg13g2_xnor2_1 _1217_ (.Y(_0553_),
    .A(_0021_),
    .B(_0552_));
 sg13g2_nor3_2 _1218_ (.A(_0090_),
    .B(_0091_),
    .C(_0540_),
    .Y(_0554_));
 sg13g2_nor2b_1 _1219_ (.A(_0554_),
    .B_N(_0021_),
    .Y(_0555_));
 sg13g2_nand2b_1 _1220_ (.Y(_0556_),
    .B(_0554_),
    .A_N(_0021_));
 sg13g2_nor2_1 _1221_ (.A(_0478_),
    .B(_0555_),
    .Y(_0557_));
 sg13g2_a221oi_1 _1222_ (.B2(_0557_),
    .C1(net113),
    .B1(_0556_),
    .A1(net108),
    .Y(_0558_),
    .A2(_0553_));
 sg13g2_o21ai_1 _1223_ (.B1(net139),
    .Y(_0559_),
    .A1(net183),
    .A2(net110));
 sg13g2_nor2_1 _1224_ (.A(_0558_),
    .B(_0559_),
    .Y(_0078_));
 sg13g2_nand3_1 _1225_ (.B(_0090_),
    .C(_0548_),
    .A(_0089_),
    .Y(_0560_));
 sg13g2_xor2_1 _1226_ (.B(_0560_),
    .A(_0010_),
    .X(_0561_));
 sg13g2_xor2_1 _1227_ (.B(_0556_),
    .A(_0010_),
    .X(_0562_));
 sg13g2_a221oi_1 _1228_ (.B2(_0477_),
    .C1(net113),
    .B1(_0562_),
    .A1(net108),
    .Y(_0563_),
    .A2(_0561_));
 sg13g2_o21ai_1 _1229_ (.B1(net139),
    .Y(_0564_),
    .A1(net188),
    .A2(net110));
 sg13g2_nor2_1 _1230_ (.A(_0563_),
    .B(_0564_),
    .Y(_0079_));
 sg13g2_nand2_1 _1231_ (.Y(_0565_),
    .A(_0232_),
    .B(_0538_));
 sg13g2_xnor2_1 _1232_ (.Y(_0566_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[14] ),
    .B(_0565_));
 sg13g2_nand3_1 _1233_ (.B(\ChiselTop.tappu.mem.tapeCounterReg[12] ),
    .C(_0554_),
    .A(\ChiselTop.tappu.mem.tapeCounterReg[13] ),
    .Y(_0567_));
 sg13g2_nand2b_1 _1234_ (.Y(_0568_),
    .B(_0105_),
    .A_N(_0567_));
 sg13g2_a21oi_1 _1235_ (.A1(_0017_),
    .A2(_0567_),
    .Y(_0569_),
    .B1(_0478_));
 sg13g2_a221oi_1 _1236_ (.B2(_0569_),
    .C1(net113),
    .B1(_0568_),
    .A1(net108),
    .Y(_0570_),
    .A2(_0566_));
 sg13g2_o21ai_1 _1237_ (.B1(net139),
    .Y(_0571_),
    .A1(net176),
    .A2(net112));
 sg13g2_nor2_1 _1238_ (.A(_0570_),
    .B(_0571_),
    .Y(_0080_));
 sg13g2_o21ai_1 _1239_ (.B1(_0011_),
    .Y(_0572_),
    .A1(_0105_),
    .A2(_0565_));
 sg13g2_or3_1 _1240_ (.A(_0105_),
    .B(_0011_),
    .C(_0565_),
    .X(_0573_));
 sg13g2_nand3_1 _1241_ (.B(_0572_),
    .C(_0573_),
    .A(net108),
    .Y(_0574_));
 sg13g2_xor2_1 _1242_ (.B(_0568_),
    .A(_0011_),
    .X(_0575_));
 sg13g2_a21oi_1 _1243_ (.A1(_0477_),
    .A2(_0575_),
    .Y(_0576_),
    .B1(net113));
 sg13g2_o21ai_1 _1244_ (.B1(net139),
    .Y(_0577_),
    .A1(net168),
    .A2(net110));
 sg13g2_a21oi_1 _1245_ (.A1(_0574_),
    .A2(_0576_),
    .Y(_0081_),
    .B1(_0577_));
 sg13g2_nand3_1 _1246_ (.B(_0171_),
    .C(_0404_),
    .A(net143),
    .Y(_0578_));
 sg13g2_a21oi_2 _1247_ (.B1(_0578_),
    .Y(_0085_),
    .A2(_0301_),
    .A1(_0246_));
 sg13g2_nor2b_1 _1248_ (.A(_0270_),
    .B_N(_0085_),
    .Y(_0084_));
 sg13g2_a21oi_1 _1249_ (.A1(_0096_),
    .A2(net127),
    .Y(_0082_),
    .B1(_0193_));
 sg13g2_mux2_1 _1250_ (.A0(net91),
    .A1(net121),
    .S(net126),
    .X(_0083_));
 sg13g2_nor2b_1 _1251_ (.A(_0270_),
    .B_N(_0085_),
    .Y(_0086_));
 sg13g2_dfrbp_1 _1252_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net24),
    .D(_0028_),
    .Q_N(_0623_),
    .Q(\ChiselTop.tappu.mem._GEN_198[1] ));
 sg13g2_dfrbp_1 _1253_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net68),
    .D(_0029_),
    .Q_N(_0622_),
    .Q(\ChiselTop.tappu.mem._GEN_198[2] ));
 sg13g2_dfrbp_1 _1254_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net66),
    .D(_0030_),
    .Q_N(_0621_),
    .Q(\ChiselTop.tappu.mem._GEN_198[3] ));
 sg13g2_dfrbp_1 _1255_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net64),
    .D(_0031_),
    .Q_N(_0620_),
    .Q(\ChiselTop.tappu.mem._GEN_198[4] ));
 sg13g2_dfrbp_1 _1256_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net25),
    .D(_0032_),
    .Q_N(_0013_),
    .Q(\ChiselTop.tappu.mem._GEN_198[5] ));
 sg13g2_dfrbp_1 _1257_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net82),
    .D(_0007_),
    .Q_N(_0624_),
    .Q(_0000_));
 sg13g2_dfrbp_1 _1258_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net62),
    .D(net92),
    .Q_N(_0619_),
    .Q(_0001_));
 sg13g2_dfrbp_1 _1259_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net60),
    .D(_0033_),
    .Q_N(_0618_),
    .Q(\ChiselTop.tappu.mem.tape[1][0] ));
 sg13g2_dfrbp_1 _1260_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net59),
    .D(_0034_),
    .Q_N(_0617_),
    .Q(\ChiselTop.tappu.mem.tape[1][1] ));
 sg13g2_dfrbp_1 _1261_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net58),
    .D(_0035_),
    .Q_N(_0616_),
    .Q(\ChiselTop.tappu.mem.tape[1][2] ));
 sg13g2_dfrbp_1 _1262_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net57),
    .D(_0036_),
    .Q_N(_0615_),
    .Q(\ChiselTop.tappu.mem.tape[1][3] ));
 sg13g2_dfrbp_1 _1263_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net56),
    .D(_0037_),
    .Q_N(_0614_),
    .Q(\ChiselTop.tappu.mem.tape[1][4] ));
 sg13g2_dfrbp_1 _1264_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net55),
    .D(_0038_),
    .Q_N(_0613_),
    .Q(\ChiselTop.tappu.mem.tape[1][5] ));
 sg13g2_dfrbp_1 _1265_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net54),
    .D(_0039_),
    .Q_N(_0612_),
    .Q(\ChiselTop.tappu.mem.tape[1][6] ));
 sg13g2_dfrbp_1 _1266_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net53),
    .D(_0040_),
    .Q_N(_0611_),
    .Q(\ChiselTop.tappu.mem.tape[1][7] ));
 sg13g2_dfrbp_1 _1267_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net52),
    .D(_0041_),
    .Q_N(_0610_),
    .Q(\ChiselTop.tappu.mem.tape[0][0] ));
 sg13g2_dfrbp_1 _1268_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net51),
    .D(_0042_),
    .Q_N(_0609_),
    .Q(\ChiselTop.tappu.mem.tape[0][1] ));
 sg13g2_dfrbp_1 _1269_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net50),
    .D(_0043_),
    .Q_N(_0608_),
    .Q(\ChiselTop.tappu.mem.tape[0][2] ));
 sg13g2_dfrbp_1 _1270_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net49),
    .D(_0044_),
    .Q_N(_0607_),
    .Q(\ChiselTop.tappu.mem.tape[0][3] ));
 sg13g2_dfrbp_1 _1271_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net48),
    .D(_0045_),
    .Q_N(_0606_),
    .Q(\ChiselTop.tappu.mem.tape[0][4] ));
 sg13g2_dfrbp_1 _1272_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net47),
    .D(_0046_),
    .Q_N(_0605_),
    .Q(\ChiselTop.tappu.mem.tape[0][5] ));
 sg13g2_dfrbp_1 _1273_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net46),
    .D(_0047_),
    .Q_N(_0604_),
    .Q(\ChiselTop.tappu.mem.tape[0][6] ));
 sg13g2_dfrbp_1 _1274_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net45),
    .D(_0048_),
    .Q_N(_0603_),
    .Q(\ChiselTop.tappu.mem.tape[0][7] ));
 sg13g2_dfrbp_1 _1275_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net44),
    .D(_0049_),
    .Q_N(_0602_),
    .Q(\ChiselTop.tappu.mem.tape[2][0] ));
 sg13g2_dfrbp_1 _1276_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net43),
    .D(_0050_),
    .Q_N(_0601_),
    .Q(\ChiselTop.tappu.mem.tape[2][1] ));
 sg13g2_dfrbp_1 _1277_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net42),
    .D(_0051_),
    .Q_N(_0600_),
    .Q(\ChiselTop.tappu.mem.tape[2][2] ));
 sg13g2_dfrbp_1 _1278_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net41),
    .D(_0052_),
    .Q_N(_0599_),
    .Q(\ChiselTop.tappu.mem.tape[2][3] ));
 sg13g2_dfrbp_1 _1279_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net40),
    .D(_0053_),
    .Q_N(_0598_),
    .Q(\ChiselTop.tappu.mem.tape[2][4] ));
 sg13g2_dfrbp_1 _1280_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net39),
    .D(_0054_),
    .Q_N(_0597_),
    .Q(\ChiselTop.tappu.mem.tape[2][5] ));
 sg13g2_dfrbp_1 _1281_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net38),
    .D(_0055_),
    .Q_N(_0596_),
    .Q(\ChiselTop.tappu.mem.tape[2][6] ));
 sg13g2_dfrbp_1 _1282_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net37),
    .D(_0056_),
    .Q_N(_0595_),
    .Q(\ChiselTop.tappu.mem.tape[2][7] ));
 sg13g2_dfrbp_1 _1283_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net36),
    .D(_0057_),
    .Q_N(_0012_),
    .Q(\ChiselTop.tappu.mem.state ));
 sg13g2_dfrbp_1 _1284_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net35),
    .D(_0058_),
    .Q_N(_0594_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _1285_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net33),
    .D(_0059_),
    .Q_N(_0593_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _1286_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net31),
    .D(_0060_),
    .Q_N(_0592_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _1287_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net29),
    .D(_0061_),
    .Q_N(_0591_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _1288_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net27),
    .D(net160),
    .Q_N(_0590_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1289_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net23),
    .D(net164),
    .Q_N(_0589_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1290_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net21),
    .D(_0064_),
    .Q_N(_0588_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1291_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net19),
    .D(_0065_),
    .Q_N(_0587_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _1292_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net80),
    .D(_0066_),
    .Q_N(_0016_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[0] ));
 sg13g2_dfrbp_1 _1293_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net78),
    .D(_0067_),
    .Q_N(_0026_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[1] ));
 sg13g2_dfrbp_1 _1294_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net76),
    .D(net180),
    .Q_N(_0025_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[2] ));
 sg13g2_dfrbp_1 _1295_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net74),
    .D(net175),
    .Q_N(_0020_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[3] ));
 sg13g2_dfrbp_1 _1296_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net72),
    .D(_0070_),
    .Q_N(_0586_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[4] ));
 sg13g2_dfrbp_1 _1297_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net70),
    .D(_0071_),
    .Q_N(_0019_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[5] ));
 sg13g2_dfrbp_1 _1298_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net67),
    .D(net182),
    .Q_N(_0024_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[6] ));
 sg13g2_dfrbp_1 _1299_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net63),
    .D(net191),
    .Q_N(_0018_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[7] ));
 sg13g2_dfrbp_1 _1300_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net34),
    .D(net203),
    .Q_N(_0023_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[8] ));
 sg13g2_dfrbp_1 _1301_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net30),
    .D(net197),
    .Q_N(_0027_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[9] ));
 sg13g2_dfrbp_1 _1302_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net26),
    .D(net201),
    .Q_N(_0022_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[10] ));
 sg13g2_dfrbp_1 _1303_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net20),
    .D(net186),
    .Q_N(_0009_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[11] ));
 sg13g2_dfrbp_1 _1304_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net79),
    .D(net184),
    .Q_N(_0021_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[12] ));
 sg13g2_dfrbp_1 _1305_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net75),
    .D(net189),
    .Q_N(_0010_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[13] ));
 sg13g2_dfrbp_1 _1306_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net71),
    .D(net177),
    .Q_N(_0017_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[14] ));
 sg13g2_dfrbp_1 _1307_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net65),
    .D(net169),
    .Q_N(_0011_),
    .Q(\ChiselTop.tappu.mem.tapeCounterReg[15] ));
 sg13g2_dfrbp_1 _1308_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net32),
    .D(net95),
    .Q_N(_0585_),
    .Q(\ChiselTop.tappu.mem.tape_readData_addr[0] ));
 sg13g2_dfrbp_1 _1309_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net28),
    .D(_0083_),
    .Q_N(_0584_),
    .Q(\ChiselTop.tappu.mem.tape_readData_addr[1] ));
 sg13g2_dfrbp_1 _1310_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net22),
    .D(_0084_),
    .Q_N(_0583_),
    .Q(\ChiselTop.tappu.instrStepReg[0] ));
 sg13g2_dfrbp_1 _1311_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net81),
    .D(_0085_),
    .Q_N(_0582_),
    .Q(\ChiselTop.tappu.instrStepReg[1] ));
 sg13g2_dfrbp_1 _1312_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net77),
    .D(_0086_),
    .Q_N(_0581_),
    .Q(\ChiselTop.tappu.instrStepReg[4] ));
 sg13g2_dfrbp_1 _1313_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net73),
    .D(net18),
    .Q_N(_0580_),
    .Q(\ChiselTop.tappu.instrStepReg[5] ));
 sg13g2_dfrbp_1 _1314_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net83),
    .D(net17),
    .Q_N(_0625_),
    .Q(\ChiselTop.tappu.instrStepReg[2] ));
 sg13g2_dfrbp_1 _1315_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net84),
    .D(net89),
    .Q_N(_0015_),
    .Q(\ChiselTop.tappu.cpuState[0] ));
 sg13g2_dfrbp_1 _1316_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net85),
    .D(_0002_),
    .Q_N(_0626_),
    .Q(\ChiselTop.tappu.cpuState[1] ));
 sg13g2_dfrbp_1 _1317_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net86),
    .D(_0003_),
    .Q_N(_0014_),
    .Q(\ChiselTop.tappu.cpuState[2] ));
 sg13g2_dfrbp_1 _1318_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net61),
    .D(_0004_),
    .Q_N(_0627_),
    .Q(\ChiselTop.tappu.cpuState[3] ));
 sg13g2_dfrbp_1 _1319_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net69),
    .D(_0006_),
    .Q_N(_0579_),
    .Q(\ChiselTop.tappu.cpuState[5] ));
 sg13g2_tiehi _1303__20 (.L_HI(net20));
 sg13g2_tiehi _1290__21 (.L_HI(net21));
 sg13g2_tiehi _1310__22 (.L_HI(net22));
 sg13g2_tiehi _1289__23 (.L_HI(net23));
 sg13g2_tiehi _1252__24 (.L_HI(net24));
 sg13g2_tiehi _1256__25 (.L_HI(net25));
 sg13g2_tiehi _1302__26 (.L_HI(net26));
 sg13g2_tiehi _1288__27 (.L_HI(net27));
 sg13g2_tiehi _1309__28 (.L_HI(net28));
 sg13g2_tiehi _1287__29 (.L_HI(net29));
 sg13g2_tiehi _1301__30 (.L_HI(net30));
 sg13g2_tiehi _1286__31 (.L_HI(net31));
 sg13g2_tiehi _1308__32 (.L_HI(net32));
 sg13g2_tiehi _1285__33 (.L_HI(net33));
 sg13g2_tiehi _1300__34 (.L_HI(net34));
 sg13g2_tiehi _1284__35 (.L_HI(net35));
 sg13g2_tiehi _1283__36 (.L_HI(net36));
 sg13g2_tiehi _1282__37 (.L_HI(net37));
 sg13g2_tiehi _1281__38 (.L_HI(net38));
 sg13g2_tiehi _1280__39 (.L_HI(net39));
 sg13g2_tiehi _1279__40 (.L_HI(net40));
 sg13g2_tiehi _1278__41 (.L_HI(net41));
 sg13g2_tiehi _1277__42 (.L_HI(net42));
 sg13g2_tiehi _1276__43 (.L_HI(net43));
 sg13g2_tiehi _1275__44 (.L_HI(net44));
 sg13g2_tiehi _1274__45 (.L_HI(net45));
 sg13g2_tiehi _1273__46 (.L_HI(net46));
 sg13g2_tiehi _1272__47 (.L_HI(net47));
 sg13g2_tiehi _1271__48 (.L_HI(net48));
 sg13g2_tiehi _1270__49 (.L_HI(net49));
 sg13g2_tiehi _1269__50 (.L_HI(net50));
 sg13g2_tiehi _1268__51 (.L_HI(net51));
 sg13g2_tiehi _1267__52 (.L_HI(net52));
 sg13g2_tiehi _1266__53 (.L_HI(net53));
 sg13g2_tiehi _1265__54 (.L_HI(net54));
 sg13g2_tiehi _1264__55 (.L_HI(net55));
 sg13g2_tiehi _1263__56 (.L_HI(net56));
 sg13g2_tiehi _1262__57 (.L_HI(net57));
 sg13g2_tiehi _1261__58 (.L_HI(net58));
 sg13g2_tiehi _1260__59 (.L_HI(net59));
 sg13g2_tiehi _1259__60 (.L_HI(net60));
 sg13g2_tiehi _1318__61 (.L_HI(net61));
 sg13g2_tiehi _1258__62 (.L_HI(net62));
 sg13g2_tiehi _1299__63 (.L_HI(net63));
 sg13g2_tiehi _1255__64 (.L_HI(net64));
 sg13g2_tiehi _1307__65 (.L_HI(net65));
 sg13g2_tiehi _1254__66 (.L_HI(net66));
 sg13g2_tiehi _1298__67 (.L_HI(net67));
 sg13g2_tiehi _1253__68 (.L_HI(net68));
 sg13g2_tiehi _1319__69 (.L_HI(net69));
 sg13g2_tiehi _1297__70 (.L_HI(net70));
 sg13g2_tiehi _1306__71 (.L_HI(net71));
 sg13g2_tiehi _1296__72 (.L_HI(net72));
 sg13g2_tiehi _1313__73 (.L_HI(net73));
 sg13g2_tiehi _1295__74 (.L_HI(net74));
 sg13g2_tiehi _1305__75 (.L_HI(net75));
 sg13g2_tiehi _1294__76 (.L_HI(net76));
 sg13g2_tiehi _1312__77 (.L_HI(net77));
 sg13g2_tiehi _1293__78 (.L_HI(net78));
 sg13g2_tiehi _1304__79 (.L_HI(net79));
 sg13g2_tiehi _1292__80 (.L_HI(net80));
 sg13g2_tiehi _1311__81 (.L_HI(net81));
 sg13g2_tiehi _1257__82 (.L_HI(net82));
 sg13g2_tiehi _1314__83 (.L_HI(net83));
 sg13g2_tiehi _1315__84 (.L_HI(net84));
 sg13g2_tiehi _1316__85 (.L_HI(net85));
 sg13g2_tiehi _1317__86 (.L_HI(net86));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_tappu_tobias1012_2 (.L_LO(net2));
 sg13g2_tielo tt_um_tappu_tobias1012_3 (.L_LO(net3));
 sg13g2_tielo tt_um_tappu_tobias1012_4 (.L_LO(net4));
 sg13g2_tielo tt_um_tappu_tobias1012_5 (.L_LO(net5));
 sg13g2_tielo tt_um_tappu_tobias1012_6 (.L_LO(net6));
 sg13g2_tielo tt_um_tappu_tobias1012_7 (.L_LO(net7));
 sg13g2_tielo tt_um_tappu_tobias1012_8 (.L_LO(net8));
 sg13g2_tielo tt_um_tappu_tobias1012_9 (.L_LO(net9));
 sg13g2_tielo tt_um_tappu_tobias1012_10 (.L_LO(net10));
 sg13g2_tielo tt_um_tappu_tobias1012_11 (.L_LO(net11));
 sg13g2_tielo tt_um_tappu_tobias1012_12 (.L_LO(net12));
 sg13g2_tielo tt_um_tappu_tobias1012_13 (.L_LO(net13));
 sg13g2_tielo tt_um_tappu_tobias1012_14 (.L_LO(net14));
 sg13g2_tielo tt_um_tappu_tobias1012_15 (.L_LO(net15));
 sg13g2_tielo tt_um_tappu_tobias1012_16 (.L_LO(net16));
 sg13g2_tielo _1314__17 (.L_LO(net17));
 sg13g2_tielo _1313__18 (.L_LO(net18));
 sg13g2_tiehi _1291__19 (.L_HI(net19));
 sg13g2_buf_2 fanout108 (.A(_0484_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0484_),
    .X(net109));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(net112));
 sg13g2_buf_2 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0410_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0409_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0409_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0402_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0392_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0392_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0291_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0096_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(\ChiselTop.tappu.mem.tapeCounterReg[8] ),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(net93),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(net123),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(net198),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(net128),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(net128),
    .X(net126));
 sg13g2_buf_1 fanout127 (.A(net128),
    .X(net127));
 sg13g2_buf_1 fanout128 (.A(\ChiselTop.tappu.mem.state ),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_0001_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0001_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_0000_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_0000_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_0013_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(net204),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_1 fanout137 (.A(net194),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net195),
    .X(net138));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net141));
 sg13g2_buf_2 fanout140 (.A(net141),
    .X(net140));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net144));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net144));
 sg13g2_buf_2 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(rst_n),
    .X(net144));
 sg13g2_tielo tt_um_tappu_tobias1012_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ChiselTop.tappu.cpuState[5] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ChiselTop.tappu.cpuState[1] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0005_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold4 (.A(\ChiselTop.tappu.cpuState[3] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold5 (.A(\ChiselTop.tappu.mem.tape_readData_addr[1] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0008_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold7 (.A(\ChiselTop.tappu.mem.tapeCounterReg[1] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold8 (.A(\ChiselTop.tappu.mem.tape_readData_addr[0] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0082_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold10 (.A(\ChiselTop.tappu.cpuState[2] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold11 (.A(\ChiselTop.tappu.mem.tape[1][5] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold12 (.A(\ChiselTop.tappu.mem.tape[1][4] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold13 (.A(\ChiselTop.tappu.mem.tape[1][0] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold14 (.A(\ChiselTop.tappu.mem.tape[2][2] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold15 (.A(\ChiselTop.tappu.mem.tape[1][2] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold16 (.A(\ChiselTop.tappu.mem.tape[0][5] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold17 (.A(\ChiselTop.tappu.mem.tape[1][1] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold18 (.A(\ChiselTop.tappu.mem.tape[1][7] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold19 (.A(\ChiselTop.tappu.mem.tape[0][0] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold20 (.A(\ChiselTop.tappu.mem.tape[2][7] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold21 (.A(\ChiselTop.tappu.mem.tape[2][4] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold22 (.A(\ChiselTop.tappu.mem.tape[2][3] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold23 (.A(\ChiselTop.tappu.mem.tape[0][6] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold24 (.A(\ChiselTop.tappu.mem.tape[2][6] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold25 (.A(\ChiselTop.tappu.mem.tape[2][5] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ChiselTop.tappu.mem.tape[0][2] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold27 (.A(\ChiselTop.tappu.mem.tape[0][4] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold28 (.A(\ChiselTop.tappu.mem.tape[0][3] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold29 (.A(\ChiselTop.tappu.mem.tape[2][0] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold30 (.A(\ChiselTop.tappu.mem.tape[1][6] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold31 (.A(\ChiselTop.tappu.mem.tape[0][1] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold32 (.A(\ChiselTop.tappu.mem.tape[0][7] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold33 (.A(\ChiselTop.tappu.mem.tape[2][1] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ChiselTop.tappu.mem.tape[1][3] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold35 (.A(uo_out[0]),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold36 (.A(uo_out[4]),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0062_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold38 (.A(uo_out[1]),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold39 (.A(uo_out[2]),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold40 (.A(uo_out[5]),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0063_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold42 (.A(uo_out[6]),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold43 (.A(uo_out[7]),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold44 (.A(uo_out[3]),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold45 (.A(\ChiselTop.tappu.mem.tapeCounterReg[15] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0081_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0014_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold48 (.A(\ChiselTop.tappu.mem.tapeCounterReg[5] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold49 (.A(\ChiselTop.tappu.mem._GEN_198[1] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0203_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold51 (.A(\ChiselTop.tappu.mem.tapeCounterReg[3] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0069_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold53 (.A(\ChiselTop.tappu.mem.tapeCounterReg[14] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0080_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold55 (.A(\ChiselTop.tappu.mem._GEN_198[5] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold56 (.A(\ChiselTop.tappu.mem.tapeCounterReg[2] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0068_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0024_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0072_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold60 (.A(\ChiselTop.tappu.mem.tapeCounterReg[12] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0078_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ChiselTop.tappu.mem.tapeCounterReg[11] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0077_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold64 (.A(\ChiselTop.tappu.mem.tapeCounterReg[4] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold65 (.A(\ChiselTop.tappu.mem.tapeCounterReg[13] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0079_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold67 (.A(\ChiselTop.tappu.mem.tapeCounterReg[7] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0073_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold69 (.A(\ChiselTop.tappu.mem.tapeCounterReg[0] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold70 (.A(\ChiselTop.tappu.cpuState[0] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ChiselTop.tappu.mem._GEN_198[3] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold72 (.A(\ChiselTop.tappu.mem._GEN_198[2] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0027_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0075_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0012_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold76 (.A(\ChiselTop.tappu.cpuState[0] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold77 (.A(\ChiselTop.tappu.mem.tapeCounterReg[10] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0076_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0023_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0074_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold81 (.A(\ChiselTop.tappu.mem._GEN_198[4] ),
    .X(net204));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_4 FILLER_11_94 ();
 sg13g2_fill_2 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_117 ();
 sg13g2_decap_8 FILLER_11_122 ();
 sg13g2_decap_8 FILLER_11_129 ();
 sg13g2_decap_8 FILLER_11_136 ();
 sg13g2_decap_8 FILLER_11_143 ();
 sg13g2_decap_8 FILLER_11_150 ();
 sg13g2_decap_4 FILLER_11_157 ();
 sg13g2_fill_2 FILLER_11_161 ();
 sg13g2_decap_4 FILLER_11_167 ();
 sg13g2_decap_8 FILLER_11_174 ();
 sg13g2_decap_8 FILLER_11_181 ();
 sg13g2_decap_8 FILLER_11_188 ();
 sg13g2_decap_8 FILLER_11_195 ();
 sg13g2_decap_8 FILLER_11_202 ();
 sg13g2_decap_8 FILLER_11_209 ();
 sg13g2_decap_8 FILLER_11_220 ();
 sg13g2_decap_8 FILLER_11_227 ();
 sg13g2_decap_8 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_241 ();
 sg13g2_decap_8 FILLER_11_248 ();
 sg13g2_decap_8 FILLER_11_255 ();
 sg13g2_decap_8 FILLER_11_262 ();
 sg13g2_decap_8 FILLER_11_269 ();
 sg13g2_decap_8 FILLER_11_276 ();
 sg13g2_decap_8 FILLER_11_283 ();
 sg13g2_decap_8 FILLER_11_290 ();
 sg13g2_decap_8 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_304 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_decap_8 FILLER_11_332 ();
 sg13g2_decap_8 FILLER_11_339 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_353 ();
 sg13g2_decap_8 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_367 ();
 sg13g2_decap_8 FILLER_11_374 ();
 sg13g2_decap_8 FILLER_11_381 ();
 sg13g2_decap_8 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_63 ();
 sg13g2_fill_1 FILLER_12_65 ();
 sg13g2_fill_2 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_fill_2 FILLER_12_78 ();
 sg13g2_fill_1 FILLER_12_80 ();
 sg13g2_fill_1 FILLER_12_97 ();
 sg13g2_fill_1 FILLER_12_124 ();
 sg13g2_fill_1 FILLER_12_151 ();
 sg13g2_decap_4 FILLER_12_185 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_fill_2 FILLER_12_200 ();
 sg13g2_fill_1 FILLER_12_202 ();
 sg13g2_decap_8 FILLER_12_246 ();
 sg13g2_decap_8 FILLER_12_253 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_decap_8 FILLER_12_274 ();
 sg13g2_decap_8 FILLER_12_281 ();
 sg13g2_decap_8 FILLER_12_288 ();
 sg13g2_decap_8 FILLER_12_295 ();
 sg13g2_decap_8 FILLER_12_302 ();
 sg13g2_decap_8 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_decap_8 FILLER_12_323 ();
 sg13g2_decap_8 FILLER_12_330 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_344 ();
 sg13g2_decap_8 FILLER_12_351 ();
 sg13g2_decap_8 FILLER_12_358 ();
 sg13g2_decap_8 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_4 FILLER_13_49 ();
 sg13g2_fill_2 FILLER_13_53 ();
 sg13g2_fill_1 FILLER_13_124 ();
 sg13g2_fill_1 FILLER_13_143 ();
 sg13g2_fill_2 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_267 ();
 sg13g2_decap_8 FILLER_13_274 ();
 sg13g2_decap_8 FILLER_13_281 ();
 sg13g2_decap_8 FILLER_13_288 ();
 sg13g2_decap_8 FILLER_13_295 ();
 sg13g2_decap_8 FILLER_13_302 ();
 sg13g2_decap_8 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_316 ();
 sg13g2_decap_8 FILLER_13_323 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_337 ();
 sg13g2_decap_8 FILLER_13_344 ();
 sg13g2_decap_8 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_56 ();
 sg13g2_fill_2 FILLER_14_163 ();
 sg13g2_fill_1 FILLER_14_165 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_201 ();
 sg13g2_fill_2 FILLER_14_233 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_4 FILLER_15_42 ();
 sg13g2_fill_2 FILLER_15_46 ();
 sg13g2_fill_2 FILLER_15_100 ();
 sg13g2_decap_4 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_decap_8 FILLER_15_162 ();
 sg13g2_fill_2 FILLER_15_169 ();
 sg13g2_fill_1 FILLER_15_171 ();
 sg13g2_decap_4 FILLER_15_178 ();
 sg13g2_fill_1 FILLER_15_182 ();
 sg13g2_fill_2 FILLER_15_188 ();
 sg13g2_fill_1 FILLER_15_195 ();
 sg13g2_decap_8 FILLER_15_209 ();
 sg13g2_decap_4 FILLER_15_216 ();
 sg13g2_fill_2 FILLER_15_230 ();
 sg13g2_fill_1 FILLER_15_249 ();
 sg13g2_decap_8 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_decap_8 FILLER_15_282 ();
 sg13g2_decap_8 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_296 ();
 sg13g2_decap_8 FILLER_15_303 ();
 sg13g2_decap_8 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_331 ();
 sg13g2_decap_8 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_345 ();
 sg13g2_decap_8 FILLER_15_352 ();
 sg13g2_decap_8 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_366 ();
 sg13g2_decap_8 FILLER_15_373 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_fill_2 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_72 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_fill_2 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_138 ();
 sg13g2_fill_1 FILLER_16_145 ();
 sg13g2_fill_2 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_173 ();
 sg13g2_fill_2 FILLER_16_188 ();
 sg13g2_fill_1 FILLER_16_190 ();
 sg13g2_decap_4 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_278 ();
 sg13g2_decap_4 FILLER_16_285 ();
 sg13g2_fill_2 FILLER_16_289 ();
 sg13g2_decap_8 FILLER_16_295 ();
 sg13g2_decap_8 FILLER_16_302 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_decap_8 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_fill_2 FILLER_17_80 ();
 sg13g2_fill_1 FILLER_17_103 ();
 sg13g2_fill_1 FILLER_17_114 ();
 sg13g2_decap_4 FILLER_17_146 ();
 sg13g2_fill_2 FILLER_17_150 ();
 sg13g2_fill_1 FILLER_17_167 ();
 sg13g2_fill_1 FILLER_17_172 ();
 sg13g2_decap_4 FILLER_17_178 ();
 sg13g2_fill_2 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_188 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_fill_2 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_fill_2 FILLER_17_217 ();
 sg13g2_fill_1 FILLER_17_219 ();
 sg13g2_fill_2 FILLER_17_230 ();
 sg13g2_fill_2 FILLER_17_248 ();
 sg13g2_fill_1 FILLER_17_250 ();
 sg13g2_decap_4 FILLER_17_261 ();
 sg13g2_fill_2 FILLER_17_277 ();
 sg13g2_fill_1 FILLER_17_279 ();
 sg13g2_decap_4 FILLER_17_306 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_decap_4 FILLER_17_320 ();
 sg13g2_fill_2 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_344 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_fill_2 FILLER_18_93 ();
 sg13g2_fill_1 FILLER_18_95 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_decap_8 FILLER_18_108 ();
 sg13g2_decap_8 FILLER_18_115 ();
 sg13g2_fill_2 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_128 ();
 sg13g2_decap_8 FILLER_18_134 ();
 sg13g2_fill_1 FILLER_18_185 ();
 sg13g2_decap_4 FILLER_18_218 ();
 sg13g2_fill_1 FILLER_18_222 ();
 sg13g2_fill_2 FILLER_18_251 ();
 sg13g2_fill_1 FILLER_18_253 ();
 sg13g2_fill_2 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_53 ();
 sg13g2_fill_2 FILLER_19_80 ();
 sg13g2_fill_1 FILLER_19_82 ();
 sg13g2_fill_2 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_125 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_4 FILLER_19_147 ();
 sg13g2_decap_4 FILLER_19_159 ();
 sg13g2_fill_2 FILLER_19_178 ();
 sg13g2_decap_4 FILLER_19_185 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_215 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_decap_4 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_246 ();
 sg13g2_fill_2 FILLER_19_263 ();
 sg13g2_decap_4 FILLER_19_269 ();
 sg13g2_fill_2 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_342 ();
 sg13g2_decap_8 FILLER_19_349 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_370 ();
 sg13g2_decap_8 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_63 ();
 sg13g2_decap_4 FILLER_20_69 ();
 sg13g2_fill_1 FILLER_20_73 ();
 sg13g2_fill_2 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_121 ();
 sg13g2_fill_2 FILLER_20_193 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_2 FILLER_20_284 ();
 sg13g2_fill_2 FILLER_20_312 ();
 sg13g2_fill_1 FILLER_20_314 ();
 sg13g2_decap_4 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_127 ();
 sg13g2_fill_2 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_152 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_decap_8 FILLER_21_215 ();
 sg13g2_fill_2 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_232 ();
 sg13g2_decap_8 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_261 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_290 ();
 sg13g2_fill_2 FILLER_21_343 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_4 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_111 ();
 sg13g2_fill_2 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_120 ();
 sg13g2_fill_1 FILLER_22_164 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_decap_4 FILLER_22_206 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_fill_1 FILLER_22_222 ();
 sg13g2_fill_1 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_249 ();
 sg13g2_fill_2 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_271 ();
 sg13g2_fill_1 FILLER_22_278 ();
 sg13g2_decap_4 FILLER_22_287 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_fill_1 FILLER_23_143 ();
 sg13g2_fill_2 FILLER_23_175 ();
 sg13g2_decap_4 FILLER_23_182 ();
 sg13g2_fill_2 FILLER_23_186 ();
 sg13g2_decap_4 FILLER_23_192 ();
 sg13g2_fill_2 FILLER_23_196 ();
 sg13g2_fill_1 FILLER_23_203 ();
 sg13g2_decap_4 FILLER_23_233 ();
 sg13g2_decap_8 FILLER_23_246 ();
 sg13g2_decap_8 FILLER_23_293 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_fill_2 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_311 ();
 sg13g2_fill_2 FILLER_23_321 ();
 sg13g2_fill_1 FILLER_23_332 ();
 sg13g2_decap_4 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_fill_1 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_82 ();
 sg13g2_decap_4 FILLER_24_89 ();
 sg13g2_fill_1 FILLER_24_145 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_198 ();
 sg13g2_fill_2 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_281 ();
 sg13g2_fill_1 FILLER_24_291 ();
 sg13g2_decap_4 FILLER_24_332 ();
 sg13g2_fill_2 FILLER_24_336 ();
 sg13g2_decap_4 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_347 ();
 sg13g2_decap_4 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_356 ();
 sg13g2_decap_4 FILLER_24_379 ();
 sg13g2_fill_2 FILLER_24_383 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_4 FILLER_25_63 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_117 ();
 sg13g2_fill_1 FILLER_25_119 ();
 sg13g2_decap_4 FILLER_25_125 ();
 sg13g2_decap_4 FILLER_25_142 ();
 sg13g2_fill_2 FILLER_25_146 ();
 sg13g2_fill_2 FILLER_25_183 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_decap_4 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_251 ();
 sg13g2_decap_4 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_2 FILLER_25_283 ();
 sg13g2_decap_4 FILLER_25_305 ();
 sg13g2_fill_1 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_fill_1 FILLER_25_380 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_62 ();
 sg13g2_decap_8 FILLER_26_116 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_fill_2 FILLER_26_170 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_212 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_decap_8 FILLER_26_225 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_decap_8 FILLER_26_293 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_324 ();
 sg13g2_decap_4 FILLER_26_341 ();
 sg13g2_fill_2 FILLER_26_345 ();
 sg13g2_fill_1 FILLER_26_356 ();
 sg13g2_fill_2 FILLER_26_379 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_42 ();
 sg13g2_fill_1 FILLER_27_107 ();
 sg13g2_decap_8 FILLER_27_115 ();
 sg13g2_fill_1 FILLER_27_122 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_160 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_fill_2 FILLER_27_234 ();
 sg13g2_fill_1 FILLER_27_247 ();
 sg13g2_decap_8 FILLER_27_256 ();
 sg13g2_decap_4 FILLER_27_263 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_decap_4 FILLER_27_381 ();
 sg13g2_fill_1 FILLER_27_385 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_4 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_fill_2 FILLER_28_96 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_decap_4 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_decap_4 FILLER_28_136 ();
 sg13g2_decap_4 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_fill_2 FILLER_28_230 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_decap_4 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_247 ();
 sg13g2_decap_4 FILLER_28_254 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_fill_1 FILLER_28_277 ();
 sg13g2_fill_1 FILLER_28_282 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_fill_2 FILLER_28_332 ();
 sg13g2_decap_8 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_fill_2 FILLER_28_379 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_83 ();
 sg13g2_decap_4 FILLER_29_132 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_decap_4 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_fill_2 FILLER_29_242 ();
 sg13g2_fill_1 FILLER_29_244 ();
 sg13g2_decap_4 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_298 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_decap_4 FILLER_29_325 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_fill_1 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_fill_2 FILLER_29_389 ();
 sg13g2_fill_1 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_4 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_86 ();
 sg13g2_fill_2 FILLER_30_97 ();
 sg13g2_fill_1 FILLER_30_99 ();
 sg13g2_decap_4 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_132 ();
 sg13g2_fill_1 FILLER_30_134 ();
 sg13g2_decap_8 FILLER_30_143 ();
 sg13g2_decap_4 FILLER_30_150 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_191 ();
 sg13g2_fill_2 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_fill_2 FILLER_30_219 ();
 sg13g2_decap_8 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_233 ();
 sg13g2_decap_4 FILLER_30_239 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_fill_1 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_265 ();
 sg13g2_decap_4 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_decap_4 FILLER_30_306 ();
 sg13g2_decap_4 FILLER_30_334 ();
 sg13g2_decap_4 FILLER_30_343 ();
 sg13g2_fill_2 FILLER_30_347 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_370 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_4 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_decap_4 FILLER_31_65 ();
 sg13g2_fill_1 FILLER_31_69 ();
 sg13g2_decap_8 FILLER_31_74 ();
 sg13g2_decap_8 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_92 ();
 sg13g2_fill_2 FILLER_31_109 ();
 sg13g2_decap_4 FILLER_31_131 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_decap_4 FILLER_31_181 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_decap_4 FILLER_31_219 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_decap_4 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_282 ();
 sg13g2_decap_4 FILLER_31_326 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_4 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_113 ();
 sg13g2_fill_2 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_135 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_fill_2 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_192 ();
 sg13g2_decap_4 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_fill_2 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_decap_4 FILLER_32_278 ();
 sg13g2_fill_2 FILLER_32_287 ();
 sg13g2_fill_1 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_313 ();
 sg13g2_fill_2 FILLER_32_318 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_fill_1 FILLER_33_100 ();
 sg13g2_decap_8 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_decap_8 FILLER_33_174 ();
 sg13g2_decap_8 FILLER_33_181 ();
 sg13g2_decap_4 FILLER_33_188 ();
 sg13g2_fill_1 FILLER_33_192 ();
 sg13g2_decap_4 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_263 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_fill_2 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_313 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_4 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_109 ();
 sg13g2_decap_8 FILLER_34_115 ();
 sg13g2_decap_8 FILLER_34_122 ();
 sg13g2_decap_8 FILLER_34_129 ();
 sg13g2_decap_8 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_143 ();
 sg13g2_decap_8 FILLER_34_149 ();
 sg13g2_decap_8 FILLER_34_156 ();
 sg13g2_decap_8 FILLER_34_163 ();
 sg13g2_decap_8 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_184 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_fill_2 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_decap_4 FILLER_34_309 ();
 sg13g2_fill_1 FILLER_34_313 ();
 sg13g2_decap_4 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_fill_2 FILLER_34_359 ();
 sg13g2_fill_2 FILLER_34_380 ();
 sg13g2_fill_1 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_4 FILLER_35_276 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_fill_1 FILLER_35_356 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_decap_4 FILLER_36_286 ();
 sg13g2_fill_2 FILLER_36_290 ();
 sg13g2_fill_2 FILLER_36_296 ();
 sg13g2_fill_2 FILLER_36_308 ();
 sg13g2_fill_1 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_decap_4 FILLER_36_376 ();
 sg13g2_fill_2 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_4 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_248 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_decap_8 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_4 FILLER_37_382 ();
 sg13g2_fill_1 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_391 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_fill_2 FILLER_38_264 ();
 sg13g2_fill_1 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_4 FILLER_38_285 ();
 sg13g2_fill_2 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_302 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule

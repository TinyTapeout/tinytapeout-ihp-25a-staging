module tt_um_ezchips_calc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \DEBUG_SIGS_GTKWAVE.@0$slideswitch[0] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$slideswitch[1] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$slideswitch[2] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$slideswitch[3] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$slideswitch[4] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$slideswitch[5] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$slideswitch[6] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$slideswitch[7] ;
 wire net44;
 wire net9;
 wire net43;
 wire net42;
 wire clknet_2_3__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_0_clk;
 wire \DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[0] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[1] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[2] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[3] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[4] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[5] ;
 wire \DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[6] ;
 wire \DEBUG_SIGS_GTKWAVE./digit[0]./leds[0].@0$viz_lit ;
 wire \DEBUG_SIGS_GTKWAVE./digit[0]./leds[1].@0$viz_lit ;
 wire \DEBUG_SIGS_GTKWAVE./digit[0]./leds[2].@0$viz_lit ;
 wire \DEBUG_SIGS_GTKWAVE./digit[0]./leds[3].@0$viz_lit ;
 wire \DEBUG_SIGS_GTKWAVE./digit[0]./leds[4].@0$viz_lit ;
 wire \DEBUG_SIGS_GTKWAVE./digit[0]./leds[5].@0$viz_lit ;
 wire \DEBUG_SIGS_GTKWAVE./digit[0]./leds[6].@0$viz_lit ;
 wire net50;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$equals_in ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$op[0] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$op[1] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$val2[0] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$val2[1] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$val2[2] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$val2[3] ;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[0] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[1] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[2] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[3] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[4] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[5] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[6] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[7] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[0] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[1] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[2] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[3] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[0] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[1] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[2] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[3] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[4] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[5] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[6] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[7] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[0] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[1] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[2] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[3] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[4] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[5] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[6] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[7] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[0] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[1] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[2] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[3] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[4] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[5] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[6] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[7] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$reset ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[0] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[1] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[2] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[3] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[4] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[5] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[6] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[7] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[0] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[1] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[2] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[3] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[4] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[5] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[6] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[7] ;
 wire \DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$valid ;
 wire \DEBUG_SIGS_GTKWAVE./switch[0].@0$viz_switch ;
 wire \DEBUG_SIGS_GTKWAVE./switch[1].@0$viz_switch ;
 wire \DEBUG_SIGS_GTKWAVE./switch[2].@0$viz_switch ;
 wire \DEBUG_SIGS_GTKWAVE./switch[3].@0$viz_switch ;
 wire \DEBUG_SIGS_GTKWAVE./switch[4].@0$viz_switch ;
 wire \DEBUG_SIGS_GTKWAVE./switch[5].@0$viz_switch ;
 wire \DEBUG_SIGS_GTKWAVE./switch[6].@0$viz_switch ;
 wire \DEBUG_SIGS_GTKWAVE./switch[7].@0$viz_switch ;
 wire FpgaPins_Fpga_CALC_equals_in_a1;
 wire FpgaPins_Fpga_CALC_equals_in_a2;
 wire \FpgaPins_Fpga_CALC_op_a1[0] ;
 wire \FpgaPins_Fpga_CALC_op_a1[1] ;
 wire \FpgaPins_Fpga_CALC_val2_a1[0] ;
 wire \FpgaPins_Fpga_CALC_val2_a1[1] ;
 wire \FpgaPins_Fpga_CALC_val2_a1[2] ;
 wire \FpgaPins_Fpga_CALC_val2_a1[3] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net45;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;

 sg13g2_inv_1 _393_ (.Y(_364_),
    .A(net44));
 sg13g2_inv_1 _394_ (.Y(_365_),
    .A(net43));
 sg13g2_inv_1 _395_ (.Y(_366_),
    .A(net46));
 sg13g2_inv_1 _396_ (.Y(_367_),
    .A(net48));
 sg13g2_inv_1 _397_ (.Y(_368_),
    .A(net70));
 sg13g2_inv_1 _398_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$reset ),
    .A(net1));
 sg13g2_inv_1 _399_ (.Y(_369_),
    .A(net65));
 sg13g2_inv_1 _400_ (.Y(_370_),
    .A(net63));
 sg13g2_inv_1 _401_ (.Y(_371_),
    .A(net62));
 sg13g2_inv_1 _402_ (.Y(_372_),
    .A(_009_));
 sg13g2_inv_1 _403_ (.Y(_016_),
    .A(_001_));
 sg13g2_inv_1 _404_ (.Y(_017_),
    .A(_003_));
 sg13g2_nand2b_2 _405_ (.Y(_018_),
    .B(net42),
    .A_N(FpgaPins_Fpga_CALC_equals_in_a2));
 sg13g2_nor2_2 _406_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$reset ),
    .B(_018_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$valid ));
 sg13g2_xor2_1 _407_ (.B(net66),
    .A(net70),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[0] ));
 sg13g2_nand2_1 _408_ (.Y(_019_),
    .A(net70),
    .B(net65));
 sg13g2_inv_1 _409_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[0] ),
    .A(_019_));
 sg13g2_and2_1 _410_ (.A(net67),
    .B(_000_),
    .X(_020_));
 sg13g2_nand2_1 _411_ (.Y(_021_),
    .A(\FpgaPins_Fpga_CALC_val2_a1[0] ),
    .B(_000_));
 sg13g2_nand2_1 _412_ (.Y(_022_),
    .A(net67),
    .B(_002_));
 sg13g2_mux2_1 _413_ (.A0(_022_),
    .A1(_002_),
    .S(_011_),
    .X(_023_));
 sg13g2_nor2_1 _414_ (.A(\FpgaPins_Fpga_CALC_val2_a1[3] ),
    .B(net62),
    .Y(_024_));
 sg13g2_o21ai_1 _415_ (.B1(_024_),
    .Y(_025_),
    .A1(_370_),
    .A2(_023_));
 sg13g2_nand2b_1 _416_ (.Y(_026_),
    .B(_010_),
    .A_N(net61));
 sg13g2_nor4_2 _417_ (.A(_364_),
    .B(net67),
    .C(net64),
    .Y(_027_),
    .D(_026_));
 sg13g2_nor2b_1 _418_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[7] ),
    .B_N(net67),
    .Y(_028_));
 sg13g2_nor2_1 _419_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[6] ),
    .B(_011_),
    .Y(_029_));
 sg13g2_or4_1 _420_ (.A(net64),
    .B(_026_),
    .C(_028_),
    .D(_029_),
    .X(_030_));
 sg13g2_nor2b_1 _421_ (.A(_027_),
    .B_N(_030_),
    .Y(_031_));
 sg13g2_inv_1 _422_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[7] ),
    .A(_031_));
 sg13g2_a21oi_1 _423_ (.A1(_372_),
    .A2(_030_),
    .Y(_032_),
    .B1(_027_));
 sg13g2_a21o_1 _424_ (.A2(_030_),
    .A1(_372_),
    .B1(_027_),
    .X(_033_));
 sg13g2_and2_1 _425_ (.A(_370_),
    .B(_023_),
    .X(_034_));
 sg13g2_a221oi_1 _426_ (.B2(_372_),
    .C1(_027_),
    .B1(_030_),
    .A1(_370_),
    .Y(_035_),
    .A2(_023_));
 sg13g2_nor2_1 _427_ (.A(_025_),
    .B(_035_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[6] ));
 sg13g2_nor3_1 _428_ (.A(_002_),
    .B(_025_),
    .C(_035_),
    .Y(_036_));
 sg13g2_xor2_1 _429_ (.B(_036_),
    .A(_011_),
    .X(_037_));
 sg13g2_inv_1 _430_ (.Y(_038_),
    .A(_037_));
 sg13g2_xnor2_1 _431_ (.Y(_039_),
    .A(_003_),
    .B(_037_));
 sg13g2_o21ai_1 _432_ (.B1(_033_),
    .Y(_040_),
    .A1(_025_),
    .A2(_034_));
 sg13g2_nor2_1 _433_ (.A(net61),
    .B(_040_),
    .Y(_041_));
 sg13g2_nand2b_1 _434_ (.Y(_042_),
    .B(_371_),
    .A_N(_040_));
 sg13g2_nand2_1 _435_ (.Y(_043_),
    .A(net61),
    .B(_032_));
 sg13g2_nand2_1 _436_ (.Y(_044_),
    .A(_042_),
    .B(_043_));
 sg13g2_mux2_2 _437_ (.A0(_016_),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[4] ),
    .S(_031_),
    .X(_045_));
 sg13g2_nor3_1 _438_ (.A(net59),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[3] ),
    .C(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[2] ),
    .Y(_046_));
 sg13g2_nor2_1 _439_ (.A(net67),
    .B(_000_),
    .Y(_047_));
 sg13g2_nor2_1 _440_ (.A(net70),
    .B(net69),
    .Y(_048_));
 sg13g2_a21oi_1 _441_ (.A1(_046_),
    .A2(_048_),
    .Y(_049_),
    .B1(net57));
 sg13g2_nor2_1 _442_ (.A(_020_),
    .B(_047_),
    .Y(_050_));
 sg13g2_or4_1 _443_ (.A(_020_),
    .B(_045_),
    .C(_047_),
    .D(_049_),
    .X(_051_));
 sg13g2_and2_1 _444_ (.A(_010_),
    .B(_021_),
    .X(_052_));
 sg13g2_o21ai_1 _445_ (.B1(_052_),
    .Y(_053_),
    .A1(_045_),
    .A2(_047_));
 sg13g2_a221oi_1 _446_ (.B2(_053_),
    .C1(_041_),
    .B1(_051_),
    .A1(net61),
    .Y(_054_),
    .A2(_032_));
 sg13g2_o21ai_1 _447_ (.B1(_042_),
    .Y(_055_),
    .A1(net64),
    .A2(_037_));
 sg13g2_and2_1 _448_ (.A(net57),
    .B(_043_),
    .X(_056_));
 sg13g2_a22oi_1 _449_ (.Y(_057_),
    .B1(_055_),
    .B2(_056_),
    .A2(_054_),
    .A1(_039_));
 sg13g2_inv_1 _450_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[5] ),
    .A(_057_));
 sg13g2_mux2_1 _451_ (.A0(_050_),
    .A1(_000_),
    .S(_057_),
    .X(_058_));
 sg13g2_nor2_1 _452_ (.A(net64),
    .B(_058_),
    .Y(_059_));
 sg13g2_xnor2_1 _453_ (.Y(_060_),
    .A(net56),
    .B(_058_));
 sg13g2_mux2_1 _454_ (.A0(_002_),
    .A1(_022_),
    .S(_045_),
    .X(_061_));
 sg13g2_a21oi_1 _455_ (.A1(_060_),
    .A2(_061_),
    .Y(_062_),
    .B1(_059_));
 sg13g2_xnor2_1 _456_ (.Y(_063_),
    .A(_020_),
    .B(_039_));
 sg13g2_nor2_1 _457_ (.A(_057_),
    .B(_063_),
    .Y(_064_));
 sg13g2_a21oi_2 _458_ (.B1(_064_),
    .Y(_065_),
    .A2(_057_),
    .A1(_037_));
 sg13g2_xnor2_1 _459_ (.Y(_066_),
    .A(_004_),
    .B(_065_));
 sg13g2_nand2_1 _460_ (.Y(_067_),
    .A(_371_),
    .B(_065_));
 sg13g2_o21ai_1 _461_ (.B1(_067_),
    .Y(_068_),
    .A1(_062_),
    .A2(_066_));
 sg13g2_a22oi_1 _462_ (.Y(_069_),
    .B1(_039_),
    .B2(_021_),
    .A2(_038_),
    .A1(net56));
 sg13g2_xnor2_1 _463_ (.Y(_070_),
    .A(_044_),
    .B(_069_));
 sg13g2_mux2_1 _464_ (.A0(_040_),
    .A1(_070_),
    .S(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[5] ),
    .X(_071_));
 sg13g2_inv_1 _465_ (.Y(_072_),
    .A(_071_));
 sg13g2_xor2_1 _466_ (.B(_071_),
    .A(net59),
    .X(_073_));
 sg13g2_a22oi_1 _467_ (.Y(_074_),
    .B1(_073_),
    .B2(_068_),
    .A2(_072_),
    .A1(net57));
 sg13g2_inv_1 _468_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[4] ),
    .A(_074_));
 sg13g2_xnor2_1 _469_ (.Y(_075_),
    .A(_062_),
    .B(_066_));
 sg13g2_nand2_1 _470_ (.Y(_076_),
    .A(_065_),
    .B(_074_));
 sg13g2_o21ai_1 _471_ (.B1(_076_),
    .Y(_077_),
    .A1(_074_),
    .A2(_075_));
 sg13g2_nand2_1 _472_ (.Y(_078_),
    .A(net57),
    .B(_077_));
 sg13g2_xor2_1 _473_ (.B(_077_),
    .A(net57),
    .X(_079_));
 sg13g2_nand2_1 _474_ (.Y(_080_),
    .A(_058_),
    .B(_074_));
 sg13g2_xor2_1 _475_ (.B(_061_),
    .A(_060_),
    .X(_081_));
 sg13g2_o21ai_1 _476_ (.B1(_080_),
    .Y(_082_),
    .A1(_074_),
    .A2(_081_));
 sg13g2_nor2_1 _477_ (.A(net61),
    .B(_082_),
    .Y(_083_));
 sg13g2_nand2_1 _478_ (.Y(_084_),
    .A(net61),
    .B(_082_));
 sg13g2_nand2_1 _479_ (.Y(_085_),
    .A(net65),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[3] ));
 sg13g2_xor2_1 _480_ (.B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[3] ),
    .A(net66),
    .X(_086_));
 sg13g2_inv_1 _481_ (.Y(_087_),
    .A(_086_));
 sg13g2_nand2_1 _482_ (.Y(_088_),
    .A(net66),
    .B(_086_));
 sg13g2_nor2_1 _483_ (.A(_002_),
    .B(_074_),
    .Y(_089_));
 sg13g2_xor2_1 _484_ (.B(_089_),
    .A(_045_),
    .X(_090_));
 sg13g2_xnor2_1 _485_ (.Y(_091_),
    .A(_017_),
    .B(_090_));
 sg13g2_and2_1 _486_ (.A(net56),
    .B(_090_),
    .X(_092_));
 sg13g2_a21o_1 _487_ (.A2(_091_),
    .A1(_088_),
    .B1(_092_),
    .X(_093_));
 sg13g2_and2_1 _488_ (.A(_084_),
    .B(_093_),
    .X(_094_));
 sg13g2_a221oi_1 _489_ (.B2(_088_),
    .C1(_083_),
    .B1(_091_),
    .A1(net56),
    .Y(_095_),
    .A2(_090_));
 sg13g2_nand3b_1 _490_ (.B(_079_),
    .C(_084_),
    .Y(_096_),
    .A_N(_095_));
 sg13g2_nand2b_1 _491_ (.Y(_097_),
    .B(net57),
    .A_N(net59));
 sg13g2_a21oi_1 _492_ (.A1(net59),
    .A2(_068_),
    .Y(_098_),
    .B1(_071_));
 sg13g2_o21ai_1 _493_ (.B1(_098_),
    .Y(_099_),
    .A1(_068_),
    .A2(_097_));
 sg13g2_nand2_1 _494_ (.Y(_100_),
    .A(_078_),
    .B(_099_));
 sg13g2_nor2b_2 _495_ (.A(_100_),
    .B_N(_096_),
    .Y(_101_));
 sg13g2_inv_1 _496_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[3] ),
    .A(_101_));
 sg13g2_mux2_1 _497_ (.A0(_087_),
    .A1(_005_),
    .S(_101_),
    .X(_102_));
 sg13g2_nor2b_1 _498_ (.A(_083_),
    .B_N(_084_),
    .Y(_103_));
 sg13g2_xnor2_1 _499_ (.Y(_104_),
    .A(_093_),
    .B(_103_));
 sg13g2_mux2_2 _500_ (.A0(_104_),
    .A1(_082_),
    .S(_101_),
    .X(_105_));
 sg13g2_inv_1 _501_ (.Y(_106_),
    .A(_105_));
 sg13g2_nor2_1 _502_ (.A(net58),
    .B(_105_),
    .Y(_107_));
 sg13g2_and2_1 _503_ (.A(net58),
    .B(_105_),
    .X(_108_));
 sg13g2_xor2_1 _504_ (.B(_091_),
    .A(_088_),
    .X(_109_));
 sg13g2_mux2_2 _505_ (.A0(_109_),
    .A1(_090_),
    .S(_101_),
    .X(_110_));
 sg13g2_or2_1 _506_ (.X(_111_),
    .B(_102_),
    .A(_017_));
 sg13g2_nor2_1 _507_ (.A(_369_),
    .B(net68),
    .Y(_112_));
 sg13g2_xnor2_1 _508_ (.Y(_113_),
    .A(net63),
    .B(_102_));
 sg13g2_o21ai_1 _509_ (.B1(_111_),
    .Y(_114_),
    .A1(_112_),
    .A2(_113_));
 sg13g2_xnor2_1 _510_ (.Y(_115_),
    .A(_004_),
    .B(_110_));
 sg13g2_xor2_1 _511_ (.B(_110_),
    .A(_004_),
    .X(_116_));
 sg13g2_a22oi_1 _512_ (.Y(_117_),
    .B1(_114_),
    .B2(_116_),
    .A2(_110_),
    .A1(_371_));
 sg13g2_a221oi_1 _513_ (.B2(_116_),
    .C1(_107_),
    .B1(_114_),
    .A1(_371_),
    .Y(_118_),
    .A2(_110_));
 sg13g2_nor2_1 _514_ (.A(_108_),
    .B(_118_),
    .Y(_119_));
 sg13g2_xnor2_1 _515_ (.Y(_120_),
    .A(net66),
    .B(net68));
 sg13g2_nand2_1 _516_ (.Y(_121_),
    .A(_048_),
    .B(_120_));
 sg13g2_xnor2_1 _517_ (.Y(_122_),
    .A(net58),
    .B(_105_));
 sg13g2_nor4_1 _518_ (.A(_113_),
    .B(_115_),
    .C(_121_),
    .D(_122_),
    .Y(_123_));
 sg13g2_nand2_1 _519_ (.Y(_124_),
    .A(_077_),
    .B(_101_));
 sg13g2_nor3_1 _520_ (.A(_079_),
    .B(_083_),
    .C(_094_),
    .Y(_125_));
 sg13g2_nand2_1 _521_ (.Y(_126_),
    .A(_096_),
    .B(_100_));
 sg13g2_o21ai_1 _522_ (.B1(_124_),
    .Y(_127_),
    .A1(_125_),
    .A2(_126_));
 sg13g2_a21oi_1 _523_ (.A1(_078_),
    .A2(_096_),
    .Y(_128_),
    .B1(_099_));
 sg13g2_nor3_1 _524_ (.A(_123_),
    .B(_127_),
    .C(_128_),
    .Y(_129_));
 sg13g2_o21ai_1 _525_ (.B1(_129_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[2] ),
    .A1(_108_),
    .A2(_118_));
 sg13g2_xnor2_1 _526_ (.Y(_130_),
    .A(_112_),
    .B(_113_));
 sg13g2_mux2_1 _527_ (.A0(_102_),
    .A1(_130_),
    .S(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[2] ),
    .X(_131_));
 sg13g2_xnor2_1 _528_ (.Y(_132_),
    .A(_114_),
    .B(_115_));
 sg13g2_mux2_1 _529_ (.A0(_110_),
    .A1(_132_),
    .S(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[2] ),
    .X(_133_));
 sg13g2_nor2_1 _530_ (.A(net57),
    .B(_133_),
    .Y(_134_));
 sg13g2_and2_1 _531_ (.A(net60),
    .B(_131_),
    .X(_135_));
 sg13g2_nor2_1 _532_ (.A(net62),
    .B(_131_),
    .Y(_136_));
 sg13g2_nand2b_2 _533_ (.Y(_137_),
    .B(net66),
    .A_N(net69));
 sg13g2_mux2_1 _534_ (.A0(_006_),
    .A1(_120_),
    .S(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[2] ),
    .X(_138_));
 sg13g2_inv_1 _535_ (.Y(_139_),
    .A(_138_));
 sg13g2_xnor2_1 _536_ (.Y(_140_),
    .A(_003_),
    .B(_138_));
 sg13g2_a22oi_1 _537_ (.Y(_141_),
    .B1(_140_),
    .B2(_137_),
    .A2(_139_),
    .A1(net56));
 sg13g2_a221oi_1 _538_ (.B2(_137_),
    .C1(_136_),
    .B1(_140_),
    .A1(net56),
    .Y(_142_),
    .A2(_139_));
 sg13g2_or2_1 _539_ (.X(_143_),
    .B(_142_),
    .A(_135_));
 sg13g2_nor3_2 _540_ (.A(_134_),
    .B(_135_),
    .C(_142_),
    .Y(_144_));
 sg13g2_or3_1 _541_ (.A(_134_),
    .B(_135_),
    .C(_142_),
    .X(_145_));
 sg13g2_o21ai_1 _542_ (.B1(_128_),
    .Y(_146_),
    .A1(_119_),
    .A2(_127_));
 sg13g2_a21oi_1 _543_ (.A1(_119_),
    .A2(_127_),
    .Y(_147_),
    .B1(_128_));
 sg13g2_xor2_1 _544_ (.B(_122_),
    .A(_117_),
    .X(_148_));
 sg13g2_mux2_1 _545_ (.A0(_106_),
    .A1(_148_),
    .S(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[2] ),
    .X(_149_));
 sg13g2_nor2_1 _546_ (.A(_133_),
    .B(_149_),
    .Y(_150_));
 sg13g2_a21oi_2 _547_ (.B1(_149_),
    .Y(_151_),
    .A2(_133_),
    .A1(net57));
 sg13g2_nand2_1 _548_ (.Y(_152_),
    .A(_147_),
    .B(_151_));
 sg13g2_inv_1 _549_ (.Y(_153_),
    .A(_152_));
 sg13g2_nor2_2 _550_ (.A(_144_),
    .B(_152_),
    .Y(_154_));
 sg13g2_inv_1 _551_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[1] ),
    .A(_154_));
 sg13g2_or2_1 _552_ (.X(_155_),
    .B(_136_),
    .A(_135_));
 sg13g2_xor2_1 _553_ (.B(_155_),
    .A(_141_),
    .X(_156_));
 sg13g2_nand2_1 _554_ (.Y(_157_),
    .A(_131_),
    .B(_154_));
 sg13g2_o21ai_1 _555_ (.B1(_157_),
    .Y(_158_),
    .A1(_154_),
    .A2(_156_));
 sg13g2_and2_1 _556_ (.A(net59),
    .B(_158_),
    .X(_159_));
 sg13g2_xnor2_1 _557_ (.Y(_160_),
    .A(_137_),
    .B(_140_));
 sg13g2_mux2_1 _558_ (.A0(_160_),
    .A1(_138_),
    .S(_154_),
    .X(_161_));
 sg13g2_nand2_1 _559_ (.Y(_162_),
    .A(net60),
    .B(_161_));
 sg13g2_nand2_1 _560_ (.Y(_163_),
    .A(_369_),
    .B(net69));
 sg13g2_nor3_1 _561_ (.A(_007_),
    .B(_144_),
    .C(_152_),
    .Y(_164_));
 sg13g2_a22oi_1 _562_ (.Y(_165_),
    .B1(_163_),
    .B2(_137_),
    .A2(_153_),
    .A1(_145_));
 sg13g2_or3_1 _563_ (.A(_017_),
    .B(_164_),
    .C(_165_),
    .X(_166_));
 sg13g2_o21ai_1 _564_ (.B1(_017_),
    .Y(_167_),
    .A1(_164_),
    .A2(_165_));
 sg13g2_a22oi_1 _565_ (.Y(_168_),
    .B1(_166_),
    .B2(_167_),
    .A2(_369_),
    .A1(net70));
 sg13g2_nor3_1 _566_ (.A(net56),
    .B(_164_),
    .C(_165_),
    .Y(_169_));
 sg13g2_xnor2_1 _567_ (.Y(_170_),
    .A(_004_),
    .B(_161_));
 sg13g2_o21ai_1 _568_ (.B1(_170_),
    .Y(_171_),
    .A1(_168_),
    .A2(_169_));
 sg13g2_nor2_1 _569_ (.A(net59),
    .B(_158_),
    .Y(_172_));
 sg13g2_a21oi_1 _570_ (.A1(_166_),
    .A2(_167_),
    .Y(_173_),
    .B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[0] ));
 sg13g2_a221oi_1 _571_ (.B2(_170_),
    .C1(_172_),
    .B1(_173_),
    .A1(_162_),
    .Y(_174_),
    .A2(_171_));
 sg13g2_nor2_1 _572_ (.A(_150_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[1] ),
    .Y(_175_));
 sg13g2_nor2b_1 _573_ (.A(_134_),
    .B_N(_149_),
    .Y(_176_));
 sg13g2_nor2_1 _574_ (.A(_151_),
    .B(_176_),
    .Y(_177_));
 sg13g2_a221oi_1 _575_ (.B2(_143_),
    .C1(_153_),
    .B1(_177_),
    .A1(_144_),
    .Y(_178_),
    .A2(_151_));
 sg13g2_and2_1 _576_ (.A(_146_),
    .B(_151_),
    .X(_179_));
 sg13g2_a21oi_1 _577_ (.A1(_143_),
    .A2(_179_),
    .Y(_180_),
    .B1(_147_));
 sg13g2_nor3_1 _578_ (.A(_175_),
    .B(_178_),
    .C(_180_),
    .Y(_181_));
 sg13g2_o21ai_1 _579_ (.B1(_181_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[0] ),
    .A1(_159_),
    .A2(_174_));
 sg13g2_and2_1 _580_ (.A(\FpgaPins_Fpga_CALC_op_a1[0] ),
    .B(\FpgaPins_Fpga_CALC_op_a1[1] ),
    .X(_182_));
 sg13g2_nand2_2 _581_ (.Y(_183_),
    .A(\FpgaPins_Fpga_CALC_op_a1[0] ),
    .B(\FpgaPins_Fpga_CALC_op_a1[1] ));
 sg13g2_nor2_1 _582_ (.A(\FpgaPins_Fpga_CALC_op_a1[1] ),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[0] ),
    .Y(_184_));
 sg13g2_nor2b_1 _583_ (.A(\FpgaPins_Fpga_CALC_op_a1[0] ),
    .B_N(\FpgaPins_Fpga_CALC_op_a1[1] ),
    .Y(_185_));
 sg13g2_nand2b_2 _584_ (.Y(_186_),
    .B(\FpgaPins_Fpga_CALC_op_a1[1] ),
    .A_N(\FpgaPins_Fpga_CALC_op_a1[0] ));
 sg13g2_o21ai_1 _585_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$valid ),
    .Y(_187_),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[0] ),
    .A2(_186_));
 sg13g2_nor2_1 _586_ (.A(_184_),
    .B(_187_),
    .Y(_188_));
 sg13g2_o21ai_1 _587_ (.B1(_188_),
    .Y(_189_),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[0] ),
    .A2(_183_));
 sg13g2_nand2_1 _588_ (.Y(_190_),
    .A(net1),
    .B(_018_));
 sg13g2_or2_1 _589_ (.X(_191_),
    .B(net54),
    .A(_008_));
 sg13g2_and2_2 _590_ (.A(_189_),
    .B(_191_),
    .X(_192_));
 sg13g2_inv_2 _591_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[0] ),
    .A(_192_));
 sg13g2_nand2b_2 _592_ (.Y(_193_),
    .B(\FpgaPins_Fpga_CALC_op_a1[0] ),
    .A_N(\FpgaPins_Fpga_CALC_op_a1[1] ));
 sg13g2_nand2_2 _593_ (.Y(_194_),
    .A(net63),
    .B(net69));
 sg13g2_xor2_1 _594_ (.B(net69),
    .A(net63),
    .X(_195_));
 sg13g2_a21oi_1 _595_ (.A1(_368_),
    .A2(net65),
    .Y(_196_),
    .B1(_195_));
 sg13g2_nand3_1 _596_ (.B(net65),
    .C(_195_),
    .A(_368_),
    .Y(_197_));
 sg13g2_nor2b_1 _597_ (.A(_196_),
    .B_N(_197_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[1] ));
 sg13g2_nor2_1 _598_ (.A(_193_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[1] ),
    .Y(_198_));
 sg13g2_or2_2 _599_ (.X(_199_),
    .B(\FpgaPins_Fpga_CALC_op_a1[1] ),
    .A(\FpgaPins_Fpga_CALC_op_a1[0] ));
 sg13g2_nand2_1 _600_ (.Y(_200_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[0] ),
    .B(_195_));
 sg13g2_xnor2_1 _601_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[1] ),
    .A(_019_),
    .B(_195_));
 sg13g2_nor2_1 _602_ (.A(_199_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[1] ),
    .Y(_201_));
 sg13g2_a22oi_1 _603_ (.Y(_202_),
    .B1(net69),
    .B2(net65),
    .A2(net63),
    .A1(net70));
 sg13g2_nor2_1 _604_ (.A(_019_),
    .B(_194_),
    .Y(_203_));
 sg13g2_nor2_1 _605_ (.A(_202_),
    .B(_203_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[1] ));
 sg13g2_o21ai_1 _606_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$valid ),
    .Y(_204_),
    .A1(_186_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[1] ));
 sg13g2_nor3_1 _607_ (.A(_198_),
    .B(_201_),
    .C(_204_),
    .Y(_205_));
 sg13g2_o21ai_1 _608_ (.B1(_205_),
    .Y(_206_),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[1] ),
    .A2(_183_));
 sg13g2_o21ai_1 _609_ (.B1(_206_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[1] ),
    .A1(net47),
    .A2(net54));
 sg13g2_inv_1 _610_ (.Y(_207_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[1] ));
 sg13g2_nor2_1 _611_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[2] ),
    .B(_183_),
    .Y(_208_));
 sg13g2_nand2_1 _612_ (.Y(_209_),
    .A(net70),
    .B(net60));
 sg13g2_nand2_1 _613_ (.Y(_210_),
    .A(net63),
    .B(net68));
 sg13g2_nand2_1 _614_ (.Y(_211_),
    .A(net65),
    .B(net68));
 sg13g2_or2_1 _615_ (.X(_212_),
    .B(_211_),
    .A(_194_));
 sg13g2_xor2_1 _616_ (.B(_211_),
    .A(_194_),
    .X(_213_));
 sg13g2_nand2b_1 _617_ (.Y(_214_),
    .B(_213_),
    .A_N(_209_));
 sg13g2_xnor2_1 _618_ (.Y(_215_),
    .A(_209_),
    .B(_213_));
 sg13g2_nand2_1 _619_ (.Y(_216_),
    .A(_203_),
    .B(_215_));
 sg13g2_xor2_1 _620_ (.B(_215_),
    .A(_203_),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[2] ));
 sg13g2_nor2_1 _621_ (.A(_186_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[2] ),
    .Y(_217_));
 sg13g2_and2_1 _622_ (.A(net60),
    .B(net68),
    .X(_218_));
 sg13g2_xnor2_1 _623_ (.Y(_219_),
    .A(net60),
    .B(net68));
 sg13g2_a21oi_1 _624_ (.A1(_194_),
    .A2(_200_),
    .Y(_220_),
    .B1(_219_));
 sg13g2_nand3_1 _625_ (.B(_200_),
    .C(_219_),
    .A(_194_),
    .Y(_221_));
 sg13g2_nor2b_1 _626_ (.A(_220_),
    .B_N(_221_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[2] ));
 sg13g2_nor2_1 _627_ (.A(_199_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[2] ),
    .Y(_222_));
 sg13g2_a21oi_1 _628_ (.A1(net56),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[1] ),
    .Y(_223_),
    .B1(_196_));
 sg13g2_inv_1 _629_ (.Y(_224_),
    .A(_223_));
 sg13g2_xnor2_1 _630_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[2] ),
    .A(_219_),
    .B(_223_));
 sg13g2_o21ai_1 _631_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$valid ),
    .Y(_225_),
    .A1(_193_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[2] ));
 sg13g2_nor4_2 _632_ (.A(_208_),
    .B(_217_),
    .C(_222_),
    .Y(_226_),
    .D(_225_));
 sg13g2_nor2_1 _633_ (.A(net50),
    .B(net54),
    .Y(_227_));
 sg13g2_nor2_2 _634_ (.A(_226_),
    .B(_227_),
    .Y(_228_));
 sg13g2_inv_1 _635_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[2] ),
    .A(_228_));
 sg13g2_nand2_1 _636_ (.Y(_229_),
    .A(net70),
    .B(net58));
 sg13g2_and2_1 _637_ (.A(_212_),
    .B(_214_),
    .X(_230_));
 sg13g2_nand2_1 _638_ (.Y(_231_),
    .A(net60),
    .B(net69));
 sg13g2_or2_1 _639_ (.X(_232_),
    .B(_210_),
    .A(_085_));
 sg13g2_xnor2_1 _640_ (.Y(_233_),
    .A(_085_),
    .B(_210_));
 sg13g2_xor2_1 _641_ (.B(_233_),
    .A(_231_),
    .X(_234_));
 sg13g2_inv_1 _642_ (.Y(_235_),
    .A(_234_));
 sg13g2_xnor2_1 _643_ (.Y(_236_),
    .A(_230_),
    .B(_234_));
 sg13g2_nand2b_1 _644_ (.Y(_237_),
    .B(_236_),
    .A_N(_229_));
 sg13g2_xnor2_1 _645_ (.Y(_238_),
    .A(_229_),
    .B(_236_));
 sg13g2_nand2b_1 _646_ (.Y(_239_),
    .B(_238_),
    .A_N(_216_));
 sg13g2_xor2_1 _647_ (.B(_238_),
    .A(_216_),
    .X(_240_));
 sg13g2_inv_1 _648_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[3] ),
    .A(_240_));
 sg13g2_nand2b_1 _649_ (.Y(_241_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[3] ),
    .A_N(net58));
 sg13g2_xor2_1 _650_ (.B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[3] ),
    .A(net58),
    .X(_242_));
 sg13g2_nor2b_1 _651_ (.A(net60),
    .B_N(net68),
    .Y(_243_));
 sg13g2_a21oi_1 _652_ (.A1(_219_),
    .A2(_224_),
    .Y(_244_),
    .B1(_243_));
 sg13g2_xor2_1 _653_ (.B(_244_),
    .A(_242_),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[3] ));
 sg13g2_o21ai_1 _654_ (.B1(_242_),
    .Y(_245_),
    .A1(_218_),
    .A2(_220_));
 sg13g2_or3_1 _655_ (.A(_218_),
    .B(_220_),
    .C(_242_),
    .X(_246_));
 sg13g2_and2_1 _656_ (.A(_245_),
    .B(_246_),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[3] ));
 sg13g2_o21ai_1 _657_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$valid ),
    .Y(_247_),
    .A1(_199_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[3] ));
 sg13g2_inv_1 _658_ (.Y(_248_),
    .A(_247_));
 sg13g2_o21ai_1 _659_ (.B1(_248_),
    .Y(_249_),
    .A1(_193_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[3] ));
 sg13g2_a221oi_1 _660_ (.B2(_240_),
    .C1(_249_),
    .B1(_185_),
    .A1(_101_),
    .Y(_250_),
    .A2(_182_));
 sg13g2_nor2_1 _661_ (.A(net49),
    .B(net54),
    .Y(_251_));
 sg13g2_nor2_2 _662_ (.A(_250_),
    .B(_251_),
    .Y(_252_));
 sg13g2_inv_2 _663_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[3] ),
    .A(_252_));
 sg13g2_o21ai_1 _664_ (.B1(_237_),
    .Y(_253_),
    .A1(_230_),
    .A2(_235_));
 sg13g2_nand2_1 _665_ (.Y(_254_),
    .A(net58),
    .B(net69));
 sg13g2_o21ai_1 _666_ (.B1(_232_),
    .Y(_255_),
    .A1(_231_),
    .A2(_233_));
 sg13g2_nand2_1 _667_ (.Y(_256_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[4] ),
    .B(net64));
 sg13g2_nor2_1 _668_ (.A(_085_),
    .B(_256_),
    .Y(_257_));
 sg13g2_a22oi_1 _669_ (.Y(_258_),
    .B1(net63),
    .B2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[3] ),
    .A2(net66),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[4] ));
 sg13g2_nor2_1 _670_ (.A(_257_),
    .B(_258_),
    .Y(_259_));
 sg13g2_xor2_1 _671_ (.B(_259_),
    .A(_218_),
    .X(_260_));
 sg13g2_nand2_1 _672_ (.Y(_261_),
    .A(_255_),
    .B(_260_));
 sg13g2_xnor2_1 _673_ (.Y(_262_),
    .A(_255_),
    .B(_260_));
 sg13g2_xor2_1 _674_ (.B(_262_),
    .A(_254_),
    .X(_263_));
 sg13g2_nand2_1 _675_ (.Y(_264_),
    .A(_253_),
    .B(_263_));
 sg13g2_xnor2_1 _676_ (.Y(_265_),
    .A(_253_),
    .B(_263_));
 sg13g2_xor2_1 _677_ (.B(_265_),
    .A(_239_),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[4] ));
 sg13g2_o21ai_1 _678_ (.B1(_264_),
    .Y(_266_),
    .A1(_239_),
    .A2(_265_));
 sg13g2_o21ai_1 _679_ (.B1(_261_),
    .Y(_267_),
    .A1(_254_),
    .A2(_262_));
 sg13g2_nand2_1 _680_ (.Y(_268_),
    .A(net58),
    .B(net68));
 sg13g2_a21o_1 _681_ (.A2(_259_),
    .A1(_218_),
    .B1(_257_),
    .X(_269_));
 sg13g2_nand2_1 _682_ (.Y(_270_),
    .A(net60),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[3] ));
 sg13g2_nand2_2 _683_ (.Y(_271_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[5] ),
    .B(net67));
 sg13g2_xor2_1 _684_ (.B(_271_),
    .A(_256_),
    .X(_272_));
 sg13g2_nand2b_1 _685_ (.Y(_273_),
    .B(_272_),
    .A_N(_270_));
 sg13g2_xnor2_1 _686_ (.Y(_274_),
    .A(_270_),
    .B(_272_));
 sg13g2_nand2_1 _687_ (.Y(_275_),
    .A(_269_),
    .B(_274_));
 sg13g2_xnor2_1 _688_ (.Y(_276_),
    .A(_269_),
    .B(_274_));
 sg13g2_xor2_1 _689_ (.B(_276_),
    .A(_268_),
    .X(_277_));
 sg13g2_xnor2_1 _690_ (.Y(_278_),
    .A(_267_),
    .B(_277_));
 sg13g2_nor2b_1 _691_ (.A(_278_),
    .B_N(_266_),
    .Y(_279_));
 sg13g2_xnor2_1 _692_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[5] ),
    .A(_266_),
    .B(_278_));
 sg13g2_a21o_1 _693_ (.A2(_277_),
    .A1(_267_),
    .B1(_279_),
    .X(_280_));
 sg13g2_o21ai_1 _694_ (.B1(_275_),
    .Y(_281_),
    .A1(_268_),
    .A2(_276_));
 sg13g2_nand2_2 _695_ (.Y(_282_),
    .A(\FpgaPins_Fpga_CALC_val2_a1[3] ),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[3] ));
 sg13g2_o21ai_1 _696_ (.B1(_273_),
    .Y(_283_),
    .A1(_256_),
    .A2(_271_));
 sg13g2_nand2_1 _697_ (.Y(_284_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[4] ),
    .B(net61));
 sg13g2_nand2_1 _698_ (.Y(_285_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[6] ),
    .B(net64));
 sg13g2_nor2_1 _699_ (.A(_271_),
    .B(_285_),
    .Y(_286_));
 sg13g2_or2_1 _700_ (.X(_287_),
    .B(_285_),
    .A(_271_));
 sg13g2_a22oi_1 _701_ (.Y(_288_),
    .B1(net63),
    .B2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[5] ),
    .A2(net67),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[6] ));
 sg13g2_nor2_1 _702_ (.A(_286_),
    .B(_288_),
    .Y(_289_));
 sg13g2_xnor2_1 _703_ (.Y(_290_),
    .A(_284_),
    .B(_289_));
 sg13g2_nand2_1 _704_ (.Y(_291_),
    .A(_283_),
    .B(_290_));
 sg13g2_xnor2_1 _705_ (.Y(_292_),
    .A(_283_),
    .B(_290_));
 sg13g2_xor2_1 _706_ (.B(_292_),
    .A(_282_),
    .X(_293_));
 sg13g2_xnor2_1 _707_ (.Y(_294_),
    .A(_281_),
    .B(_293_));
 sg13g2_nor2b_1 _708_ (.A(_294_),
    .B_N(_280_),
    .Y(_295_));
 sg13g2_xnor2_1 _709_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[6] ),
    .A(_280_),
    .B(_294_));
 sg13g2_a21oi_1 _710_ (.A1(_281_),
    .A2(_293_),
    .Y(_296_),
    .B1(_295_));
 sg13g2_o21ai_1 _711_ (.B1(_291_),
    .Y(_297_),
    .A1(_282_),
    .A2(_292_));
 sg13g2_o21ai_1 _712_ (.B1(_287_),
    .Y(_298_),
    .A1(_284_),
    .A2(_288_));
 sg13g2_nand2_1 _713_ (.Y(_299_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[4] ),
    .B(net59));
 sg13g2_nand2_1 _714_ (.Y(_300_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[5] ),
    .B(net61));
 sg13g2_xnor2_1 _715_ (.Y(_301_),
    .A(_299_),
    .B(_300_));
 sg13g2_nand2_1 _716_ (.Y(_302_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[7] ),
    .B(net67));
 sg13g2_xor2_1 _717_ (.B(_302_),
    .A(_285_),
    .X(_303_));
 sg13g2_xnor2_1 _718_ (.Y(_304_),
    .A(_301_),
    .B(_303_));
 sg13g2_xnor2_1 _719_ (.Y(_305_),
    .A(_298_),
    .B(_304_));
 sg13g2_xnor2_1 _720_ (.Y(_306_),
    .A(_297_),
    .B(_305_));
 sg13g2_xnor2_1 _721_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[7] ),
    .A(_296_),
    .B(_306_));
 sg13g2_o21ai_1 _722_ (.B1(_241_),
    .Y(_307_),
    .A1(_242_),
    .A2(_244_));
 sg13g2_xnor2_1 _723_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[4] ),
    .A(_016_),
    .B(_307_));
 sg13g2_nor2_1 _724_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[4] ),
    .B(_307_),
    .Y(_308_));
 sg13g2_xnor2_1 _725_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[5] ),
    .A(_000_),
    .B(_308_));
 sg13g2_nor3_1 _726_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[5] ),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[4] ),
    .C(_307_),
    .Y(_309_));
 sg13g2_xnor2_1 _727_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[6] ),
    .A(_011_),
    .B(_309_));
 sg13g2_and2_1 _728_ (.A(_365_),
    .B(_309_),
    .X(_310_));
 sg13g2_xnor2_1 _729_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[7] ),
    .A(_009_),
    .B(_310_));
 sg13g2_nand2_1 _730_ (.Y(_311_),
    .A(_245_),
    .B(_282_));
 sg13g2_a21oi_1 _731_ (.A1(_245_),
    .A2(_282_),
    .Y(_312_),
    .B1(_367_));
 sg13g2_xnor2_1 _732_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[4] ),
    .A(_367_),
    .B(_311_));
 sg13g2_xnor2_1 _733_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[5] ),
    .A(_000_),
    .B(_312_));
 sg13g2_nand2_1 _734_ (.Y(_313_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[5] ),
    .B(_312_));
 sg13g2_nor2_1 _735_ (.A(_011_),
    .B(_313_),
    .Y(_314_));
 sg13g2_xor2_1 _736_ (.B(_313_),
    .A(_011_),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[6] ));
 sg13g2_xnor2_1 _737_ (.Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[7] ),
    .A(_009_),
    .B(_314_));
 sg13g2_o21ai_1 _738_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$valid ),
    .Y(_315_),
    .A1(_199_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[4] ));
 sg13g2_inv_1 _739_ (.Y(_316_),
    .A(_315_));
 sg13g2_o21ai_1 _740_ (.B1(_316_),
    .Y(_317_),
    .A1(_193_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[4] ));
 sg13g2_a21oi_1 _741_ (.A1(_074_),
    .A2(_182_),
    .Y(_318_),
    .B1(_317_));
 sg13g2_o21ai_1 _742_ (.B1(_318_),
    .Y(_319_),
    .A1(_186_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[4] ));
 sg13g2_o21ai_1 _743_ (.B1(_319_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[4] ),
    .A1(_001_),
    .A2(net55));
 sg13g2_nand2_1 _744_ (.Y(_320_),
    .A(_057_),
    .B(_182_));
 sg13g2_o21ai_1 _745_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$valid ),
    .Y(_321_),
    .A1(_199_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[5] ));
 sg13g2_o21ai_1 _746_ (.B1(_320_),
    .Y(_322_),
    .A1(_193_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[5] ));
 sg13g2_nor2_1 _747_ (.A(_321_),
    .B(_322_),
    .Y(_323_));
 sg13g2_o21ai_1 _748_ (.B1(_323_),
    .Y(_324_),
    .A1(_186_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[5] ));
 sg13g2_o21ai_1 _749_ (.B1(_324_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[5] ),
    .A1(_000_),
    .A2(net55));
 sg13g2_nor2_1 _750_ (.A(_186_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[6] ),
    .Y(_325_));
 sg13g2_nor2_1 _751_ (.A(_199_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[6] ),
    .Y(_326_));
 sg13g2_o21ai_1 _752_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$valid ),
    .Y(_327_),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$quot[6] ),
    .A2(_183_));
 sg13g2_nor2_1 _753_ (.A(_193_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[6] ),
    .Y(_328_));
 sg13g2_nor4_1 _754_ (.A(_325_),
    .B(_326_),
    .C(_327_),
    .D(_328_),
    .Y(_329_));
 sg13g2_inv_1 _755_ (.Y(_330_),
    .A(_329_));
 sg13g2_o21ai_1 _756_ (.B1(_330_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[6] ),
    .A1(_011_),
    .A2(net55));
 sg13g2_nor2_1 _757_ (.A(_199_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[7] ),
    .Y(_331_));
 sg13g2_a21oi_1 _758_ (.A1(_031_),
    .A2(_182_),
    .Y(_332_),
    .B1(_331_));
 sg13g2_o21ai_1 _759_ (.B1(_332_),
    .Y(_333_),
    .A1(_193_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$diff[7] ));
 sg13g2_nor3_1 _760_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$reset ),
    .B(_018_),
    .C(_333_),
    .Y(_334_));
 sg13g2_o21ai_1 _761_ (.B1(_334_),
    .Y(_335_),
    .A1(_186_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$prod[7] ));
 sg13g2_o21ai_1 _762_ (.B1(_335_),
    .Y(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[7] ),
    .A1(_009_),
    .A2(net55));
 sg13g2_a21oi_2 _763_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[1] ),
    .Y(_336_),
    .A2(_191_),
    .A1(_189_));
 sg13g2_nor2_2 _764_ (.A(_228_),
    .B(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[3] ),
    .Y(_337_));
 sg13g2_nor2_1 _765_ (.A(_228_),
    .B(_252_),
    .Y(_338_));
 sg13g2_nand2_1 _766_ (.Y(_339_),
    .A(_228_),
    .B(_252_));
 sg13g2_nor2b_1 _767_ (.A(_338_),
    .B_N(_339_),
    .Y(_340_));
 sg13g2_nand2_1 _768_ (.Y(_341_),
    .A(_336_),
    .B(_340_));
 sg13g2_o21ai_1 _769_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[1] ),
    .Y(_342_),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[2] ),
    .A2(_252_));
 sg13g2_o21ai_1 _770_ (.B1(_342_),
    .Y(_343_),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[0] ),
    .A2(_337_));
 sg13g2_nor2b_1 _771_ (.A(_343_),
    .B_N(_341_),
    .Y(\DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[0] ));
 sg13g2_nand2b_1 _772_ (.Y(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[0].@0$viz_lit ),
    .B(_341_),
    .A_N(_343_));
 sg13g2_nand2_2 _773_ (.Y(_344_),
    .A(_207_),
    .B(_252_));
 sg13g2_inv_1 _774_ (.Y(_345_),
    .A(_344_));
 sg13g2_a21oi_1 _775_ (.A1(_192_),
    .A2(_345_),
    .Y(_346_),
    .B1(_228_));
 sg13g2_o21ai_1 _776_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[2] ),
    .Y(_347_),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[0] ),
    .A2(_344_));
 sg13g2_a21oi_2 _777_ (.B1(_207_),
    .Y(_348_),
    .A2(_191_),
    .A1(_189_));
 sg13g2_and2_1 _778_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[3] ),
    .B(_348_),
    .X(_349_));
 sg13g2_nand2_1 _779_ (.Y(_350_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[3] ),
    .B(_348_));
 sg13g2_nand2_1 _780_ (.Y(_351_),
    .A(_337_),
    .B(_348_));
 sg13g2_and2_1 _781_ (.A(_336_),
    .B(_338_),
    .X(_352_));
 sg13g2_a22oi_1 _782_ (.Y(_353_),
    .B1(_348_),
    .B2(_337_),
    .A2(_338_),
    .A1(_336_));
 sg13g2_a221oi_1 _783_ (.B2(_347_),
    .C1(_352_),
    .B1(_350_),
    .A1(_337_),
    .Y(\DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[1] ),
    .A2(_348_));
 sg13g2_o21ai_1 _784_ (.B1(_353_),
    .Y(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[1].@0$viz_lit ),
    .A1(_346_),
    .A2(_349_));
 sg13g2_nand2_1 _785_ (.Y(_354_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[1] ),
    .B(_339_));
 sg13g2_inv_1 _786_ (.Y(_355_),
    .A(_354_));
 sg13g2_o21ai_1 _787_ (.B1(_344_),
    .Y(_356_),
    .A1(_192_),
    .A2(_355_));
 sg13g2_nor2_1 _788_ (.A(_340_),
    .B(_356_),
    .Y(\DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[2] ));
 sg13g2_or2_1 _789_ (.X(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[2].@0$viz_lit ),
    .B(_356_),
    .A(_340_));
 sg13g2_xnor2_1 _790_ (.Y(_357_),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[0] ),
    .B(_228_));
 sg13g2_mux2_1 _791_ (.A0(_355_),
    .A1(_345_),
    .S(_357_),
    .X(\DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[3] ));
 sg13g2_mux2_1 _792_ (.A0(_354_),
    .A1(_344_),
    .S(_357_),
    .X(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[3].@0$viz_lit ));
 sg13g2_a21o_1 _793_ (.A2(_228_),
    .A1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[0] ),
    .B1(_337_),
    .X(_358_));
 sg13g2_o21ai_1 _794_ (.B1(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[1] ),
    .Y(_359_),
    .A1(_192_),
    .A2(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[3] ));
 sg13g2_and2_1 _795_ (.A(_358_),
    .B(_359_),
    .X(\DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[4] ));
 sg13g2_nand2_1 _796_ (.Y(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[4].@0$viz_lit ),
    .A(_358_),
    .B(_359_));
 sg13g2_nor2_1 _797_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[2] ),
    .B(_344_),
    .Y(_360_));
 sg13g2_inv_1 _798_ (.Y(_361_),
    .A(_360_));
 sg13g2_nor2_1 _799_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[0] ),
    .B(_361_),
    .Y(_362_));
 sg13g2_a21oi_1 _800_ (.A1(_339_),
    .A2(_353_),
    .Y(\DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[5] ),
    .B1(_362_));
 sg13g2_a21o_1 _801_ (.A2(_353_),
    .A1(_339_),
    .B1(_362_),
    .X(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[5].@0$viz_lit ));
 sg13g2_nand3_1 _802_ (.B(_207_),
    .C(_338_),
    .A(_192_),
    .Y(_363_));
 sg13g2_and3_1 _803_ (.X(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[6].@0$viz_lit ),
    .A(_351_),
    .B(_361_),
    .C(_363_));
 sg13g2_nand3_1 _804_ (.B(_361_),
    .C(_363_),
    .A(_351_),
    .Y(\DEBUG_SIGS_GTKWAVE.@0$sseg_segment_n[6] ));
 sg13g2_o21ai_1 _805_ (.B1(_319_),
    .Y(_012_),
    .A1(_367_),
    .A2(net54));
 sg13g2_o21ai_1 _806_ (.B1(_324_),
    .Y(_013_),
    .A1(_366_),
    .A2(net54));
 sg13g2_o21ai_1 _807_ (.B1(_330_),
    .Y(_014_),
    .A1(_365_),
    .A2(net54));
 sg13g2_o21ai_1 _808_ (.B1(_335_),
    .Y(_015_),
    .A1(_364_),
    .A2(net54));
 sg13g2_xor2_1 _809_ (.B(net65),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[0] ),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$sum[0] ));
 sg13g2_dfrbp_1 _810_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net30),
    .D(_012_),
    .Q_N(_001_),
    .Q(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[4] ));
 sg13g2_dfrbp_1 _811_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net26),
    .D(_013_),
    .Q_N(_000_),
    .Q(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[5] ));
 sg13g2_dfrbp_1 _812_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net28),
    .D(_014_),
    .Q_N(_011_),
    .Q(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[6] ));
 sg13g2_dfrbp_1 _813_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net31),
    .D(net45),
    .Q_N(_009_),
    .Q(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[7] ));
 sg13g2_dfrbp_1 _814_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net32),
    .D(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[0] ),
    .Q_N(_008_),
    .Q(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[0] ));
 sg13g2_dfrbp_1 _815_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net33),
    .D(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[1] ),
    .Q_N(_007_),
    .Q(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[1] ));
 sg13g2_dfrbp_1 _816_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net34),
    .D(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[2] ),
    .Q_N(_006_),
    .Q(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[2] ));
 sg13g2_dfrbp_1 _817_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net35),
    .D(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[3] ),
    .Q_N(_005_),
    .Q(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[3] ));
 sg13g2_dfrbp_1 _818_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net36),
    .D(net2),
    .Q_N(_002_),
    .Q(\FpgaPins_Fpga_CALC_val2_a1[0] ));
 sg13g2_dfrbp_1 _819_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net37),
    .D(net3),
    .Q_N(_003_),
    .Q(\FpgaPins_Fpga_CALC_val2_a1[1] ));
 sg13g2_dfrbp_1 _820_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net38),
    .D(net4),
    .Q_N(_004_),
    .Q(\FpgaPins_Fpga_CALC_val2_a1[2] ));
 sg13g2_dfrbp_1 _821_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net39),
    .D(net5),
    .Q_N(_010_),
    .Q(\FpgaPins_Fpga_CALC_val2_a1[3] ));
 sg13g2_dfrbp_1 _822_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net40),
    .D(net6),
    .Q_N(_374_),
    .Q(\FpgaPins_Fpga_CALC_op_a1[0] ));
 sg13g2_dfrbp_1 _823_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net41),
    .D(net7),
    .Q_N(_375_),
    .Q(\FpgaPins_Fpga_CALC_op_a1[1] ));
 sg13g2_dfrbp_1 _824_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net27),
    .D(net42),
    .Q_N(_376_),
    .Q(FpgaPins_Fpga_CALC_equals_in_a2));
 sg13g2_dfrbp_1 _825_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net29),
    .D(net8),
    .Q_N(_373_),
    .Q(FpgaPins_Fpga_CALC_equals_in_a1));
 sg13g2_tiehi _824__27 (.L_HI(net27));
 sg13g2_tiehi _812__28 (.L_HI(net28));
 sg13g2_tiehi _825__29 (.L_HI(net29));
 sg13g2_tiehi _810__30 (.L_HI(net30));
 sg13g2_tiehi _813__31 (.L_HI(net31));
 sg13g2_tiehi _814__32 (.L_HI(net32));
 sg13g2_tiehi _815__33 (.L_HI(net33));
 sg13g2_tiehi _816__34 (.L_HI(net34));
 sg13g2_tiehi _817__35 (.L_HI(net35));
 sg13g2_tiehi _818__36 (.L_HI(net36));
 sg13g2_tiehi _819__37 (.L_HI(net37));
 sg13g2_tiehi _820__38 (.L_HI(net38));
 sg13g2_tiehi _821__39 (.L_HI(net39));
 sg13g2_tiehi _822__40 (.L_HI(net40));
 sg13g2_tiehi _823__41 (.L_HI(net41));
 sg13g2_dlygate4sd3_1 hold4 (.A(_015_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold3 (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[7] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold2 (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[6] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold1 (.A(FpgaPins_Fpga_CALC_equals_in_a1),
    .X(net42));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold9 (.A(_006_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold8 (.A(_005_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold7 (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[4] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold6 (.A(_007_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold5 (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[5] ),
    .X(net46));
 sg13g2_tielo tt_um_ezchips_calc_9 (.L_LO(net9));
 sg13g2_tielo tt_um_ezchips_calc_10 (.L_LO(net10));
 sg13g2_tielo tt_um_ezchips_calc_11 (.L_LO(net11));
 sg13g2_tielo tt_um_ezchips_calc_12 (.L_LO(net12));
 sg13g2_tielo tt_um_ezchips_calc_13 (.L_LO(net13));
 sg13g2_tielo tt_um_ezchips_calc_14 (.L_LO(net14));
 sg13g2_tielo tt_um_ezchips_calc_15 (.L_LO(net15));
 sg13g2_tielo tt_um_ezchips_calc_16 (.L_LO(net16));
 sg13g2_tielo tt_um_ezchips_calc_17 (.L_LO(net17));
 sg13g2_tielo tt_um_ezchips_calc_18 (.L_LO(net18));
 sg13g2_tielo tt_um_ezchips_calc_19 (.L_LO(net19));
 sg13g2_tielo tt_um_ezchips_calc_20 (.L_LO(net20));
 sg13g2_tielo tt_um_ezchips_calc_21 (.L_LO(net21));
 sg13g2_tielo tt_um_ezchips_calc_22 (.L_LO(net22));
 sg13g2_tielo tt_um_ezchips_calc_23 (.L_LO(net23));
 sg13g2_tielo tt_um_ezchips_calc_24 (.L_LO(net24));
 sg13g2_tielo tt_um_ezchips_calc_25 (.L_LO(net25));
 sg13g2_tiehi _811__26 (.L_HI(net26));
 sg13g2_buf_1 _873_ (.A(net2),
    .X(\DEBUG_SIGS_GTKWAVE.@0$slideswitch[0] ));
 sg13g2_buf_1 _874_ (.A(net3),
    .X(\DEBUG_SIGS_GTKWAVE.@0$slideswitch[1] ));
 sg13g2_buf_1 _875_ (.A(net4),
    .X(\DEBUG_SIGS_GTKWAVE.@0$slideswitch[2] ));
 sg13g2_buf_1 _876_ (.A(net5),
    .X(\DEBUG_SIGS_GTKWAVE.@0$slideswitch[3] ));
 sg13g2_buf_1 _877_ (.A(net6),
    .X(\DEBUG_SIGS_GTKWAVE.@0$slideswitch[4] ));
 sg13g2_buf_1 _878_ (.A(net7),
    .X(\DEBUG_SIGS_GTKWAVE.@0$slideswitch[5] ));
 sg13g2_buf_1 _879_ (.A(ui_in[6]),
    .X(\DEBUG_SIGS_GTKWAVE.@0$slideswitch[6] ));
 sg13g2_buf_1 _880_ (.A(net8),
    .X(\DEBUG_SIGS_GTKWAVE.@0$slideswitch[7] ));
 sg13g2_buf_1 _881_ (.A(net2),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$val2[0] ));
 sg13g2_buf_1 _882_ (.A(net3),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$val2[1] ));
 sg13g2_buf_1 _883_ (.A(net4),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$val2[2] ));
 sg13g2_buf_1 _884_ (.A(net5),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$val2[3] ));
 sg13g2_buf_1 _885_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[0] ),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[0] ));
 sg13g2_buf_1 _886_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[1] ),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[1] ));
 sg13g2_buf_1 _887_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[2] ),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[2] ));
 sg13g2_buf_1 _888_ (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$digit[3] ),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$out[3] ));
 sg13g2_buf_1 _889_ (.A(net6),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$op[0] ));
 sg13g2_buf_1 _890_ (.A(net7),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$op[1] ));
 sg13g2_buf_1 _891_ (.A(net8),
    .X(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@0$equals_in ));
 sg13g2_buf_1 _892_ (.A(net2),
    .X(\DEBUG_SIGS_GTKWAVE./switch[0].@0$viz_switch ));
 sg13g2_buf_1 _893_ (.A(net3),
    .X(\DEBUG_SIGS_GTKWAVE./switch[1].@0$viz_switch ));
 sg13g2_buf_1 _894_ (.A(net4),
    .X(\DEBUG_SIGS_GTKWAVE./switch[2].@0$viz_switch ));
 sg13g2_buf_1 _895_ (.A(net5),
    .X(\DEBUG_SIGS_GTKWAVE./switch[3].@0$viz_switch ));
 sg13g2_buf_1 _896_ (.A(net6),
    .X(\DEBUG_SIGS_GTKWAVE./switch[4].@0$viz_switch ));
 sg13g2_buf_1 _897_ (.A(net7),
    .X(\DEBUG_SIGS_GTKWAVE./switch[5].@0$viz_switch ));
 sg13g2_buf_1 _898_ (.A(ui_in[6]),
    .X(\DEBUG_SIGS_GTKWAVE./switch[6].@0$viz_switch ));
 sg13g2_buf_1 _899_ (.A(net8),
    .X(\DEBUG_SIGS_GTKWAVE./switch[7].@0$viz_switch ));
 sg13g2_buf_1 _900_ (.A(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[0].@0$viz_lit ),
    .X(uo_out[0]));
 sg13g2_buf_2 _901_ (.A(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[1].@0$viz_lit ),
    .X(uo_out[1]));
 sg13g2_buf_1 _902_ (.A(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[2].@0$viz_lit ),
    .X(uo_out[2]));
 sg13g2_buf_2 _903_ (.A(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[3].@0$viz_lit ),
    .X(uo_out[3]));
 sg13g2_buf_1 _904_ (.A(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[4].@0$viz_lit ),
    .X(uo_out[4]));
 sg13g2_buf_2 _905_ (.A(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[5].@0$viz_lit ),
    .X(uo_out[5]));
 sg13g2_buf_1 _906_ (.A(\DEBUG_SIGS_GTKWAVE./digit[0]./leds[6].@0$viz_lit ),
    .X(uo_out[6]));
 sg13g2_buf_2 fanout54 (.A(_190_),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(_190_),
    .X(net55));
 sg13g2_buf_4 fanout56 (.X(net56),
    .A(_370_));
 sg13g2_buf_4 fanout57 (.X(net57),
    .A(_010_));
 sg13g2_buf_4 fanout58 (.X(net58),
    .A(net59));
 sg13g2_buf_4 fanout59 (.X(net59),
    .A(\FpgaPins_Fpga_CALC_val2_a1[3] ));
 sg13g2_buf_2 fanout60 (.A(net62),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(net62),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(\FpgaPins_Fpga_CALC_val2_a1[2] ),
    .X(net62));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(\FpgaPins_Fpga_CALC_val2_a1[1] ));
 sg13g2_buf_2 fanout64 (.A(\FpgaPins_Fpga_CALC_val2_a1[1] ),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(net66),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(\FpgaPins_Fpga_CALC_val2_a1[0] ),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(\FpgaPins_Fpga_CALC_val2_a1[0] ),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[2] ),
    .X(net68));
 sg13g2_buf_4 fanout69 (.X(net69),
    .A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[1] ));
 sg13g2_buf_2 fanout70 (.A(\DEBUG_SIGS_GTKWAVE./fpga_pins./fpga.P_calc.@1$val1[0] ),
    .X(net70));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_4 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_233 ();
 sg13g2_decap_8 FILLER_22_240 ();
 sg13g2_decap_8 FILLER_22_247 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_261 ();
 sg13g2_decap_8 FILLER_22_268 ();
 sg13g2_decap_8 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_decap_8 FILLER_22_289 ();
 sg13g2_decap_8 FILLER_22_296 ();
 sg13g2_decap_8 FILLER_22_303 ();
 sg13g2_decap_8 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_decap_8 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_338 ();
 sg13g2_decap_8 FILLER_22_345 ();
 sg13g2_decap_8 FILLER_22_352 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_decap_4 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_decap_8 FILLER_23_243 ();
 sg13g2_fill_2 FILLER_23_250 ();
 sg13g2_fill_1 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_fill_2 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_282 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_decap_8 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_337 ();
 sg13g2_decap_8 FILLER_23_344 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_108 ();
 sg13g2_decap_4 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_116 ();
 sg13g2_fill_2 FILLER_24_122 ();
 sg13g2_decap_8 FILLER_24_128 ();
 sg13g2_decap_4 FILLER_24_135 ();
 sg13g2_fill_2 FILLER_24_139 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_decap_8 FILLER_24_152 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_166 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_206 ();
 sg13g2_decap_4 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_decap_4 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_decap_4 FILLER_24_271 ();
 sg13g2_decap_4 FILLER_24_299 ();
 sg13g2_decap_8 FILLER_24_324 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_88 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_188 ();
 sg13g2_fill_2 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_216 ();
 sg13g2_fill_2 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_fill_2 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_decap_8 FILLER_25_286 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_318 ();
 sg13g2_decap_4 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_79 ();
 sg13g2_decap_4 FILLER_26_93 ();
 sg13g2_decap_4 FILLER_26_102 ();
 sg13g2_decap_4 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_138 ();
 sg13g2_decap_4 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_153 ();
 sg13g2_fill_2 FILLER_26_160 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_fill_2 FILLER_26_168 ();
 sg13g2_fill_1 FILLER_26_170 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_4 FILLER_26_182 ();
 sg13g2_fill_2 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_201 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_245 ();
 sg13g2_fill_1 FILLER_26_247 ();
 sg13g2_decap_4 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_275 ();
 sg13g2_fill_2 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_decap_4 FILLER_26_330 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_4 FILLER_27_70 ();
 sg13g2_fill_2 FILLER_27_100 ();
 sg13g2_fill_2 FILLER_27_106 ();
 sg13g2_fill_2 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_125 ();
 sg13g2_fill_2 FILLER_27_154 ();
 sg13g2_decap_4 FILLER_27_165 ();
 sg13g2_fill_1 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_202 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_fill_1 FILLER_27_234 ();
 sg13g2_decap_8 FILLER_27_243 ();
 sg13g2_decap_8 FILLER_27_250 ();
 sg13g2_decap_8 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_268 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_292 ();
 sg13g2_decap_4 FILLER_27_299 ();
 sg13g2_fill_1 FILLER_27_332 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_fill_1 FILLER_27_348 ();
 sg13g2_fill_2 FILLER_27_363 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_fill_2 FILLER_28_84 ();
 sg13g2_fill_1 FILLER_28_86 ();
 sg13g2_decap_8 FILLER_28_97 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_fill_2 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_fill_2 FILLER_28_159 ();
 sg13g2_decap_4 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_207 ();
 sg13g2_decap_4 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_228 ();
 sg13g2_decap_4 FILLER_28_237 ();
 sg13g2_decap_4 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_257 ();
 sg13g2_decap_4 FILLER_28_290 ();
 sg13g2_decap_4 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_4 FILLER_28_342 ();
 sg13g2_fill_2 FILLER_28_353 ();
 sg13g2_decap_4 FILLER_28_363 ();
 sg13g2_fill_2 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_99 ();
 sg13g2_fill_1 FILLER_29_101 ();
 sg13g2_decap_8 FILLER_29_120 ();
 sg13g2_decap_8 FILLER_29_127 ();
 sg13g2_decap_8 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_175 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_1 FILLER_29_205 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_fill_2 FILLER_29_260 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_decap_4 FILLER_29_298 ();
 sg13g2_fill_1 FILLER_29_302 ();
 sg13g2_fill_2 FILLER_29_325 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_fill_2 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_107 ();
 sg13g2_fill_2 FILLER_30_111 ();
 sg13g2_fill_1 FILLER_30_113 ();
 sg13g2_decap_8 FILLER_30_118 ();
 sg13g2_fill_2 FILLER_30_125 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_fill_2 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_decap_8 FILLER_30_195 ();
 sg13g2_fill_1 FILLER_30_219 ();
 sg13g2_decap_8 FILLER_30_255 ();
 sg13g2_decap_4 FILLER_30_262 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_282 ();
 sg13g2_decap_4 FILLER_30_287 ();
 sg13g2_decap_4 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_316 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_2 FILLER_30_324 ();
 sg13g2_decap_4 FILLER_30_330 ();
 sg13g2_fill_2 FILLER_30_334 ();
 sg13g2_fill_2 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_361 ();
 sg13g2_fill_1 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_fill_2 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_199 ();
 sg13g2_fill_2 FILLER_31_204 ();
 sg13g2_decap_4 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_223 ();
 sg13g2_decap_4 FILLER_31_230 ();
 sg13g2_fill_2 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_257 ();
 sg13g2_fill_2 FILLER_31_283 ();
 sg13g2_fill_2 FILLER_31_302 ();
 sg13g2_fill_1 FILLER_31_304 ();
 sg13g2_decap_4 FILLER_31_353 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_372 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_fill_2 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_118 ();
 sg13g2_decap_4 FILLER_32_125 ();
 sg13g2_fill_2 FILLER_32_129 ();
 sg13g2_decap_8 FILLER_32_135 ();
 sg13g2_decap_8 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_decap_4 FILLER_32_200 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_fill_2 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_2 FILLER_32_282 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_309 ();
 sg13g2_decap_4 FILLER_32_320 ();
 sg13g2_fill_2 FILLER_32_324 ();
 sg13g2_decap_8 FILLER_32_330 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_decap_4 FILLER_32_342 ();
 sg13g2_fill_2 FILLER_32_346 ();
 sg13g2_fill_2 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_4 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_109 ();
 sg13g2_fill_2 FILLER_33_118 ();
 sg13g2_decap_4 FILLER_33_146 ();
 sg13g2_fill_2 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_174 ();
 sg13g2_decap_8 FILLER_33_190 ();
 sg13g2_decap_8 FILLER_33_197 ();
 sg13g2_decap_8 FILLER_33_204 ();
 sg13g2_fill_2 FILLER_33_211 ();
 sg13g2_decap_4 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_247 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_decap_4 FILLER_33_294 ();
 sg13g2_fill_1 FILLER_33_298 ();
 sg13g2_decap_4 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_352 ();
 sg13g2_fill_2 FILLER_33_373 ();
 sg13g2_fill_1 FILLER_33_375 ();
 sg13g2_decap_4 FILLER_33_381 ();
 sg13g2_fill_1 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_4 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_130 ();
 sg13g2_decap_8 FILLER_34_135 ();
 sg13g2_decap_8 FILLER_34_142 ();
 sg13g2_fill_2 FILLER_34_149 ();
 sg13g2_fill_1 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_169 ();
 sg13g2_decap_8 FILLER_34_200 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_decap_4 FILLER_34_231 ();
 sg13g2_fill_2 FILLER_34_235 ();
 sg13g2_decap_8 FILLER_34_240 ();
 sg13g2_decap_4 FILLER_34_247 ();
 sg13g2_fill_2 FILLER_34_251 ();
 sg13g2_decap_8 FILLER_34_261 ();
 sg13g2_decap_8 FILLER_34_268 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_decap_4 FILLER_34_301 ();
 sg13g2_decap_4 FILLER_34_313 ();
 sg13g2_fill_2 FILLER_34_317 ();
 sg13g2_decap_4 FILLER_34_341 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_174 ();
 sg13g2_fill_2 FILLER_35_206 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_fill_1 FILLER_35_217 ();
 sg13g2_decap_4 FILLER_35_224 ();
 sg13g2_fill_1 FILLER_35_228 ();
 sg13g2_decap_4 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_decap_8 FILLER_35_275 ();
 sg13g2_decap_4 FILLER_35_282 ();
 sg13g2_decap_4 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_1 FILLER_35_320 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_fill_2 FILLER_35_372 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_138 ();
 sg13g2_decap_8 FILLER_36_145 ();
 sg13g2_decap_4 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_171 ();
 sg13g2_decap_4 FILLER_36_177 ();
 sg13g2_fill_2 FILLER_36_181 ();
 sg13g2_fill_1 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_226 ();
 sg13g2_decap_8 FILLER_36_233 ();
 sg13g2_fill_2 FILLER_36_240 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_2 FILLER_36_248 ();
 sg13g2_decap_8 FILLER_36_267 ();
 sg13g2_fill_2 FILLER_36_274 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_fill_2 FILLER_36_317 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_4 FILLER_36_362 ();
 sg13g2_fill_2 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_4 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_121 ();
 sg13g2_fill_2 FILLER_37_156 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_fill_1 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_183 ();
 sg13g2_fill_1 FILLER_37_190 ();
 sg13g2_fill_1 FILLER_37_264 ();
 sg13g2_decap_4 FILLER_37_269 ();
 sg13g2_fill_2 FILLER_37_273 ();
 sg13g2_decap_4 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_283 ();
 sg13g2_decap_8 FILLER_37_289 ();
 sg13g2_fill_1 FILLER_37_296 ();
 sg13g2_fill_2 FILLER_37_316 ();
 sg13g2_fill_1 FILLER_37_318 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_4 FILLER_37_333 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_decap_8 FILLER_38_188 ();
 sg13g2_fill_1 FILLER_38_195 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_4 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_255 ();
 sg13g2_decap_8 FILLER_38_295 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_320 ();
 sg13g2_fill_2 FILLER_38_394 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
 assign uo_out[7] = net25;
endmodule
